

module b17_C_2inp_gates_syn ( P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, 
        DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, 
        DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, 
        DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, 
        DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, 
        DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, 
        READY1, READY2, P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN, 
        P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN, 
        P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN, 
        P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN, 
        P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN, 
        P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN, 
        P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN, 
        P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN, 
        P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN, 
        P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN, 
        P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN, 
        P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN, 
        P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN, 
        P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN, 
        P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN, 
        P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN, 
        P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN, 
        P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, 
        P1_REIP_REG_6__SCAN_IN, P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, 
        P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, 
        P1_REIP_REG_0__SCAN_IN, P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, 
        P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, 
        P1_EBX_REG_26__SCAN_IN, P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, 
        P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, 
        P1_EBX_REG_20__SCAN_IN, P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, 
        P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, 
        P1_EBX_REG_14__SCAN_IN, P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, 
        P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, 
        P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, 
        P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, 
        P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, 
        P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, 
        P1_EAX_REG_28__SCAN_IN, P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, 
        P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, 
        P1_EAX_REG_22__SCAN_IN, P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, 
        P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, 
        P1_EAX_REG_16__SCAN_IN, P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, 
        P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, 
        P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, 
        P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, 
        P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, 
        P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, U355, 
        U356, U357, U358, U359, U360, U361, U362, U363, U364, U366, U367, U368, 
        U369, U370, U371, U372, U373, U374, U375, U347, U348, U349, U350, U351, 
        U352, U353, U354, U365, U376, U247, U246, U245, U244, U243, U242, U241, 
        U240, U239, U238, U237, U236, U235, U234, U233, U232, U231, U230, U229, 
        U228, U227, U226, U225, U224, U223, U222, U221, U220, U219, U218, U217, 
        U216, U251, U252, U253, U254, U255, U256, U257, U258, U259, U260, U261, 
        U262, U263, U264, U265, U266, U267, U268, U269, U270, U271, U272, U273, 
        U274, U275, U276, U277, U278, U279, U280, U281, U282, U212, U215, U213, 
        U214, P3_U3274, P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, 
        P3_U3059, P3_U3058, P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, 
        P3_U3052, P3_U3051, P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, 
        P3_U3045, P3_U3044, P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, 
        P3_U3038, P3_U3037, P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, 
        P3_U3031, P3_U3030, P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, 
        P3_U3026, P3_U3025, P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, 
        P3_U3019, P3_U3018, P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, 
        P3_U3012, P3_U3011, P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, 
        P3_U3005, P3_U3004, P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, 
        P3_U3282, P3_U2998, P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, 
        P3_U2992, P3_U2991, P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, 
        P3_U2985, P3_U2984, P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, 
        P3_U2978, P3_U2977, P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, 
        P3_U2971, P3_U2970, P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, 
        P3_U2964, P3_U2963, P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, 
        P3_U2957, P3_U2956, P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, 
        P3_U2950, P3_U2949, P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, 
        P3_U2943, P3_U2942, P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, 
        P3_U2936, P3_U2935, P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, 
        P3_U2929, P3_U2928, P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, 
        P3_U2922, P3_U2921, P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, 
        P3_U2915, P3_U2914, P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, 
        P3_U2908, P3_U2907, P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, 
        P3_U2901, P3_U2900, P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, 
        P3_U2894, P3_U2893, P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, 
        P3_U2887, P3_U2886, P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, 
        P3_U2880, P3_U2879, P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, 
        P3_U2873, P3_U2872, P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, 
        P3_U3285, P3_U3288, P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, 
        P3_U2864, P3_U2863, P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, 
        P3_U2857, P3_U2856, P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, 
        P3_U2850, P3_U2849, P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, 
        P3_U2843, P3_U2842, P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, 
        P3_U2836, P3_U2835, P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, 
        P3_U2829, P3_U2828, P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, 
        P3_U2822, P3_U2821, P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, 
        P3_U2815, P3_U2814, P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, 
        P3_U2808, P3_U2807, P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, 
        P3_U2801, P3_U2800, P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, 
        P3_U2794, P3_U2793, P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, 
        P3_U2787, P3_U2786, P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, 
        P3_U2780, P3_U2779, P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, 
        P3_U2773, P3_U2772, P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, 
        P3_U2766, P3_U2765, P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, 
        P3_U2759, P3_U2758, P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, 
        P3_U2752, P3_U2751, P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, 
        P3_U2745, P3_U2744, P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, 
        P3_U2738, P3_U2737, P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, 
        P3_U2731, P3_U2730, P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, 
        P3_U2724, P3_U2723, P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, 
        P3_U2717, P3_U2716, P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, 
        P3_U2710, P3_U2709, P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, 
        P3_U2703, P3_U2702, P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, 
        P3_U2696, P3_U2695, P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, 
        P3_U2689, P3_U2688, P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, 
        P3_U2682, P3_U2681, P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, 
        P3_U2675, P3_U2674, P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, 
        P3_U2668, P3_U2667, P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, 
        P3_U2661, P3_U2660, P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, 
        P3_U2654, P3_U2653, P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, 
        P3_U2647, P3_U2646, P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, 
        P3_U2640, P3_U2639, P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, 
        P3_U3295, P3_U2636, P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, 
        P3_U3298, P3_U3299, P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, 
        P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, 
        P2_U3179, P2_U3593, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, 
        P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, 
        P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, 
        P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, 
        P2_U3152, P2_U3151, P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, 
        P2_U3145, P2_U3144, P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, 
        P2_U3138, P2_U3137, P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, 
        P2_U3131, P2_U3130, P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, 
        P2_U3124, P2_U3123, P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, 
        P2_U3117, P2_U3116, P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, 
        P2_U3110, P2_U3109, P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, 
        P2_U3103, P2_U3102, P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, 
        P2_U3096, P2_U3095, P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, 
        P2_U3089, P2_U3088, P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, 
        P2_U3082, P2_U3081, P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, 
        P2_U3075, P2_U3074, P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, 
        P2_U3068, P2_U3067, P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, 
        P2_U3061, P2_U3060, P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, 
        P2_U3054, P2_U3053, P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, 
        P2_U3595, P2_U3596, P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, 
        P2_U3603, P2_U3604, P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, 
        P2_U3042, P2_U3041, P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, 
        P2_U3035, P2_U3034, P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, 
        P2_U3028, P2_U3027, P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, 
        P2_U3021, P2_U3020, P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, 
        P2_U3014, P2_U3013, P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, 
        P2_U3007, P2_U3006, P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, 
        P2_U3000, P2_U2999, P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, 
        P2_U2993, P2_U2992, P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, 
        P2_U2986, P2_U2985, P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, 
        P2_U2979, P2_U2978, P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, 
        P2_U2972, P2_U2971, P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, 
        P2_U2965, P2_U2964, P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, 
        P2_U2958, P2_U2957, P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, 
        P2_U2951, P2_U2950, P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, 
        P2_U2944, P2_U2943, P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, 
        P2_U2937, P2_U2936, P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, 
        P2_U2930, P2_U2929, P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, 
        P2_U2923, P2_U2922, P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, 
        P2_U2916, P2_U2915, P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, 
        P2_U2909, P2_U2908, P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, 
        P2_U2902, P2_U2901, P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, 
        P2_U2895, P2_U2894, P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, 
        P2_U2888, P2_U2887, P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, 
        P2_U2881, P2_U2880, P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, 
        P2_U2874, P2_U2873, P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, 
        P2_U2867, P2_U2866, P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, 
        P2_U2860, P2_U2859, P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, 
        P2_U2853, P2_U2852, P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, 
        P2_U2846, P2_U2845, P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, 
        P2_U2839, P2_U2838, P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, 
        P2_U2832, P2_U2831, P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, 
        P2_U2825, P2_U2824, P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, 
        P2_U2819, P2_U3609, P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, 
        P2_U2815, P2_U3612, P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, 
        P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, 
        P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, 
        P1_U3212, P1_U3211, P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, 
        P1_U3205, P1_U3204, P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, 
        P1_U3198, P1_U3197, P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, 
        P1_U3193, P1_U3192, P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, 
        P1_U3186, P1_U3185, P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, 
        P1_U3179, P1_U3178, P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, 
        P1_U3172, P1_U3171, P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, 
        P1_U3165, P1_U3164, P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, 
        P1_U3159, P1_U3158, P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, 
        P1_U3152, P1_U3151, P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, 
        P1_U3145, P1_U3144, P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, 
        P1_U3138, P1_U3137, P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, 
        P1_U3131, P1_U3130, P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, 
        P1_U3124, P1_U3123, P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, 
        P1_U3117, P1_U3116, P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, 
        P1_U3110, P1_U3109, P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, 
        P1_U3103, P1_U3102, P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, 
        P1_U3096, P1_U3095, P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, 
        P1_U3089, P1_U3088, P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, 
        P1_U3082, P1_U3081, P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, 
        P1_U3075, P1_U3074, P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, 
        P1_U3068, P1_U3067, P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, 
        P1_U3061, P1_U3060, P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, 
        P1_U3054, P1_U3053, P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, 
        P1_U3047, P1_U3046, P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, 
        P1_U3040, P1_U3039, P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, 
        P1_U3033, P1_U3468, P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, 
        P1_U3475, P1_U3476, P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, 
        P1_U3028, P1_U3027, P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, 
        P1_U3021, P1_U3020, P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, 
        P1_U3014, P1_U3013, P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, 
        P1_U3007, P1_U3006, P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, 
        P1_U3000, P1_U2999, P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, 
        P1_U2993, P1_U2992, P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, 
        P1_U2986, P1_U2985, P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, 
        P1_U2979, P1_U2978, P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, 
        P1_U2972, P1_U2971, P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, 
        P1_U2965, P1_U2964, P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, 
        P1_U2958, P1_U2957, P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, 
        P1_U2951, P1_U2950, P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, 
        P1_U2944, P1_U2943, P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, 
        P1_U2937, P1_U2936, P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, 
        P1_U2930, P1_U2929, P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, 
        P1_U2923, P1_U2922, P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, 
        P1_U2916, P1_U2915, P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, 
        P1_U2909, P1_U2908, P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, 
        P1_U2902, P1_U2901, P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, 
        P1_U2895, P1_U2894, P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, 
        P1_U2888, P1_U2887, P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, 
        P1_U2881, P1_U2880, P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, 
        P1_U2874, P1_U2873, P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, 
        P1_U2867, P1_U2866, P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, 
        P1_U2860, P1_U2859, P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, 
        P1_U2853, P1_U2852, P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, 
        P1_U2846, P1_U2845, P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, 
        P1_U2839, P1_U2838, P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, 
        P1_U2832, P1_U2831, P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, 
        P1_U2825, P1_U2824, P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, 
        P1_U2818, P1_U2817, P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, 
        P1_U2811, P1_U2810, P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, 
        P1_U3483, P1_U2806, P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, 
        P1_U2803, P1_U2802, P1_U3487, P1_U2801, keyinput127, keyinput126, 
        keyinput125, keyinput124, keyinput123, keyinput122, keyinput121, 
        keyinput120, keyinput119, keyinput118, keyinput117, keyinput116, 
        keyinput115, keyinput114, keyinput113, keyinput112, keyinput111, 
        keyinput110, keyinput109, keyinput108, keyinput107, keyinput106, 
        keyinput105, keyinput104, keyinput103, keyinput102, keyinput101, 
        keyinput100, keyinput99, keyinput98, keyinput97, keyinput96, 
        keyinput95, keyinput94, keyinput93, keyinput92, keyinput91, keyinput90, 
        keyinput89, keyinput88, keyinput87, keyinput86, keyinput85, keyinput84, 
        keyinput83, keyinput82, keyinput81, keyinput80, keyinput79, keyinput78, 
        keyinput77, keyinput76, keyinput75, keyinput74, keyinput73, keyinput72, 
        keyinput71, keyinput70, keyinput69, keyinput68, keyinput67, keyinput66, 
        keyinput65, keyinput64, keyinput63, keyinput62, keyinput61, keyinput60, 
        keyinput59, keyinput58, keyinput57, keyinput56, keyinput55, keyinput54, 
        keyinput53, keyinput52, keyinput51, keyinput50, keyinput49, keyinput48, 
        keyinput47, keyinput46, keyinput45, keyinput44, keyinput43, keyinput42, 
        keyinput41, keyinput40, keyinput39, keyinput38, keyinput37, keyinput36, 
        keyinput35, keyinput34, keyinput33, keyinput32, keyinput31, keyinput30, 
        keyinput29, keyinput28, keyinput27, keyinput26, keyinput25, keyinput24, 
        keyinput23, keyinput22, keyinput21, keyinput20, keyinput19, keyinput18, 
        keyinput17, keyinput16, keyinput15, keyinput14, keyinput13, keyinput12, 
        keyinput11, keyinput10, keyinput9, keyinput8, keyinput7, keyinput6, 
        keyinput5, keyinput4, keyinput3, keyinput2, keyinput1, keyinput0 );
  input P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_,
         DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_,
         DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_,
         DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_,
         DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_,
         DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2,
         P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN, keyinput127, keyinput126, keyinput125,
         keyinput124, keyinput123, keyinput122, keyinput121, keyinput120,
         keyinput119, keyinput118, keyinput117, keyinput116, keyinput115,
         keyinput114, keyinput113, keyinput112, keyinput111, keyinput110,
         keyinput109, keyinput108, keyinput107, keyinput106, keyinput105,
         keyinput104, keyinput103, keyinput102, keyinput101, keyinput100,
         keyinput99, keyinput98, keyinput97, keyinput96, keyinput95,
         keyinput94, keyinput93, keyinput92, keyinput91, keyinput90,
         keyinput89, keyinput88, keyinput87, keyinput86, keyinput85,
         keyinput84, keyinput83, keyinput82, keyinput81, keyinput80,
         keyinput79, keyinput78, keyinput77, keyinput76, keyinput75,
         keyinput74, keyinput73, keyinput72, keyinput71, keyinput70,
         keyinput69, keyinput68, keyinput67, keyinput66, keyinput65,
         keyinput64, keyinput63, keyinput62, keyinput61, keyinput60,
         keyinput59, keyinput58, keyinput57, keyinput56, keyinput55,
         keyinput54, keyinput53, keyinput52, keyinput51, keyinput50,
         keyinput49, keyinput48, keyinput47, keyinput46, keyinput45,
         keyinput44, keyinput43, keyinput42, keyinput41, keyinput40,
         keyinput39, keyinput38, keyinput37, keyinput36, keyinput35,
         keyinput34, keyinput33, keyinput32, keyinput31, keyinput30,
         keyinput29, keyinput28, keyinput27, keyinput26, keyinput25,
         keyinput24, keyinput23, keyinput22, keyinput21, keyinput20,
         keyinput19, keyinput18, keyinput17, keyinput16, keyinput15,
         keyinput14, keyinput13, keyinput12, keyinput11, keyinput10, keyinput9,
         keyinput8, keyinput7, keyinput6, keyinput5, keyinput4, keyinput3,
         keyinput2, keyinput1, keyinput0;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n9719, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9729, n9730,
         n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740,
         n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750,
         n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760,
         n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770,
         n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780,
         n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790,
         n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800,
         n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810,
         n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820,
         n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830,
         n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840,
         n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850,
         n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860,
         n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870,
         n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880,
         n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890,
         n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900,
         n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910,
         n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920,
         n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930,
         n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940,
         n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950,
         n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960,
         n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970,
         n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980,
         n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990,
         n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
         n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
         n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296,
         n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304,
         n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
         n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320,
         n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328,
         n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336,
         n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344,
         n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352,
         n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360,
         n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368,
         n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376,
         n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384,
         n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392,
         n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400,
         n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408,
         n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416,
         n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424,
         n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432,
         n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440,
         n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448,
         n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456,
         n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464,
         n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472,
         n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480,
         n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488,
         n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496,
         n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504,
         n10505, n10507, n10508, n10509, n10510, n10511, n10512, n10513,
         n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521,
         n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529,
         n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537,
         n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545,
         n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553,
         n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561,
         n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569,
         n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577,
         n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585,
         n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593,
         n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601,
         n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609,
         n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617,
         n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625,
         n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633,
         n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641,
         n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649,
         n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657,
         n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665,
         n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673,
         n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681,
         n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689,
         n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697,
         n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705,
         n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713,
         n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721,
         n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729,
         n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737,
         n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745,
         n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753,
         n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761,
         n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769,
         n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777,
         n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785,
         n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793,
         n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801,
         n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809,
         n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817,
         n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825,
         n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833,
         n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841,
         n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849,
         n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857,
         n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865,
         n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873,
         n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881,
         n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889,
         n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897,
         n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905,
         n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913,
         n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921,
         n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929,
         n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937,
         n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945,
         n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953,
         n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961,
         n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969,
         n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977,
         n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985,
         n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993,
         n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001,
         n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009,
         n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017,
         n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025,
         n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033,
         n11034, n11035, n11036, n11037, n11039, n11040, n11041, n11042,
         n11043, n11044, n11045, n11046, n11047, n11048, n11049, n11050,
         n11051, n11052, n11053, n11054, n11055, n11056, n11057, n11058,
         n11059, n11060, n11061, n11062, n11063, n11064, n11065, n11066,
         n11067, n11068, n11069, n11070, n11071, n11072, n11073, n11074,
         n11075, n11076, n11077, n11078, n11079, n11080, n11081, n11082,
         n11083, n11084, n11085, n11086, n11087, n11088, n11089, n11090,
         n11091, n11092, n11093, n11094, n11095, n11096, n11097, n11098,
         n11099, n11100, n11101, n11102, n11103, n11104, n11105, n11106,
         n11107, n11108, n11109, n11110, n11111, n11112, n11113, n11114,
         n11115, n11116, n11117, n11118, n11119, n11120, n11121, n11122,
         n11123, n11124, n11125, n11126, n11127, n11128, n11129, n11130,
         n11131, n11132, n11133, n11134, n11135, n11136, n11137, n11138,
         n11139, n11140, n11141, n11142, n11143, n11144, n11145, n11146,
         n11147, n11148, n11149, n11150, n11151, n11152, n11153, n11154,
         n11155, n11156, n11157, n11158, n11159, n11160, n11161, n11162,
         n11163, n11164, n11165, n11166, n11167, n11168, n11169, n11170,
         n11171, n11172, n11173, n11174, n11175, n11176, n11177, n11178,
         n11179, n11180, n11181, n11182, n11183, n11184, n11185, n11186,
         n11187, n11188, n11189, n11190, n11191, n11192, n11193, n11194,
         n11195, n11196, n11197, n11198, n11199, n11200, n11201, n11202,
         n11203, n11204, n11205, n11206, n11207, n11208, n11209, n11210,
         n11211, n11212, n11213, n11214, n11215, n11216, n11217, n11218,
         n11219, n11220, n11221, n11222, n11223, n11224, n11225, n11226,
         n11227, n11228, n11229, n11230, n11231, n11232, n11233, n11234,
         n11235, n11236, n11237, n11238, n11239, n11240, n11241, n11242,
         n11243, n11244, n11245, n11246, n11247, n11248, n11249, n11250,
         n11251, n11252, n11253, n11254, n11255, n11256, n11257, n11258,
         n11259, n11260, n11261, n11262, n11263, n11264, n11265, n11266,
         n11267, n11268, n11269, n11270, n11271, n11272, n11273, n11274,
         n11275, n11276, n11277, n11278, n11279, n11280, n11281, n11282,
         n11283, n11284, n11285, n11286, n11287, n11288, n11289, n11290,
         n11291, n11292, n11293, n11294, n11295, n11296, n11297, n11298,
         n11299, n11300, n11301, n11302, n11303, n11304, n11305, n11306,
         n11307, n11308, n11309, n11310, n11311, n11312, n11313, n11314,
         n11315, n11316, n11317, n11318, n11319, n11320, n11321, n11322,
         n11323, n11324, n11325, n11326, n11327, n11328, n11329, n11330,
         n11331, n11332, n11333, n11334, n11335, n11336, n11337, n11338,
         n11339, n11340, n11341, n11342, n11343, n11344, n11345, n11346,
         n11347, n11348, n11349, n11350, n11351, n11352, n11353, n11354,
         n11355, n11356, n11357, n11358, n11359, n11360, n11361, n11362,
         n11363, n11364, n11365, n11366, n11367, n11368, n11369, n11370,
         n11371, n11372, n11373, n11374, n11375, n11376, n11377, n11378,
         n11379, n11380, n11381, n11382, n11383, n11384, n11385, n11386,
         n11387, n11388, n11389, n11390, n11391, n11392, n11393, n11394,
         n11395, n11396, n11397, n11398, n11399, n11400, n11401, n11402,
         n11403, n11404, n11405, n11406, n11407, n11408, n11409, n11410,
         n11411, n11412, n11413, n11414, n11415, n11416, n11417, n11418,
         n11419, n11420, n11421, n11422, n11423, n11424, n11425, n11426,
         n11427, n11428, n11429, n11430, n11431, n11432, n11433, n11434,
         n11435, n11436, n11437, n11438, n11439, n11440, n11441, n11442,
         n11443, n11444, n11445, n11446, n11447, n11448, n11449, n11450,
         n11451, n11452, n11453, n11454, n11455, n11456, n11457, n11458,
         n11459, n11460, n11461, n11462, n11463, n11464, n11465, n11466,
         n11467, n11468, n11469, n11470, n11471, n11472, n11473, n11474,
         n11475, n11476, n11477, n11478, n11479, n11480, n11481, n11482,
         n11483, n11484, n11485, n11486, n11487, n11488, n11489, n11490,
         n11491, n11492, n11493, n11494, n11495, n11496, n11497, n11498,
         n11499, n11500, n11501, n11502, n11503, n11504, n11505, n11506,
         n11507, n11508, n11509, n11510, n11511, n11512, n11513, n11514,
         n11515, n11516, n11517, n11518, n11519, n11520, n11521, n11522,
         n11523, n11524, n11525, n11526, n11527, n11528, n11529, n11530,
         n11531, n11532, n11533, n11534, n11535, n11536, n11537, n11538,
         n11539, n11540, n11541, n11542, n11543, n11544, n11545, n11546,
         n11547, n11548, n11549, n11550, n11551, n11552, n11553, n11554,
         n11555, n11556, n11557, n11558, n11559, n11560, n11561, n11562,
         n11563, n11564, n11565, n11566, n11567, n11568, n11569, n11570,
         n11571, n11572, n11573, n11574, n11575, n11576, n11577, n11578,
         n11579, n11580, n11581, n11582, n11583, n11584, n11585, n11586,
         n11587, n11588, n11589, n11590, n11591, n11592, n11593, n11594,
         n11595, n11596, n11597, n11598, n11599, n11600, n11601, n11602,
         n11603, n11604, n11605, n11606, n11607, n11608, n11609, n11610,
         n11611, n11612, n11613, n11614, n11615, n11616, n11617, n11618,
         n11619, n11620, n11621, n11622, n11623, n11624, n11625, n11626,
         n11627, n11628, n11629, n11630, n11631, n11632, n11633, n11634,
         n11635, n11636, n11637, n11638, n11639, n11640, n11641, n11642,
         n11643, n11644, n11645, n11646, n11647, n11648, n11649, n11650,
         n11651, n11652, n11653, n11654, n11655, n11656, n11657, n11658,
         n11659, n11660, n11661, n11662, n11663, n11664, n11665, n11666,
         n11667, n11668, n11669, n11670, n11671, n11672, n11673, n11674,
         n11675, n11676, n11677, n11678, n11679, n11680, n11681, n11682,
         n11683, n11684, n11685, n11686, n11687, n11688, n11689, n11690,
         n11691, n11692, n11693, n11694, n11695, n11696, n11697, n11698,
         n11699, n11700, n11701, n11702, n11703, n11704, n11705, n11706,
         n11707, n11708, n11709, n11710, n11711, n11712, n11713, n11714,
         n11715, n11716, n11717, n11718, n11719, n11720, n11721, n11722,
         n11723, n11724, n11725, n11726, n11727, n11728, n11729, n11730,
         n11731, n11732, n11733, n11734, n11735, n11736, n11737, n11738,
         n11739, n11740, n11741, n11742, n11743, n11744, n11745, n11746,
         n11747, n11748, n11749, n11750, n11751, n11752, n11753, n11754,
         n11755, n11756, n11757, n11758, n11759, n11760, n11761, n11762,
         n11763, n11764, n11765, n11766, n11767, n11768, n11769, n11770,
         n11771, n11772, n11773, n11774, n11775, n11776, n11777, n11778,
         n11779, n11780, n11781, n11782, n11783, n11784, n11785, n11786,
         n11787, n11788, n11789, n11790, n11791, n11792, n11793, n11794,
         n11795, n11796, n11797, n11798, n11799, n11800, n11801, n11802,
         n11803, n11804, n11805, n11806, n11807, n11808, n11809, n11810,
         n11811, n11812, n11813, n11814, n11815, n11816, n11817, n11818,
         n11819, n11820, n11821, n11822, n11823, n11824, n11825, n11826,
         n11827, n11828, n11829, n11830, n11831, n11832, n11833, n11834,
         n11835, n11836, n11837, n11838, n11839, n11840, n11841, n11842,
         n11843, n11844, n11845, n11846, n11847, n11848, n11849, n11850,
         n11851, n11852, n11853, n11854, n11855, n11856, n11857, n11858,
         n11859, n11860, n11861, n11862, n11863, n11864, n11865, n11866,
         n11867, n11868, n11869, n11870, n11871, n11872, n11873, n11874,
         n11875, n11876, n11877, n11878, n11879, n11880, n11881, n11882,
         n11883, n11884, n11885, n11886, n11887, n11888, n11889, n11890,
         n11891, n11892, n11893, n11894, n11895, n11896, n11897, n11898,
         n11899, n11900, n11901, n11902, n11903, n11904, n11905, n11906,
         n11907, n11908, n11909, n11910, n11911, n11912, n11913, n11914,
         n11915, n11916, n11917, n11918, n11919, n11920, n11921, n11922,
         n11923, n11924, n11925, n11926, n11927, n11928, n11929, n11930,
         n11931, n11932, n11933, n11934, n11935, n11936, n11937, n11938,
         n11939, n11940, n11941, n11942, n11943, n11944, n11945, n11946,
         n11947, n11948, n11949, n11950, n11951, n11952, n11953, n11954,
         n11955, n11956, n11957, n11958, n11959, n11960, n11961, n11962,
         n11963, n11964, n11965, n11966, n11967, n11968, n11969, n11970,
         n11971, n11972, n11973, n11974, n11975, n11976, n11977, n11978,
         n11979, n11980, n11981, n11982, n11983, n11984, n11985, n11986,
         n11987, n11988, n11989, n11990, n11991, n11992, n11993, n11994,
         n11995, n11996, n11997, n11998, n11999, n12000, n12001, n12002,
         n12003, n12004, n12005, n12006, n12007, n12008, n12009, n12010,
         n12011, n12012, n12013, n12014, n12015, n12016, n12017, n12018,
         n12019, n12020, n12021, n12022, n12023, n12024, n12025, n12026,
         n12027, n12028, n12029, n12030, n12031, n12032, n12033, n12034,
         n12035, n12036, n12037, n12038, n12039, n12040, n12041, n12042,
         n12043, n12044, n12045, n12046, n12047, n12048, n12049, n12050,
         n12051, n12052, n12053, n12054, n12055, n12056, n12057, n12058,
         n12059, n12060, n12061, n12062, n12063, n12064, n12065, n12066,
         n12067, n12068, n12069, n12070, n12071, n12072, n12073, n12074,
         n12075, n12076, n12077, n12078, n12079, n12080, n12081, n12082,
         n12083, n12084, n12085, n12086, n12087, n12088, n12089, n12090,
         n12091, n12092, n12093, n12094, n12095, n12096, n12097, n12098,
         n12099, n12100, n12101, n12102, n12103, n12104, n12105, n12106,
         n12107, n12108, n12109, n12110, n12111, n12112, n12113, n12114,
         n12115, n12116, n12117, n12118, n12119, n12120, n12121, n12122,
         n12123, n12124, n12125, n12126, n12127, n12128, n12129, n12130,
         n12131, n12132, n12133, n12134, n12135, n12136, n12137, n12138,
         n12139, n12140, n12141, n12142, n12143, n12144, n12145, n12146,
         n12147, n12148, n12149, n12150, n12151, n12152, n12153, n12154,
         n12155, n12156, n12157, n12158, n12159, n12160, n12161, n12162,
         n12163, n12164, n12165, n12166, n12167, n12168, n12169, n12170,
         n12171, n12172, n12173, n12174, n12175, n12176, n12177, n12178,
         n12179, n12180, n12181, n12182, n12183, n12184, n12185, n12186,
         n12187, n12188, n12189, n12190, n12191, n12192, n12193, n12194,
         n12195, n12196, n12197, n12198, n12199, n12200, n12201, n12202,
         n12203, n12204, n12205, n12206, n12207, n12208, n12209, n12210,
         n12211, n12212, n12213, n12214, n12215, n12216, n12217, n12218,
         n12219, n12220, n12221, n12222, n12223, n12224, n12225, n12226,
         n12227, n12228, n12229, n12230, n12231, n12232, n12233, n12234,
         n12235, n12236, n12237, n12238, n12239, n12240, n12241, n12242,
         n12243, n12244, n12245, n12246, n12247, n12248, n12249, n12250,
         n12251, n12252, n12253, n12254, n12255, n12256, n12257, n12258,
         n12259, n12260, n12261, n12262, n12263, n12264, n12265, n12266,
         n12267, n12268, n12269, n12270, n12271, n12272, n12273, n12274,
         n12275, n12276, n12277, n12278, n12279, n12280, n12281, n12282,
         n12283, n12284, n12285, n12286, n12287, n12288, n12289, n12290,
         n12291, n12292, n12293, n12294, n12295, n12296, n12297, n12298,
         n12299, n12300, n12301, n12302, n12303, n12304, n12305, n12306,
         n12307, n12308, n12309, n12310, n12311, n12312, n12313, n12314,
         n12315, n12316, n12317, n12318, n12319, n12320, n12321, n12322,
         n12323, n12324, n12325, n12326, n12327, n12328, n12329, n12330,
         n12331, n12332, n12333, n12334, n12335, n12336, n12337, n12338,
         n12339, n12340, n12341, n12342, n12343, n12344, n12345, n12346,
         n12347, n12348, n12349, n12350, n12351, n12352, n12353, n12354,
         n12355, n12356, n12357, n12358, n12359, n12360, n12361, n12362,
         n12363, n12364, n12365, n12366, n12367, n12368, n12369, n12370,
         n12371, n12372, n12373, n12374, n12375, n12376, n12377, n12378,
         n12379, n12380, n12381, n12382, n12383, n12384, n12385, n12386,
         n12387, n12388, n12389, n12390, n12391, n12392, n12393, n12394,
         n12395, n12396, n12397, n12398, n12399, n12400, n12401, n12402,
         n12403, n12404, n12405, n12406, n12407, n12408, n12409, n12410,
         n12411, n12412, n12413, n12414, n12415, n12416, n12417, n12418,
         n12419, n12420, n12421, n12422, n12423, n12424, n12425, n12426,
         n12427, n12428, n12429, n12430, n12431, n12432, n12433, n12434,
         n12435, n12436, n12437, n12438, n12439, n12440, n12441, n12442,
         n12443, n12444, n12445, n12446, n12447, n12448, n12449, n12450,
         n12451, n12452, n12453, n12454, n12455, n12456, n12457, n12458,
         n12459, n12460, n12461, n12462, n12463, n12464, n12465, n12466,
         n12467, n12468, n12469, n12470, n12471, n12472, n12473, n12474,
         n12475, n12476, n12477, n12478, n12479, n12480, n12481, n12482,
         n12483, n12484, n12485, n12486, n12487, n12488, n12489, n12490,
         n12491, n12492, n12493, n12494, n12495, n12496, n12497, n12498,
         n12499, n12500, n12501, n12502, n12503, n12504, n12505, n12506,
         n12507, n12508, n12509, n12510, n12511, n12512, n12513, n12514,
         n12515, n12516, n12517, n12518, n12519, n12520, n12521, n12522,
         n12523, n12524, n12525, n12526, n12527, n12528, n12529, n12530,
         n12531, n12532, n12533, n12534, n12535, n12536, n12537, n12538,
         n12539, n12540, n12541, n12542, n12543, n12544, n12545, n12546,
         n12547, n12548, n12549, n12550, n12551, n12552, n12553, n12554,
         n12555, n12556, n12557, n12558, n12559, n12560, n12561, n12562,
         n12563, n12564, n12565, n12566, n12567, n12568, n12569, n12570,
         n12571, n12572, n12573, n12574, n12575, n12576, n12577, n12578,
         n12579, n12580, n12581, n12582, n12583, n12584, n12585, n12586,
         n12587, n12588, n12589, n12590, n12591, n12592, n12593, n12594,
         n12595, n12596, n12597, n12598, n12599, n12600, n12601, n12602,
         n12603, n12604, n12605, n12606, n12607, n12608, n12609, n12610,
         n12611, n12612, n12613, n12614, n12615, n12616, n12617, n12618,
         n12619, n12620, n12621, n12622, n12623, n12624, n12625, n12626,
         n12627, n12628, n12629, n12630, n12631, n12632, n12633, n12634,
         n12635, n12636, n12637, n12638, n12639, n12640, n12641, n12642,
         n12643, n12644, n12645, n12646, n12647, n12648, n12649, n12650,
         n12651, n12652, n12653, n12654, n12655, n12656, n12657, n12658,
         n12659, n12660, n12661, n12662, n12663, n12664, n12665, n12666,
         n12667, n12668, n12669, n12670, n12671, n12672, n12673, n12674,
         n12675, n12676, n12677, n12678, n12679, n12680, n12681, n12682,
         n12683, n12684, n12685, n12686, n12687, n12688, n12689, n12690,
         n12691, n12692, n12693, n12694, n12695, n12696, n12697, n12698,
         n12699, n12700, n12701, n12702, n12703, n12704, n12705, n12706,
         n12707, n12708, n12709, n12710, n12711, n12712, n12713, n12714,
         n12715, n12716, n12717, n12718, n12719, n12720, n12721, n12722,
         n12723, n12724, n12725, n12726, n12727, n12728, n12729, n12730,
         n12731, n12732, n12733, n12734, n12735, n12736, n12737, n12738,
         n12739, n12740, n12741, n12742, n12743, n12744, n12745, n12746,
         n12747, n12748, n12749, n12750, n12751, n12752, n12753, n12754,
         n12755, n12756, n12757, n12758, n12759, n12760, n12761, n12762,
         n12763, n12764, n12765, n12766, n12767, n12768, n12769, n12770,
         n12771, n12772, n12773, n12774, n12775, n12776, n12777, n12778,
         n12779, n12780, n12781, n12782, n12783, n12784, n12785, n12786,
         n12787, n12788, n12789, n12790, n12791, n12792, n12793, n12794,
         n12795, n12796, n12797, n12798, n12799, n12800, n12801, n12802,
         n12803, n12804, n12805, n12806, n12807, n12808, n12809, n12810,
         n12811, n12812, n12813, n12814, n12815, n12816, n12817, n12818,
         n12819, n12820, n12821, n12822, n12823, n12824, n12825, n12826,
         n12827, n12828, n12829, n12830, n12831, n12832, n12833, n12834,
         n12835, n12836, n12837, n12838, n12839, n12840, n12841, n12842,
         n12843, n12844, n12845, n12846, n12847, n12848, n12849, n12850,
         n12851, n12852, n12853, n12854, n12855, n12856, n12857, n12858,
         n12859, n12860, n12861, n12862, n12863, n12864, n12865, n12866,
         n12867, n12868, n12869, n12870, n12871, n12872, n12873, n12874,
         n12875, n12876, n12877, n12878, n12879, n12880, n12881, n12882,
         n12883, n12884, n12885, n12886, n12887, n12888, n12889, n12890,
         n12891, n12892, n12893, n12894, n12895, n12896, n12897, n12898,
         n12899, n12900, n12901, n12902, n12903, n12904, n12905, n12906,
         n12907, n12908, n12909, n12910, n12911, n12912, n12913, n12914,
         n12915, n12916, n12917, n12918, n12919, n12920, n12921, n12922,
         n12923, n12924, n12925, n12926, n12927, n12928, n12929, n12930,
         n12931, n12932, n12933, n12934, n12935, n12936, n12937, n12938,
         n12939, n12940, n12941, n12942, n12943, n12944, n12945, n12946,
         n12947, n12948, n12949, n12950, n12951, n12952, n12953, n12954,
         n12955, n12956, n12957, n12958, n12959, n12960, n12961, n12962,
         n12963, n12964, n12965, n12966, n12967, n12968, n12969, n12970,
         n12971, n12972, n12973, n12974, n12975, n12976, n12977, n12978,
         n12979, n12980, n12981, n12982, n12983, n12984, n12985, n12986,
         n12987, n12988, n12989, n12990, n12991, n12992, n12993, n12994,
         n12995, n12996, n12997, n12998, n12999, n13000, n13001, n13002,
         n13003, n13004, n13005, n13006, n13007, n13008, n13009, n13010,
         n13011, n13012, n13013, n13014, n13015, n13016, n13017, n13018,
         n13019, n13020, n13021, n13022, n13023, n13024, n13025, n13026,
         n13027, n13028, n13029, n13030, n13031, n13032, n13033, n13034,
         n13035, n13036, n13037, n13038, n13039, n13040, n13041, n13042,
         n13043, n13044, n13045, n13046, n13047, n13048, n13049, n13050,
         n13051, n13052, n13053, n13054, n13055, n13056, n13057, n13058,
         n13059, n13060, n13061, n13062, n13063, n13064, n13065, n13066,
         n13067, n13068, n13069, n13070, n13071, n13072, n13073, n13074,
         n13075, n13076, n13077, n13078, n13079, n13080, n13081, n13082,
         n13083, n13084, n13085, n13086, n13087, n13088, n13089, n13090,
         n13091, n13092, n13093, n13094, n13095, n13096, n13097, n13098,
         n13099, n13100, n13101, n13102, n13103, n13104, n13105, n13106,
         n13107, n13108, n13109, n13110, n13111, n13112, n13113, n13114,
         n13115, n13116, n13117, n13118, n13119, n13120, n13121, n13122,
         n13123, n13124, n13125, n13126, n13127, n13128, n13129, n13130,
         n13131, n13132, n13133, n13134, n13135, n13136, n13137, n13138,
         n13139, n13140, n13141, n13142, n13143, n13144, n13145, n13146,
         n13147, n13148, n13149, n13150, n13151, n13152, n13153, n13154,
         n13155, n13156, n13157, n13158, n13159, n13160, n13161, n13162,
         n13163, n13164, n13165, n13166, n13167, n13168, n13169, n13170,
         n13171, n13172, n13173, n13174, n13175, n13176, n13177, n13178,
         n13179, n13180, n13181, n13182, n13183, n13184, n13185, n13186,
         n13187, n13188, n13189, n13190, n13191, n13192, n13193, n13194,
         n13195, n13196, n13197, n13198, n13199, n13200, n13201, n13202,
         n13203, n13204, n13205, n13206, n13207, n13208, n13209, n13210,
         n13211, n13212, n13213, n13214, n13215, n13216, n13217, n13218,
         n13219, n13220, n13221, n13222, n13223, n13224, n13225, n13226,
         n13227, n13228, n13229, n13230, n13231, n13232, n13233, n13234,
         n13235, n13236, n13237, n13238, n13239, n13240, n13241, n13242,
         n13243, n13244, n13245, n13246, n13247, n13248, n13249, n13250,
         n13251, n13252, n13253, n13254, n13255, n13256, n13257, n13258,
         n13259, n13260, n13261, n13262, n13263, n13264, n13265, n13266,
         n13267, n13268, n13269, n13270, n13271, n13272, n13273, n13274,
         n13275, n13276, n13277, n13278, n13279, n13280, n13281, n13282,
         n13283, n13284, n13285, n13286, n13287, n13288, n13289, n13290,
         n13291, n13292, n13293, n13294, n13295, n13296, n13297, n13298,
         n13299, n13300, n13301, n13302, n13303, n13304, n13305, n13306,
         n13307, n13308, n13309, n13310, n13311, n13312, n13313, n13314,
         n13315, n13316, n13317, n13318, n13319, n13320, n13321, n13322,
         n13323, n13324, n13325, n13326, n13327, n13328, n13329, n13330,
         n13331, n13332, n13333, n13334, n13335, n13336, n13337, n13338,
         n13339, n13340, n13341, n13342, n13343, n13344, n13345, n13346,
         n13347, n13348, n13349, n13350, n13351, n13352, n13353, n13354,
         n13355, n13356, n13357, n13358, n13359, n13360, n13361, n13362,
         n13363, n13364, n13365, n13366, n13367, n13368, n13369, n13370,
         n13371, n13372, n13373, n13374, n13375, n13376, n13377, n13378,
         n13379, n13380, n13381, n13382, n13383, n13384, n13385, n13386,
         n13387, n13388, n13389, n13390, n13391, n13392, n13393, n13394,
         n13395, n13396, n13397, n13398, n13399, n13400, n13401, n13402,
         n13403, n13404, n13405, n13406, n13407, n13408, n13409, n13410,
         n13411, n13412, n13413, n13414, n13415, n13416, n13417, n13418,
         n13419, n13420, n13421, n13422, n13423, n13424, n13425, n13426,
         n13427, n13428, n13429, n13430, n13431, n13432, n13433, n13434,
         n13435, n13436, n13437, n13438, n13439, n13440, n13441, n13442,
         n13443, n13444, n13445, n13446, n13447, n13448, n13449, n13450,
         n13451, n13452, n13453, n13454, n13455, n13456, n13457, n13458,
         n13459, n13460, n13461, n13462, n13463, n13464, n13465, n13466,
         n13467, n13468, n13469, n13470, n13471, n13472, n13473, n13474,
         n13475, n13476, n13477, n13478, n13479, n13480, n13481, n13482,
         n13483, n13484, n13485, n13486, n13487, n13488, n13489, n13490,
         n13491, n13492, n13493, n13494, n13495, n13496, n13497, n13498,
         n13499, n13500, n13501, n13502, n13503, n13504, n13505, n13506,
         n13507, n13508, n13509, n13510, n13511, n13512, n13513, n13514,
         n13515, n13516, n13517, n13518, n13519, n13520, n13521, n13522,
         n13523, n13524, n13525, n13526, n13527, n13528, n13529, n13530,
         n13531, n13532, n13533, n13534, n13535, n13536, n13537, n13538,
         n13539, n13540, n13541, n13542, n13543, n13544, n13545, n13546,
         n13547, n13548, n13549, n13550, n13551, n13552, n13553, n13554,
         n13555, n13556, n13557, n13558, n13559, n13560, n13561, n13562,
         n13563, n13564, n13565, n13566, n13567, n13568, n13569, n13570,
         n13571, n13572, n13573, n13574, n13575, n13576, n13577, n13578,
         n13579, n13580, n13581, n13582, n13583, n13584, n13585, n13586,
         n13587, n13588, n13589, n13590, n13591, n13592, n13593, n13594,
         n13595, n13596, n13597, n13598, n13599, n13600, n13601, n13602,
         n13603, n13604, n13605, n13606, n13607, n13608, n13609, n13610,
         n13611, n13612, n13613, n13614, n13615, n13616, n13617, n13618,
         n13619, n13620, n13621, n13622, n13623, n13624, n13625, n13626,
         n13627, n13628, n13629, n13630, n13631, n13632, n13633, n13634,
         n13635, n13636, n13637, n13638, n13639, n13640, n13641, n13642,
         n13643, n13644, n13645, n13646, n13647, n13648, n13649, n13650,
         n13651, n13652, n13653, n13654, n13655, n13656, n13657, n13658,
         n13659, n13660, n13661, n13662, n13663, n13664, n13665, n13666,
         n13667, n13668, n13669, n13670, n13671, n13672, n13673, n13674,
         n13675, n13676, n13677, n13678, n13679, n13680, n13681, n13682,
         n13683, n13684, n13685, n13686, n13687, n13688, n13689, n13690,
         n13691, n13692, n13693, n13694, n13695, n13696, n13697, n13698,
         n13699, n13700, n13701, n13702, n13703, n13704, n13705, n13706,
         n13707, n13708, n13709, n13710, n13711, n13712, n13713, n13714,
         n13715, n13716, n13717, n13718, n13719, n13720, n13721, n13722,
         n13723, n13724, n13725, n13726, n13727, n13728, n13729, n13730,
         n13731, n13732, n13733, n13734, n13735, n13736, n13737, n13738,
         n13739, n13740, n13741, n13742, n13743, n13744, n13745, n13746,
         n13747, n13748, n13749, n13750, n13751, n13752, n13753, n13754,
         n13755, n13756, n13757, n13758, n13759, n13760, n13761, n13762,
         n13763, n13765, n13766, n13767, n13768, n13769, n13770, n13771,
         n13772, n13773, n13774, n13775, n13776, n13777, n13778, n13779,
         n13780, n13781, n13782, n13783, n13784, n13785, n13786, n13787,
         n13788, n13789, n13790, n13791, n13792, n13793, n13794, n13795,
         n13796, n13797, n13798, n13799, n13800, n13801, n13802, n13803,
         n13804, n13805, n13806, n13807, n13808, n13809, n13810, n13811,
         n13812, n13813, n13814, n13815, n13816, n13817, n13818, n13819,
         n13820, n13821, n13822, n13823, n13824, n13825, n13826, n13827,
         n13828, n13829, n13830, n13831, n13832, n13833, n13834, n13835,
         n13837, n13838, n13839, n13840, n13841, n13842, n13843, n13844,
         n13845, n13846, n13847, n13848, n13849, n13850, n13851, n13852,
         n13853, n13854, n13855, n13856, n13857, n13858, n13859, n13860,
         n13861, n13862, n13863, n13864, n13865, n13866, n13867, n13868,
         n13869, n13870, n13871, n13872, n13873, n13874, n13875, n13876,
         n13877, n13878, n13879, n13880, n13881, n13882, n13883, n13884,
         n13885, n13886, n13887, n13888, n13889, n13890, n13891, n13892,
         n13893, n13894, n13895, n13896, n13897, n13898, n13899, n13900,
         n13901, n13902, n13903, n13904, n13905, n13906, n13907, n13908,
         n13909, n13910, n13911, n13912, n13913, n13914, n13915, n13916,
         n13917, n13918, n13919, n13920, n13921, n13922, n13923, n13924,
         n13925, n13926, n13927, n13928, n13929, n13930, n13931, n13932,
         n13933, n13934, n13935, n13936, n13937, n13938, n13939, n13940,
         n13941, n13942, n13943, n13944, n13945, n13946, n13947, n13948,
         n13949, n13950, n13951, n13952, n13953, n13954, n13955, n13956,
         n13957, n13958, n13959, n13960, n13961, n13962, n13963, n13964,
         n13965, n13966, n13967, n13968, n13969, n13970, n13971, n13972,
         n13973, n13974, n13975, n13976, n13977, n13978, n13979, n13980,
         n13981, n13982, n13983, n13984, n13985, n13986, n13987, n13988,
         n13989, n13990, n13991, n13992, n13993, n13994, n13995, n13996,
         n13997, n13998, n13999, n14000, n14001, n14002, n14003, n14004,
         n14005, n14006, n14007, n14008, n14009, n14010, n14011, n14012,
         n14013, n14014, n14015, n14016, n14017, n14018, n14019, n14020,
         n14021, n14022, n14023, n14024, n14025, n14026, n14027, n14028,
         n14029, n14030, n14031, n14032, n14033, n14034, n14035, n14036,
         n14037, n14038, n14039, n14040, n14041, n14042, n14043, n14044,
         n14045, n14046, n14047, n14048, n14049, n14050, n14051, n14052,
         n14053, n14054, n14055, n14056, n14057, n14058, n14059, n14060,
         n14061, n14062, n14063, n14064, n14065, n14066, n14067, n14068,
         n14069, n14070, n14071, n14072, n14073, n14074, n14075, n14076,
         n14077, n14078, n14079, n14080, n14081, n14082, n14083, n14084,
         n14085, n14086, n14087, n14088, n14089, n14090, n14091, n14092,
         n14093, n14094, n14095, n14096, n14097, n14098, n14099, n14100,
         n14101, n14102, n14103, n14104, n14105, n14106, n14107, n14108,
         n14109, n14110, n14111, n14112, n14113, n14114, n14115, n14116,
         n14117, n14118, n14119, n14120, n14121, n14122, n14123, n14124,
         n14125, n14126, n14127, n14128, n14129, n14130, n14131, n14132,
         n14133, n14134, n14135, n14136, n14137, n14138, n14139, n14140,
         n14141, n14142, n14143, n14144, n14145, n14146, n14147, n14148,
         n14149, n14150, n14151, n14152, n14153, n14154, n14155, n14156,
         n14157, n14158, n14159, n14160, n14161, n14162, n14163, n14164,
         n14165, n14166, n14167, n14168, n14169, n14170, n14171, n14172,
         n14173, n14174, n14175, n14176, n14177, n14178, n14179, n14180,
         n14181, n14182, n14183, n14184, n14185, n14186, n14187, n14188,
         n14189, n14190, n14191, n14192, n14193, n14194, n14195, n14196,
         n14197, n14198, n14199, n14200, n14201, n14202, n14203, n14204,
         n14205, n14206, n14207, n14208, n14209, n14210, n14211, n14212,
         n14213, n14214, n14215, n14216, n14217, n14218, n14219, n14220,
         n14221, n14222, n14223, n14224, n14225, n14226, n14227, n14228,
         n14229, n14230, n14231, n14232, n14233, n14234, n14235, n14236,
         n14237, n14238, n14239, n14240, n14241, n14242, n14243, n14244,
         n14245, n14246, n14247, n14248, n14249, n14250, n14251, n14252,
         n14253, n14254, n14255, n14256, n14257, n14258, n14259, n14260,
         n14261, n14262, n14263, n14264, n14265, n14266, n14267, n14268,
         n14269, n14270, n14271, n14272, n14273, n14274, n14275, n14276,
         n14277, n14278, n14279, n14280, n14281, n14282, n14283, n14284,
         n14285, n14286, n14287, n14288, n14289, n14290, n14291, n14292,
         n14293, n14294, n14295, n14296, n14297, n14298, n14299, n14300,
         n14301, n14302, n14303, n14304, n14305, n14306, n14307, n14308,
         n14309, n14310, n14311, n14312, n14313, n14314, n14315, n14316,
         n14317, n14318, n14319, n14320, n14321, n14322, n14323, n14324,
         n14325, n14326, n14327, n14328, n14329, n14330, n14331, n14332,
         n14333, n14334, n14335, n14336, n14337, n14338, n14339, n14340,
         n14341, n14342, n14343, n14344, n14345, n14346, n14347, n14348,
         n14349, n14350, n14351, n14352, n14353, n14354, n14355, n14356,
         n14357, n14358, n14359, n14360, n14361, n14362, n14363, n14364,
         n14365, n14366, n14367, n14368, n14369, n14370, n14371, n14372,
         n14373, n14374, n14375, n14376, n14377, n14378, n14379, n14380,
         n14381, n14382, n14383, n14384, n14385, n14386, n14387, n14388,
         n14389, n14390, n14391, n14392, n14393, n14394, n14395, n14396,
         n14397, n14398, n14399, n14400, n14401, n14402, n14403, n14404,
         n14405, n14406, n14407, n14408, n14409, n14410, n14411, n14412,
         n14413, n14414, n14415, n14416, n14417, n14418, n14419, n14420,
         n14421, n14422, n14423, n14424, n14425, n14426, n14427, n14428,
         n14429, n14430, n14431, n14432, n14433, n14434, n14435, n14436,
         n14437, n14438, n14439, n14440, n14441, n14442, n14443, n14444,
         n14445, n14446, n14447, n14448, n14449, n14450, n14451, n14452,
         n14453, n14454, n14455, n14456, n14457, n14458, n14459, n14460,
         n14461, n14462, n14463, n14464, n14465, n14466, n14467, n14468,
         n14469, n14470, n14471, n14472, n14473, n14474, n14475, n14476,
         n14477, n14478, n14479, n14480, n14481, n14482, n14483, n14484,
         n14485, n14486, n14487, n14488, n14489, n14490, n14491, n14492,
         n14493, n14494, n14495, n14496, n14497, n14498, n14499, n14500,
         n14501, n14502, n14503, n14504, n14505, n14506, n14507, n14508,
         n14509, n14510, n14511, n14512, n14513, n14514, n14515, n14516,
         n14517, n14518, n14519, n14520, n14521, n14522, n14523, n14524,
         n14525, n14526, n14527, n14528, n14529, n14530, n14531, n14532,
         n14533, n14534, n14535, n14536, n14537, n14538, n14539, n14540,
         n14541, n14542, n14543, n14544, n14545, n14546, n14547, n14548,
         n14549, n14550, n14551, n14552, n14553, n14554, n14555, n14556,
         n14557, n14558, n14559, n14560, n14561, n14562, n14563, n14564,
         n14565, n14566, n14567, n14568, n14569, n14570, n14571, n14572,
         n14573, n14574, n14575, n14576, n14577, n14578, n14579, n14580,
         n14581, n14582, n14583, n14584, n14585, n14586, n14587, n14588,
         n14589, n14590, n14591, n14592, n14593, n14594, n14595, n14596,
         n14597, n14598, n14599, n14600, n14601, n14602, n14603, n14604,
         n14605, n14606, n14607, n14608, n14609, n14610, n14611, n14612,
         n14613, n14614, n14615, n14616, n14617, n14618, n14619, n14620,
         n14621, n14622, n14623, n14624, n14625, n14626, n14627, n14628,
         n14629, n14630, n14631, n14632, n14633, n14634, n14635, n14636,
         n14637, n14638, n14639, n14640, n14641, n14642, n14643, n14644,
         n14645, n14646, n14647, n14648, n14649, n14650, n14651, n14652,
         n14653, n14654, n14655, n14656, n14657, n14658, n14659, n14660,
         n14661, n14662, n14663, n14664, n14665, n14666, n14667, n14668,
         n14669, n14670, n14671, n14672, n14673, n14674, n14675, n14676,
         n14677, n14678, n14679, n14680, n14681, n14682, n14683, n14684,
         n14685, n14686, n14687, n14688, n14689, n14690, n14691, n14692,
         n14693, n14694, n14695, n14696, n14697, n14698, n14699, n14700,
         n14701, n14702, n14703, n14704, n14705, n14706, n14707, n14708,
         n14709, n14710, n14711, n14712, n14713, n14714, n14715, n14716,
         n14717, n14718, n14719, n14720, n14721, n14722, n14723, n14724,
         n14725, n14726, n14727, n14728, n14729, n14730, n14731, n14732,
         n14733, n14734, n14735, n14736, n14737, n14738, n14739, n14740,
         n14741, n14742, n14743, n14744, n14745, n14746, n14747, n14748,
         n14749, n14750, n14751, n14752, n14753, n14754, n14755, n14756,
         n14757, n14758, n14759, n14760, n14761, n14762, n14763, n14764,
         n14765, n14766, n14767, n14768, n14769, n14770, n14771, n14772,
         n14773, n14774, n14775, n14776, n14777, n14778, n14779, n14780,
         n14781, n14782, n14783, n14784, n14785, n14786, n14787, n14788,
         n14789, n14790, n14791, n14792, n14793, n14794, n14795, n14796,
         n14797, n14798, n14799, n14800, n14801, n14802, n14803, n14804,
         n14805, n14806, n14807, n14808, n14809, n14810, n14811, n14812,
         n14813, n14814, n14815, n14816, n14817, n14818, n14819, n14820,
         n14821, n14822, n14823, n14824, n14825, n14826, n14827, n14828,
         n14829, n14830, n14831, n14832, n14833, n14834, n14835, n14836,
         n14837, n14838, n14839, n14840, n14841, n14842, n14843, n14844,
         n14845, n14846, n14847, n14848, n14849, n14850, n14851, n14852,
         n14853, n14854, n14855, n14856, n14857, n14858, n14859, n14860,
         n14861, n14862, n14863, n14864, n14865, n14866, n14867, n14868,
         n14869, n14870, n14871, n14872, n14873, n14874, n14875, n14876,
         n14877, n14878, n14879, n14880, n14881, n14882, n14883, n14884,
         n14885, n14886, n14887, n14888, n14889, n14890, n14891, n14892,
         n14893, n14894, n14895, n14896, n14897, n14898, n14899, n14900,
         n14901, n14902, n14903, n14904, n14905, n14906, n14907, n14908,
         n14909, n14910, n14911, n14912, n14913, n14914, n14915, n14916,
         n14917, n14918, n14919, n14920, n14921, n14922, n14923, n14924,
         n14925, n14926, n14927, n14928, n14929, n14930, n14931, n14932,
         n14933, n14934, n14935, n14936, n14937, n14938, n14939, n14940,
         n14941, n14942, n14943, n14944, n14945, n14946, n14947, n14948,
         n14949, n14950, n14951, n14952, n14953, n14954, n14955, n14956,
         n14957, n14958, n14959, n14960, n14961, n14962, n14963, n14964,
         n14965, n14966, n14967, n14968, n14969, n14970, n14971, n14972,
         n14973, n14974, n14975, n14976, n14977, n14978, n14979, n14980,
         n14981, n14982, n14983, n14984, n14985, n14986, n14987, n14988,
         n14989, n14990, n14991, n14992, n14993, n14994, n14995, n14996,
         n14997, n14998, n14999, n15000, n15001, n15002, n15003, n15004,
         n15005, n15006, n15007, n15008, n15009, n15010, n15011, n15012,
         n15013, n15014, n15015, n15016, n15017, n15018, n15019, n15020,
         n15021, n15022, n15023, n15024, n15025, n15026, n15027, n15028,
         n15029, n15030, n15031, n15032, n15033, n15034, n15035, n15036,
         n15037, n15038, n15039, n15040, n15041, n15042, n15043, n15044,
         n15045, n15046, n15047, n15048, n15049, n15050, n15051, n15052,
         n15053, n15054, n15055, n15056, n15057, n15058, n15059, n15060,
         n15061, n15062, n15063, n15064, n15065, n15066, n15067, n15068,
         n15069, n15070, n15071, n15072, n15073, n15074, n15075, n15076,
         n15077, n15078, n15079, n15080, n15081, n15082, n15083, n15084,
         n15085, n15086, n15087, n15088, n15089, n15090, n15091, n15092,
         n15093, n15094, n15095, n15096, n15097, n15098, n15099, n15100,
         n15101, n15102, n15103, n15104, n15105, n15106, n15107, n15108,
         n15109, n15110, n15111, n15112, n15113, n15114, n15115, n15116,
         n15117, n15118, n15119, n15120, n15121, n15122, n15123, n15124,
         n15125, n15126, n15127, n15128, n15129, n15130, n15131, n15132,
         n15133, n15134, n15135, n15136, n15137, n15138, n15139, n15140,
         n15141, n15142, n15143, n15144, n15145, n15146, n15147, n15148,
         n15149, n15150, n15151, n15152, n15153, n15154, n15155, n15156,
         n15157, n15158, n15159, n15160, n15161, n15162, n15163, n15164,
         n15165, n15166, n15167, n15168, n15169, n15170, n15171, n15172,
         n15173, n15174, n15175, n15176, n15177, n15178, n15179, n15180,
         n15181, n15182, n15183, n15184, n15185, n15186, n15187, n15188,
         n15189, n15190, n15191, n15192, n15193, n15194, n15195, n15196,
         n15197, n15198, n15199, n15200, n15201, n15202, n15203, n15204,
         n15205, n15206, n15207, n15208, n15209, n15210, n15211, n15212,
         n15213, n15214, n15215, n15216, n15217, n15218, n15219, n15220,
         n15221, n15222, n15223, n15224, n15225, n15226, n15227, n15228,
         n15229, n15230, n15231, n15232, n15233, n15234, n15235, n15236,
         n15237, n15238, n15239, n15240, n15241, n15242, n15243, n15244,
         n15245, n15246, n15247, n15248, n15249, n15250, n15251, n15252,
         n15253, n15254, n15255, n15256, n15257, n15258, n15259, n15260,
         n15261, n15262, n15263, n15264, n15265, n15266, n15267, n15268,
         n15269, n15270, n15271, n15272, n15273, n15274, n15275, n15276,
         n15277, n15278, n15279, n15280, n15281, n15282, n15283, n15284,
         n15285, n15286, n15287, n15288, n15289, n15290, n15291, n15292,
         n15293, n15294, n15295, n15296, n15297, n15298, n15299, n15300,
         n15301, n15302, n15303, n15304, n15305, n15306, n15307, n15308,
         n15309, n15310, n15311, n15312, n15313, n15314, n15315, n15316,
         n15317, n15318, n15319, n15320, n15321, n15322, n15323, n15324,
         n15325, n15326, n15327, n15328, n15329, n15330, n15331, n15332,
         n15333, n15334, n15335, n15336, n15337, n15338, n15339, n15340,
         n15341, n15342, n15343, n15344, n15345, n15346, n15347, n15348,
         n15349, n15350, n15351, n15352, n15353, n15354, n15355, n15356,
         n15357, n15358, n15359, n15360, n15361, n15362, n15363, n15364,
         n15365, n15366, n15367, n15368, n15369, n15370, n15371, n15372,
         n15373, n15374, n15375, n15376, n15377, n15378, n15379, n15380,
         n15381, n15382, n15383, n15384, n15385, n15386, n15387, n15388,
         n15389, n15390, n15391, n15392, n15393, n15394, n15395, n15396,
         n15397, n15398, n15399, n15400, n15401, n15402, n15403, n15404,
         n15405, n15406, n15407, n15408, n15409, n15410, n15411, n15412,
         n15413, n15414, n15415, n15416, n15417, n15418, n15419, n15420,
         n15421, n15422, n15423, n15424, n15425, n15426, n15427, n15428,
         n15429, n15430, n15431, n15432, n15433, n15434, n15435, n15436,
         n15437, n15438, n15439, n15440, n15441, n15442, n15443, n15444,
         n15445, n15446, n15447, n15448, n15449, n15450, n15451, n15452,
         n15453, n15454, n15455, n15456, n15457, n15458, n15459, n15460,
         n15461, n15462, n15463, n15464, n15465, n15466, n15467, n15468,
         n15469, n15470, n15471, n15472, n15473, n15474, n15475, n15476,
         n15477, n15478, n15479, n15480, n15481, n15482, n15483, n15484,
         n15485, n15486, n15487, n15488, n15489, n15490, n15491, n15492,
         n15493, n15494, n15495, n15496, n15497, n15498, n15499, n15500,
         n15501, n15502, n15503, n15504, n15505, n15506, n15507, n15508,
         n15509, n15510, n15511, n15512, n15513, n15514, n15515, n15516,
         n15517, n15518, n15519, n15520, n15521, n15522, n15523, n15524,
         n15525, n15526, n15527, n15528, n15529, n15530, n15531, n15532,
         n15533, n15534, n15535, n15536, n15537, n15538, n15539, n15540,
         n15541, n15542, n15543, n15544, n15545, n15546, n15547, n15548,
         n15549, n15550, n15551, n15552, n15553, n15554, n15555, n15556,
         n15557, n15558, n15559, n15560, n15561, n15562, n15563, n15564,
         n15565, n15566, n15567, n15568, n15569, n15570, n15571, n15572,
         n15573, n15574, n15575, n15576, n15577, n15578, n15579, n15580,
         n15581, n15582, n15583, n15584, n15585, n15586, n15587, n15588,
         n15589, n15590, n15591, n15592, n15593, n15594, n15595, n15596,
         n15597, n15598, n15599, n15600, n15601, n15602, n15603, n15604,
         n15605, n15606, n15607, n15608, n15609, n15610, n15611, n15612,
         n15613, n15614, n15615, n15616, n15617, n15618, n15619, n15620,
         n15621, n15622, n15623, n15624, n15625, n15626, n15627, n15628,
         n15629, n15630, n15631, n15632, n15633, n15634, n15635, n15636,
         n15637, n15638, n15639, n15640, n15641, n15642, n15643, n15644,
         n15645, n15646, n15647, n15648, n15649, n15650, n15651, n15652,
         n15653, n15654, n15655, n15656, n15657, n15658, n15659, n15660,
         n15661, n15662, n15663, n15664, n15665, n15666, n15667, n15668,
         n15669, n15670, n15671, n15672, n15673, n15674, n15675, n15676,
         n15677, n15678, n15679, n15680, n15681, n15682, n15683, n15684,
         n15685, n15686, n15687, n15688, n15689, n15690, n15691, n15692,
         n15693, n15694, n15695, n15696, n15697, n15698, n15699, n15700,
         n15701, n15702, n15703, n15704, n15705, n15706, n15707, n15708,
         n15709, n15710, n15711, n15712, n15713, n15714, n15715, n15716,
         n15717, n15718, n15719, n15720, n15721, n15722, n15723, n15724,
         n15725, n15726, n15727, n15728, n15729, n15730, n15731, n15732,
         n15733, n15734, n15735, n15736, n15737, n15738, n15739, n15740,
         n15741, n15742, n15743, n15744, n15745, n15746, n15747, n15748,
         n15749, n15750, n15751, n15752, n15753, n15754, n15755, n15756,
         n15757, n15758, n15759, n15760, n15761, n15762, n15763, n15764,
         n15765, n15766, n15767, n15768, n15769, n15770, n15771, n15772,
         n15773, n15774, n15775, n15776, n15777, n15778, n15779, n15780,
         n15781, n15782, n15783, n15784, n15785, n15786, n15787, n15788,
         n15789, n15790, n15791, n15792, n15793, n15794, n15795, n15796,
         n15797, n15798, n15799, n15800, n15801, n15802, n15803, n15804,
         n15805, n15806, n15807, n15808, n15809, n15810, n15811, n15812,
         n15813, n15814, n15815, n15816, n15817, n15818, n15819, n15820,
         n15821, n15822, n15823, n15824, n15825, n15826, n15827, n15828,
         n15829, n15830, n15831, n15832, n15833, n15834, n15835, n15836,
         n15837, n15838, n15839, n15840, n15841, n15842, n15843, n15844,
         n15845, n15846, n15847, n15848, n15849, n15850, n15851, n15852,
         n15853, n15854, n15855, n15856, n15857, n15858, n15859, n15860,
         n15861, n15862, n15863, n15864, n15865, n15866, n15867, n15868,
         n15869, n15870, n15871, n15872, n15873, n15874, n15875, n15876,
         n15877, n15878, n15879, n15880, n15881, n15882, n15883, n15884,
         n15885, n15886, n15887, n15888, n15889, n15890, n15891, n15892,
         n15893, n15894, n15895, n15896, n15897, n15898, n15899, n15900,
         n15901, n15902, n15903, n15904, n15905, n15906, n15907, n15908,
         n15909, n15910, n15911, n15912, n15913, n15914, n15915, n15916,
         n15917, n15918, n15919, n15920, n15921, n15922, n15923, n15924,
         n15925, n15926, n15927, n15928, n15929, n15930, n15931, n15932,
         n15933, n15934, n15935, n15936, n15937, n15938, n15939, n15940,
         n15941, n15942, n15943, n15944, n15945, n15946, n15947, n15948,
         n15949, n15950, n15951, n15952, n15953, n15954, n15955, n15956,
         n15957, n15958, n15959, n15960, n15961, n15962, n15963, n15964,
         n15965, n15966, n15967, n15968, n15969, n15970, n15971, n15972,
         n15973, n15974, n15975, n15976, n15977, n15978, n15979, n15980,
         n15981, n15982, n15983, n15984, n15985, n15986, n15987, n15988,
         n15989, n15990, n15991, n15992, n15993, n15994, n15995, n15996,
         n15997, n15998, n15999, n16000, n16001, n16002, n16003, n16004,
         n16005, n16006, n16007, n16008, n16009, n16010, n16011, n16012,
         n16013, n16014, n16015, n16016, n16017, n16018, n16019, n16020,
         n16021, n16022, n16023, n16024, n16025, n16026, n16027, n16028,
         n16029, n16030, n16031, n16032, n16033, n16034, n16035, n16036,
         n16037, n16038, n16039, n16040, n16041, n16042, n16043, n16044,
         n16045, n16046, n16047, n16048, n16049, n16050, n16051, n16052,
         n16053, n16054, n16055, n16056, n16057, n16058, n16059, n16060,
         n16061, n16062, n16063, n16064, n16065, n16066, n16067, n16068,
         n16069, n16070, n16071, n16072, n16073, n16074, n16075, n16076,
         n16077, n16078, n16079, n16080, n16081, n16082, n16083, n16084,
         n16085, n16086, n16087, n16088, n16089, n16090, n16091, n16092,
         n16093, n16094, n16095, n16096, n16097, n16098, n16099, n16100,
         n16101, n16102, n16103, n16104, n16105, n16106, n16107, n16108,
         n16109, n16110, n16111, n16112, n16113, n16114, n16115, n16116,
         n16117, n16118, n16119, n16120, n16121, n16122, n16123, n16124,
         n16125, n16126, n16127, n16128, n16129, n16130, n16131, n16132,
         n16133, n16134, n16135, n16136, n16137, n16138, n16139, n16140,
         n16141, n16142, n16143, n16144, n16145, n16146, n16147, n16148,
         n16149, n16150, n16151, n16152, n16153, n16154, n16155, n16156,
         n16157, n16158, n16159, n16160, n16161, n16162, n16163, n16164,
         n16165, n16166, n16167, n16168, n16169, n16170, n16171, n16172,
         n16173, n16174, n16175, n16176, n16177, n16178, n16179, n16180,
         n16181, n16182, n16183, n16184, n16185, n16186, n16187, n16188,
         n16189, n16190, n16191, n16192, n16193, n16194, n16195, n16196,
         n16197, n16198, n16199, n16200, n16201, n16202, n16203, n16204,
         n16205, n16206, n16207, n16208, n16209, n16210, n16211, n16212,
         n16213, n16214, n16215, n16216, n16217, n16218, n16219, n16220,
         n16221, n16222, n16223, n16224, n16225, n16226, n16227, n16228,
         n16229, n16230, n16231, n16232, n16233, n16234, n16235, n16236,
         n16237, n16238, n16239, n16240, n16241, n16242, n16243, n16244,
         n16245, n16246, n16247, n16248, n16249, n16250, n16251, n16252,
         n16253, n16254, n16255, n16256, n16257, n16258, n16259, n16260,
         n16261, n16262, n16263, n16264, n16265, n16266, n16267, n16268,
         n16269, n16270, n16271, n16272, n16273, n16274, n16275, n16276,
         n16277, n16278, n16279, n16280, n16281, n16282, n16283, n16284,
         n16285, n16286, n16287, n16288, n16289, n16290, n16291, n16292,
         n16293, n16294, n16295, n16296, n16297, n16298, n16299, n16300,
         n16301, n16302, n16303, n16304, n16305, n16306, n16307, n16308,
         n16309, n16310, n16311, n16312, n16313, n16314, n16315, n16316,
         n16317, n16318, n16319, n16320, n16321, n16322, n16323, n16324,
         n16325, n16326, n16327, n16328, n16329, n16330, n16331, n16332,
         n16333, n16334, n16335, n16336, n16337, n16338, n16339, n16340,
         n16341, n16342, n16343, n16344, n16345, n16346, n16347, n16348,
         n16349, n16350, n16351, n16352, n16353, n16354, n16355, n16356,
         n16357, n16358, n16359, n16360, n16361, n16362, n16363, n16364,
         n16365, n16366, n16367, n16368, n16369, n16370, n16371, n16372,
         n16373, n16374, n16375, n16376, n16377, n16378, n16379, n16380,
         n16381, n16382, n16383, n16384, n16385, n16386, n16387, n16388,
         n16389, n16390, n16391, n16392, n16393, n16394, n16395, n16396,
         n16397, n16398, n16399, n16400, n16401, n16402, n16403, n16404,
         n16405, n16406, n16407, n16408, n16409, n16410, n16411, n16412,
         n16413, n16414, n16415, n16416, n16417, n16418, n16419, n16420,
         n16421, n16422, n16423, n16424, n16425, n16426, n16427, n16428,
         n16429, n16430, n16431, n16432, n16433, n16434, n16435, n16436,
         n16437, n16438, n16439, n16440, n16441, n16442, n16443, n16444,
         n16445, n16446, n16447, n16448, n16449, n16450, n16451, n16452,
         n16453, n16454, n16455, n16456, n16457, n16458, n16459, n16460,
         n16461, n16462, n16463, n16464, n16465, n16466, n16467, n16468,
         n16469, n16470, n16471, n16472, n16473, n16474, n16475, n16476,
         n16477, n16478, n16479, n16480, n16481, n16482, n16483, n16484,
         n16485, n16486, n16487, n16488, n16489, n16490, n16491, n16492,
         n16493, n16494, n16495, n16496, n16497, n16498, n16499, n16500,
         n16501, n16502, n16503, n16504, n16505, n16506, n16507, n16508,
         n16509, n16510, n16511, n16512, n16513, n16514, n16515, n16516,
         n16517, n16518, n16519, n16520, n16521, n16522, n16523, n16524,
         n16525, n16526, n16527, n16528, n16529, n16530, n16531, n16532,
         n16533, n16534, n16535, n16536, n16537, n16538, n16539, n16540,
         n16541, n16542, n16543, n16544, n16545, n16546, n16547, n16548,
         n16549, n16550, n16551, n16552, n16553, n16554, n16555, n16556,
         n16557, n16558, n16559, n16560, n16561, n16562, n16563, n16564,
         n16565, n16566, n16567, n16568, n16569, n16570, n16571, n16572,
         n16573, n16574, n16575, n16576, n16577, n16578, n16579, n16580,
         n16581, n16582, n16583, n16584, n16585, n16586, n16587, n16588,
         n16589, n16590, n16591, n16592, n16593, n16594, n16595, n16596,
         n16597, n16598, n16599, n16600, n16601, n16602, n16603, n16604,
         n16605, n16606, n16607, n16608, n16609, n16610, n16611, n16612,
         n16613, n16614, n16615, n16616, n16617, n16618, n16619, n16620,
         n16621, n16622, n16623, n16624, n16625, n16626, n16627, n16628,
         n16629, n16630, n16631, n16632, n16633, n16634, n16635, n16636,
         n16637, n16638, n16639, n16640, n16641, n16642, n16643, n16644,
         n16645, n16646, n16647, n16648, n16649, n16650, n16651, n16652,
         n16653, n16654, n16655, n16656, n16657, n16658, n16659, n16660,
         n16661, n16662, n16663, n16664, n16665, n16666, n16667, n16668,
         n16669, n16670, n16671, n16672, n16673, n16674, n16675, n16676,
         n16677, n16678, n16679, n16680, n16681, n16682, n16683, n16684,
         n16685, n16686, n16687, n16688, n16689, n16690, n16691, n16692,
         n16693, n16694, n16695, n16696, n16697, n16698, n16699, n16700,
         n16701, n16702, n16703, n16704, n16705, n16706, n16707, n16708,
         n16709, n16710, n16711, n16712, n16713, n16714, n16715, n16716,
         n16717, n16718, n16719, n16720, n16721, n16722, n16723, n16724,
         n16725, n16726, n16727, n16728, n16729, n16730, n16731, n16732,
         n16733, n16734, n16735, n16736, n16737, n16738, n16739, n16740,
         n16741, n16742, n16743, n16744, n16745, n16746, n16747, n16748,
         n16749, n16750, n16751, n16752, n16753, n16754, n16755, n16756,
         n16757, n16758, n16759, n16760, n16761, n16762, n16763, n16764,
         n16765, n16766, n16767, n16768, n16769, n16770, n16771, n16772,
         n16773, n16774, n16775, n16776, n16777, n16778, n16779, n16780,
         n16781, n16782, n16783, n16784, n16785, n16786, n16787, n16788,
         n16789, n16790, n16791, n16792, n16793, n16794, n16795, n16796,
         n16797, n16798, n16799, n16800, n16801, n16802, n16803, n16804,
         n16805, n16806, n16807, n16808, n16809, n16810, n16811, n16812,
         n16813, n16814, n16815, n16816, n16817, n16818, n16819, n16820,
         n16821, n16822, n16823, n16824, n16825, n16826, n16827, n16828,
         n16829, n16830, n16831, n16832, n16833, n16834, n16835, n16836,
         n16837, n16838, n16839, n16840, n16841, n16842, n16843, n16844,
         n16845, n16846, n16847, n16848, n16849, n16850, n16851, n16852,
         n16853, n16854, n16855, n16856, n16857, n16858, n16859, n16860,
         n16861, n16862, n16863, n16864, n16865, n16866, n16867, n16868,
         n16869, n16870, n16871, n16872, n16873, n16874, n16875, n16876,
         n16877, n16878, n16879, n16880, n16881, n16882, n16883, n16884,
         n16885, n16886, n16887, n16888, n16889, n16890, n16891, n16892,
         n16893, n16894, n16895, n16896, n16897, n16898, n16899, n16900,
         n16901, n16902, n16903, n16904, n16905, n16906, n16907, n16908,
         n16909, n16910, n16911, n16912, n16913, n16914, n16915, n16916,
         n16917, n16918, n16919, n16920, n16921, n16922, n16923, n16924,
         n16925, n16926, n16927, n16928, n16929, n16930, n16931, n16932,
         n16933, n16934, n16935, n16936, n16937, n16938, n16939, n16940,
         n16941, n16942, n16943, n16944, n16945, n16946, n16947, n16948,
         n16949, n16950, n16951, n16952, n16953, n16954, n16955, n16956,
         n16957, n16958, n16959, n16960, n16961, n16962, n16963, n16964,
         n16965, n16966, n16967, n16968, n16969, n16970, n16971, n16972,
         n16973, n16974, n16975, n16976, n16977, n16978, n16979, n16980,
         n16981, n16982, n16983, n16984, n16985, n16986, n16987, n16988,
         n16989, n16990, n16991, n16992, n16993, n16994, n16995, n16996,
         n16997, n16998, n16999, n17000, n17001, n17002, n17003, n17004,
         n17005, n17006, n17007, n17008, n17009, n17010, n17011, n17012,
         n17013, n17014, n17015, n17016, n17017, n17018, n17019, n17020,
         n17021, n17022, n17023, n17024, n17025, n17026, n17027, n17028,
         n17029, n17030, n17031, n17032, n17033, n17034, n17035, n17036,
         n17037, n17038, n17039, n17040, n17041, n17042, n17043, n17044,
         n17045, n17046, n17047, n17048, n17049, n17050, n17051, n17052,
         n17053, n17054, n17055, n17056, n17057, n17058, n17059, n17060,
         n17061, n17062, n17063, n17064, n17065, n17066, n17067, n17068,
         n17069, n17070, n17071, n17072, n17073, n17074, n17075, n17076,
         n17077, n17078, n17079, n17080, n17081, n17082, n17083, n17084,
         n17085, n17086, n17087, n17088, n17089, n17090, n17091, n17092,
         n17093, n17094, n17095, n17096, n17097, n17098, n17099, n17100,
         n17101, n17102, n17103, n17104, n17105, n17106, n17107, n17108,
         n17109, n17110, n17111, n17112, n17113, n17114, n17115, n17116,
         n17117, n17118, n17119, n17120, n17121, n17122, n17123, n17124,
         n17125, n17126, n17127, n17128, n17129, n17130, n17131, n17132,
         n17133, n17134, n17135, n17136, n17137, n17138, n17139, n17140,
         n17141, n17142, n17143, n17144, n17145, n17146, n17147, n17148,
         n17149, n17150, n17151, n17152, n17153, n17154, n17155, n17156,
         n17157, n17158, n17159, n17160, n17161, n17162, n17163, n17164,
         n17165, n17166, n17167, n17168, n17169, n17170, n17171, n17172,
         n17173, n17174, n17175, n17176, n17177, n17178, n17179, n17180,
         n17181, n17182, n17183, n17184, n17185, n17186, n17187, n17188,
         n17189, n17190, n17191, n17192, n17193, n17194, n17195, n17196,
         n17197, n17198, n17199, n17200, n17201, n17202, n17203, n17204,
         n17205, n17206, n17207, n17208, n17209, n17210, n17211, n17212,
         n17213, n17214, n17215, n17216, n17217, n17218, n17219, n17220,
         n17221, n17222, n17223, n17224, n17225, n17226, n17227, n17228,
         n17229, n17230, n17231, n17232, n17233, n17234, n17235, n17236,
         n17237, n17238, n17239, n17240, n17241, n17242, n17243, n17244,
         n17245, n17246, n17247, n17248, n17249, n17250, n17251, n17252,
         n17253, n17254, n17255, n17256, n17257, n17258, n17259, n17260,
         n17261, n17262, n17263, n17264, n17265, n17266, n17267, n17268,
         n17269, n17270, n17271, n17272, n17273, n17274, n17275, n17276,
         n17277, n17278, n17279, n17280, n17281, n17282, n17283, n17284,
         n17285, n17286, n17287, n17288, n17289, n17290, n17291, n17292,
         n17293, n17294, n17295, n17296, n17297, n17298, n17299, n17300,
         n17301, n17302, n17303, n17304, n17305, n17306, n17307, n17308,
         n17309, n17310, n17311, n17312, n17313, n17314, n17315, n17316,
         n17317, n17318, n17319, n17320, n17321, n17322, n17323, n17324,
         n17325, n17326, n17327, n17328, n17329, n17330, n17331, n17332,
         n17333, n17334, n17335, n17336, n17337, n17338, n17339, n17340,
         n17341, n17342, n17343, n17344, n17345, n17346, n17347, n17348,
         n17349, n17350, n17351, n17352, n17353, n17354, n17355, n17356,
         n17357, n17358, n17359, n17360, n17361, n17362, n17363, n17364,
         n17365, n17366, n17367, n17368, n17369, n17370, n17371, n17372,
         n17373, n17374, n17375, n17376, n17377, n17378, n17379, n17380,
         n17381, n17382, n17383, n17384, n17385, n17386, n17387, n17388,
         n17389, n17390, n17391, n17392, n17393, n17394, n17395, n17396,
         n17397, n17398, n17399, n17400, n17401, n17402, n17403, n17404,
         n17405, n17406, n17407, n17408, n17409, n17410, n17411, n17412,
         n17413, n17414, n17415, n17416, n17417, n17418, n17419, n17420,
         n17421, n17422, n17423, n17424, n17425, n17426, n17427, n17428,
         n17429, n17430, n17431, n17432, n17433, n17434, n17435, n17436,
         n17437, n17438, n17439, n17440, n17441, n17442, n17443, n17444,
         n17445, n17446, n17447, n17448, n17449, n17450, n17451, n17452,
         n17453, n17454, n17455, n17456, n17457, n17458, n17459, n17460,
         n17461, n17462, n17463, n17464, n17465, n17466, n17467, n17468,
         n17469, n17470, n17471, n17472, n17473, n17474, n17475, n17476,
         n17477, n17478, n17479, n17480, n17481, n17482, n17483, n17484,
         n17485, n17486, n17487, n17488, n17489, n17490, n17491, n17492,
         n17493, n17494, n17495, n17496, n17497, n17498, n17499, n17500,
         n17501, n17502, n17503, n17504, n17505, n17506, n17507, n17508,
         n17509, n17510, n17511, n17512, n17513, n17514, n17515, n17516,
         n17517, n17518, n17519, n17520, n17521, n17522, n17523, n17524,
         n17525, n17526, n17527, n17528, n17529, n17530, n17531, n17532,
         n17533, n17534, n17535, n17536, n17537, n17538, n17539, n17540,
         n17541, n17542, n17543, n17544, n17545, n17546, n17547, n17548,
         n17549, n17550, n17551, n17552, n17553, n17554, n17555, n17556,
         n17557, n17558, n17559, n17560, n17561, n17562, n17563, n17564,
         n17565, n17566, n17567, n17568, n17569, n17570, n17571, n17572,
         n17573, n17574, n17575, n17576, n17577, n17578, n17579, n17580,
         n17581, n17582, n17583, n17584, n17585, n17586, n17587, n17588,
         n17589, n17590, n17591, n17592, n17593, n17594, n17595, n17596,
         n17597, n17598, n17599, n17600, n17601, n17602, n17603, n17604,
         n17605, n17606, n17607, n17608, n17609, n17610, n17611, n17612,
         n17613, n17614, n17615, n17616, n17617, n17618, n17619, n17620,
         n17621, n17622, n17623, n17624, n17625, n17626, n17627, n17628,
         n17629, n17630, n17631, n17632, n17633, n17634, n17635, n17636,
         n17637, n17638, n17639, n17640, n17641, n17642, n17643, n17644,
         n17645, n17646, n17647, n17648, n17649, n17650, n17651, n17652,
         n17653, n17654, n17655, n17656, n17657, n17658, n17659, n17660,
         n17661, n17662, n17663, n17664, n17665, n17666, n17667, n17668,
         n17669, n17670, n17671, n17672, n17673, n17674, n17675, n17676,
         n17677, n17678, n17679, n17680, n17681, n17682, n17683, n17684,
         n17685, n17686, n17687, n17688, n17689, n17690, n17691, n17692,
         n17693, n17694, n17695, n17696, n17697, n17698, n17699, n17700,
         n17701, n17702, n17703, n17704, n17705, n17706, n17707, n17708,
         n17709, n17710, n17711, n17712, n17713, n17714, n17715, n17716,
         n17717, n17718, n17719, n17720, n17721, n17722, n17723, n17724,
         n17725, n17726, n17727, n17728, n17729, n17730, n17731, n17732,
         n17733, n17734, n17735, n17736, n17737, n17738, n17739, n17740,
         n17741, n17742, n17743, n17744, n17745, n17746, n17747, n17748,
         n17749, n17750, n17751, n17752, n17753, n17754, n17755, n17756,
         n17757, n17758, n17759, n17760, n17761, n17762, n17763, n17764,
         n17765, n17766, n17767, n17768, n17769, n17770, n17771, n17772,
         n17773, n17774, n17775, n17776, n17777, n17778, n17779, n17780,
         n17781, n17782, n17783, n17784, n17785, n17786, n17787, n17788,
         n17789, n17790, n17791, n17792, n17793, n17794, n17795, n17796,
         n17797, n17798, n17799, n17800, n17801, n17802, n17803, n17804,
         n17805, n17806, n17807, n17808, n17809, n17810, n17811, n17812,
         n17813, n17814, n17815, n17816, n17817, n17818, n17819, n17820,
         n17821, n17822, n17823, n17824, n17825, n17826, n17827, n17828,
         n17829, n17830, n17831, n17832, n17833, n17834, n17835, n17836,
         n17837, n17838, n17839, n17840, n17841, n17842, n17843, n17844,
         n17845, n17846, n17847, n17848, n17849, n17850, n17851, n17852,
         n17853, n17854, n17855, n17856, n17857, n17858, n17859, n17860,
         n17861, n17862, n17863, n17864, n17865, n17866, n17867, n17868,
         n17869, n17870, n17871, n17872, n17873, n17874, n17875, n17876,
         n17877, n17878, n17879, n17880, n17881, n17882, n17883, n17884,
         n17885, n17886, n17887, n17888, n17889, n17890, n17891, n17892,
         n17893, n17894, n17895, n17896, n17897, n17898, n17899, n17900,
         n17901, n17902, n17903, n17904, n17905, n17906, n17907, n17908,
         n17909, n17910, n17911, n17912, n17913, n17914, n17915, n17916,
         n17917, n17918, n17919, n17920, n17921, n17922, n17923, n17924,
         n17925, n17926, n17927, n17928, n17929, n17930, n17931, n17932,
         n17933, n17934, n17935, n17936, n17937, n17938, n17939, n17940,
         n17941, n17942, n17943, n17944, n17945, n17946, n17947, n17948,
         n17949, n17950, n17951, n17952, n17953, n17954, n17955, n17956,
         n17957, n17958, n17959, n17960, n17961, n17962, n17963, n17964,
         n17965, n17966, n17967, n17968, n17969, n17970, n17971, n17972,
         n17973, n17974, n17975, n17976, n17977, n17978, n17979, n17980,
         n17981, n17982, n17983, n17984, n17985, n17986, n17987, n17988,
         n17989, n17990, n17991, n17992, n17993, n17994, n17995, n17996,
         n17997, n17998, n17999, n18000, n18001, n18002, n18003, n18004,
         n18005, n18006, n18007, n18008, n18009, n18010, n18011, n18012,
         n18013, n18014, n18015, n18016, n18017, n18018, n18019, n18020,
         n18021, n18022, n18023, n18024, n18025, n18026, n18027, n18028,
         n18029, n18030, n18031, n18032, n18033, n18034, n18035, n18036,
         n18037, n18038, n18039, n18040, n18041, n18042, n18043, n18044,
         n18045, n18046, n18047, n18048, n18049, n18050, n18051, n18052,
         n18053, n18054, n18055, n18056, n18057, n18058, n18059, n18060,
         n18061, n18062, n18063, n18064, n18065, n18066, n18067, n18068,
         n18069, n18070, n18071, n18072, n18073, n18074, n18075, n18076,
         n18077, n18078, n18079, n18080, n18081, n18082, n18083, n18084,
         n18085, n18086, n18087, n18088, n18089, n18090, n18091, n18092,
         n18093, n18094, n18095, n18096, n18097, n18098, n18099, n18100,
         n18101, n18102, n18103, n18104, n18105, n18106, n18107, n18108,
         n18109, n18110, n18111, n18112, n18113, n18114, n18115, n18116,
         n18117, n18118, n18119, n18120, n18121, n18122, n18123, n18124,
         n18125, n18126, n18127, n18128, n18129, n18130, n18131, n18132,
         n18133, n18134, n18135, n18136, n18137, n18138, n18139, n18140,
         n18141, n18142, n18143, n18144, n18145, n18146, n18147, n18148,
         n18149, n18150, n18151, n18152, n18153, n18154, n18155, n18156,
         n18157, n18158, n18159, n18160, n18161, n18162, n18163, n18164,
         n18165, n18166, n18167, n18168, n18169, n18170, n18171, n18172,
         n18173, n18174, n18175, n18176, n18177, n18178, n18179, n18180,
         n18181, n18182, n18183, n18184, n18185, n18186, n18187, n18188,
         n18189, n18190, n18191, n18192, n18193, n18194, n18195, n18196,
         n18197, n18198, n18199, n18200, n18201, n18202, n18203, n18204,
         n18205, n18206, n18207, n18208, n18209, n18210, n18211, n18212,
         n18213, n18214, n18215, n18216, n18217, n18218, n18219, n18220,
         n18221, n18222, n18223, n18224, n18225, n18226, n18227, n18228,
         n18229, n18230, n18231, n18232, n18233, n18234, n18235, n18236,
         n18237, n18238, n18239, n18240, n18241, n18242, n18243, n18244,
         n18245, n18246, n18247, n18248, n18249, n18250, n18251, n18252,
         n18253, n18254, n18255, n18256, n18257, n18258, n18259, n18260,
         n18261, n18262, n18263, n18264, n18265, n18266, n18267, n18268,
         n18269, n18270, n18271, n18272, n18273, n18274, n18275, n18276,
         n18277, n18278, n18279, n18280, n18281, n18282, n18283, n18284,
         n18285, n18286, n18287, n18288, n18289, n18290, n18291, n18292,
         n18293, n18294, n18295, n18296, n18297, n18298, n18299, n18300,
         n18301, n18302, n18303, n18304, n18305, n18306, n18307, n18308,
         n18309, n18310, n18311, n18312, n18313, n18314, n18315, n18316,
         n18317, n18318, n18319, n18320, n18321, n18322, n18323, n18324,
         n18325, n18326, n18327, n18328, n18329, n18330, n18331, n18332,
         n18333, n18334, n18335, n18336, n18337, n18338, n18339, n18340,
         n18341, n18342, n18343, n18344, n18345, n18346, n18347, n18348,
         n18349, n18350, n18351, n18352, n18353, n18354, n18355, n18356,
         n18357, n18358, n18359, n18360, n18361, n18362, n18363, n18364,
         n18365, n18366, n18367, n18368, n18369, n18370, n18371, n18372,
         n18373, n18374, n18375, n18376, n18377, n18378, n18379, n18380,
         n18381, n18382, n18383, n18384, n18385, n18386, n18387, n18388,
         n18389, n18390, n18391, n18392, n18393, n18394, n18395, n18396,
         n18397, n18398, n18399, n18400, n18401, n18402, n18403, n18404,
         n18405, n18406, n18407, n18408, n18409, n18410, n18411, n18412,
         n18413, n18414, n18415, n18416, n18417, n18418, n18419, n18420,
         n18421, n18422, n18423, n18424, n18425, n18426, n18427, n18428,
         n18429, n18430, n18431, n18432, n18433, n18434, n18435, n18436,
         n18437, n18438, n18439, n18440, n18441, n18442, n18443, n18444,
         n18445, n18446, n18447, n18448, n18449, n18450, n18451, n18452,
         n18453, n18454, n18455, n18456, n18457, n18458, n18459, n18460,
         n18461, n18462, n18463, n18464, n18465, n18466, n18467, n18468,
         n18469, n18470, n18471, n18472, n18473, n18474, n18475, n18476,
         n18477, n18478, n18479, n18480, n18481, n18482, n18483, n18484,
         n18485, n18486, n18487, n18488, n18489, n18490, n18491, n18492,
         n18493, n18494, n18495, n18496, n18497, n18498, n18499, n18500,
         n18501, n18502, n18503, n18504, n18505, n18506, n18507, n18508,
         n18509, n18510, n18511, n18512, n18513, n18514, n18515, n18516,
         n18517, n18518, n18519, n18520, n18521, n18522, n18523, n18524,
         n18525, n18526, n18527, n18528, n18529, n18530, n18531, n18532,
         n18533, n18534, n18535, n18536, n18537, n18538, n18539, n18540,
         n18541, n18542, n18543, n18544, n18545, n18546, n18547, n18548,
         n18549, n18550, n18551, n18552, n18553, n18554, n18555, n18556,
         n18557, n18558, n18559, n18560, n18561, n18562, n18563, n18564,
         n18565, n18566, n18567, n18568, n18569, n18570, n18571, n18572,
         n18573, n18574, n18575, n18576, n18577, n18578, n18579, n18580,
         n18581, n18582, n18583, n18584, n18585, n18586, n18587, n18588,
         n18589, n18590, n18591, n18592, n18593, n18594, n18595, n18596,
         n18597, n18598, n18599, n18600, n18601, n18602, n18603, n18604,
         n18605, n18606, n18607, n18608, n18609, n18610, n18611, n18612,
         n18613, n18614, n18615, n18616, n18617, n18618, n18619, n18620,
         n18621, n18622, n18623, n18624, n18625, n18626, n18627, n18628,
         n18629, n18630, n18631, n18632, n18633, n18634, n18635, n18636,
         n18637, n18638, n18639, n18640, n18641, n18642, n18643, n18644,
         n18645, n18646, n18647, n18648, n18649, n18650, n18651, n18652,
         n18653, n18654, n18655, n18656, n18657, n18658, n18659, n18660,
         n18661, n18662, n18663, n18664, n18665, n18666, n18667, n18668,
         n18669, n18670, n18671, n18672, n18673, n18674, n18675, n18676,
         n18677, n18678, n18679, n18680, n18681, n18682, n18683, n18684,
         n18685, n18686, n18687, n18688, n18689, n18690, n18691, n18692,
         n18693, n18694, n18695, n18696, n18697, n18698, n18699, n18700,
         n18701, n18702, n18703, n18704, n18705, n18706, n18707, n18708,
         n18709, n18710, n18711, n18712, n18713, n18714, n18715, n18716,
         n18717, n18718, n18719, n18720, n18721, n18722, n18723, n18724,
         n18725, n18726, n18727, n18728, n18729, n18730, n18731, n18732,
         n18733, n18734, n18735, n18736, n18737, n18738, n18739, n18740,
         n18741, n18742, n18743, n18744, n18745, n18746, n18747, n18748,
         n18749, n18750, n18751, n18752, n18753, n18754, n18755, n18756,
         n18757, n18758, n18759, n18760, n18761, n18762, n18763, n18764,
         n18765, n18766, n18767, n18768, n18769, n18770, n18771, n18772,
         n18773, n18774, n18775, n18776, n18777, n18778, n18779, n18780,
         n18781, n18782, n18783, n18784, n18785, n18786, n18787, n18788,
         n18789, n18790, n18791, n18792, n18793, n18794, n18795, n18796,
         n18797, n18798, n18799, n18800, n18801, n18802, n18803, n18804,
         n18805, n18806, n18807, n18808, n18809, n18810, n18811, n18812,
         n18813, n18814, n18815, n18816, n18817, n18818, n18819, n18820,
         n18821, n18822, n18823, n18824, n18825, n18826, n18827, n18828,
         n18829, n18830, n18831, n18832, n18833, n18834, n18835, n18836,
         n18837, n18838, n18839, n18840, n18841, n18842, n18843, n18844,
         n18845, n18846, n18847, n18848, n18849, n18850, n18851, n18852,
         n18853, n18854, n18855, n18856, n18857, n18858, n18859, n18860,
         n18861, n18862, n18863, n18864, n18865, n18866, n18867, n18868,
         n18869, n18870, n18871, n18872, n18873, n18874, n18875, n18876,
         n18877, n18878, n18879, n18880, n18881, n18882, n18883, n18884,
         n18885, n18886, n18887, n18888, n18889, n18890, n18891, n18892,
         n18893, n18894, n18895, n18896, n18897, n18898, n18899, n18900,
         n18901, n18902, n18903, n18904, n18905, n18906, n18907, n18908,
         n18909, n18910, n18911, n18912, n18913, n18914, n18915, n18916,
         n18917, n18918, n18919, n18920, n18921, n18922, n18923, n18924,
         n18925, n18926, n18927, n18928, n18929, n18930, n18931, n18932,
         n18933, n18934, n18935, n18936, n18937, n18938, n18939, n18940,
         n18941, n18942, n18943, n18944, n18945, n18946, n18947, n18948,
         n18949, n18950, n18951, n18952, n18953, n18954, n18955, n18956,
         n18957, n18958, n18959, n18960, n18961, n18962, n18963, n18964,
         n18965, n18966, n18967, n18968, n18969, n18970, n18971, n18972,
         n18973, n18974, n18975, n18976, n18977, n18978, n18979, n18980,
         n18981, n18982, n18983, n18984, n18985, n18986, n18987, n18988,
         n18989, n18990, n18991, n18992, n18993, n18994, n18995, n18996,
         n18997, n18998, n18999, n19000, n19001, n19002, n19003, n19004,
         n19005, n19006, n19007, n19008, n19009, n19010, n19011, n19012,
         n19013, n19014, n19015, n19016, n19017, n19018, n19019, n19020,
         n19021, n19022, n19023, n19024, n19025, n19026, n19027, n19028,
         n19029, n19030, n19031, n19032, n19033, n19034, n19035, n19036,
         n19037, n19038, n19039, n19040, n19041, n19042, n19043, n19044,
         n19045, n19046, n19047, n19048, n19049, n19050, n19051, n19052,
         n19053, n19054, n19055, n19056, n19057, n19058, n19059, n19060,
         n19061, n19062, n19063, n19064, n19065, n19066, n19067, n19068,
         n19069, n19070, n19071, n19072, n19073, n19074, n19075, n19076,
         n19077, n19078, n19079, n19080, n19081, n19082, n19083, n19084,
         n19085, n19086, n19087, n19088, n19089, n19090, n19091, n19092,
         n19093, n19094, n19095, n19096, n19097, n19098, n19099, n19100,
         n19101, n19102, n19103, n19104, n19105, n19106, n19107, n19108,
         n19109, n19110, n19111, n19112, n19113, n19114, n19115, n19116,
         n19117, n19118, n19119, n19120, n19121, n19122, n19123, n19124,
         n19125, n19126, n19127, n19128, n19129, n19130, n19131, n19132,
         n19133, n19134, n19135, n19136, n19137, n19138, n19139, n19140,
         n19141, n19142, n19143, n19144, n19145, n19146, n19147, n19148,
         n19149, n19150, n19151, n19152, n19153, n19154, n19155, n19156,
         n19157, n19158, n19159, n19160, n19161, n19162, n19163, n19164,
         n19165, n19166, n19167, n19168, n19169, n19170, n19171, n19172,
         n19173, n19174, n19175, n19176, n19177, n19178, n19179, n19180,
         n19181, n19182, n19183, n19184, n19185, n19186, n19187, n19188,
         n19189, n19190, n19191, n19192, n19193, n19194, n19195, n19196,
         n19197, n19198, n19199, n19200, n19201, n19202, n19203, n19204,
         n19205, n19206, n19207, n19208, n19209, n19210, n19211, n19212,
         n19213, n19214, n19215, n19216, n19217, n19218, n19219, n19220,
         n19221, n19222, n19223, n19224, n19225, n19226, n19227, n19228,
         n19229, n19230, n19231, n19232, n19233, n19234, n19235, n19236,
         n19237, n19238, n19239, n19240, n19241, n19242, n19243, n19244,
         n19245, n19246, n19247, n19248, n19249, n19250, n19251, n19252,
         n19253, n19254, n19255, n19256, n19257, n19258, n19259, n19260,
         n19261, n19262, n19263, n19264, n19265, n19266, n19267, n19268,
         n19269, n19270, n19271, n19272, n19273, n19274, n19275, n19276,
         n19277, n19278, n19279, n19280, n19281, n19282, n19283, n19284,
         n19285, n19286, n19287, n19288, n19289, n19290, n19291, n19292,
         n19293, n19294, n19295, n19296, n19297, n19298, n19299, n19300,
         n19301, n19302, n19303, n19304, n19305, n19306, n19307, n19308,
         n19309, n19310, n19311, n19312, n19313, n19314, n19315, n19316,
         n19317, n19318, n19319, n19320, n19321, n19322, n19323, n19324,
         n19325, n19326, n19327, n19328, n19329, n19330, n19331, n19332,
         n19333, n19334, n19335, n19336, n19337, n19338, n19339, n19340,
         n19341, n19342, n19343, n19344, n19345, n19346, n19347, n19348,
         n19349, n19350, n19351, n19352, n19353, n19354, n19355, n19356,
         n19357, n19358, n19359, n19360, n19361, n19362, n19363, n19364,
         n19365, n19366, n19367, n19368, n19369, n19370, n19371, n19372,
         n19373, n19374, n19375, n19376, n19377, n19378, n19379, n19380,
         n19381, n19382, n19383, n19384, n19385, n19386, n19387, n19388,
         n19389, n19390, n19391, n19392, n19393, n19394, n19395, n19396,
         n19397, n19398, n19399, n19400, n19401, n19402, n19403, n19404,
         n19405, n19406, n19407, n19408, n19409, n19410, n19411, n19412,
         n19413, n19414, n19415, n19416, n19417, n19418, n19419, n19420,
         n19421, n19422, n19423, n19424, n19425, n19426, n19427, n19428,
         n19429, n19430, n19431, n19432, n19433, n19434, n19435, n19436,
         n19437, n19438, n19439, n19440, n19441, n19442, n19443, n19444,
         n19445, n19446, n19447, n19448, n19449, n19450, n19451, n19452,
         n19453, n19454, n19455, n19456, n19457, n19458, n19459, n19460,
         n19461, n19462, n19463, n19464, n19465, n19466, n19467, n19468,
         n19469, n19470, n19471, n19472, n19473, n19474, n19475, n19476,
         n19477, n19478, n19479, n19480, n19481, n19482, n19483, n19484,
         n19485, n19486, n19487, n19488, n19489, n19490, n19491, n19492,
         n19493, n19494, n19495, n19496, n19497, n19498, n19499, n19500,
         n19501, n19502, n19503, n19504, n19505, n19506, n19507, n19508,
         n19509, n19510, n19511, n19512, n19513, n19514, n19515, n19516,
         n19517, n19518, n19519, n19520, n19521, n19522, n19523, n19524,
         n19525, n19526, n19527, n19528, n19529, n19530, n19531, n19532,
         n19533, n19534, n19535, n19536, n19537, n19538, n19539, n19540,
         n19541, n19542, n19543, n19544, n19545, n19546, n19547, n19548,
         n19549, n19550, n19551, n19552, n19553, n19554, n19555, n19556,
         n19557, n19558, n19559, n19560, n19561, n19562, n19563, n19564,
         n19565, n19566, n19567, n19568, n19569, n19570, n19571, n19572,
         n19573, n19574, n19575, n19576, n19577, n19578, n19579, n19580,
         n19581, n19582, n19583, n19584, n19585, n19586, n19587, n19588,
         n19589, n19590, n19591, n19592, n19593, n19594, n19595, n19596,
         n19597, n19598, n19599, n19600, n19601, n19602, n19603, n19604,
         n19605, n19606, n19607, n19608, n19609, n19610, n19611, n19612,
         n19613, n19614, n19615, n19616, n19617, n19618, n19619, n19620,
         n19621, n19622, n19623, n19624, n19625, n19626, n19627, n19628,
         n19629, n19630, n19631, n19632, n19633, n19634, n19635, n19636,
         n19637, n19638, n19639, n19640, n19641, n19642, n19643, n19644,
         n19645, n19646, n19647, n19648, n19649, n19650, n19651, n19652,
         n19653, n19654, n19655, n19656, n19657, n19658, n19659, n19660,
         n19661, n19662, n19663, n19664, n19665, n19666, n19667, n19668,
         n19669, n19670, n19671, n19672, n19673, n19674, n19675, n19676,
         n19677, n19678, n19679, n19680, n19681, n19682, n19683, n19684,
         n19685, n19686, n19687, n19688, n19689, n19690, n19691, n19692,
         n19693, n19694, n19695, n19696, n19697, n19698, n19699, n19700,
         n19701, n19702, n19703, n19704, n19705, n19706, n19707, n19708,
         n19709, n19710, n19711, n19712, n19713, n19714, n19715, n19716,
         n19717, n19718, n19719, n19720, n19721, n19722, n19723, n19724,
         n19725, n19726, n19727, n19728, n19729, n19730, n19731, n19732,
         n19733, n19734, n19735, n19736, n19737, n19738, n19739, n19740,
         n19741, n19742, n19743, n19744, n19745, n19746, n19747, n19748,
         n19749, n19750, n19751, n19752, n19753, n19754, n19755, n19756,
         n19757, n19758, n19759, n19760, n19761, n19762, n19763, n19764,
         n19765, n19766, n19767, n19768, n19769, n19770, n19771, n19772,
         n19773, n19774, n19775, n19776, n19777, n19778, n19779, n19780,
         n19781, n19782, n19783, n19784, n19785, n19786, n19787, n19788,
         n19789, n19790, n19791, n19792, n19793, n19794, n19795, n19796,
         n19797, n19798, n19799, n19800, n19801, n19802, n19803, n19804,
         n19805, n19806, n19807, n19808, n19809, n19810, n19811, n19812,
         n19813, n19814, n19815, n19816, n19817, n19818, n19819, n19820,
         n19821, n19822, n19823, n19824, n19825, n19826, n19827, n19828,
         n19829, n19830, n19831, n19832, n19833, n19834, n19835, n19836,
         n19837, n19838, n19839, n19840, n19841, n19842, n19843, n19844,
         n19845, n19846, n19847, n19848, n19849, n19850, n19851, n19852,
         n19853, n19854, n19855, n19856, n19857, n19858, n19859, n19860,
         n19861, n19862, n19863, n19864, n19865, n19866, n19867, n19868,
         n19869, n19870, n19871, n19872, n19873, n19874, n19875, n19876,
         n19877, n19878, n19879, n19880, n19881, n19882, n19883, n19884,
         n19885, n19886, n19887, n19888, n19889, n19890, n19891, n19892,
         n19893, n19894, n19895, n19896, n19897, n19898, n19899, n19900,
         n19901, n19902, n19903, n19904, n19905, n19906, n19907, n19908,
         n19909, n19910, n19911, n19912, n19913, n19914, n19915, n19916,
         n19917, n19918, n19919, n19920, n19921, n19922, n19923, n19924,
         n19925, n19926, n19927, n19928, n19929, n19930, n19931, n19932,
         n19933, n19934, n19935, n19936, n19937, n19938, n19939, n19940,
         n19941, n19942, n19943, n19944, n19945, n19946, n19947, n19948,
         n19949, n19950, n19951, n19952, n19953, n19954, n19955, n19956,
         n19957, n19958, n19959, n19960, n19961, n19962, n19963, n19964,
         n19965, n19967, n19968, n19969, n19970, n19971, n19972, n19973,
         n19974, n19975, n19976, n19977, n19978, n19979, n19980, n19981,
         n19982, n19983, n19984, n19985, n19986, n19987, n19988, n19989,
         n19990, n19991, n19992, n19993, n19994, n19995, n19996, n19997,
         n19998, n19999, n20000, n20001, n20002, n20003, n20004, n20005,
         n20006, n20007, n20008, n20009, n20010, n20011, n20012, n20013,
         n20014, n20015, n20016, n20017, n20018, n20019, n20020, n20021,
         n20022, n20023, n20024, n20025, n20026, n20027, n20028, n20029,
         n20030, n20031, n20032, n20033, n20034, n20035, n20036, n20037,
         n20038, n20039, n20040, n20041, n20042, n20043, n20044, n20045,
         n20046, n20047, n20048, n20049, n20050, n20051, n20052, n20053,
         n20054, n20055, n20056, n20057, n20058, n20059, n20060, n20061,
         n20062, n20063, n20064, n20065, n20066, n20067, n20068, n20069,
         n20070, n20071, n20072, n20073, n20074, n20075, n20076, n20077,
         n20078, n20079, n20080, n20081, n20082, n20083, n20084, n20085,
         n20086, n20087, n20088, n20089, n20090, n20091, n20092, n20093,
         n20094, n20095, n20096, n20097, n20098, n20099, n20100, n20101,
         n20102, n20103, n20104, n20105, n20106, n20107, n20108, n20109,
         n20110, n20111, n20112, n20113, n20114, n20115, n20116, n20117,
         n20118, n20119, n20120, n20121, n20122, n20123, n20124, n20125,
         n20126, n20127, n20128, n20129, n20130, n20131, n20132, n20133,
         n20134, n20135, n20136, n20137, n20138, n20139, n20140, n20141,
         n20142, n20143, n20144, n20145, n20146, n20147, n20148, n20149,
         n20150, n20151, n20152, n20153, n20154, n20155, n20156, n20157,
         n20158, n20159, n20160, n20161, n20162, n20163, n20164, n20165,
         n20166, n20167, n20168, n20169, n20170, n20171, n20172, n20173,
         n20174, n20175, n20176, n20177, n20178, n20179, n20180, n20181,
         n20182, n20183, n20184, n20185, n20186, n20187, n20188, n20189,
         n20190, n20191, n20192, n20193, n20194, n20195, n20196, n20197,
         n20198, n20199, n20200, n20201, n20202, n20203, n20204, n20205,
         n20206, n20207, n20208, n20209, n20210, n20211, n20212, n20213,
         n20214, n20215, n20216, n20217, n20218, n20219, n20220, n20221,
         n20222, n20223, n20224, n20225, n20226, n20227, n20228, n20229,
         n20230, n20231, n20232, n20233, n20234, n20235, n20236, n20237,
         n20238, n20239, n20240, n20241, n20242, n20243, n20244, n20245,
         n20246, n20247, n20248, n20249, n20250, n20251, n20252, n20253,
         n20254, n20255, n20256, n20257, n20258, n20259, n20260, n20261,
         n20262, n20263, n20264, n20265, n20266, n20267, n20268, n20269,
         n20270, n20271, n20272, n20273, n20274, n20275, n20276, n20277,
         n20278, n20279, n20280, n20281, n20282, n20283, n20284, n20285,
         n20286, n20287, n20288, n20289, n20290, n20291, n20292, n20293,
         n20294, n20295, n20296, n20297, n20298, n20299, n20300, n20301,
         n20302, n20303, n20304, n20305, n20306, n20307, n20308, n20309,
         n20310, n20311, n20312, n20313, n20314, n20315, n20316, n20317,
         n20318, n20319, n20320, n20321, n20322, n20323, n20324, n20325,
         n20326, n20327, n20328, n20329, n20330, n20331, n20332, n20333,
         n20334, n20335, n20336, n20337, n20338, n20339, n20340, n20341,
         n20342, n20343, n20344, n20345, n20346, n20347, n20348, n20349,
         n20350, n20351, n20352, n20353, n20354, n20355, n20356, n20357,
         n20358, n20359, n20360, n20361, n20362, n20363, n20364, n20365,
         n20366, n20367, n20368, n20369, n20370, n20371, n20372, n20373,
         n20374, n20375, n20376, n20377, n20378, n20379, n20380, n20381,
         n20382, n20383, n20384, n20385, n20386, n20387, n20388, n20389,
         n20390, n20391, n20392, n20393, n20394, n20395, n20396, n20397,
         n20398, n20399, n20400, n20401, n20402, n20403, n20404, n20405,
         n20406, n20407, n20408, n20409, n20410, n20411, n20412, n20413,
         n20414, n20415, n20416, n20417, n20418, n20419, n20420, n20421,
         n20422, n20423, n20424, n20425, n20426, n20427, n20428, n20429,
         n20430, n20431, n20432, n20433, n20434, n20435, n20436, n20437,
         n20438, n20439, n20440, n20441, n20442, n20443, n20444, n20445,
         n20446, n20447, n20448, n20449, n20450, n20451, n20452, n20453,
         n20454, n20455, n20456, n20457, n20458, n20459, n20460, n20461,
         n20462, n20463, n20464, n20465, n20466, n20467, n20468, n20469,
         n20470, n20471, n20472, n20473, n20474, n20475, n20476, n20477,
         n20478, n20479, n20480, n20481, n20482, n20483, n20484, n20485,
         n20486, n20487, n20488, n20489, n20490, n20491, n20492, n20493,
         n20494, n20495, n20496, n20497, n20498, n20499, n20500, n20501,
         n20502, n20503, n20504, n20505, n20506, n20507, n20508, n20509,
         n20510, n20511, n20512, n20513, n20514, n20515, n20516, n20517,
         n20518, n20519, n20520, n20521, n20522, n20523, n20524, n20525,
         n20526, n20527, n20528, n20529, n20530, n20531, n20532, n20533,
         n20534, n20535, n20536, n20537, n20538, n20539, n20540, n20541,
         n20542, n20543, n20544, n20545, n20546, n20547, n20548, n20549,
         n20550, n20551, n20552, n20553, n20554, n20555, n20556, n20557,
         n20558, n20559, n20560, n20561, n20562, n20563, n20564, n20565,
         n20566, n20567, n20568, n20569, n20570, n20571, n20572, n20573,
         n20574, n20575, n20576, n20577, n20578, n20579, n20580, n20581,
         n20582, n20583, n20584, n20585, n20586, n20587, n20588, n20589,
         n20590, n20591, n20592, n20593, n20594, n20595, n20596, n20597,
         n20598, n20599, n20600, n20601, n20602, n20603, n20604, n20605,
         n20606, n20607, n20608, n20609, n20610, n20611, n20612, n20613,
         n20614, n20615, n20616, n20617, n20618, n20619, n20620, n20621,
         n20622, n20623, n20624, n20625, n20626, n20627, n20628, n20629,
         n20630, n20631, n20632, n20633, n20634, n20635, n20636, n20637,
         n20638, n20639, n20640, n20641, n20642, n20643, n20644, n20645,
         n20646, n20647, n20648, n20649, n20650, n20651, n20652, n20653,
         n20654, n20655, n20656, n20657, n20658, n20659, n20660, n20661,
         n20662, n20663, n20664, n20665, n20666, n20667, n20668, n20669,
         n20670, n20671, n20672, n20673, n20674, n20675, n20676, n20677,
         n20678, n20679, n20680, n20681, n20682, n20683, n20684, n20685,
         n20686, n20687, n20688, n20689, n20690, n20691, n20692, n20693,
         n20694, n20695, n20696, n20697, n20698, n20699, n20700, n20701,
         n20702, n20703, n20704, n20705, n20706, n20707, n20708, n20709,
         n20710, n20711, n20712, n20713, n20714, n20715, n20716, n20717,
         n20718, n20719, n20720, n20721, n20722, n20723, n20724, n20725,
         n20726, n20727, n20728, n20729, n20730, n20731, n20732, n20733,
         n20734, n20735, n20736, n20737, n20738, n20739, n20740, n20741,
         n20742, n20743, n20744, n20745, n20746, n20747, n20748, n20749,
         n20750, n20751, n20752, n20753, n20754, n20755, n20756, n20757,
         n20758, n20759, n20760, n20761, n20762, n20763, n20764, n20765,
         n20766, n20767, n20768, n20769, n20770, n20771, n20772, n20773,
         n20774, n20775, n20776, n20777, n20778, n20779, n20780, n20781,
         n20782, n20783, n20784, n20785, n20786, n20787, n20788, n20789,
         n20790, n20791, n20792, n20793, n20794, n20795, n20796, n20797,
         n20798, n20799, n20800, n20801, n20802, n20803, n20804, n20805,
         n20806, n20807, n20808, n20809, n20810, n20811, n20812, n20813,
         n20814, n20815, n20816, n20817, n20818, n20819, n20820, n20821,
         n20822, n20823, n20824, n20825, n20826, n20827, n20828, n20829,
         n20830, n20831, n20832, n20833, n20834, n20835, n20836, n20837,
         n20838, n20839, n20840, n20841, n20842, n20843, n20844, n20845,
         n20846, n20847, n20848, n20849, n20850, n20851, n20852, n20853,
         n20854, n20855, n20856, n20857, n20858, n20859, n20860, n20861,
         n20862, n20863, n20864, n20865, n20866, n20867, n20868, n20869,
         n20870, n20871, n20872, n20873, n20874, n20875, n20876, n20877,
         n20878, n20879, n20880, n20881, n20882, n20883, n20884, n20885,
         n20886, n20887, n20888, n20889, n20890, n20891, n20892, n20893,
         n20894, n20895, n20896, n20897, n20898, n20899, n20900, n20901,
         n20902, n20903, n20904, n20905, n20906, n20907, n20908, n20909,
         n20910, n20911, n20912, n20913, n20914, n20915, n20916, n20917,
         n20918, n20919, n20920, n20921, n20922, n20923, n20924, n20925,
         n20926, n20927, n20928, n20929, n20930, n20931, n20932, n20933,
         n20934, n20935, n20936, n20937, n20938, n20939, n20940, n20941,
         n20942, n20943, n20944, n20945, n20946, n20947, n20948, n20949,
         n20950, n20951, n20952, n20953, n20954, n20955, n20956, n20957,
         n20958, n20959, n20960, n20961, n20962, n20963, n20964, n20965,
         n20966, n20967, n20968, n20969, n20970, n20971, n20972, n20973,
         n20974, n20975, n20976, n20977, n20978, n20979, n20980, n20981,
         n20982, n20983;

  AOI21_X2 U11163 ( .B1(n18453), .B2(n18458), .A(n18452), .ZN(n18465) );
  INV_X1 U11164 ( .A(n9750), .ZN(n14354) );
  NOR2_X1 U11165 ( .A1(n16098), .A2(n16099), .ZN(n16097) );
  INV_X2 U11167 ( .A(n17551), .ZN(n17585) );
  CLKBUF_X2 U11168 ( .A(n10456), .Z(n11599) );
  NAND2_X1 U11169 ( .A1(n13015), .A2(n13014), .ZN(n13234) );
  NAND2_X1 U11170 ( .A1(n12454), .A2(n12453), .ZN(n12693) );
  CLKBUF_X1 U11171 ( .A(n12330), .Z(n13944) );
  XNOR2_X1 U11172 ( .A(n12636), .B(n12635), .ZN(n10216) );
  OAI22_X1 U11173 ( .A1(n12631), .A2(P1_STATE2_REG_0__SCAN_IN), .B1(n13238), 
        .B2(n12630), .ZN(n12636) );
  INV_X2 U11174 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n12396) );
  CLKBUF_X2 U11175 ( .A(n10981), .Z(n11515) );
  NAND2_X1 U11176 ( .A1(n11136), .A2(n11116), .ZN(n11221) );
  NAND2_X1 U11177 ( .A1(n20119), .A2(n12433), .ZN(n12528) );
  INV_X1 U11180 ( .A(n16837), .ZN(n16954) );
  BUF_X1 U11181 ( .A(n16986), .Z(n15286) );
  BUF_X1 U11182 ( .A(n15264), .Z(n15254) );
  CLKBUF_X2 U11183 ( .A(n15149), .Z(n17000) );
  CLKBUF_X2 U11184 ( .A(n13869), .Z(n9732) );
  AND2_X2 U11185 ( .A1(n10833), .A2(n10359), .ZN(n10581) );
  INV_X1 U11186 ( .A(n16837), .ZN(n16987) );
  INV_X1 U11187 ( .A(n9785), .ZN(n11806) );
  NAND2_X2 U11188 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18624), .ZN(
        n11736) );
  INV_X1 U11189 ( .A(n12564), .ZN(n20026) );
  AND2_X4 U11190 ( .A1(n10112), .A2(n12783), .ZN(n12709) );
  INV_X1 U11191 ( .A(n9737), .ZN(n9739) );
  AND2_X1 U11192 ( .A1(n12781), .A2(n14515), .ZN(n12658) );
  AND2_X2 U11193 ( .A1(n9900), .A2(n12778), .ZN(n12783) );
  NAND2_X1 U11194 ( .A1(n10317), .A2(n10316), .ZN(n10391) );
  NAND2_X1 U11195 ( .A1(n10339), .A2(n10340), .ZN(n10426) );
  AND2_X2 U11196 ( .A1(n13185), .A2(n10876), .ZN(n10375) );
  AND2_X1 U11197 ( .A1(n10507), .A2(n9955), .ZN(n10500) );
  NOR2_X1 U11198 ( .A1(n18449), .A2(n18469), .ZN(n17887) );
  NOR2_X1 U11199 ( .A1(n12545), .A2(n12344), .ZN(n12349) );
  INV_X1 U11200 ( .A(n9737), .ZN(n9741) );
  BUF_X2 U11201 ( .A(n12127), .Z(n9755) );
  INV_X1 U11202 ( .A(n10391), .ZN(n10910) );
  AND2_X1 U11203 ( .A1(n12014), .A2(n12783), .ZN(n12127) );
  AND2_X1 U11204 ( .A1(n12783), .A2(n14515), .ZN(n13718) );
  INV_X2 U11205 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n9900) );
  NOR2_X1 U11206 ( .A1(n11354), .A2(n10383), .ZN(n10925) );
  CLKBUF_X3 U11207 ( .A(n10499), .Z(n10843) );
  NAND2_X1 U11208 ( .A1(n10056), .A2(n10054), .ZN(n12430) );
  INV_X1 U11209 ( .A(n20669), .ZN(n13383) );
  NAND2_X1 U11211 ( .A1(n12387), .A2(n12386), .ZN(n10111) );
  NAND2_X1 U11212 ( .A1(n11491), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n16047) );
  INV_X1 U11213 ( .A(n9793), .ZN(n16988) );
  NAND2_X1 U11214 ( .A1(n9917), .A2(n12535), .ZN(n12804) );
  AND2_X1 U11215 ( .A1(n12681), .A2(n12680), .ZN(n12775) );
  CLKBUF_X2 U11216 ( .A(n13402), .Z(n9750) );
  NAND2_X1 U11217 ( .A1(n19740), .A2(n10927), .ZN(n10869) );
  BUF_X1 U11218 ( .A(n10418), .Z(n19085) );
  OR2_X1 U11219 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n16736) );
  AOI21_X1 U11221 ( .B1(n14548), .B2(n10807), .A(n14540), .ZN(n14534) );
  OAI21_X1 U11222 ( .B1(n15511), .B2(n15510), .A(n18648), .ZN(n17192) );
  INV_X1 U11223 ( .A(n19860), .ZN(n19829) );
  INV_X1 U11224 ( .A(n11986), .ZN(n11148) );
  INV_X1 U11225 ( .A(n15084), .ZN(n11154) );
  AND4_X1 U11226 ( .A1(n10126), .A2(n10125), .A3(n13132), .A4(n10124), .ZN(
        n13265) );
  NAND2_X1 U11227 ( .A1(n10843), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9719) );
  NAND2_X2 U11228 ( .A1(n11196), .A2(n11487), .ZN(n11490) );
  NAND2_X2 U11229 ( .A1(n10352), .A2(n10351), .ZN(n10353) );
  AND2_X4 U11230 ( .A1(n10401), .A2(n10330), .ZN(n10368) );
  AND2_X2 U11231 ( .A1(n17419), .A2(n9896), .ZN(n17357) );
  NAND2_X2 U11232 ( .A1(n17458), .A2(n17551), .ZN(n17419) );
  NAND2_X2 U11233 ( .A1(n10345), .A2(n9791), .ZN(n10354) );
  NAND3_X2 U11234 ( .A1(n11816), .A2(n11815), .A3(n11814), .ZN(n18046) );
  NOR2_X1 U11236 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n17332), .ZN(
        n17331) );
  MUX2_X2 U11237 ( .A(n12093), .B(n12096), .S(n12564), .Z(n12094) );
  OR2_X2 U11238 ( .A1(n12092), .A2(n12091), .ZN(n12564) );
  NAND2_X2 U11239 ( .A1(n14534), .A2(n14533), .ZN(n14535) );
  XNOR2_X2 U11240 ( .A(n11439), .B(n11438), .ZN(n11690) );
  AND2_X4 U11241 ( .A1(n10501), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10517) );
  BUF_X1 U11242 ( .A(n12067), .Z(n9721) );
  CLKBUF_X1 U11243 ( .A(n12067), .Z(n9722) );
  AND2_X1 U11244 ( .A1(n12783), .A2(n14516), .ZN(n12067) );
  AND2_X4 U11245 ( .A1(n10843), .A2(n10359), .ZN(n10542) );
  NOR2_X4 U11246 ( .A1(n11736), .A2(n11735), .ZN(n15162) );
  NAND2_X2 U11247 ( .A1(n18617), .A2(n18607), .ZN(n11735) );
  AND2_X1 U11248 ( .A1(n12781), .A2(n14516), .ZN(n13869) );
  INV_X4 U11249 ( .A(n9719), .ZN(n9723) );
  XNOR2_X2 U11250 ( .A(n12430), .B(n12362), .ZN(n12394) );
  NOR2_X2 U11251 ( .A1(n17574), .A2(n16238), .ZN(n17460) );
  AOI211_X1 U11252 ( .C1(n16054), .C2(n15837), .A(n14763), .B(n14762), .ZN(
        n14764) );
  OR2_X1 U11253 ( .A1(n14761), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n9935) );
  XNOR2_X1 U11254 ( .A(n13974), .B(n13889), .ZN(n14229) );
  AND2_X1 U11255 ( .A1(n14279), .A2(n10002), .ZN(n14263) );
  CLKBUF_X1 U11256 ( .A(n13997), .Z(n14011) );
  OR2_X1 U11257 ( .A1(n14200), .A2(n14199), .ZN(n15676) );
  AND2_X1 U11258 ( .A1(n9894), .A2(n9893), .ZN(n17309) );
  CLKBUF_X1 U11259 ( .A(n11503), .Z(n11504) );
  NAND2_X1 U11260 ( .A1(n9895), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n17321) );
  NAND2_X1 U11261 ( .A1(n11248), .A2(n9891), .ZN(n11477) );
  AND2_X1 U11262 ( .A1(n13289), .A2(n10184), .ZN(n14612) );
  OR2_X1 U11263 ( .A1(n17357), .A2(n17719), .ZN(n9897) );
  BUF_X2 U11264 ( .A(n13402), .Z(n9749) );
  NAND2_X1 U11265 ( .A1(n13380), .A2(n13379), .ZN(n13402) );
  OR2_X1 U11266 ( .A1(n14103), .A2(n14093), .ZN(n14095) );
  NAND2_X1 U11267 ( .A1(n11126), .A2(n11154), .ZN(n19308) );
  NAND2_X1 U11268 ( .A1(n11126), .A2(n15084), .ZN(n19374) );
  NAND2_X1 U11269 ( .A1(n11149), .A2(n11148), .ZN(n12999) );
  NAND2_X1 U11270 ( .A1(n9794), .A2(n11148), .ZN(n19340) );
  BUF_X1 U11271 ( .A(n12813), .Z(n9751) );
  OR3_X2 U11272 ( .A1(n11146), .A2(n11153), .A3(n11133), .ZN(n19167) );
  AND2_X1 U11273 ( .A1(n11146), .A2(n11145), .ZN(n11149) );
  INV_X2 U11274 ( .A(n17674), .ZN(n17646) );
  CLKBUF_X2 U11275 ( .A(n11113), .Z(n11153) );
  OR2_X1 U11276 ( .A1(n17599), .A2(n17902), .ZN(n15341) );
  CLKBUF_X2 U11277 ( .A(n11115), .Z(n15084) );
  CLKBUF_X2 U11278 ( .A(n16219), .Z(n9742) );
  OR2_X1 U11279 ( .A1(n12425), .A2(n12427), .ZN(n12428) );
  AOI21_X1 U11280 ( .B1(n18032), .B2(n11828), .A(n15208), .ZN(n15222) );
  NAND4_X1 U11281 ( .A1(n9789), .A2(n12349), .A3(n10203), .A4(n10204), .ZN(
        n10202) );
  NOR2_X1 U11282 ( .A1(n12342), .A2(n12537), .ZN(n10204) );
  AND3_X1 U11283 ( .A1(n10264), .A2(n12118), .A3(n12539), .ZN(n13415) );
  NAND2_X1 U11284 ( .A1(n20026), .A2(n12469), .ZN(n12909) );
  BUF_X1 U11285 ( .A(n12187), .Z(n20034) );
  CLKBUF_X3 U11286 ( .A(n13936), .Z(n9724) );
  OR2_X2 U11287 ( .A1(n12030), .A2(n12029), .ZN(n12121) );
  INV_X1 U11288 ( .A(n10389), .ZN(n10406) );
  INV_X2 U11289 ( .A(n20010), .ZN(n9725) );
  CLKBUF_X2 U11290 ( .A(n12658), .Z(n12367) );
  CLKBUF_X2 U11291 ( .A(n13843), .Z(n13868) );
  CLKBUF_X2 U11292 ( .A(n12126), .Z(n12619) );
  CLKBUF_X2 U11294 ( .A(n13862), .Z(n13707) );
  CLKBUF_X2 U11296 ( .A(n15149), .Z(n15294) );
  BUF_X4 U11297 ( .A(n15118), .Z(n9726) );
  OR2_X1 U11298 ( .A1(n11735), .A2(n18478), .ZN(n10274) );
  AND2_X1 U11299 ( .A1(n11447), .A2(n10876), .ZN(n10376) );
  INV_X2 U11301 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n15822) );
  NAND3_X2 U11302 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10286) );
  CLKBUF_X2 U11303 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n16164) );
  OR2_X1 U11304 ( .A1(n14909), .A2(n16139), .ZN(n9936) );
  AND2_X1 U11305 ( .A1(n11685), .A2(n11684), .ZN(n11686) );
  XNOR2_X1 U11306 ( .A(n14745), .B(n14747), .ZN(n14757) );
  NAND2_X1 U11307 ( .A1(n14751), .A2(n9935), .ZN(n14906) );
  OR2_X1 U11308 ( .A1(n14938), .A2(n14939), .ZN(n10241) );
  OR2_X1 U11309 ( .A1(n15005), .A2(n20745), .ZN(n15981) );
  AND2_X1 U11310 ( .A1(n15950), .A2(n10258), .ZN(n14926) );
  NAND2_X1 U11311 ( .A1(n15953), .A2(n11406), .ZN(n14938) );
  OR2_X1 U11312 ( .A1(n14780), .A2(n9981), .ZN(n9978) );
  OR2_X1 U11313 ( .A1(n15990), .A2(n14778), .ZN(n14780) );
  OR2_X1 U11314 ( .A1(n15992), .A2(n14820), .ZN(n15005) );
  OR2_X1 U11315 ( .A1(n14448), .A2(n19964), .ZN(n10067) );
  AOI21_X1 U11316 ( .B1(n14376), .B2(n14297), .A(n14280), .ZN(n14281) );
  OAI21_X1 U11317 ( .B1(n9976), .B2(n9975), .A(n9974), .ZN(n14836) );
  AND2_X1 U11318 ( .A1(n10791), .A2(n10790), .ZN(n14539) );
  OR2_X1 U11319 ( .A1(n10791), .A2(n10790), .ZN(n10173) );
  XNOR2_X1 U11320 ( .A(n11505), .B(n15066), .ZN(n15060) );
  NAND2_X1 U11321 ( .A1(n10245), .A2(n10243), .ZN(n16007) );
  AOI21_X1 U11322 ( .B1(n14166), .B2(n14165), .A(n14164), .ZN(n15652) );
  NAND2_X1 U11323 ( .A1(n14217), .A2(n10262), .ZN(n14303) );
  NOR2_X1 U11324 ( .A1(n14043), .A2(n14046), .ZN(n13738) );
  OR2_X1 U11325 ( .A1(n14076), .A2(n14086), .ZN(n14165) );
  INV_X1 U11326 ( .A(n15844), .ZN(n14874) );
  OR2_X1 U11327 ( .A1(n14076), .A2(n14077), .ZN(n14163) );
  NAND2_X1 U11328 ( .A1(n14563), .A2(n10751), .ZN(n10769) );
  NAND2_X1 U11329 ( .A1(n10212), .A2(n10214), .ZN(n14323) );
  NAND2_X1 U11330 ( .A1(n15676), .A2(n14201), .ZN(n15677) );
  XNOR2_X1 U11331 ( .A(n11507), .B(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n15041) );
  AND2_X1 U11332 ( .A1(n14557), .A2(n14558), .ZN(n14560) );
  OR2_X1 U11333 ( .A1(n11504), .A2(n11235), .ZN(n11507) );
  OR2_X1 U11334 ( .A1(n9961), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12922) );
  NOR2_X2 U11335 ( .A1(n14598), .A2(n14600), .ZN(n14599) );
  AOI21_X1 U11336 ( .B1(n14338), .B2(n14329), .A(n10004), .ZN(n10003) );
  OAI21_X1 U11337 ( .B1(n11477), .B2(n11307), .A(n12965), .ZN(n9961) );
  NAND2_X1 U11338 ( .A1(n14612), .A2(n14605), .ZN(n14598) );
  OR2_X1 U11339 ( .A1(n14648), .A2(n14641), .ZN(n14639) );
  NOR2_X1 U11340 ( .A1(n13376), .A2(n10063), .ZN(n10062) );
  NAND2_X1 U11341 ( .A1(n13245), .A2(n13244), .ZN(n13341) );
  NAND2_X1 U11342 ( .A1(n10219), .A2(n11195), .ZN(n11247) );
  NOR2_X1 U11343 ( .A1(n14688), .A2(n14698), .ZN(n14680) );
  XNOR2_X1 U11344 ( .A(n13339), .B(n13237), .ZN(n13245) );
  AND2_X1 U11345 ( .A1(n11294), .A2(n11293), .ZN(n11296) );
  AOI21_X1 U11346 ( .B1(n13360), .B2(n13505), .A(n13069), .ZN(n13096) );
  NAND2_X1 U11347 ( .A1(n13022), .A2(n13021), .ZN(n13236) );
  AND2_X1 U11348 ( .A1(n13380), .A2(n13063), .ZN(n13360) );
  XNOR2_X1 U11349 ( .A(n13380), .B(n13090), .ZN(n13369) );
  NAND2_X1 U11350 ( .A1(n10495), .A2(n10494), .ZN(n12216) );
  AND2_X1 U11351 ( .A1(n10470), .A2(n12231), .ZN(n12215) );
  NAND2_X1 U11352 ( .A1(n13059), .A2(n13060), .ZN(n13380) );
  INV_X1 U11353 ( .A(n19135), .ZN(n11218) );
  OR2_X1 U11354 ( .A1(n11985), .A2(n11983), .ZN(n10495) );
  CLKBUF_X1 U11355 ( .A(n11219), .Z(n13078) );
  CLKBUF_X1 U11356 ( .A(n13892), .Z(n14188) );
  INV_X1 U11357 ( .A(n12723), .ZN(n12743) );
  AND2_X1 U11358 ( .A1(n11136), .A2(n9963), .ZN(n19135) );
  INV_X1 U11359 ( .A(n19167), .ZN(n19170) );
  NAND2_X1 U11360 ( .A1(n11155), .A2(n11154), .ZN(n19420) );
  NAND2_X1 U11361 ( .A1(n10468), .A2(n10467), .ZN(n10497) );
  OR2_X1 U11362 ( .A1(n12236), .A2(n12237), .ZN(n12235) );
  NAND2_X1 U11363 ( .A1(n10479), .A2(n10478), .ZN(n10494) );
  NOR2_X1 U11364 ( .A1(n12668), .A2(n12866), .ZN(n12723) );
  OR2_X1 U11365 ( .A1(n20008), .A2(n13345), .ZN(n13020) );
  OR2_X2 U11366 ( .A1(n19938), .A2(n12916), .ZN(n15701) );
  AND2_X1 U11367 ( .A1(n12667), .A2(n12666), .ZN(n12866) );
  NAND2_X1 U11368 ( .A1(n11331), .A2(n10024), .ZN(n11364) );
  AOI221_X1 U11369 ( .B1(n18449), .B2(n18448), .C1(n18447), .C2(n18448), .A(
        n18446), .ZN(n18645) );
  NAND2_X1 U11370 ( .A1(n11418), .A2(n11333), .ZN(n11331) );
  XNOR2_X1 U11371 ( .A(n12804), .B(n20156), .ZN(n20269) );
  NAND2_X1 U11372 ( .A1(n10485), .A2(n10484), .ZN(n15077) );
  NAND2_X1 U11373 ( .A1(n17613), .A2(n15362), .ZN(n15364) );
  NOR2_X2 U11374 ( .A1(n12990), .A2(n19426), .ZN(n12991) );
  NAND2_X1 U11375 ( .A1(n18926), .A2(n11694), .ZN(n10485) );
  NAND2_X1 U11376 ( .A1(n10924), .A2(n10923), .ZN(n18948) );
  NAND2_X1 U11377 ( .A1(n12528), .A2(n12527), .ZN(n9917) );
  XNOR2_X1 U11378 ( .A(n11544), .B(n11545), .ZN(n11543) );
  NOR2_X1 U11379 ( .A1(n17605), .A2(n17604), .ZN(n17603) );
  NAND2_X1 U11380 ( .A1(n10454), .A2(n10453), .ZN(n11544) );
  NAND2_X1 U11381 ( .A1(n10441), .A2(n10440), .ZN(n10447) );
  NOR2_X1 U11382 ( .A1(n12460), .A2(n12462), .ZN(n12486) );
  NAND2_X1 U11383 ( .A1(n12653), .A2(n12652), .ZN(n20156) );
  OAI21_X1 U11384 ( .B1(n10455), .B2(n19067), .A(n10445), .ZN(n10446) );
  AND2_X1 U11385 ( .A1(n10083), .A2(n10082), .ZN(n17617) );
  XNOR2_X1 U11386 ( .A(n11853), .B(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n16219) );
  NAND2_X1 U11387 ( .A1(n11316), .A2(n11354), .ZN(n11418) );
  AND2_X1 U11388 ( .A1(n11311), .A2(n11309), .ZN(n11316) );
  NOR2_X2 U11389 ( .A1(n18654), .A2(n17293), .ZN(n17294) );
  NAND2_X1 U11390 ( .A1(n17639), .A2(n15358), .ZN(n15359) );
  AND2_X1 U11391 ( .A1(n10084), .A2(n9819), .ZN(n10082) );
  AND2_X1 U11392 ( .A1(n11301), .A2(n11300), .ZN(n11311) );
  AOI21_X1 U11393 ( .B1(n12425), .B2(n10057), .A(n10055), .ZN(n10054) );
  NAND2_X1 U11394 ( .A1(n12191), .A2(n9805), .ZN(n12537) );
  NAND2_X1 U11395 ( .A1(n10164), .A2(n10163), .ZN(n10917) );
  AND2_X1 U11396 ( .A1(n11520), .A2(n11525), .ZN(n10412) );
  AND2_X1 U11397 ( .A1(n12189), .A2(n12350), .ZN(n12191) );
  NAND2_X1 U11398 ( .A1(n10419), .A2(n10744), .ZN(n11548) );
  INV_X1 U11399 ( .A(n12909), .ZN(n12118) );
  AND2_X1 U11400 ( .A1(n15356), .A2(n17673), .ZN(n15352) );
  NOR4_X1 U11401 ( .A1(n18032), .A2(n18037), .A3(n11830), .A4(n15230), .ZN(
        n11829) );
  AND2_X1 U11402 ( .A1(n13951), .A2(n12909), .ZN(n12342) );
  NAND2_X2 U11403 ( .A1(n10930), .A2(n10925), .ZN(n11089) );
  AND2_X1 U11404 ( .A1(n10159), .A2(n11164), .ZN(n9966) );
  NAND2_X1 U11405 ( .A1(n20026), .A2(n20030), .ZN(n12780) );
  AND2_X1 U11406 ( .A1(n11526), .A2(n10909), .ZN(n11519) );
  CLKBUF_X1 U11407 ( .A(n10869), .Z(n11476) );
  AND2_X2 U11408 ( .A1(n10930), .A2(n11354), .ZN(n11071) );
  NAND2_X1 U11409 ( .A1(n12469), .A2(n13438), .ZN(n13936) );
  AND3_X1 U11410 ( .A1(n19085), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n10927), 
        .ZN(n10744) );
  INV_X2 U11411 ( .A(n10426), .ZN(n11354) );
  NAND4_X1 U11412 ( .A1(n12079), .A2(n12078), .A3(n12077), .A4(n12076), .ZN(
        n12119) );
  AND4_X2 U11413 ( .A1(n12116), .A2(n12115), .A3(n12114), .A4(n12113), .ZN(
        n20010) );
  NAND2_X1 U11414 ( .A1(n10071), .A2(n10070), .ZN(n17506) );
  NAND2_X1 U11415 ( .A1(n10329), .A2(n10328), .ZN(n19077) );
  NAND2_X2 U11416 ( .A1(n10222), .A2(n10221), .ZN(n19740) );
  AND4_X1 U11417 ( .A1(n12042), .A2(n12041), .A3(n12040), .A4(n12039), .ZN(
        n12058) );
  AND4_X1 U11418 ( .A1(n12066), .A2(n12065), .A3(n12064), .A4(n12063), .ZN(
        n12078) );
  AND4_X1 U11419 ( .A1(n12131), .A2(n12130), .A3(n12129), .A4(n12128), .ZN(
        n12142) );
  AND4_X1 U11420 ( .A1(n12112), .A2(n12111), .A3(n12110), .A4(n12109), .ZN(
        n12113) );
  AND4_X1 U11421 ( .A1(n12100), .A2(n12099), .A3(n12098), .A4(n12097), .ZN(
        n12116) );
  AND4_X1 U11422 ( .A1(n12135), .A2(n12134), .A3(n12133), .A4(n12132), .ZN(
        n12141) );
  NAND2_X1 U11423 ( .A1(n10381), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10221) );
  AND4_X1 U11424 ( .A1(n12104), .A2(n12103), .A3(n12102), .A4(n12101), .ZN(
        n12115) );
  AND4_X1 U11425 ( .A1(n12108), .A2(n12107), .A3(n12106), .A4(n12105), .ZN(
        n12114) );
  NOR2_X2 U11426 ( .A1(n20006), .A2(n20005), .ZN(n20007) );
  NAND2_X1 U11427 ( .A1(n10382), .A2(n10359), .ZN(n10222) );
  AND4_X1 U11428 ( .A1(n12071), .A2(n12070), .A3(n12069), .A4(n12068), .ZN(
        n12077) );
  AND4_X1 U11429 ( .A1(n12125), .A2(n12124), .A3(n12123), .A4(n12122), .ZN(
        n12143) );
  AND4_X1 U11430 ( .A1(n12062), .A2(n12061), .A3(n12060), .A4(n12059), .ZN(
        n12079) );
  AND4_X1 U11431 ( .A1(n12054), .A2(n12053), .A3(n12052), .A4(n12051), .ZN(
        n12055) );
  AND4_X1 U11432 ( .A1(n12050), .A2(n12049), .A3(n12048), .A4(n12047), .ZN(
        n12056) );
  NAND2_X1 U11433 ( .A1(n10315), .A2(n10359), .ZN(n10316) );
  NAND2_X1 U11434 ( .A1(n10266), .A2(n9792), .ZN(n10339) );
  NAND2_X2 U11435 ( .A1(n18665), .A2(n20947), .ZN(n18582) );
  AND2_X4 U11436 ( .A1(n9736), .A2(n10359), .ZN(n10522) );
  AND2_X4 U11437 ( .A1(n9736), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10576) );
  INV_X2 U11438 ( .A(n20005), .ZN(n9727) );
  AND4_X1 U11439 ( .A1(n12046), .A2(n12045), .A3(n12044), .A4(n12043), .ZN(
        n12057) );
  AND2_X1 U11440 ( .A1(n10344), .A2(n10343), .ZN(n9791) );
  AND3_X1 U11441 ( .A1(n10342), .A2(n10359), .A3(n10341), .ZN(n10345) );
  AND3_X1 U11442 ( .A1(n10348), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        n10347), .ZN(n10352) );
  AND2_X1 U11443 ( .A1(n10350), .A2(n10349), .ZN(n10351) );
  INV_X2 U11444 ( .A(n18956), .ZN(n19017) );
  BUF_X2 U11445 ( .A(n15264), .Z(n16991) );
  INV_X2 U11446 ( .A(n16371), .ZN(U215) );
  AND3_X1 U11447 ( .A1(n9958), .A2(n10359), .A3(n9957), .ZN(n10334) );
  BUF_X2 U11448 ( .A(n11788), .Z(n16777) );
  NAND2_X2 U11449 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(n19665), .ZN(n19669) );
  INV_X2 U11450 ( .A(n10673), .ZN(n10501) );
  INV_X4 U11451 ( .A(n10274), .ZN(n16974) );
  BUF_X2 U11452 ( .A(n12127), .Z(n9756) );
  BUF_X4 U11453 ( .A(n15151), .Z(n9729) );
  OR2_X1 U11454 ( .A1(n11736), .A2(n13568), .ZN(n9785) );
  INV_X4 U11455 ( .A(n9787), .ZN(n16968) );
  NAND2_X1 U11456 ( .A1(n9898), .A2(n9937), .ZN(n16990) );
  AND2_X2 U11457 ( .A1(n10509), .A2(n10674), .ZN(n10524) );
  AND2_X1 U11458 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n12690), .ZN(
        n10112) );
  AND2_X2 U11459 ( .A1(n13185), .A2(n10876), .ZN(n9753) );
  NAND2_X1 U11460 ( .A1(n18607), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11733) );
  NOR2_X2 U11461 ( .A1(n12778), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12781) );
  NAND2_X1 U11462 ( .A1(n18617), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11737) );
  NAND3_X2 U11463 ( .A1(n18667), .A2(n18596), .A3(n18666), .ZN(n17993) );
  AND2_X2 U11464 ( .A1(n12553), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12014) );
  OR2_X1 U11465 ( .A1(n18478), .A2(n13568), .ZN(n9787) );
  NAND2_X1 U11466 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n18630), .ZN(
        n11734) );
  AND2_X2 U11467 ( .A1(n11447), .A2(n10876), .ZN(n9735) );
  AND2_X1 U11468 ( .A1(n10507), .A2(n9955), .ZN(n9734) );
  INV_X2 U11469 ( .A(n10286), .ZN(n13188) );
  INV_X1 U11470 ( .A(n10376), .ZN(n9730) );
  AND2_X2 U11471 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14515) );
  AND2_X1 U11472 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12784) );
  NOR2_X1 U11473 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19685) );
  INV_X1 U11474 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n9955) );
  NOR2_X2 U11475 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10508) );
  NAND2_X1 U11476 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n18478) );
  NAND2_X1 U11477 ( .A1(n11149), .A2(n11986), .ZN(n11204) );
  AOI21_X1 U11478 ( .B1(n10241), .B2(n10236), .A(n14739), .ZN(n14745) );
  NAND4_X1 U11479 ( .A1(n10334), .A2(n10333), .A3(n10332), .A4(n10331), .ZN(
        n10340) );
  NOR2_X4 U11480 ( .A1(n11735), .A2(n16736), .ZN(n11754) );
  XNOR2_X1 U11481 ( .A(n9973), .B(n9788), .ZN(n11132) );
  NAND2_X1 U11482 ( .A1(n9971), .A2(n10437), .ZN(n9973) );
  INV_X1 U11483 ( .A(n10424), .ZN(n9965) );
  AND2_X1 U11484 ( .A1(n10509), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n9731) );
  AND2_X1 U11485 ( .A1(n10509), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n9745) );
  NAND2_X1 U11486 ( .A1(n10384), .A2(n10402), .ZN(n10415) );
  INV_X1 U11487 ( .A(n10402), .ZN(n10408) );
  NAND2_X1 U11488 ( .A1(n9887), .A2(n10383), .ZN(n10402) );
  NOR3_X2 U11489 ( .A1(n12900), .A2(n10192), .A3(n13230), .ZN(n13297) );
  INV_X2 U11490 ( .A(n11146), .ZN(n11119) );
  AND2_X1 U11491 ( .A1(n11109), .A2(n11146), .ZN(n11126) );
  AND2_X2 U11492 ( .A1(n14106), .A2(n13605), .ZN(n14097) );
  AND2_X1 U11493 ( .A1(n10507), .A2(n9955), .ZN(n9733) );
  XNOR2_X2 U11494 ( .A(n13234), .B(n20722), .ZN(n13022) );
  AND2_X2 U11495 ( .A1(n10435), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10452) );
  OR3_X2 U11496 ( .A1(n14938), .A2(n14939), .A3(n10269), .ZN(n10234) );
  AND2_X1 U11497 ( .A1(n11447), .A2(n10876), .ZN(n9736) );
  INV_X2 U11498 ( .A(n12618), .ZN(n9737) );
  INV_X2 U11499 ( .A(n9737), .ZN(n9738) );
  INV_X2 U11500 ( .A(n9737), .ZN(n9740) );
  AND2_X1 U11501 ( .A1(n12782), .A2(n10112), .ZN(n12618) );
  AND2_X4 U11502 ( .A1(n11538), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10456) );
  AND2_X2 U11503 ( .A1(n9956), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10510) );
  NAND2_X1 U11504 ( .A1(n10293), .A2(n10292), .ZN(n10389) );
  AND2_X1 U11505 ( .A1(n10480), .A2(n10483), .ZN(n18926) );
  NAND2_X1 U11506 ( .A1(n9959), .A2(n10418), .ZN(n10908) );
  NAND2_X2 U11507 ( .A1(n10246), .A2(n11232), .ZN(n11297) );
  NAND2_X1 U11508 ( .A1(n10210), .A2(n15645), .ZN(n14297) );
  INV_X2 U11509 ( .A(n10286), .ZN(n9743) );
  AND2_X1 U11510 ( .A1(n10509), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n9744) );
  BUF_X4 U11511 ( .A(n10346), .Z(n9746) );
  BUF_X4 U11512 ( .A(n10346), .Z(n9747) );
  BUF_X4 U11513 ( .A(n10346), .Z(n9748) );
  NOR2_X4 U11514 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13185) );
  OAI211_X2 U11515 ( .C1(n10432), .C2(n18954), .A(n10431), .B(n10430), .ZN(
        n10482) );
  OAI211_X2 U11516 ( .C1(n11522), .C2(n16176), .A(n10395), .B(n11530), .ZN(
        n10417) );
  AOI21_X2 U11517 ( .B1(n14722), .B2(n14719), .A(n14718), .ZN(n11439) );
  NAND2_X1 U11518 ( .A1(n11119), .A2(n11128), .ZN(n11284) );
  AND2_X1 U11519 ( .A1(n11119), .A2(n9886), .ZN(n11138) );
  AND2_X2 U11520 ( .A1(n13985), .A2(n10127), .ZN(n13974) );
  NOR2_X4 U11521 ( .A1(n13997), .A2(n13998), .ZN(n13985) );
  XNOR2_X1 U11522 ( .A(n12439), .B(n12438), .ZN(n12813) );
  AND2_X2 U11523 ( .A1(n13185), .A2(n10876), .ZN(n9752) );
  OAI21_X1 U11524 ( .B1(n9917), .B2(n12535), .A(n12804), .ZN(n12631) );
  NOR2_X1 U11525 ( .A1(n18654), .A2(n17293), .ZN(n9758) );
  INV_X4 U11526 ( .A(n18023), .ZN(n18654) );
  INV_X1 U11527 ( .A(n10385), .ZN(n9887) );
  NOR2_X1 U11528 ( .A1(n10927), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n10930) );
  AND2_X1 U11529 ( .A1(n18954), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n11694) );
  NAND2_X1 U11530 ( .A1(n11138), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n9885) );
  OAI21_X1 U11531 ( .B1(n11221), .B2(n11167), .A(n9962), .ZN(n11171) );
  NAND2_X1 U11532 ( .A1(n19135), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n9962) );
  NAND2_X1 U11533 ( .A1(n10426), .A2(n10418), .ZN(n10396) );
  NAND2_X1 U11534 ( .A1(n12723), .A2(n9765), .ZN(n13062) );
  INV_X1 U11535 ( .A(n9844), .ZN(n10001) );
  OAI21_X1 U11536 ( .B1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n9900), .A(
        n12003), .ZN(n12005) );
  AND2_X1 U11537 ( .A1(n11331), .A2(n10020), .ZN(n11374) );
  NOR2_X1 U11538 ( .A1(n10021), .A2(n11341), .ZN(n10020) );
  INV_X1 U11539 ( .A(n10022), .ZN(n10021) );
  NAND2_X1 U11540 ( .A1(n10007), .A2(n10006), .ZN(n10233) );
  NOR2_X1 U11541 ( .A1(n14923), .A2(n10237), .ZN(n10006) );
  INV_X1 U11542 ( .A(n14940), .ZN(n10237) );
  INV_X1 U11543 ( .A(n11233), .ZN(n11232) );
  INV_X1 U11544 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n9883) );
  NAND2_X1 U11545 ( .A1(n9825), .A2(n10116), .ZN(n10115) );
  INV_X1 U11546 ( .A(n14023), .ZN(n10116) );
  INV_X1 U11547 ( .A(n13096), .ZN(n10124) );
  INV_X1 U11548 ( .A(n13095), .ZN(n10125) );
  OR2_X1 U11549 ( .A1(n12539), .A2(n12396), .ZN(n13753) );
  INV_X1 U11550 ( .A(n13586), .ZN(n13505) );
  NAND2_X1 U11551 ( .A1(n14199), .A2(n14201), .ZN(n10213) );
  AND2_X1 U11552 ( .A1(n12191), .A2(n12190), .ZN(n12566) );
  INV_X1 U11553 ( .A(n13368), .ZN(n10063) );
  OR2_X1 U11554 ( .A1(n12373), .A2(n12372), .ZN(n13382) );
  OR2_X1 U11555 ( .A1(n12384), .A2(n12383), .ZN(n12907) );
  INV_X1 U11556 ( .A(n12665), .ZN(n13089) );
  INV_X1 U11557 ( .A(n12119), .ZN(n12187) );
  AND2_X1 U11558 ( .A1(n12120), .A2(n13437), .ZN(n12665) );
  NOR2_X1 U11559 ( .A1(n20010), .A2(n15822), .ZN(n12120) );
  AND2_X1 U11560 ( .A1(n12121), .A2(n13438), .ZN(n13377) );
  NAND2_X1 U11561 ( .A1(n11400), .A2(n11418), .ZN(n11398) );
  NOR2_X1 U11562 ( .A1(n16164), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10674) );
  INV_X1 U11563 ( .A(n10744), .ZN(n10788) );
  NAND2_X1 U11564 ( .A1(n10408), .A2(n10406), .ZN(n10163) );
  AND2_X1 U11565 ( .A1(n14859), .A2(n9831), .ZN(n10243) );
  INV_X1 U11566 ( .A(n16118), .ZN(n10156) );
  INV_X1 U11567 ( .A(n11506), .ZN(n9926) );
  AOI21_X1 U11568 ( .B1(n11506), .B2(n9925), .A(n9924), .ZN(n9922) );
  INV_X1 U11569 ( .A(n15059), .ZN(n9925) );
  INV_X1 U11570 ( .A(n15041), .ZN(n9924) );
  NOR2_X1 U11571 ( .A1(n11018), .A2(n11017), .ZN(n11242) );
  NAND2_X1 U11572 ( .A1(n9997), .A2(n9996), .ZN(n16837) );
  INV_X1 U11573 ( .A(n11735), .ZN(n9996) );
  INV_X1 U11574 ( .A(n11734), .ZN(n9997) );
  OR2_X1 U11575 ( .A1(n11733), .A2(n16736), .ZN(n9793) );
  OR2_X1 U11576 ( .A1(n15462), .A2(n12502), .ZN(n12506) );
  NOR2_X1 U11577 ( .A1(n14450), .A2(n9830), .ZN(n14412) );
  AND2_X1 U11578 ( .A1(n13422), .A2(n13421), .ZN(n13440) );
  NAND2_X1 U11579 ( .A1(n9913), .A2(n9912), .ZN(n13420) );
  NAND2_X1 U11580 ( .A1(n13417), .A2(n12564), .ZN(n9912) );
  AND2_X1 U11581 ( .A1(n12665), .A2(n13377), .ZN(n12173) );
  NOR2_X1 U11582 ( .A1(n14752), .A2(n11697), .ZN(n14734) );
  AND2_X1 U11584 ( .A1(n12301), .A2(n12298), .ZN(n12299) );
  NOR2_X1 U11585 ( .A1(n10498), .A2(n10183), .ZN(n10182) );
  INV_X1 U11586 ( .A(n10496), .ZN(n10183) );
  AND2_X1 U11587 ( .A1(n10497), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n10498) );
  INV_X1 U11588 ( .A(n11089), .ZN(n11516) );
  NAND2_X1 U11589 ( .A1(n15395), .A2(n9773), .ZN(n15411) );
  AND4_X1 U11590 ( .A1(n11042), .A2(n11041), .A3(n11040), .A4(n11039), .ZN(
        n11049) );
  AND4_X1 U11591 ( .A1(n11037), .A2(n11036), .A3(n11035), .A4(n11034), .ZN(
        n11050) );
  XNOR2_X1 U11592 ( .A(n11542), .B(n11543), .ZN(n10462) );
  AND2_X1 U11593 ( .A1(n11475), .A2(n18949), .ZN(n11668) );
  AOI21_X1 U11594 ( .B1(n15084), .B2(n11694), .A(n10489), .ZN(n12201) );
  XNOR2_X1 U11595 ( .A(n15077), .B(n10490), .ZN(n12202) );
  OR3_X1 U11596 ( .A1(n15462), .A2(n19757), .A3(n12340), .ZN(n13904) );
  OR3_X1 U11597 ( .A1(n15462), .A2(n19757), .A3(n15447), .ZN(n19764) );
  NOR2_X1 U11598 ( .A1(n16064), .A2(n15979), .ZN(n9987) );
  AND2_X1 U11599 ( .A1(n16064), .A2(n19706), .ZN(n19041) );
  OAI22_X1 U11600 ( .A1(n11185), .A2(n19340), .B1(n19420), .B2(n11184), .ZN(
        n11189) );
  OAI21_X1 U11601 ( .B1(n11214), .B2(n11178), .A(n9885), .ZN(n11183) );
  INV_X1 U11602 ( .A(n11211), .ZN(n11121) );
  AOI21_X1 U11603 ( .B1(n13464), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A(n9826), .ZN(n12714) );
  NAND2_X1 U11604 ( .A1(n19135), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n11140) );
  OAI22_X1 U11605 ( .A1(n11157), .A2(n19340), .B1(n19420), .B2(n11156), .ZN(
        n11158) );
  OAI211_X1 U11606 ( .C1(n11548), .C2(n13175), .A(n10434), .B(n10433), .ZN(
        n9970) );
  NAND2_X1 U11607 ( .A1(n10397), .A2(n10396), .ZN(n10902) );
  AND2_X1 U11608 ( .A1(n18926), .A2(n11110), .ZN(n11118) );
  CLKBUF_X1 U11609 ( .A(n13477), .Z(n13464) );
  AND2_X1 U11610 ( .A1(n12721), .A2(n12720), .ZN(n12742) );
  AOI21_X1 U11611 ( .B1(n13769), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .A(n9839), .ZN(n12411) );
  NOR2_X1 U11612 ( .A1(n12146), .A2(n12160), .ZN(n12166) );
  INV_X1 U11613 ( .A(n13086), .ZN(n12146) );
  NOR2_X1 U11614 ( .A1(n10023), .A2(n11338), .ZN(n10022) );
  INV_X1 U11615 ( .A(n10024), .ZN(n10023) );
  INV_X1 U11616 ( .A(n14589), .ZN(n10175) );
  INV_X1 U11617 ( .A(n10426), .ZN(n9959) );
  NAND2_X1 U11618 ( .A1(n10411), .A2(n10220), .ZN(n11520) );
  INV_X1 U11619 ( .A(n11118), .ZN(n11137) );
  NOR2_X1 U11620 ( .A1(n15330), .A2(n17181), .ZN(n15316) );
  NAND2_X1 U11621 ( .A1(n17187), .A2(n15356), .ZN(n15330) );
  NOR2_X1 U11622 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18630), .ZN(
        n13558) );
  INV_X1 U11623 ( .A(n14146), .ZN(n10117) );
  NAND2_X1 U11624 ( .A1(n9851), .A2(n10141), .ZN(n10140) );
  NOR2_X1 U11625 ( .A1(n10143), .A2(n10142), .ZN(n10141) );
  INV_X1 U11626 ( .A(n13508), .ZN(n10142) );
  NOR2_X1 U11627 ( .A1(n13511), .A2(n10144), .ZN(n10143) );
  INV_X1 U11628 ( .A(n13534), .ZN(n10144) );
  NAND2_X1 U11629 ( .A1(n10123), .A2(n10122), .ZN(n10126) );
  INV_X1 U11630 ( .A(n13094), .ZN(n10122) );
  AND2_X1 U11631 ( .A1(n9861), .A2(n10109), .ZN(n10108) );
  INV_X1 U11632 ( .A(n13999), .ZN(n10109) );
  NAND2_X1 U11633 ( .A1(n10106), .A2(n14081), .ZN(n10105) );
  INV_X1 U11634 ( .A(n14087), .ZN(n10106) );
  INV_X1 U11635 ( .A(n14323), .ZN(n14217) );
  INV_X1 U11636 ( .A(n15656), .ZN(n10004) );
  NAND2_X1 U11637 ( .A1(n9724), .A2(n9759), .ZN(n13948) );
  INV_X1 U11638 ( .A(n13144), .ZN(n10101) );
  INV_X1 U11639 ( .A(n13948), .ZN(n13940) );
  NAND2_X1 U11640 ( .A1(n13236), .A2(n13235), .ZN(n13339) );
  NAND2_X1 U11641 ( .A1(n12913), .A2(n12912), .ZN(n13011) );
  NAND2_X1 U11642 ( .A1(n10202), .A2(n10057), .ZN(n10056) );
  NOR2_X1 U11643 ( .A1(n12690), .A2(n15822), .ZN(n10057) );
  INV_X1 U11644 ( .A(n12633), .ZN(n13238) );
  AND2_X1 U11645 ( .A1(n12422), .A2(n12421), .ZN(n12637) );
  AND2_X1 U11646 ( .A1(n12419), .A2(n12418), .ZN(n12422) );
  NAND2_X1 U11647 ( .A1(n10111), .A2(n12403), .ZN(n12405) );
  NAND2_X1 U11648 ( .A1(n12425), .A2(n10201), .ZN(n10199) );
  AND2_X1 U11649 ( .A1(n20511), .A2(n12650), .ZN(n20270) );
  NOR2_X1 U11650 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n20009), .ZN(n20161) );
  NAND2_X1 U11651 ( .A1(n13089), .A2(n12167), .ZN(n9903) );
  NOR3_X1 U11652 ( .A1(n12170), .A2(n12169), .A3(n13089), .ZN(n12171) );
  AND2_X1 U11653 ( .A1(n12173), .A2(n12172), .ZN(n9901) );
  AOI21_X1 U11654 ( .B1(n10872), .B2(n10870), .A(n10867), .ZN(n10889) );
  INV_X1 U11655 ( .A(n10397), .ZN(n10393) );
  AND2_X1 U11656 ( .A1(n11414), .A2(n11436), .ZN(n11416) );
  NOR2_X1 U11657 ( .A1(n10018), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n10017) );
  NAND2_X1 U11658 ( .A1(n11347), .A2(n11346), .ZN(n11400) );
  NAND2_X1 U11659 ( .A1(n11331), .A2(n10022), .ZN(n11366) );
  NOR2_X1 U11660 ( .A1(n11321), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n11323) );
  NAND2_X1 U11661 ( .A1(n11318), .A2(n12245), .ZN(n11321) );
  INV_X1 U11662 ( .A(n10409), .ZN(n9931) );
  AOI21_X1 U11663 ( .B1(n9929), .B2(n15092), .A(n18954), .ZN(n9927) );
  NOR2_X1 U11664 ( .A1(n11538), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n9929) );
  NAND2_X1 U11665 ( .A1(n10439), .A2(n10438), .ZN(n10472) );
  INV_X1 U11666 ( .A(n9973), .ZN(n10486) );
  OR2_X1 U11667 ( .A1(n18788), .A2(n11235), .ZN(n11387) );
  AND2_X1 U11668 ( .A1(n10053), .A2(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n10051) );
  NOR2_X1 U11669 ( .A1(n16052), .A2(n10050), .ZN(n10053) );
  NAND2_X1 U11670 ( .A1(n11297), .A2(n11234), .ZN(n11492) );
  AND4_X1 U11671 ( .A1(n11046), .A2(n11045), .A3(n11044), .A4(n11043), .ZN(
        n11047) );
  AND2_X1 U11672 ( .A1(n11418), .A2(n14741), .ZN(n11436) );
  AOI21_X1 U11673 ( .B1(n10233), .B2(n10240), .A(n14748), .ZN(n10232) );
  INV_X1 U11674 ( .A(n9881), .ZN(n10235) );
  OR2_X1 U11675 ( .A1(n15905), .A2(n11235), .ZN(n11412) );
  NOR2_X1 U11676 ( .A1(n10148), .A2(n10147), .ZN(n10146) );
  INV_X1 U11677 ( .A(n13333), .ZN(n10147) );
  INV_X1 U11678 ( .A(n9982), .ZN(n9981) );
  NAND2_X1 U11679 ( .A1(n12893), .A2(n10193), .ZN(n10192) );
  NOR2_X1 U11680 ( .A1(n12899), .A2(n13041), .ZN(n10193) );
  NOR2_X1 U11681 ( .A1(n11059), .A2(n10158), .ZN(n10157) );
  INV_X1 U11682 ( .A(n12227), .ZN(n10158) );
  OR2_X1 U11683 ( .A1(n18821), .A2(n11235), .ZN(n11329) );
  NOR2_X1 U11684 ( .A1(n10189), .A2(n12243), .ZN(n10188) );
  INV_X1 U11685 ( .A(n12286), .ZN(n10189) );
  NAND2_X1 U11686 ( .A1(n11502), .A2(n11501), .ZN(n11505) );
  OR2_X1 U11687 ( .A1(n10861), .A2(n10860), .ZN(n11487) );
  OR2_X1 U11688 ( .A1(n10997), .A2(n10996), .ZN(n11240) );
  INV_X1 U11689 ( .A(n10415), .ZN(n10416) );
  NAND2_X1 U11690 ( .A1(n10476), .A2(n10475), .ZN(n10479) );
  AOI22_X1 U11691 ( .A1(n10672), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n9733), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10283) );
  AND2_X1 U11692 ( .A1(n10191), .A2(n10190), .ZN(n10281) );
  INV_X1 U11693 ( .A(n10279), .ZN(n10285) );
  NAND2_X1 U11694 ( .A1(n9951), .A2(n9950), .ZN(n11805) );
  INV_X1 U11695 ( .A(n18478), .ZN(n9950) );
  INV_X1 U11696 ( .A(n11733), .ZN(n9951) );
  INV_X1 U11697 ( .A(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n20912) );
  AND2_X1 U11698 ( .A1(n18630), .A2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n9937) );
  NAND2_X1 U11699 ( .A1(n11833), .A2(n15214), .ZN(n15202) );
  NOR2_X1 U11700 ( .A1(n16736), .A2(n11737), .ZN(n15264) );
  NOR2_X1 U11701 ( .A1(n17331), .A2(n15381), .ZN(n9895) );
  OR2_X1 U11702 ( .A1(n15380), .A2(n10268), .ZN(n15381) );
  INV_X1 U11703 ( .A(n16281), .ZN(n15338) );
  AND2_X1 U11704 ( .A1(n10261), .A2(n17907), .ZN(n10094) );
  NOR2_X1 U11705 ( .A1(n17594), .A2(n17902), .ZN(n15366) );
  NOR2_X1 U11706 ( .A1(n17603), .A2(n15336), .ZN(n15339) );
  AND2_X1 U11707 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n15335), .ZN(
        n15336) );
  XNOR2_X1 U11708 ( .A(n15316), .B(n17176), .ZN(n15333) );
  INV_X1 U11709 ( .A(n17628), .ZN(n10087) );
  NAND2_X1 U11710 ( .A1(n18459), .A2(n18458), .ZN(n15214) );
  OR2_X1 U11711 ( .A1(n13129), .A2(n19793), .ZN(n13251) );
  OR2_X1 U11712 ( .A1(n20664), .A2(n12835), .ZN(n15545) );
  INV_X1 U11713 ( .A(n19757), .ZN(n13421) );
  INV_X1 U11714 ( .A(n13753), .ZN(n13888) );
  NOR2_X1 U11715 ( .A1(n13975), .A2(n10128), .ZN(n10127) );
  INV_X1 U11716 ( .A(n13987), .ZN(n10128) );
  AND2_X1 U11717 ( .A1(n10130), .A2(n14156), .ZN(n10129) );
  AND2_X1 U11718 ( .A1(n13302), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n13444) );
  OR2_X1 U11719 ( .A1(n13095), .A2(n13096), .ZN(n13097) );
  AOI21_X1 U11720 ( .B1(n13350), .B2(n13505), .A(n12741), .ZN(n12755) );
  NAND2_X1 U11721 ( .A1(n12747), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12746) );
  NAND2_X1 U11722 ( .A1(n12688), .A2(n12647), .ZN(n12681) );
  AOI21_X1 U11723 ( .B1(n12645), .B2(n13586), .A(n10121), .ZN(n10120) );
  INV_X1 U11724 ( .A(n12647), .ZN(n10121) );
  INV_X1 U11725 ( .A(n15645), .ZN(n10209) );
  NOR2_X1 U11726 ( .A1(n10069), .A2(n9879), .ZN(n10068) );
  NAND2_X1 U11727 ( .A1(n13327), .A2(n13326), .ZN(n13536) );
  AOI21_X1 U11728 ( .B1(n10062), .B2(n10060), .A(n9807), .ZN(n10059) );
  INV_X1 U11729 ( .A(n13367), .ZN(n10060) );
  INV_X1 U11730 ( .A(n10062), .ZN(n10061) );
  INV_X1 U11731 ( .A(n19839), .ZN(n12761) );
  OAI21_X1 U11732 ( .B1(n20083), .B2(n13345), .A(n12471), .ZN(n12472) );
  NAND2_X1 U11733 ( .A1(n13440), .A2(n13433), .ZN(n19985) );
  OR2_X1 U11734 ( .A1(n9751), .A2(n20083), .ZN(n20434) );
  AND2_X1 U11735 ( .A1(n20330), .A2(n20161), .ZN(n20473) );
  NAND2_X1 U11736 ( .A1(n9751), .A2(n20400), .ZN(n20376) );
  OR2_X1 U11737 ( .A1(n11431), .A2(n11430), .ZN(n11434) );
  OR2_X1 U11738 ( .A1(n11422), .A2(n11421), .ZN(n15896) );
  INV_X1 U11739 ( .A(n11249), .ZN(n10011) );
  AND2_X1 U11740 ( .A1(n11250), .A2(n10012), .ZN(n11301) );
  AND3_X1 U11741 ( .A1(n10009), .A2(n11249), .A3(n10008), .ZN(n10012) );
  INV_X1 U11742 ( .A(n11243), .ZN(n10008) );
  XNOR2_X1 U11743 ( .A(n14599), .B(n10726), .ZN(n14590) );
  NAND2_X1 U11744 ( .A1(n12483), .A2(n11032), .ZN(n11968) );
  XNOR2_X1 U11745 ( .A(n11699), .B(n11698), .ZN(n12950) );
  OR2_X1 U11746 ( .A1(n14836), .A2(n14832), .ZN(n14777) );
  NOR2_X1 U11747 ( .A1(n15406), .A2(n18836), .ZN(n15400) );
  AND2_X1 U11748 ( .A1(n11573), .A2(n11572), .ZN(n12295) );
  NAND2_X1 U11749 ( .A1(n10257), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10254) );
  INV_X1 U11750 ( .A(n12824), .ZN(n10257) );
  OAI21_X1 U11751 ( .B1(n14751), .B2(n10249), .A(n12949), .ZN(n10248) );
  OR2_X1 U11752 ( .A1(n10251), .A2(n14717), .ZN(n10249) );
  AND2_X1 U11753 ( .A1(n14543), .A2(n14542), .ZN(n14545) );
  NOR2_X1 U11754 ( .A1(n10231), .A2(n10229), .ZN(n10228) );
  INV_X1 U11755 ( .A(n14845), .ZN(n10229) );
  OR2_X1 U11756 ( .A1(n11379), .A2(n14787), .ZN(n10231) );
  NOR2_X1 U11757 ( .A1(n14789), .A2(n14786), .ZN(n11396) );
  NAND2_X1 U11758 ( .A1(n13332), .A2(n13333), .ZN(n14707) );
  AND2_X1 U11759 ( .A1(n14624), .A2(n14623), .ZN(n14626) );
  NOR2_X1 U11760 ( .A1(n15418), .A2(n9983), .ZN(n9982) );
  INV_X1 U11761 ( .A(n14781), .ZN(n9983) );
  NAND2_X1 U11762 ( .A1(n14780), .A2(n9760), .ZN(n9984) );
  NAND2_X1 U11763 ( .A1(n13110), .A2(n13111), .ZN(n13290) );
  NAND2_X1 U11764 ( .A1(n16097), .A2(n15014), .ZN(n15015) );
  OR2_X1 U11765 ( .A1(n15025), .A2(n16122), .ZN(n16015) );
  AND2_X1 U11766 ( .A1(n11063), .A2(n11062), .ZN(n16118) );
  OR2_X1 U11767 ( .A1(n15025), .A2(n16134), .ZN(n16014) );
  AND2_X1 U11768 ( .A1(n11588), .A2(n11587), .ZN(n12304) );
  INV_X1 U11769 ( .A(n15027), .ZN(n10244) );
  NAND2_X1 U11770 ( .A1(n14819), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n15025) );
  NAND2_X1 U11771 ( .A1(n16044), .A2(n16045), .ZN(n9889) );
  NAND2_X1 U11772 ( .A1(n12921), .A2(n12924), .ZN(n9960) );
  AND2_X1 U11773 ( .A1(n10983), .A2(n10982), .ZN(n12251) );
  NAND2_X1 U11774 ( .A1(n10493), .A2(n10492), .ZN(n11983) );
  OR2_X1 U11775 ( .A1(n10497), .A2(n10469), .ZN(n10470) );
  NOR2_X1 U11776 ( .A1(n15084), .A2(n11127), .ZN(n11116) );
  AND2_X1 U11777 ( .A1(n15105), .A2(n18912), .ZN(n19225) );
  OR2_X1 U11778 ( .A1(n13215), .A2(n19710), .ZN(n19302) );
  INV_X1 U11779 ( .A(n19302), .ZN(n19338) );
  INV_X1 U11780 ( .A(n19686), .ZN(n19162) );
  NAND2_X1 U11781 ( .A1(n19690), .A2(n19716), .ZN(n19424) );
  AND2_X1 U11782 ( .A1(n13215), .A2(n19710), .ZN(n19553) );
  INV_X1 U11783 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n19744) );
  NAND2_X1 U11784 ( .A1(n16526), .A2(n10081), .ZN(n16507) );
  NAND2_X1 U11785 ( .A1(n9742), .A2(n17431), .ZN(n10081) );
  INV_X1 U11786 ( .A(n18046), .ZN(n17048) );
  NAND2_X1 U11787 ( .A1(n9726), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n10091) );
  AOI21_X1 U11788 ( .B1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B2(n16993), .A(n9942), .ZN(n9941) );
  INV_X1 U11789 ( .A(n15326), .ZN(n9942) );
  INV_X1 U11790 ( .A(n15324), .ZN(n9943) );
  NOR2_X1 U11791 ( .A1(n17544), .A2(n17534), .ZN(n10070) );
  INV_X1 U11792 ( .A(n17577), .ZN(n10071) );
  NAND2_X1 U11793 ( .A1(n17807), .A2(n9876), .ZN(n17346) );
  INV_X1 U11794 ( .A(n17465), .ZN(n15375) );
  AND2_X1 U11795 ( .A1(n15378), .A2(n17367), .ZN(n9896) );
  NAND3_X1 U11796 ( .A1(n15252), .A2(n15251), .A3(n15250), .ZN(n16273) );
  NOR2_X1 U11797 ( .A1(n15242), .A2(n15241), .ZN(n17919) );
  AND2_X1 U11798 ( .A1(n10088), .A2(n9954), .ZN(n17459) );
  AOI21_X1 U11799 ( .B1(n17802), .B2(n17585), .A(n17464), .ZN(n10088) );
  NAND2_X1 U11800 ( .A1(n17465), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n9954) );
  NAND2_X1 U11801 ( .A1(n17459), .A2(n17782), .ZN(n17458) );
  NOR2_X1 U11802 ( .A1(n18032), .A2(n18027), .ZN(n18453) );
  NAND2_X1 U11803 ( .A1(n17854), .A2(n17868), .ZN(n17848) );
  NOR2_X1 U11804 ( .A1(n17596), .A2(n17595), .ZN(n17594) );
  XNOR2_X1 U11805 ( .A(n15339), .B(n15340), .ZN(n17599) );
  NAND2_X1 U11806 ( .A1(n10087), .A2(n15332), .ZN(n10084) );
  OR2_X1 U11807 ( .A1(n17644), .A2(n10085), .ZN(n10083) );
  NAND2_X1 U11808 ( .A1(n10087), .A2(n10086), .ZN(n10085) );
  INV_X1 U11809 ( .A(n17643), .ZN(n10086) );
  NOR2_X1 U11810 ( .A1(n17644), .A2(n17643), .ZN(n17642) );
  XNOR2_X1 U11811 ( .A(n17199), .B(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n17665) );
  NAND2_X1 U11812 ( .A1(n18046), .A2(n18041), .ZN(n15230) );
  OR2_X1 U11813 ( .A1(n20578), .A2(n15822), .ZN(n19757) );
  NAND2_X1 U11814 ( .A1(n13903), .A2(n13904), .ZN(n20664) );
  NOR2_X1 U11815 ( .A1(n19885), .A2(n20667), .ZN(n15492) );
  NOR2_X1 U11816 ( .A1(n14409), .A2(n9915), .ZN(n14396) );
  NAND2_X1 U11817 ( .A1(n9916), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n9915) );
  NAND2_X1 U11818 ( .A1(n19988), .A2(n14221), .ZN(n9916) );
  NAND2_X1 U11819 ( .A1(n14460), .A2(n14380), .ZN(n14450) );
  INV_X1 U11820 ( .A(n14449), .ZN(n10065) );
  XNOR2_X1 U11821 ( .A(n14281), .B(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14448) );
  NAND2_X1 U11822 ( .A1(n9843), .A2(n9907), .ZN(n15702) );
  INV_X1 U11823 ( .A(n15711), .ZN(n9907) );
  NAND2_X1 U11824 ( .A1(n13440), .A2(n13426), .ZN(n15751) );
  NAND2_X1 U11825 ( .A1(n13440), .A2(n13425), .ZN(n19964) );
  AND2_X1 U11826 ( .A1(n9914), .A2(n12177), .ZN(n15462) );
  NAND2_X1 U11827 ( .A1(n12175), .A2(n12176), .ZN(n9914) );
  OR2_X1 U11828 ( .A1(n15866), .A2(n15838), .ZN(n10039) );
  NAND2_X1 U11829 ( .A1(n10033), .A2(n10034), .ZN(n10032) );
  NAND2_X1 U11830 ( .A1(n9769), .A2(n15838), .ZN(n10033) );
  INV_X1 U11831 ( .A(n10035), .ZN(n10034) );
  OR3_X1 U11832 ( .A1(n15866), .A2(n10038), .A3(n15838), .ZN(n10037) );
  NAND2_X1 U11833 ( .A1(n15867), .A2(n15868), .ZN(n15866) );
  OR2_X1 U11834 ( .A1(n15909), .A2(n15933), .ZN(n10027) );
  NAND2_X1 U11835 ( .A1(n10030), .A2(n10028), .ZN(n15890) );
  AOI21_X1 U11836 ( .B1(n18863), .B2(n15933), .A(n10029), .ZN(n10028) );
  INV_X1 U11837 ( .A(n15892), .ZN(n10029) );
  NAND2_X1 U11838 ( .A1(n15909), .A2(n18863), .ZN(n15901) );
  NAND2_X1 U11839 ( .A1(n15910), .A2(n15948), .ZN(n15909) );
  NAND2_X1 U11840 ( .A1(n12951), .A2(n10273), .ZN(n18736) );
  OR2_X1 U11841 ( .A1(n19735), .A2(n12959), .ZN(n18848) );
  INV_X1 U11842 ( .A(n18848), .ZN(n18918) );
  AND2_X1 U11843 ( .A1(n19024), .A2(n12954), .ZN(n18925) );
  OAI21_X1 U11844 ( .B1(n14874), .B2(n14602), .A(n11711), .ZN(n11712) );
  NAND2_X1 U11845 ( .A1(n10170), .A2(n10172), .ZN(n10168) );
  AND2_X1 U11846 ( .A1(n10565), .A2(n10588), .ZN(n10181) );
  AND2_X1 U11847 ( .A1(n12898), .A2(n12891), .ZN(n10588) );
  AND2_X1 U11848 ( .A1(n14621), .A2(n10390), .ZN(n14601) );
  NOR3_X1 U11849 ( .A1(n14648), .A2(n10160), .A3(n11514), .ZN(n11518) );
  INV_X1 U11850 ( .A(n15978), .ZN(n9988) );
  INV_X1 U11851 ( .A(n19035), .ZN(n16055) );
  NAND2_X1 U11852 ( .A1(n11867), .A2(n11693), .ZN(n16064) );
  AND2_X1 U11853 ( .A1(n11689), .A2(n10407), .ZN(n16060) );
  OR2_X1 U11854 ( .A1(n11691), .A2(n19056), .ZN(n11685) );
  AOI21_X1 U11855 ( .B1(n14908), .B2(n16154), .A(n14907), .ZN(n9934) );
  XNOR2_X1 U11856 ( .A(n14757), .B(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14909) );
  XNOR2_X1 U11857 ( .A(n15974), .B(n15973), .ZN(n16085) );
  INV_X1 U11858 ( .A(n19061), .ZN(n16154) );
  AND2_X1 U11859 ( .A1(n11668), .A2(n19724), .ZN(n16157) );
  AND2_X1 U11860 ( .A1(n11668), .A2(n19730), .ZN(n19065) );
  INV_X1 U11861 ( .A(n19707), .ZN(n19710) );
  INV_X1 U11862 ( .A(n16199), .ZN(n15104) );
  AND2_X1 U11863 ( .A1(n19225), .A2(n19162), .ZN(n19216) );
  INV_X1 U11864 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n19714) );
  AND2_X1 U11865 ( .A1(P3_EBX_REG_9__SCAN_IN), .A2(n17006), .ZN(n16982) );
  AND4_X1 U11866 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(P3_EBX_REG_5__SCAN_IN), 
        .A3(n17015), .A4(n16985), .ZN(n17006) );
  NAND2_X1 U11867 ( .A1(P3_EAX_REG_16__SCAN_IN), .A2(n17128), .ZN(n17124) );
  OR2_X1 U11868 ( .A1(n17691), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n9949) );
  NOR2_X1 U11869 ( .A1(n9946), .A2(n17928), .ZN(n9945) );
  NOR2_X1 U11870 ( .A1(n17696), .A2(n9947), .ZN(n9946) );
  NAND2_X1 U11871 ( .A1(n9948), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n9947) );
  NAND2_X1 U11872 ( .A1(n18469), .A2(n20821), .ZN(n9948) );
  AOI21_X1 U11873 ( .B1(n12658), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .A(
        n9871), .ZN(n13870) );
  AOI21_X1 U11874 ( .B1(n13477), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .A(n9870), .ZN(n13830) );
  AOI21_X1 U11875 ( .B1(n13477), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .A(n9869), .ZN(n13791) );
  AOI21_X1 U11876 ( .B1(n13769), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .A(n9856), .ZN(n13770) );
  AOI21_X1 U11877 ( .B1(n13477), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .A(n9857), .ZN(n13745) );
  INV_X1 U11878 ( .A(n12742), .ZN(n12722) );
  AOI21_X1 U11879 ( .B1(n13464), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .A(n9827), .ZN(n12729) );
  NOR2_X1 U11880 ( .A1(n20669), .A2(n20034), .ZN(n12344) );
  AOI21_X1 U11881 ( .B1(n13464), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .A(n9841), .ZN(n12659) );
  NAND2_X1 U11882 ( .A1(n12148), .A2(n9904), .ZN(n12149) );
  OR2_X1 U11883 ( .A1(n12096), .A2(n20010), .ZN(n9904) );
  AND2_X1 U11884 ( .A1(n9906), .A2(n9905), .ZN(n12148) );
  NAND2_X1 U11885 ( .A1(n12121), .A2(n12180), .ZN(n9905) );
  NAND2_X1 U11886 ( .A1(n9735), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n9958) );
  NAND2_X1 U11887 ( .A1(n9743), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n9957) );
  NAND2_X1 U11888 ( .A1(n10368), .A2(n10410), .ZN(n10369) );
  AOI21_X1 U11889 ( .B1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B2(n18013), .A(
        n11836), .ZN(n11837) );
  AOI21_X1 U11890 ( .B1(n13848), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .A(n9868), .ZN(n13696) );
  AOI21_X1 U11891 ( .B1(n13769), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .A(n9855), .ZN(n13498) );
  AOI21_X1 U11892 ( .B1(n13464), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A(n9859), .ZN(n13478) );
  AOI21_X1 U11893 ( .B1(n13769), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .A(n9853), .ZN(n13307) );
  AOI21_X1 U11894 ( .B1(n13464), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .A(n9858), .ZN(n13252) );
  NAND2_X1 U11895 ( .A1(n12723), .A2(n12722), .ZN(n12745) );
  INV_X1 U11896 ( .A(n12341), .ZN(n12188) );
  AOI21_X1 U11897 ( .B1(n13464), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .A(n9828), .ZN(n13051) );
  OR2_X1 U11898 ( .A1(n12719), .A2(n12718), .ZN(n13351) );
  NAND2_X1 U11899 ( .A1(n13848), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n12069) );
  NAND2_X1 U11900 ( .A1(n13867), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n12070) );
  NAND2_X1 U11901 ( .A1(n13843), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n12071) );
  AOI21_X1 U11902 ( .B1(n13769), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A(n9838), .ZN(n12379) );
  INV_X1 U11903 ( .A(n12348), .ZN(n10055) );
  AOI21_X1 U11904 ( .B1(n13464), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .A(n9840), .ZN(n12624) );
  NOR2_X1 U11905 ( .A1(n20047), .A2(n12339), .ZN(n9920) );
  NAND2_X1 U11906 ( .A1(n12780), .A2(n9918), .ZN(n12540) );
  NOR2_X1 U11907 ( .A1(n12553), .A2(n15822), .ZN(n10201) );
  NAND2_X1 U11908 ( .A1(n10202), .A2(n10201), .ZN(n10200) );
  AOI21_X1 U11909 ( .B1(n13477), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .A(
        n10198), .ZN(n12035) );
  AND2_X1 U11910 ( .A1(n12082), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n10198) );
  NOR2_X1 U11911 ( .A1(n10016), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n10015) );
  INV_X1 U11912 ( .A(n10017), .ZN(n10016) );
  AND2_X1 U11913 ( .A1(n11374), .A2(n11344), .ZN(n11369) );
  NOR2_X1 U11914 ( .A1(n10247), .A2(n10869), .ZN(n10409) );
  CLKBUF_X1 U11915 ( .A(n10672), .Z(n10844) );
  NAND2_X1 U11916 ( .A1(n10405), .A2(n10404), .ZN(n10435) );
  OR2_X1 U11917 ( .A1(n10978), .A2(n10977), .ZN(n11165) );
  NAND2_X1 U11918 ( .A1(n10400), .A2(n10399), .ZN(n11531) );
  NAND2_X1 U11919 ( .A1(n11666), .A2(n9968), .ZN(n9967) );
  INV_X1 U11920 ( .A(n9970), .ZN(n9969) );
  NOR2_X1 U11921 ( .A1(n9972), .A2(n18954), .ZN(n9968) );
  AND2_X1 U11922 ( .A1(n10908), .A2(n11164), .ZN(n10384) );
  AOI22_X1 U11923 ( .A1(n9743), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n9735), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10361) );
  AOI22_X1 U11924 ( .A1(n9743), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(n9735), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10355) );
  NOR2_X1 U11925 ( .A1(n11153), .A2(n11137), .ZN(n9886) );
  NOR2_X1 U11926 ( .A1(n11127), .A2(n11154), .ZN(n11128) );
  INV_X1 U11927 ( .A(n11127), .ZN(n11114) );
  NAND2_X1 U11928 ( .A1(n13188), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n10191) );
  NAND2_X1 U11929 ( .A1(n9735), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n10190) );
  INV_X1 U11930 ( .A(n10369), .ZN(n11468) );
  AND2_X1 U11931 ( .A1(n19722), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10880) );
  NOR2_X1 U11932 ( .A1(n15352), .A2(n17187), .ZN(n15350) );
  AOI21_X1 U11933 ( .B1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n18288), .A(
        n11835), .ZN(n11840) );
  AND2_X1 U11934 ( .A1(n11834), .A2(n13558), .ZN(n11835) );
  AND2_X1 U11935 ( .A1(n12550), .A2(n12501), .ZN(n12502) );
  NAND2_X1 U11936 ( .A1(n10114), .A2(n14012), .ZN(n10113) );
  INV_X1 U11937 ( .A(n10115), .ZN(n10114) );
  NOR2_X1 U11938 ( .A1(n13688), .A2(n10131), .ZN(n10130) );
  INV_X1 U11939 ( .A(n10132), .ZN(n10131) );
  OR2_X1 U11940 ( .A1(n14078), .A2(n14077), .ZN(n13688) );
  OR2_X1 U11941 ( .A1(n14166), .A2(n14086), .ZN(n14077) );
  NOR2_X1 U11942 ( .A1(n10134), .A2(n10133), .ZN(n10132) );
  INV_X1 U11943 ( .A(n14098), .ZN(n10134) );
  INV_X1 U11944 ( .A(n14091), .ZN(n10133) );
  AOI21_X1 U11945 ( .B1(n13769), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .A(n9854), .ZN(n13451) );
  OR2_X1 U11946 ( .A1(n13458), .A2(n13446), .ZN(n13513) );
  AOI21_X1 U11947 ( .B1(n13769), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A(n9852), .ZN(n13122) );
  NOR2_X1 U11948 ( .A1(n12746), .A2(n19822), .ZN(n12836) );
  NAND2_X1 U11949 ( .A1(n20042), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13586) );
  AND2_X1 U11950 ( .A1(n12395), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12677) );
  INV_X1 U11951 ( .A(n14007), .ZN(n10110) );
  NOR2_X1 U11952 ( .A1(n13536), .A2(n13535), .ZN(n10097) );
  INV_X1 U11953 ( .A(n13062), .ZN(n13059) );
  OAI21_X1 U11954 ( .B1(n15462), .B2(n13416), .A(n20026), .ZN(n9913) );
  NOR2_X1 U11955 ( .A1(n12390), .A2(n15822), .ZN(n13378) );
  OR2_X1 U11956 ( .A1(n12416), .A2(n12415), .ZN(n12908) );
  OAI21_X1 U11957 ( .B1(n10202), .B2(n12425), .A(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n12648) );
  NAND2_X1 U11958 ( .A1(n10216), .A2(n10217), .ZN(n12668) );
  AND2_X2 U11959 ( .A1(n12778), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12782) );
  INV_X1 U11960 ( .A(n12094), .ZN(n9999) );
  INV_X1 U11961 ( .A(n12095), .ZN(n10000) );
  OR3_X1 U11962 ( .A1(n12574), .A2(n12573), .A3(n12572), .ZN(n12806) );
  AOI21_X1 U11963 ( .B1(n15820), .B2(n15824), .A(n12811), .ZN(n20009) );
  NAND2_X1 U11964 ( .A1(n20010), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12632) );
  OR2_X1 U11965 ( .A1(n13437), .A2(n15822), .ZN(n12630) );
  AOI21_X1 U11966 ( .B1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n20368), .A(
        n11998), .ZN(n12007) );
  NOR2_X1 U11967 ( .A1(n11997), .A2(n12006), .ZN(n11998) );
  INV_X1 U11968 ( .A(n11165), .ZN(n11481) );
  AND2_X1 U11969 ( .A1(n11476), .A2(n11443), .ZN(n11237) );
  AND2_X1 U11970 ( .A1(n11398), .A2(n10013), .ZN(n11422) );
  NOR2_X1 U11971 ( .A1(n10014), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n10013) );
  INV_X1 U11972 ( .A(n10015), .ZN(n10014) );
  AND2_X1 U11973 ( .A1(n11369), .A2(n11345), .ZN(n11347) );
  NOR2_X1 U11974 ( .A1(n11361), .A2(n10025), .ZN(n10024) );
  NAND2_X1 U11975 ( .A1(n11418), .A2(n10005), .ZN(n11318) );
  NAND2_X1 U11976 ( .A1(n11250), .A2(n11249), .ZN(n11262) );
  INV_X1 U11977 ( .A(n10178), .ZN(n10750) );
  OAI211_X1 U11978 ( .C1(n14590), .C2(n10174), .A(n9863), .B(n10177), .ZN(
        n10178) );
  NAND2_X1 U11979 ( .A1(n10176), .A2(n10175), .ZN(n10174) );
  NOR2_X1 U11980 ( .A1(n11354), .A2(n10391), .ZN(n10159) );
  OR2_X1 U11981 ( .A1(n11031), .A2(n11030), .ZN(n11299) );
  NOR2_X1 U11982 ( .A1(n15940), .A2(n10048), .ZN(n10047) );
  AND2_X1 U11983 ( .A1(n10228), .A2(n9796), .ZN(n10227) );
  AND2_X1 U11984 ( .A1(n14585), .A2(n14587), .ZN(n14579) );
  AND2_X1 U11985 ( .A1(n14624), .A2(n10195), .ZN(n14593) );
  AND2_X1 U11986 ( .A1(n9832), .A2(n14606), .ZN(n10195) );
  NOR2_X1 U11987 ( .A1(n15409), .A2(n10045), .ZN(n10044) );
  NOR2_X1 U11988 ( .A1(n16021), .A2(n10042), .ZN(n10041) );
  INV_X1 U11989 ( .A(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n10042) );
  NAND2_X1 U11990 ( .A1(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n10250) );
  NAND2_X1 U11991 ( .A1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n10251) );
  AND2_X1 U11992 ( .A1(n10151), .A2(n10150), .ZN(n10149) );
  INV_X1 U11993 ( .A(n14664), .ZN(n10150) );
  NOR2_X1 U11994 ( .A1(n10259), .A2(n14930), .ZN(n10258) );
  INV_X1 U11995 ( .A(n10260), .ZN(n10259) );
  NOR2_X1 U11996 ( .A1(n14946), .A2(n15952), .ZN(n10260) );
  NOR2_X1 U11997 ( .A1(n10152), .A2(n14670), .ZN(n10151) );
  INV_X1 U11998 ( .A(n15916), .ZN(n10152) );
  AND2_X1 U11999 ( .A1(n11672), .A2(n10253), .ZN(n10252) );
  INV_X1 U12000 ( .A(n11675), .ZN(n10253) );
  OR2_X1 U12001 ( .A1(n18719), .A2(n11235), .ZN(n11382) );
  INV_X1 U12002 ( .A(n10461), .ZN(n11545) );
  OAI21_X1 U12003 ( .B1(n12927), .B2(n10455), .A(n10460), .ZN(n10461) );
  NAND2_X1 U12004 ( .A1(n10451), .A2(n10450), .ZN(n11542) );
  AND2_X1 U12005 ( .A1(n9800), .A2(n10948), .ZN(n10967) );
  NOR2_X1 U12006 ( .A1(n10960), .A2(n10959), .ZN(n11478) );
  NAND3_X1 U12007 ( .A1(n10393), .A2(n10428), .A3(n10392), .ZN(n10424) );
  NAND3_X1 U12008 ( .A1(n11119), .A2(n11109), .A3(n11154), .ZN(n11219) );
  INV_X1 U12009 ( .A(n11138), .ZN(n19098) );
  NOR2_X1 U12010 ( .A1(n11148), .A2(n11137), .ZN(n11120) );
  NAND2_X1 U12011 ( .A1(n9794), .A2(n11986), .ZN(n19453) );
  NAND3_X1 U12012 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n19685), .A3(n19549), 
        .ZN(n12979) );
  NAND2_X1 U12013 ( .A1(n9899), .A2(n9898), .ZN(n16767) );
  INV_X1 U12014 ( .A(n16736), .ZN(n9899) );
  NOR2_X1 U12015 ( .A1(n11734), .A2(n11733), .ZN(n15151) );
  INV_X1 U12016 ( .A(n17621), .ZN(n16679) );
  XNOR2_X1 U12017 ( .A(n17187), .B(n15356), .ZN(n15328) );
  NOR2_X1 U12018 ( .A1(n18448), .A2(n15217), .ZN(n15212) );
  OAI21_X1 U12019 ( .B1(n11845), .B2(n13560), .A(n13559), .ZN(n15233) );
  AND3_X1 U12020 ( .A1(n10000), .A2(n12117), .A3(n9999), .ZN(n12347) );
  NAND2_X1 U12021 ( .A1(n10264), .A2(n12118), .ZN(n12193) );
  AND2_X1 U12022 ( .A1(n12452), .A2(n12451), .ZN(n12453) );
  NOR2_X1 U12023 ( .A1(n14451), .A2(n13935), .ZN(n14454) );
  INV_X1 U12024 ( .A(n12772), .ZN(n19920) );
  AND2_X1 U12025 ( .A1(n12396), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n13887) );
  OR2_X1 U12026 ( .A1(n13858), .A2(n13989), .ZN(n13861) );
  NAND2_X1 U12027 ( .A1(n13820), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n13858) );
  NOR2_X1 U12028 ( .A1(n13779), .A2(n13777), .ZN(n13782) );
  OAI21_X1 U12029 ( .B1(n13886), .B2(n14275), .A(n13800), .ZN(n14023) );
  OR2_X1 U12030 ( .A1(n13761), .A2(n13760), .ZN(n14146) );
  AND2_X1 U12031 ( .A1(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n13734), .ZN(
        n13756) );
  NOR2_X1 U12032 ( .A1(n13655), .A2(n12840), .ZN(n13689) );
  NAND2_X1 U12033 ( .A1(n13654), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n13655) );
  AND2_X1 U12034 ( .A1(n14097), .A2(n14098), .ZN(n14100) );
  NOR2_X1 U12035 ( .A1(n13572), .A2(n12838), .ZN(n13589) );
  NAND2_X1 U12036 ( .A1(n13589), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n13616) );
  NAND2_X1 U12037 ( .A1(n10137), .A2(n10136), .ZN(n10135) );
  INV_X1 U12038 ( .A(n14114), .ZN(n10136) );
  INV_X1 U12039 ( .A(n10140), .ZN(n10137) );
  AND2_X1 U12040 ( .A1(n13459), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n13493) );
  NAND2_X1 U12041 ( .A1(n9851), .A2(n10139), .ZN(n10138) );
  INV_X1 U12042 ( .A(n10143), .ZN(n10139) );
  NOR2_X1 U12043 ( .A1(n13251), .A2(n12837), .ZN(n13302) );
  INV_X1 U12044 ( .A(n10126), .ZN(n13098) );
  NOR2_X1 U12045 ( .A1(n13097), .A2(n13098), .ZN(n13133) );
  AND2_X1 U12046 ( .A1(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n12836), .ZN(
        n13091) );
  INV_X1 U12047 ( .A(n12755), .ZN(n12754) );
  NOR2_X1 U12048 ( .A1(n12671), .A2(n12670), .ZN(n12747) );
  INV_X1 U12049 ( .A(n12685), .ZN(n12646) );
  NAND2_X1 U12050 ( .A1(n14262), .A2(n9921), .ZN(n14232) );
  NOR2_X1 U12051 ( .A1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n9921) );
  NAND2_X1 U12052 ( .A1(n14039), .A2(n9861), .ZN(n14009) );
  NOR2_X1 U12053 ( .A1(n14430), .A2(n14438), .ZN(n10002) );
  AND3_X1 U12054 ( .A1(n10210), .A2(n15645), .A3(n10206), .ZN(n14262) );
  INV_X1 U12055 ( .A(n10207), .ZN(n10206) );
  OAI21_X1 U12056 ( .B1(n9750), .B2(n14438), .A(n10208), .ZN(n10207) );
  INV_X1 U12057 ( .A(n14219), .ZN(n10208) );
  AND2_X1 U12058 ( .A1(n14454), .A2(n14037), .ZN(n14039) );
  NAND2_X1 U12059 ( .A1(n14039), .A2(n14019), .ZN(n14021) );
  NAND2_X1 U12060 ( .A1(n10104), .A2(n10103), .ZN(n10102) );
  NOR2_X1 U12061 ( .A1(n9874), .A2(n15526), .ZN(n10103) );
  INV_X1 U12062 ( .A(n10105), .ZN(n10104) );
  NOR3_X1 U12063 ( .A1(n14095), .A2(n9874), .A3(n14087), .ZN(n15502) );
  NOR2_X1 U12064 ( .A1(n14095), .A2(n14087), .ZN(n15501) );
  INV_X1 U12065 ( .A(n14215), .ZN(n10215) );
  NOR2_X1 U12066 ( .A1(n14118), .A2(n14110), .ZN(n14109) );
  AND2_X1 U12067 ( .A1(n13909), .A2(n13908), .ZN(n14115) );
  OR2_X1 U12068 ( .A1(n14116), .A2(n14115), .ZN(n14118) );
  AND2_X1 U12069 ( .A1(n14461), .A2(n14385), .ZN(n15726) );
  OR2_X1 U12070 ( .A1(n9749), .A2(n15744), .ZN(n14341) );
  NAND2_X1 U12071 ( .A1(n14058), .A2(n13531), .ZN(n14116) );
  NOR2_X1 U12072 ( .A1(n14503), .A2(n14059), .ZN(n14058) );
  NAND2_X1 U12073 ( .A1(n10097), .A2(n10096), .ZN(n14503) );
  INV_X1 U12074 ( .A(n14500), .ZN(n10096) );
  INV_X1 U12075 ( .A(n10097), .ZN(n14501) );
  AND2_X1 U12076 ( .A1(n15789), .A2(n9846), .ZN(n13327) );
  NAND2_X1 U12077 ( .A1(n15789), .A2(n9761), .ZN(n13145) );
  AND2_X1 U12078 ( .A1(n13101), .A2(n13100), .ZN(n15788) );
  NAND2_X1 U12079 ( .A1(n12761), .A2(n10272), .ZN(n19842) );
  NAND2_X1 U12080 ( .A1(n12392), .A2(n12391), .ZN(n12403) );
  AND3_X1 U12081 ( .A1(n12390), .A2(n12389), .A3(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n12391) );
  NAND2_X1 U12082 ( .A1(n12432), .A2(n12431), .ZN(n20055) );
  OR2_X1 U12083 ( .A1(n20008), .A2(n12867), .ZN(n20239) );
  INV_X1 U12084 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20368) );
  OR2_X1 U12085 ( .A1(n12864), .A2(n12865), .ZN(n20377) );
  INV_X1 U12086 ( .A(n20083), .ZN(n20400) );
  INV_X1 U12087 ( .A(n12121), .ZN(n20038) );
  INV_X2 U12088 ( .A(n9919), .ZN(n20042) );
  AOI21_X1 U12089 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n20435), .A(n20057), 
        .ZN(n20523) );
  OR3_X1 U12090 ( .A1(n20275), .A2(P1_STATE2_REG_0__SCAN_IN), .A3(n20009), 
        .ZN(n20048) );
  NAND2_X1 U12091 ( .A1(n12632), .A2(n12630), .ZN(n13086) );
  AOI21_X1 U12092 ( .B1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n15822), .A(
        n12174), .ZN(n12175) );
  NAND2_X1 U12093 ( .A1(n9902), .A2(n9801), .ZN(n12174) );
  OAI21_X1 U12094 ( .B1(n12164), .B2(n9837), .A(n9903), .ZN(n9902) );
  INV_X1 U12095 ( .A(n13438), .ZN(n12180) );
  AOI21_X1 U12096 ( .B1(n10892), .B2(n10891), .A(n10890), .ZN(n11459) );
  AND2_X1 U12097 ( .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n15508), .ZN(
        n10890) );
  OAI21_X1 U12098 ( .B1(n18863), .B2(n10038), .A(n10036), .ZN(n10035) );
  INV_X1 U12099 ( .A(n15846), .ZN(n10038) );
  NAND2_X1 U12100 ( .A1(n11424), .A2(n14740), .ZN(n14744) );
  NAND2_X1 U12101 ( .A1(n11398), .A2(n10017), .ZN(n11410) );
  AND2_X1 U12102 ( .A1(n15395), .A2(n10043), .ZN(n15410) );
  AND2_X1 U12103 ( .A1(n9773), .A2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n10043) );
  AND2_X1 U12104 ( .A1(n11353), .A2(n11373), .ZN(n18744) );
  AND2_X1 U12105 ( .A1(n11368), .A2(n11367), .ZN(n18753) );
  AND2_X1 U12106 ( .A1(n12986), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n11361) );
  NAND2_X1 U12107 ( .A1(n11323), .A2(n18809), .ZN(n11333) );
  NAND2_X1 U12108 ( .A1(n11331), .A2(n11332), .ZN(n11362) );
  AND2_X1 U12109 ( .A1(n11970), .A2(n11051), .ZN(n11991) );
  AND2_X1 U12110 ( .A1(n11053), .A2(n11052), .ZN(n11990) );
  INV_X1 U12111 ( .A(n15092), .ZN(n9930) );
  AND2_X1 U12112 ( .A1(n14560), .A2(n14551), .ZN(n14543) );
  AND2_X1 U12113 ( .A1(n11056), .A2(n12241), .ZN(n12298) );
  NAND2_X1 U12114 ( .A1(n10162), .A2(n10161), .ZN(n10160) );
  INV_X1 U12115 ( .A(n14633), .ZN(n10161) );
  INV_X1 U12116 ( .A(n14641), .ZN(n10162) );
  INV_X1 U12117 ( .A(n10851), .ZN(n10172) );
  NOR2_X1 U12118 ( .A1(n10829), .A2(n10851), .ZN(n10169) );
  NAND2_X1 U12119 ( .A1(n13332), .A2(n9775), .ZN(n14698) );
  AND2_X1 U12120 ( .A1(n9774), .A2(n10185), .ZN(n10184) );
  INV_X1 U12121 ( .A(n14614), .ZN(n10185) );
  NAND2_X1 U12122 ( .A1(n13289), .A2(n9774), .ZN(n14613) );
  OR2_X1 U12123 ( .A1(n10630), .A2(n10629), .ZN(n13330) );
  NAND2_X1 U12124 ( .A1(n13289), .A2(n9771), .ZN(n13391) );
  NOR2_X1 U12125 ( .A1(n11991), .A2(n11990), .ZN(n11989) );
  OAI21_X1 U12126 ( .B1(n11104), .B2(n11103), .A(P2_ADDRESS_REG_29__SCAN_IN), 
        .ZN(n11897) );
  INV_X1 U12127 ( .A(n11897), .ZN(n12980) );
  NAND2_X1 U12128 ( .A1(n14758), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14752) );
  AND2_X1 U12129 ( .A1(n15835), .A2(n10046), .ZN(n14758) );
  AND2_X1 U12130 ( .A1(n9777), .A2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n10046) );
  NAND2_X1 U12131 ( .A1(n15835), .A2(n9777), .ZN(n14768) );
  AND2_X1 U12132 ( .A1(n14580), .A2(n14566), .ZN(n14557) );
  NAND2_X1 U12133 ( .A1(n15835), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15836) );
  AND2_X1 U12134 ( .A1(n14579), .A2(n14578), .ZN(n14580) );
  NOR2_X1 U12135 ( .A1(n15834), .A2(n15959), .ZN(n15835) );
  NAND2_X1 U12136 ( .A1(n10226), .A2(n10225), .ZN(n15955) );
  OAI21_X1 U12137 ( .B1(n10224), .B2(n11397), .A(n9796), .ZN(n10225) );
  NAND2_X1 U12138 ( .A1(n10230), .A2(n10227), .ZN(n10226) );
  INV_X1 U12139 ( .A(n14953), .ZN(n10224) );
  NAND2_X1 U12140 ( .A1(n15410), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n14808) );
  NOR2_X1 U12141 ( .A1(n14808), .A2(n18695), .ZN(n15394) );
  AND2_X1 U12142 ( .A1(n14624), .A2(n9832), .ZN(n14619) );
  NAND2_X1 U12143 ( .A1(n15395), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15408) );
  NOR2_X1 U12144 ( .A1(n15396), .A2(n15996), .ZN(n15395) );
  NAND2_X1 U12145 ( .A1(n15397), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n15396) );
  AND2_X1 U12146 ( .A1(n15400), .A2(n10040), .ZN(n15397) );
  AND2_X1 U12147 ( .A1(n9772), .A2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n10040) );
  AND2_X1 U12148 ( .A1(n11605), .A2(n11604), .ZN(n12899) );
  NAND2_X1 U12149 ( .A1(n15400), .A2(n9772), .ZN(n15398) );
  NAND2_X1 U12150 ( .A1(n15400), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n15399) );
  NAND2_X1 U12151 ( .A1(n9813), .A2(n10052), .ZN(n15406) );
  AND2_X1 U12152 ( .A1(n10052), .A2(n10051), .ZN(n15407) );
  NAND2_X1 U12153 ( .A1(n10052), .A2(n10053), .ZN(n15404) );
  NOR2_X1 U12154 ( .A1(n15402), .A2(n16052), .ZN(n15405) );
  INV_X1 U12155 ( .A(n11492), .ZN(n11491) );
  INV_X1 U12156 ( .A(n12822), .ZN(n9888) );
  NOR2_X1 U12157 ( .A1(n11957), .A2(n16065), .ZN(n15403) );
  OR2_X1 U12158 ( .A1(n10941), .A2(n10940), .ZN(n11923) );
  INV_X1 U12159 ( .A(n14739), .ZN(n10239) );
  NAND2_X1 U12160 ( .A1(n10234), .A2(n10232), .ZN(n9884) );
  OR2_X1 U12161 ( .A1(n14658), .A2(n14650), .ZN(n14648) );
  OAI21_X1 U12162 ( .B1(n11417), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n11426), .ZN(n14765) );
  NAND2_X1 U12163 ( .A1(n10241), .A2(n14940), .ZN(n14925) );
  NAND2_X1 U12164 ( .A1(n15950), .A2(n10260), .ZN(n14937) );
  NAND2_X1 U12165 ( .A1(n14679), .A2(n10151), .ZN(n14672) );
  NAND2_X1 U12166 ( .A1(n14679), .A2(n15916), .ZN(n15915) );
  AND2_X1 U12167 ( .A1(n14624), .A2(n9829), .ZN(n14616) );
  NAND2_X1 U12168 ( .A1(n13332), .A2(n10146), .ZN(n14705) );
  AND2_X1 U12169 ( .A1(n13297), .A2(n13298), .ZN(n14624) );
  INV_X1 U12170 ( .A(n9980), .ZN(n9979) );
  OAI21_X1 U12171 ( .B1(n9760), .B2(n9981), .A(n14785), .ZN(n9980) );
  NOR2_X1 U12172 ( .A1(n13290), .A2(n13291), .ZN(n13332) );
  NOR2_X1 U12173 ( .A1(n15015), .A2(n11074), .ZN(n13110) );
  AOI21_X1 U12174 ( .B1(n14776), .B2(n9977), .A(n15997), .ZN(n9974) );
  INV_X1 U12175 ( .A(n14776), .ZN(n9975) );
  NAND2_X1 U12176 ( .A1(n16010), .A2(n14845), .ZN(n9977) );
  AND2_X1 U12177 ( .A1(n11067), .A2(n11066), .ZN(n16099) );
  AND2_X1 U12178 ( .A1(n11597), .A2(n11596), .ZN(n12515) );
  OR2_X1 U12179 ( .A1(n12514), .A2(n12515), .ZN(n12900) );
  NOR2_X1 U12180 ( .A1(n9824), .A2(n10155), .ZN(n10154) );
  INV_X1 U12181 ( .A(n12261), .ZN(n10155) );
  NOR2_X1 U12182 ( .A1(n15031), .A2(n9824), .ZN(n16116) );
  AND2_X1 U12183 ( .A1(n12293), .A2(n9817), .ZN(n12496) );
  INV_X1 U12184 ( .A(n12304), .ZN(n10187) );
  NOR2_X1 U12185 ( .A1(n15031), .A2(n11059), .ZN(n15033) );
  NAND2_X1 U12186 ( .A1(n10153), .A2(n10157), .ZN(n16117) );
  OR2_X1 U12187 ( .A1(n11504), .A2(n11509), .ZN(n11510) );
  NAND2_X1 U12188 ( .A1(n12293), .A2(n10188), .ZN(n12303) );
  NOR2_X1 U12189 ( .A1(n12294), .A2(n12295), .ZN(n12293) );
  NAND2_X1 U12190 ( .A1(n12293), .A2(n12286), .ZN(n12287) );
  CLKBUF_X1 U12191 ( .A(n15042), .Z(n15043) );
  OR2_X1 U12192 ( .A1(n12235), .A2(n12264), .ZN(n12275) );
  AND2_X1 U12193 ( .A1(n11567), .A2(n11566), .ZN(n12276) );
  OR2_X1 U12194 ( .A1(n12275), .A2(n12276), .ZN(n12294) );
  AND2_X1 U12195 ( .A1(n12487), .A2(n12482), .ZN(n10145) );
  NAND2_X1 U12196 ( .A1(n9891), .A2(n11488), .ZN(n11489) );
  NAND2_X1 U12197 ( .A1(n12486), .A2(n12487), .ZN(n12488) );
  AND2_X1 U12198 ( .A1(n11554), .A2(n11553), .ZN(n12237) );
  NAND2_X1 U12199 ( .A1(n19047), .A2(n19048), .ZN(n14998) );
  NAND2_X1 U12200 ( .A1(n12253), .A2(n10987), .ZN(n12460) );
  AND2_X1 U12201 ( .A1(n11005), .A2(n11004), .ZN(n12462) );
  INV_X1 U12202 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n9956) );
  CLKBUF_X1 U12203 ( .A(n10436), .Z(n15091) );
  INV_X1 U12204 ( .A(n19607), .ZN(n18949) );
  AND2_X1 U12205 ( .A1(n15105), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19226) );
  NOR2_X1 U12206 ( .A1(n11154), .A2(n11135), .ZN(n9963) );
  NAND2_X1 U12207 ( .A1(n15105), .A2(n19716), .ZN(n19199) );
  INV_X1 U12208 ( .A(n19423), .ZN(n19459) );
  OAI21_X1 U12209 ( .B1(n10285), .B2(n10284), .A(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10293) );
  NOR2_X1 U12210 ( .A1(n12980), .A2(n12979), .ZN(n19089) );
  NOR2_X1 U12211 ( .A1(n14634), .A2(n12979), .ZN(n19090) );
  INV_X1 U12212 ( .A(n19089), .ZN(n19079) );
  INV_X1 U12213 ( .A(n19090), .ZN(n19080) );
  INV_X1 U12214 ( .A(n19084), .ZN(n19076) );
  INV_X1 U12215 ( .A(n16167), .ZN(n11861) );
  NOR2_X1 U12216 ( .A1(n15220), .A2(n15202), .ZN(n18442) );
  NOR2_X1 U12217 ( .A1(n16445), .A2(n16444), .ZN(n16443) );
  NOR2_X1 U12218 ( .A1(n17344), .A2(n16464), .ZN(n16463) );
  NOR2_X1 U12219 ( .A1(P3_EBX_REG_19__SCAN_IN), .A2(n16529), .ZN(n16520) );
  AND2_X1 U12220 ( .A1(n16888), .A2(n9990), .ZN(n16835) );
  AND2_X1 U12221 ( .A1(n9784), .A2(P3_EBX_REG_20__SCAN_IN), .ZN(n9990) );
  NOR2_X1 U12222 ( .A1(n11743), .A2(n11742), .ZN(n16694) );
  OR2_X1 U12223 ( .A1(n13565), .A2(n15212), .ZN(n9994) );
  NOR3_X1 U12224 ( .A1(n13556), .A2(n18037), .A3(n18052), .ZN(n13565) );
  AND3_X1 U12225 ( .A1(n18443), .A2(n18655), .A3(n15202), .ZN(n15511) );
  NOR3_X1 U12226 ( .A1(n17200), .A2(n18652), .A3(n17238), .ZN(n17218) );
  NAND2_X1 U12227 ( .A1(n17333), .A2(n9770), .ZN(n16253) );
  AND2_X1 U12228 ( .A1(n17333), .A2(n9776), .ZN(n16252) );
  NOR2_X1 U12229 ( .A1(n17314), .A2(n10073), .ZN(n10072) );
  NAND2_X1 U12230 ( .A1(n17321), .A2(n17585), .ZN(n9894) );
  NAND2_X1 U12231 ( .A1(n17333), .A2(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n17313) );
  NOR2_X1 U12232 ( .A1(n17352), .A2(n17353), .ZN(n17333) );
  NAND2_X1 U12233 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n17376), .ZN(
        n17352) );
  NOR2_X1 U12234 ( .A1(n17467), .A2(n17473), .ZN(n17453) );
  NAND2_X1 U12235 ( .A1(n17584), .A2(n15373), .ZN(n17480) );
  OR2_X1 U12236 ( .A1(n17509), .A2(n17498), .ZN(n17472) );
  OR2_X1 U12237 ( .A1(n17506), .A2(n17472), .ZN(n17467) );
  INV_X1 U12238 ( .A(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n17534) );
  NAND4_X1 U12239 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A4(
        P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n17544) );
  OR2_X1 U12240 ( .A1(n17533), .A2(n20957), .ZN(n17577) );
  NAND2_X1 U12241 ( .A1(n16679), .A2(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n17533) );
  AND2_X1 U12242 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17631) );
  AOI22_X1 U12243 ( .A1(n16207), .A2(n18447), .B1(n18445), .B2(n17919), .ZN(
        n16218) );
  NOR2_X1 U12244 ( .A1(n15479), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16209) );
  NAND2_X1 U12245 ( .A1(n16282), .A2(n10092), .ZN(n15479) );
  INV_X1 U12246 ( .A(n16272), .ZN(n10092) );
  NOR2_X1 U12247 ( .A1(n17345), .A2(n17679), .ZN(n17686) );
  NOR2_X1 U12248 ( .A1(n17346), .A2(n20821), .ZN(n17690) );
  OR2_X1 U12249 ( .A1(n17367), .A2(n17715), .ZN(n17345) );
  NAND2_X1 U12250 ( .A1(n17807), .A2(n17366), .ZN(n17716) );
  OR2_X1 U12251 ( .A1(n17778), .A2(n17465), .ZN(n17403) );
  NOR2_X1 U12252 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17585), .ZN(
        n17447) );
  INV_X1 U12253 ( .A(n9952), .ZN(n17464) );
  OAI21_X1 U12254 ( .B1(n15373), .B2(n9953), .A(n17551), .ZN(n9952) );
  NOR2_X1 U12255 ( .A1(n17848), .A2(n17517), .ZN(n17495) );
  NAND2_X1 U12256 ( .A1(n15371), .A2(n17575), .ZN(n17868) );
  INV_X1 U12257 ( .A(n15373), .ZN(n17552) );
  INV_X1 U12258 ( .A(n10095), .ZN(n17874) );
  NAND2_X1 U12259 ( .A1(n17607), .A2(n15365), .ZN(n17595) );
  XNOR2_X1 U12260 ( .A(n15364), .B(n9939), .ZN(n17608) );
  INV_X1 U12261 ( .A(n15363), .ZN(n9939) );
  NAND2_X1 U12262 ( .A1(n17608), .A2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n17607) );
  NAND2_X1 U12263 ( .A1(n9892), .A2(n17616), .ZN(n17605) );
  OAI21_X1 U12264 ( .B1(n17617), .B2(n17618), .A(n17936), .ZN(n9892) );
  NAND2_X1 U12265 ( .A1(n17617), .A2(n17618), .ZN(n17616) );
  NAND2_X1 U12266 ( .A1(n17632), .A2(n15361), .ZN(n17614) );
  XNOR2_X1 U12267 ( .A(n15359), .B(n9938), .ZN(n17633) );
  INV_X1 U12268 ( .A(n15360), .ZN(n9938) );
  NAND2_X1 U12269 ( .A1(n17633), .A2(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n17632) );
  NOR2_X1 U12270 ( .A1(n18668), .A2(n15217), .ZN(n18449) );
  XNOR2_X1 U12271 ( .A(n15328), .B(n20894), .ZN(n17653) );
  NOR2_X1 U12272 ( .A1(n17654), .A2(n17653), .ZN(n17652) );
  NOR2_X1 U12273 ( .A1(n11804), .A2(n11803), .ZN(n15229) );
  INV_X1 U12274 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n18288) );
  NAND3_X2 U12275 ( .A1(n11753), .A2(n11752), .A3(n11751), .ZN(n18023) );
  AOI22_X1 U12276 ( .A1(n15294), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n15162), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11752) );
  AOI22_X1 U12277 ( .A1(n16993), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_5__1__SCAN_IN), .B2(n9726), .ZN(n11753) );
  AOI211_X1 U12278 ( .C1(n16975), .C2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A(
        n11750), .B(n11749), .ZN(n11751) );
  NAND3_X1 U12279 ( .A1(n11764), .A2(n11763), .A3(n11762), .ZN(n18027) );
  AOI211_X1 U12280 ( .C1(n16992), .C2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A(
        n11761), .B(n11760), .ZN(n11762) );
  OR2_X1 U12281 ( .A1(n11783), .A2(n11782), .ZN(n18032) );
  INV_X1 U12282 ( .A(n15229), .ZN(n18037) );
  NOR2_X1 U12283 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18011), .ZN(n18362) );
  INV_X1 U12284 ( .A(n13564), .ZN(n18041) );
  AOI211_X1 U12285 ( .C1(n16993), .C2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A(
        n11813), .B(n11812), .ZN(n11814) );
  CLKBUF_X1 U12286 ( .A(n11897), .Z(n14634) );
  AND2_X1 U12287 ( .A1(n15545), .A2(n12843), .ZN(n19816) );
  AND2_X1 U12288 ( .A1(n15545), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n19861) );
  NAND2_X1 U12289 ( .A1(n20664), .A2(n12852), .ZN(n19838) );
  AND2_X1 U12290 ( .A1(n15545), .A2(n12857), .ZN(n19860) );
  AND2_X1 U12291 ( .A1(n20664), .A2(n12856), .ZN(n19850) );
  INV_X1 U12292 ( .A(n14120), .ZN(n19875) );
  NAND2_X2 U12293 ( .A1(n12338), .A2(n12337), .ZN(n19879) );
  INV_X1 U12294 ( .A(n14184), .ZN(n14179) );
  NOR2_X1 U12295 ( .A1(n14194), .A2(n12510), .ZN(n14195) );
  NAND2_X1 U12296 ( .A1(n12509), .A2(n12508), .ZN(n14191) );
  INV_X1 U12297 ( .A(n14195), .ZN(n14193) );
  AND2_X1 U12298 ( .A1(n12311), .A2(n12310), .ZN(n19885) );
  OR3_X1 U12299 ( .A1(n15462), .A2(n19757), .A3(n12790), .ZN(n12309) );
  BUF_X1 U12300 ( .A(n15492), .Z(n19903) );
  INV_X1 U12301 ( .A(n19909), .ZN(n13149) );
  NAND2_X1 U12302 ( .A1(n14412), .A2(n9835), .ZN(n14409) );
  AND2_X1 U12303 ( .A1(n10210), .A2(n10205), .ZN(n14272) );
  AOI21_X1 U12304 ( .B1(n14374), .B2(n15719), .A(n14373), .ZN(n15711) );
  NAND2_X1 U12305 ( .A1(n9911), .A2(n19984), .ZN(n9909) );
  NAND2_X1 U12306 ( .A1(n19963), .A2(n15474), .ZN(n9911) );
  OR2_X1 U12307 ( .A1(n15734), .A2(n15726), .ZN(n15745) );
  NAND2_X1 U12308 ( .A1(n10058), .A2(n10059), .ZN(n13398) );
  NAND2_X1 U12309 ( .A1(n10064), .A2(n13368), .ZN(n15687) );
  NAND2_X1 U12310 ( .A1(n15692), .A2(n13367), .ZN(n10064) );
  OR2_X1 U12311 ( .A1(n13440), .A2(n13009), .ZN(n9910) );
  NAND2_X1 U12312 ( .A1(n15751), .A2(n15472), .ZN(n19963) );
  AND2_X1 U12313 ( .A1(n13440), .A2(n13439), .ZN(n19993) );
  INV_X1 U12314 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20757) );
  INV_X1 U12315 ( .A(n12641), .ZN(n12439) );
  NOR2_X1 U12316 ( .A1(n20275), .A2(n15462), .ZN(n12811) );
  INV_X1 U12317 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n15813) );
  INV_X1 U12318 ( .A(n20203), .ZN(n20206) );
  NOR2_X1 U12319 ( .A1(n20435), .A2(n20241), .ZN(n20261) );
  INV_X1 U12320 ( .A(n20258), .ZN(n20292) );
  OAI211_X1 U12321 ( .C1(n20409), .C2(n12396), .A(n20473), .B(n20408), .ZN(
        n20430) );
  OAI211_X1 U12322 ( .C1(n20503), .C2(n20474), .A(n20473), .B(n20472), .ZN(
        n20507) );
  INV_X1 U12323 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n20898) );
  INV_X1 U12324 ( .A(n15818), .ZN(n15824) );
  AOI221_X1 U12325 ( .B1(n15822), .B2(n20898), .C1(n15458), .C2(n20898), .A(
        n15817), .ZN(n15823) );
  AND2_X1 U12326 ( .A1(n11939), .A2(n18949), .ZN(n19735) );
  NAND2_X1 U12327 ( .A1(n15879), .A2(n18863), .ZN(n15867) );
  NAND2_X1 U12328 ( .A1(n15890), .A2(n18863), .ZN(n15880) );
  NAND2_X1 U12329 ( .A1(n15880), .A2(n15881), .ZN(n15879) );
  NAND2_X1 U12330 ( .A1(n15919), .A2(n18863), .ZN(n15910) );
  NAND2_X1 U12331 ( .A1(n15833), .A2(n18863), .ZN(n15920) );
  NAND2_X1 U12332 ( .A1(n15920), .A2(n15921), .ZN(n15919) );
  NAND2_X1 U12333 ( .A1(n18701), .A2(n18863), .ZN(n15413) );
  NAND2_X1 U12334 ( .A1(n15413), .A2(n15960), .ZN(n15833) );
  NAND2_X1 U12335 ( .A1(n18702), .A2(n18703), .ZN(n18701) );
  NAND2_X1 U12336 ( .A1(n12951), .A2(n9836), .ZN(n18724) );
  INV_X1 U12337 ( .A(n18737), .ZN(n10026) );
  NAND2_X1 U12338 ( .A1(n18724), .A2(n18725), .ZN(n18723) );
  NAND2_X1 U12339 ( .A1(n10010), .A2(n11250), .ZN(n11244) );
  NOR2_X1 U12340 ( .A1(n11261), .A2(n10011), .ZN(n10010) );
  INV_X1 U12341 ( .A(n19614), .ZN(n10036) );
  OR2_X1 U12342 ( .A1(n10587), .A2(n10586), .ZN(n12891) );
  OR2_X1 U12343 ( .A1(n10516), .A2(n10515), .ZN(n12518) );
  OR2_X1 U12344 ( .A1(n10541), .A2(n10540), .ZN(n12301) );
  NAND2_X1 U12345 ( .A1(n12214), .A2(n10496), .ZN(n12233) );
  INV_X1 U12346 ( .A(n14601), .ZN(n14630) );
  AND2_X1 U12347 ( .A1(n10807), .A2(n10173), .ZN(n14550) );
  NOR2_X1 U12348 ( .A1(n14575), .A2(n14574), .ZN(n14573) );
  AND2_X1 U12349 ( .A1(n10180), .A2(n10179), .ZN(n14575) );
  INV_X1 U12350 ( .A(n10180), .ZN(n14588) );
  INV_X1 U12351 ( .A(n18930), .ZN(n14709) );
  AND2_X1 U12352 ( .A1(n18948), .A2(n10383), .ZN(n18930) );
  NOR2_X1 U12353 ( .A1(n15077), .A2(n11972), .ZN(n18912) );
  AND2_X1 U12354 ( .A1(n18948), .A2(n11965), .ZN(n15928) );
  NAND2_X1 U12355 ( .A1(n10223), .A2(n14845), .ZN(n16000) );
  INV_X1 U12356 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n16021) );
  INV_X1 U12357 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n16065) );
  INV_X1 U12358 ( .A(n16054), .ZN(n19045) );
  INV_X1 U12359 ( .A(n16064), .ZN(n19032) );
  AOI211_X1 U12360 ( .C1(n15843), .C2(n19059), .A(n14870), .B(n14869), .ZN(
        n14873) );
  AOI21_X1 U12361 ( .B1(n10223), .B2(n10228), .A(n11397), .ZN(n14954) );
  NAND2_X1 U12362 ( .A1(n9984), .A2(n9982), .ZN(n15421) );
  NAND2_X1 U12363 ( .A1(n9984), .A2(n14781), .ZN(n15419) );
  NAND2_X1 U12364 ( .A1(n14780), .A2(n15988), .ZN(n14826) );
  AND2_X1 U12365 ( .A1(n10242), .A2(n9831), .ZN(n14857) );
  NAND2_X1 U12366 ( .A1(n10242), .A2(n11315), .ZN(n15029) );
  NAND2_X1 U12367 ( .A1(n15060), .A2(n15059), .ZN(n9923) );
  NAND2_X1 U12368 ( .A1(n9960), .A2(n12922), .ZN(n12823) );
  INV_X1 U12369 ( .A(n19059), .ZN(n16131) );
  INV_X1 U12370 ( .A(n14998), .ZN(n16163) );
  INV_X1 U12371 ( .A(n18912), .ZN(n19716) );
  INV_X1 U12372 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19704) );
  INV_X1 U12373 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n15508) );
  XNOR2_X1 U12374 ( .A(n12203), .B(n12202), .ZN(n19707) );
  AND2_X1 U12375 ( .A1(n12976), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n16199) );
  INV_X1 U12376 ( .A(n11983), .ZN(n11984) );
  OAI21_X1 U12377 ( .B1(n19219), .B2(n19203), .A(n19202), .ZN(n19221) );
  OR3_X1 U12378 ( .A1(n19262), .A2(n19261), .A3(n19426), .ZN(n19281) );
  OAI21_X1 U12379 ( .B1(n19312), .B2(n19311), .A(n19310), .ZN(n19330) );
  OAI21_X1 U12380 ( .B1(n19377), .B2(n19393), .A(n19549), .ZN(n19396) );
  AND2_X1 U12381 ( .A1(n19334), .A2(n19338), .ZN(n19395) );
  OAI22_X1 U12382 ( .A1(n16315), .A2(n19080), .B1(n18018), .B2(n19079), .ZN(
        n19465) );
  OR2_X1 U12383 ( .A1(n19424), .A2(n13214), .ZN(n13224) );
  OAI22_X1 U12384 ( .A1(n16308), .A2(n19080), .B1(n18042), .B2(n19079), .ZN(
        n19529) );
  AND2_X1 U12385 ( .A1(n19334), .A2(n19459), .ZN(n19537) );
  AND2_X1 U12386 ( .A1(n10944), .A2(n19076), .ZN(n19559) );
  AND2_X1 U12387 ( .A1(n10389), .A2(n19076), .ZN(n19571) );
  INV_X1 U12388 ( .A(n19504), .ZN(n19591) );
  OAI22_X1 U12389 ( .A1(n16291), .A2(n19080), .B1(n18058), .B2(n19079), .ZN(
        n19599) );
  INV_X1 U12390 ( .A(n13224), .ZN(n19600) );
  OR2_X1 U12391 ( .A1(n12957), .A2(n19744), .ZN(n19607) );
  NAND2_X1 U12392 ( .A1(n18648), .A2(n18443), .ZN(n17238) );
  NOR2_X1 U12393 ( .A1(n18442), .A2(n17238), .ZN(n18669) );
  NOR2_X1 U12394 ( .A1(n16425), .A2(n16426), .ZN(n16424) );
  AOI21_X1 U12395 ( .B1(n16428), .B2(P3_REIP_REG_29__SCAN_IN), .A(n10077), 
        .ZN(n10076) );
  NAND2_X1 U12396 ( .A1(n16429), .A2(n10078), .ZN(n10077) );
  OR2_X1 U12397 ( .A1(n16740), .A2(n16430), .ZN(n10078) );
  AOI21_X1 U12398 ( .B1(n16425), .B2(n16426), .A(n9780), .ZN(n10080) );
  NOR2_X1 U12399 ( .A1(n17374), .A2(n11855), .ZN(n16406) );
  NOR2_X1 U12400 ( .A1(n17412), .A2(n16495), .ZN(n16494) );
  NAND2_X1 U12401 ( .A1(n9742), .A2(n9834), .ZN(n16526) );
  INV_X1 U12402 ( .A(n16751), .ZN(n16711) );
  NOR2_X1 U12403 ( .A1(P3_EBX_REG_7__SCAN_IN), .A2(n16673), .ZN(n16658) );
  NOR2_X2 U12404 ( .A1(n16737), .A2(n18599), .ZN(n16709) );
  INV_X1 U12405 ( .A(n16743), .ZN(n16750) );
  NOR2_X1 U12406 ( .A1(n16806), .A2(n16805), .ZN(n15183) );
  INV_X1 U12407 ( .A(n15183), .ZN(n16801) );
  NAND2_X1 U12408 ( .A1(n16815), .A2(P3_EBX_REG_25__SCAN_IN), .ZN(n16806) );
  NOR3_X1 U12409 ( .A1(n16816), .A2(n16758), .A3(n16812), .ZN(n16815) );
  NOR2_X1 U12410 ( .A1(n16497), .A2(n16848), .ZN(n16822) );
  NOR2_X1 U12411 ( .A1(n16887), .A2(n9992), .ZN(n9991) );
  INV_X1 U12412 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n9992) );
  NAND2_X1 U12413 ( .A1(n16888), .A2(n9784), .ZN(n16872) );
  NAND2_X1 U12414 ( .A1(n16888), .A2(P3_EBX_REG_17__SCAN_IN), .ZN(n16884) );
  NOR2_X1 U12415 ( .A1(n16914), .A2(n16902), .ZN(n16888) );
  NOR2_X1 U12416 ( .A1(n15195), .A2(n16579), .ZN(n9995) );
  NAND2_X1 U12417 ( .A1(n16982), .A2(n9781), .ZN(n15196) );
  AND2_X1 U12418 ( .A1(n16982), .A2(n9872), .ZN(n16939) );
  NOR2_X1 U12419 ( .A1(n17020), .A2(n17019), .ZN(n17015) );
  NOR2_X1 U12420 ( .A1(n16726), .A2(n17027), .ZN(n17023) );
  INV_X1 U12421 ( .A(n18052), .ZN(n17047) );
  NAND2_X1 U12422 ( .A1(P3_EBX_REG_1__SCAN_IN), .A2(n17041), .ZN(n17027) );
  AND2_X1 U12423 ( .A1(n9994), .A2(n9993), .ZN(n17034) );
  NOR2_X1 U12424 ( .A1(n16208), .A2(n16694), .ZN(n9993) );
  AND2_X1 U12425 ( .A1(n17034), .A2(P3_EBX_REG_0__SCAN_IN), .ZN(n17041) );
  INV_X1 U12426 ( .A(n17056), .ZN(n17052) );
  NAND2_X1 U12427 ( .A1(P3_EAX_REG_27__SCAN_IN), .A2(n17073), .ZN(n17068) );
  NOR2_X1 U12428 ( .A1(n20918), .A2(n17077), .ZN(n17073) );
  INV_X1 U12429 ( .A(n17082), .ZN(n17078) );
  NAND2_X1 U12430 ( .A1(P3_EAX_REG_25__SCAN_IN), .A2(n17078), .ZN(n17077) );
  INV_X1 U12431 ( .A(n17102), .ZN(n17099) );
  NOR2_X1 U12432 ( .A1(n17092), .A2(n17117), .ZN(n17106) );
  NOR2_X1 U12433 ( .A1(n17160), .A2(n17044), .ZN(n17045) );
  NAND2_X1 U12434 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(n17167), .ZN(n17160) );
  NOR2_X1 U12435 ( .A1(n15285), .A2(n15284), .ZN(n17181) );
  NOR2_X1 U12436 ( .A1(n17047), .A2(n17192), .ZN(n17185) );
  NOR2_X1 U12437 ( .A1(n15303), .A2(n10090), .ZN(n10089) );
  NOR3_X1 U12438 ( .A1(n15509), .A2(n18012), .A3(n18023), .ZN(n15510) );
  INV_X1 U12439 ( .A(n9994), .ZN(n15509) );
  OR2_X1 U12440 ( .A1(n9940), .A2(n15323), .ZN(n17673) );
  NOR2_X1 U12441 ( .A1(n18464), .A2(n17192), .ZN(n17188) );
  NOR2_X1 U12442 ( .A1(n17235), .A2(n17218), .ZN(n17215) );
  CLKBUF_X1 U12444 ( .A(n17300), .Z(n17293) );
  NOR2_X1 U12445 ( .A1(n17385), .A2(n11849), .ZN(n17376) );
  NOR2_X1 U12446 ( .A1(n17430), .A2(n17431), .ZN(n17423) );
  INV_X1 U12447 ( .A(n17506), .ZN(n17496) );
  INV_X1 U12448 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n20957) );
  INV_X1 U12449 ( .A(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17645) );
  INV_X1 U12450 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n17662) );
  NAND2_X1 U12451 ( .A1(n18362), .A2(n18083), .ZN(n18057) );
  INV_X1 U12452 ( .A(n17667), .ZN(n17678) );
  INV_X1 U12453 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n18610) );
  AND2_X1 U12454 ( .A1(n17807), .A2(n9782), .ZN(n17347) );
  NAND2_X1 U12455 ( .A1(n17419), .A2(n15378), .ZN(n17358) );
  AND2_X1 U12456 ( .A1(n16279), .A2(n17786), .ZN(n17741) );
  NOR2_X1 U12457 ( .A1(n17741), .A2(n17928), .ZN(n17769) );
  INV_X1 U12458 ( .A(n17815), .ZN(n17910) );
  INV_X1 U12459 ( .A(n15341), .ZN(n17598) );
  NAND2_X1 U12460 ( .A1(n10083), .A2(n10084), .ZN(n17627) );
  INV_X1 U12461 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18013) );
  INV_X1 U12462 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18487) );
  INV_X1 U12463 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n16695) );
  NOR2_X1 U12464 ( .A1(n18504), .A2(n18666), .ZN(n18648) );
  CLKBUF_X1 U12465 ( .A(n18587), .Z(n18579) );
  NOR2_X1 U12466 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n20812), .ZN(n18584) );
  INV_X1 U12467 ( .A(n18584), .ZN(n18663) );
  AOI21_X1 U12469 ( .B1(n14229), .B2(n9727), .A(n14228), .ZN(n14230) );
  OAI21_X1 U12470 ( .B1(n14402), .B2(n19964), .A(n10098), .ZN(P1_U3001) );
  AND2_X1 U12471 ( .A1(n10100), .A2(n10099), .ZN(n10098) );
  AOI21_X1 U12472 ( .B1(n14401), .B2(n14400), .A(n14399), .ZN(n10099) );
  OR2_X1 U12473 ( .A1(n14398), .A2(n15807), .ZN(n10100) );
  NAND2_X1 U12474 ( .A1(n10067), .A2(n9806), .ZN(P1_U3006) );
  NAND2_X1 U12475 ( .A1(n14450), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n10066) );
  NAND2_X1 U12476 ( .A1(n10039), .A2(n18863), .ZN(n15845) );
  NAND2_X1 U12477 ( .A1(n10037), .A2(n10031), .ZN(n15847) );
  NAND2_X1 U12478 ( .A1(n15858), .A2(n15859), .ZN(n15857) );
  NAND2_X1 U12479 ( .A1(n10027), .A2(n18863), .ZN(n15891) );
  NAND2_X1 U12480 ( .A1(n15901), .A2(n15902), .ZN(n15900) );
  NAND2_X1 U12481 ( .A1(n18736), .A2(n18737), .ZN(n18735) );
  NAND2_X1 U12482 ( .A1(n14601), .A2(n10168), .ZN(n10166) );
  AND2_X1 U12483 ( .A1(n11705), .A2(n11704), .ZN(n11706) );
  INV_X1 U12484 ( .A(n11703), .ZN(n11704) );
  OAI21_X1 U12485 ( .B1(n16085), .B2(n19037), .A(n9985), .ZN(P2_U2995) );
  AND2_X1 U12486 ( .A1(n15977), .A2(n9986), .ZN(n9985) );
  NOR2_X1 U12487 ( .A1(n9988), .A2(n9987), .ZN(n9986) );
  AND2_X1 U12488 ( .A1(n11683), .A2(n11682), .ZN(n11684) );
  INV_X1 U12489 ( .A(n9933), .ZN(n9932) );
  OAI21_X1 U12490 ( .B1(n14906), .B2(n19056), .A(n9934), .ZN(n9933) );
  OAI21_X1 U12491 ( .B1(n10079), .B2(n16424), .A(n10074), .ZN(P3_U2642) );
  NOR2_X1 U12492 ( .A1(n16427), .A2(n10075), .ZN(n10074) );
  INV_X1 U12493 ( .A(n10080), .ZN(n10079) );
  INV_X1 U12494 ( .A(n10076), .ZN(n10075) );
  AND2_X1 U12495 ( .A1(n16982), .A2(P3_EBX_REG_10__SCAN_IN), .ZN(n16952) );
  AOI21_X1 U12496 ( .B1(n9949), .B2(n9945), .A(n9944), .ZN(n17693) );
  AND2_X1 U12497 ( .A1(n17918), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n9944) );
  BUF_X1 U12498 ( .A(n11788), .Z(n16992) );
  NAND2_X1 U12499 ( .A1(n14045), .A2(n9825), .ZN(n14022) );
  INV_X1 U12500 ( .A(n10869), .ZN(n10407) );
  AND2_X1 U12501 ( .A1(n9725), .A2(n13438), .ZN(n9759) );
  INV_X1 U12502 ( .A(n12951), .ZN(n18903) );
  AOI22_X1 U12503 ( .A1(n12950), .A2(n18954), .B1(P2_STATE2_REG_0__SCAN_IN), 
        .B2(n12949), .ZN(n12951) );
  OR2_X1 U12504 ( .A1(n13458), .A2(n10140), .ZN(n13588) );
  NOR2_X1 U12505 ( .A1(n14751), .A2(n14895), .ZN(n14727) );
  AND2_X1 U12506 ( .A1(n14825), .A2(n15988), .ZN(n9760) );
  AND2_X1 U12507 ( .A1(n15788), .A2(n9877), .ZN(n9761) );
  AND4_X1 U12508 ( .A1(n12038), .A2(n12037), .A3(n12036), .A4(n12035), .ZN(
        n9762) );
  AND2_X1 U12509 ( .A1(n14097), .A2(n10130), .ZN(n14079) );
  AND2_X1 U12510 ( .A1(n16982), .A2(n9875), .ZN(n9763) );
  AND2_X1 U12511 ( .A1(n10089), .A2(n9802), .ZN(n17199) );
  OR3_X1 U12512 ( .A1(n14095), .A2(n10105), .A3(n9874), .ZN(n9764) );
  AND2_X1 U12513 ( .A1(n10001), .A2(n12722), .ZN(n9765) );
  AND2_X1 U12514 ( .A1(n12117), .A2(n12180), .ZN(n9766) );
  AND2_X1 U12515 ( .A1(n9761), .A2(n10101), .ZN(n9767) );
  NOR3_X1 U12516 ( .A1(n12900), .A2(n10194), .A3(n12899), .ZN(n9768) );
  AND2_X1 U12517 ( .A1(n18863), .A2(n10038), .ZN(n9769) );
  AND2_X1 U12518 ( .A1(n10072), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n9770) );
  AND2_X1 U12519 ( .A1(n13288), .A2(n13330), .ZN(n9771) );
  AND2_X1 U12520 ( .A1(n10041), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n9772) );
  AND2_X1 U12521 ( .A1(n10044), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n9773) );
  AND2_X1 U12522 ( .A1(n9771), .A2(n9878), .ZN(n9774) );
  AND2_X1 U12523 ( .A1(n10146), .A2(n11079), .ZN(n9775) );
  AND2_X1 U12524 ( .A1(n9770), .A2(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n9776) );
  AND2_X1 U12525 ( .A1(n10047), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n9777) );
  AND2_X1 U12526 ( .A1(n10108), .A2(n13984), .ZN(n9778) );
  OR2_X1 U12527 ( .A1(n10169), .A2(n10171), .ZN(n9779) );
  OR4_X1 U12528 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(P3_STATE2_REG_0__SCAN_IN), 
        .A3(P3_STATEBS16_REG_SCAN_IN), .A4(n18610), .ZN(n9780) );
  AND2_X1 U12529 ( .A1(n9872), .A2(P3_EBX_REG_12__SCAN_IN), .ZN(n9781) );
  AND2_X1 U12530 ( .A1(n17366), .A2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n9782) );
  AND2_X1 U12531 ( .A1(n10252), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n9783) );
  AND2_X1 U12532 ( .A1(n9991), .A2(P3_EBX_REG_19__SCAN_IN), .ZN(n9784) );
  AND2_X2 U12533 ( .A1(n10510), .A2(n10674), .ZN(n10535) );
  AND2_X2 U12534 ( .A1(n10833), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10935) );
  AND2_X2 U12535 ( .A1(n10508), .A2(n10674), .ZN(n10523) );
  NAND2_X1 U12536 ( .A1(n16273), .A2(n15338), .ZN(n17551) );
  AND2_X1 U12537 ( .A1(n14039), .A2(n10108), .ZN(n9786) );
  OR2_X1 U12538 ( .A1(n14590), .A2(n14589), .ZN(n10180) );
  NAND2_X1 U12539 ( .A1(n14761), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14751) );
  NAND2_X1 U12540 ( .A1(n15644), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n10210) );
  NAND2_X1 U12541 ( .A1(n14819), .A2(n11672), .ZN(n14802) );
  AND2_X1 U12542 ( .A1(n9969), .A2(n9967), .ZN(n9788) );
  INV_X2 U12543 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10359) );
  NAND4_X1 U12544 ( .A1(n9725), .A2(n10264), .A3(n12118), .A4(n9920), .ZN(
        n9789) );
  NAND2_X1 U12545 ( .A1(n14819), .A2(n10252), .ZN(n14797) );
  INV_X1 U12546 ( .A(n10233), .ZN(n10236) );
  XNOR2_X1 U12547 ( .A(n13973), .B(n13972), .ZN(n14398) );
  AND2_X1 U12548 ( .A1(n15950), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n9790) );
  AND3_X1 U12549 ( .A1(n10338), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        n10337), .ZN(n9792) );
  INV_X2 U12550 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12778) );
  NOR2_X1 U12551 ( .A1(n14044), .A2(n14146), .ZN(n14031) );
  AND2_X1 U12552 ( .A1(n11146), .A2(n11118), .ZN(n9794) );
  AND2_X1 U12553 ( .A1(n14679), .A2(n10149), .ZN(n9795) );
  NAND2_X1 U12554 ( .A1(n14097), .A2(n10132), .ZN(n14076) );
  NAND2_X1 U12555 ( .A1(n9923), .A2(n11506), .ZN(n15040) );
  NAND2_X1 U12556 ( .A1(n11403), .A2(n14956), .ZN(n9796) );
  NAND2_X1 U12557 ( .A1(n12743), .A2(n12669), .ZN(n12864) );
  AND4_X1 U12558 ( .A1(n12034), .A2(n12033), .A3(n12032), .A4(n12031), .ZN(
        n9797) );
  NAND2_X1 U12559 ( .A1(n11155), .A2(n15084), .ZN(n11199) );
  NAND2_X2 U12560 ( .A1(n10366), .A2(n10367), .ZN(n10927) );
  AND2_X1 U12561 ( .A1(n16176), .A2(n10427), .ZN(n9798) );
  NOR2_X1 U12562 ( .A1(n13458), .A2(n10138), .ZN(n9799) );
  OR2_X1 U12563 ( .A1(n11089), .A2(n13175), .ZN(n9800) );
  AND2_X1 U12564 ( .A1(n14680), .A2(n14681), .ZN(n14679) );
  NOR2_X1 U12565 ( .A1(n12171), .A2(n9901), .ZN(n9801) );
  OR2_X1 U12566 ( .A1(n14751), .A2(n10251), .ZN(n14716) );
  AND4_X1 U12567 ( .A1(n15302), .A2(n15301), .A3(n15300), .A4(n15299), .ZN(
        n9802) );
  OR2_X1 U12568 ( .A1(n13399), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n9803) );
  OR2_X1 U12569 ( .A1(n10771), .A2(n10770), .ZN(n9804) );
  NAND2_X1 U12570 ( .A1(n12341), .A2(n13437), .ZN(n9805) );
  OR2_X1 U12571 ( .A1(n11113), .A2(n18926), .ZN(n11135) );
  NOR2_X1 U12572 ( .A1(n13458), .A2(n10135), .ZN(n14106) );
  AND2_X1 U12573 ( .A1(n10066), .A2(n10065), .ZN(n9806) );
  NOR2_X1 U12574 ( .A1(n15685), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n9807) );
  NAND2_X1 U12575 ( .A1(n10003), .A2(n15659), .ZN(n9808) );
  OR3_X1 U12576 ( .A1(n14751), .A2(n10251), .A3(n10250), .ZN(n9809) );
  NAND2_X1 U12577 ( .A1(n10218), .A2(n11166), .ZN(n9810) );
  INV_X2 U12578 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n12690) );
  NAND2_X1 U12579 ( .A1(n11398), .A2(n10015), .ZN(n10019) );
  NOR2_X1 U12580 ( .A1(n11773), .A2(n9989), .ZN(n9811) );
  INV_X1 U12581 ( .A(n13563), .ZN(n15219) );
  NAND2_X1 U12582 ( .A1(n18032), .A2(n18052), .ZN(n13563) );
  OR2_X1 U12583 ( .A1(n11199), .A2(n20884), .ZN(n9812) );
  NAND2_X1 U12584 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13568) );
  INV_X1 U12585 ( .A(n13568), .ZN(n9898) );
  AND2_X1 U12586 ( .A1(n10051), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n9813) );
  OR2_X1 U12587 ( .A1(n15657), .A2(n14214), .ZN(n9814) );
  OR2_X1 U12588 ( .A1(n14354), .A2(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n9815) );
  INV_X1 U12589 ( .A(n16007), .ZN(n9976) );
  AND2_X1 U12590 ( .A1(n10059), .A2(n9803), .ZN(n9816) );
  AND2_X1 U12591 ( .A1(n10188), .A2(n10187), .ZN(n9817) );
  AND2_X1 U12592 ( .A1(n12082), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n9818) );
  NAND2_X1 U12593 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n15333), .ZN(
        n9819) );
  AND2_X1 U12594 ( .A1(n10236), .A2(n10235), .ZN(n9820) );
  INV_X1 U12595 ( .A(n9893), .ZN(n16282) );
  OR2_X1 U12596 ( .A1(n9895), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n9893) );
  AND2_X1 U12597 ( .A1(n14515), .A2(n12784), .ZN(n12082) );
  NAND4_X2 U12598 ( .A1(n11050), .A2(n11049), .A3(n11048), .A4(n11047), .ZN(
        n11307) );
  INV_X1 U12599 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n10862) );
  OAI21_X1 U12600 ( .B1(n15472), .B2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n9910), .ZN(n19962) );
  NOR2_X1 U12601 ( .A1(n20269), .A2(n20013), .ZN(n9821) );
  NOR2_X1 U12602 ( .A1(n11251), .A2(n11256), .ZN(n11250) );
  INV_X1 U12603 ( .A(n10926), .ZN(n11000) );
  INV_X1 U12604 ( .A(n11000), .ZN(n11085) );
  NOR2_X2 U12605 ( .A1(n10390), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n10926) );
  INV_X1 U12606 ( .A(n15402), .ZN(n10052) );
  NAND2_X1 U12607 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n11957) );
  NOR2_X1 U12608 ( .A1(n14095), .A2(n10102), .ZN(n10107) );
  XOR2_X1 U12609 ( .A(n11483), .B(n19067), .Z(n9822) );
  AND2_X1 U12610 ( .A1(n15400), .A2(n10041), .ZN(n9823) );
  NAND2_X1 U12611 ( .A1(n10156), .A2(n10157), .ZN(n9824) );
  AND2_X1 U12612 ( .A1(n14032), .A2(n10117), .ZN(n9825) );
  AND2_X1 U12613 ( .A1(n13265), .A2(n13266), .ZN(n13320) );
  AND2_X1 U12614 ( .A1(n10197), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n9826) );
  AND2_X1 U12615 ( .A1(n10197), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n9827) );
  AND2_X1 U12616 ( .A1(n10197), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n9828) );
  NAND2_X1 U12617 ( .A1(n9890), .A2(n11264), .ZN(n16044) );
  AND2_X1 U12618 ( .A1(n13393), .A2(n14623), .ZN(n9829) );
  NAND2_X1 U12619 ( .A1(n9961), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12921) );
  AND2_X1 U12620 ( .A1(n9966), .A2(n9798), .ZN(n10916) );
  AND2_X1 U12621 ( .A1(n19988), .A2(n14381), .ZN(n9830) );
  AND2_X1 U12622 ( .A1(n10244), .A2(n11315), .ZN(n9831) );
  AND2_X1 U12623 ( .A1(n9829), .A2(n14617), .ZN(n9832) );
  INV_X1 U12624 ( .A(n9724), .ZN(n13931) );
  AND2_X1 U12625 ( .A1(n16888), .A2(n9991), .ZN(n9833) );
  OR2_X1 U12626 ( .A1(n16536), .A2(n16549), .ZN(n9834) );
  INV_X1 U12627 ( .A(n9908), .ZN(n15719) );
  OR2_X1 U12628 ( .A1(n14372), .A2(n9909), .ZN(n9908) );
  OR2_X1 U12629 ( .A1(n14468), .A2(n14389), .ZN(n9835) );
  OR2_X1 U12630 ( .A1(n10273), .A2(n10026), .ZN(n9836) );
  INV_X1 U12631 ( .A(n10186), .ZN(n13331) );
  NAND2_X1 U12632 ( .A1(n13289), .A2(n13288), .ZN(n10186) );
  AND2_X1 U12633 ( .A1(n12165), .A2(n12166), .ZN(n9837) );
  INV_X1 U12634 ( .A(n10247), .ZN(n11525) );
  NAND2_X1 U12635 ( .A1(n10910), .A2(n10406), .ZN(n10247) );
  AND2_X1 U12636 ( .A1(n12082), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n9838) );
  AND2_X1 U12637 ( .A1(n12082), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n9839) );
  AND2_X1 U12638 ( .A1(n12082), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n9840) );
  AND2_X1 U12639 ( .A1(n12082), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n9841) );
  AND2_X1 U12640 ( .A1(n14593), .A2(n14594), .ZN(n14585) );
  OR2_X1 U12641 ( .A1(n12900), .A2(n10192), .ZN(n9842) );
  NAND2_X1 U12642 ( .A1(n19988), .A2(n15714), .ZN(n9843) );
  AND2_X1 U12643 ( .A1(n11387), .A2(n11598), .ZN(n15997) );
  NAND2_X1 U12644 ( .A1(n10276), .A2(n11396), .ZN(n11397) );
  INV_X1 U12645 ( .A(n16010), .ZN(n11327) );
  AND2_X1 U12646 ( .A1(n12736), .A2(n12735), .ZN(n9844) );
  AND2_X1 U12647 ( .A1(n11166), .A2(n11195), .ZN(n9845) );
  AND2_X1 U12648 ( .A1(n9767), .A2(n13286), .ZN(n9846) );
  INV_X1 U12649 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n18860) );
  INV_X1 U12650 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n9972) );
  AND2_X1 U12651 ( .A1(n12230), .A2(n10565), .ZN(n12516) );
  AND2_X1 U12652 ( .A1(n15789), .A2(n9767), .ZN(n9847) );
  INV_X1 U12653 ( .A(n11332), .ZN(n10025) );
  INV_X1 U12654 ( .A(n11399), .ZN(n10018) );
  AND2_X1 U12655 ( .A1(n15789), .A2(n15788), .ZN(n9848) );
  AND2_X1 U12656 ( .A1(n15395), .A2(n10044), .ZN(n9849) );
  AND2_X1 U12657 ( .A1(n15835), .A2(n10047), .ZN(n9850) );
  AND2_X1 U12658 ( .A1(n14054), .A2(n13514), .ZN(n9851) );
  AND2_X1 U12659 ( .A1(n10197), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n9852) );
  AND2_X1 U12660 ( .A1(n10197), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n9853) );
  AND2_X1 U12661 ( .A1(n10197), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n9854) );
  AND2_X1 U12662 ( .A1(n10197), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n9855) );
  AND2_X1 U12663 ( .A1(n10197), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n9856) );
  AND2_X1 U12664 ( .A1(n10197), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n9857) );
  AND2_X1 U12665 ( .A1(n10197), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n9858) );
  AND2_X1 U12666 ( .A1(n10197), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n9859) );
  AND2_X1 U12667 ( .A1(n14542), .A2(n14532), .ZN(n9860) );
  AND2_X1 U12668 ( .A1(n10110), .A2(n14019), .ZN(n9861) );
  AND2_X1 U12669 ( .A1(n10197), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n9862) );
  INV_X1 U12670 ( .A(n14574), .ZN(n10176) );
  NAND4_X2 U12671 ( .A1(n12058), .A2(n12057), .A3(n12056), .A4(n12055), .ZN(
        n12539) );
  INV_X1 U12672 ( .A(n12539), .ZN(n20047) );
  AND2_X1 U12673 ( .A1(n10907), .A2(n10425), .ZN(n10919) );
  NAND2_X1 U12674 ( .A1(n11989), .A2(n11980), .ZN(n15031) );
  INV_X1 U12675 ( .A(n10171), .ZN(n10170) );
  NOR2_X1 U12676 ( .A1(n10830), .A2(n10172), .ZN(n10171) );
  NAND2_X1 U12677 ( .A1(n10726), .A2(n10725), .ZN(n9863) );
  AND2_X1 U12678 ( .A1(n14601), .A2(n9779), .ZN(n9864) );
  AND2_X1 U12679 ( .A1(n10149), .A2(n14656), .ZN(n9865) );
  AND2_X1 U12680 ( .A1(n9860), .A2(n11710), .ZN(n9866) );
  INV_X1 U12681 ( .A(n14704), .ZN(n10148) );
  INV_X1 U12682 ( .A(n12844), .ZN(n9906) );
  AND2_X1 U12683 ( .A1(n17333), .A2(n10072), .ZN(n9867) );
  INV_X1 U12684 ( .A(n11548), .ZN(n11561) );
  AND2_X1 U12685 ( .A1(n10197), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n9868) );
  AND2_X1 U12686 ( .A1(n10197), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n9869) );
  AND2_X1 U12687 ( .A1(n10197), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n9870) );
  AND2_X1 U12688 ( .A1(n10197), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n9871) );
  AND2_X1 U12689 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(P3_EBX_REG_11__SCAN_IN), 
        .ZN(n9872) );
  NOR2_X1 U12690 ( .A1(n17642), .A2(n15332), .ZN(n9873) );
  NAND2_X1 U12691 ( .A1(n13922), .A2(n13921), .ZN(n9874) );
  AND2_X1 U12692 ( .A1(n9781), .A2(n9995), .ZN(n9875) );
  AND2_X1 U12693 ( .A1(n9782), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n9876) );
  NAND2_X1 U12694 ( .A1(n13105), .A2(n13104), .ZN(n9877) );
  INV_X1 U12695 ( .A(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n10073) );
  INV_X1 U12696 ( .A(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n10050) );
  OR2_X1 U12697 ( .A1(n10640), .A2(n10639), .ZN(n9878) );
  NAND3_X1 U12698 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n9879) );
  INV_X1 U12699 ( .A(n10269), .ZN(n10240) );
  AND2_X1 U12700 ( .A1(n10258), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n9880) );
  NAND2_X1 U12701 ( .A1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n9881) );
  INV_X1 U12702 ( .A(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n10045) );
  INV_X1 U12703 ( .A(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n10049) );
  INV_X1 U12704 ( .A(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n10048) );
  INV_X1 U12705 ( .A(n9780), .ZN(n9882) );
  AOI22_X2 U12706 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n20046), .B1(DATAI_28_), 
        .B2(n20007), .ZN(n20553) );
  AOI22_X2 U12707 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n20046), .B1(DATAI_18_), 
        .B2(n20007), .ZN(n20486) );
  NOR3_X2 U12708 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18357), .A3(
        n18240), .ZN(n18210) );
  NOR3_X2 U12709 ( .A1(n18357), .A2(n18288), .A3(n18149), .ZN(n18120) );
  AOI22_X2 U12710 ( .A1(DATAI_17_), .A2(n20007), .B1(BUF1_REG_17__SCAN_IN), 
        .B2(n20046), .ZN(n20482) );
  AOI22_X1 U12711 ( .A1(n13867), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10197), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13844) );
  AOI22_X1 U12712 ( .A1(n13843), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n10197), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n13804) );
  AOI22_X1 U12713 ( .A1(n13867), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10197), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n13460) );
  AND3_X2 U12714 ( .A1(n10280), .A2(n9883), .A3(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10346) );
  OAI21_X2 U12715 ( .B1(n14732), .B2(n14730), .A(n14728), .ZN(n14722) );
  AND3_X2 U12716 ( .A1(n9884), .A2(n10239), .A3(n10238), .ZN(n14732) );
  AND2_X2 U12717 ( .A1(n10408), .A2(n10409), .ZN(n11538) );
  NAND3_X1 U12718 ( .A1(n9960), .A2(n12922), .A3(n9888), .ZN(n9890) );
  NAND2_X1 U12719 ( .A1(n9889), .A2(n11266), .ZN(n13273) );
  INV_X1 U12720 ( .A(n11196), .ZN(n9891) );
  NAND2_X1 U12721 ( .A1(n9936), .A2(n9932), .ZN(P2_U3019) );
  OR2_X2 U12722 ( .A1(n14846), .A2(n14775), .ZN(n10230) );
  NOR2_X1 U12723 ( .A1(n16007), .A2(n11327), .ZN(n14846) );
  NAND2_X1 U12724 ( .A1(n11312), .A2(n10277), .ZN(n10245) );
  NOR2_X2 U12725 ( .A1(n17309), .A2(n17308), .ZN(n17307) );
  NOR2_X2 U12726 ( .A1(n17370), .A2(n9897), .ZN(n17349) );
  NAND3_X1 U12727 ( .A1(n15295), .A2(n15296), .A3(n15297), .ZN(n17187) );
  OR2_X2 U12728 ( .A1(n17480), .A2(n16238), .ZN(n17465) );
  INV_X2 U12729 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n18630) );
  AND2_X4 U12730 ( .A1(n12690), .A2(n12553), .ZN(n14516) );
  NOR2_X2 U12731 ( .A1(n9725), .A2(n13438), .ZN(n12844) );
  NAND2_X1 U12732 ( .A1(n12539), .A2(n9919), .ZN(n13891) );
  AND2_X1 U12733 ( .A1(n12121), .A2(n9919), .ZN(n12093) );
  NAND2_X1 U12734 ( .A1(n20038), .A2(n9919), .ZN(n12334) );
  AOI21_X1 U12735 ( .B1(n12564), .B2(n20042), .A(n20047), .ZN(n9918) );
  OR2_X2 U12736 ( .A1(n12019), .A2(n12020), .ZN(n9919) );
  NAND4_X1 U12737 ( .A1(n9725), .A2(n10264), .A3(n12118), .A4(n12539), .ZN(
        n12340) );
  XNOR2_X1 U12738 ( .A(n9750), .B(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15659) );
  NAND3_X1 U12739 ( .A1(n10003), .A2(n9815), .A3(n15659), .ZN(n14215) );
  NOR2_X1 U12740 ( .A1(n14215), .A2(n10213), .ZN(n10211) );
  AND2_X2 U12741 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11447) );
  NAND3_X1 U12742 ( .A1(n10427), .A2(n10426), .A3(n10398), .ZN(n10385) );
  INV_X2 U12743 ( .A(n19077), .ZN(n10398) );
  INV_X2 U12744 ( .A(n10418), .ZN(n10427) );
  AND2_X2 U12745 ( .A1(n15950), .A2(n9880), .ZN(n14761) );
  NOR2_X4 U12746 ( .A1(n14952), .A2(n14956), .ZN(n15950) );
  NAND2_X2 U12747 ( .A1(n14819), .A2(n9783), .ZN(n14952) );
  OAI21_X1 U12748 ( .B1(n9926), .B2(n15060), .A(n9922), .ZN(n11511) );
  OAI21_X1 U12749 ( .B1(n9928), .B2(n9930), .A(n9927), .ZN(n10414) );
  NAND3_X1 U12750 ( .A1(n10405), .A2(n9931), .A3(n10404), .ZN(n9928) );
  AND3_X2 U12751 ( .A1(n10218), .A2(n10219), .A3(n9845), .ZN(n11196) );
  NAND3_X1 U12752 ( .A1(n9943), .A2(n9941), .A3(n15325), .ZN(n9940) );
  INV_X2 U12753 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n18607) );
  NAND3_X1 U12754 ( .A1(n15374), .A2(n17831), .A3(n17864), .ZN(n9953) );
  NAND2_X2 U12755 ( .A1(n15341), .A2(n10094), .ZN(n15373) );
  AND2_X2 U12756 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10507) );
  AND2_X4 U12757 ( .A1(n10510), .A2(n9955), .ZN(n10672) );
  INV_X2 U12758 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10876) );
  NAND3_X1 U12759 ( .A1(n9959), .A2(n10418), .A3(n10909), .ZN(n10399) );
  INV_X1 U12760 ( .A(n11146), .ZN(n11136) );
  NAND3_X1 U12761 ( .A1(n10368), .A2(n10410), .A3(n19740), .ZN(n10425) );
  NAND3_X1 U12762 ( .A1(n10907), .A2(n10425), .A3(n9964), .ZN(n10436) );
  NAND3_X1 U12763 ( .A1(n9966), .A2(n9798), .A3(n10428), .ZN(n9964) );
  NAND2_X2 U12764 ( .A1(n9965), .A2(n16176), .ZN(n10907) );
  NAND2_X1 U12765 ( .A1(n10452), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n9971) );
  NAND2_X2 U12766 ( .A1(n11666), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10455) );
  NAND2_X1 U12767 ( .A1(n9978), .A2(n9979), .ZN(n14815) );
  NAND2_X2 U12768 ( .A1(n9811), .A2(n11771), .ZN(n18052) );
  NAND3_X1 U12769 ( .A1(n11769), .A2(n11770), .A3(n11772), .ZN(n9989) );
  INV_X2 U12770 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n18617) );
  XNOR2_X2 U12771 ( .A(n9998), .B(n12523), .ZN(n20119) );
  NAND2_X2 U12772 ( .A1(n12428), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12523) );
  NAND3_X1 U12773 ( .A1(n10200), .A2(n10199), .A3(n12424), .ZN(n9998) );
  NAND3_X1 U12774 ( .A1(n10000), .A2(n9766), .A3(n9999), .ZN(n12503) );
  NOR2_X2 U12775 ( .A1(n12095), .A2(n12094), .ZN(n12345) );
  NAND2_X2 U12776 ( .A1(n12503), .A2(n12500), .ZN(n12425) );
  NAND2_X1 U12777 ( .A1(n13415), .A2(n9759), .ZN(n12500) );
  NAND2_X1 U12778 ( .A1(n10210), .A2(n9749), .ZN(n14279) );
  NAND2_X1 U12779 ( .A1(n11316), .A2(n12291), .ZN(n10005) );
  INV_X1 U12780 ( .A(n14765), .ZN(n10007) );
  INV_X1 U12781 ( .A(n11261), .ZN(n10009) );
  NAND2_X1 U12782 ( .A1(n11398), .A2(n11399), .ZN(n11407) );
  INV_X1 U12783 ( .A(n10019), .ZN(n11420) );
  NAND2_X1 U12784 ( .A1(n15909), .A2(n18863), .ZN(n10030) );
  AOI21_X1 U12785 ( .B1(n15866), .B2(n9769), .A(n10032), .ZN(n10031) );
  NAND2_X1 U12786 ( .A1(n15866), .A2(n18863), .ZN(n15858) );
  NAND2_X1 U12787 ( .A1(n10058), .A2(n9816), .ZN(n13401) );
  OR2_X2 U12788 ( .A1(n15692), .A2(n10061), .ZN(n10058) );
  NAND2_X1 U12789 ( .A1(n14323), .A2(n10068), .ZN(n14216) );
  NAND2_X1 U12790 ( .A1(n14323), .A2(n14322), .ZN(n14321) );
  INV_X1 U12791 ( .A(n14322), .ZN(n10069) );
  XNOR2_X2 U12792 ( .A(n10111), .B(n12403), .ZN(n20083) );
  INV_X2 U12793 ( .A(n9742), .ZN(n16667) );
  INV_X2 U12794 ( .A(n17199), .ZN(n15356) );
  NAND3_X1 U12795 ( .A1(n15304), .A2(n15305), .A3(n10091), .ZN(n10090) );
  NAND2_X1 U12796 ( .A1(n15341), .A2(n10261), .ZN(n10093) );
  NAND2_X1 U12797 ( .A1(n10093), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10095) );
  NAND3_X1 U12798 ( .A1(n15373), .A2(n10095), .A3(n17585), .ZN(n17584) );
  NOR2_X1 U12799 ( .A1(n17552), .A2(n17874), .ZN(n17912) );
  AND2_X2 U12800 ( .A1(n12782), .A2(n14516), .ZN(n13477) );
  INV_X1 U12801 ( .A(n10107), .ZN(n14451) );
  NAND2_X1 U12802 ( .A1(n14039), .A2(n9778), .ZN(n13983) );
  AND2_X2 U12803 ( .A1(n10112), .A2(n12784), .ZN(n13862) );
  AND2_X2 U12804 ( .A1(n10112), .A2(n12781), .ZN(n13843) );
  NOR2_X1 U12805 ( .A1(n14044), .A2(n10115), .ZN(n14010) );
  OR2_X2 U12806 ( .A1(n14044), .A2(n10113), .ZN(n13997) );
  NAND2_X1 U12807 ( .A1(n20008), .A2(n12645), .ZN(n10118) );
  NAND2_X1 U12808 ( .A1(n10118), .A2(n10120), .ZN(n12686) );
  INV_X1 U12809 ( .A(n12686), .ZN(n10119) );
  NAND2_X1 U12810 ( .A1(n10119), .A2(n12646), .ZN(n12688) );
  NAND2_X2 U12811 ( .A1(n20042), .A2(n12121), .ZN(n12341) );
  NAND2_X1 U12812 ( .A1(n13369), .A2(n13505), .ZN(n10123) );
  NAND2_X1 U12813 ( .A1(n13985), .A2(n13987), .ZN(n13986) );
  NAND2_X1 U12814 ( .A1(n14097), .A2(n10129), .ZN(n14043) );
  NAND2_X1 U12815 ( .A1(n12486), .A2(n10145), .ZN(n12483) );
  NAND2_X1 U12816 ( .A1(n14679), .A2(n9865), .ZN(n14658) );
  INV_X1 U12817 ( .A(n15031), .ZN(n10153) );
  NAND2_X1 U12818 ( .A1(n10153), .A2(n10154), .ZN(n16098) );
  INV_X2 U12819 ( .A(n11354), .ZN(n12986) );
  NOR2_X1 U12820 ( .A1(n14648), .A2(n10160), .ZN(n14632) );
  INV_X1 U12821 ( .A(n10917), .ZN(n10403) );
  NAND2_X1 U12822 ( .A1(n11531), .A2(n10401), .ZN(n10164) );
  NAND2_X1 U12823 ( .A1(n14535), .A2(n10169), .ZN(n10167) );
  OAI211_X1 U12824 ( .C1(n14535), .C2(n10166), .A(n10165), .B(n11713), .ZN(
        P2_U2857) );
  NAND2_X1 U12825 ( .A1(n14535), .A2(n9864), .ZN(n10165) );
  OAI211_X1 U12826 ( .C1(n14535), .C2(n10172), .A(n10167), .B(n10170), .ZN(
        n11709) );
  NAND3_X1 U12827 ( .A1(n10807), .A2(n10173), .A3(n14549), .ZN(n14548) );
  INV_X1 U12828 ( .A(n10704), .ZN(n10179) );
  NAND2_X1 U12829 ( .A1(n10704), .A2(n10176), .ZN(n10177) );
  NAND2_X1 U12830 ( .A1(n12230), .A2(n10181), .ZN(n13040) );
  NAND2_X2 U12831 ( .A1(n12214), .A2(n10182), .ZN(n12230) );
  NAND2_X2 U12832 ( .A1(n10353), .A2(n10354), .ZN(n10418) );
  NAND4_X1 U12833 ( .A1(n10339), .A2(n10353), .A3(n10340), .A4(n10354), .ZN(
        n10397) );
  NOR2_X1 U12834 ( .A1(n12900), .A2(n12899), .ZN(n12901) );
  INV_X1 U12835 ( .A(n12893), .ZN(n10194) );
  NAND2_X1 U12836 ( .A1(n14543), .A2(n9860), .ZN(n14531) );
  NAND2_X1 U12837 ( .A1(n14543), .A2(n9866), .ZN(n11665) );
  NAND2_X1 U12838 ( .A1(n10196), .A2(n11547), .ZN(n12236) );
  NAND2_X1 U12839 ( .A1(n11542), .A2(n11543), .ZN(n10196) );
  CLKBUF_X1 U12840 ( .A(n12082), .Z(n10197) );
  AOI21_X1 U12841 ( .B1(n13477), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A(n9818), .ZN(n12368) );
  AOI21_X1 U12842 ( .B1(n13477), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A(n9862), .ZN(n13723) );
  OAI21_X2 U12843 ( .B1(n12357), .B2(n12346), .A(n20010), .ZN(n10203) );
  NAND2_X2 U12844 ( .A1(n9762), .A2(n9797), .ZN(n12469) );
  NAND2_X1 U12845 ( .A1(n12474), .A2(n13971), .ZN(n13427) );
  NOR2_X1 U12846 ( .A1(n10209), .A2(n14219), .ZN(n10205) );
  NOR2_X1 U12847 ( .A1(n10211), .A2(n9814), .ZN(n10212) );
  NAND3_X1 U12848 ( .A1(n10215), .A2(n14200), .A3(n14201), .ZN(n10214) );
  XNOR2_X2 U12849 ( .A(n10216), .B(n10217), .ZN(n20008) );
  AOI21_X2 U12850 ( .B1(n12906), .B2(n12641), .A(n12640), .ZN(n10217) );
  NAND4_X1 U12851 ( .A1(n11193), .A2(n11191), .A3(n11192), .A4(n11190), .ZN(
        n10219) );
  NAND3_X1 U12852 ( .A1(n11162), .A2(n11161), .A3(n11160), .ZN(n10218) );
  NAND3_X1 U12853 ( .A1(n10428), .A2(n10410), .A3(n10869), .ZN(n10220) );
  CLKBUF_X1 U12854 ( .A(n10230), .Z(n10223) );
  NAND2_X1 U12855 ( .A1(n10241), .A2(n9820), .ZN(n10238) );
  CLKBUF_X1 U12856 ( .A(n10245), .Z(n10242) );
  NAND3_X1 U12857 ( .A1(n11297), .A2(n11234), .A3(n11235), .ZN(n11246) );
  INV_X1 U12858 ( .A(n11490), .ZN(n10246) );
  AND2_X2 U12859 ( .A1(n11114), .A2(n11146), .ZN(n11155) );
  NAND2_X1 U12860 ( .A1(n9809), .A2(n10248), .ZN(n11691) );
  NAND2_X1 U12861 ( .A1(n16046), .A2(n16049), .ZN(n11493) );
  NAND2_X1 U12862 ( .A1(n10255), .A2(n10254), .ZN(n16049) );
  NAND2_X1 U12863 ( .A1(n12826), .A2(n10256), .ZN(n10255) );
  NAND2_X1 U12864 ( .A1(n12824), .A2(n16147), .ZN(n10256) );
  NAND2_X1 U12865 ( .A1(n13320), .A2(n13319), .ZN(n13458) );
  AOI22_X1 U12866 ( .A1(n9743), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(n9735), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n10302) );
  INV_X2 U12867 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n12553) );
  OAI21_X2 U12868 ( .B1(n14303), .B2(n14218), .A(n14354), .ZN(n15645) );
  OAI21_X1 U12869 ( .B1(n10479), .B2(n10478), .A(n10494), .ZN(n11985) );
  CLKBUF_X1 U12870 ( .A(n11146), .Z(n15103) );
  NAND2_X1 U12871 ( .A1(n11146), .A2(n11694), .ZN(n10468) );
  NAND2_X1 U12872 ( .A1(n14554), .A2(n9804), .ZN(n10791) );
  NAND2_X1 U12873 ( .A1(n14556), .A2(n14555), .ZN(n14554) );
  NAND2_X1 U12874 ( .A1(n12864), .A2(n20008), .ZN(n20122) );
  OR2_X1 U12875 ( .A1(n20008), .A2(n12866), .ZN(n20462) );
  NAND2_X1 U12876 ( .A1(n11666), .A2(n10275), .ZN(n10430) );
  OR2_X1 U12877 ( .A1(n10482), .A2(n10481), .ZN(n10483) );
  NAND2_X2 U12878 ( .A1(n10481), .A2(n10482), .ZN(n10480) );
  NAND2_X1 U12879 ( .A1(n11121), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n11122) );
  NAND2_X1 U12880 ( .A1(n10472), .A2(n10471), .ZN(n10451) );
  INV_X1 U12881 ( .A(n14106), .ZN(n14113) );
  NAND2_X1 U12882 ( .A1(n13869), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n12110) );
  OR2_X1 U12883 ( .A1(n10750), .A2(n10749), .ZN(n10751) );
  NAND2_X1 U12884 ( .A1(n11113), .A2(n12221), .ZN(n11127) );
  OR2_X1 U12885 ( .A1(n11691), .A2(n19035), .ZN(n11705) );
  AND2_X2 U12886 ( .A1(n19764), .A2(n12476), .ZN(n19938) );
  OR2_X1 U12887 ( .A1(n15339), .A2(n15340), .ZN(n10261) );
  INV_X1 U12888 ( .A(n17200), .ZN(n15220) );
  AND2_X1 U12889 ( .A1(n14312), .A2(n15721), .ZN(n10262) );
  AND2_X1 U12890 ( .A1(n10910), .A2(n10927), .ZN(n10263) );
  INV_X1 U12891 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n15605) );
  AND3_X1 U12892 ( .A1(n20038), .A2(n20042), .A3(n12187), .ZN(n10264) );
  AND2_X1 U12893 ( .A1(n11495), .A2(n11494), .ZN(n10265) );
  INV_X1 U12894 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n12449) );
  AND2_X1 U12895 ( .A1(n10336), .A2(n10335), .ZN(n10266) );
  NAND2_X1 U12896 ( .A1(n9743), .A2(n10359), .ZN(n10267) );
  AND2_X1 U12897 ( .A1(n17585), .A2(n17679), .ZN(n10268) );
  NOR2_X1 U12898 ( .A1(n17390), .A2(n17470), .ZN(n17659) );
  INV_X1 U12899 ( .A(n14602), .ZN(n14582) );
  XNOR2_X1 U12900 ( .A(n11132), .B(n10480), .ZN(n11115) );
  AND2_X1 U12901 ( .A1(n17034), .A2(n18052), .ZN(n17024) );
  OR2_X1 U12902 ( .A1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n10269) );
  INV_X1 U12903 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14221) );
  AND3_X1 U12904 ( .A1(n11107), .A2(n11106), .A3(n11105), .ZN(n10270) );
  OR3_X1 U12905 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(n17398), .ZN(n10271) );
  AND2_X1 U12906 ( .A1(n19840), .A2(n19841), .ZN(n10272) );
  INV_X1 U12907 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n19793) );
  NAND2_X1 U12908 ( .A1(n17387), .A2(n17674), .ZN(n17424) );
  INV_X1 U12909 ( .A(n17424), .ZN(n17390) );
  INV_X2 U12910 ( .A(n18962), .ZN(n19006) );
  NAND2_X1 U12911 ( .A1(n12215), .A2(n12216), .ZN(n12214) );
  OR2_X1 U12912 ( .A1(n18741), .A2(n18743), .ZN(n10273) );
  OR2_X1 U12913 ( .A1(n12532), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n19845) );
  AND2_X1 U12914 ( .A1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P2_STATE2_REG_0__SCAN_IN), .ZN(n10275) );
  AND3_X1 U12915 ( .A1(n14793), .A2(n11392), .A3(n14833), .ZN(n10276) );
  NAND2_X1 U12916 ( .A1(n15955), .A2(n15954), .ZN(n15953) );
  AND2_X1 U12917 ( .A1(n15045), .A2(n15062), .ZN(n10277) );
  INV_X1 U12918 ( .A(n10390), .ZN(n10383) );
  AND2_X1 U12919 ( .A1(n12084), .A2(n12083), .ZN(n10278) );
  INV_X1 U12920 ( .A(n13951), .ZN(n12450) );
  INV_X1 U12921 ( .A(n11204), .ZN(n11150) );
  NAND2_X1 U12922 ( .A1(n11150), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n11151) );
  INV_X1 U12923 ( .A(n12147), .ZN(n11994) );
  AOI21_X1 U12924 ( .B1(n12000), .B2(n11994), .A(n11993), .ZN(n12002) );
  NOR3_X1 U12925 ( .A1(n12180), .A2(n12156), .A3(n13086), .ZN(n12168) );
  NAND2_X1 U12926 ( .A1(n11996), .A2(n11995), .ZN(n12003) );
  OR2_X1 U12927 ( .A1(n13089), .A2(n12708), .ZN(n12721) );
  OR2_X1 U12928 ( .A1(n12734), .A2(n12733), .ZN(n13362) );
  AOI22_X1 U12929 ( .A1(n13188), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n10376), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10337) );
  NAND2_X1 U12930 ( .A1(n10415), .A2(n16176), .ZN(n10395) );
  NAND2_X1 U12931 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n20435), .ZN(
        n12147) );
  BUF_X1 U12932 ( .A(n12374), .Z(n13803) );
  OR2_X1 U12933 ( .A1(n12629), .A2(n12628), .ZN(n12633) );
  OR2_X1 U12934 ( .A1(n13056), .A2(n13055), .ZN(n13371) );
  NOR2_X1 U12935 ( .A1(n12639), .A2(n12638), .ZN(n12640) );
  NAND2_X1 U12936 ( .A1(n12067), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n12068) );
  INV_X1 U12937 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10280) );
  AND2_X2 U12938 ( .A1(n10406), .A2(n10390), .ZN(n10428) );
  AOI22_X1 U12939 ( .A1(n13188), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n10376), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10341) );
  NAND2_X1 U12940 ( .A1(n20034), .A2(n13382), .ZN(n12390) );
  AND4_X1 U12941 ( .A1(n12075), .A2(n12074), .A3(n12073), .A4(n12072), .ZN(
        n12076) );
  INV_X1 U12942 ( .A(n10396), .ZN(n10410) );
  NAND2_X1 U12943 ( .A1(n14734), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11699) );
  NAND2_X1 U12944 ( .A1(n12450), .A2(n12449), .ZN(n12451) );
  AND2_X1 U12945 ( .A1(n12841), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n13820) );
  INV_X1 U12946 ( .A(n12756), .ZN(n12753) );
  INV_X1 U12947 ( .A(n12906), .ZN(n12438) );
  AND2_X1 U12948 ( .A1(n12430), .A2(n12429), .ZN(n12433) );
  OR2_X1 U12949 ( .A1(n12664), .A2(n12663), .ZN(n13352) );
  NAND2_X1 U12950 ( .A1(n11153), .A2(n11694), .ZN(n10476) );
  INV_X1 U12951 ( .A(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n20798) );
  INV_X1 U12952 ( .A(n13690), .ZN(n13734) );
  NAND2_X1 U12953 ( .A1(n12534), .A2(n12533), .ZN(n12535) );
  INV_X1 U12954 ( .A(n13883), .ZN(n13855) );
  OR2_X1 U12955 ( .A1(n13412), .A2(n12504), .ZN(n12505) );
  NAND2_X1 U12956 ( .A1(n13782), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n13817) );
  OR2_X1 U12957 ( .A1(n12341), .A2(n15822), .ZN(n13883) );
  INV_X1 U12958 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n12837) );
  NAND2_X1 U12959 ( .A1(n12754), .A2(n12753), .ZN(n13095) );
  INV_X1 U12960 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20321) );
  NAND2_X1 U12961 ( .A1(n20269), .A2(n15822), .ZN(n12667) );
  INV_X1 U12962 ( .A(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n11697) );
  AND2_X1 U12963 ( .A1(n10564), .A2(n12299), .ZN(n10565) );
  AND2_X1 U12964 ( .A1(n14599), .A2(n10726), .ZN(n10704) );
  OR2_X1 U12965 ( .A1(n15896), .A2(n11425), .ZN(n14921) );
  AND2_X1 U12966 ( .A1(n11619), .A2(n11618), .ZN(n13230) );
  AND2_X1 U12967 ( .A1(n11390), .A2(n14839), .ZN(n14832) );
  NOR2_X1 U12968 ( .A1(n11467), .A2(n10915), .ZN(n16169) );
  NAND2_X1 U12969 ( .A1(n10463), .A2(n19714), .ZN(n10487) );
  INV_X1 U12970 ( .A(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n20836) );
  INV_X1 U12971 ( .A(n18027), .ZN(n15231) );
  NOR2_X1 U12972 ( .A1(n15346), .A2(n15334), .ZN(n15337) );
  AND2_X1 U12973 ( .A1(n14025), .A2(n13958), .ZN(n14004) );
  NOR2_X1 U12974 ( .A1(n13616), .A2(n15568), .ZN(n13621) );
  NAND2_X1 U12975 ( .A1(n13493), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n13572) );
  INV_X1 U12976 ( .A(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n19822) );
  INV_X1 U12977 ( .A(n19861), .ZN(n19823) );
  OR2_X1 U12978 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n13886) );
  NAND2_X1 U12979 ( .A1(n12506), .A2(n12505), .ZN(n12574) );
  AND4_X1 U12980 ( .A1(n12139), .A2(n12138), .A3(n12137), .A4(n12136), .ZN(
        n12140) );
  NOR2_X1 U12981 ( .A1(n13685), .A2(n12839), .ZN(n13654) );
  NAND2_X1 U12982 ( .A1(n14243), .A2(n14221), .ZN(n14223) );
  AND2_X1 U12983 ( .A1(n13919), .A2(n13918), .ZN(n14087) );
  AND2_X1 U12984 ( .A1(n13528), .A2(n13527), .ZN(n14059) );
  AND2_X1 U12985 ( .A1(n13522), .A2(n13521), .ZN(n13535) );
  AND2_X1 U12986 ( .A1(n12765), .A2(n12764), .ZN(n12766) );
  NAND2_X1 U12987 ( .A1(n13440), .A2(n13432), .ZN(n15472) );
  INV_X1 U12988 ( .A(n12806), .ZN(n15430) );
  NOR2_X1 U12989 ( .A1(n20155), .A2(n20057), .ZN(n20328) );
  AND2_X1 U12990 ( .A1(n11614), .A2(n11613), .ZN(n13041) );
  AND2_X1 U12991 ( .A1(n11582), .A2(n11581), .ZN(n12243) );
  AND2_X1 U12992 ( .A1(n11560), .A2(n11559), .ZN(n12264) );
  OR3_X1 U12993 ( .A1(n12967), .A2(n11164), .A3(n15830), .ZN(n18923) );
  INV_X1 U12994 ( .A(n18882), .ZN(n18911) );
  INV_X2 U12995 ( .A(n11561), .ZN(n11659) );
  OR2_X1 U12996 ( .A1(n10530), .A2(n10529), .ZN(n12517) );
  INV_X1 U12997 ( .A(n14616), .ZN(n13394) );
  AND2_X1 U12998 ( .A1(n16119), .A2(n11674), .ZN(n16079) );
  AND2_X1 U12999 ( .A1(n15065), .A2(n11671), .ZN(n16119) );
  INV_X1 U13000 ( .A(n19033), .ZN(n18823) );
  NAND2_X1 U13001 ( .A1(n11440), .A2(n10899), .ZN(n12976) );
  OR2_X1 U13002 ( .A1(n19103), .A2(n19101), .ZN(n19129) );
  INV_X1 U13003 ( .A(n15105), .ZN(n19690) );
  OR2_X1 U13004 ( .A1(n19460), .A2(n19455), .ZN(n19508) );
  INV_X1 U13005 ( .A(n15233), .ZN(n18443) );
  NOR2_X1 U13006 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n16556), .ZN(n16540) );
  NOR2_X1 U13007 ( .A1(P3_EBX_REG_11__SCAN_IN), .A2(n16628), .ZN(n16611) );
  NAND2_X1 U13008 ( .A1(n11846), .A2(n18497), .ZN(n16710) );
  INV_X2 U13009 ( .A(n9793), .ZN(n16975) );
  INV_X1 U13010 ( .A(P3_EBX_REG_4__SCAN_IN), .ZN(n17020) );
  NAND2_X1 U13011 ( .A1(n17043), .A2(n17174), .ZN(n17168) );
  NOR2_X1 U13012 ( .A1(n15274), .A2(n15273), .ZN(n15346) );
  AOI21_X1 U13013 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n17390), .A(
        n18390), .ZN(n17471) );
  NOR2_X1 U13014 ( .A1(n17822), .A2(n17501), .ZN(n17808) );
  INV_X1 U13015 ( .A(n17671), .ZN(n17567) );
  NAND2_X1 U13016 ( .A1(n15377), .A2(n10271), .ZN(n15378) );
  NOR2_X1 U13017 ( .A1(n15329), .A2(n17652), .ZN(n17644) );
  INV_X1 U13018 ( .A(n17989), .ZN(n17928) );
  NOR2_X1 U13019 ( .A1(n11794), .A2(n11793), .ZN(n13564) );
  NAND2_X1 U13020 ( .A1(n13756), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n13779) );
  NAND2_X1 U13021 ( .A1(n13621), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n13685) );
  NOR2_X1 U13022 ( .A1(n13489), .A2(n15605), .ZN(n13459) );
  INV_X1 U13023 ( .A(n19838), .ZN(n19857) );
  AND2_X1 U13024 ( .A1(n20664), .A2(n12848), .ZN(n19856) );
  INV_X1 U13025 ( .A(n15631), .ZN(n19876) );
  OR3_X1 U13026 ( .A1(n13419), .A2(n19757), .A3(n12538), .ZN(n12338) );
  INV_X1 U13027 ( .A(n14191), .ZN(n14194) );
  NAND2_X1 U13028 ( .A1(n12574), .A2(n13421), .ZN(n12509) );
  INV_X1 U13029 ( .A(n13150), .ZN(n19912) );
  INV_X1 U13030 ( .A(n13150), .ZN(n19932) );
  INV_X1 U13031 ( .A(n13149), .ZN(n19935) );
  NAND2_X1 U13032 ( .A1(n13689), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n13690) );
  NAND2_X1 U13033 ( .A1(n13444), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n13489) );
  NAND2_X1 U13034 ( .A1(n13091), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n13129) );
  NOR2_X1 U13035 ( .A1(n15726), .A2(n14388), .ZN(n15703) );
  OR2_X1 U13036 ( .A1(n19996), .A2(n19998), .ZN(n19988) );
  INV_X1 U13037 ( .A(n19964), .ZN(n19994) );
  INV_X1 U13038 ( .A(n20161), .ZN(n20057) );
  INV_X1 U13039 ( .A(n20076), .ZN(n20079) );
  OAI21_X1 U13040 ( .B1(n20178), .B2(n20162), .A(n20473), .ZN(n20180) );
  OR2_X1 U13041 ( .A1(n9751), .A2(n20400), .ZN(n20267) );
  INV_X1 U13042 ( .A(n20266), .ZN(n20255) );
  INV_X1 U13043 ( .A(n20366), .ZN(n20316) );
  OAI22_X1 U13044 ( .A1(n20413), .A2(n20412), .B1(n20466), .B2(n20411), .ZN(
        n20429) );
  NOR2_X2 U13045 ( .A1(n20401), .A2(n20400), .ZN(n20458) );
  INV_X1 U13046 ( .A(n20468), .ZN(n20506) );
  NOR2_X2 U13047 ( .A1(n20462), .A2(n20376), .ZN(n20571) );
  INV_X2 U13048 ( .A(n19740), .ZN(n16176) );
  AND2_X1 U13049 ( .A1(n16198), .A2(n12963), .ZN(n18917) );
  OR2_X1 U13050 ( .A1(n10575), .A2(n10574), .ZN(n12898) );
  OR2_X1 U13051 ( .A1(n10562), .A2(n10561), .ZN(n12284) );
  OR2_X1 U13052 ( .A1(n12216), .A2(n12215), .ZN(n12217) );
  OR2_X1 U13053 ( .A1(n15928), .A2(n18930), .ZN(n18944) );
  INV_X1 U13054 ( .A(n18948), .ZN(n18934) );
  INV_X1 U13055 ( .A(n11882), .ZN(n19028) );
  INV_X1 U13056 ( .A(n15006), .ZN(n18761) );
  AND2_X1 U13057 ( .A1(n16064), .A2(n11925), .ZN(n16054) );
  AND2_X1 U13058 ( .A1(n11668), .A2(n11523), .ZN(n19059) );
  XNOR2_X1 U13059 ( .A(n11985), .B(n11984), .ZN(n13215) );
  NOR2_X2 U13060 ( .A1(n19302), .A2(n19199), .ZN(n19131) );
  INV_X1 U13061 ( .A(n19194), .ZN(n19186) );
  OR2_X1 U13062 ( .A1(n13215), .A2(n19707), .ZN(n19686) );
  INV_X1 U13063 ( .A(n19254), .ZN(n19247) );
  AND2_X1 U13064 ( .A1(n19225), .A2(n19459), .ZN(n19280) );
  NOR2_X1 U13065 ( .A1(n13214), .A2(n19199), .ZN(n19297) );
  AND2_X1 U13066 ( .A1(n19225), .A2(n19553), .ZN(n19329) );
  INV_X1 U13067 ( .A(n19362), .ZN(n19363) );
  AND2_X1 U13068 ( .A1(n13005), .A2(n13004), .ZN(n19414) );
  OAI21_X1 U13069 ( .B1(n19445), .B2(n19714), .A(n19430), .ZN(n19447) );
  NOR2_X1 U13070 ( .A1(n19424), .A2(n19423), .ZN(n19451) );
  INV_X1 U13071 ( .A(n19576), .ZN(n19522) );
  INV_X1 U13072 ( .A(n19549), .ZN(n19426) );
  AND2_X1 U13073 ( .A1(n10391), .A2(n19076), .ZN(n19565) );
  NOR2_X1 U13074 ( .A1(n15105), .A2(n19716), .ZN(n19334) );
  XNOR2_X1 U13075 ( .A(n18654), .B(n16694), .ZN(n18657) );
  OAI211_X1 U13076 ( .C1(n13562), .C2(n13561), .A(n13560), .B(n13559), .ZN(
        n18448) );
  NOR2_X1 U13077 ( .A1(P3_EBX_REG_15__SCAN_IN), .A2(n16578), .ZN(n16560) );
  NOR2_X1 U13078 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(n16602), .ZN(n16590) );
  NOR2_X1 U13079 ( .A1(P3_EBX_REG_9__SCAN_IN), .A2(n16649), .ZN(n16631) );
  INV_X1 U13080 ( .A(n16710), .ZN(n16739) );
  NAND2_X1 U13081 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n16822), .ZN(n16816) );
  NAND2_X1 U13082 ( .A1(P3_EBX_REG_15__SCAN_IN), .A2(n9763), .ZN(n16902) );
  NOR2_X1 U13083 ( .A1(n17266), .A2(n17068), .ZN(n17060) );
  NOR2_X1 U13084 ( .A1(n18052), .A2(n17087), .ZN(n17083) );
  NOR3_X1 U13085 ( .A1(n18052), .A2(n17124), .A3(n17245), .ZN(n17113) );
  NOR2_X1 U13086 ( .A1(n17284), .A2(n17168), .ZN(n17167) );
  INV_X1 U13087 ( .A(n17185), .ZN(n17180) );
  OAI211_X1 U13088 ( .C1(n18654), .C2(n18655), .A(n17241), .B(n17240), .ZN(
        n17300) );
  INV_X1 U13089 ( .A(n18057), .ZN(n18390) );
  INV_X1 U13090 ( .A(n17493), .ZN(n17586) );
  NOR2_X2 U13091 ( .A1(n18610), .A2(n17567), .ZN(n17470) );
  NOR2_X1 U13092 ( .A1(n16218), .A2(n16208), .ZN(n17664) );
  NOR3_X1 U13093 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17307), .A3(
        n16281), .ZN(n16283) );
  NAND2_X1 U13094 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n17495), .ZN(
        n17494) );
  NOR2_X1 U13095 ( .A1(n17995), .A2(n17989), .ZN(n17918) );
  NOR2_X1 U13096 ( .A1(n17972), .A2(n17928), .ZN(n17982) );
  INV_X1 U13097 ( .A(n18362), .ZN(n18054) );
  NOR2_X1 U13098 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18599), .ZN(
        n18626) );
  INV_X1 U13099 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n18666) );
  INV_X1 U13100 ( .A(P3_STATE_REG_1__SCAN_IN), .ZN(n20812) );
  INV_X1 U13101 ( .A(U212), .ZN(n16332) );
  OR2_X1 U13102 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n19755), .ZN(n20662) );
  INV_X1 U13103 ( .A(n19816), .ZN(n15589) );
  INV_X1 U13104 ( .A(n19856), .ZN(n19836) );
  INV_X1 U13105 ( .A(n19850), .ZN(n19870) );
  NAND2_X1 U13106 ( .A1(n19879), .A2(n12539), .ZN(n15631) );
  NAND2_X1 U13107 ( .A1(n19885), .A2(n9725), .ZN(n12616) );
  INV_X1 U13108 ( .A(n19885), .ZN(n19905) );
  NOR2_X1 U13109 ( .A1(n13904), .A2(n12592), .ZN(n13150) );
  INV_X1 U13110 ( .A(n19993), .ZN(n15807) );
  INV_X1 U13111 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20435) );
  OR2_X1 U13112 ( .A1(n20122), .A2(n20267), .ZN(n20076) );
  OR2_X1 U13113 ( .A1(n20122), .A2(n20434), .ZN(n20117) );
  OR2_X1 U13114 ( .A1(n20122), .A2(n20463), .ZN(n20149) );
  OR2_X1 U13115 ( .A1(n20122), .A2(n20376), .ZN(n20183) );
  OR2_X1 U13116 ( .A1(n20239), .A2(n20267), .ZN(n20203) );
  OR2_X1 U13117 ( .A1(n20239), .A2(n20434), .ZN(n20238) );
  OR2_X1 U13118 ( .A1(n20239), .A2(n20376), .ZN(n20258) );
  OR2_X1 U13119 ( .A1(n20239), .A2(n20463), .ZN(n20266) );
  NAND2_X1 U13120 ( .A1(n20371), .A2(n20268), .ZN(n20320) );
  OR2_X1 U13121 ( .A1(n20377), .A2(n20434), .ZN(n20366) );
  OR2_X1 U13122 ( .A1(n20377), .A2(n20463), .ZN(n20391) );
  OR2_X1 U13123 ( .A1(n20377), .A2(n20376), .ZN(n20433) );
  OR2_X1 U13124 ( .A1(n20462), .A2(n20434), .ZN(n20468) );
  NAND2_X1 U13125 ( .A1(n20519), .A2(n20464), .ZN(n20575) );
  INV_X1 U13126 ( .A(n20654), .ZN(n20580) );
  INV_X1 U13127 ( .A(n18917), .ZN(n18898) );
  INV_X1 U13128 ( .A(n11712), .ZN(n11713) );
  AND2_X1 U13129 ( .A1(n11708), .A2(n18949), .ZN(n14621) );
  NAND2_X1 U13130 ( .A1(n12214), .A2(n12217), .ZN(n15105) );
  INV_X1 U13131 ( .A(n18944), .ZN(n18937) );
  NAND2_X1 U13132 ( .A1(n19019), .A2(n18956), .ZN(n18962) );
  NAND2_X1 U13133 ( .A1(n18953), .A2(n19741), .ZN(n19019) );
  OR2_X1 U13134 ( .A1(n11692), .A2(n10944), .ZN(n19035) );
  INV_X1 U13135 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n16006) );
  INV_X1 U13136 ( .A(n16060), .ZN(n19037) );
  INV_X1 U13137 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n16052) );
  INV_X1 U13138 ( .A(n19041), .ZN(n16058) );
  INV_X1 U13139 ( .A(n16157), .ZN(n19056) );
  INV_X1 U13140 ( .A(n19065), .ZN(n16139) );
  INV_X1 U13141 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19722) );
  AOI21_X1 U13142 ( .B1(n13082), .B2(n13081), .A(n13080), .ZN(n19095) );
  NAND2_X1 U13143 ( .A1(n19338), .A2(n19225), .ZN(n19153) );
  OR2_X1 U13144 ( .A1(n19199), .A2(n19686), .ZN(n19194) );
  INV_X1 U13145 ( .A(n19216), .ZN(n19224) );
  OR2_X1 U13146 ( .A1(n19199), .A2(n19423), .ZN(n19254) );
  INV_X1 U13147 ( .A(n19280), .ZN(n19275) );
  INV_X1 U13148 ( .A(n19297), .ZN(n19295) );
  INV_X1 U13149 ( .A(n19292), .ZN(n19301) );
  INV_X1 U13150 ( .A(n19329), .ZN(n19325) );
  OR2_X1 U13151 ( .A1(n19424), .A2(n19302), .ZN(n19362) );
  INV_X1 U13152 ( .A(n19395), .ZN(n19390) );
  NAND2_X1 U13153 ( .A1(n19334), .A2(n19162), .ZN(n19450) );
  INV_X1 U13154 ( .A(n19451), .ZN(n19513) );
  INV_X1 U13155 ( .A(n19525), .ZN(n19582) );
  NAND2_X1 U13156 ( .A1(n19334), .A2(n19553), .ZN(n19604) );
  INV_X1 U13157 ( .A(n18657), .ZN(n18668) );
  NAND2_X1 U13158 ( .A1(n18648), .A2(n18450), .ZN(n16381) );
  INV_X1 U13159 ( .A(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n17498) );
  INV_X1 U13160 ( .A(n16681), .ZN(n16743) );
  INV_X1 U13161 ( .A(n16709), .ZN(n16740) );
  NOR2_X1 U13162 ( .A1(n16764), .A2(n16763), .ZN(n16791) );
  INV_X1 U13163 ( .A(n15343), .ZN(n17171) );
  INV_X1 U13164 ( .A(n17188), .ZN(n17198) );
  INV_X1 U13165 ( .A(n17218), .ZN(n17237) );
  INV_X1 U13166 ( .A(n17470), .ZN(n17521) );
  NAND2_X1 U13167 ( .A1(n17664), .A2(n16273), .ZN(n17493) );
  AOI22_X1 U13168 ( .A1(n17667), .A2(n17868), .B1(n17587), .B2(n17874), .ZN(
        n17574) );
  OAI21_X1 U13169 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n18647), .A(n16381), 
        .ZN(n17674) );
  NOR2_X1 U13170 ( .A1(n17646), .A2(n17629), .ZN(n17671) );
  INV_X1 U13171 ( .A(n17993), .ZN(n17979) );
  INV_X1 U13172 ( .A(n17918), .ZN(n17980) );
  INV_X1 U13173 ( .A(n17982), .ZN(n17999) );
  INV_X1 U13174 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n18599) );
  INV_X1 U13175 ( .A(n18595), .ZN(n18516) );
  NAND2_X1 U13176 ( .A1(P3_STATE_REG_2__SCAN_IN), .A2(n18665), .ZN(n18587) );
  INV_X1 U13177 ( .A(n16339), .ZN(n16329) );
  CLKBUF_X1 U13178 ( .A(n16373), .Z(n20676) );
  AOI22_X1 U13179 ( .A1(n9746), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n10375), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10279) );
  AND2_X2 U13180 ( .A1(n10280), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10509) );
  AND2_X4 U13181 ( .A1(n10509), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10499) );
  AND2_X4 U13182 ( .A1(n10508), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10833) );
  AOI22_X1 U13183 ( .A1(n9745), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n10833), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10282) );
  NAND3_X1 U13184 ( .A1(n10283), .A2(n10282), .A3(n10281), .ZN(n10284) );
  AOI22_X1 U13185 ( .A1(n9747), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(n9753), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10290) );
  AOI22_X1 U13186 ( .A1(n9745), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n10833), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10289) );
  AOI22_X1 U13187 ( .A1(n10672), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n10500), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10288) );
  AOI22_X1 U13188 ( .A1(n9743), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n10376), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10287) );
  NAND4_X1 U13189 ( .A1(n10290), .A2(n10289), .A3(n10288), .A4(n10287), .ZN(
        n10291) );
  NAND2_X1 U13190 ( .A1(n10291), .A2(n10359), .ZN(n10292) );
  AOI22_X1 U13191 ( .A1(n13188), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n9735), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10297) );
  AOI22_X1 U13192 ( .A1(n9744), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n10833), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n10296) );
  AOI22_X1 U13193 ( .A1(n9748), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(n9734), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n10295) );
  AOI22_X1 U13194 ( .A1(n10672), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n9752), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n10294) );
  NAND4_X1 U13195 ( .A1(n10297), .A2(n10296), .A3(n10295), .A4(n10294), .ZN(
        n10298) );
  NAND2_X1 U13196 ( .A1(n10298), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10305) );
  AOI22_X1 U13197 ( .A1(n9731), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n10833), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10301) );
  AOI22_X1 U13198 ( .A1(n10672), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n9734), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10300) );
  AOI22_X1 U13199 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n9746), .B1(n9753), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10299) );
  NAND4_X1 U13200 ( .A1(n10302), .A2(n10301), .A3(n10300), .A4(n10299), .ZN(
        n10303) );
  NAND2_X1 U13201 ( .A1(n10303), .A2(n10359), .ZN(n10304) );
  NAND2_X4 U13202 ( .A1(n10305), .A2(n10304), .ZN(n10390) );
  AND2_X2 U13203 ( .A1(n10389), .A2(n10390), .ZN(n10401) );
  AOI22_X1 U13204 ( .A1(n9746), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n10375), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10309) );
  AOI22_X1 U13205 ( .A1(n9744), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n10833), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10308) );
  AOI22_X1 U13206 ( .A1(n10672), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n10500), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10307) );
  AOI22_X1 U13207 ( .A1(n9743), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n9735), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10306) );
  NAND4_X1 U13208 ( .A1(n10309), .A2(n10308), .A3(n10307), .A4(n10306), .ZN(
        n10310) );
  NAND2_X1 U13209 ( .A1(n10310), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10317) );
  AOI22_X1 U13210 ( .A1(n9747), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n10375), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10314) );
  AOI22_X1 U13211 ( .A1(n10499), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n10833), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10313) );
  AOI22_X1 U13212 ( .A1(n10672), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n9734), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10312) );
  AOI22_X1 U13213 ( .A1(n13188), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n9735), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10311) );
  NAND4_X1 U13214 ( .A1(n10314), .A2(n10313), .A3(n10312), .A4(n10311), .ZN(
        n10315) );
  AOI22_X1 U13215 ( .A1(n9743), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n10376), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10321) );
  AOI22_X1 U13216 ( .A1(n10672), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n10500), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10320) );
  AOI22_X1 U13217 ( .A1(n9744), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n10833), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10319) );
  AOI22_X1 U13218 ( .A1(n9746), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(n9753), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10318) );
  NAND4_X1 U13219 ( .A1(n10321), .A2(n10320), .A3(n10319), .A4(n10318), .ZN(
        n10322) );
  NAND2_X1 U13220 ( .A1(n10322), .A2(n10359), .ZN(n10329) );
  AOI22_X1 U13221 ( .A1(n9743), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n9735), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10326) );
  AOI22_X1 U13222 ( .A1(n10499), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n10833), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10325) );
  AOI22_X1 U13223 ( .A1(n9747), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(n9752), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10324) );
  AOI22_X1 U13224 ( .A1(n10672), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n10500), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n10323) );
  NAND4_X1 U13225 ( .A1(n10326), .A2(n10325), .A3(n10324), .A4(n10323), .ZN(
        n10327) );
  NAND2_X1 U13226 ( .A1(n10327), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10328) );
  NOR2_X1 U13227 ( .A1(n10391), .A2(n19077), .ZN(n10330) );
  AOI22_X1 U13228 ( .A1(n9753), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(n9734), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10333) );
  AOI22_X1 U13229 ( .A1(n10672), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n9748), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10332) );
  AOI22_X1 U13230 ( .A1(n9731), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10833), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10331) );
  AOI22_X1 U13231 ( .A1(n9744), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n9748), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10336) );
  AOI22_X1 U13232 ( .A1(n9753), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(n9734), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10335) );
  AOI22_X1 U13233 ( .A1(n10672), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n10833), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10338) );
  AOI22_X1 U13234 ( .A1(n10499), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n10833), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10342) );
  AOI22_X1 U13235 ( .A1(n10672), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n9733), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10344) );
  AOI22_X1 U13236 ( .A1(n9747), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(n9752), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10343) );
  AOI22_X1 U13237 ( .A1(n10499), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n10833), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10348) );
  AOI22_X1 U13238 ( .A1(n9748), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(n9752), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10347) );
  AOI22_X1 U13239 ( .A1(n9743), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n10376), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10350) );
  AOI22_X1 U13240 ( .A1(n10672), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n9734), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10349) );
  NAND2_X2 U13241 ( .A1(n10368), .A2(n10393), .ZN(n11451) );
  AOI22_X1 U13242 ( .A1(n10672), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n9746), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10358) );
  AOI22_X1 U13243 ( .A1(n9752), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n10500), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10357) );
  AOI22_X1 U13244 ( .A1(n10499), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n10833), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10356) );
  NAND4_X1 U13245 ( .A1(n10358), .A2(n10357), .A3(n10356), .A4(n10355), .ZN(
        n10360) );
  NAND2_X1 U13246 ( .A1(n10360), .A2(n10359), .ZN(n10367) );
  AOI22_X1 U13247 ( .A1(n10672), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n9747), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10364) );
  AOI22_X1 U13248 ( .A1(n9731), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n10833), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10363) );
  AOI22_X1 U13249 ( .A1(n10375), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n9733), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10362) );
  NAND4_X1 U13250 ( .A1(n10364), .A2(n10363), .A3(n10362), .A4(n10361), .ZN(
        n10365) );
  NAND2_X1 U13251 ( .A1(n10365), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10366) );
  NAND2_X1 U13252 ( .A1(n11451), .A2(n10263), .ZN(n10370) );
  NAND2_X1 U13253 ( .A1(n10370), .A2(n10369), .ZN(n11522) );
  AOI22_X1 U13254 ( .A1(n10672), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n9748), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10374) );
  AOI22_X1 U13255 ( .A1(n10499), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10833), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10373) );
  AOI22_X1 U13256 ( .A1(n9752), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n10500), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10372) );
  AOI22_X1 U13257 ( .A1(n13188), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n9735), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10371) );
  NAND4_X1 U13258 ( .A1(n10374), .A2(n10373), .A3(n10372), .A4(n10371), .ZN(
        n10382) );
  AOI22_X1 U13259 ( .A1(n10499), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10833), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10380) );
  AOI22_X1 U13260 ( .A1(n10672), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n9752), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10379) );
  AOI22_X1 U13261 ( .A1(n9746), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(n9733), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10378) );
  AOI22_X1 U13262 ( .A1(n9743), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n9735), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10377) );
  NAND4_X1 U13263 ( .A1(n10380), .A2(n10379), .A3(n10378), .A4(n10377), .ZN(
        n10381) );
  INV_X2 U13264 ( .A(n10398), .ZN(n10909) );
  NAND3_X1 U13265 ( .A1(n10397), .A2(n10909), .A3(n10390), .ZN(n10386) );
  NAND2_X1 U13266 ( .A1(n10385), .A2(n10386), .ZN(n10388) );
  NAND2_X1 U13267 ( .A1(n10908), .A2(n10389), .ZN(n10387) );
  NAND3_X1 U13268 ( .A1(n10388), .A2(n10387), .A3(n10910), .ZN(n10394) );
  AND2_X1 U13269 ( .A1(n10391), .A2(n10398), .ZN(n10392) );
  NAND3_X1 U13270 ( .A1(n10394), .A2(n16176), .A3(n10424), .ZN(n11530) );
  INV_X1 U13271 ( .A(n10417), .ZN(n10405) );
  NAND2_X1 U13272 ( .A1(n10902), .A2(n10398), .ZN(n10400) );
  NAND2_X1 U13273 ( .A1(n10403), .A2(n10407), .ZN(n10404) );
  INV_X1 U13274 ( .A(n10908), .ZN(n11965) );
  NAND2_X1 U13275 ( .A1(n11965), .A2(n10401), .ZN(n10411) );
  OAI21_X1 U13276 ( .B1(n10927), .B2(n19740), .A(n10869), .ZN(n11526) );
  NAND2_X2 U13277 ( .A1(n10412), .A2(n11519), .ZN(n15092) );
  NOR2_X1 U13278 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n19734) );
  NAND2_X1 U13279 ( .A1(n19734), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n10413) );
  NAND2_X1 U13280 ( .A1(n10414), .A2(n10413), .ZN(n10481) );
  NOR2_X1 U13281 ( .A1(n10917), .A2(n10416), .ZN(n11524) );
  NOR2_X1 U13282 ( .A1(n11524), .A2(n10417), .ZN(n10432) );
  INV_X1 U13283 ( .A(n10425), .ZN(n10419) );
  INV_X1 U13284 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n10947) );
  NAND2_X1 U13285 ( .A1(n10456), .A2(P2_EBX_REG_0__SCAN_IN), .ZN(n10422) );
  AND2_X1 U13286 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n10420) );
  NOR2_X1 U13287 ( .A1(n19734), .A2(n10420), .ZN(n10421) );
  OAI211_X1 U13288 ( .C1(n11548), .C2(n10947), .A(n10422), .B(n10421), .ZN(
        n10423) );
  INV_X1 U13289 ( .A(n10423), .ZN(n10431) );
  INV_X4 U13290 ( .A(n10927), .ZN(n11164) );
  NAND2_X1 U13291 ( .A1(n10436), .A2(n11164), .ZN(n10429) );
  NAND2_X2 U13292 ( .A1(n10429), .A2(n15092), .ZN(n11666) );
  INV_X1 U13293 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n13175) );
  NAND2_X1 U13294 ( .A1(n10456), .A2(P2_EBX_REG_1__SCAN_IN), .ZN(n10434) );
  NAND2_X1 U13295 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n10433) );
  AOI22_X1 U13296 ( .A1(n10436), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(n19734), 
        .B2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n10437) );
  OAI21_X2 U13297 ( .B1(n10480), .B2(n9788), .A(n10486), .ZN(n10439) );
  NAND2_X1 U13298 ( .A1(n10480), .A2(n9788), .ZN(n10438) );
  NAND2_X1 U13299 ( .A1(n10452), .A2(n16164), .ZN(n10441) );
  AOI21_X1 U13300 ( .B1(n18954), .B2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n10440) );
  INV_X1 U13301 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n19067) );
  INV_X1 U13302 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n11958) );
  NAND2_X1 U13303 ( .A1(n10456), .A2(P2_EBX_REG_2__SCAN_IN), .ZN(n10443) );
  NAND2_X1 U13304 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n10442) );
  OAI211_X1 U13305 ( .C1(n11548), .C2(n11958), .A(n10443), .B(n10442), .ZN(
        n10444) );
  INV_X1 U13306 ( .A(n10444), .ZN(n10445) );
  INV_X1 U13307 ( .A(n10446), .ZN(n10448) );
  XNOR2_X2 U13308 ( .A(n10447), .B(n10448), .ZN(n10471) );
  INV_X1 U13309 ( .A(n10447), .ZN(n10449) );
  NAND2_X1 U13310 ( .A1(n10449), .A2(n10448), .ZN(n10450) );
  NAND2_X1 U13311 ( .A1(n10452), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10454) );
  NAND2_X1 U13312 ( .A1(n19734), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n10453) );
  INV_X1 U13313 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n12927) );
  INV_X1 U13314 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n11002) );
  NAND2_X1 U13315 ( .A1(n10456), .A2(P2_EBX_REG_3__SCAN_IN), .ZN(n10458) );
  NAND2_X1 U13316 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n10457) );
  OAI211_X1 U13317 ( .C1(n11548), .C2(n11002), .A(n10458), .B(n10457), .ZN(
        n10459) );
  INV_X1 U13318 ( .A(n10459), .ZN(n10460) );
  BUF_X4 U13319 ( .A(n10462), .Z(n11146) );
  NAND2_X1 U13320 ( .A1(n10427), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10463) );
  NAND2_X1 U13321 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19544) );
  INV_X1 U13322 ( .A(n19544), .ZN(n10464) );
  NAND2_X1 U13323 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n10464), .ZN(
        n13072) );
  NAND2_X1 U13324 ( .A1(n13072), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n10465) );
  NOR2_X1 U13325 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19544), .ZN(
        n12981) );
  NAND2_X1 U13326 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n12981), .ZN(
        n12985) );
  NAND2_X1 U13327 ( .A1(n10465), .A2(n12985), .ZN(n10466) );
  AOI22_X1 U13328 ( .A1(n10487), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n19685), .B2(n10466), .ZN(n10467) );
  INV_X1 U13329 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11169) );
  NOR2_X1 U13330 ( .A1(n10788), .A2(n11169), .ZN(n10469) );
  NAND2_X1 U13331 ( .A1(n10497), .A2(n10469), .ZN(n12231) );
  XNOR2_X2 U13332 ( .A(n10472), .B(n10471), .ZN(n11113) );
  INV_X1 U13333 ( .A(n19685), .ZN(n19337) );
  NAND2_X1 U13334 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19163) );
  NAND2_X1 U13335 ( .A1(n19163), .A2(n19704), .ZN(n10473) );
  NAND2_X1 U13336 ( .A1(n10473), .A2(n13072), .ZN(n19196) );
  NOR2_X1 U13337 ( .A1(n19337), .A2(n19196), .ZN(n10474) );
  AOI21_X1 U13338 ( .B1(n10487), .B2(n16164), .A(n10474), .ZN(n10475) );
  INV_X1 U13339 ( .A(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10477) );
  NOR2_X1 U13340 ( .A1(n10788), .A2(n10477), .ZN(n10478) );
  AOI22_X1 U13341 ( .A1(n10487), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n19685), .B2(n19722), .ZN(n10484) );
  NAND2_X1 U13342 ( .A1(n10744), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n10490) );
  NAND2_X1 U13343 ( .A1(n10487), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10488) );
  NAND2_X1 U13344 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n10862), .ZN(
        n19336) );
  NAND2_X1 U13345 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19722), .ZN(
        n19368) );
  NAND2_X1 U13346 ( .A1(n19336), .A2(n19368), .ZN(n19195) );
  NAND2_X1 U13347 ( .A1(n19685), .A2(n19195), .ZN(n19371) );
  NAND2_X1 U13348 ( .A1(n10488), .A2(n19371), .ZN(n10489) );
  NAND2_X1 U13349 ( .A1(n12202), .A2(n12201), .ZN(n10493) );
  INV_X1 U13350 ( .A(n15077), .ZN(n10491) );
  NAND2_X1 U13351 ( .A1(n10491), .A2(n10490), .ZN(n10492) );
  NAND2_X1 U13352 ( .A1(n10427), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n10496) );
  AOI22_X1 U13353 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n10542), .B1(
        n9723), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10505) );
  AND2_X2 U13354 ( .A1(n10672), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10600) );
  INV_X1 U13355 ( .A(n10500), .ZN(n10673) );
  AOI22_X1 U13356 ( .A1(n10600), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n10517), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10504) );
  AND2_X2 U13357 ( .A1(n9747), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10949) );
  AND2_X2 U13358 ( .A1(n9752), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10651) );
  AOI22_X1 U13359 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n10949), .B1(
        n10651), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10503) );
  AOI22_X1 U13360 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n10576), .B1(
        n11008), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10502) );
  NAND4_X1 U13361 ( .A1(n10505), .A2(n10504), .A3(n10503), .A4(n10502), .ZN(
        n10516) );
  AOI22_X1 U13362 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n10581), .B1(
        n10935), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10514) );
  AND2_X2 U13363 ( .A1(n13188), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10593) );
  AOI22_X1 U13364 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n10522), .B1(
        n10593), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10513) );
  AND2_X2 U13365 ( .A1(n10674), .A2(n10507), .ZN(n10954) );
  AOI22_X1 U13366 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n10954), .B1(
        n10523), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10512) );
  AOI22_X1 U13367 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n10524), .B1(
        n10535), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10511) );
  NAND4_X1 U13368 ( .A1(n10514), .A2(n10513), .A3(n10512), .A4(n10511), .ZN(
        n10515) );
  AOI22_X1 U13369 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n10542), .B1(
        n9723), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10521) );
  AOI22_X1 U13370 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n10949), .B1(
        n10651), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n10520) );
  AOI22_X1 U13371 ( .A1(n10600), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n10517), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10519) );
  AOI22_X1 U13372 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n10576), .B1(
        n11008), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10518) );
  NAND4_X1 U13373 ( .A1(n10521), .A2(n10520), .A3(n10519), .A4(n10518), .ZN(
        n10530) );
  AOI22_X1 U13374 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n10581), .B1(
        n10935), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10528) );
  AOI22_X1 U13375 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n10593), .B1(
        n10522), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10527) );
  AOI22_X1 U13376 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n10954), .B1(
        n10523), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10526) );
  AOI22_X1 U13377 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n10535), .B1(
        n10524), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10525) );
  NAND4_X1 U13378 ( .A1(n10528), .A2(n10527), .A3(n10526), .A4(n10525), .ZN(
        n10529) );
  AND2_X1 U13379 ( .A1(n12518), .A2(n12517), .ZN(n10564) );
  AOI22_X1 U13380 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n10600), .B1(
        n10949), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10534) );
  AOI22_X1 U13381 ( .A1(n10542), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n10651), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10533) );
  AOI22_X1 U13382 ( .A1(n9723), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n10517), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10532) );
  AOI22_X1 U13383 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n10593), .B1(
        n10576), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10531) );
  NAND4_X1 U13384 ( .A1(n10534), .A2(n10533), .A3(n10532), .A4(n10531), .ZN(
        n10541) );
  AOI22_X1 U13385 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n10581), .B1(
        n10935), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10539) );
  INV_X2 U13386 ( .A(n10267), .ZN(n11008) );
  AOI22_X1 U13387 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n11008), .B1(
        n10522), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10538) );
  AOI22_X1 U13388 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n10954), .B1(
        n10523), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10537) );
  AOI22_X1 U13389 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n10535), .B1(
        n10524), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10536) );
  NAND4_X1 U13390 ( .A1(n10539), .A2(n10538), .A3(n10537), .A4(n10536), .ZN(
        n10540) );
  INV_X1 U13391 ( .A(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n20859) );
  AOI22_X1 U13392 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n9723), .B1(
        n10542), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10546) );
  AOI22_X1 U13393 ( .A1(n10600), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n10517), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10545) );
  AOI22_X1 U13394 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n10949), .B1(
        n10651), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10544) );
  AOI22_X1 U13395 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n10576), .B1(
        n11008), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10543) );
  NAND4_X1 U13396 ( .A1(n10546), .A2(n10545), .A3(n10544), .A4(n10543), .ZN(
        n10552) );
  AOI22_X1 U13397 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n10581), .B1(
        n10935), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10550) );
  AOI22_X1 U13398 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n10593), .B1(
        n10522), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10549) );
  AOI22_X1 U13399 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n10954), .B1(
        n10523), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10548) );
  AOI22_X1 U13400 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n10524), .B1(
        n10535), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10547) );
  NAND4_X1 U13401 ( .A1(n10550), .A2(n10549), .A3(n10548), .A4(n10547), .ZN(
        n10551) );
  NOR2_X1 U13402 ( .A1(n10552), .A2(n10551), .ZN(n12242) );
  INV_X1 U13403 ( .A(n12242), .ZN(n11056) );
  AOI22_X1 U13404 ( .A1(n9723), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n10600), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10556) );
  AOI22_X1 U13405 ( .A1(n10542), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n10517), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10555) );
  AOI22_X1 U13406 ( .A1(n10949), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n10651), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10554) );
  AOI22_X1 U13407 ( .A1(n10522), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n10576), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10553) );
  NAND4_X1 U13408 ( .A1(n10556), .A2(n10555), .A3(n10554), .A4(n10553), .ZN(
        n10562) );
  AOI22_X1 U13409 ( .A1(n10935), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n10581), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10560) );
  AOI22_X1 U13410 ( .A1(n11008), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10593), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10559) );
  AOI22_X1 U13411 ( .A1(n10954), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10523), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10558) );
  AOI22_X1 U13412 ( .A1(n10535), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n10524), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10557) );
  NAND4_X1 U13413 ( .A1(n10560), .A2(n10559), .A3(n10558), .A4(n10557), .ZN(
        n10561) );
  INV_X1 U13414 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10838) );
  NAND2_X1 U13415 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12271) );
  NOR2_X1 U13416 ( .A1(n10838), .A2(n12271), .ZN(n12281) );
  AND2_X1 U13417 ( .A1(n12284), .A2(n12281), .ZN(n10563) );
  INV_X1 U13418 ( .A(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10773) );
  NOR2_X1 U13419 ( .A1(n10788), .A2(n10773), .ZN(n12280) );
  AND2_X1 U13420 ( .A1(n10563), .A2(n12280), .ZN(n12241) );
  AOI22_X1 U13421 ( .A1(n9723), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n10542), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10569) );
  AOI22_X1 U13422 ( .A1(n10600), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n10517), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10568) );
  AOI22_X1 U13423 ( .A1(n10949), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n10651), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10567) );
  AOI22_X1 U13424 ( .A1(n11008), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10576), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10566) );
  NAND4_X1 U13425 ( .A1(n10569), .A2(n10568), .A3(n10567), .A4(n10566), .ZN(
        n10575) );
  AOI22_X1 U13426 ( .A1(n10935), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n10581), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10573) );
  AOI22_X1 U13427 ( .A1(n10522), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10593), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10572) );
  AOI22_X1 U13428 ( .A1(n10954), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10523), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10571) );
  AOI22_X1 U13429 ( .A1(n10535), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10524), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10570) );
  NAND4_X1 U13430 ( .A1(n10573), .A2(n10572), .A3(n10571), .A4(n10570), .ZN(
        n10574) );
  AOI22_X1 U13431 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n10542), .B1(
        n10651), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10580) );
  AOI22_X1 U13432 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n9723), .B1(
        n10949), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10579) );
  AOI22_X1 U13433 ( .A1(n10600), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n10517), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10578) );
  AOI22_X1 U13434 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n10593), .B1(
        n10576), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10577) );
  NAND4_X1 U13435 ( .A1(n10580), .A2(n10579), .A3(n10578), .A4(n10577), .ZN(
        n10587) );
  AOI22_X1 U13436 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n10581), .B1(
        n10935), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10585) );
  AOI22_X1 U13437 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n11008), .B1(
        n10522), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10584) );
  AOI22_X1 U13438 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n10954), .B1(
        n10523), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10583) );
  AOI22_X1 U13439 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n10524), .B1(
        n10535), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10582) );
  NAND4_X1 U13440 ( .A1(n10585), .A2(n10584), .A3(n10583), .A4(n10582), .ZN(
        n10586) );
  AOI22_X1 U13441 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n10542), .B1(
        n9723), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10592) );
  AOI22_X1 U13442 ( .A1(n10600), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n10517), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10591) );
  AOI22_X1 U13443 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n10949), .B1(
        n10651), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n10590) );
  AOI22_X1 U13444 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n10576), .B1(
        n11008), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n10589) );
  NAND4_X1 U13445 ( .A1(n10592), .A2(n10591), .A3(n10590), .A4(n10589), .ZN(
        n10599) );
  AOI22_X1 U13446 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n10581), .B1(
        n10935), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10597) );
  AOI22_X1 U13447 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n10593), .B1(
        n10522), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n10596) );
  AOI22_X1 U13448 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n10954), .B1(
        n10523), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10595) );
  AOI22_X1 U13449 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n10535), .B1(
        n10524), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10594) );
  NAND4_X1 U13450 ( .A1(n10597), .A2(n10596), .A3(n10595), .A4(n10594), .ZN(
        n10598) );
  NOR2_X1 U13451 ( .A1(n10599), .A2(n10598), .ZN(n13039) );
  OR2_X2 U13452 ( .A1(n13040), .A2(n13039), .ZN(n13108) );
  AOI22_X1 U13453 ( .A1(n9723), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n10542), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10604) );
  AOI22_X1 U13454 ( .A1(n10600), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10517), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10603) );
  AOI22_X1 U13455 ( .A1(n10949), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10651), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10602) );
  AOI22_X1 U13456 ( .A1(n11008), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n10576), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10601) );
  NAND4_X1 U13457 ( .A1(n10604), .A2(n10603), .A3(n10602), .A4(n10601), .ZN(
        n10610) );
  AOI22_X1 U13458 ( .A1(n10935), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n10581), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10608) );
  AOI22_X1 U13459 ( .A1(n10522), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10593), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10607) );
  AOI22_X1 U13460 ( .A1(n10954), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10523), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10606) );
  AOI22_X1 U13461 ( .A1(n10535), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10524), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10605) );
  NAND4_X1 U13462 ( .A1(n10608), .A2(n10607), .A3(n10606), .A4(n10605), .ZN(
        n10609) );
  NOR2_X1 U13463 ( .A1(n10610), .A2(n10609), .ZN(n13109) );
  NOR2_X4 U13464 ( .A1(n13108), .A2(n13109), .ZN(n13289) );
  AOI22_X1 U13465 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n9723), .B1(
        n10542), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10614) );
  INV_X1 U13466 ( .A(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n20884) );
  AOI22_X1 U13467 ( .A1(n10600), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n10517), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10613) );
  AOI22_X1 U13468 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n10651), .B1(
        n10949), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10612) );
  AOI22_X1 U13469 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n10576), .B1(
        n11008), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10611) );
  NAND4_X1 U13470 ( .A1(n10614), .A2(n10613), .A3(n10612), .A4(n10611), .ZN(
        n10620) );
  AOI22_X1 U13471 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n10581), .B1(
        n10935), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10618) );
  AOI22_X1 U13472 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n10593), .B1(
        n10522), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10617) );
  AOI22_X1 U13473 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n10954), .B1(
        n10523), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10616) );
  AOI22_X1 U13474 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n10535), .B1(
        n10524), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10615) );
  NAND4_X1 U13475 ( .A1(n10618), .A2(n10617), .A3(n10616), .A4(n10615), .ZN(
        n10619) );
  OR2_X1 U13476 ( .A1(n10620), .A2(n10619), .ZN(n13288) );
  AOI22_X1 U13477 ( .A1(n9723), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n10542), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10624) );
  AOI22_X1 U13478 ( .A1(n10600), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n10517), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10623) );
  AOI22_X1 U13479 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n10949), .B1(
        n10651), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10622) );
  AOI22_X1 U13480 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n10576), .B1(
        n11008), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10621) );
  NAND4_X1 U13481 ( .A1(n10624), .A2(n10623), .A3(n10622), .A4(n10621), .ZN(
        n10630) );
  AOI22_X1 U13482 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n10935), .B1(
        n10581), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10628) );
  AOI22_X1 U13483 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n10593), .B1(
        n10522), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10627) );
  AOI22_X1 U13484 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n10954), .B1(
        n10523), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10626) );
  AOI22_X1 U13485 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n10535), .B1(
        n10524), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10625) );
  NAND4_X1 U13486 ( .A1(n10628), .A2(n10627), .A3(n10626), .A4(n10625), .ZN(
        n10629) );
  AOI22_X1 U13487 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n9723), .B1(
        n10542), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10634) );
  AOI22_X1 U13488 ( .A1(n10600), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n10517), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10633) );
  AOI22_X1 U13489 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n10651), .B1(
        n10949), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10632) );
  AOI22_X1 U13490 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n11008), .B1(
        n10576), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10631) );
  NAND4_X1 U13491 ( .A1(n10634), .A2(n10633), .A3(n10632), .A4(n10631), .ZN(
        n10640) );
  AOI22_X1 U13492 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n10581), .B1(
        n10935), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10638) );
  AOI22_X1 U13493 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n10593), .B1(
        n10522), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10637) );
  AOI22_X1 U13494 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n10954), .B1(
        n10523), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10636) );
  AOI22_X1 U13495 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n10535), .B1(
        n10524), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10635) );
  NAND4_X1 U13496 ( .A1(n10638), .A2(n10637), .A3(n10636), .A4(n10635), .ZN(
        n10639) );
  AOI22_X1 U13497 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n9723), .B1(
        n10542), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10644) );
  AOI22_X1 U13498 ( .A1(n10600), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n10517), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10643) );
  AOI22_X1 U13499 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n10651), .B1(
        n10949), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10642) );
  AOI22_X1 U13500 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n10576), .B1(
        n11008), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n10641) );
  NAND4_X1 U13501 ( .A1(n10644), .A2(n10643), .A3(n10642), .A4(n10641), .ZN(
        n10650) );
  AOI22_X1 U13502 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n10581), .B1(
        n10935), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10648) );
  AOI22_X1 U13503 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n10593), .B1(
        n10522), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10647) );
  AOI22_X1 U13504 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n10954), .B1(
        n10523), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10646) );
  AOI22_X1 U13505 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n10524), .B1(
        n10535), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10645) );
  NAND4_X1 U13506 ( .A1(n10648), .A2(n10647), .A3(n10646), .A4(n10645), .ZN(
        n10649) );
  NOR2_X1 U13507 ( .A1(n10650), .A2(n10649), .ZN(n14614) );
  AOI22_X1 U13508 ( .A1(n9723), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n10542), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10655) );
  AOI22_X1 U13509 ( .A1(n10600), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n10517), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10654) );
  AOI22_X1 U13510 ( .A1(n10949), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n10651), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10653) );
  AOI22_X1 U13511 ( .A1(n11008), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n10576), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10652) );
  NAND4_X1 U13512 ( .A1(n10655), .A2(n10654), .A3(n10653), .A4(n10652), .ZN(
        n10661) );
  AOI22_X1 U13513 ( .A1(n10935), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n10581), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10659) );
  AOI22_X1 U13514 ( .A1(n10522), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10593), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10658) );
  AOI22_X1 U13515 ( .A1(n10954), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10523), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10657) );
  AOI22_X1 U13516 ( .A1(n10535), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10524), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10656) );
  NAND4_X1 U13517 ( .A1(n10659), .A2(n10658), .A3(n10657), .A4(n10656), .ZN(
        n10660) );
  OR2_X1 U13518 ( .A1(n10661), .A2(n10660), .ZN(n14605) );
  AOI22_X1 U13519 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n9723), .B1(
        n10542), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10665) );
  AOI22_X1 U13520 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n10576), .B1(
        n11008), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10664) );
  AOI22_X1 U13521 ( .A1(n10600), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n10517), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10663) );
  AOI22_X1 U13522 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n10949), .B1(
        n10651), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10662) );
  NAND4_X1 U13523 ( .A1(n10665), .A2(n10664), .A3(n10663), .A4(n10662), .ZN(
        n10671) );
  AOI22_X1 U13524 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n10522), .B1(
        n10593), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10669) );
  AOI22_X1 U13525 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n10581), .B1(
        n10935), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10668) );
  AOI22_X1 U13526 ( .A1(n10954), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_3__6__SCAN_IN), .B2(n10523), .ZN(n10667) );
  AOI22_X1 U13527 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n10535), .B1(
        n10524), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10666) );
  NAND4_X1 U13528 ( .A1(n10669), .A2(n10668), .A3(n10667), .A4(n10666), .ZN(
        n10670) );
  NOR2_X1 U13529 ( .A1(n10671), .A2(n10670), .ZN(n14600) );
  AOI22_X1 U13530 ( .A1(n10844), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10843), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10683) );
  AOI22_X1 U13531 ( .A1(n9748), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(n9753), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10682) );
  AOI22_X1 U13532 ( .A1(n9743), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n10501), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10681) );
  INV_X1 U13533 ( .A(n10833), .ZN(n10839) );
  INV_X1 U13534 ( .A(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10678) );
  NAND2_X1 U13535 ( .A1(n9736), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n10677) );
  INV_X1 U13536 ( .A(n10674), .ZN(n10676) );
  NAND2_X1 U13537 ( .A1(n16164), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10675) );
  NAND2_X1 U13538 ( .A1(n10676), .A2(n10675), .ZN(n10837) );
  OAI211_X1 U13539 ( .C1(n10839), .C2(n10678), .A(n10677), .B(n10837), .ZN(
        n10679) );
  INV_X1 U13540 ( .A(n10679), .ZN(n10680) );
  NAND4_X1 U13541 ( .A1(n10683), .A2(n10682), .A3(n10681), .A4(n10680), .ZN(
        n10692) );
  AOI22_X1 U13542 ( .A1(n9746), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10375), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10690) );
  AOI22_X1 U13543 ( .A1(n10843), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10501), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10689) );
  AOI22_X1 U13544 ( .A1(n10844), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n9743), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10688) );
  INV_X1 U13545 ( .A(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10685) );
  NAND2_X1 U13546 ( .A1(n9736), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n10684) );
  INV_X1 U13547 ( .A(n10837), .ZN(n10808) );
  OAI211_X1 U13548 ( .C1(n10839), .C2(n10685), .A(n10684), .B(n10808), .ZN(
        n10686) );
  INV_X1 U13549 ( .A(n10686), .ZN(n10687) );
  NAND4_X1 U13550 ( .A1(n10690), .A2(n10689), .A3(n10688), .A4(n10687), .ZN(
        n10691) );
  AND2_X1 U13551 ( .A1(n10692), .A2(n10691), .ZN(n10723) );
  NAND2_X1 U13552 ( .A1(n10944), .A2(n10723), .ZN(n10703) );
  AOI22_X1 U13553 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n10600), .B1(
        n10542), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n10696) );
  AOI22_X1 U13554 ( .A1(n9723), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n10517), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10695) );
  AOI22_X1 U13555 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n10949), .B1(
        n10651), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n10694) );
  AOI22_X1 U13556 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n10576), .B1(
        n10593), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10693) );
  NAND4_X1 U13557 ( .A1(n10696), .A2(n10695), .A3(n10694), .A4(n10693), .ZN(
        n10702) );
  AOI22_X1 U13558 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n10581), .B1(
        n10935), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10700) );
  AOI22_X1 U13559 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n10522), .B1(
        n11008), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n10699) );
  AOI22_X1 U13560 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n10535), .B1(
        n10954), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n10698) );
  AOI22_X1 U13561 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n10524), .B1(
        n10523), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10697) );
  NAND4_X1 U13562 ( .A1(n10700), .A2(n10699), .A3(n10698), .A4(n10697), .ZN(
        n10701) );
  OR2_X1 U13563 ( .A1(n10702), .A2(n10701), .ZN(n10705) );
  XNOR2_X1 U13564 ( .A(n10703), .B(n10705), .ZN(n10726) );
  NAND2_X1 U13565 ( .A1(n11164), .A2(n10723), .ZN(n14589) );
  NAND2_X1 U13566 ( .A1(n10705), .A2(n10723), .ZN(n10728) );
  AOI22_X1 U13567 ( .A1(n10844), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n10843), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10712) );
  AOI22_X1 U13568 ( .A1(n9748), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n10501), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10711) );
  AOI22_X1 U13569 ( .A1(n10375), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n13188), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10710) );
  INV_X1 U13570 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10707) );
  NAND2_X1 U13571 ( .A1(n9736), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n10706) );
  OAI211_X1 U13572 ( .C1(n10839), .C2(n10707), .A(n10706), .B(n10837), .ZN(
        n10708) );
  INV_X1 U13573 ( .A(n10708), .ZN(n10709) );
  NAND4_X1 U13574 ( .A1(n10712), .A2(n10711), .A3(n10710), .A4(n10709), .ZN(
        n10720) );
  AOI22_X1 U13575 ( .A1(n10844), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n10843), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10718) );
  AOI22_X1 U13576 ( .A1(n9747), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n10501), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10717) );
  AOI22_X1 U13577 ( .A1(n9752), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n13188), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10716) );
  INV_X1 U13578 ( .A(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11112) );
  NAND2_X1 U13579 ( .A1(n9736), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n10713) );
  OAI211_X1 U13580 ( .C1(n10839), .C2(n11112), .A(n10713), .B(n10808), .ZN(
        n10714) );
  INV_X1 U13581 ( .A(n10714), .ZN(n10715) );
  NAND4_X1 U13582 ( .A1(n10718), .A2(n10717), .A3(n10716), .A4(n10715), .ZN(
        n10719) );
  NAND2_X1 U13583 ( .A1(n10720), .A2(n10719), .ZN(n10727) );
  XOR2_X1 U13584 ( .A(n10728), .B(n10727), .Z(n10721) );
  NAND2_X1 U13585 ( .A1(n10721), .A2(n10744), .ZN(n14574) );
  INV_X1 U13586 ( .A(n10727), .ZN(n10722) );
  NAND2_X1 U13587 ( .A1(n11164), .A2(n10722), .ZN(n14577) );
  INV_X1 U13588 ( .A(n10723), .ZN(n10724) );
  NOR2_X1 U13589 ( .A1(n14577), .A2(n10724), .ZN(n10725) );
  NOR2_X1 U13590 ( .A1(n10728), .A2(n10727), .ZN(n10745) );
  AOI22_X1 U13591 ( .A1(n10844), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n10843), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10734) );
  AOI22_X1 U13592 ( .A1(n9747), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n10375), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10733) );
  INV_X1 U13593 ( .A(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n20774) );
  AOI22_X1 U13594 ( .A1(n9743), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n10501), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10732) );
  NAND2_X1 U13595 ( .A1(n9736), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n10729) );
  OAI211_X1 U13596 ( .C1(n10839), .C2(n10477), .A(n10729), .B(n10837), .ZN(
        n10730) );
  INV_X1 U13597 ( .A(n10730), .ZN(n10731) );
  NAND4_X1 U13598 ( .A1(n10734), .A2(n10733), .A3(n10732), .A4(n10731), .ZN(
        n10743) );
  AOI22_X1 U13599 ( .A1(n10844), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n10843), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10741) );
  AOI22_X1 U13600 ( .A1(n9746), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n9753), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10740) );
  AOI22_X1 U13601 ( .A1(n13188), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n10501), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10739) );
  INV_X1 U13602 ( .A(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10736) );
  INV_X1 U13603 ( .A(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n20881) );
  NAND2_X1 U13604 ( .A1(n9736), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n10735) );
  OAI211_X1 U13605 ( .C1(n10839), .C2(n10736), .A(n10735), .B(n10808), .ZN(
        n10737) );
  INV_X1 U13606 ( .A(n10737), .ZN(n10738) );
  NAND4_X1 U13607 ( .A1(n10741), .A2(n10740), .A3(n10739), .A4(n10738), .ZN(
        n10742) );
  AND2_X1 U13608 ( .A1(n10743), .A2(n10742), .ZN(n10747) );
  NAND2_X1 U13609 ( .A1(n10745), .A2(n10747), .ZN(n10766) );
  OAI211_X1 U13610 ( .C1(n10745), .C2(n10747), .A(n10744), .B(n10766), .ZN(
        n10749) );
  INV_X1 U13611 ( .A(n10749), .ZN(n10746) );
  XNOR2_X1 U13612 ( .A(n10750), .B(n10746), .ZN(n14565) );
  INV_X1 U13613 ( .A(n10747), .ZN(n10748) );
  NOR2_X1 U13614 ( .A1(n10944), .A2(n10748), .ZN(n14564) );
  NAND2_X1 U13615 ( .A1(n14565), .A2(n14564), .ZN(n14563) );
  AOI22_X1 U13616 ( .A1(n10844), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n10843), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10757) );
  AOI22_X1 U13617 ( .A1(n9746), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n10501), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10756) );
  AOI22_X1 U13618 ( .A1(n9752), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(n9743), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10755) );
  NAND2_X1 U13619 ( .A1(n9736), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n10752) );
  OAI211_X1 U13620 ( .C1(n10839), .C2(n11169), .A(n10752), .B(n10837), .ZN(
        n10753) );
  INV_X1 U13621 ( .A(n10753), .ZN(n10754) );
  NAND4_X1 U13622 ( .A1(n10757), .A2(n10756), .A3(n10755), .A4(n10754), .ZN(
        n10765) );
  AOI22_X1 U13623 ( .A1(n10844), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n10843), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10763) );
  AOI22_X1 U13624 ( .A1(n9748), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n10501), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10762) );
  AOI22_X1 U13625 ( .A1(n10375), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n13188), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10761) );
  INV_X1 U13626 ( .A(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11175) );
  NAND2_X1 U13627 ( .A1(n9736), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n10758) );
  OAI211_X1 U13628 ( .C1(n10839), .C2(n11175), .A(n10758), .B(n10808), .ZN(
        n10759) );
  INV_X1 U13629 ( .A(n10759), .ZN(n10760) );
  NAND4_X1 U13630 ( .A1(n10763), .A2(n10762), .A3(n10761), .A4(n10760), .ZN(
        n10764) );
  NAND2_X1 U13631 ( .A1(n10765), .A2(n10764), .ZN(n10768) );
  AOI21_X1 U13632 ( .B1(n10766), .B2(n10768), .A(n10788), .ZN(n10767) );
  OR2_X1 U13633 ( .A1(n10766), .A2(n10768), .ZN(n10789) );
  NAND2_X1 U13634 ( .A1(n10767), .A2(n10789), .ZN(n10770) );
  XNOR2_X1 U13635 ( .A(n10769), .B(n10770), .ZN(n14556) );
  NOR2_X1 U13636 ( .A1(n10944), .A2(n10768), .ZN(n14555) );
  INV_X1 U13637 ( .A(n10769), .ZN(n10771) );
  AOI22_X1 U13638 ( .A1(n10843), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n9753), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10778) );
  AOI22_X1 U13639 ( .A1(n10844), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n9747), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10777) );
  AOI22_X1 U13640 ( .A1(n9743), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n10501), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10776) );
  NAND2_X1 U13641 ( .A1(n9736), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n10772) );
  OAI211_X1 U13642 ( .C1(n10839), .C2(n10773), .A(n10772), .B(n10837), .ZN(
        n10774) );
  INV_X1 U13643 ( .A(n10774), .ZN(n10775) );
  NAND4_X1 U13644 ( .A1(n10778), .A2(n10777), .A3(n10776), .A4(n10775), .ZN(
        n10787) );
  AOI22_X1 U13645 ( .A1(n10843), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n9748), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10785) );
  INV_X1 U13646 ( .A(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n20961) );
  AOI22_X1 U13647 ( .A1(n9753), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n10501), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10784) );
  INV_X1 U13648 ( .A(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n19528) );
  AOI22_X1 U13649 ( .A1(n10844), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n13188), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n10783) );
  INV_X1 U13650 ( .A(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10780) );
  NAND2_X1 U13651 ( .A1(n9736), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n10779) );
  OAI211_X1 U13652 ( .C1(n10839), .C2(n10780), .A(n10779), .B(n10808), .ZN(
        n10781) );
  INV_X1 U13653 ( .A(n10781), .ZN(n10782) );
  NAND4_X1 U13654 ( .A1(n10785), .A2(n10784), .A3(n10783), .A4(n10782), .ZN(
        n10786) );
  NAND2_X1 U13655 ( .A1(n10787), .A2(n10786), .ZN(n10792) );
  NOR2_X1 U13656 ( .A1(n10789), .A2(n10792), .ZN(n14538) );
  AOI211_X1 U13657 ( .C1(n10792), .C2(n10789), .A(n10788), .B(n14538), .ZN(
        n10790) );
  NOR2_X1 U13658 ( .A1(n10944), .A2(n10792), .ZN(n14549) );
  INV_X1 U13659 ( .A(n14539), .ZN(n10807) );
  AOI22_X1 U13660 ( .A1(n10844), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10843), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10798) );
  AOI22_X1 U13661 ( .A1(n9747), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10501), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10797) );
  AOI22_X1 U13662 ( .A1(n9752), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(n9743), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10796) );
  INV_X1 U13663 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12270) );
  NAND2_X1 U13664 ( .A1(n9736), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n10793) );
  OAI211_X1 U13665 ( .C1(n10839), .C2(n12270), .A(n10793), .B(n10837), .ZN(
        n10794) );
  INV_X1 U13666 ( .A(n10794), .ZN(n10795) );
  NAND4_X1 U13667 ( .A1(n10798), .A2(n10797), .A3(n10796), .A4(n10795), .ZN(
        n10806) );
  AOI22_X1 U13668 ( .A1(n10844), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n10843), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10804) );
  AOI22_X1 U13669 ( .A1(n9746), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n10501), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10803) );
  AOI22_X1 U13670 ( .A1(n10375), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n13188), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10802) );
  INV_X1 U13671 ( .A(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11197) );
  NAND2_X1 U13672 ( .A1(n9736), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n10799) );
  OAI211_X1 U13673 ( .C1(n10839), .C2(n11197), .A(n10799), .B(n10808), .ZN(
        n10800) );
  INV_X1 U13674 ( .A(n10800), .ZN(n10801) );
  NAND4_X1 U13675 ( .A1(n10804), .A2(n10803), .A3(n10802), .A4(n10801), .ZN(
        n10805) );
  NAND2_X1 U13676 ( .A1(n10806), .A2(n10805), .ZN(n14540) );
  INV_X1 U13677 ( .A(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11272) );
  INV_X1 U13678 ( .A(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n20775) );
  NAND2_X1 U13679 ( .A1(n13188), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n10809) );
  OAI211_X1 U13680 ( .C1(n10839), .C2(n11272), .A(n10809), .B(n10808), .ZN(
        n10812) );
  INV_X1 U13681 ( .A(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10810) );
  INV_X1 U13682 ( .A(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11267) );
  OAI22_X1 U13683 ( .A1(n10810), .A2(n9730), .B1(n10673), .B2(n11267), .ZN(
        n10811) );
  NOR2_X1 U13684 ( .A1(n10812), .A2(n10811), .ZN(n10815) );
  AOI22_X1 U13685 ( .A1(n10843), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n9746), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10814) );
  AOI22_X1 U13686 ( .A1(n10844), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n9753), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10813) );
  NAND3_X1 U13687 ( .A1(n10815), .A2(n10814), .A3(n10813), .ZN(n10824) );
  AOI22_X1 U13688 ( .A1(n10844), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n10843), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10822) );
  AOI22_X1 U13689 ( .A1(n9748), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n10501), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10821) );
  AOI22_X1 U13690 ( .A1(n9753), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n13188), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10820) );
  INV_X1 U13691 ( .A(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10817) );
  INV_X1 U13692 ( .A(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n19094) );
  OR2_X1 U13693 ( .A1(n10839), .A2(n19094), .ZN(n10816) );
  OAI211_X1 U13694 ( .C1(n10817), .C2(n9730), .A(n10816), .B(n10837), .ZN(
        n10818) );
  INV_X1 U13695 ( .A(n10818), .ZN(n10819) );
  NAND4_X1 U13696 ( .A1(n10822), .A2(n10821), .A3(n10820), .A4(n10819), .ZN(
        n10823) );
  NAND2_X1 U13697 ( .A1(n10824), .A2(n10823), .ZN(n10828) );
  INV_X1 U13698 ( .A(n14540), .ZN(n10825) );
  AND2_X1 U13699 ( .A1(n10944), .A2(n10825), .ZN(n10826) );
  NAND2_X1 U13700 ( .A1(n14538), .A2(n10826), .ZN(n10827) );
  NOR2_X1 U13701 ( .A1(n10827), .A2(n10828), .ZN(n10829) );
  AOI21_X1 U13702 ( .B1(n10828), .B2(n10827), .A(n10829), .ZN(n14533) );
  INV_X1 U13703 ( .A(n10829), .ZN(n10830) );
  AOI22_X1 U13704 ( .A1(n10844), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n10843), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n10832) );
  AOI22_X1 U13705 ( .A1(n9747), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n9752), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n10831) );
  NAND2_X1 U13706 ( .A1(n10832), .A2(n10831), .ZN(n10850) );
  INV_X1 U13707 ( .A(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n10836) );
  AOI22_X1 U13708 ( .A1(n13188), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n10501), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10835) );
  AOI21_X1 U13709 ( .B1(n10833), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A(
        n10837), .ZN(n10834) );
  OAI211_X1 U13710 ( .C1(n9730), .C2(n10836), .A(n10835), .B(n10834), .ZN(
        n10849) );
  OAI21_X1 U13711 ( .B1(n10839), .B2(n10838), .A(n10837), .ZN(n10842) );
  INV_X1 U13712 ( .A(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10840) );
  INV_X1 U13713 ( .A(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n19300) );
  OAI22_X1 U13714 ( .A1(n10286), .A2(n10840), .B1(n10673), .B2(n19300), .ZN(
        n10841) );
  AOI211_X1 U13715 ( .C1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .C2(n9736), .A(
        n10842), .B(n10841), .ZN(n10847) );
  AOI22_X1 U13716 ( .A1(n10844), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n10843), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10846) );
  AOI22_X1 U13717 ( .A1(n9748), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n10375), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10845) );
  NAND3_X1 U13718 ( .A1(n10847), .A2(n10846), .A3(n10845), .ZN(n10848) );
  OAI21_X1 U13719 ( .B1(n10850), .B2(n10849), .A(n10848), .ZN(n10851) );
  AOI22_X1 U13720 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n10542), .B1(
        n9723), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10855) );
  AOI22_X1 U13721 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n10600), .B1(
        n10949), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n10854) );
  AOI22_X1 U13722 ( .A1(n10651), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n10517), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10853) );
  AOI22_X1 U13723 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n10522), .B1(
        n10593), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10852) );
  NAND4_X1 U13724 ( .A1(n10855), .A2(n10854), .A3(n10853), .A4(n10852), .ZN(
        n10861) );
  AOI22_X1 U13725 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n10581), .B1(
        n10935), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10859) );
  AOI22_X1 U13726 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n10576), .B1(
        n11008), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10858) );
  AOI22_X1 U13727 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n10954), .B1(
        n10523), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10857) );
  AOI22_X1 U13728 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n10535), .B1(
        n10524), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10856) );
  NAND4_X1 U13729 ( .A1(n10859), .A2(n10858), .A3(n10857), .A4(n10856), .ZN(
        n10860) );
  MUX2_X1 U13730 ( .A(n10862), .B(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .S(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Z(n10879) );
  NAND2_X1 U13731 ( .A1(n10879), .A2(n10880), .ZN(n10864) );
  NAND2_X1 U13732 ( .A1(n10862), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10863) );
  NAND2_X1 U13733 ( .A1(n10864), .A2(n10863), .ZN(n10875) );
  XNOR2_X1 U13734 ( .A(n16164), .B(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n10873) );
  NAND2_X1 U13735 ( .A1(n10875), .A2(n10873), .ZN(n10866) );
  NAND2_X1 U13736 ( .A1(n19704), .A2(n16164), .ZN(n10865) );
  NAND2_X1 U13737 ( .A1(n10866), .A2(n10865), .ZN(n10872) );
  XNOR2_X1 U13738 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n10870) );
  NOR2_X1 U13739 ( .A1(n10359), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n10867) );
  NOR2_X1 U13740 ( .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n15508), .ZN(
        n10868) );
  NAND2_X1 U13741 ( .A1(n10889), .A2(n10868), .ZN(n10888) );
  MUX2_X1 U13742 ( .A(n11487), .B(n10888), .S(n11476), .Z(n11456) );
  INV_X1 U13743 ( .A(n10870), .ZN(n10871) );
  XNOR2_X1 U13744 ( .A(n10872), .B(n10871), .ZN(n11239) );
  AOI21_X1 U13745 ( .B1(n11456), .B2(n11239), .A(n10407), .ZN(n10895) );
  INV_X1 U13746 ( .A(n10873), .ZN(n10874) );
  XNOR2_X1 U13747 ( .A(n10875), .B(n10874), .ZN(n11443) );
  NAND2_X1 U13748 ( .A1(n19740), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n19739) );
  AOI21_X1 U13749 ( .B1(n19739), .B2(n10944), .A(n11443), .ZN(n10887) );
  INV_X1 U13750 ( .A(n11443), .ZN(n10882) );
  INV_X1 U13751 ( .A(n10880), .ZN(n10878) );
  NAND2_X1 U13752 ( .A1(n10876), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n10877) );
  AND2_X1 U13753 ( .A1(n10878), .A2(n10877), .ZN(n11442) );
  INV_X1 U13754 ( .A(n10879), .ZN(n11454) );
  XNOR2_X1 U13755 ( .A(n11454), .B(n10880), .ZN(n10920) );
  OAI21_X1 U13756 ( .B1(n10944), .B2(n11442), .A(n10920), .ZN(n10881) );
  OAI21_X1 U13757 ( .B1(n10882), .B2(n10944), .A(n10881), .ZN(n10883) );
  NAND2_X1 U13758 ( .A1(n10883), .A2(n16176), .ZN(n10885) );
  INV_X1 U13759 ( .A(n11442), .ZN(n11252) );
  OAI21_X1 U13760 ( .B1(n11454), .B2(n11252), .A(n10407), .ZN(n10884) );
  NAND2_X1 U13761 ( .A1(n10885), .A2(n10884), .ZN(n10886) );
  OAI21_X1 U13762 ( .B1(n11237), .B2(n10887), .A(n10886), .ZN(n10894) );
  NAND2_X1 U13763 ( .A1(n10888), .A2(n11239), .ZN(n11445) );
  INV_X1 U13764 ( .A(n10889), .ZN(n10892) );
  INV_X1 U13765 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n16179) );
  NAND2_X1 U13766 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n16179), .ZN(
        n10891) );
  INV_X1 U13767 ( .A(n11459), .ZN(n10897) );
  AOI21_X1 U13768 ( .B1(n10407), .B2(n11445), .A(n10897), .ZN(n10893) );
  OAI21_X1 U13769 ( .B1(n10895), .B2(n10894), .A(n10893), .ZN(n10896) );
  MUX2_X1 U13770 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B(n10896), .S(
        P2_STATE2_REG_0__SCAN_IN), .Z(n11440) );
  INV_X1 U13771 ( .A(n19739), .ZN(n10898) );
  NAND2_X1 U13772 ( .A1(n10898), .A2(n10897), .ZN(n10899) );
  NAND2_X1 U13773 ( .A1(n11164), .A2(n10909), .ZN(n10915) );
  INV_X1 U13774 ( .A(n10401), .ZN(n10900) );
  AOI21_X1 U13775 ( .B1(n10915), .B2(n16176), .A(n10900), .ZN(n10905) );
  NAND2_X1 U13776 ( .A1(n10902), .A2(n10390), .ZN(n10901) );
  AND2_X1 U13777 ( .A1(n11164), .A2(n19740), .ZN(n11461) );
  NAND2_X1 U13778 ( .A1(n10901), .A2(n11461), .ZN(n11533) );
  INV_X1 U13779 ( .A(n10902), .ZN(n10903) );
  NAND2_X1 U13780 ( .A1(n10903), .A2(n10398), .ZN(n10904) );
  OAI211_X1 U13781 ( .C1(n10905), .C2(n10391), .A(n11533), .B(n10904), .ZN(
        n10906) );
  INV_X1 U13782 ( .A(n10906), .ZN(n10914) );
  NAND2_X1 U13783 ( .A1(n10908), .A2(n10909), .ZN(n10911) );
  NAND2_X1 U13784 ( .A1(n10911), .A2(n10910), .ZN(n10912) );
  NAND2_X1 U13785 ( .A1(n10907), .A2(n10912), .ZN(n10913) );
  NAND2_X1 U13786 ( .A1(n10914), .A2(n10913), .ZN(n11467) );
  NAND2_X1 U13787 ( .A1(n12976), .A2(n16169), .ZN(n11941) );
  NAND2_X1 U13788 ( .A1(n10917), .A2(n10916), .ZN(n11528) );
  NAND2_X1 U13789 ( .A1(n11941), .A2(n11528), .ZN(n10918) );
  NAND2_X1 U13790 ( .A1(n13196), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12957) );
  NAND2_X1 U13791 ( .A1(n10918), .A2(n18949), .ZN(n10924) );
  INV_X1 U13792 ( .A(n10919), .ZN(n16168) );
  NAND2_X1 U13793 ( .A1(n11443), .A2(n10920), .ZN(n10921) );
  OR2_X1 U13794 ( .A1(n11445), .A2(n10921), .ZN(n10922) );
  NAND2_X1 U13795 ( .A1(n10922), .A2(n11459), .ZN(n16167) );
  AND2_X1 U13796 ( .A1(n16168), .A2(n11861), .ZN(n11939) );
  NAND2_X1 U13797 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n19736) );
  AND2_X1 U13798 ( .A1(n11526), .A2(n19736), .ZN(n11938) );
  NAND2_X1 U13799 ( .A1(n19735), .A2(n11938), .ZN(n10923) );
  NAND2_X1 U13800 ( .A1(n11709), .A2(n15928), .ZN(n11108) );
  NAND2_X1 U13801 ( .A1(n11516), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n10929) );
  AND2_X1 U13802 ( .A1(n10927), .A2(n19714), .ZN(n10981) );
  AOI22_X1 U13803 ( .A1(n10926), .A2(P2_EAX_REG_21__SCAN_IN), .B1(n11515), 
        .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n10928) );
  AND2_X1 U13804 ( .A1(n10929), .A2(n10928), .ZN(n14688) );
  AOI22_X1 U13805 ( .A1(n9723), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n10542), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10934) );
  AOI22_X1 U13806 ( .A1(n10600), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n10517), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10933) );
  AOI22_X1 U13807 ( .A1(n10949), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n10651), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10932) );
  AOI22_X1 U13808 ( .A1(n11008), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n10576), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10931) );
  NAND4_X1 U13809 ( .A1(n10934), .A2(n10933), .A3(n10932), .A4(n10931), .ZN(
        n10941) );
  AOI22_X1 U13810 ( .A1(n10935), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10581), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10939) );
  AOI22_X1 U13811 ( .A1(n10522), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n10593), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10938) );
  AOI22_X1 U13812 ( .A1(n10954), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n10523), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10937) );
  AOI22_X1 U13813 ( .A1(n10535), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n10524), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10936) );
  NAND4_X1 U13814 ( .A1(n10939), .A2(n10938), .A3(n10937), .A4(n10936), .ZN(
        n10940) );
  NAND2_X1 U13815 ( .A1(n11071), .A2(n11923), .ZN(n10943) );
  NAND2_X1 U13816 ( .A1(n11965), .A2(n10981), .ZN(n10979) );
  NAND2_X1 U13817 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n10942) );
  NAND4_X1 U13818 ( .A1(n10943), .A2(n11000), .A3(n10979), .A4(n10942), .ZN(
        n11974) );
  AOI21_X1 U13819 ( .B1(n10383), .B2(P2_EAX_REG_0__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n10946) );
  NAND2_X1 U13820 ( .A1(n10944), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n10945) );
  OAI211_X1 U13821 ( .C1(n11089), .C2(n10947), .A(n10946), .B(n10945), .ZN(
        n11973) );
  NAND2_X1 U13822 ( .A1(n11974), .A2(n11973), .ZN(n10966) );
  AOI22_X1 U13823 ( .A1(n10926), .A2(P2_EAX_REG_1__SCAN_IN), .B1(n10981), .B2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n10948) );
  XNOR2_X1 U13824 ( .A(n10966), .B(n10967), .ZN(n12205) );
  AOI22_X1 U13825 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n10542), .B1(
        n9723), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10953) );
  AOI22_X1 U13826 ( .A1(n10600), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n10935), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10952) );
  AOI22_X1 U13827 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n10576), .B1(
        n11008), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10951) );
  AOI22_X1 U13828 ( .A1(n10949), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n10517), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10950) );
  NAND4_X1 U13829 ( .A1(n10953), .A2(n10952), .A3(n10951), .A4(n10950), .ZN(
        n10960) );
  AOI22_X1 U13830 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n10523), .B1(
        n10954), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10958) );
  AOI22_X1 U13831 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n10535), .B1(
        n10524), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10957) );
  AOI22_X1 U13832 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n10522), .B1(
        n10593), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10956) );
  AOI22_X1 U13833 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n10651), .B1(
        n10581), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10955) );
  NAND4_X1 U13834 ( .A1(n10958), .A2(n10957), .A3(n10956), .A4(n10955), .ZN(
        n10959) );
  INV_X1 U13835 ( .A(n11071), .ZN(n10961) );
  OR2_X1 U13836 ( .A1(n11478), .A2(n10961), .ZN(n10965) );
  AND2_X1 U13837 ( .A1(n10390), .A2(n19714), .ZN(n10963) );
  NOR2_X1 U13838 ( .A1(n19714), .A2(n10862), .ZN(n10962) );
  AOI21_X1 U13839 ( .B1(n10908), .B2(n10963), .A(n10962), .ZN(n10964) );
  NAND2_X1 U13840 ( .A1(n10965), .A2(n10964), .ZN(n12204) );
  NAND2_X1 U13841 ( .A1(n10967), .A2(n10966), .ZN(n10968) );
  OAI21_X1 U13842 ( .B1(n12205), .B2(n12204), .A(n10968), .ZN(n10985) );
  AOI22_X1 U13843 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n9723), .B1(
        n10600), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10972) );
  AOI22_X1 U13844 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n10542), .B1(
        n10651), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10971) );
  AOI22_X1 U13845 ( .A1(n10949), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n10517), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10970) );
  AOI22_X1 U13846 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n10576), .B1(
        n10522), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10969) );
  NAND4_X1 U13847 ( .A1(n10972), .A2(n10971), .A3(n10970), .A4(n10969), .ZN(
        n10978) );
  AOI22_X1 U13848 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n10581), .B1(
        n10935), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10976) );
  AOI22_X1 U13849 ( .A1(n11008), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n10593), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10975) );
  AOI22_X1 U13850 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n10535), .B1(
        n10954), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10974) );
  AOI22_X1 U13851 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n10524), .B1(
        n10523), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10973) );
  NAND4_X1 U13852 ( .A1(n10976), .A2(n10975), .A3(n10974), .A4(n10973), .ZN(
        n10977) );
  NAND2_X1 U13853 ( .A1(n11071), .A2(n11165), .ZN(n10980) );
  OAI211_X1 U13854 ( .C1(n19714), .C2(n19704), .A(n10980), .B(n10979), .ZN(
        n10984) );
  XNOR2_X1 U13855 ( .A(n10985), .B(n10984), .ZN(n12252) );
  NAND2_X1 U13856 ( .A1(n11516), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n10983) );
  AOI22_X1 U13857 ( .A1(n11085), .A2(P2_EAX_REG_2__SCAN_IN), .B1(n11515), .B2(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n10982) );
  NAND2_X1 U13858 ( .A1(n12252), .A2(n12251), .ZN(n12253) );
  INV_X1 U13859 ( .A(n10984), .ZN(n10986) );
  NAND2_X1 U13860 ( .A1(n10986), .A2(n10985), .ZN(n10987) );
  AOI22_X1 U13861 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n9723), .B1(
        n10600), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10991) );
  AOI22_X1 U13862 ( .A1(n10542), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n10517), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10990) );
  AOI22_X1 U13863 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n10651), .B1(
        n10949), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10989) );
  AOI22_X1 U13864 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n10522), .B1(
        n11008), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10988) );
  NAND4_X1 U13865 ( .A1(n10991), .A2(n10990), .A3(n10989), .A4(n10988), .ZN(
        n10997) );
  AOI22_X1 U13866 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n10581), .B1(
        n10935), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10995) );
  AOI22_X1 U13867 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n10593), .B1(
        n10576), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10994) );
  AOI22_X1 U13868 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n10523), .B1(
        n10954), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10993) );
  AOI22_X1 U13869 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n10535), .B1(
        n10524), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10992) );
  NAND4_X1 U13870 ( .A1(n10995), .A2(n10994), .A3(n10993), .A4(n10992), .ZN(
        n10996) );
  INV_X1 U13871 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19697) );
  NAND2_X1 U13872 ( .A1(n11515), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10998) );
  OAI21_X1 U13873 ( .B1(n19714), .B2(n19697), .A(n10998), .ZN(n10999) );
  AOI21_X1 U13874 ( .B1(n11071), .B2(n11240), .A(n10999), .ZN(n11005) );
  NAND2_X1 U13875 ( .A1(n11085), .A2(P2_EAX_REG_3__SCAN_IN), .ZN(n11001) );
  OAI21_X1 U13876 ( .B1(n11089), .B2(n11002), .A(n11001), .ZN(n11003) );
  INV_X1 U13877 ( .A(n11003), .ZN(n11004) );
  INV_X1 U13878 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n11551) );
  AOI22_X1 U13879 ( .A1(n11085), .A2(P2_EAX_REG_4__SCAN_IN), .B1(n11515), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n11007) );
  NAND2_X1 U13880 ( .A1(n11071), .A2(n11487), .ZN(n11006) );
  OAI211_X1 U13881 ( .C1(n11089), .C2(n11551), .A(n11007), .B(n11006), .ZN(
        n12487) );
  INV_X1 U13882 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n11557) );
  AOI22_X1 U13883 ( .A1(n9723), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n10542), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11012) );
  AOI22_X1 U13884 ( .A1(n10600), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n10517), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11011) );
  AOI22_X1 U13885 ( .A1(n10949), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n10651), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11010) );
  AOI22_X1 U13886 ( .A1(n11008), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10576), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11009) );
  NAND4_X1 U13887 ( .A1(n11012), .A2(n11011), .A3(n11010), .A4(n11009), .ZN(
        n11018) );
  AOI22_X1 U13888 ( .A1(n10935), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n10581), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11016) );
  AOI22_X1 U13889 ( .A1(n10522), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n10593), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11015) );
  AOI22_X1 U13890 ( .A1(n10954), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10523), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11014) );
  AOI22_X1 U13891 ( .A1(n10535), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n10524), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11013) );
  NAND4_X1 U13892 ( .A1(n11016), .A2(n11015), .A3(n11014), .A4(n11013), .ZN(
        n11017) );
  INV_X1 U13893 ( .A(n11242), .ZN(n11019) );
  NAND2_X1 U13894 ( .A1(n11071), .A2(n11019), .ZN(n11021) );
  AOI22_X1 U13895 ( .A1(n11085), .A2(P2_EAX_REG_5__SCAN_IN), .B1(n11515), .B2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n11020) );
  OAI211_X1 U13896 ( .C1(n11089), .C2(n11557), .A(n11021), .B(n11020), .ZN(
        n12482) );
  AOI22_X1 U13897 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n10542), .B1(
        n9723), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11025) );
  AOI22_X1 U13898 ( .A1(n10600), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10517), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11024) );
  AOI22_X1 U13899 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n10651), .B1(
        n10949), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11023) );
  AOI22_X1 U13900 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n10576), .B1(
        n11008), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11022) );
  NAND4_X1 U13901 ( .A1(n11025), .A2(n11024), .A3(n11023), .A4(n11022), .ZN(
        n11031) );
  AOI22_X1 U13902 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n10581), .B1(
        n10935), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11029) );
  AOI22_X1 U13903 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n10522), .B1(
        n10593), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11028) );
  AOI22_X1 U13904 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n10523), .B1(
        n10954), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11027) );
  AOI22_X1 U13905 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n10535), .B1(
        n10524), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11026) );
  NAND4_X1 U13906 ( .A1(n11029), .A2(n11028), .A3(n11027), .A4(n11026), .ZN(
        n11030) );
  NAND2_X1 U13907 ( .A1(n11071), .A2(n11299), .ZN(n11032) );
  INV_X1 U13908 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n11564) );
  AOI22_X1 U13909 ( .A1(n11085), .A2(P2_EAX_REG_6__SCAN_IN), .B1(n11515), .B2(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n11033) );
  OAI21_X1 U13910 ( .B1(n11089), .B2(n11564), .A(n11033), .ZN(n11967) );
  NAND2_X1 U13911 ( .A1(n11968), .A2(n11967), .ZN(n11970) );
  NAND2_X1 U13912 ( .A1(n10542), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n11037) );
  NAND2_X1 U13913 ( .A1(n9723), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n11036) );
  NAND2_X1 U13914 ( .A1(n10600), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n11035) );
  NAND2_X1 U13915 ( .A1(n10517), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n11034) );
  AOI22_X1 U13916 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n10535), .B1(
        n10524), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11042) );
  AOI22_X1 U13917 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n10523), .B1(
        n10954), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11041) );
  NAND2_X1 U13918 ( .A1(n10935), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n11040) );
  NAND2_X1 U13919 ( .A1(n10581), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n11039) );
  AOI22_X1 U13920 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n10522), .B1(
        n10593), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11048) );
  NAND2_X1 U13921 ( .A1(n10949), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n11046) );
  NAND2_X1 U13922 ( .A1(n10651), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n11045) );
  NAND2_X1 U13923 ( .A1(n11008), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n11044) );
  NAND2_X1 U13924 ( .A1(n10576), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n11043) );
  NAND2_X1 U13925 ( .A1(n11071), .A2(n11307), .ZN(n11051) );
  NAND2_X1 U13926 ( .A1(n11516), .A2(P2_REIP_REG_7__SCAN_IN), .ZN(n11053) );
  AOI22_X1 U13927 ( .A1(n11085), .A2(P2_EAX_REG_7__SCAN_IN), .B1(n11515), .B2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n11052) );
  INV_X1 U13928 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n11576) );
  AOI22_X1 U13929 ( .A1(n11085), .A2(P2_EAX_REG_8__SCAN_IN), .B1(n11515), .B2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n11055) );
  NAND2_X1 U13930 ( .A1(n11071), .A2(n12284), .ZN(n11054) );
  OAI211_X1 U13931 ( .C1(n11089), .C2(n11576), .A(n11055), .B(n11054), .ZN(
        n11980) );
  INV_X1 U13932 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n11579) );
  AOI22_X1 U13933 ( .A1(n11085), .A2(P2_EAX_REG_9__SCAN_IN), .B1(n11515), .B2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n11058) );
  NAND2_X1 U13934 ( .A1(n11071), .A2(n11056), .ZN(n11057) );
  OAI211_X1 U13935 ( .C1(n11089), .C2(n11579), .A(n11058), .B(n11057), .ZN(
        n15032) );
  INV_X1 U13936 ( .A(n15032), .ZN(n11059) );
  INV_X1 U13937 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n11585) );
  AOI22_X1 U13938 ( .A1(n11085), .A2(P2_EAX_REG_10__SCAN_IN), .B1(n11515), 
        .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n11061) );
  NAND2_X1 U13939 ( .A1(n11071), .A2(n12301), .ZN(n11060) );
  OAI211_X1 U13940 ( .C1(n11089), .C2(n11585), .A(n11061), .B(n11060), .ZN(
        n12227) );
  AOI22_X1 U13941 ( .A1(n11516), .A2(P2_REIP_REG_11__SCAN_IN), .B1(n11071), 
        .B2(n12518), .ZN(n11063) );
  AOI22_X1 U13942 ( .A1(n11085), .A2(P2_EAX_REG_11__SCAN_IN), .B1(n11515), 
        .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n11062) );
  INV_X1 U13943 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n11594) );
  AOI22_X1 U13944 ( .A1(n11085), .A2(P2_EAX_REG_12__SCAN_IN), .B1(n11515), 
        .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n11065) );
  NAND2_X1 U13945 ( .A1(n11071), .A2(n12517), .ZN(n11064) );
  OAI211_X1 U13946 ( .C1(n11089), .C2(n11594), .A(n11065), .B(n11064), .ZN(
        n12261) );
  AOI22_X1 U13947 ( .A1(n11516), .A2(P2_REIP_REG_13__SCAN_IN), .B1(n11071), 
        .B2(n12898), .ZN(n11067) );
  AOI22_X1 U13948 ( .A1(n11085), .A2(P2_EAX_REG_13__SCAN_IN), .B1(n11515), 
        .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n11066) );
  INV_X1 U13949 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n11608) );
  AOI22_X1 U13950 ( .A1(n11085), .A2(P2_EAX_REG_14__SCAN_IN), .B1(n11515), 
        .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n11069) );
  NAND2_X1 U13951 ( .A1(n11071), .A2(n12891), .ZN(n11068) );
  OAI211_X1 U13952 ( .C1(n11089), .C2(n11608), .A(n11069), .B(n11068), .ZN(
        n15014) );
  INV_X1 U13953 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n11611) );
  AOI22_X1 U13954 ( .A1(n11085), .A2(P2_EAX_REG_15__SCAN_IN), .B1(n11515), 
        .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n11073) );
  INV_X1 U13955 ( .A(n13039), .ZN(n11070) );
  NAND2_X1 U13956 ( .A1(n11071), .A2(n11070), .ZN(n11072) );
  OAI211_X1 U13957 ( .C1(n11089), .C2(n11611), .A(n11073), .B(n11072), .ZN(
        n12884) );
  INV_X1 U13958 ( .A(n12884), .ZN(n11074) );
  INV_X1 U13959 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n19647) );
  AOI22_X1 U13960 ( .A1(n11085), .A2(P2_EAX_REG_16__SCAN_IN), .B1(n11515), 
        .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n11075) );
  OAI21_X1 U13961 ( .B1(n11089), .B2(n19647), .A(n11075), .ZN(n13111) );
  AOI222_X1 U13962 ( .A1(n11516), .A2(P2_REIP_REG_17__SCAN_IN), .B1(n11085), 
        .B2(P2_EAX_REG_17__SCAN_IN), .C1(n11515), .C2(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n13291) );
  INV_X1 U13963 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n19650) );
  AOI22_X1 U13964 ( .A1(n11085), .A2(P2_EAX_REG_18__SCAN_IN), .B1(n11515), 
        .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n11076) );
  OAI21_X1 U13965 ( .B1(n11089), .B2(n19650), .A(n11076), .ZN(n13333) );
  INV_X1 U13966 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n11628) );
  AOI22_X1 U13967 ( .A1(n11085), .A2(P2_EAX_REG_19__SCAN_IN), .B1(n11515), 
        .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n11077) );
  OAI21_X1 U13968 ( .B1(n11089), .B2(n11628), .A(n11077), .ZN(n14704) );
  INV_X1 U13969 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n20777) );
  AOI22_X1 U13970 ( .A1(n10926), .A2(P2_EAX_REG_20__SCAN_IN), .B1(n11515), 
        .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n11078) );
  OAI21_X1 U13971 ( .B1(n11089), .B2(n20777), .A(n11078), .ZN(n11079) );
  INV_X1 U13972 ( .A(n11079), .ZN(n14696) );
  INV_X1 U13973 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n19656) );
  AOI22_X1 U13974 ( .A1(n10926), .A2(P2_EAX_REG_22__SCAN_IN), .B1(n11515), 
        .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n11080) );
  OAI21_X1 U13975 ( .B1(n11089), .B2(n19656), .A(n11080), .ZN(n14681) );
  NAND2_X1 U13976 ( .A1(n11516), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n11082) );
  AOI22_X1 U13977 ( .A1(n10926), .A2(P2_EAX_REG_23__SCAN_IN), .B1(n11515), 
        .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n11081) );
  NAND2_X1 U13978 ( .A1(n11082), .A2(n11081), .ZN(n15916) );
  NAND2_X1 U13979 ( .A1(n11516), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n11084) );
  AOI22_X1 U13980 ( .A1(n10926), .A2(P2_EAX_REG_24__SCAN_IN), .B1(n11515), 
        .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n11083) );
  AND2_X1 U13981 ( .A1(n11084), .A2(n11083), .ZN(n14670) );
  NAND2_X1 U13982 ( .A1(n11516), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n11087) );
  AOI22_X1 U13983 ( .A1(n11085), .A2(P2_EAX_REG_25__SCAN_IN), .B1(n11515), 
        .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n11086) );
  AND2_X1 U13984 ( .A1(n11087), .A2(n11086), .ZN(n14664) );
  INV_X1 U13985 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n20880) );
  AOI22_X1 U13986 ( .A1(n10926), .A2(P2_EAX_REG_26__SCAN_IN), .B1(n11515), 
        .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n11088) );
  OAI21_X1 U13987 ( .B1(n11089), .B2(n20880), .A(n11088), .ZN(n14656) );
  NAND2_X1 U13988 ( .A1(n11516), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n11091) );
  AOI22_X1 U13989 ( .A1(n10926), .A2(P2_EAX_REG_27__SCAN_IN), .B1(n11515), 
        .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n11090) );
  AND2_X1 U13990 ( .A1(n11091), .A2(n11090), .ZN(n14650) );
  NAND2_X1 U13991 ( .A1(n11516), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n11093) );
  AOI22_X1 U13992 ( .A1(n10926), .A2(P2_EAX_REG_28__SCAN_IN), .B1(n11515), 
        .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n11092) );
  AND2_X1 U13993 ( .A1(n11093), .A2(n11092), .ZN(n14641) );
  NAND2_X1 U13994 ( .A1(n11516), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n11095) );
  AOI22_X1 U13995 ( .A1(n10926), .A2(P2_EAX_REG_29__SCAN_IN), .B1(n11515), 
        .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n11094) );
  AND2_X1 U13996 ( .A1(n11095), .A2(n11094), .ZN(n14633) );
  AOI222_X1 U13997 ( .A1(n11516), .A2(P2_REIP_REG_30__SCAN_IN), .B1(n11085), 
        .B2(P2_EAX_REG_30__SCAN_IN), .C1(n11515), .C2(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n11514) );
  XNOR2_X1 U13998 ( .A(n14632), .B(n11514), .ZN(n15843) );
  AOI22_X1 U13999 ( .A1(n15843), .A2(n18930), .B1(n18934), .B2(
        P2_EAX_REG_30__SCAN_IN), .ZN(n11107) );
  NAND2_X1 U14000 ( .A1(n18948), .A2(n10390), .ZN(n11966) );
  NOR2_X2 U14001 ( .A1(n11966), .A2(n11354), .ZN(n15927) );
  NOR4_X1 U14002 ( .A1(P2_ADDRESS_REG_16__SCAN_IN), .A2(
        P2_ADDRESS_REG_15__SCAN_IN), .A3(P2_ADDRESS_REG_14__SCAN_IN), .A4(
        P2_ADDRESS_REG_13__SCAN_IN), .ZN(n11099) );
  NOR4_X1 U14003 ( .A1(P2_ADDRESS_REG_20__SCAN_IN), .A2(
        P2_ADDRESS_REG_19__SCAN_IN), .A3(P2_ADDRESS_REG_18__SCAN_IN), .A4(
        P2_ADDRESS_REG_17__SCAN_IN), .ZN(n11098) );
  NOR4_X1 U14004 ( .A1(P2_ADDRESS_REG_7__SCAN_IN), .A2(
        P2_ADDRESS_REG_5__SCAN_IN), .A3(P2_ADDRESS_REG_4__SCAN_IN), .A4(
        P2_ADDRESS_REG_3__SCAN_IN), .ZN(n11097) );
  NOR4_X1 U14005 ( .A1(P2_ADDRESS_REG_12__SCAN_IN), .A2(
        P2_ADDRESS_REG_11__SCAN_IN), .A3(P2_ADDRESS_REG_9__SCAN_IN), .A4(
        P2_ADDRESS_REG_8__SCAN_IN), .ZN(n11096) );
  NAND4_X1 U14006 ( .A1(n11099), .A2(n11098), .A3(n11097), .A4(n11096), .ZN(
        n11104) );
  NOR4_X1 U14007 ( .A1(P2_ADDRESS_REG_1__SCAN_IN), .A2(
        P2_ADDRESS_REG_0__SCAN_IN), .A3(P2_ADDRESS_REG_6__SCAN_IN), .A4(
        P2_ADDRESS_REG_10__SCAN_IN), .ZN(n11102) );
  NOR4_X1 U14008 ( .A1(P2_ADDRESS_REG_24__SCAN_IN), .A2(
        P2_ADDRESS_REG_23__SCAN_IN), .A3(P2_ADDRESS_REG_22__SCAN_IN), .A4(
        P2_ADDRESS_REG_21__SCAN_IN), .ZN(n11101) );
  NOR4_X1 U14009 ( .A1(P2_ADDRESS_REG_28__SCAN_IN), .A2(
        P2_ADDRESS_REG_27__SCAN_IN), .A3(P2_ADDRESS_REG_26__SCAN_IN), .A4(
        P2_ADDRESS_REG_25__SCAN_IN), .ZN(n11100) );
  INV_X1 U14010 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n19636) );
  NAND4_X1 U14011 ( .A1(n11102), .A2(n11101), .A3(n11100), .A4(n19636), .ZN(
        n11103) );
  MUX2_X1 U14012 ( .A(BUF1_REG_14__SCAN_IN), .B(BUF2_REG_14__SCAN_IN), .S(
        n14634), .Z(n19023) );
  NAND2_X1 U14013 ( .A1(n15927), .A2(n19023), .ZN(n11106) );
  NOR3_X4 U14014 ( .A1(n11966), .A2(n19085), .A3(n12980), .ZN(n18929) );
  NOR3_X4 U14015 ( .A1(n11966), .A2(n19085), .A3(n14634), .ZN(n18931) );
  AOI22_X1 U14016 ( .A1(n18929), .A2(BUF2_REG_30__SCAN_IN), .B1(n18931), .B2(
        BUF1_REG_30__SCAN_IN), .ZN(n11105) );
  NAND2_X1 U14017 ( .A1(n11108), .A2(n10270), .ZN(P2_U2889) );
  INV_X1 U14018 ( .A(n11135), .ZN(n11109) );
  INV_X1 U14019 ( .A(n11132), .ZN(n11110) );
  BUF_X2 U14020 ( .A(n11113), .Z(n11986) );
  INV_X1 U14021 ( .A(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11111) );
  OAI22_X1 U14022 ( .A1(n11112), .A2(n19308), .B1(n19453), .B2(n11111), .ZN(
        n11125) );
  INV_X1 U14023 ( .A(n18926), .ZN(n12221) );
  INV_X1 U14024 ( .A(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11117) );
  OR2_X1 U14025 ( .A1(n11221), .A2(n11117), .ZN(n11123) );
  NAND2_X2 U14026 ( .A1(n11120), .A2(n11119), .ZN(n11211) );
  NAND4_X1 U14027 ( .A1(n9812), .A2(n11123), .A3(n11122), .A4(n10944), .ZN(
        n11124) );
  NOR2_X1 U14028 ( .A1(n11125), .A2(n11124), .ZN(n11162) );
  INV_X1 U14029 ( .A(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11131) );
  INV_X1 U14030 ( .A(n11284), .ZN(n19256) );
  NAND2_X1 U14031 ( .A1(n19256), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n11130) );
  INV_X1 U14032 ( .A(n11219), .ZN(n13074) );
  NAND2_X1 U14033 ( .A1(n13074), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11129) );
  OAI211_X1 U14034 ( .C1(n19374), .C2(n11131), .A(n11130), .B(n11129), .ZN(
        n11144) );
  AND2_X1 U14035 ( .A1(n18926), .A2(n11132), .ZN(n11145) );
  INV_X1 U14036 ( .A(n11145), .ZN(n11133) );
  NAND2_X1 U14037 ( .A1(n19170), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n11142) );
  OR3_X2 U14038 ( .A1(n11146), .A2(n11148), .A3(n11133), .ZN(n11214) );
  INV_X1 U14039 ( .A(n11214), .ZN(n11134) );
  NAND2_X1 U14040 ( .A1(n11134), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n11141) );
  NAND2_X1 U14041 ( .A1(n11138), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n11139) );
  NAND4_X1 U14042 ( .A1(n11142), .A2(n11141), .A3(n11140), .A4(n11139), .ZN(
        n11143) );
  NOR2_X1 U14043 ( .A1(n11144), .A2(n11143), .ZN(n11161) );
  INV_X1 U14044 ( .A(n12999), .ZN(n11147) );
  NAND2_X1 U14045 ( .A1(n11147), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n11152) );
  NAND2_X1 U14046 ( .A1(n11152), .A2(n11151), .ZN(n11159) );
  INV_X1 U14047 ( .A(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11157) );
  INV_X1 U14048 ( .A(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11156) );
  NOR2_X1 U14049 ( .A1(n11159), .A2(n11158), .ZN(n11160) );
  INV_X1 U14050 ( .A(n11923), .ZN(n11922) );
  NOR2_X1 U14051 ( .A1(n11922), .A2(n11478), .ZN(n11163) );
  NAND2_X1 U14052 ( .A1(n11164), .A2(n11163), .ZN(n11482) );
  NAND2_X1 U14053 ( .A1(n11482), .A2(n11481), .ZN(n11166) );
  INV_X1 U14054 ( .A(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11167) );
  INV_X1 U14055 ( .A(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11168) );
  OAI22_X1 U14056 ( .A1(n11169), .A2(n11219), .B1(n11284), .B2(n11168), .ZN(
        n11170) );
  NOR2_X1 U14057 ( .A1(n11171), .A2(n11170), .ZN(n11193) );
  INV_X1 U14058 ( .A(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11173) );
  INV_X1 U14059 ( .A(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11172) );
  OAI22_X1 U14060 ( .A1(n11173), .A2(n19453), .B1(n12999), .B2(n11172), .ZN(
        n11177) );
  INV_X1 U14061 ( .A(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11174) );
  OAI22_X1 U14062 ( .A1(n11175), .A2(n19308), .B1(n11199), .B2(n11174), .ZN(
        n11176) );
  NOR2_X1 U14063 ( .A1(n11177), .A2(n11176), .ZN(n11192) );
  INV_X1 U14064 ( .A(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11179) );
  INV_X1 U14065 ( .A(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11178) );
  INV_X1 U14066 ( .A(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11181) );
  INV_X1 U14067 ( .A(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11180) );
  OAI22_X1 U14068 ( .A1(n11181), .A2(n11211), .B1(n19167), .B2(n11180), .ZN(
        n11182) );
  NOR2_X1 U14069 ( .A1(n11183), .A2(n11182), .ZN(n11191) );
  INV_X1 U14070 ( .A(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11185) );
  INV_X1 U14071 ( .A(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11184) );
  INV_X1 U14072 ( .A(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11187) );
  INV_X1 U14073 ( .A(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11186) );
  OAI22_X1 U14074 ( .A1(n11187), .A2(n19374), .B1(n11204), .B2(n11186), .ZN(
        n11188) );
  NOR2_X1 U14075 ( .A1(n11189), .A2(n11188), .ZN(n11190) );
  INV_X1 U14076 ( .A(n11240), .ZN(n11194) );
  NAND2_X1 U14077 ( .A1(n11194), .A2(n11164), .ZN(n11195) );
  INV_X1 U14078 ( .A(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11198) );
  OAI22_X1 U14079 ( .A1(n11198), .A2(n19374), .B1(n19308), .B2(n11197), .ZN(
        n11203) );
  INV_X1 U14080 ( .A(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11201) );
  INV_X1 U14081 ( .A(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11200) );
  OAI22_X1 U14082 ( .A1(n11201), .A2(n11199), .B1(n12999), .B2(n11200), .ZN(
        n11202) );
  NOR2_X1 U14083 ( .A1(n11203), .A2(n11202), .ZN(n11229) );
  INV_X1 U14084 ( .A(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11206) );
  INV_X1 U14085 ( .A(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11205) );
  OAI22_X1 U14086 ( .A1(n11206), .A2(n11204), .B1(n19420), .B2(n11205), .ZN(
        n11210) );
  INV_X1 U14087 ( .A(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11208) );
  INV_X1 U14088 ( .A(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11207) );
  OAI22_X1 U14089 ( .A1(n11208), .A2(n19340), .B1(n19453), .B2(n11207), .ZN(
        n11209) );
  NOR2_X1 U14090 ( .A1(n11210), .A2(n11209), .ZN(n11228) );
  INV_X1 U14091 ( .A(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11213) );
  INV_X1 U14092 ( .A(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11212) );
  OAI22_X1 U14093 ( .A1(n11213), .A2(n11211), .B1(n19167), .B2(n11212), .ZN(
        n11217) );
  INV_X1 U14094 ( .A(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11215) );
  INV_X1 U14095 ( .A(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12989) );
  OAI22_X1 U14096 ( .A1(n11215), .A2(n19098), .B1(n11214), .B2(n12989), .ZN(
        n11216) );
  NOR2_X1 U14097 ( .A1(n11217), .A2(n11216), .ZN(n11227) );
  INV_X1 U14098 ( .A(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11220) );
  OAI22_X1 U14099 ( .A1(n11220), .A2(n11218), .B1(n13078), .B2(n12270), .ZN(
        n11225) );
  INV_X1 U14100 ( .A(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11223) );
  INV_X1 U14101 ( .A(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11222) );
  OAI22_X1 U14102 ( .A1(n11223), .A2(n11284), .B1(n11221), .B2(n11222), .ZN(
        n11224) );
  NOR2_X1 U14103 ( .A1(n11225), .A2(n11224), .ZN(n11226) );
  NAND4_X1 U14104 ( .A1(n11229), .A2(n11228), .A3(n11227), .A4(n11226), .ZN(
        n11231) );
  NAND2_X1 U14105 ( .A1(n11242), .A2(n11164), .ZN(n11230) );
  NAND2_X1 U14106 ( .A1(n11231), .A2(n11230), .ZN(n11233) );
  NAND2_X1 U14107 ( .A1(n11490), .A2(n11233), .ZN(n11234) );
  INV_X1 U14108 ( .A(n11307), .ZN(n11235) );
  INV_X1 U14109 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n12220) );
  INV_X1 U14110 ( .A(P2_EBX_REG_1__SCAN_IN), .ZN(n12212) );
  NAND2_X1 U14111 ( .A1(n12220), .A2(n12212), .ZN(n11236) );
  MUX2_X1 U14112 ( .A(n11478), .B(n11236), .S(n12986), .Z(n11256) );
  NOR2_X1 U14113 ( .A1(n11481), .A2(n11476), .ZN(n11238) );
  NOR2_X1 U14114 ( .A1(n11238), .A2(n11237), .ZN(n11453) );
  MUX2_X1 U14115 ( .A(P2_EBX_REG_2__SCAN_IN), .B(n11453), .S(n11354), .Z(
        n11251) );
  MUX2_X1 U14116 ( .A(n11240), .B(n11239), .S(n11476), .Z(n11457) );
  INV_X1 U14117 ( .A(P2_EBX_REG_3__SCAN_IN), .ZN(n12969) );
  MUX2_X1 U14118 ( .A(n11457), .B(n12969), .S(n12986), .Z(n11249) );
  INV_X1 U14119 ( .A(n11456), .ZN(n11241) );
  MUX2_X1 U14120 ( .A(n11241), .B(P2_EBX_REG_4__SCAN_IN), .S(n12986), .Z(
        n11261) );
  MUX2_X1 U14121 ( .A(n11242), .B(P2_EBX_REG_5__SCAN_IN), .S(n12986), .Z(
        n11243) );
  AND2_X1 U14122 ( .A1(n11244), .A2(n11243), .ZN(n11245) );
  OR2_X1 U14123 ( .A1(n11245), .A2(n11301), .ZN(n18884) );
  NAND2_X1 U14124 ( .A1(n11246), .A2(n18884), .ZN(n11265) );
  INV_X1 U14125 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n16146) );
  XNOR2_X1 U14126 ( .A(n11265), .B(n16146), .ZN(n16045) );
  NAND2_X1 U14127 ( .A1(n9810), .A2(n11247), .ZN(n11248) );
  OAI21_X1 U14128 ( .B1(n11250), .B2(n11249), .A(n11262), .ZN(n12965) );
  XNOR2_X1 U14129 ( .A(n11256), .B(n11251), .ZN(n13029) );
  XNOR2_X1 U14130 ( .A(n13029), .B(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11955) );
  MUX2_X1 U14131 ( .A(n11922), .B(n11252), .S(n11476), .Z(n11455) );
  INV_X1 U14132 ( .A(n11455), .ZN(n11253) );
  MUX2_X1 U14133 ( .A(n11253), .B(P2_EBX_REG_0__SCAN_IN), .S(n12986), .Z(
        n18915) );
  NAND2_X1 U14134 ( .A1(n18915), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n11928) );
  AND2_X1 U14135 ( .A1(P2_EBX_REG_1__SCAN_IN), .A2(P2_EBX_REG_0__SCAN_IN), 
        .ZN(n11254) );
  NAND2_X1 U14136 ( .A1(n12986), .A2(n11254), .ZN(n11255) );
  NAND2_X1 U14137 ( .A1(n11256), .A2(n11255), .ZN(n13173) );
  OAI21_X1 U14138 ( .B1(n9972), .B2(n11928), .A(n13173), .ZN(n11258) );
  NAND2_X1 U14139 ( .A1(n11928), .A2(n9972), .ZN(n11257) );
  AND2_X1 U14140 ( .A1(n11258), .A2(n11257), .ZN(n11954) );
  NAND2_X1 U14141 ( .A1(n11955), .A2(n11954), .ZN(n11953) );
  INV_X1 U14142 ( .A(n13029), .ZN(n11259) );
  NAND2_X1 U14143 ( .A1(n11259), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11260) );
  AND2_X1 U14144 ( .A1(n11953), .A2(n11260), .ZN(n12924) );
  XNOR2_X1 U14145 ( .A(n11262), .B(n11261), .ZN(n11263) );
  INV_X1 U14146 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n16147) );
  XNOR2_X1 U14147 ( .A(n11263), .B(n16147), .ZN(n12822) );
  INV_X1 U14148 ( .A(n11263), .ZN(n18896) );
  NAND2_X1 U14149 ( .A1(n18896), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11264) );
  NAND2_X1 U14150 ( .A1(n11265), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11266) );
  INV_X1 U14151 ( .A(n11297), .ZN(n11295) );
  OAI22_X1 U14152 ( .A1(n10810), .A2(n19374), .B1(n11204), .B2(n11267), .ZN(
        n11270) );
  INV_X1 U14153 ( .A(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11268) );
  OAI22_X1 U14154 ( .A1(n11268), .A2(n19340), .B1(n12999), .B2(n20775), .ZN(
        n11269) );
  NOR2_X1 U14155 ( .A1(n11270), .A2(n11269), .ZN(n11291) );
  INV_X1 U14156 ( .A(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11271) );
  OAI22_X1 U14157 ( .A1(n11272), .A2(n19308), .B1(n19453), .B2(n11271), .ZN(
        n11276) );
  INV_X1 U14158 ( .A(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11274) );
  INV_X1 U14159 ( .A(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11273) );
  OAI22_X1 U14160 ( .A1(n11274), .A2(n11199), .B1(n19420), .B2(n11273), .ZN(
        n11275) );
  NOR2_X1 U14161 ( .A1(n11276), .A2(n11275), .ZN(n11290) );
  INV_X1 U14162 ( .A(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11278) );
  INV_X1 U14163 ( .A(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11277) );
  OAI22_X1 U14164 ( .A1(n11278), .A2(n11211), .B1(n19167), .B2(n11277), .ZN(
        n11282) );
  INV_X1 U14165 ( .A(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11280) );
  INV_X1 U14166 ( .A(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11279) );
  OAI22_X1 U14167 ( .A1(n11280), .A2(n19098), .B1(n11214), .B2(n11279), .ZN(
        n11281) );
  NOR2_X1 U14168 ( .A1(n11282), .A2(n11281), .ZN(n11289) );
  OAI22_X1 U14169 ( .A1(n19094), .A2(n13078), .B1(n11218), .B2(n10817), .ZN(
        n11287) );
  INV_X1 U14170 ( .A(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11285) );
  INV_X1 U14171 ( .A(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11283) );
  OAI22_X1 U14172 ( .A1(n11285), .A2(n11284), .B1(n11221), .B2(n11283), .ZN(
        n11286) );
  NOR2_X1 U14173 ( .A1(n11287), .A2(n11286), .ZN(n11288) );
  NAND4_X1 U14174 ( .A1(n11291), .A2(n11290), .A3(n11289), .A4(n11288), .ZN(
        n11294) );
  INV_X1 U14175 ( .A(n11299), .ZN(n11292) );
  NAND2_X1 U14176 ( .A1(n11292), .A2(n11164), .ZN(n11293) );
  NAND2_X1 U14177 ( .A1(n11295), .A2(n11296), .ZN(n11503) );
  INV_X1 U14178 ( .A(n11296), .ZN(n11494) );
  NAND2_X1 U14179 ( .A1(n11297), .A2(n11494), .ZN(n11298) );
  NAND2_X2 U14180 ( .A1(n11503), .A2(n11298), .ZN(n11498) );
  INV_X1 U14181 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n12279) );
  MUX2_X1 U14182 ( .A(n11299), .B(n12279), .S(n12986), .Z(n11300) );
  NOR2_X1 U14183 ( .A1(n11301), .A2(n11300), .ZN(n11302) );
  OR2_X1 U14184 ( .A1(n11311), .A2(n11302), .ZN(n18872) );
  OAI21_X2 U14185 ( .B1(n11498), .B2(n11307), .A(n18872), .ZN(n11303) );
  INV_X1 U14186 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n20739) );
  XNOR2_X1 U14187 ( .A(n11303), .B(n20739), .ZN(n13272) );
  NAND2_X1 U14188 ( .A1(n13273), .A2(n13272), .ZN(n11305) );
  NAND2_X1 U14189 ( .A1(n11303), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11304) );
  NAND2_X1 U14190 ( .A1(n11305), .A2(n11304), .ZN(n15042) );
  INV_X1 U14191 ( .A(n15042), .ZN(n11312) );
  INV_X1 U14192 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n11306) );
  MUX2_X1 U14193 ( .A(n11307), .B(n11306), .S(n12986), .Z(n11309) );
  AND2_X1 U14194 ( .A1(n12986), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n11308) );
  XNOR2_X1 U14195 ( .A(n11316), .B(n11308), .ZN(n18845) );
  AND2_X1 U14196 ( .A1(n11307), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11508) );
  NAND2_X1 U14197 ( .A1(n18845), .A2(n11508), .ZN(n15045) );
  INV_X1 U14198 ( .A(n11309), .ZN(n11310) );
  XNOR2_X1 U14199 ( .A(n11311), .B(n11310), .ZN(n18858) );
  NAND2_X1 U14200 ( .A1(n18858), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15062) );
  NAND2_X1 U14201 ( .A1(n18845), .A2(n11307), .ZN(n11313) );
  INV_X1 U14202 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n20738) );
  NAND2_X1 U14203 ( .A1(n11313), .A2(n20738), .ZN(n15046) );
  INV_X1 U14204 ( .A(n18858), .ZN(n11314) );
  INV_X1 U14205 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n15066) );
  NAND2_X1 U14206 ( .A1(n11314), .A2(n15066), .ZN(n15061) );
  AND2_X1 U14207 ( .A1(n15046), .A2(n15061), .ZN(n11315) );
  INV_X1 U14208 ( .A(P2_EBX_REG_8__SCAN_IN), .ZN(n12291) );
  AND2_X1 U14209 ( .A1(n12986), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n11317) );
  XNOR2_X1 U14210 ( .A(n11318), .B(n11317), .ZN(n18834) );
  AOI21_X1 U14211 ( .B1(n18834), .B2(n11307), .A(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15027) );
  NAND2_X1 U14212 ( .A1(n12986), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n11319) );
  INV_X1 U14213 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n12245) );
  MUX2_X1 U14214 ( .A(P2_EBX_REG_10__SCAN_IN), .B(n11319), .S(n11321), .Z(
        n11320) );
  NAND2_X1 U14215 ( .A1(n11320), .A2(n11418), .ZN(n18821) );
  INV_X1 U14216 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16134) );
  NAND2_X1 U14217 ( .A1(n11329), .A2(n16134), .ZN(n14859) );
  NAND2_X1 U14218 ( .A1(n12986), .A2(P2_EBX_REG_11__SCAN_IN), .ZN(n11322) );
  OR2_X1 U14219 ( .A1(n11323), .A2(n11322), .ZN(n11325) );
  INV_X1 U14220 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n18809) );
  INV_X1 U14221 ( .A(n11331), .ZN(n11324) );
  NAND2_X1 U14222 ( .A1(n11325), .A2(n11324), .ZN(n18811) );
  OR2_X1 U14223 ( .A1(n18811), .A2(n11235), .ZN(n11326) );
  INV_X1 U14224 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16013) );
  NAND2_X1 U14225 ( .A1(n11326), .A2(n16013), .ZN(n16010) );
  OR3_X1 U14226 ( .A1(n18811), .A2(n11235), .A3(n16013), .ZN(n16009) );
  AND2_X1 U14227 ( .A1(n11307), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11328) );
  NAND2_X1 U14228 ( .A1(n18834), .A2(n11328), .ZN(n14856) );
  OR2_X1 U14229 ( .A1(n16134), .A2(n11329), .ZN(n14858) );
  NAND2_X1 U14230 ( .A1(n14856), .A2(n14858), .ZN(n16008) );
  INV_X1 U14231 ( .A(n16008), .ZN(n11330) );
  AND2_X1 U14232 ( .A1(n16009), .A2(n11330), .ZN(n14847) );
  NAND2_X1 U14233 ( .A1(n12986), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n11332) );
  NAND2_X1 U14234 ( .A1(n10025), .A2(n11333), .ZN(n11334) );
  NAND2_X1 U14235 ( .A1(n11362), .A2(n11334), .ZN(n18799) );
  INV_X1 U14236 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n11335) );
  OR3_X1 U14237 ( .A1(n18799), .A2(n11235), .A3(n11335), .ZN(n14844) );
  NAND2_X1 U14238 ( .A1(n14847), .A2(n14844), .ZN(n14775) );
  OR2_X1 U14239 ( .A1(n18799), .A2(n11235), .ZN(n11336) );
  NAND2_X1 U14240 ( .A1(n11336), .A2(n11335), .ZN(n14845) );
  INV_X1 U14241 ( .A(P2_EBX_REG_14__SCAN_IN), .ZN(n12897) );
  INV_X1 U14242 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n13043) );
  NAND2_X1 U14243 ( .A1(n12897), .A2(n13043), .ZN(n11337) );
  AND2_X1 U14244 ( .A1(n12986), .A2(n11337), .ZN(n11338) );
  INV_X1 U14245 ( .A(P2_EBX_REG_16__SCAN_IN), .ZN(n11351) );
  INV_X1 U14246 ( .A(P2_EBX_REG_17__SCAN_IN), .ZN(n11339) );
  NAND2_X1 U14247 ( .A1(n11351), .A2(n11339), .ZN(n11340) );
  AND2_X1 U14248 ( .A1(n12986), .A2(n11340), .ZN(n11341) );
  INV_X1 U14249 ( .A(P2_EBX_REG_18__SCAN_IN), .ZN(n14627) );
  INV_X1 U14250 ( .A(P2_EBX_REG_19__SCAN_IN), .ZN(n11342) );
  NAND2_X1 U14251 ( .A1(n14627), .A2(n11342), .ZN(n11343) );
  NAND2_X1 U14252 ( .A1(n12986), .A2(n11343), .ZN(n11344) );
  INV_X1 U14253 ( .A(P2_EBX_REG_20__SCAN_IN), .ZN(n11345) );
  INV_X1 U14254 ( .A(P2_EBX_REG_21__SCAN_IN), .ZN(n11346) );
  INV_X1 U14255 ( .A(n11398), .ZN(n11350) );
  INV_X1 U14256 ( .A(n11347), .ZN(n11348) );
  NAND3_X1 U14257 ( .A1(n11348), .A2(P2_EBX_REG_21__SCAN_IN), .A3(n12986), 
        .ZN(n11349) );
  AND2_X1 U14258 ( .A1(n11350), .A2(n11349), .ZN(n18696) );
  NAND2_X1 U14259 ( .A1(n18696), .A2(n11307), .ZN(n11380) );
  INV_X1 U14260 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n14966) );
  NAND2_X1 U14261 ( .A1(n11380), .A2(n14966), .ZN(n14792) );
  INV_X1 U14262 ( .A(n11366), .ZN(n11352) );
  NAND2_X1 U14263 ( .A1(n11352), .A2(n11351), .ZN(n11368) );
  NAND3_X1 U14264 ( .A1(n11368), .A2(n12986), .A3(P2_EBX_REG_17__SCAN_IN), 
        .ZN(n11353) );
  INV_X1 U14265 ( .A(n11374), .ZN(n11373) );
  AOI21_X1 U14266 ( .B1(n18744), .B2(n11307), .A(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n14784) );
  NAND2_X1 U14267 ( .A1(n11364), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n11355) );
  MUX2_X1 U14268 ( .A(n11355), .B(n11364), .S(n11354), .Z(n11356) );
  OR2_X1 U14269 ( .A1(n11364), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n11359) );
  NAND2_X1 U14270 ( .A1(n11356), .A2(n11359), .ZN(n18778) );
  INV_X1 U14271 ( .A(n18778), .ZN(n11357) );
  NAND2_X1 U14272 ( .A1(n11357), .A2(n11307), .ZN(n11390) );
  AND2_X1 U14273 ( .A1(n12986), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n11358) );
  NAND2_X1 U14274 ( .A1(n11359), .A2(n11358), .ZN(n11360) );
  AND2_X1 U14275 ( .A1(n11360), .A2(n11366), .ZN(n18765) );
  AOI21_X1 U14276 ( .B1(n18765), .B2(n11307), .A(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n14779) );
  NAND2_X1 U14277 ( .A1(n11362), .A2(n11361), .ZN(n11363) );
  NAND2_X1 U14278 ( .A1(n11364), .A2(n11363), .ZN(n18788) );
  INV_X1 U14279 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n11598) );
  NOR4_X1 U14280 ( .A1(n14784), .A2(n14832), .A3(n14779), .A4(n15997), .ZN(
        n11371) );
  AND2_X1 U14281 ( .A1(n12986), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n11365) );
  INV_X1 U14282 ( .A(n11418), .ZN(n11408) );
  AOI21_X1 U14283 ( .B1(n11366), .B2(n11365), .A(n11408), .ZN(n11367) );
  NAND2_X1 U14284 ( .A1(n18753), .A2(n11307), .ZN(n11383) );
  XNOR2_X1 U14285 ( .A(n11383), .B(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n14825) );
  INV_X1 U14286 ( .A(n11369), .ZN(n11377) );
  AND2_X1 U14287 ( .A1(n12986), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n11370) );
  XNOR2_X1 U14288 ( .A(n11377), .B(n11370), .ZN(n11393) );
  INV_X1 U14289 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n11629) );
  OAI21_X1 U14290 ( .B1(n11393), .B2(n11235), .A(n11629), .ZN(n14791) );
  NAND4_X1 U14291 ( .A1(n14792), .A2(n11371), .A3(n14825), .A4(n14791), .ZN(
        n11379) );
  NAND2_X1 U14292 ( .A1(n11373), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n11372) );
  MUX2_X1 U14293 ( .A(n11373), .B(n11372), .S(n12986), .Z(n11375) );
  NAND2_X1 U14294 ( .A1(n11374), .A2(n14627), .ZN(n11376) );
  NAND2_X1 U14295 ( .A1(n11375), .A2(n11376), .ZN(n18732) );
  INV_X1 U14296 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n14989) );
  OAI21_X1 U14297 ( .B1(n18732), .B2(n11235), .A(n14989), .ZN(n15968) );
  NAND3_X1 U14298 ( .A1(n11376), .A2(n12986), .A3(P2_EBX_REG_19__SCAN_IN), 
        .ZN(n11378) );
  NAND2_X1 U14299 ( .A1(n11378), .A2(n11377), .ZN(n18719) );
  INV_X1 U14300 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n11625) );
  NAND2_X1 U14301 ( .A1(n11382), .A2(n11625), .ZN(n15970) );
  NAND2_X1 U14302 ( .A1(n15968), .A2(n15970), .ZN(n14787) );
  INV_X1 U14303 ( .A(n11380), .ZN(n11381) );
  NAND2_X1 U14304 ( .A1(n11381), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n14793) );
  NOR2_X1 U14305 ( .A1(n11382), .A2(n11625), .ZN(n15971) );
  INV_X1 U14306 ( .A(n11383), .ZN(n11384) );
  NAND2_X1 U14307 ( .A1(n11384), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n14781) );
  AND2_X1 U14308 ( .A1(n11307), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n11385) );
  NAND2_X1 U14309 ( .A1(n18744), .A2(n11385), .ZN(n14782) );
  AND2_X1 U14310 ( .A1(n11307), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n11386) );
  NAND2_X1 U14311 ( .A1(n18765), .A2(n11386), .ZN(n15987) );
  INV_X1 U14312 ( .A(n11387), .ZN(n11388) );
  NAND2_X1 U14313 ( .A1(n11388), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n14774) );
  NAND4_X1 U14314 ( .A1(n14781), .A2(n14782), .A3(n15987), .A4(n14774), .ZN(
        n11389) );
  NOR2_X1 U14315 ( .A1(n15971), .A2(n11389), .ZN(n11392) );
  INV_X1 U14316 ( .A(n11390), .ZN(n11391) );
  NAND2_X1 U14317 ( .A1(n11391), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n14833) );
  INV_X1 U14318 ( .A(n11393), .ZN(n18707) );
  AND2_X1 U14319 ( .A1(n11307), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n11394) );
  AND2_X1 U14320 ( .A1(n18707), .A2(n11394), .ZN(n14789) );
  NAND2_X1 U14321 ( .A1(n11307), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n11395) );
  NOR2_X1 U14322 ( .A1(n18732), .A2(n11395), .ZN(n14786) );
  NAND2_X1 U14323 ( .A1(n12986), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n11399) );
  NAND2_X1 U14324 ( .A1(n11400), .A2(n10018), .ZN(n11401) );
  NAND2_X1 U14325 ( .A1(n11407), .A2(n11401), .ZN(n15390) );
  NOR2_X1 U14326 ( .A1(n15390), .A2(n11235), .ZN(n11402) );
  XOR2_X1 U14327 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .B(n11402), .Z(
        n14953) );
  INV_X1 U14328 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n14956) );
  INV_X1 U14329 ( .A(n11402), .ZN(n11403) );
  NAND2_X1 U14330 ( .A1(n12986), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n11404) );
  XNOR2_X1 U14331 ( .A(n11407), .B(n11404), .ZN(n15914) );
  NAND2_X1 U14332 ( .A1(n15914), .A2(n11307), .ZN(n11405) );
  XNOR2_X1 U14333 ( .A(n11405), .B(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15954) );
  INV_X1 U14334 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15952) );
  OR2_X1 U14335 ( .A1(n11405), .A2(n15952), .ZN(n11406) );
  AND2_X1 U14336 ( .A1(n12986), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n11409) );
  AOI21_X1 U14337 ( .B1(n11410), .B2(n11409), .A(n11408), .ZN(n11411) );
  NAND2_X1 U14338 ( .A1(n10019), .A2(n11411), .ZN(n15905) );
  INV_X1 U14339 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14946) );
  NOR2_X1 U14340 ( .A1(n11412), .A2(n14946), .ZN(n14939) );
  NAND2_X1 U14341 ( .A1(n11412), .A2(n14946), .ZN(n14940) );
  INV_X1 U14342 ( .A(P2_EBX_REG_25__SCAN_IN), .ZN(n14571) );
  NAND2_X1 U14343 ( .A1(n12986), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n11413) );
  OR2_X1 U14344 ( .A1(n11422), .A2(n11413), .ZN(n11414) );
  INV_X1 U14345 ( .A(P2_EBX_REG_26__SCAN_IN), .ZN(n15886) );
  NAND2_X1 U14346 ( .A1(n15886), .A2(n11422), .ZN(n14741) );
  INV_X1 U14347 ( .A(n11416), .ZN(n15885) );
  NOR2_X1 U14348 ( .A1(n15885), .A2(n11235), .ZN(n11417) );
  AND2_X1 U14349 ( .A1(n11307), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11415) );
  NAND2_X1 U14350 ( .A1(n11416), .A2(n11415), .ZN(n11426) );
  NAND2_X1 U14351 ( .A1(n12986), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n11419) );
  OAI21_X1 U14352 ( .B1(n11420), .B2(n11419), .A(n11418), .ZN(n11421) );
  INV_X1 U14353 ( .A(n15896), .ZN(n11423) );
  AOI21_X1 U14354 ( .B1(n11423), .B2(n11307), .A(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n14923) );
  INV_X1 U14355 ( .A(n11436), .ZN(n11424) );
  NAND2_X1 U14356 ( .A1(n12986), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n14740) );
  NAND2_X1 U14357 ( .A1(n12986), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n11427) );
  XNOR2_X1 U14358 ( .A(n14744), .B(n11427), .ZN(n15863) );
  NAND2_X1 U14359 ( .A1(n15863), .A2(n11307), .ZN(n14748) );
  NAND2_X1 U14360 ( .A1(n11307), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n11425) );
  NAND2_X1 U14361 ( .A1(n11426), .A2(n14921), .ZN(n14739) );
  INV_X1 U14362 ( .A(n14744), .ZN(n11428) );
  NAND2_X1 U14363 ( .A1(n11428), .A2(n11427), .ZN(n11431) );
  NAND2_X1 U14364 ( .A1(n12986), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n11429) );
  XNOR2_X1 U14365 ( .A(n11431), .B(n11429), .ZN(n15851) );
  AOI21_X1 U14366 ( .B1(n15851), .B2(n11307), .A(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14730) );
  NAND3_X1 U14367 ( .A1(n15851), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n11307), .ZN(n14728) );
  AND2_X1 U14368 ( .A1(n12986), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n11430) );
  NAND2_X1 U14369 ( .A1(n12986), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n11432) );
  XNOR2_X1 U14370 ( .A(n11434), .B(n11432), .ZN(n15842) );
  NAND2_X1 U14371 ( .A1(n15842), .A2(n11307), .ZN(n11433) );
  INV_X1 U14372 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14717) );
  NAND2_X1 U14373 ( .A1(n11433), .A2(n14717), .ZN(n14719) );
  NOR2_X1 U14374 ( .A1(n11433), .A2(n14717), .ZN(n14718) );
  NOR2_X1 U14375 ( .A1(n11434), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n11435) );
  MUX2_X1 U14376 ( .A(n11436), .B(n11435), .S(n12986), .Z(n15827) );
  NAND2_X1 U14377 ( .A1(n15827), .A2(n11307), .ZN(n11437) );
  XNOR2_X1 U14378 ( .A(n11437), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n11438) );
  NAND2_X1 U14379 ( .A1(n12976), .A2(n10944), .ZN(n11936) );
  NOR2_X1 U14380 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(P2_STATE_REG_2__SCAN_IN), 
        .ZN(n19625) );
  AOI211_X1 U14381 ( .C1(P2_STATE_REG_1__SCAN_IN), .C2(P2_STATE_REG_2__SCAN_IN), .A(P2_STATE_REG_0__SCAN_IN), .B(n19625), .ZN(n19741) );
  NAND2_X1 U14382 ( .A1(n19741), .A2(n19736), .ZN(n12960) );
  INV_X1 U14383 ( .A(n12960), .ZN(n11937) );
  NAND2_X1 U14384 ( .A1(n10391), .A2(n11937), .ZN(n11474) );
  AOI21_X1 U14385 ( .B1(n11440), .B2(n16176), .A(n10398), .ZN(n11441) );
  NAND2_X1 U14386 ( .A1(n11936), .A2(n11441), .ZN(n11473) );
  NAND2_X1 U14387 ( .A1(n11443), .A2(n11442), .ZN(n11444) );
  OR2_X1 U14388 ( .A1(n11445), .A2(n11444), .ZN(n11446) );
  NAND2_X1 U14389 ( .A1(n11861), .A2(n11446), .ZN(n11450) );
  NAND2_X1 U14390 ( .A1(n11447), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11448) );
  NAND2_X1 U14391 ( .A1(n11448), .A2(n16179), .ZN(n11950) );
  INV_X1 U14392 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n11946) );
  OAI21_X1 U14393 ( .B1(n9723), .B2(n11950), .A(n11946), .ZN(n19718) );
  INV_X1 U14394 ( .A(n19718), .ZN(n11449) );
  MUX2_X1 U14395 ( .A(n11450), .B(n11449), .S(P2_STATE2_REG_1__SCAN_IN), .Z(
        n19729) );
  INV_X1 U14396 ( .A(n11451), .ZN(n11452) );
  NAND2_X1 U14397 ( .A1(n11452), .A2(n10944), .ZN(n11464) );
  OAI21_X1 U14398 ( .B1(n11455), .B2(n11454), .A(n11453), .ZN(n11458) );
  NAND3_X1 U14399 ( .A1(n11458), .A2(n11457), .A3(n11456), .ZN(n11460) );
  AND2_X1 U14400 ( .A1(n11460), .A2(n11459), .ZN(n19726) );
  INV_X1 U14401 ( .A(n11461), .ZN(n11462) );
  NOR2_X1 U14402 ( .A1(n11451), .A2(n11462), .ZN(n19724) );
  NAND2_X1 U14403 ( .A1(n19726), .A2(n19724), .ZN(n11463) );
  OAI21_X1 U14404 ( .B1(n19729), .B2(n11464), .A(n11463), .ZN(n11688) );
  NOR2_X1 U14405 ( .A1(n16167), .A2(n12960), .ZN(n11465) );
  AND2_X1 U14406 ( .A1(n11468), .A2(n11465), .ZN(n11466) );
  NOR2_X1 U14407 ( .A1(n11467), .A2(n11466), .ZN(n11942) );
  MUX2_X1 U14408 ( .A(n11468), .B(n10391), .S(n11164), .Z(n11469) );
  NAND3_X1 U14409 ( .A1(n11469), .A2(n11861), .A3(n19736), .ZN(n11470) );
  NAND2_X1 U14410 ( .A1(n11942), .A2(n11470), .ZN(n11471) );
  NOR2_X1 U14411 ( .A1(n11688), .A2(n11471), .ZN(n11472) );
  OAI211_X1 U14412 ( .C1(n11936), .C2(n11474), .A(n11473), .B(n11472), .ZN(
        n11475) );
  NOR2_X1 U14413 ( .A1(n11451), .A2(n11476), .ZN(n19730) );
  NAND2_X1 U14414 ( .A1(n11690), .A2(n19065), .ZN(n11687) );
  INV_X1 U14415 ( .A(n11477), .ZN(n12933) );
  INV_X1 U14416 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n13195) );
  NOR3_X1 U14417 ( .A1(n11478), .A2(n11923), .A3(n13195), .ZN(n11480) );
  NOR2_X1 U14418 ( .A1(n11923), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n11479) );
  XNOR2_X1 U14419 ( .A(n11479), .B(n11478), .ZN(n11931) );
  NOR2_X1 U14420 ( .A1(n9972), .A2(n11931), .ZN(n11930) );
  NOR2_X1 U14421 ( .A1(n11480), .A2(n11930), .ZN(n11483) );
  XNOR2_X1 U14422 ( .A(n11482), .B(n11481), .ZN(n11960) );
  NAND2_X1 U14423 ( .A1(n9822), .A2(n11960), .ZN(n11959) );
  OR2_X1 U14424 ( .A1(n11483), .A2(n19067), .ZN(n11484) );
  NAND2_X1 U14425 ( .A1(n11959), .A2(n11484), .ZN(n11485) );
  XNOR2_X1 U14426 ( .A(n11485), .B(n12927), .ZN(n12932) );
  NAND2_X1 U14427 ( .A1(n12933), .A2(n12932), .ZN(n12934) );
  NAND2_X1 U14428 ( .A1(n11485), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11486) );
  NAND2_X1 U14429 ( .A1(n12934), .A2(n11486), .ZN(n12826) );
  INV_X1 U14430 ( .A(n11487), .ZN(n11488) );
  NAND2_X1 U14431 ( .A1(n11490), .A2(n11489), .ZN(n12824) );
  NAND2_X1 U14432 ( .A1(n11492), .A2(n16146), .ZN(n16046) );
  NAND2_X1 U14433 ( .A1(n11493), .A2(n16047), .ZN(n11500) );
  INV_X1 U14434 ( .A(n11493), .ZN(n11496) );
  INV_X1 U14435 ( .A(n16047), .ZN(n11495) );
  AOI21_X1 U14436 ( .B1(n11496), .B2(n11498), .A(n10265), .ZN(n11497) );
  OAI21_X1 U14437 ( .B1(n11500), .B2(n11498), .A(n11497), .ZN(n13271) );
  NAND2_X1 U14438 ( .A1(n13271), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11502) );
  INV_X1 U14439 ( .A(n11498), .ZN(n11499) );
  NAND2_X1 U14440 ( .A1(n11500), .A2(n11499), .ZN(n11501) );
  XNOR2_X1 U14441 ( .A(n11504), .B(n11307), .ZN(n15059) );
  NAND2_X1 U14442 ( .A1(n11505), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11506) );
  INV_X1 U14443 ( .A(n11508), .ZN(n11509) );
  NAND2_X2 U14444 ( .A1(n11511), .A2(n11510), .ZN(n14819) );
  INV_X1 U14445 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n16121) );
  NAND2_X1 U14446 ( .A1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16122) );
  NOR2_X1 U14447 ( .A1(n16121), .A2(n16122), .ZN(n15012) );
  INV_X1 U14448 ( .A(n15012), .ZN(n15013) );
  NOR2_X1 U14449 ( .A1(n11335), .A2(n11598), .ZN(n16103) );
  NAND2_X1 U14450 ( .A1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n16103), .ZN(
        n16091) );
  NOR2_X1 U14451 ( .A1(n15013), .A2(n16091), .ZN(n14996) );
  NAND2_X1 U14452 ( .A1(n14996), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15004) );
  NAND2_X1 U14453 ( .A1(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n14985) );
  INV_X1 U14454 ( .A(n14985), .ZN(n11512) );
  NAND2_X1 U14455 ( .A1(n11512), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n11513) );
  NOR2_X1 U14456 ( .A1(n15004), .A2(n11513), .ZN(n11672) );
  NAND2_X1 U14457 ( .A1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n11675) );
  INV_X1 U14458 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n14930) );
  INV_X1 U14459 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14895) );
  AOI222_X1 U14460 ( .A1(n11516), .A2(P2_REIP_REG_31__SCAN_IN), .B1(n11085), 
        .B2(P2_EAX_REG_31__SCAN_IN), .C1(n11515), .C2(
        P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n11517) );
  XNOR2_X1 U14461 ( .A(n11518), .B(n11517), .ZN(n15826) );
  NAND2_X1 U14462 ( .A1(n11520), .A2(n11519), .ZN(n15073) );
  INV_X1 U14463 ( .A(n15073), .ZN(n11521) );
  AND2_X1 U14464 ( .A1(n11522), .A2(n11521), .ZN(n13187) );
  INV_X1 U14465 ( .A(n13187), .ZN(n16171) );
  OAI21_X1 U14466 ( .B1(n10919), .B2(n11164), .A(n16171), .ZN(n11523) );
  NOR2_X1 U14467 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19606) );
  NAND2_X1 U14468 ( .A1(n19606), .A2(n19744), .ZN(n18675) );
  INV_X1 U14469 ( .A(n18675), .ZN(n11862) );
  AND2_X2 U14470 ( .A1(n11862), .A2(n18954), .ZN(n19033) );
  INV_X1 U14471 ( .A(n19033), .ZN(n18846) );
  INV_X1 U14472 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n19672) );
  NOR2_X1 U14473 ( .A1(n18846), .A2(n19672), .ZN(n11701) );
  NAND2_X1 U14474 ( .A1(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14911) );
  NAND2_X1 U14475 ( .A1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n16072) );
  NAND2_X1 U14476 ( .A1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n15049) );
  NAND2_X1 U14477 ( .A1(n11668), .A2(n16169), .ZN(n19047) );
  INV_X1 U14478 ( .A(n19047), .ZN(n14995) );
  NOR2_X1 U14479 ( .A1(n9972), .A2(n13195), .ZN(n19052) );
  INV_X1 U14480 ( .A(n19052), .ZN(n19046) );
  NAND2_X1 U14481 ( .A1(n19067), .A2(n19046), .ZN(n11540) );
  NAND2_X1 U14482 ( .A1(n11524), .A2(n11525), .ZN(n11537) );
  NAND2_X1 U14483 ( .A1(n10247), .A2(n10398), .ZN(n11527) );
  INV_X1 U14484 ( .A(n11526), .ZN(n11863) );
  AOI22_X1 U14485 ( .A1(n11527), .A2(n11863), .B1(n10391), .B2(n19740), .ZN(
        n11529) );
  AND3_X1 U14486 ( .A1(n11530), .A2(n11529), .A3(n11528), .ZN(n11536) );
  NAND2_X1 U14487 ( .A1(n11531), .A2(n10390), .ZN(n11532) );
  NAND2_X1 U14488 ( .A1(n11532), .A2(n10944), .ZN(n15074) );
  NAND2_X1 U14489 ( .A1(n15074), .A2(n11533), .ZN(n11534) );
  NAND2_X1 U14490 ( .A1(n11534), .A2(n10389), .ZN(n11535) );
  AND3_X1 U14491 ( .A1(n11537), .A2(n11536), .A3(n11535), .ZN(n15072) );
  INV_X1 U14492 ( .A(n11538), .ZN(n15093) );
  NAND2_X1 U14493 ( .A1(n15072), .A2(n15093), .ZN(n11539) );
  NAND2_X1 U14494 ( .A1(n11668), .A2(n11539), .ZN(n19048) );
  INV_X1 U14495 ( .A(n19048), .ZN(n19053) );
  AND2_X1 U14496 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n19052), .ZN(
        n11667) );
  AOI22_X1 U14497 ( .A1(n14995), .A2(n11540), .B1(n19053), .B2(n11667), .ZN(
        n12926) );
  NAND3_X1 U14498 ( .A1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n11670) );
  NOR2_X1 U14499 ( .A1(n12926), .A2(n11670), .ZN(n13275) );
  NAND2_X1 U14500 ( .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n13275), .ZN(
        n15067) );
  NOR2_X1 U14501 ( .A1(n15049), .A2(n15067), .ZN(n14984) );
  NAND2_X1 U14502 ( .A1(n14984), .A2(n11672), .ZN(n16080) );
  NOR2_X1 U14503 ( .A1(n16080), .A2(n11675), .ZN(n14967) );
  NAND2_X1 U14504 ( .A1(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n14967), .ZN(
        n14955) );
  NOR2_X1 U14505 ( .A1(n16072), .A2(n14955), .ZN(n14945) );
  NAND2_X1 U14506 ( .A1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n14945), .ZN(
        n14931) );
  NOR2_X1 U14507 ( .A1(n14911), .A2(n14931), .ZN(n14883) );
  INV_X1 U14508 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14904) );
  INV_X1 U14509 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n11656) );
  NOR3_X1 U14510 ( .A1(n14895), .A2(n14904), .A3(n11656), .ZN(n11678) );
  NAND2_X1 U14511 ( .A1(n14883), .A2(n11678), .ZN(n14868) );
  NOR3_X1 U14512 ( .A1(n14717), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n14868), .ZN(n11541) );
  AOI211_X1 U14513 ( .C1(n15826), .C2(n19059), .A(n11701), .B(n11541), .ZN(
        n11683) );
  INV_X1 U14514 ( .A(n11544), .ZN(n11546) );
  NAND2_X1 U14515 ( .A1(n11546), .A2(n11545), .ZN(n11547) );
  OR2_X1 U14516 ( .A1(n10455), .A2(n16147), .ZN(n11554) );
  NAND2_X1 U14517 ( .A1(n10456), .A2(P2_EBX_REG_4__SCAN_IN), .ZN(n11550) );
  NAND2_X1 U14518 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n11549) );
  OAI211_X1 U14519 ( .C1(n11659), .C2(n11551), .A(n11550), .B(n11549), .ZN(
        n11552) );
  INV_X1 U14520 ( .A(n11552), .ZN(n11553) );
  OR2_X1 U14521 ( .A1(n10455), .A2(n16146), .ZN(n11560) );
  NAND2_X1 U14522 ( .A1(n10456), .A2(P2_EBX_REG_5__SCAN_IN), .ZN(n11556) );
  NAND2_X1 U14523 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n11555) );
  OAI211_X1 U14524 ( .C1(n11659), .C2(n11557), .A(n11556), .B(n11555), .ZN(
        n11558) );
  INV_X1 U14525 ( .A(n11558), .ZN(n11559) );
  OR2_X1 U14526 ( .A1(n10455), .A2(n20739), .ZN(n11567) );
  NAND2_X1 U14527 ( .A1(n11599), .A2(P2_EBX_REG_6__SCAN_IN), .ZN(n11563) );
  NAND2_X1 U14528 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n11562) );
  OAI211_X1 U14529 ( .C1(n11659), .C2(n11564), .A(n11563), .B(n11562), .ZN(
        n11565) );
  INV_X1 U14530 ( .A(n11565), .ZN(n11566) );
  OR2_X1 U14531 ( .A1(n10455), .A2(n15066), .ZN(n11573) );
  INV_X1 U14532 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n11570) );
  NAND2_X1 U14533 ( .A1(n11599), .A2(P2_EBX_REG_7__SCAN_IN), .ZN(n11569) );
  NAND2_X1 U14534 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n11568) );
  OAI211_X1 U14535 ( .C1(n11659), .C2(n11570), .A(n11569), .B(n11568), .ZN(
        n11571) );
  INV_X1 U14536 ( .A(n11571), .ZN(n11572) );
  OR2_X1 U14537 ( .A1(n11662), .A2(n20738), .ZN(n11575) );
  AOI22_X1 U14538 ( .A1(n11599), .A2(P2_EBX_REG_8__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11574) );
  OAI211_X1 U14539 ( .C1(n11659), .C2(n11576), .A(n11575), .B(n11574), .ZN(
        n12286) );
  OR2_X1 U14540 ( .A1(n11662), .A2(n16121), .ZN(n11582) );
  NAND2_X1 U14541 ( .A1(n11599), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n11578) );
  NAND2_X1 U14542 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n11577) );
  OAI211_X1 U14543 ( .C1(n11659), .C2(n11579), .A(n11578), .B(n11577), .ZN(
        n11580) );
  INV_X1 U14544 ( .A(n11580), .ZN(n11581) );
  OR2_X1 U14545 ( .A1(n11662), .A2(n16134), .ZN(n11588) );
  NAND2_X1 U14546 ( .A1(n11599), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n11584) );
  NAND2_X1 U14547 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n11583) );
  OAI211_X1 U14548 ( .C1(n11659), .C2(n11585), .A(n11584), .B(n11583), .ZN(
        n11586) );
  INV_X1 U14549 ( .A(n11586), .ZN(n11587) );
  INV_X1 U14550 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n11591) );
  OR2_X1 U14551 ( .A1(n11662), .A2(n16013), .ZN(n11590) );
  AOI22_X1 U14552 ( .A1(n11599), .A2(P2_EBX_REG_11__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), 
        .ZN(n11589) );
  OAI211_X1 U14553 ( .C1(n11659), .C2(n11591), .A(n11590), .B(n11589), .ZN(
        n12495) );
  NAND2_X1 U14554 ( .A1(n12496), .A2(n12495), .ZN(n12514) );
  OR2_X1 U14555 ( .A1(n11662), .A2(n11335), .ZN(n11597) );
  NAND2_X1 U14556 ( .A1(n11599), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n11593) );
  NAND2_X1 U14557 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n11592) );
  OAI211_X1 U14558 ( .C1(n11659), .C2(n11594), .A(n11593), .B(n11592), .ZN(
        n11595) );
  INV_X1 U14559 ( .A(n11595), .ZN(n11596) );
  OR2_X1 U14560 ( .A1(n11662), .A2(n11598), .ZN(n11605) );
  INV_X1 U14561 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n11602) );
  NAND2_X1 U14562 ( .A1(n11599), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n11601) );
  NAND2_X1 U14563 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n11600) );
  OAI211_X1 U14564 ( .C1(n11659), .C2(n11602), .A(n11601), .B(n11600), .ZN(
        n11603) );
  INV_X1 U14565 ( .A(n11603), .ZN(n11604) );
  INV_X1 U14566 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n14839) );
  OR2_X1 U14567 ( .A1(n11662), .A2(n14839), .ZN(n11607) );
  AOI22_X1 U14568 ( .A1(n11599), .A2(P2_EBX_REG_14__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), 
        .ZN(n11606) );
  OAI211_X1 U14569 ( .C1(n11659), .C2(n11608), .A(n11607), .B(n11606), .ZN(
        n12893) );
  INV_X1 U14570 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n14820) );
  OR2_X1 U14571 ( .A1(n11662), .A2(n14820), .ZN(n11614) );
  NAND2_X1 U14572 ( .A1(n11599), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n11610) );
  NAND2_X1 U14573 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n11609) );
  OAI211_X1 U14574 ( .C1(n11659), .C2(n11611), .A(n11610), .B(n11609), .ZN(
        n11612) );
  INV_X1 U14575 ( .A(n11612), .ZN(n11613) );
  INV_X1 U14576 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n20745) );
  OR2_X1 U14577 ( .A1(n11662), .A2(n20745), .ZN(n11619) );
  NAND2_X1 U14578 ( .A1(n11599), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n11616) );
  NAND2_X1 U14579 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n11615) );
  OAI211_X1 U14580 ( .C1(n11659), .C2(n19647), .A(n11616), .B(n11615), .ZN(
        n11617) );
  INV_X1 U14581 ( .A(n11617), .ZN(n11618) );
  INV_X1 U14582 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n11622) );
  INV_X1 U14583 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n14821) );
  OR2_X1 U14584 ( .A1(n11662), .A2(n14821), .ZN(n11621) );
  AOI22_X1 U14585 ( .A1(n11599), .A2(P2_EBX_REG_17__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), 
        .ZN(n11620) );
  OAI211_X1 U14586 ( .C1(n11659), .C2(n11622), .A(n11621), .B(n11620), .ZN(
        n13298) );
  OR2_X1 U14587 ( .A1(n11662), .A2(n14989), .ZN(n11624) );
  AOI22_X1 U14588 ( .A1(n11599), .A2(P2_EBX_REG_18__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), 
        .ZN(n11623) );
  OAI211_X1 U14589 ( .C1(n11659), .C2(n19650), .A(n11624), .B(n11623), .ZN(
        n14623) );
  OR2_X1 U14590 ( .A1(n11662), .A2(n11625), .ZN(n11627) );
  AOI22_X1 U14591 ( .A1(n11599), .A2(P2_EBX_REG_19__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), 
        .ZN(n11626) );
  OAI211_X1 U14592 ( .C1(n11628), .C2(n11659), .A(n11627), .B(n11626), .ZN(
        n13393) );
  OR2_X1 U14593 ( .A1(n11662), .A2(n11629), .ZN(n11634) );
  NAND2_X1 U14594 ( .A1(n11599), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n11631) );
  NAND2_X1 U14595 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n11630) );
  OAI211_X1 U14596 ( .C1(n11659), .C2(n20777), .A(n11631), .B(n11630), .ZN(
        n11632) );
  INV_X1 U14597 ( .A(n11632), .ZN(n11633) );
  NAND2_X1 U14598 ( .A1(n11634), .A2(n11633), .ZN(n14617) );
  INV_X1 U14599 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n19654) );
  OR2_X1 U14600 ( .A1(n11662), .A2(n14966), .ZN(n11636) );
  AOI22_X1 U14601 ( .A1(n11599), .A2(P2_EBX_REG_21__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), 
        .ZN(n11635) );
  OAI211_X1 U14602 ( .C1(n11659), .C2(n19654), .A(n11636), .B(n11635), .ZN(
        n14606) );
  OR2_X1 U14603 ( .A1(n11662), .A2(n14956), .ZN(n11638) );
  AOI22_X1 U14604 ( .A1(n11599), .A2(P2_EBX_REG_22__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), 
        .ZN(n11637) );
  OAI211_X1 U14605 ( .C1(n11659), .C2(n19656), .A(n11638), .B(n11637), .ZN(
        n14594) );
  INV_X1 U14606 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n11641) );
  OR2_X1 U14607 ( .A1(n11662), .A2(n15952), .ZN(n11640) );
  AOI22_X1 U14608 ( .A1(n11599), .A2(P2_EBX_REG_23__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), 
        .ZN(n11639) );
  OAI211_X1 U14609 ( .C1(n11659), .C2(n11641), .A(n11640), .B(n11639), .ZN(
        n14587) );
  INV_X1 U14610 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n19659) );
  OR2_X1 U14611 ( .A1(n11662), .A2(n14946), .ZN(n11643) );
  AOI22_X1 U14612 ( .A1(n11599), .A2(P2_EBX_REG_24__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), 
        .ZN(n11642) );
  OAI211_X1 U14613 ( .C1(n11659), .C2(n19659), .A(n11643), .B(n11642), .ZN(
        n14578) );
  INV_X1 U14614 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n11646) );
  OR2_X1 U14615 ( .A1(n11662), .A2(n14930), .ZN(n11645) );
  AOI22_X1 U14616 ( .A1(n11599), .A2(P2_EBX_REG_25__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), 
        .ZN(n11644) );
  OAI211_X1 U14617 ( .C1(n11659), .C2(n11646), .A(n11645), .B(n11644), .ZN(
        n14566) );
  INV_X1 U14618 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n11647) );
  OR2_X1 U14619 ( .A1(n11662), .A2(n11647), .ZN(n11649) );
  AOI22_X1 U14620 ( .A1(n11599), .A2(P2_EBX_REG_26__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), 
        .ZN(n11648) );
  OAI211_X1 U14621 ( .C1(n11659), .C2(n20880), .A(n11649), .B(n11648), .ZN(
        n14558) );
  INV_X1 U14622 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n14759) );
  OR2_X1 U14623 ( .A1(n11662), .A2(n14904), .ZN(n11651) );
  AOI22_X1 U14624 ( .A1(n11599), .A2(P2_EBX_REG_27__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), 
        .ZN(n11650) );
  OAI211_X1 U14625 ( .C1(n11659), .C2(n14759), .A(n11651), .B(n11650), .ZN(
        n14551) );
  INV_X1 U14626 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n19664) );
  OR2_X1 U14627 ( .A1(n11662), .A2(n14895), .ZN(n11653) );
  AOI22_X1 U14628 ( .A1(n11599), .A2(P2_EBX_REG_28__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), 
        .ZN(n11652) );
  OAI211_X1 U14629 ( .C1(n11659), .C2(n19664), .A(n11653), .B(n11652), .ZN(
        n14542) );
  AOI22_X1 U14630 ( .A1(n11599), .A2(P2_EBX_REG_29__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), 
        .ZN(n11655) );
  NAND2_X1 U14631 ( .A1(n11561), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n11654) );
  OAI211_X1 U14632 ( .C1(n11662), .C2(n11656), .A(n11655), .B(n11654), .ZN(
        n14532) );
  INV_X1 U14633 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n19670) );
  OR2_X1 U14634 ( .A1(n11662), .A2(n14717), .ZN(n11658) );
  AOI22_X1 U14635 ( .A1(n11599), .A2(P2_EBX_REG_30__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), 
        .ZN(n11657) );
  OAI211_X1 U14636 ( .C1(n11659), .C2(n19670), .A(n11658), .B(n11657), .ZN(
        n11710) );
  INV_X1 U14637 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n12949) );
  AOI22_X1 U14638 ( .A1(n11599), .A2(P2_EBX_REG_31__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n11661) );
  NAND2_X1 U14639 ( .A1(n11561), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n11660) );
  OAI211_X1 U14640 ( .C1(n11662), .C2(n12949), .A(n11661), .B(n11660), .ZN(
        n11663) );
  INV_X1 U14641 ( .A(n11663), .ZN(n11664) );
  XNOR2_X2 U14642 ( .A(n11665), .B(n11664), .ZN(n15841) );
  NAND2_X1 U14643 ( .A1(n11668), .A2(n11666), .ZN(n19061) );
  NOR2_X1 U14644 ( .A1(n19048), .A2(n11667), .ZN(n11669) );
  NOR2_X1 U14645 ( .A1(n11668), .A2(n19033), .ZN(n19049) );
  NOR3_X1 U14646 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n19052), .A3(
        n19047), .ZN(n19063) );
  OR3_X1 U14647 ( .A1(n11669), .A2(n19049), .A3(n19063), .ZN(n12929) );
  AOI221_X1 U14648 ( .B1(n14998), .B2(n20739), .C1(n14998), .C2(n11670), .A(
        n12929), .ZN(n15065) );
  NAND2_X1 U14649 ( .A1(n14998), .A2(n15049), .ZN(n11671) );
  INV_X1 U14650 ( .A(n11672), .ZN(n11673) );
  NAND2_X1 U14651 ( .A1(n14998), .A2(n11673), .ZN(n11674) );
  OAI21_X1 U14652 ( .B1(n11675), .B2(n14966), .A(n14998), .ZN(n11676) );
  NAND2_X1 U14653 ( .A1(n16079), .A2(n11676), .ZN(n16067) );
  AND2_X1 U14654 ( .A1(n14998), .A2(n16072), .ZN(n11677) );
  NOR2_X1 U14655 ( .A1(n16067), .A2(n11677), .ZN(n14943) );
  OAI21_X1 U14656 ( .B1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n16163), .A(
        n14943), .ZN(n14927) );
  AOI21_X1 U14657 ( .B1(n14998), .B2(n14911), .A(n14927), .ZN(n14905) );
  OAI21_X1 U14658 ( .B1(n16163), .B2(n11678), .A(n14905), .ZN(n14871) );
  NOR2_X1 U14659 ( .A1(n16163), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11679) );
  OAI21_X1 U14660 ( .B1(n14871), .B2(n11679), .A(
        P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n11680) );
  OAI21_X1 U14661 ( .B1(n15841), .B2(n19061), .A(n11680), .ZN(n11681) );
  INV_X1 U14662 ( .A(n11681), .ZN(n11682) );
  NAND2_X1 U14663 ( .A1(n11687), .A2(n11686), .ZN(P2_U3015) );
  NAND2_X1 U14664 ( .A1(n11688), .A2(n18949), .ZN(n11692) );
  INV_X1 U14665 ( .A(n11692), .ZN(n11689) );
  NAND2_X1 U14666 ( .A1(n11690), .A2(n16060), .ZN(n11707) );
  OR2_X1 U14667 ( .A1(n11692), .A2(n16176), .ZN(n11867) );
  OR2_X1 U14668 ( .A1(n19685), .A2(n19606), .ZN(n19705) );
  NAND2_X1 U14669 ( .A1(n19705), .A2(n18954), .ZN(n11693) );
  AND2_X1 U14670 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19706) );
  INV_X1 U14671 ( .A(n11694), .ZN(n11696) );
  INV_X1 U14672 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n12954) );
  NAND2_X1 U14673 ( .A1(n12954), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n11695) );
  NAND2_X1 U14674 ( .A1(n11696), .A2(n11695), .ZN(n11925) );
  NAND2_X1 U14675 ( .A1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n15403), .ZN(
        n15402) );
  INV_X1 U14676 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n18836) );
  INV_X1 U14677 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n15996) );
  INV_X1 U14678 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n15409) );
  INV_X1 U14679 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n15979) );
  INV_X1 U14680 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n18695) );
  NAND2_X1 U14681 ( .A1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n15394), .ZN(
        n15834) );
  INV_X1 U14682 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n15959) );
  INV_X1 U14683 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n15940) );
  INV_X1 U14684 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n15874) );
  INV_X1 U14685 ( .A(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n11698) );
  NOR2_X1 U14686 ( .A1(n19045), .A2(n12950), .ZN(n11700) );
  AOI211_X1 U14687 ( .C1(n19032), .C2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n11701), .B(n11700), .ZN(n11702) );
  OAI21_X1 U14688 ( .B1(n15841), .B2(n16058), .A(n11702), .ZN(n11703) );
  NAND2_X1 U14689 ( .A1(n11707), .A2(n11706), .ZN(P2_U2983) );
  INV_X1 U14690 ( .A(n12976), .ZN(n16172) );
  NAND2_X1 U14691 ( .A1(n16172), .A2(n13187), .ZN(n11943) );
  NAND2_X1 U14692 ( .A1(n11943), .A2(n15093), .ZN(n11708) );
  XNOR2_X1 U14693 ( .A(n14531), .B(n11710), .ZN(n15844) );
  INV_X2 U14694 ( .A(n14621), .ZN(n14602) );
  NAND2_X1 U14695 ( .A1(n14602), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n11711) );
  NOR2_X1 U14696 ( .A1(P2_BE_N_REG_0__SCAN_IN), .A2(P2_BE_N_REG_1__SCAN_IN), 
        .ZN(n11715) );
  NOR4_X1 U14697 ( .A1(P2_BE_N_REG_2__SCAN_IN), .A2(P2_BE_N_REG_3__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n11714) );
  NAND4_X1 U14698 ( .A1(P2_M_IO_N_REG_SCAN_IN), .A2(P2_W_R_N_REG_SCAN_IN), 
        .A3(n11715), .A4(n11714), .ZN(n11728) );
  NOR2_X1 U14699 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n11728), .ZN(n16367)
         );
  NOR4_X1 U14700 ( .A1(P1_ADDRESS_REG_14__SCAN_IN), .A2(
        P1_ADDRESS_REG_13__SCAN_IN), .A3(P1_ADDRESS_REG_12__SCAN_IN), .A4(
        P1_ADDRESS_REG_11__SCAN_IN), .ZN(n11719) );
  NOR4_X1 U14701 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(
        P1_ADDRESS_REG_17__SCAN_IN), .A3(P1_ADDRESS_REG_16__SCAN_IN), .A4(
        P1_ADDRESS_REG_15__SCAN_IN), .ZN(n11718) );
  NOR4_X1 U14702 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(
        P1_ADDRESS_REG_5__SCAN_IN), .A3(P1_ADDRESS_REG_4__SCAN_IN), .A4(
        P1_ADDRESS_REG_3__SCAN_IN), .ZN(n11717) );
  NOR4_X1 U14703 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(
        P1_ADDRESS_REG_9__SCAN_IN), .A3(P1_ADDRESS_REG_8__SCAN_IN), .A4(
        P1_ADDRESS_REG_7__SCAN_IN), .ZN(n11716) );
  AND4_X1 U14704 ( .A1(n11719), .A2(n11718), .A3(n11717), .A4(n11716), .ZN(
        n11724) );
  NOR4_X1 U14705 ( .A1(P1_ADDRESS_REG_1__SCAN_IN), .A2(
        P1_ADDRESS_REG_0__SCAN_IN), .A3(P1_ADDRESS_REG_20__SCAN_IN), .A4(
        P1_ADDRESS_REG_21__SCAN_IN), .ZN(n11722) );
  NOR4_X1 U14706 ( .A1(P1_ADDRESS_REG_24__SCAN_IN), .A2(
        P1_ADDRESS_REG_23__SCAN_IN), .A3(P1_ADDRESS_REG_22__SCAN_IN), .A4(
        P1_ADDRESS_REG_19__SCAN_IN), .ZN(n11721) );
  NOR4_X1 U14707 ( .A1(P1_ADDRESS_REG_28__SCAN_IN), .A2(
        P1_ADDRESS_REG_27__SCAN_IN), .A3(P1_ADDRESS_REG_26__SCAN_IN), .A4(
        P1_ADDRESS_REG_25__SCAN_IN), .ZN(n11720) );
  INV_X1 U14708 ( .A(P1_ADDRESS_REG_2__SCAN_IN), .ZN(n20601) );
  AND4_X1 U14709 ( .A1(n11722), .A2(n11721), .A3(n11720), .A4(n20601), .ZN(
        n11723) );
  NAND2_X1 U14710 ( .A1(n11724), .A2(n11723), .ZN(n11725) );
  AND2_X2 U14711 ( .A1(n11725), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n20006)
         );
  INV_X1 U14712 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n20663) );
  NOR3_X1 U14713 ( .A1(P1_BE_N_REG_0__SCAN_IN), .A2(P1_BE_N_REG_1__SCAN_IN), 
        .A3(n20663), .ZN(n11727) );
  NOR4_X1 U14714 ( .A1(P1_BE_N_REG_2__SCAN_IN), .A2(P1_BE_N_REG_3__SCAN_IN), 
        .A3(P1_D_C_N_REG_SCAN_IN), .A4(P1_ADS_N_REG_SCAN_IN), .ZN(n11726) );
  NAND4_X1 U14715 ( .A1(n20006), .A2(P1_M_IO_N_REG_SCAN_IN), .A3(n11727), .A4(
        n11726), .ZN(U214) );
  NOR2_X1 U14716 ( .A1(n14634), .A2(n11728), .ZN(n16290) );
  NAND2_X1 U14717 ( .A1(n16290), .A2(U214), .ZN(U212) );
  NAND2_X1 U14718 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(P3_REIP_REG_21__SCAN_IN), 
        .ZN(n16490) );
  INV_X1 U14719 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n18570) );
  INV_X1 U14720 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n18564) );
  INV_X1 U14721 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n18558) );
  NAND2_X1 U14722 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(P3_REIP_REG_15__SCAN_IN), 
        .ZN(n16547) );
  NOR2_X1 U14723 ( .A1(n18558), .A2(n16547), .ZN(n16519) );
  NAND3_X1 U14724 ( .A1(n16519), .A2(P3_REIP_REG_19__SCAN_IN), .A3(
        P3_REIP_REG_18__SCAN_IN), .ZN(n16508) );
  NOR2_X1 U14725 ( .A1(n18564), .A2(n16508), .ZN(n11847) );
  INV_X2 U14726 ( .A(n11805), .ZN(n16993) );
  AOI22_X1 U14727 ( .A1(n16993), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n16975), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11732) );
  NOR2_X2 U14728 ( .A1(n11736), .A2(n11733), .ZN(n15118) );
  AOI22_X1 U14729 ( .A1(n9726), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n16987), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11731) );
  AOI22_X1 U14730 ( .A1(n15318), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n16991), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11730) );
  INV_X2 U14731 ( .A(n16990), .ZN(n16969) );
  AOI22_X1 U14732 ( .A1(n16969), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n16974), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11729) );
  NAND4_X1 U14733 ( .A1(n11732), .A2(n11731), .A3(n11730), .A4(n11729), .ZN(
        n11743) );
  NOR2_X2 U14734 ( .A1(n11734), .A2(n11737), .ZN(n15149) );
  AOI22_X1 U14735 ( .A1(n17000), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n15162), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11741) );
  AOI22_X1 U14736 ( .A1(n9729), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n15279), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11740) );
  NOR2_X2 U14737 ( .A1(n11737), .A2(n18478), .ZN(n16986) );
  BUF_X2 U14738 ( .A(n16986), .Z(n16959) );
  AOI22_X1 U14739 ( .A1(n16968), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n16959), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11739) );
  NOR2_X2 U14740 ( .A1(n11737), .A2(n11736), .ZN(n11788) );
  AOI22_X1 U14741 ( .A1(n11754), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n16777), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11738) );
  NAND4_X1 U14742 ( .A1(n11741), .A2(n11740), .A3(n11739), .A4(n11738), .ZN(
        n11742) );
  INV_X1 U14743 ( .A(n16694), .ZN(n18012) );
  AOI22_X1 U14744 ( .A1(n9729), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n11754), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11744) );
  OAI21_X1 U14745 ( .B1(n20912), .B2(n9787), .A(n11744), .ZN(n11750) );
  INV_X2 U14746 ( .A(n16767), .ZN(n15279) );
  AOI22_X1 U14747 ( .A1(n16992), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n15279), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11748) );
  AOI22_X1 U14748 ( .A1(n16954), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n15286), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11747) );
  AOI22_X1 U14749 ( .A1(n16974), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n15254), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11746) );
  AOI22_X1 U14751 ( .A1(n16969), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n15318), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11745) );
  NAND4_X1 U14752 ( .A1(n11748), .A2(n11747), .A3(n11746), .A4(n11745), .ZN(
        n11749) );
  AOI22_X1 U14753 ( .A1(n15162), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n9726), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11764) );
  AOI22_X1 U14754 ( .A1(n11754), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n15254), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11763) );
  AOI22_X1 U14755 ( .A1(n15318), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n16974), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11755) );
  OAI21_X1 U14756 ( .B1(n11805), .B2(n20798), .A(n11755), .ZN(n11761) );
  AOI22_X1 U14757 ( .A1(n16954), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n16959), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11759) );
  AOI22_X1 U14758 ( .A1(n16988), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n9729), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11758) );
  AOI22_X1 U14759 ( .A1(n16968), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n15279), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11757) );
  AOI22_X1 U14760 ( .A1(n15294), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n16969), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11756) );
  NAND4_X1 U14761 ( .A1(n11759), .A2(n11758), .A3(n11757), .A4(n11756), .ZN(
        n11760) );
  AOI22_X1 U14762 ( .A1(n9726), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n16959), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11768) );
  AOI22_X1 U14763 ( .A1(n16993), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n9729), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11767) );
  AOI22_X1 U14764 ( .A1(n11754), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n16974), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11766) );
  AOI22_X1 U14765 ( .A1(n15162), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n16969), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11765) );
  NAND4_X1 U14766 ( .A1(n11768), .A2(n11767), .A3(n11766), .A4(n11765), .ZN(
        n11773) );
  AOI22_X1 U14767 ( .A1(n15294), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n16968), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11772) );
  AOI22_X1 U14768 ( .A1(n16954), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n15318), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11771) );
  AOI22_X1 U14769 ( .A1(n16992), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n15254), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11770) );
  AOI22_X1 U14770 ( .A1(n16988), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n15279), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11769) );
  AOI22_X1 U14771 ( .A1(n16993), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n11754), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11777) );
  AOI22_X1 U14772 ( .A1(n15162), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n9726), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11776) );
  AOI22_X1 U14773 ( .A1(n16992), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n16969), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11775) );
  AOI22_X1 U14774 ( .A1(n15294), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n15279), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11774) );
  NAND4_X1 U14775 ( .A1(n11777), .A2(n11776), .A3(n11775), .A4(n11774), .ZN(
        n11783) );
  AOI22_X1 U14776 ( .A1(n16959), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n16974), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11781) );
  AOI22_X1 U14777 ( .A1(n16988), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n9729), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11780) );
  AOI22_X1 U14778 ( .A1(n16968), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n15254), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11779) );
  AOI22_X1 U14779 ( .A1(n16954), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n11806), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11778) );
  NAND4_X1 U14780 ( .A1(n11781), .A2(n11780), .A3(n11779), .A4(n11778), .ZN(
        n11782) );
  AOI22_X1 U14781 ( .A1(n9729), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n15254), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11787) );
  AOI22_X1 U14782 ( .A1(n15162), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11806), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11786) );
  AOI22_X1 U14783 ( .A1(n16959), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n16974), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11785) );
  AOI22_X1 U14784 ( .A1(n16968), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n16969), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11784) );
  NAND4_X1 U14785 ( .A1(n11787), .A2(n11786), .A3(n11785), .A4(n11784), .ZN(
        n11794) );
  AOI22_X1 U14786 ( .A1(n16993), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n16987), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11792) );
  AOI22_X1 U14787 ( .A1(n11754), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n16777), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11791) );
  AOI22_X1 U14788 ( .A1(n9726), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n16975), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11790) );
  AOI22_X1 U14789 ( .A1(n15294), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n15279), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11789) );
  NAND4_X1 U14790 ( .A1(n11792), .A2(n11791), .A3(n11790), .A4(n11789), .ZN(
        n11793) );
  AOI22_X1 U14791 ( .A1(n11754), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n16987), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11798) );
  AOI22_X1 U14792 ( .A1(n15162), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n16974), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11797) );
  AOI22_X1 U14793 ( .A1(n16959), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n16777), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11796) );
  AOI22_X1 U14794 ( .A1(n16969), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n15318), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11795) );
  NAND4_X1 U14795 ( .A1(n11798), .A2(n11797), .A3(n11796), .A4(n11795), .ZN(
        n11804) );
  AOI22_X1 U14796 ( .A1(n15279), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n15254), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11802) );
  AOI22_X1 U14797 ( .A1(n15294), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n16968), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11801) );
  AOI22_X1 U14798 ( .A1(n9726), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n16975), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11800) );
  AOI22_X1 U14799 ( .A1(n16993), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n9729), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11799) );
  NAND4_X1 U14800 ( .A1(n11802), .A2(n11801), .A3(n11800), .A4(n11799), .ZN(
        n11803) );
  AOI22_X1 U14801 ( .A1(n16968), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n16987), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11816) );
  AOI22_X1 U14802 ( .A1(n15279), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n15254), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11815) );
  AOI22_X1 U14803 ( .A1(n16988), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11806), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11807) );
  OAI21_X1 U14804 ( .B1(n16990), .B2(n20836), .A(n11807), .ZN(n11813) );
  AOI22_X1 U14805 ( .A1(n9729), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n16777), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11811) );
  AOI22_X1 U14806 ( .A1(n15162), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n9726), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11810) );
  AOI22_X1 U14807 ( .A1(n15294), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n16974), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11809) );
  AOI22_X1 U14808 ( .A1(n11754), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n16986), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11808) );
  NAND4_X1 U14809 ( .A1(n11811), .A2(n11810), .A3(n11809), .A4(n11808), .ZN(
        n11812) );
  NAND2_X1 U14810 ( .A1(n15229), .A2(n17048), .ZN(n11822) );
  NOR4_X1 U14811 ( .A1(n16694), .A2(n13563), .A3(n18041), .A4(n11822), .ZN(
        n11817) );
  NAND2_X1 U14812 ( .A1(n15231), .A2(n11817), .ZN(n17239) );
  NAND2_X1 U14813 ( .A1(n16694), .A2(n18052), .ZN(n11830) );
  NAND2_X1 U14814 ( .A1(n11829), .A2(n18027), .ZN(n15207) );
  NAND2_X1 U14815 ( .A1(n17239), .A2(n15207), .ZN(n16380) );
  NAND2_X2 U14816 ( .A1(n18668), .A2(n16380), .ZN(n17200) );
  INV_X1 U14817 ( .A(n17239), .ZN(n17241) );
  NAND2_X1 U14818 ( .A1(n17241), .A2(n18023), .ZN(n11833) );
  NOR2_X1 U14819 ( .A1(n16694), .A2(n18023), .ZN(n11818) );
  NAND2_X1 U14820 ( .A1(n17048), .A2(n18041), .ZN(n18464) );
  NAND2_X1 U14821 ( .A1(n18052), .A2(n18464), .ZN(n15512) );
  NAND2_X1 U14822 ( .A1(n11818), .A2(n15512), .ZN(n15209) );
  NAND2_X1 U14823 ( .A1(n13564), .A2(n11822), .ZN(n15203) );
  NAND3_X1 U14824 ( .A1(n15231), .A2(n15209), .A3(n15203), .ZN(n11828) );
  INV_X1 U14825 ( .A(n11830), .ZN(n11827) );
  NAND2_X1 U14826 ( .A1(n16694), .A2(n18023), .ZN(n11819) );
  NAND2_X1 U14827 ( .A1(n15231), .A2(n11819), .ZN(n15204) );
  OAI21_X1 U14828 ( .B1(n18027), .B2(n18012), .A(n18464), .ZN(n11820) );
  INV_X1 U14829 ( .A(n11820), .ZN(n11821) );
  AOI21_X1 U14830 ( .B1(n11822), .B2(n15230), .A(n11821), .ZN(n11823) );
  AOI21_X1 U14831 ( .B1(n15230), .B2(n15204), .A(n11823), .ZN(n11826) );
  AOI21_X1 U14832 ( .B1(n18052), .B2(n15230), .A(n15229), .ZN(n11824) );
  INV_X1 U14833 ( .A(n11824), .ZN(n11825) );
  OAI211_X1 U14834 ( .C1(n11827), .C2(n18032), .A(n11826), .B(n11825), .ZN(
        n15208) );
  NAND2_X1 U14835 ( .A1(n11829), .A2(n15222), .ZN(n15218) );
  INV_X1 U14836 ( .A(n15218), .ZN(n18459) );
  NAND3_X1 U14837 ( .A1(n13564), .A2(n18453), .A3(n18046), .ZN(n13556) );
  NOR2_X1 U14838 ( .A1(n11830), .A2(n13556), .ZN(n11832) );
  NAND2_X1 U14839 ( .A1(n17200), .A2(n11833), .ZN(n11831) );
  AOI21_X4 U14840 ( .B1(n11832), .B2(n18654), .A(n11831), .ZN(n18458) );
  NAND2_X1 U14841 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18610), .ZN(n18504) );
  AOI22_X1 U14842 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n18288), .B1(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n18624), .ZN(n11834) );
  INV_X1 U14843 ( .A(n11834), .ZN(n13562) );
  XOR2_X1 U14844 ( .A(n13562), .B(n13558), .Z(n11845) );
  AOI22_X1 U14845 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B1(n18013), .B2(n18617), .ZN(
        n11839) );
  NOR2_X1 U14846 ( .A1(n11840), .A2(n11839), .ZN(n11836) );
  AOI22_X1 U14847 ( .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n16695), .B1(
        n11837), .B2(n18607), .ZN(n11843) );
  NOR2_X1 U14848 ( .A1(n11837), .A2(n18607), .ZN(n11842) );
  NAND2_X1 U14849 ( .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n16695), .ZN(
        n11838) );
  OAI22_X1 U14850 ( .A1(n11843), .A2(n18487), .B1(n11842), .B2(n11838), .ZN(
        n13557) );
  INV_X1 U14851 ( .A(n13557), .ZN(n11841) );
  XOR2_X1 U14852 ( .A(n11840), .B(n11839), .Z(n15228) );
  NAND2_X1 U14853 ( .A1(n11841), .A2(n15228), .ZN(n13560) );
  INV_X1 U14854 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n18009) );
  OR2_X1 U14855 ( .A1(n11842), .A2(n18487), .ZN(n11844) );
  AOI22_X1 U14856 ( .A1(n18009), .A2(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B1(
        n11844), .B2(n11843), .ZN(n13559) );
  NAND2_X1 U14857 ( .A1(n18012), .A2(n18669), .ZN(n11856) );
  INV_X1 U14858 ( .A(n11856), .ZN(n11846) );
  INV_X1 U14859 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n18519) );
  INV_X2 U14860 ( .A(n18663), .ZN(n18665) );
  OAI211_X1 U14861 ( .C1(P3_STATE_REG_2__SCAN_IN), .C2(P3_STATE_REG_1__SCAN_IN), .A(n18519), .B(n18579), .ZN(n18652) );
  NAND2_X1 U14862 ( .A1(READY22_REG_SCAN_IN), .A2(READY2), .ZN(n18655) );
  INV_X1 U14863 ( .A(n18655), .ZN(n18650) );
  AOI211_X1 U14864 ( .C1(n18654), .C2(n18652), .A(n18650), .B(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n18497) );
  INV_X1 U14865 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n18552) );
  INV_X1 U14866 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n18549) );
  INV_X1 U14867 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n18545) );
  INV_X1 U14868 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n18539) );
  INV_X1 U14869 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n18535) );
  INV_X1 U14870 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n18532) );
  NAND2_X1 U14871 ( .A1(P3_REIP_REG_2__SCAN_IN), .A2(P3_REIP_REG_1__SCAN_IN), 
        .ZN(n16732) );
  NOR2_X1 U14872 ( .A1(n18532), .A2(n16732), .ZN(n16699) );
  NAND2_X1 U14873 ( .A1(P3_REIP_REG_4__SCAN_IN), .A2(n16699), .ZN(n16684) );
  NOR2_X1 U14874 ( .A1(n18535), .A2(n16684), .ZN(n16672) );
  NAND2_X1 U14875 ( .A1(P3_REIP_REG_6__SCAN_IN), .A2(n16672), .ZN(n16653) );
  NOR2_X1 U14876 ( .A1(n18539), .A2(n16653), .ZN(n16642) );
  NAND2_X1 U14877 ( .A1(P3_REIP_REG_8__SCAN_IN), .A2(n16642), .ZN(n16617) );
  NAND2_X1 U14878 ( .A1(P3_REIP_REG_10__SCAN_IN), .A2(P3_REIP_REG_9__SCAN_IN), 
        .ZN(n16610) );
  NOR3_X1 U14879 ( .A1(n18545), .A2(n16617), .A3(n16610), .ZN(n16600) );
  NAND2_X1 U14880 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n16600), .ZN(n16586) );
  NOR3_X1 U14881 ( .A1(n18552), .A2(n18549), .A3(n16586), .ZN(n16572) );
  NAND2_X1 U14882 ( .A1(n16739), .A2(n16572), .ZN(n16566) );
  INV_X1 U14883 ( .A(n16566), .ZN(n16548) );
  NAND2_X1 U14884 ( .A1(n11847), .A2(n16548), .ZN(n16502) );
  NAND2_X1 U14885 ( .A1(n16572), .A2(n11847), .ZN(n16482) );
  NOR3_X1 U14886 ( .A1(n18570), .A2(n16482), .A3(n16490), .ZN(n16394) );
  INV_X1 U14887 ( .A(n16394), .ZN(n16474) );
  NOR2_X1 U14888 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n18667) );
  INV_X1 U14889 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n18596) );
  INV_X2 U14890 ( .A(n17993), .ZN(n17995) );
  NAND2_X1 U14891 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n18666), .ZN(n18505) );
  NOR2_X1 U14892 ( .A1(n18504), .A2(n18505), .ZN(n18499) );
  NOR4_X4 U14893 ( .A1(n17995), .A2(n18669), .A3(n9882), .A4(n18499), .ZN(
        n16737) );
  AOI21_X1 U14894 ( .B1(n16739), .B2(n16474), .A(n16737), .ZN(n16481) );
  AOI221_X1 U14895 ( .B1(n16490), .B2(n18570), .C1(n16502), .C2(n18570), .A(
        n16481), .ZN(n11860) );
  NOR2_X1 U14896 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n16738) );
  INV_X1 U14897 ( .A(P3_EBX_REG_2__SCAN_IN), .ZN(n16726) );
  NAND2_X1 U14898 ( .A1(n16738), .A2(n16726), .ZN(n16725) );
  NOR2_X1 U14899 ( .A1(P3_EBX_REG_3__SCAN_IN), .A2(n16725), .ZN(n16712) );
  NAND2_X1 U14900 ( .A1(n16712), .A2(n17020), .ZN(n16700) );
  NOR2_X1 U14901 ( .A1(P3_EBX_REG_5__SCAN_IN), .A2(n16700), .ZN(n16685) );
  INV_X1 U14902 ( .A(P3_EBX_REG_6__SCAN_IN), .ZN(n16674) );
  NAND2_X1 U14903 ( .A1(n16685), .A2(n16674), .ZN(n16673) );
  INV_X1 U14904 ( .A(P3_EBX_REG_8__SCAN_IN), .ZN(n16650) );
  NAND2_X1 U14905 ( .A1(n16658), .A2(n16650), .ZN(n16649) );
  INV_X1 U14906 ( .A(P3_EBX_REG_10__SCAN_IN), .ZN(n20809) );
  NAND2_X1 U14907 ( .A1(n16631), .A2(n20809), .ZN(n16628) );
  INV_X1 U14908 ( .A(P3_EBX_REG_12__SCAN_IN), .ZN(n16938) );
  NAND2_X1 U14909 ( .A1(n16611), .A2(n16938), .ZN(n16602) );
  INV_X1 U14910 ( .A(P3_EBX_REG_14__SCAN_IN), .ZN(n16579) );
  NAND2_X1 U14911 ( .A1(n16590), .A2(n16579), .ZN(n16578) );
  INV_X1 U14912 ( .A(P3_EBX_REG_16__SCAN_IN), .ZN(n16914) );
  NAND2_X1 U14913 ( .A1(n16560), .A2(n16914), .ZN(n16556) );
  INV_X1 U14914 ( .A(P3_EBX_REG_18__SCAN_IN), .ZN(n16887) );
  NAND2_X1 U14915 ( .A1(n16540), .A2(n16887), .ZN(n16529) );
  INV_X1 U14916 ( .A(P3_EBX_REG_20__SCAN_IN), .ZN(n15182) );
  NAND2_X1 U14917 ( .A1(n16520), .A2(n15182), .ZN(n16504) );
  NOR2_X1 U14918 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n16504), .ZN(n16496) );
  INV_X1 U14919 ( .A(P3_EBX_REG_22__SCAN_IN), .ZN(n16487) );
  NAND2_X1 U14920 ( .A1(n16496), .A2(n16487), .ZN(n16485) );
  NOR2_X1 U14921 ( .A1(P3_EBX_REG_23__SCAN_IN), .A2(n16485), .ZN(n16478) );
  INV_X1 U14922 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n18653) );
  NAND2_X1 U14923 ( .A1(P3_EBX_REG_31__SCAN_IN), .A2(n18023), .ZN(n11848) );
  AOI211_X4 U14924 ( .C1(n18653), .C2(n18655), .A(n11856), .B(n11848), .ZN(
        n16751) );
  AOI211_X1 U14925 ( .C1(P3_EBX_REG_23__SCAN_IN), .C2(n16485), .A(n16478), .B(
        n16711), .ZN(n11859) );
  INV_X1 U14926 ( .A(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n17378) );
  NAND2_X1 U14927 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n11849) );
  INV_X1 U14928 ( .A(n11849), .ZN(n17384) );
  INV_X1 U14929 ( .A(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n17389) );
  NAND2_X1 U14930 ( .A1(n17631), .A2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n17621) );
  NAND2_X1 U14931 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n17509) );
  NAND2_X1 U14932 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n17473) );
  NAND2_X1 U14933 ( .A1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n17453), .ZN(
        n17430) );
  NAND2_X1 U14934 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n17431) );
  NAND2_X1 U14935 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17423), .ZN(
        n17386) );
  NOR2_X1 U14936 ( .A1(n17389), .A2(n17386), .ZN(n11852) );
  NAND2_X1 U14937 ( .A1(n17384), .A2(n11852), .ZN(n17343) );
  INV_X1 U14938 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n17670) );
  NAND2_X1 U14939 ( .A1(n17423), .A2(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n17385) );
  NOR2_X1 U14940 ( .A1(n17670), .A2(n17352), .ZN(n16405) );
  AOI21_X1 U14941 ( .B1(n17378), .B2(n17343), .A(n16405), .ZN(n17374) );
  INV_X1 U14942 ( .A(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n17391) );
  NAND2_X1 U14943 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n11852), .ZN(
        n11851) );
  INV_X1 U14944 ( .A(n17343), .ZN(n11850) );
  AOI21_X1 U14945 ( .B1(n17391), .B2(n11851), .A(n11850), .ZN(n17394) );
  INV_X1 U14946 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n17409) );
  XNOR2_X1 U14947 ( .A(n17409), .B(n11852), .ZN(n17412) );
  AOI21_X1 U14948 ( .B1(n17389), .B2(n17386), .A(n11852), .ZN(n17425) );
  INV_X1 U14949 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n16430) );
  NAND2_X1 U14950 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n17353) );
  NAND2_X1 U14951 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n17314) );
  NAND2_X1 U14952 ( .A1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n16252), .ZN(
        n11853) );
  NOR2_X1 U14953 ( .A1(n17670), .A2(n17467), .ZN(n17468) );
  INV_X1 U14954 ( .A(n17468), .ZN(n11854) );
  NOR2_X1 U14955 ( .A1(n17473), .A2(n11854), .ZN(n16537) );
  NAND2_X1 U14956 ( .A1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n16537), .ZN(
        n16536) );
  NOR2_X1 U14957 ( .A1(n17670), .A2(n17533), .ZN(n16680) );
  NAND2_X1 U14958 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n16680), .ZN(
        n16666) );
  NOR3_X1 U14959 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n17544), .A3(
        n16666), .ZN(n16608) );
  NAND2_X1 U14960 ( .A1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n16608), .ZN(
        n16597) );
  NOR2_X1 U14961 ( .A1(n17472), .A2(n16597), .ZN(n16562) );
  NAND2_X1 U14962 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n16562), .ZN(
        n16549) );
  NOR2_X1 U14963 ( .A1(n17425), .A2(n16507), .ZN(n16506) );
  NOR2_X1 U14964 ( .A1(n16506), .A2(n16667), .ZN(n16495) );
  NOR2_X1 U14965 ( .A1(n16494), .A2(n16667), .ZN(n16484) );
  NOR2_X1 U14966 ( .A1(n17394), .A2(n16484), .ZN(n16483) );
  NOR2_X1 U14967 ( .A1(n16483), .A2(n16667), .ZN(n11855) );
  AOI211_X1 U14968 ( .C1(n17374), .C2(n11855), .A(n16406), .B(n9780), .ZN(
        n11858) );
  AOI211_X1 U14969 ( .C1(P3_EBX_REG_31__SCAN_IN), .C2(n18023), .A(n18497), .B(
        n11856), .ZN(n16681) );
  INV_X1 U14970 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n16812) );
  OAI22_X1 U14971 ( .A1(n17378), .A2(n16740), .B1(n16743), .B2(n16812), .ZN(
        n11857) );
  OR4_X1 U14972 ( .A1(n11860), .A2(n11859), .A3(n11858), .A4(n11857), .ZN(
        P3_U2648) );
  NAND2_X1 U14973 ( .A1(n11861), .A2(n18949), .ZN(n12962) );
  NOR2_X1 U14974 ( .A1(n12962), .A2(n10907), .ZN(n18913) );
  INV_X1 U14975 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .ZN(n19754) );
  NOR2_X1 U14976 ( .A1(n10425), .A2(n12962), .ZN(n12956) );
  NOR2_X1 U14977 ( .A1(n12956), .A2(n11862), .ZN(n11865) );
  OAI21_X1 U14978 ( .B1(n18913), .B2(n19754), .A(n11865), .ZN(P2_U2814) );
  NOR2_X1 U14979 ( .A1(n18913), .A2(P2_READREQUEST_REG_SCAN_IN), .ZN(n11864)
         );
  AOI22_X1 U14980 ( .A1(n11865), .A2(n11864), .B1(n19735), .B2(n11863), .ZN(
        P2_U3612) );
  INV_X1 U14981 ( .A(n11939), .ZN(n11866) );
  NOR3_X1 U14982 ( .A1(n11866), .A2(n11938), .A3(n11937), .ZN(n16173) );
  NOR2_X1 U14983 ( .A1(n16173), .A2(n19607), .ZN(n19733) );
  OAI21_X1 U14984 ( .B1(n19733), .B2(n11946), .A(n11867), .ZN(P2_U2819) );
  INV_X1 U14985 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n12890) );
  NAND2_X1 U14986 ( .A1(n12956), .A2(n11164), .ZN(n18951) );
  INV_X1 U14987 ( .A(P2_LWORD_REG_15__SCAN_IN), .ZN(n11870) );
  OAI21_X1 U14988 ( .B1(n11164), .B2(n19736), .A(n12956), .ZN(n11880) );
  INV_X1 U14989 ( .A(n11880), .ZN(n11882) );
  AND2_X1 U14990 ( .A1(n10944), .A2(n19736), .ZN(n11868) );
  AND2_X1 U14991 ( .A1(n12956), .A2(n11868), .ZN(n19024) );
  INV_X1 U14992 ( .A(n19024), .ZN(n11869) );
  AOI22_X1 U14993 ( .A1(n12980), .A2(BUF1_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n11897), .ZN(n12887) );
  OAI222_X1 U14994 ( .A1(n12890), .A2(n18951), .B1(n11870), .B2(n11882), .C1(
        n11869), .C2(n12887), .ZN(P2_U2982) );
  INV_X2 U14995 ( .A(n18951), .ZN(n19029) );
  AOI22_X1 U14996 ( .A1(n19029), .A2(P2_EAX_REG_26__SCAN_IN), .B1(n11880), 
        .B2(P2_UWORD_REG_10__SCAN_IN), .ZN(n11874) );
  INV_X1 U14997 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n11871) );
  OR2_X1 U14998 ( .A1(n11897), .A2(n11871), .ZN(n11873) );
  NAND2_X1 U14999 ( .A1(n11897), .A2(BUF2_REG_10__SCAN_IN), .ZN(n11872) );
  NAND2_X1 U15000 ( .A1(n11873), .A2(n11872), .ZN(n14660) );
  NAND2_X1 U15001 ( .A1(n19024), .A2(n14660), .ZN(n11917) );
  NAND2_X1 U15002 ( .A1(n11874), .A2(n11917), .ZN(P2_U2962) );
  AOI22_X1 U15003 ( .A1(n19029), .A2(P2_EAX_REG_28__SCAN_IN), .B1(n11880), 
        .B2(P2_UWORD_REG_12__SCAN_IN), .ZN(n11875) );
  AOI22_X1 U15004 ( .A1(n12980), .A2(BUF1_REG_12__SCAN_IN), .B1(
        BUF2_REG_12__SCAN_IN), .B2(n14634), .ZN(n12263) );
  INV_X1 U15005 ( .A(n12263), .ZN(n14644) );
  NAND2_X1 U15006 ( .A1(n19024), .A2(n14644), .ZN(n11876) );
  NAND2_X1 U15007 ( .A1(n11875), .A2(n11876), .ZN(P2_U2964) );
  AOI22_X1 U15008 ( .A1(n19029), .A2(P2_EAX_REG_12__SCAN_IN), .B1(n11880), 
        .B2(P2_LWORD_REG_12__SCAN_IN), .ZN(n11877) );
  NAND2_X1 U15009 ( .A1(n11877), .A2(n11876), .ZN(P2_U2979) );
  AOI22_X1 U15010 ( .A1(n19029), .A2(P2_EAX_REG_1__SCAN_IN), .B1(n11880), .B2(
        P2_LWORD_REG_1__SCAN_IN), .ZN(n11878) );
  AOI22_X1 U15011 ( .A1(n12980), .A2(BUF1_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n14634), .ZN(n13076) );
  INV_X1 U15012 ( .A(n13076), .ZN(n13294) );
  NAND2_X1 U15013 ( .A1(n19024), .A2(n13294), .ZN(n11913) );
  NAND2_X1 U15014 ( .A1(n11878), .A2(n11913), .ZN(P2_U2968) );
  AOI22_X1 U15015 ( .A1(n19029), .A2(P2_EAX_REG_3__SCAN_IN), .B1(n11880), .B2(
        P2_LWORD_REG_3__SCAN_IN), .ZN(n11879) );
  AOI22_X1 U15016 ( .A1(n12980), .A2(BUF1_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n14634), .ZN(n19073) );
  INV_X1 U15017 ( .A(n19073), .ZN(n14711) );
  NAND2_X1 U15018 ( .A1(n19024), .A2(n14711), .ZN(n11902) );
  NAND2_X1 U15019 ( .A1(n11879), .A2(n11902), .ZN(P2_U2970) );
  AOI22_X1 U15020 ( .A1(n19029), .A2(P2_EAX_REG_0__SCAN_IN), .B1(n11880), .B2(
        P2_LWORD_REG_0__SCAN_IN), .ZN(n11881) );
  AOI22_X1 U15021 ( .A1(n12980), .A2(BUF1_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n14634), .ZN(n12990) );
  INV_X1 U15022 ( .A(n12990), .ZN(n13114) );
  NAND2_X1 U15023 ( .A1(n19024), .A2(n13114), .ZN(n11919) );
  NAND2_X1 U15024 ( .A1(n11881), .A2(n11919), .ZN(P2_U2967) );
  INV_X1 U15025 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n20931) );
  MUX2_X1 U15026 ( .A(BUF1_REG_11__SCAN_IN), .B(BUF2_REG_11__SCAN_IN), .S(
        n14634), .Z(n18941) );
  NAND2_X1 U15027 ( .A1(n19024), .A2(n18941), .ZN(n11890) );
  NAND2_X1 U15028 ( .A1(n19028), .A2(P2_LWORD_REG_11__SCAN_IN), .ZN(n11883) );
  OAI211_X1 U15029 ( .C1(n20931), .C2(n18951), .A(n11890), .B(n11883), .ZN(
        P2_U2978) );
  INV_X1 U15030 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n18970) );
  INV_X1 U15031 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n16326) );
  OR2_X1 U15032 ( .A1(n14634), .A2(n16326), .ZN(n11885) );
  NAND2_X1 U15033 ( .A1(n11897), .A2(BUF2_REG_9__SCAN_IN), .ZN(n11884) );
  NAND2_X1 U15034 ( .A1(n11885), .A2(n11884), .ZN(n18945) );
  NAND2_X1 U15035 ( .A1(n19024), .A2(n18945), .ZN(n11888) );
  NAND2_X1 U15036 ( .A1(n19028), .A2(P2_UWORD_REG_9__SCAN_IN), .ZN(n11886) );
  OAI211_X1 U15037 ( .C1(n18970), .C2(n18951), .A(n11888), .B(n11886), .ZN(
        P2_U2961) );
  INV_X1 U15038 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n19000) );
  NAND2_X1 U15039 ( .A1(n19028), .A2(P2_LWORD_REG_9__SCAN_IN), .ZN(n11887) );
  OAI211_X1 U15040 ( .C1(n19000), .C2(n18951), .A(n11888), .B(n11887), .ZN(
        P2_U2976) );
  INV_X1 U15041 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n18966) );
  NAND2_X1 U15042 ( .A1(n19028), .A2(P2_UWORD_REG_11__SCAN_IN), .ZN(n11889) );
  OAI211_X1 U15043 ( .C1(n18966), .C2(n18951), .A(n11890), .B(n11889), .ZN(
        P2_U2963) );
  AOI22_X1 U15044 ( .A1(n19029), .A2(P2_EAX_REG_21__SCAN_IN), .B1(n19028), 
        .B2(P2_UWORD_REG_5__SCAN_IN), .ZN(n11891) );
  AOI22_X1 U15045 ( .A1(n12980), .A2(BUF1_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n14634), .ZN(n12984) );
  INV_X1 U15046 ( .A(n12984), .ZN(n14692) );
  NAND2_X1 U15047 ( .A1(n19024), .A2(n14692), .ZN(n11892) );
  NAND2_X1 U15048 ( .A1(n11891), .A2(n11892), .ZN(P2_U2957) );
  AOI22_X1 U15049 ( .A1(n19029), .A2(P2_EAX_REG_5__SCAN_IN), .B1(n19028), .B2(
        P2_LWORD_REG_5__SCAN_IN), .ZN(n11893) );
  NAND2_X1 U15050 ( .A1(n11893), .A2(n11892), .ZN(P2_U2972) );
  AOI22_X1 U15051 ( .A1(n19029), .A2(P2_EAX_REG_20__SCAN_IN), .B1(n19028), 
        .B2(P2_UWORD_REG_4__SCAN_IN), .ZN(n11894) );
  AOI22_X1 U15052 ( .A1(n12980), .A2(BUF1_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n14634), .ZN(n19078) );
  INV_X1 U15053 ( .A(n19078), .ZN(n14700) );
  NAND2_X1 U15054 ( .A1(n19024), .A2(n14700), .ZN(n11915) );
  NAND2_X1 U15055 ( .A1(n11894), .A2(n11915), .ZN(P2_U2956) );
  AOI22_X1 U15056 ( .A1(n19029), .A2(P2_EAX_REG_22__SCAN_IN), .B1(n19028), 
        .B2(P2_UWORD_REG_6__SCAN_IN), .ZN(n11895) );
  AOI22_X1 U15057 ( .A1(n12980), .A2(BUF1_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n14634), .ZN(n19088) );
  INV_X1 U15058 ( .A(n19088), .ZN(n14684) );
  NAND2_X1 U15059 ( .A1(n19024), .A2(n14684), .ZN(n11911) );
  NAND2_X1 U15060 ( .A1(n11895), .A2(n11911), .ZN(P2_U2958) );
  AOI22_X1 U15061 ( .A1(n19029), .A2(P2_EAX_REG_8__SCAN_IN), .B1(n19028), .B2(
        P2_LWORD_REG_8__SCAN_IN), .ZN(n11900) );
  INV_X1 U15062 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n11896) );
  OR2_X1 U15063 ( .A1(n11897), .A2(n11896), .ZN(n11899) );
  NAND2_X1 U15064 ( .A1(n14634), .A2(BUF2_REG_8__SCAN_IN), .ZN(n11898) );
  NAND2_X1 U15065 ( .A1(n11899), .A2(n11898), .ZN(n14674) );
  NAND2_X1 U15066 ( .A1(n19024), .A2(n14674), .ZN(n11906) );
  NAND2_X1 U15067 ( .A1(n11900), .A2(n11906), .ZN(P2_U2975) );
  AOI22_X1 U15068 ( .A1(n19029), .A2(P2_EAX_REG_7__SCAN_IN), .B1(n19028), .B2(
        P2_LWORD_REG_7__SCAN_IN), .ZN(n11901) );
  OAI22_X1 U15069 ( .A1(n14634), .A2(BUF1_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n12980), .ZN(n13201) );
  INV_X1 U15070 ( .A(n13201), .ZN(n15926) );
  NAND2_X1 U15071 ( .A1(n19024), .A2(n15926), .ZN(n11904) );
  NAND2_X1 U15072 ( .A1(n11901), .A2(n11904), .ZN(P2_U2974) );
  AOI22_X1 U15073 ( .A1(n19029), .A2(P2_EAX_REG_19__SCAN_IN), .B1(n19028), 
        .B2(P2_UWORD_REG_3__SCAN_IN), .ZN(n11903) );
  NAND2_X1 U15074 ( .A1(n11903), .A2(n11902), .ZN(P2_U2955) );
  AOI22_X1 U15075 ( .A1(n19029), .A2(P2_EAX_REG_23__SCAN_IN), .B1(n19028), 
        .B2(P2_UWORD_REG_7__SCAN_IN), .ZN(n11905) );
  NAND2_X1 U15076 ( .A1(n11905), .A2(n11904), .ZN(P2_U2959) );
  AOI22_X1 U15077 ( .A1(n19029), .A2(P2_EAX_REG_24__SCAN_IN), .B1(n19028), 
        .B2(P2_UWORD_REG_8__SCAN_IN), .ZN(n11907) );
  NAND2_X1 U15078 ( .A1(n11907), .A2(n11906), .ZN(P2_U2960) );
  AOI22_X1 U15079 ( .A1(n19029), .A2(P2_EAX_REG_18__SCAN_IN), .B1(n19028), 
        .B2(P2_UWORD_REG_2__SCAN_IN), .ZN(n11908) );
  AOI22_X1 U15080 ( .A1(n12980), .A2(BUF1_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n14634), .ZN(n19069) );
  INV_X1 U15081 ( .A(n19069), .ZN(n13336) );
  NAND2_X1 U15082 ( .A1(n19024), .A2(n13336), .ZN(n11909) );
  NAND2_X1 U15083 ( .A1(n11908), .A2(n11909), .ZN(P2_U2954) );
  AOI22_X1 U15084 ( .A1(n19029), .A2(P2_EAX_REG_2__SCAN_IN), .B1(n19028), .B2(
        P2_LWORD_REG_2__SCAN_IN), .ZN(n11910) );
  NAND2_X1 U15085 ( .A1(n11910), .A2(n11909), .ZN(P2_U2969) );
  AOI22_X1 U15086 ( .A1(n19029), .A2(P2_EAX_REG_6__SCAN_IN), .B1(n19028), .B2(
        P2_LWORD_REG_6__SCAN_IN), .ZN(n11912) );
  NAND2_X1 U15087 ( .A1(n11912), .A2(n11911), .ZN(P2_U2973) );
  AOI22_X1 U15088 ( .A1(n19029), .A2(P2_EAX_REG_17__SCAN_IN), .B1(n19028), 
        .B2(P2_UWORD_REG_1__SCAN_IN), .ZN(n11914) );
  NAND2_X1 U15089 ( .A1(n11914), .A2(n11913), .ZN(P2_U2953) );
  AOI22_X1 U15090 ( .A1(n19029), .A2(P2_EAX_REG_4__SCAN_IN), .B1(n19028), .B2(
        P2_LWORD_REG_4__SCAN_IN), .ZN(n11916) );
  NAND2_X1 U15091 ( .A1(n11916), .A2(n11915), .ZN(P2_U2971) );
  AOI22_X1 U15092 ( .A1(n19029), .A2(P2_EAX_REG_10__SCAN_IN), .B1(n19028), 
        .B2(P2_LWORD_REG_10__SCAN_IN), .ZN(n11918) );
  NAND2_X1 U15093 ( .A1(n11918), .A2(n11917), .ZN(P2_U2977) );
  AOI22_X1 U15094 ( .A1(n19029), .A2(P2_EAX_REG_16__SCAN_IN), .B1(n19028), 
        .B2(P2_UWORD_REG_0__SCAN_IN), .ZN(n11920) );
  NAND2_X1 U15095 ( .A1(n11920), .A2(n11919), .ZN(P2_U2952) );
  OAI21_X1 U15096 ( .B1(n18915), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n11928), .ZN(n11921) );
  INV_X1 U15097 ( .A(n11921), .ZN(n16152) );
  AND2_X1 U15098 ( .A1(n19033), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n16153) );
  AOI22_X1 U15099 ( .A1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n11923), .B1(
        n11922), .B2(n13195), .ZN(n16155) );
  NOR2_X1 U15100 ( .A1(n19035), .A2(n16155), .ZN(n11924) );
  AOI211_X1 U15101 ( .C1(n16060), .C2(n16152), .A(n16153), .B(n11924), .ZN(
        n11927) );
  OAI21_X1 U15102 ( .B1(n19032), .B2(n11925), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n11926) );
  OAI211_X1 U15103 ( .C1(n12221), .C2(n16058), .A(n11927), .B(n11926), .ZN(
        P2_U3014) );
  XNOR2_X1 U15104 ( .A(n11928), .B(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n11929) );
  XNOR2_X1 U15105 ( .A(n11929), .B(n13173), .ZN(n13897) );
  INV_X1 U15106 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13174) );
  NAND2_X1 U15107 ( .A1(n16054), .A2(n13174), .ZN(n11933) );
  AOI21_X1 U15108 ( .B1(n9972), .B2(n11931), .A(n11930), .ZN(n13895) );
  AND2_X1 U15109 ( .A1(n19033), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n13896) );
  AOI21_X1 U15110 ( .B1(n16055), .B2(n13895), .A(n13896), .ZN(n11932) );
  OAI211_X1 U15111 ( .C1(n16064), .C2(n13174), .A(n11933), .B(n11932), .ZN(
        n11934) );
  AOI21_X1 U15112 ( .B1(n16060), .B2(n13897), .A(n11934), .ZN(n11935) );
  OAI21_X1 U15113 ( .B1(n11154), .B2(n16058), .A(n11935), .ZN(P2_U3013) );
  NOR2_X1 U15114 ( .A1(n11936), .A2(n10907), .ZN(n18950) );
  NAND2_X1 U15115 ( .A1(n18950), .A2(n11937), .ZN(n11945) );
  NAND2_X1 U15116 ( .A1(n11939), .A2(n11938), .ZN(n11940) );
  AND4_X1 U15117 ( .A1(n11943), .A2(n11942), .A3(n11941), .A4(n11940), .ZN(
        n11944) );
  NAND2_X1 U15118 ( .A1(n11945), .A2(n11944), .ZN(n16180) );
  NAND2_X1 U15119 ( .A1(n16180), .A2(n18949), .ZN(n11949) );
  INV_X1 U15120 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n18954) );
  INV_X1 U15121 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n13196) );
  NOR2_X1 U15122 ( .A1(n19744), .A2(n13196), .ZN(n19719) );
  AND2_X1 U15123 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19719), .ZN(n16196) );
  AOI21_X1 U15124 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n18954), .A(n16196), 
        .ZN(n16206) );
  AOI21_X1 U15125 ( .B1(n11946), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n16206), 
        .ZN(n11947) );
  INV_X1 U15126 ( .A(n11947), .ZN(n11948) );
  NAND2_X1 U15127 ( .A1(n11949), .A2(n11948), .ZN(n15106) );
  INV_X1 U15128 ( .A(n15106), .ZN(n13199) );
  INV_X1 U15129 ( .A(n19606), .ZN(n19687) );
  INV_X1 U15130 ( .A(n10907), .ZN(n11951) );
  NAND3_X1 U15131 ( .A1(n11951), .A2(n11164), .A3(n11950), .ZN(n16174) );
  OR3_X1 U15132 ( .A1(n13199), .A2(n19687), .A3(n16174), .ZN(n11952) );
  OAI21_X1 U15133 ( .B1(n16179), .B2(n15106), .A(n11952), .ZN(P2_U3595) );
  OAI21_X1 U15134 ( .B1(n11955), .B2(n11954), .A(n11953), .ZN(n11956) );
  INV_X1 U15135 ( .A(n11956), .ZN(n19064) );
  OAI21_X1 U15136 ( .B1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A(n11957), .ZN(n13034) );
  NOR2_X1 U15137 ( .A1(n18846), .A2(n11958), .ZN(n19058) );
  OAI21_X1 U15138 ( .B1(n9822), .B2(n11960), .A(n11959), .ZN(n19055) );
  NOR2_X1 U15139 ( .A1(n19055), .A2(n19035), .ZN(n11961) );
  AOI211_X1 U15140 ( .C1(n19032), .C2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A(
        n19058), .B(n11961), .ZN(n11962) );
  OAI21_X1 U15141 ( .B1(n19045), .B2(n13034), .A(n11962), .ZN(n11963) );
  AOI21_X1 U15142 ( .B1(n16060), .B2(n19064), .A(n11963), .ZN(n11964) );
  OAI21_X1 U15143 ( .B1(n11148), .B2(n16058), .A(n11964), .ZN(P2_U3012) );
  OR2_X1 U15144 ( .A1(n11966), .A2(n11965), .ZN(n12888) );
  OR2_X1 U15145 ( .A1(n11968), .A2(n11967), .ZN(n11969) );
  NAND2_X1 U15146 ( .A1(n11970), .A2(n11969), .ZN(n18881) );
  INV_X1 U15147 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n19005) );
  OAI222_X1 U15148 ( .A1(n12888), .A2(n19088), .B1(n18881), .B2(n18937), .C1(
        n18948), .C2(n19005), .ZN(P2_U2913) );
  NAND2_X1 U15149 ( .A1(n10944), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n11971) );
  AND4_X1 U15150 ( .A1(n11971), .A2(n19085), .A3(P2_STATE2_REG_0__SCAN_IN), 
        .A4(n19714), .ZN(n11972) );
  OR2_X1 U15151 ( .A1(n11974), .A2(n11973), .ZN(n11975) );
  NAND2_X1 U15152 ( .A1(n10966), .A2(n11975), .ZN(n11976) );
  INV_X1 U15153 ( .A(n11976), .ZN(n18916) );
  NOR2_X1 U15154 ( .A1(n19716), .A2(n11976), .ZN(n12208) );
  INV_X1 U15155 ( .A(n12208), .ZN(n11977) );
  OAI211_X1 U15156 ( .C1(n18912), .C2(n18916), .A(n11977), .B(n15928), .ZN(
        n11979) );
  AOI22_X1 U15157 ( .A1(n18930), .A2(n18916), .B1(n18934), .B2(
        P2_EAX_REG_0__SCAN_IN), .ZN(n11978) );
  OAI211_X1 U15158 ( .C1(n12990), .C2(n12888), .A(n11979), .B(n11978), .ZN(
        P2_U2919) );
  INV_X1 U15159 ( .A(n14674), .ZN(n11982) );
  OR2_X1 U15160 ( .A1(n11980), .A2(n11989), .ZN(n11981) );
  NAND2_X1 U15161 ( .A1(n11981), .A2(n15031), .ZN(n18857) );
  INV_X1 U15162 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n19002) );
  OAI222_X1 U15163 ( .A1(n12888), .A2(n11982), .B1(n18857), .B2(n18937), .C1(
        n18948), .C2(n19002), .ZN(P2_U2911) );
  MUX2_X1 U15164 ( .A(P2_EBX_REG_2__SCAN_IN), .B(n11986), .S(n14621), .Z(
        n11987) );
  AOI21_X1 U15165 ( .B1(n13215), .B2(n14601), .A(n11987), .ZN(n11988) );
  INV_X1 U15166 ( .A(n11988), .ZN(P2_U2885) );
  INV_X1 U15167 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n11992) );
  AOI21_X1 U15168 ( .B1(n11991), .B2(n11990), .A(n11989), .ZN(n18867) );
  INV_X1 U15169 ( .A(n18867), .ZN(n15068) );
  OAI222_X1 U15170 ( .A1(n11992), .A2(n18948), .B1(n12888), .B2(n13201), .C1(
        n15068), .C2(n18937), .ZN(P2_U2912) );
  MUX2_X1 U15171 ( .A(n20757), .B(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .S(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Z(n12000) );
  NOR2_X1 U15172 ( .A1(n12553), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n11993) );
  INV_X1 U15173 ( .A(n12002), .ZN(n11996) );
  XNOR2_X1 U15174 ( .A(n9900), .B(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n12001) );
  INV_X1 U15175 ( .A(n12001), .ZN(n11995) );
  INV_X1 U15176 ( .A(n12005), .ZN(n11997) );
  XNOR2_X1 U15177 ( .A(n12778), .B(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n12006) );
  INV_X1 U15178 ( .A(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n20003) );
  NOR2_X1 U15179 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n20003), .ZN(
        n11999) );
  AOI221_X1 U15180 ( .B1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(n12007), 
        .C1(n15813), .C2(n12007), .A(n11999), .ZN(n12144) );
  XNOR2_X1 U15181 ( .A(n12000), .B(n12147), .ZN(n12159) );
  NAND2_X1 U15182 ( .A1(n12002), .A2(n12001), .ZN(n12004) );
  NAND2_X1 U15183 ( .A1(n12004), .A2(n12003), .ZN(n12160) );
  XNOR2_X1 U15184 ( .A(n12006), .B(n12005), .ZN(n12145) );
  NAND3_X1 U15185 ( .A1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n12007), .A3(
        n15813), .ZN(n12170) );
  NAND2_X1 U15186 ( .A1(n12145), .A2(n12170), .ZN(n12167) );
  NOR2_X1 U15187 ( .A1(n12160), .A2(n12167), .ZN(n12008) );
  AND2_X1 U15188 ( .A1(n12159), .A2(n12008), .ZN(n12009) );
  OR2_X1 U15189 ( .A1(n12144), .A2(n12009), .ZN(n13412) );
  AND2_X4 U15190 ( .A1(n12782), .A2(n14515), .ZN(n13867) );
  AOI22_X1 U15191 ( .A1(n13477), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n13867), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12013) );
  AND2_X2 U15192 ( .A1(n12782), .A2(n12014), .ZN(n12374) );
  AOI22_X1 U15193 ( .A1(n12374), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n9755), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12012) );
  AOI22_X1 U15194 ( .A1(n13843), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12067), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12011) );
  AND2_X2 U15195 ( .A1(n12781), .A2(n12014), .ZN(n12126) );
  AOI22_X1 U15196 ( .A1(n12126), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n13718), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12010) );
  NAND4_X1 U15197 ( .A1(n12013), .A2(n12012), .A3(n12011), .A4(n12010), .ZN(
        n12020) );
  AOI22_X1 U15198 ( .A1(n12709), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n13869), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12018) );
  AOI22_X1 U15199 ( .A1(n9738), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12658), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12017) );
  AND2_X4 U15200 ( .A1(n14516), .A2(n12784), .ZN(n13825) );
  AOI22_X1 U15201 ( .A1(n13862), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n13825), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12016) );
  AND2_X4 U15202 ( .A1(n12014), .A2(n12784), .ZN(n13848) );
  AOI22_X1 U15203 ( .A1(n13848), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12082), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12015) );
  NAND4_X1 U15204 ( .A1(n12018), .A2(n12017), .A3(n12016), .A4(n12015), .ZN(
        n12019) );
  AOI22_X1 U15205 ( .A1(n13477), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n13867), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12024) );
  AOI22_X1 U15206 ( .A1(n12709), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n13869), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12023) );
  AOI22_X1 U15207 ( .A1(n13848), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12067), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12022) );
  AOI22_X1 U15208 ( .A1(n12658), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n13718), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12021) );
  NAND4_X1 U15209 ( .A1(n12024), .A2(n12023), .A3(n12022), .A4(n12021), .ZN(
        n12030) );
  AOI22_X1 U15210 ( .A1(n9740), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12126), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12028) );
  AOI22_X1 U15211 ( .A1(n12374), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n9756), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12027) );
  AOI22_X1 U15212 ( .A1(n13862), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n13825), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12026) );
  AOI22_X1 U15213 ( .A1(n13843), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12082), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12025) );
  NAND4_X1 U15214 ( .A1(n12028), .A2(n12027), .A3(n12026), .A4(n12025), .ZN(
        n12029) );
  AOI22_X1 U15215 ( .A1(n12709), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n13869), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12034) );
  AOI22_X1 U15216 ( .A1(n9741), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12126), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12033) );
  AOI22_X1 U15217 ( .A1(n12374), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n9755), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12032) );
  AOI22_X1 U15218 ( .A1(n13862), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n13825), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12031) );
  AOI22_X1 U15219 ( .A1(n13843), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n13867), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12038) );
  AOI22_X1 U15220 ( .A1(n12658), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n13718), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12037) );
  AOI22_X1 U15221 ( .A1(n13848), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n9721), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12036) );
  NAND2_X1 U15222 ( .A1(n12341), .A2(n12469), .ZN(n12358) );
  NAND2_X1 U15223 ( .A1(n12709), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n12042) );
  NAND2_X1 U15224 ( .A1(n9740), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n12041) );
  NAND2_X1 U15225 ( .A1(n13862), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n12040) );
  NAND2_X1 U15226 ( .A1(n12126), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n12039) );
  NAND2_X1 U15227 ( .A1(n13477), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n12046) );
  NAND2_X1 U15228 ( .A1(n13843), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n12045) );
  NAND2_X1 U15229 ( .A1(n13867), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n12044) );
  NAND2_X1 U15230 ( .A1(n12082), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n12043) );
  NAND2_X1 U15231 ( .A1(n13869), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n12050) );
  NAND2_X1 U15232 ( .A1(n12374), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n12049) );
  NAND2_X1 U15233 ( .A1(n9757), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n12048) );
  NAND2_X1 U15234 ( .A1(n13825), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n12047) );
  NAND2_X1 U15235 ( .A1(n12658), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n12054) );
  NAND2_X1 U15236 ( .A1(n13848), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n12053) );
  NAND2_X1 U15237 ( .A1(n12067), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n12052) );
  NAND2_X1 U15238 ( .A1(n13718), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n12051) );
  NAND2_X1 U15239 ( .A1(n13862), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n12062) );
  NAND2_X1 U15240 ( .A1(n12709), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n12061) );
  NAND2_X1 U15241 ( .A1(n13869), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n12060) );
  NAND2_X1 U15242 ( .A1(n13825), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n12059) );
  NAND2_X1 U15243 ( .A1(n12374), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n12066) );
  NAND2_X1 U15244 ( .A1(n9741), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n12065) );
  NAND2_X1 U15245 ( .A1(n12126), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n12064) );
  NAND2_X1 U15246 ( .A1(n9757), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n12063) );
  NAND2_X1 U15247 ( .A1(n13477), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n12075) );
  NAND2_X1 U15248 ( .A1(n12658), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n12074) );
  NAND2_X1 U15249 ( .A1(n13718), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n12073) );
  NAND2_X1 U15250 ( .A1(n12082), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n12072) );
  NAND2_X1 U15251 ( .A1(n12539), .A2(n12119), .ZN(n12080) );
  NAND2_X1 U15252 ( .A1(n13891), .A2(n12080), .ZN(n12081) );
  NAND2_X1 U15253 ( .A1(n12358), .A2(n12081), .ZN(n12095) );
  NAND2_X2 U15254 ( .A1(n12187), .A2(n12121), .ZN(n12096) );
  AOI22_X1 U15255 ( .A1(n13848), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12067), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12086) );
  AOI22_X1 U15256 ( .A1(n13477), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n12082), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12085) );
  AOI22_X1 U15257 ( .A1(n13862), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n13825), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12084) );
  AOI22_X1 U15258 ( .A1(n9755), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n12658), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12083) );
  NAND3_X1 U15259 ( .A1(n12086), .A2(n12085), .A3(n10278), .ZN(n12092) );
  AOI22_X1 U15260 ( .A1(n12374), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12126), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12090) );
  AOI22_X1 U15261 ( .A1(n13843), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n13867), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12089) );
  AOI22_X1 U15262 ( .A1(n12709), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n13869), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12088) );
  AOI22_X1 U15263 ( .A1(n9739), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n13718), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12087) );
  NAND4_X1 U15264 ( .A1(n12090), .A2(n12089), .A3(n12088), .A4(n12087), .ZN(
        n12091) );
  NAND2_X1 U15265 ( .A1(n13862), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n12100) );
  NAND2_X1 U15266 ( .A1(n12709), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n12099) );
  NAND2_X1 U15267 ( .A1(n9756), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n12098) );
  NAND2_X1 U15268 ( .A1(n13825), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n12097) );
  NAND2_X1 U15269 ( .A1(n13867), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n12104) );
  NAND2_X1 U15270 ( .A1(n13477), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n12103) );
  NAND2_X1 U15271 ( .A1(n13843), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n12102) );
  NAND2_X1 U15272 ( .A1(n12067), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n12101) );
  NAND2_X1 U15273 ( .A1(n12658), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n12108) );
  NAND2_X1 U15274 ( .A1(n12374), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n12107) );
  NAND2_X1 U15275 ( .A1(n13848), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n12106) );
  NAND2_X1 U15276 ( .A1(n13718), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n12105) );
  NAND2_X1 U15277 ( .A1(n9739), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n12112) );
  NAND2_X1 U15278 ( .A1(n12126), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n12111) );
  NAND2_X1 U15279 ( .A1(n12082), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n12109) );
  NOR2_X1 U15280 ( .A1(n12096), .A2(n9725), .ZN(n12117) );
  INV_X1 U15281 ( .A(n12347), .ZN(n12568) );
  NOR2_X1 U15282 ( .A1(n13412), .A2(n12568), .ZN(n12224) );
  INV_X1 U15283 ( .A(n12340), .ZN(n15453) );
  OR2_X1 U15284 ( .A1(n12224), .A2(n15453), .ZN(n12179) );
  NAND2_X1 U15285 ( .A1(n13862), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n12125) );
  NAND2_X1 U15286 ( .A1(n12709), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n12124) );
  NAND2_X1 U15287 ( .A1(n13869), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n12123) );
  NAND2_X1 U15288 ( .A1(n13825), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n12122) );
  NAND2_X1 U15289 ( .A1(n12374), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n12131) );
  NAND2_X1 U15290 ( .A1(n9738), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n12130) );
  NAND2_X1 U15291 ( .A1(n12126), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n12129) );
  NAND2_X1 U15292 ( .A1(n9756), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n12128) );
  NAND2_X1 U15293 ( .A1(n13843), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n12135) );
  NAND2_X1 U15294 ( .A1(n13867), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n12134) );
  NAND2_X1 U15295 ( .A1(n13848), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n12133) );
  NAND2_X1 U15296 ( .A1(n12067), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n12132) );
  NAND2_X1 U15297 ( .A1(n13477), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n12139) );
  NAND2_X1 U15298 ( .A1(n12658), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n12138) );
  NAND2_X1 U15299 ( .A1(n13718), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n12137) );
  NAND2_X1 U15300 ( .A1(n12082), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n12136) );
  NAND4_X4 U15301 ( .A1(n12143), .A2(n12142), .A3(n12141), .A4(n12140), .ZN(
        n13438) );
  NAND2_X1 U15302 ( .A1(n12144), .A2(n12173), .ZN(n12177) );
  NAND2_X1 U15303 ( .A1(n12144), .A2(n13086), .ZN(n12176) );
  INV_X1 U15304 ( .A(n12145), .ZN(n12172) );
  INV_X1 U15305 ( .A(n12148), .ZN(n12165) );
  OAI21_X1 U15306 ( .B1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n20435), .A(
        n12147), .ZN(n12150) );
  NOR2_X1 U15307 ( .A1(n12150), .A2(n12149), .ZN(n12153) );
  INV_X1 U15308 ( .A(n12150), .ZN(n12151) );
  AOI21_X1 U15309 ( .B1(n12151), .B2(n13086), .A(n12173), .ZN(n12152) );
  NOR2_X1 U15310 ( .A1(n12153), .A2(n12152), .ZN(n12158) );
  NAND2_X1 U15311 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n20038), .ZN(n12155) );
  NAND2_X1 U15312 ( .A1(n13086), .A2(n13438), .ZN(n12154) );
  OAI211_X1 U15313 ( .C1(n12159), .C2(n13089), .A(n12155), .B(n12154), .ZN(
        n12157) );
  NAND2_X1 U15314 ( .A1(n12158), .A2(n12157), .ZN(n12163) );
  INV_X1 U15315 ( .A(n12155), .ZN(n12156) );
  OAI22_X1 U15316 ( .A1(n12168), .A2(n12159), .B1(n12158), .B2(n12157), .ZN(
        n12162) );
  AOI211_X1 U15317 ( .C1(n12665), .C2(n12160), .A(n12166), .B(n12165), .ZN(
        n12161) );
  AOI21_X1 U15318 ( .B1(n12163), .B2(n12162), .A(n12161), .ZN(n12164) );
  INV_X1 U15319 ( .A(n12168), .ZN(n12169) );
  NAND2_X1 U15320 ( .A1(n15462), .A2(n9906), .ZN(n12178) );
  NAND2_X1 U15321 ( .A1(n12179), .A2(n12178), .ZN(n19758) );
  XNOR2_X1 U15322 ( .A(P1_STATE_REG_1__SCAN_IN), .B(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n12339) );
  INV_X1 U15323 ( .A(n12339), .ZN(n12181) );
  INV_X1 U15324 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n20585) );
  NAND2_X1 U15325 ( .A1(n12181), .A2(n20585), .ZN(n15490) );
  NAND3_X1 U15326 ( .A1(n9906), .A2(n13950), .A3(n15490), .ZN(n12182) );
  NAND2_X1 U15327 ( .A1(READY1), .A2(READY11_REG_SCAN_IN), .ZN(n20666) );
  AND2_X1 U15328 ( .A1(n12182), .A2(n20666), .ZN(n20668) );
  NOR2_X1 U15329 ( .A1(n19758), .A2(n20668), .ZN(n15444) );
  NAND2_X1 U15330 ( .A1(n20898), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20578) );
  OR2_X1 U15331 ( .A1(n15444), .A2(n19757), .ZN(n12198) );
  INV_X1 U15332 ( .A(n12198), .ZN(n19766) );
  INV_X1 U15333 ( .A(P1_MORE_REG_SCAN_IN), .ZN(n12200) );
  OR2_X1 U15334 ( .A1(n12469), .A2(n20010), .ZN(n12330) );
  NAND2_X2 U15335 ( .A1(n12330), .A2(n13936), .ZN(n13951) );
  INV_X1 U15336 ( .A(n12342), .ZN(n12184) );
  NAND2_X1 U15337 ( .A1(n20010), .A2(n13438), .ZN(n12565) );
  INV_X1 U15338 ( .A(n12565), .ZN(n12846) );
  NAND2_X1 U15339 ( .A1(n12846), .A2(n12096), .ZN(n12183) );
  NAND2_X1 U15340 ( .A1(n12184), .A2(n12183), .ZN(n12538) );
  NAND3_X1 U15341 ( .A1(n13437), .A2(n13438), .A3(n12539), .ZN(n12185) );
  NOR2_X1 U15342 ( .A1(n12341), .A2(n12185), .ZN(n12333) );
  INV_X1 U15343 ( .A(n12333), .ZN(n12186) );
  NOR2_X1 U15344 ( .A1(n12538), .A2(n12186), .ZN(n13433) );
  INV_X1 U15345 ( .A(n13433), .ZN(n12196) );
  AND2_X1 U15346 ( .A1(n12334), .A2(n12539), .ZN(n12350) );
  NAND2_X1 U15347 ( .A1(n12188), .A2(n20034), .ZN(n12189) );
  AOI21_X1 U15348 ( .B1(n20010), .B2(n12341), .A(n12909), .ZN(n12190) );
  INV_X1 U15349 ( .A(n12096), .ZN(n12474) );
  OR2_X1 U15350 ( .A1(n12844), .A2(n12474), .ZN(n12192) );
  NAND2_X1 U15351 ( .A1(n12566), .A2(n12192), .ZN(n13423) );
  OAI21_X1 U15352 ( .B1(n20010), .B2(n12193), .A(n13423), .ZN(n12194) );
  AOI22_X1 U15353 ( .A1(n15462), .A2(n12194), .B1(n12347), .B2(n13412), .ZN(
        n12195) );
  OAI21_X1 U15354 ( .B1(n15462), .B2(n12196), .A(n12195), .ZN(n12197) );
  NAND2_X1 U15355 ( .A1(n12197), .A2(n12539), .ZN(n15445) );
  OR2_X1 U15356 ( .A1(n12198), .A2(n15445), .ZN(n12199) );
  OAI21_X1 U15357 ( .B1(n19766), .B2(n12200), .A(n12199), .ZN(P1_U3484) );
  INV_X1 U15358 ( .A(n12201), .ZN(n12203) );
  XNOR2_X1 U15359 ( .A(n12205), .B(n12204), .ZN(n19712) );
  INV_X1 U15360 ( .A(n19712), .ZN(n12206) );
  NAND2_X1 U15361 ( .A1(n19707), .A2(n12206), .ZN(n12248) );
  OAI21_X1 U15362 ( .B1(n19707), .B2(n12206), .A(n12248), .ZN(n12207) );
  NOR2_X1 U15363 ( .A1(n12207), .A2(n12208), .ZN(n12250) );
  AOI21_X1 U15364 ( .B1(n12208), .B2(n12207), .A(n12250), .ZN(n12211) );
  INV_X1 U15365 ( .A(n15928), .ZN(n14714) );
  AOI22_X1 U15366 ( .A1(n18930), .A2(n19712), .B1(n18934), .B2(
        P2_EAX_REG_1__SCAN_IN), .ZN(n12210) );
  INV_X1 U15367 ( .A(n12888), .ZN(n18946) );
  NAND2_X1 U15368 ( .A1(n18946), .A2(n13294), .ZN(n12209) );
  OAI211_X1 U15369 ( .C1(n12211), .C2(n14714), .A(n12210), .B(n12209), .ZN(
        P2_U2918) );
  MUX2_X1 U15370 ( .A(n12212), .B(n11154), .S(n14582), .Z(n12213) );
  OAI21_X1 U15371 ( .B1(n19707), .B2(n14630), .A(n12213), .ZN(P2_U2886) );
  NOR2_X1 U15372 ( .A1(n11119), .A2(n14602), .ZN(n12218) );
  AOI21_X1 U15373 ( .B1(P2_EBX_REG_3__SCAN_IN), .B2(n14602), .A(n12218), .ZN(
        n12219) );
  OAI21_X1 U15374 ( .B1(n15105), .B2(n14630), .A(n12219), .ZN(P2_U2884) );
  MUX2_X1 U15375 ( .A(n12221), .B(n12220), .S(n14602), .Z(n12222) );
  OAI21_X1 U15376 ( .B1(n19716), .B2(n14630), .A(n12222), .ZN(P2_U2887) );
  NOR2_X2 U15377 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20524) );
  NAND2_X1 U15378 ( .A1(n20524), .A2(n20898), .ZN(n19760) );
  INV_X1 U15379 ( .A(n19760), .ZN(n12223) );
  NOR2_X1 U15380 ( .A1(n12223), .A2(P1_READREQUEST_REG_SCAN_IN), .ZN(n12226)
         );
  NAND2_X1 U15381 ( .A1(n12224), .A2(n13421), .ZN(n13903) );
  OAI21_X1 U15382 ( .B1(n12844), .B2(n13971), .A(n20664), .ZN(n12225) );
  OAI21_X1 U15383 ( .B1(n12226), .B2(n20664), .A(n12225), .ZN(P1_U3487) );
  INV_X1 U15384 ( .A(n14660), .ZN(n12229) );
  OR2_X1 U15385 ( .A1(n12227), .A2(n15033), .ZN(n12228) );
  NAND2_X1 U15386 ( .A1(n12228), .A2(n16117), .ZN(n18833) );
  INV_X1 U15387 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n18998) );
  OAI222_X1 U15388 ( .A1(n12888), .A2(n12229), .B1(n18833), .B2(n18937), .C1(
        n18948), .C2(n18998), .ZN(P2_U2909) );
  NAND2_X1 U15389 ( .A1(n12230), .A2(n12280), .ZN(n12272) );
  INV_X1 U15390 ( .A(n12231), .ZN(n12232) );
  OR3_X1 U15391 ( .A1(n12233), .A2(n12232), .A3(n12280), .ZN(n12234) );
  NAND2_X1 U15392 ( .A1(n12272), .A2(n12234), .ZN(n12578) );
  INV_X1 U15393 ( .A(n12235), .ZN(n12266) );
  AOI21_X1 U15394 ( .B1(n12237), .B2(n12236), .A(n12266), .ZN(n19040) );
  INV_X1 U15395 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n12238) );
  NOR2_X1 U15396 ( .A1(n14582), .A2(n12238), .ZN(n12239) );
  AOI21_X1 U15397 ( .B1(n19040), .B2(n14621), .A(n12239), .ZN(n12240) );
  OAI21_X1 U15398 ( .B1(n12578), .B2(n14630), .A(n12240), .ZN(P2_U2883) );
  NAND2_X1 U15399 ( .A1(n12230), .A2(n12241), .ZN(n12283) );
  XNOR2_X1 U15400 ( .A(n12283), .B(n12242), .ZN(n12247) );
  NAND2_X1 U15401 ( .A1(n12287), .A2(n12243), .ZN(n12244) );
  NAND2_X1 U15402 ( .A1(n12303), .A2(n12244), .ZN(n18844) );
  MUX2_X1 U15403 ( .A(n18844), .B(n12245), .S(n14602), .Z(n12246) );
  OAI21_X1 U15404 ( .B1(n12247), .B2(n14630), .A(n12246), .ZN(P2_U2878) );
  INV_X1 U15405 ( .A(n12248), .ZN(n12249) );
  NOR2_X1 U15406 ( .A1(n12250), .A2(n12249), .ZN(n12257) );
  INV_X1 U15407 ( .A(n13215), .ZN(n19700) );
  OR2_X1 U15408 ( .A1(n12252), .A2(n12251), .ZN(n12254) );
  NAND2_X1 U15409 ( .A1(n12254), .A2(n12253), .ZN(n19702) );
  INV_X1 U15410 ( .A(n19702), .ZN(n12255) );
  NAND2_X1 U15411 ( .A1(n19700), .A2(n12255), .ZN(n12457) );
  OAI21_X1 U15412 ( .B1(n19700), .B2(n12255), .A(n12457), .ZN(n12256) );
  NOR2_X1 U15413 ( .A1(n12257), .A2(n12256), .ZN(n12459) );
  AOI21_X1 U15414 ( .B1(n12257), .B2(n12256), .A(n12459), .ZN(n12260) );
  AOI22_X1 U15415 ( .A1(n18930), .A2(n19702), .B1(n18934), .B2(
        P2_EAX_REG_2__SCAN_IN), .ZN(n12259) );
  NAND2_X1 U15416 ( .A1(n18946), .A2(n13336), .ZN(n12258) );
  OAI211_X1 U15417 ( .C1(n12260), .C2(n14714), .A(n12259), .B(n12258), .ZN(
        P2_U2917) );
  OR2_X1 U15418 ( .A1(n12261), .A2(n16116), .ZN(n12262) );
  NAND2_X1 U15419 ( .A1(n12262), .A2(n16098), .ZN(n18808) );
  INV_X1 U15420 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n18995) );
  OAI222_X1 U15421 ( .A1(n12888), .A2(n12263), .B1(n18808), .B2(n18937), .C1(
        n18948), .C2(n18995), .ZN(P2_U2907) );
  XOR2_X1 U15422 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B(n12272), .Z(n12269)
         );
  INV_X1 U15423 ( .A(n12264), .ZN(n12265) );
  OAI21_X1 U15424 ( .B1(n12266), .B2(n12265), .A(n12275), .ZN(n18893) );
  NOR2_X1 U15425 ( .A1(n18893), .A2(n14602), .ZN(n12267) );
  AOI21_X1 U15426 ( .B1(P2_EBX_REG_5__SCAN_IN), .B2(n14602), .A(n12267), .ZN(
        n12268) );
  OAI21_X1 U15427 ( .B1(n12269), .B2(n14630), .A(n12268), .ZN(P2_U2882) );
  NOR2_X1 U15428 ( .A1(n12272), .A2(n12270), .ZN(n12273) );
  OR2_X1 U15429 ( .A1(n12272), .A2(n12271), .ZN(n12292) );
  OAI211_X1 U15430 ( .C1(n12273), .C2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A(
        n14601), .B(n12292), .ZN(n12278) );
  INV_X1 U15431 ( .A(n12294), .ZN(n12274) );
  AOI21_X1 U15432 ( .B1(n12276), .B2(n12275), .A(n12274), .ZN(n18877) );
  NAND2_X1 U15433 ( .A1(n18877), .A2(n14582), .ZN(n12277) );
  OAI211_X1 U15434 ( .C1(n14621), .C2(n12279), .A(n12278), .B(n12277), .ZN(
        P2_U2881) );
  AND2_X1 U15435 ( .A1(n12230), .A2(n12280), .ZN(n12282) );
  AND2_X1 U15436 ( .A1(n12282), .A2(n12281), .ZN(n12285) );
  OAI211_X1 U15437 ( .C1(n12285), .C2(n12284), .A(n12283), .B(n14601), .ZN(
        n12290) );
  OR2_X1 U15438 ( .A1(n12293), .A2(n12286), .ZN(n12288) );
  AND2_X1 U15439 ( .A1(n12288), .A2(n12287), .ZN(n18853) );
  NAND2_X1 U15440 ( .A1(n18853), .A2(n14582), .ZN(n12289) );
  OAI211_X1 U15441 ( .C1(n14621), .C2(n12291), .A(n12290), .B(n12289), .ZN(
        P2_U2879) );
  XOR2_X1 U15442 ( .A(n12292), .B(P2_INSTQUEUE_REG_0__7__SCAN_IN), .Z(n12297)
         );
  AOI21_X1 U15443 ( .B1(n12295), .B2(n12294), .A(n12293), .ZN(n16035) );
  INV_X1 U15444 ( .A(n16035), .ZN(n18870) );
  MUX2_X1 U15445 ( .A(n11306), .B(n18870), .S(n14582), .Z(n12296) );
  OAI21_X1 U15446 ( .B1(n12297), .B2(n14630), .A(n12296), .ZN(P2_U2880) );
  INV_X1 U15447 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n12307) );
  AND2_X1 U15448 ( .A1(n12230), .A2(n12298), .ZN(n12302) );
  AND2_X1 U15449 ( .A1(n12230), .A2(n12299), .ZN(n12519) );
  INV_X1 U15450 ( .A(n12519), .ZN(n12300) );
  OAI211_X1 U15451 ( .C1(n12302), .C2(n12301), .A(n12300), .B(n14601), .ZN(
        n12306) );
  AOI21_X1 U15452 ( .B1(n12304), .B2(n12303), .A(n12496), .ZN(n18830) );
  NAND2_X1 U15453 ( .A1(n18830), .A2(n14582), .ZN(n12305) );
  OAI211_X1 U15454 ( .C1(n14621), .C2(n12307), .A(n12306), .B(n12305), .ZN(
        P2_U2877) );
  INV_X1 U15455 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n12313) );
  NOR2_X1 U15456 ( .A1(n12565), .A2(n12096), .ZN(n12308) );
  AND2_X1 U15457 ( .A1(n12345), .A2(n12308), .ZN(n13426) );
  INV_X1 U15458 ( .A(n13426), .ZN(n12790) );
  OAI21_X1 U15459 ( .B1(n13904), .B2(n13438), .A(n12309), .ZN(n12311) );
  INV_X1 U15460 ( .A(n15490), .ZN(n12310) );
  NOR2_X1 U15461 ( .A1(n20898), .A2(n12396), .ZN(n15818) );
  OR2_X1 U15462 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n15824), .ZN(n19887) );
  INV_X2 U15463 ( .A(n19887), .ZN(n20667) );
  AOI22_X1 U15464 ( .A1(P1_UWORD_REG_3__SCAN_IN), .A2(n20667), .B1(n15492), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n12312) );
  OAI21_X1 U15465 ( .B1(n12313), .B2(n12616), .A(n12312), .ZN(P1_U2917) );
  INV_X1 U15466 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n12315) );
  AOI22_X1 U15467 ( .A1(P1_UWORD_REG_1__SCAN_IN), .A2(n20667), .B1(n15492), 
        .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n12314) );
  OAI21_X1 U15468 ( .B1(n12315), .B2(n12616), .A(n12314), .ZN(P1_U2919) );
  INV_X1 U15469 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n12317) );
  AOI22_X1 U15470 ( .A1(P1_UWORD_REG_9__SCAN_IN), .A2(n20667), .B1(n15492), 
        .B2(P1_DATAO_REG_25__SCAN_IN), .ZN(n12316) );
  OAI21_X1 U15471 ( .B1(n12317), .B2(n12616), .A(n12316), .ZN(P1_U2911) );
  INV_X1 U15472 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n12319) );
  AOI22_X1 U15473 ( .A1(P1_UWORD_REG_8__SCAN_IN), .A2(n20667), .B1(n15492), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n12318) );
  OAI21_X1 U15474 ( .B1(n12319), .B2(n12616), .A(n12318), .ZN(P1_U2912) );
  INV_X1 U15475 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n20934) );
  AOI22_X1 U15476 ( .A1(P1_UWORD_REG_2__SCAN_IN), .A2(n20667), .B1(n15492), 
        .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n12320) );
  OAI21_X1 U15477 ( .B1(n20934), .B2(n12616), .A(n12320), .ZN(P1_U2918) );
  INV_X1 U15478 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n12322) );
  AOI22_X1 U15479 ( .A1(P1_UWORD_REG_12__SCAN_IN), .A2(n20667), .B1(n15492), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n12321) );
  OAI21_X1 U15480 ( .B1(n12322), .B2(n12616), .A(n12321), .ZN(P1_U2908) );
  INV_X1 U15481 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n12324) );
  AOI22_X1 U15482 ( .A1(P1_UWORD_REG_0__SCAN_IN), .A2(n20667), .B1(n15492), 
        .B2(P1_DATAO_REG_16__SCAN_IN), .ZN(n12323) );
  OAI21_X1 U15483 ( .B1(n12324), .B2(n12616), .A(n12323), .ZN(P1_U2920) );
  INV_X1 U15484 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n12326) );
  AOI22_X1 U15485 ( .A1(P1_UWORD_REG_13__SCAN_IN), .A2(n20667), .B1(n15492), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n12325) );
  OAI21_X1 U15486 ( .B1(n12326), .B2(n12616), .A(n12325), .ZN(P1_U2907) );
  INV_X1 U15487 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n20835) );
  AOI22_X1 U15488 ( .A1(P1_UWORD_REG_7__SCAN_IN), .A2(n20667), .B1(n15492), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n12327) );
  OAI21_X1 U15489 ( .B1(n20835), .B2(n12616), .A(n12327), .ZN(P1_U2913) );
  INV_X1 U15490 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n12329) );
  AOI22_X1 U15491 ( .A1(P1_UWORD_REG_11__SCAN_IN), .A2(n20667), .B1(n15492), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n12328) );
  OAI21_X1 U15492 ( .B1(n12329), .B2(n12616), .A(n12328), .ZN(P1_U2909) );
  NOR2_X1 U15493 ( .A1(n13951), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12332) );
  INV_X1 U15494 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n12331) );
  OAI22_X1 U15495 ( .A1(n13944), .A2(n12331), .B1(n9724), .B2(
        P1_EBX_REG_0__SCAN_IN), .ZN(n12455) );
  OR2_X1 U15496 ( .A1(n12332), .A2(n12455), .ZN(n12849) );
  NAND2_X1 U15497 ( .A1(n15462), .A2(n12333), .ZN(n13419) );
  INV_X1 U15498 ( .A(n12334), .ZN(n12336) );
  INV_X1 U15499 ( .A(n12469), .ZN(n20030) );
  INV_X1 U15500 ( .A(n12780), .ZN(n12352) );
  NOR2_X1 U15501 ( .A1(n13437), .A2(n19757), .ZN(n12335) );
  AND4_X1 U15502 ( .A1(n12336), .A2(n20047), .A3(n12352), .A4(n12335), .ZN(
        n12507) );
  NAND2_X1 U15503 ( .A1(n12507), .A2(n9759), .ZN(n12337) );
  NAND2_X1 U15504 ( .A1(n19879), .A2(n20047), .ZN(n14120) );
  NAND2_X1 U15505 ( .A1(n9725), .A2(n12564), .ZN(n12343) );
  NAND2_X1 U15506 ( .A1(n13427), .A2(n12343), .ZN(n12545) );
  OR2_X1 U15507 ( .A1(n20010), .A2(n13438), .ZN(n20669) );
  INV_X1 U15508 ( .A(n12345), .ZN(n12357) );
  NAND2_X1 U15509 ( .A1(n12780), .A2(n12180), .ZN(n12346) );
  INV_X1 U15510 ( .A(n20578), .ZN(n15459) );
  NOR2_X1 U15511 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n15810) );
  NAND2_X1 U15512 ( .A1(n15810), .A2(n15822), .ZN(n12532) );
  MUX2_X1 U15513 ( .A(n15459), .B(n12532), .S(n20435), .Z(n12348) );
  INV_X1 U15514 ( .A(n12349), .ZN(n12356) );
  INV_X1 U15515 ( .A(n12350), .ZN(n12351) );
  NAND2_X1 U15516 ( .A1(n13383), .A2(n12351), .ZN(n12354) );
  INV_X1 U15517 ( .A(n15810), .ZN(n14526) );
  NOR2_X1 U15518 ( .A1(n14526), .A2(n15822), .ZN(n12353) );
  NAND2_X1 U15519 ( .A1(n12352), .A2(n20042), .ZN(n13428) );
  NAND4_X1 U15520 ( .A1(n12354), .A2(n12353), .A3(n13428), .A4(n12565), .ZN(
        n12355) );
  NOR2_X1 U15521 ( .A1(n12356), .A2(n12355), .ZN(n12361) );
  OAI21_X1 U15522 ( .B1(n12844), .B2(n12358), .A(n12357), .ZN(n12360) );
  NAND2_X1 U15523 ( .A1(n12537), .A2(n13438), .ZN(n12359) );
  NAND3_X1 U15524 ( .A1(n12361), .A2(n12360), .A3(n12359), .ZN(n12429) );
  INV_X1 U15525 ( .A(n12429), .ZN(n12362) );
  NAND2_X1 U15526 ( .A1(n12394), .A2(n15822), .ZN(n12387) );
  AOI22_X1 U15527 ( .A1(n12709), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n9732), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12366) );
  AOI22_X1 U15528 ( .A1(n9738), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12619), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12365) );
  AOI22_X1 U15529 ( .A1(n13803), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n9757), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12364) );
  AOI22_X1 U15530 ( .A1(n13707), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n13825), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12363) );
  NAND4_X1 U15531 ( .A1(n12366), .A2(n12365), .A3(n12364), .A4(n12363), .ZN(
        n12373) );
  AOI22_X1 U15532 ( .A1(n13843), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n13867), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12371) );
  AOI22_X1 U15533 ( .A1(n12367), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n13718), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12370) );
  AOI22_X1 U15534 ( .A1(n13848), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n9722), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12369) );
  NAND4_X1 U15535 ( .A1(n12371), .A2(n12370), .A3(n12369), .A4(n12368), .ZN(
        n12372) );
  NOR2_X1 U15536 ( .A1(n12630), .A2(n13382), .ZN(n12406) );
  AOI22_X1 U15537 ( .A1(n13803), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12619), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12378) );
  AOI22_X1 U15538 ( .A1(n13868), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n13867), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12377) );
  AOI22_X1 U15539 ( .A1(n13477), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12367), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12376) );
  AOI22_X1 U15540 ( .A1(n13848), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n9722), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12375) );
  NAND4_X1 U15541 ( .A1(n12378), .A2(n12377), .A3(n12376), .A4(n12375), .ZN(
        n12384) );
  AOI22_X1 U15542 ( .A1(n12709), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n9732), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12382) );
  AOI22_X1 U15543 ( .A1(n9739), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(n9755), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12381) );
  AOI22_X1 U15544 ( .A1(n13707), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n13825), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12380) );
  NAND4_X1 U15545 ( .A1(n12382), .A2(n12381), .A3(n12380), .A4(n12379), .ZN(
        n12383) );
  MUX2_X1 U15546 ( .A(n13378), .B(n12406), .S(n12907), .Z(n12385) );
  INV_X1 U15547 ( .A(n12385), .ZN(n12386) );
  INV_X1 U15548 ( .A(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12388) );
  OR2_X1 U15549 ( .A1(n13089), .A2(n12388), .ZN(n12392) );
  NAND2_X1 U15550 ( .A1(n20010), .A2(n12907), .ZN(n12389) );
  NAND2_X1 U15551 ( .A1(n20083), .A2(n20042), .ZN(n12393) );
  NAND2_X1 U15552 ( .A1(n12393), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12401) );
  INV_X1 U15553 ( .A(n12401), .ZN(n12402) );
  INV_X1 U15554 ( .A(n13891), .ZN(n12395) );
  INV_X1 U15555 ( .A(n12677), .ZN(n12750) );
  NAND2_X1 U15556 ( .A1(n12396), .A2(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12398) );
  NAND2_X1 U15557 ( .A1(n13888), .A2(P1_EAX_REG_0__SCAN_IN), .ZN(n12397) );
  OAI211_X1 U15558 ( .C1(n12750), .C2(n12690), .A(n12398), .B(n12397), .ZN(
        n12399) );
  AOI21_X1 U15559 ( .B1(n12394), .B2(n13505), .A(n12399), .ZN(n12400) );
  INV_X1 U15560 ( .A(n12400), .ZN(n12444) );
  OR2_X1 U15561 ( .A1(n12401), .A2(n12400), .ZN(n12446) );
  OAI21_X1 U15562 ( .B1(n12402), .B2(n12444), .A(n12446), .ZN(n12863) );
  OAI222_X1 U15563 ( .A1(n12849), .A2(n14120), .B1(n19879), .B2(n12331), .C1(
        n12863), .C2(n15631), .ZN(P1_U2872) );
  INV_X1 U15564 ( .A(n13378), .ZN(n12404) );
  NAND2_X2 U15565 ( .A1(n12405), .A2(n12404), .ZN(n12639) );
  INV_X1 U15566 ( .A(n12406), .ZN(n12419) );
  AOI22_X1 U15567 ( .A1(n13803), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12619), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12410) );
  AOI22_X1 U15568 ( .A1(n9740), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n13868), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12409) );
  AOI22_X1 U15569 ( .A1(n12709), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n9756), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12408) );
  AOI22_X1 U15570 ( .A1(n13707), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n13825), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12407) );
  NAND4_X1 U15571 ( .A1(n12410), .A2(n12409), .A3(n12408), .A4(n12407), .ZN(
        n12416) );
  AOI22_X1 U15572 ( .A1(n13477), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n13867), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12414) );
  AOI22_X1 U15573 ( .A1(n9732), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12367), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12413) );
  AOI22_X1 U15574 ( .A1(n13848), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n9722), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12412) );
  NAND4_X1 U15575 ( .A1(n12414), .A2(n12413), .A3(n12412), .A4(n12411), .ZN(
        n12415) );
  INV_X1 U15576 ( .A(n12908), .ZN(n12417) );
  OR2_X1 U15577 ( .A1(n12417), .A2(n12632), .ZN(n12418) );
  INV_X1 U15578 ( .A(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12420) );
  OR2_X1 U15579 ( .A1(n13089), .A2(n12420), .ZN(n12421) );
  XNOR2_X2 U15580 ( .A(n12639), .B(n12637), .ZN(n12641) );
  NAND2_X1 U15581 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n12530) );
  OAI21_X1 U15582 ( .B1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n12530), .ZN(n20326) );
  NAND2_X1 U15583 ( .A1(n20578), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n12524) );
  OAI21_X1 U15584 ( .B1(n12532), .B2(n20326), .A(n12524), .ZN(n12423) );
  INV_X1 U15585 ( .A(n12423), .ZN(n12424) );
  AND2_X1 U15586 ( .A1(n12844), .A2(n20038), .ZN(n12544) );
  NOR2_X1 U15587 ( .A1(n12780), .A2(n13891), .ZN(n12426) );
  NAND2_X1 U15588 ( .A1(n12544), .A2(n12426), .ZN(n13436) );
  NAND2_X1 U15589 ( .A1(n9789), .A2(n13436), .ZN(n12427) );
  INV_X1 U15590 ( .A(n20119), .ZN(n12432) );
  INV_X1 U15591 ( .A(n12433), .ZN(n12431) );
  NAND2_X2 U15592 ( .A1(n20055), .A2(n12528), .ZN(n20406) );
  INV_X1 U15593 ( .A(n20406), .ZN(n12434) );
  NAND2_X1 U15594 ( .A1(n12434), .A2(n15822), .ZN(n12437) );
  INV_X1 U15595 ( .A(n12630), .ZN(n12435) );
  NAND2_X1 U15596 ( .A1(n12435), .A2(n12908), .ZN(n12436) );
  AND2_X2 U15597 ( .A1(n12437), .A2(n12436), .ZN(n12906) );
  NAND2_X1 U15598 ( .A1(n12813), .A2(n13505), .ZN(n12443) );
  INV_X1 U15599 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n12440) );
  INV_X1 U15600 ( .A(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n12944) );
  OAI22_X1 U15601 ( .A1(n13753), .A2(n12440), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n12944), .ZN(n12441) );
  AOI21_X1 U15602 ( .B1(n12677), .B2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n12441), .ZN(n12442) );
  NAND2_X1 U15603 ( .A1(n12443), .A2(n12442), .ZN(n12448) );
  OR2_X1 U15604 ( .A1(n12444), .A2(n13886), .ZN(n12445) );
  NAND2_X1 U15605 ( .A1(n12446), .A2(n12445), .ZN(n12447) );
  NAND2_X1 U15606 ( .A1(n12448), .A2(n12447), .ZN(n12685) );
  OAI21_X1 U15607 ( .B1(n12448), .B2(n12447), .A(n12685), .ZN(n12948) );
  INV_X1 U15608 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n12456) );
  MUX2_X1 U15609 ( .A(n13948), .B(n9724), .S(P1_EBX_REG_1__SCAN_IN), .Z(n12454) );
  INV_X2 U15610 ( .A(n9759), .ZN(n13950) );
  NAND2_X1 U15611 ( .A1(n13950), .A2(n13971), .ZN(n12452) );
  XNOR2_X1 U15612 ( .A(n12693), .B(n12455), .ZN(n12938) );
  XNOR2_X1 U15613 ( .A(n12938), .B(n13950), .ZN(n19981) );
  OAI222_X1 U15614 ( .A1(n12948), .A2(n15631), .B1(n19879), .B2(n12456), .C1(
        n14120), .C2(n19981), .ZN(P1_U2871) );
  INV_X1 U15615 ( .A(n12457), .ZN(n12458) );
  NOR2_X1 U15616 ( .A1(n12459), .A2(n12458), .ZN(n12464) );
  INV_X1 U15617 ( .A(n12460), .ZN(n12461) );
  XNOR2_X1 U15618 ( .A(n12462), .B(n12461), .ZN(n19692) );
  INV_X1 U15619 ( .A(n19692), .ZN(n12925) );
  XNOR2_X1 U15620 ( .A(n15105), .B(n12925), .ZN(n12463) );
  NOR2_X1 U15621 ( .A1(n12464), .A2(n12463), .ZN(n12491) );
  AOI21_X1 U15622 ( .B1(n12464), .B2(n12463), .A(n12491), .ZN(n12467) );
  AOI22_X1 U15623 ( .A1(n18930), .A2(n19692), .B1(n18934), .B2(
        P2_EAX_REG_3__SCAN_IN), .ZN(n12466) );
  NAND2_X1 U15624 ( .A1(n18946), .A2(n14711), .ZN(n12465) );
  OAI211_X1 U15625 ( .C1(n12467), .C2(n14714), .A(n12466), .B(n12465), .ZN(
        P2_U2916) );
  AND2_X1 U15626 ( .A1(n20524), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n12868) );
  NAND2_X1 U15627 ( .A1(n15822), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n15816) );
  INV_X1 U15628 ( .A(n15816), .ZN(n12468) );
  NAND2_X1 U15629 ( .A1(n12868), .A2(n12468), .ZN(n20005) );
  INV_X1 U15630 ( .A(n13377), .ZN(n13345) );
  NAND2_X1 U15631 ( .A1(n20010), .A2(n12469), .ZN(n13016) );
  OAI21_X1 U15632 ( .B1(n20669), .B2(n12907), .A(n13016), .ZN(n12470) );
  INV_X1 U15633 ( .A(n12470), .ZN(n12471) );
  OR2_X1 U15634 ( .A1(n12472), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12473) );
  NAND2_X1 U15635 ( .A1(n12472), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13013) );
  AND2_X1 U15636 ( .A1(n12473), .A2(n13013), .ZN(n19995) );
  NAND2_X1 U15637 ( .A1(n12566), .A2(n12474), .ZN(n15447) );
  INV_X1 U15638 ( .A(n19764), .ZN(n19944) );
  INV_X1 U15639 ( .A(P1_REIP_REG_0__SCAN_IN), .ZN(n12475) );
  OR2_X1 U15640 ( .A1(n19845), .A2(n12475), .ZN(n20000) );
  INV_X1 U15641 ( .A(n20000), .ZN(n12480) );
  INV_X1 U15642 ( .A(n20524), .ZN(n20518) );
  NAND2_X1 U15643 ( .A1(n20518), .A2(n12532), .ZN(n20665) );
  NAND2_X1 U15644 ( .A1(n20665), .A2(n15822), .ZN(n12476) );
  INV_X1 U15645 ( .A(n19938), .ZN(n14334) );
  NAND2_X1 U15646 ( .A1(n15822), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n15454) );
  INV_X1 U15647 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n20439) );
  NAND2_X1 U15648 ( .A1(n20439), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n12477) );
  AND2_X1 U15649 ( .A1(n15454), .A2(n12477), .ZN(n12916) );
  INV_X1 U15650 ( .A(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n12478) );
  AOI21_X1 U15651 ( .B1(n14334), .B2(n12916), .A(n12478), .ZN(n12479) );
  AOI211_X1 U15652 ( .C1(n19995), .C2(n19944), .A(n12480), .B(n12479), .ZN(
        n12481) );
  OAI21_X1 U15653 ( .B1(n20005), .B2(n12863), .A(n12481), .ZN(P1_U2999) );
  INV_X1 U15654 ( .A(n12482), .ZN(n12485) );
  INV_X1 U15655 ( .A(n12483), .ZN(n12484) );
  AOI21_X1 U15656 ( .B1(n12485), .B2(n12488), .A(n12484), .ZN(n18890) );
  INV_X1 U15657 ( .A(n18890), .ZN(n12494) );
  NOR2_X1 U15658 ( .A1(n19690), .A2(n19692), .ZN(n12490) );
  OR2_X1 U15659 ( .A1(n12487), .A2(n12486), .ZN(n12489) );
  NAND2_X1 U15660 ( .A1(n12489), .A2(n12488), .ZN(n18897) );
  OAI21_X1 U15661 ( .B1(n12491), .B2(n12490), .A(n18897), .ZN(n12579) );
  INV_X1 U15662 ( .A(n12578), .ZN(n18901) );
  NAND3_X1 U15663 ( .A1(n12579), .A2(n18901), .A3(n15928), .ZN(n12493) );
  AOI22_X1 U15664 ( .A1(n18946), .A2(n14692), .B1(n18934), .B2(
        P2_EAX_REG_5__SCAN_IN), .ZN(n12492) );
  OAI211_X1 U15665 ( .C1(n18937), .C2(n12494), .A(n12493), .B(n12492), .ZN(
        P2_U2914) );
  XNOR2_X1 U15666 ( .A(n12519), .B(n12518), .ZN(n12499) );
  OR2_X1 U15667 ( .A1(n12496), .A2(n12495), .ZN(n12497) );
  NAND2_X1 U15668 ( .A1(n12514), .A2(n12497), .ZN(n18820) );
  MUX2_X1 U15669 ( .A(n18820), .B(n18809), .S(n14602), .Z(n12498) );
  OAI21_X1 U15670 ( .B1(n12499), .B2(n14630), .A(n12498), .ZN(P2_U2876) );
  NAND2_X1 U15671 ( .A1(n12566), .A2(n12844), .ZN(n12550) );
  INV_X1 U15672 ( .A(n20666), .ZN(n20590) );
  OR2_X1 U15673 ( .A1(n12500), .A2(n20590), .ZN(n12501) );
  INV_X1 U15674 ( .A(n12503), .ZN(n15809) );
  NAND2_X1 U15675 ( .A1(n15809), .A2(n20666), .ZN(n12504) );
  NAND2_X1 U15676 ( .A1(n12507), .A2(n12844), .ZN(n12508) );
  NAND2_X1 U15677 ( .A1(n12341), .A2(n12539), .ZN(n12510) );
  NAND2_X2 U15678 ( .A1(n14191), .A2(n12510), .ZN(n14197) );
  INV_X1 U15679 ( .A(n20006), .ZN(n20004) );
  NAND2_X1 U15680 ( .A1(n20004), .A2(DATAI_0_), .ZN(n12512) );
  NAND2_X1 U15681 ( .A1(n20006), .A2(BUF1_REG_0__SCAN_IN), .ZN(n12511) );
  AND2_X1 U15682 ( .A1(n12512), .A2(n12511), .ZN(n20017) );
  INV_X1 U15683 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n19906) );
  OAI222_X1 U15684 ( .A1(n12863), .A2(n14197), .B1(n14193), .B2(n20017), .C1(
        n14191), .C2(n19906), .ZN(P1_U2904) );
  INV_X1 U15685 ( .A(n12900), .ZN(n12513) );
  AOI21_X1 U15686 ( .B1(n12515), .B2(n12514), .A(n12513), .ZN(n18805) );
  INV_X1 U15687 ( .A(n18805), .ZN(n14851) );
  AOI21_X1 U15688 ( .B1(n12519), .B2(n12518), .A(n12517), .ZN(n12520) );
  OR3_X1 U15689 ( .A1(n12516), .A2(n12520), .A3(n14630), .ZN(n12522) );
  NAND2_X1 U15690 ( .A1(n14602), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n12521) );
  OAI211_X1 U15691 ( .C1(n14851), .C2(n14602), .A(n12522), .B(n12521), .ZN(
        P2_U2875) );
  INV_X1 U15692 ( .A(n12523), .ZN(n12526) );
  NAND2_X1 U15693 ( .A1(n12524), .A2(n12553), .ZN(n12525) );
  NAND2_X1 U15694 ( .A1(n12526), .A2(n12525), .ZN(n12527) );
  OR2_X1 U15695 ( .A1(n12648), .A2(n9900), .ZN(n12534) );
  INV_X1 U15696 ( .A(n12530), .ZN(n12529) );
  NAND2_X1 U15697 ( .A1(n12529), .A2(n20321), .ZN(n20367) );
  NAND2_X1 U15698 ( .A1(n12530), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n12531) );
  NAND2_X1 U15699 ( .A1(n20367), .A2(n12531), .ZN(n20018) );
  INV_X1 U15700 ( .A(n12532), .ZN(n12651) );
  AOI22_X1 U15701 ( .A1(n20018), .A2(n12651), .B1(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n20578), .ZN(n12533) );
  NOR2_X1 U15702 ( .A1(n12341), .A2(n13438), .ZN(n12536) );
  OAI21_X1 U15703 ( .B1(n12537), .B2(n12536), .A(n9725), .ZN(n12567) );
  NAND2_X1 U15704 ( .A1(n12357), .A2(n12844), .ZN(n12543) );
  INV_X1 U15705 ( .A(n12538), .ZN(n12542) );
  NAND2_X1 U15706 ( .A1(n12540), .A2(n13438), .ZN(n12541) );
  NAND4_X1 U15707 ( .A1(n12567), .A2(n12543), .A3(n12542), .A4(n12541), .ZN(
        n13431) );
  INV_X1 U15708 ( .A(n13415), .ZN(n12547) );
  NOR2_X1 U15709 ( .A1(n12545), .A2(n12544), .ZN(n12546) );
  NAND2_X1 U15710 ( .A1(n12547), .A2(n12546), .ZN(n12548) );
  NOR2_X1 U15711 ( .A1(n13431), .A2(n12548), .ZN(n12549) );
  NAND2_X1 U15712 ( .A1(n12549), .A2(n12503), .ZN(n14513) );
  INV_X1 U15713 ( .A(n14513), .ZN(n12794) );
  OR2_X1 U15714 ( .A1(n9754), .A2(n12794), .ZN(n12561) );
  INV_X1 U15715 ( .A(n12550), .ZN(n12551) );
  OR2_X1 U15716 ( .A1(n13433), .A2(n12551), .ZN(n12787) );
  INV_X1 U15717 ( .A(n12787), .ZN(n12558) );
  XNOR2_X1 U15718 ( .A(n14515), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12552) );
  INV_X1 U15719 ( .A(n12552), .ZN(n12563) );
  OR3_X1 U15720 ( .A1(n14513), .A2(n12780), .A3(n12552), .ZN(n12557) );
  NAND2_X1 U15721 ( .A1(n13426), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12555) );
  AND2_X1 U15722 ( .A1(n13426), .A2(n12553), .ZN(n14512) );
  INV_X1 U15723 ( .A(n14512), .ZN(n12554) );
  MUX2_X1 U15724 ( .A(n12555), .B(n12554), .S(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n12556) );
  OAI211_X1 U15725 ( .C1(n12558), .C2(n12563), .A(n12557), .B(n12556), .ZN(
        n12559) );
  INV_X1 U15726 ( .A(n12559), .ZN(n12560) );
  NAND2_X1 U15727 ( .A1(n12561), .A2(n12560), .ZN(n12800) );
  INV_X1 U15728 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n19968) );
  NOR2_X1 U15729 ( .A1(n20898), .A2(n19968), .ZN(n14518) );
  INV_X1 U15730 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n12562) );
  AOI22_X1 U15731 ( .A1(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n12449), .B2(n12562), .ZN(
        n14514) );
  INV_X1 U15732 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n20275) );
  AOI222_X1 U15733 ( .A1(n12800), .A2(n15810), .B1(n14518), .B2(n14514), .C1(
        n12563), .C2(n12811), .ZN(n12577) );
  INV_X1 U15734 ( .A(n13419), .ZN(n12573) );
  OR2_X1 U15735 ( .A1(n15490), .A2(n20590), .ZN(n12850) );
  INV_X1 U15736 ( .A(n12850), .ZN(n15452) );
  OAI21_X1 U15737 ( .B1(n13426), .B2(n13415), .A(n15452), .ZN(n12571) );
  OR2_X1 U15738 ( .A1(n12565), .A2(n12564), .ZN(n12570) );
  NAND2_X1 U15739 ( .A1(n12567), .A2(n12566), .ZN(n12569) );
  NAND2_X1 U15740 ( .A1(n12569), .A2(n12568), .ZN(n13418) );
  OAI211_X1 U15741 ( .C1(n15462), .C2(n12571), .A(n12570), .B(n13418), .ZN(
        n12572) );
  NOR2_X1 U15742 ( .A1(n15822), .A2(n15824), .ZN(n12810) );
  NAND2_X1 U15743 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n12810), .ZN(n12575) );
  OAI21_X1 U15744 ( .B1(n15430), .B2(n19757), .A(n12575), .ZN(n15808) );
  AOI21_X1 U15745 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n15822), .A(n15808), 
        .ZN(n14521) );
  NAND2_X1 U15746 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n14521), .ZN(
        n12576) );
  OAI21_X1 U15747 ( .B1(n12577), .B2(n14521), .A(n12576), .ZN(P1_U3472) );
  XNOR2_X1 U15748 ( .A(n12579), .B(n12578), .ZN(n12580) );
  NAND2_X1 U15749 ( .A1(n12580), .A2(n15928), .ZN(n12583) );
  INV_X1 U15750 ( .A(n18897), .ZN(n12581) );
  AOI22_X1 U15751 ( .A1(n18930), .A2(n12581), .B1(n18934), .B2(
        P2_EAX_REG_4__SCAN_IN), .ZN(n12582) );
  OAI211_X1 U15752 ( .C1(n19078), .C2(n12888), .A(n12583), .B(n12582), .ZN(
        P2_U2915) );
  INV_X1 U15753 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n12585) );
  AOI22_X1 U15754 ( .A1(P1_UWORD_REG_6__SCAN_IN), .A2(n20667), .B1(n19903), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n12584) );
  OAI21_X1 U15755 ( .B1(n12585), .B2(n12616), .A(n12584), .ZN(P1_U2914) );
  INV_X1 U15756 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n12587) );
  AOI22_X1 U15757 ( .A1(P1_UWORD_REG_10__SCAN_IN), .A2(n20667), .B1(n19903), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n12586) );
  OAI21_X1 U15758 ( .B1(n12587), .B2(n12616), .A(n12586), .ZN(P1_U2910) );
  INV_X1 U15759 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n12589) );
  AOI22_X1 U15760 ( .A1(P1_UWORD_REG_4__SCAN_IN), .A2(n20667), .B1(n19903), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n12588) );
  OAI21_X1 U15761 ( .B1(n12589), .B2(n12616), .A(n12588), .ZN(P1_U2916) );
  INV_X1 U15762 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n12591) );
  AOI22_X1 U15763 ( .A1(P1_UWORD_REG_5__SCAN_IN), .A2(n20667), .B1(n19903), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n12590) );
  OAI21_X1 U15764 ( .B1(n12591), .B2(n12616), .A(n12590), .ZN(P1_U2915) );
  AND2_X1 U15765 ( .A1(n20669), .A2(n20590), .ZN(n12592) );
  NOR2_X1 U15766 ( .A1(n19912), .A2(n13438), .ZN(n19909) );
  AOI22_X1 U15767 ( .A1(n19909), .A2(P1_EAX_REG_5__SCAN_IN), .B1(
        P1_LWORD_REG_5__SCAN_IN), .B2(n19932), .ZN(n12595) );
  NAND2_X1 U15768 ( .A1(n13150), .A2(n13438), .ZN(n12772) );
  NAND2_X1 U15769 ( .A1(n20004), .A2(DATAI_5_), .ZN(n12594) );
  NAND2_X1 U15770 ( .A1(n20006), .A2(BUF1_REG_5__SCAN_IN), .ZN(n12593) );
  AND2_X1 U15771 ( .A1(n12594), .A2(n12593), .ZN(n20039) );
  INV_X1 U15772 ( .A(n20039), .ZN(n14160) );
  NAND2_X1 U15773 ( .A1(n19920), .A2(n14160), .ZN(n13151) );
  NAND2_X1 U15774 ( .A1(n12595), .A2(n13151), .ZN(P1_U2957) );
  AOI22_X1 U15775 ( .A1(n19909), .A2(P1_EAX_REG_7__SCAN_IN), .B1(
        P1_LWORD_REG_7__SCAN_IN), .B2(n19932), .ZN(n12599) );
  NAND2_X1 U15776 ( .A1(n20004), .A2(DATAI_7_), .ZN(n12597) );
  NAND2_X1 U15777 ( .A1(n20006), .A2(BUF1_REG_7__SCAN_IN), .ZN(n12596) );
  AND2_X1 U15778 ( .A1(n12597), .A2(n12596), .ZN(n20050) );
  INV_X1 U15779 ( .A(n20050), .ZN(n12598) );
  NAND2_X1 U15780 ( .A1(n19920), .A2(n12598), .ZN(n13159) );
  NAND2_X1 U15781 ( .A1(n12599), .A2(n13159), .ZN(P1_U2959) );
  AOI22_X1 U15782 ( .A1(n19909), .A2(P1_EAX_REG_6__SCAN_IN), .B1(
        P1_LWORD_REG_6__SCAN_IN), .B2(n19932), .ZN(n12603) );
  NAND2_X1 U15783 ( .A1(n20004), .A2(DATAI_6_), .ZN(n12601) );
  NAND2_X1 U15784 ( .A1(n20006), .A2(BUF1_REG_6__SCAN_IN), .ZN(n12600) );
  AND2_X1 U15785 ( .A1(n12601), .A2(n12600), .ZN(n20043) );
  INV_X1 U15786 ( .A(n20043), .ZN(n12602) );
  NAND2_X1 U15787 ( .A1(n19920), .A2(n12602), .ZN(n13157) );
  NAND2_X1 U15788 ( .A1(n12603), .A2(n13157), .ZN(P1_U2958) );
  AOI22_X1 U15789 ( .A1(n19909), .A2(P1_EAX_REG_2__SCAN_IN), .B1(
        P1_LWORD_REG_2__SCAN_IN), .B2(n19932), .ZN(n12607) );
  NAND2_X1 U15790 ( .A1(n20004), .A2(DATAI_2_), .ZN(n12605) );
  NAND2_X1 U15791 ( .A1(n20006), .A2(BUF1_REG_2__SCAN_IN), .ZN(n12604) );
  AND2_X1 U15792 ( .A1(n12605), .A2(n12604), .ZN(n20027) );
  INV_X1 U15793 ( .A(n20027), .ZN(n12606) );
  NAND2_X1 U15794 ( .A1(n19920), .A2(n12606), .ZN(n13161) );
  NAND2_X1 U15795 ( .A1(n12607), .A2(n13161), .ZN(P1_U2954) );
  AOI22_X1 U15796 ( .A1(n19909), .A2(P1_EAX_REG_3__SCAN_IN), .B1(
        P1_LWORD_REG_3__SCAN_IN), .B2(n19932), .ZN(n12610) );
  NAND2_X1 U15797 ( .A1(n20004), .A2(DATAI_3_), .ZN(n12609) );
  NAND2_X1 U15798 ( .A1(n20006), .A2(BUF1_REG_3__SCAN_IN), .ZN(n12608) );
  AND2_X1 U15799 ( .A1(n12609), .A2(n12608), .ZN(n20031) );
  INV_X1 U15800 ( .A(n20031), .ZN(n14171) );
  NAND2_X1 U15801 ( .A1(n19920), .A2(n14171), .ZN(n13155) );
  NAND2_X1 U15802 ( .A1(n12610), .A2(n13155), .ZN(P1_U2955) );
  AOI22_X1 U15803 ( .A1(n19909), .A2(P1_EAX_REG_4__SCAN_IN), .B1(
        P1_LWORD_REG_4__SCAN_IN), .B2(n19932), .ZN(n12614) );
  NAND2_X1 U15804 ( .A1(n20004), .A2(DATAI_4_), .ZN(n12612) );
  NAND2_X1 U15805 ( .A1(n20006), .A2(BUF1_REG_4__SCAN_IN), .ZN(n12611) );
  AND2_X1 U15806 ( .A1(n12612), .A2(n12611), .ZN(n20035) );
  INV_X1 U15807 ( .A(n20035), .ZN(n12613) );
  NAND2_X1 U15808 ( .A1(n19920), .A2(n12613), .ZN(n13168) );
  NAND2_X1 U15809 ( .A1(n12614), .A2(n13168), .ZN(P1_U2956) );
  INV_X1 U15810 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n12617) );
  AOI22_X1 U15811 ( .A1(P1_UWORD_REG_14__SCAN_IN), .A2(n20667), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n19903), .ZN(n12615) );
  OAI21_X1 U15812 ( .B1(n12617), .B2(n12616), .A(n12615), .ZN(P1_U2906) );
  AOI22_X1 U15813 ( .A1(n12709), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n9732), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12623) );
  AOI22_X1 U15814 ( .A1(n9741), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12619), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12622) );
  INV_X1 U15815 ( .A(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n20966) );
  AOI22_X1 U15816 ( .A1(n13803), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n9757), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12621) );
  AOI22_X1 U15817 ( .A1(n13707), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n13825), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12620) );
  NAND4_X1 U15818 ( .A1(n12623), .A2(n12622), .A3(n12621), .A4(n12620), .ZN(
        n12629) );
  AOI22_X1 U15819 ( .A1(n13868), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n13867), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12627) );
  AOI22_X1 U15820 ( .A1(n12367), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n13769), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12626) );
  AOI22_X1 U15821 ( .A1(n13848), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n9722), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12625) );
  NAND4_X1 U15822 ( .A1(n12627), .A2(n12626), .A3(n12625), .A4(n12624), .ZN(
        n12628) );
  INV_X1 U15823 ( .A(n12632), .ZN(n12634) );
  AOI22_X1 U15824 ( .A1(n12665), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n12634), .B2(n12633), .ZN(n12635) );
  INV_X1 U15825 ( .A(n12637), .ZN(n12638) );
  INV_X1 U15826 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n12643) );
  INV_X1 U15827 ( .A(n13886), .ZN(n13880) );
  XNOR2_X1 U15828 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n19858) );
  AOI21_X1 U15829 ( .B1(n13880), .B2(n19858), .A(n13887), .ZN(n12642) );
  OAI21_X1 U15830 ( .B1(n13753), .B2(n12643), .A(n12642), .ZN(n12644) );
  AOI21_X1 U15831 ( .B1(n12677), .B2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n12644), .ZN(n12645) );
  NAND2_X1 U15832 ( .A1(n13887), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12647) );
  OR2_X1 U15833 ( .A1(n12648), .A2(n12778), .ZN(n12653) );
  NAND3_X1 U15834 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20514) );
  INV_X1 U15835 ( .A(n20514), .ZN(n20525) );
  NAND2_X1 U15836 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20525), .ZN(
        n20511) );
  NOR3_X1 U15837 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n20321), .A3(
        n20757), .ZN(n20244) );
  INV_X1 U15838 ( .A(n20244), .ZN(n20241) );
  INV_X1 U15839 ( .A(n20261), .ZN(n12649) );
  NAND2_X1 U15840 ( .A1(n20368), .A2(n12649), .ZN(n12650) );
  AOI22_X1 U15841 ( .A1(n20270), .A2(n12651), .B1(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n20578), .ZN(n12652) );
  AOI22_X1 U15842 ( .A1(n12709), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n9732), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12657) );
  AOI22_X1 U15843 ( .A1(n9738), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12619), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12656) );
  AOI22_X1 U15844 ( .A1(n13803), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n9755), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12655) );
  AOI22_X1 U15845 ( .A1(n13707), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n13825), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12654) );
  NAND4_X1 U15846 ( .A1(n12657), .A2(n12656), .A3(n12655), .A4(n12654), .ZN(
        n12664) );
  AOI22_X1 U15847 ( .A1(n13868), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n13867), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12662) );
  AOI22_X1 U15848 ( .A1(n12367), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n13769), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12661) );
  AOI22_X1 U15849 ( .A1(n13848), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n9722), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12660) );
  NAND4_X1 U15850 ( .A1(n12662), .A2(n12661), .A3(n12660), .A4(n12659), .ZN(
        n12663) );
  AOI22_X1 U15851 ( .A1(n12665), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n13086), .B2(n13352), .ZN(n12666) );
  NAND2_X1 U15852 ( .A1(n12668), .A2(n12866), .ZN(n12669) );
  OR2_X1 U15853 ( .A1(n12864), .A2(n13586), .ZN(n12679) );
  INV_X1 U15854 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n12675) );
  NAND2_X1 U15855 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n12671) );
  INV_X1 U15856 ( .A(n12671), .ZN(n12673) );
  INV_X1 U15857 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n12670) );
  INV_X1 U15858 ( .A(n12747), .ZN(n12672) );
  OAI21_X1 U15859 ( .B1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n12673), .A(
        n12672), .ZN(n13247) );
  AOI22_X1 U15860 ( .A1(n13880), .A2(n13247), .B1(n13887), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n12674) );
  OAI21_X1 U15861 ( .B1(n13753), .B2(n12675), .A(n12674), .ZN(n12676) );
  AOI21_X1 U15862 ( .B1(n12677), .B2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n12676), .ZN(n12678) );
  NAND2_X1 U15863 ( .A1(n12679), .A2(n12678), .ZN(n12680) );
  NOR2_X1 U15864 ( .A1(n12681), .A2(n12680), .ZN(n12682) );
  NOR2_X1 U15865 ( .A1(n12775), .A2(n12682), .ZN(n13249) );
  INV_X1 U15866 ( .A(n13249), .ZN(n12702) );
  OAI222_X1 U15867 ( .A1(n12702), .A2(n14197), .B1(n14193), .B2(n20031), .C1(
        n14191), .C2(n12675), .ZN(P1_U2901) );
  NAND2_X1 U15868 ( .A1(n20004), .A2(DATAI_1_), .ZN(n12684) );
  NAND2_X1 U15869 ( .A1(n20006), .A2(BUF1_REG_1__SCAN_IN), .ZN(n12683) );
  AND2_X1 U15870 ( .A1(n12684), .A2(n12683), .ZN(n20023) );
  OAI222_X1 U15871 ( .A1(n12948), .A2(n14197), .B1(n14193), .B2(n20023), .C1(
        n14191), .C2(n12440), .ZN(P1_U2903) );
  NAND2_X1 U15872 ( .A1(n12686), .A2(n12685), .ZN(n12687) );
  AND2_X1 U15873 ( .A1(n12688), .A2(n12687), .ZN(n19867) );
  INV_X1 U15874 ( .A(n19867), .ZN(n12707) );
  OAI222_X1 U15875 ( .A1(n12707), .A2(n14197), .B1(n14193), .B2(n20027), .C1(
        n14191), .C2(n12643), .ZN(P1_U2902) );
  INV_X1 U15876 ( .A(n12394), .ZN(n12819) );
  OAI22_X1 U15877 ( .A1(n12819), .A2(n12794), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n12341), .ZN(n15428) );
  INV_X1 U15878 ( .A(n12811), .ZN(n14524) );
  OAI22_X1 U15879 ( .A1(n20898), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n14524), .ZN(n12689) );
  AOI21_X1 U15880 ( .B1(n15428), .B2(n15810), .A(n12689), .ZN(n12692) );
  NOR2_X1 U15881 ( .A1(n12790), .A2(n12690), .ZN(n15429) );
  AOI22_X1 U15882 ( .A1(n15429), .A2(n15810), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n14521), .ZN(n12691) );
  OAI21_X1 U15883 ( .B1(n12692), .B2(n14521), .A(n12691), .ZN(P1_U3474) );
  AOI21_X1 U15884 ( .B1(n12938), .B2(n9759), .A(n12693), .ZN(n12704) );
  INV_X1 U15885 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n20857) );
  NAND2_X1 U15886 ( .A1(n13940), .A2(n20857), .ZN(n12696) );
  NAND2_X1 U15887 ( .A1(n9724), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12694) );
  OAI211_X1 U15888 ( .C1(n13950), .C2(P1_EBX_REG_2__SCAN_IN), .A(n13944), .B(
        n12694), .ZN(n12695) );
  AND2_X1 U15889 ( .A1(n12696), .A2(n12695), .ZN(n12703) );
  NAND2_X1 U15890 ( .A1(n12704), .A2(n12703), .ZN(n19839) );
  INV_X1 U15891 ( .A(P1_EBX_REG_3__SCAN_IN), .ZN(n12697) );
  NAND2_X1 U15892 ( .A1(n13931), .A2(n12697), .ZN(n12700) );
  INV_X1 U15893 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n13237) );
  NAND2_X1 U15894 ( .A1(n13944), .A2(n13237), .ZN(n12698) );
  OAI211_X1 U15895 ( .C1(n13950), .C2(P1_EBX_REG_3__SCAN_IN), .A(n12698), .B(
        n9724), .ZN(n12699) );
  NAND2_X1 U15896 ( .A1(n12700), .A2(n12699), .ZN(n19841) );
  XNOR2_X1 U15897 ( .A(n19839), .B(n19841), .ZN(n19954) );
  INV_X1 U15898 ( .A(n19879), .ZN(n14111) );
  AOI22_X1 U15899 ( .A1(n19875), .A2(n19954), .B1(n14111), .B2(
        P1_EBX_REG_3__SCAN_IN), .ZN(n12701) );
  OAI21_X1 U15900 ( .B1(n12702), .B2(n15631), .A(n12701), .ZN(P1_U2869) );
  OR2_X1 U15901 ( .A1(n12704), .A2(n12703), .ZN(n12705) );
  AND2_X1 U15902 ( .A1(n12705), .A2(n19839), .ZN(n19967) );
  AOI22_X1 U15903 ( .A1(n19875), .A2(n19967), .B1(n14111), .B2(
        P1_EBX_REG_2__SCAN_IN), .ZN(n12706) );
  OAI21_X1 U15904 ( .B1(n12707), .B2(n15631), .A(n12706), .ZN(P1_U2870) );
  INV_X1 U15905 ( .A(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12708) );
  AOI22_X1 U15906 ( .A1(n12709), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n9732), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12713) );
  AOI22_X1 U15907 ( .A1(n9739), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n12619), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12712) );
  AOI22_X1 U15908 ( .A1(n13803), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n9756), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12711) );
  AOI22_X1 U15909 ( .A1(n13707), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n13825), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12710) );
  NAND4_X1 U15910 ( .A1(n12713), .A2(n12712), .A3(n12711), .A4(n12710), .ZN(
        n12719) );
  AOI22_X1 U15911 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n13867), .B1(
        n13868), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12717) );
  AOI22_X1 U15912 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n12367), .B1(
        n13769), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12716) );
  AOI22_X1 U15913 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n13848), .B1(
        n9722), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12715) );
  NAND4_X1 U15914 ( .A1(n12717), .A2(n12716), .A3(n12715), .A4(n12714), .ZN(
        n12718) );
  NAND2_X1 U15915 ( .A1(n13086), .A2(n13351), .ZN(n12720) );
  INV_X1 U15916 ( .A(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12724) );
  OR2_X1 U15917 ( .A1(n13089), .A2(n12724), .ZN(n12736) );
  AOI22_X1 U15918 ( .A1(n12709), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n9732), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12728) );
  AOI22_X1 U15919 ( .A1(n9740), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12619), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12727) );
  AOI22_X1 U15920 ( .A1(n13803), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n9757), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12726) );
  AOI22_X1 U15921 ( .A1(n13707), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n13825), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12725) );
  NAND4_X1 U15922 ( .A1(n12728), .A2(n12727), .A3(n12726), .A4(n12725), .ZN(
        n12734) );
  AOI22_X1 U15923 ( .A1(n13868), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n13867), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12732) );
  AOI22_X1 U15924 ( .A1(n12367), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n13769), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12731) );
  AOI22_X1 U15925 ( .A1(n13848), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n9722), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12730) );
  NAND4_X1 U15926 ( .A1(n12732), .A2(n12731), .A3(n12730), .A4(n12729), .ZN(
        n12733) );
  NAND2_X1 U15927 ( .A1(n13086), .A2(n13362), .ZN(n12735) );
  NAND2_X1 U15928 ( .A1(n12745), .A2(n9844), .ZN(n12737) );
  AND2_X1 U15929 ( .A1(n13062), .A2(n12737), .ZN(n13350) );
  INV_X1 U15930 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n12740) );
  INV_X1 U15931 ( .A(n12746), .ZN(n12738) );
  INV_X1 U15932 ( .A(n12836), .ZN(n13064) );
  OAI21_X1 U15933 ( .B1(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n12738), .A(
        n13064), .ZN(n19830) );
  AOI22_X1 U15934 ( .A1(n13880), .A2(n19830), .B1(n13887), .B2(
        P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n12739) );
  OAI21_X1 U15935 ( .B1(n13753), .B2(n12740), .A(n12739), .ZN(n12741) );
  NAND2_X1 U15936 ( .A1(n12743), .A2(n12742), .ZN(n12744) );
  NAND2_X1 U15937 ( .A1(n12745), .A2(n12744), .ZN(n13346) );
  OAI21_X1 U15938 ( .B1(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n12747), .A(
        n12746), .ZN(n19947) );
  OAI21_X1 U15939 ( .B1(n20439), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n12396), .ZN(n12749) );
  NAND2_X1 U15940 ( .A1(n13888), .A2(P1_EAX_REG_4__SCAN_IN), .ZN(n12748) );
  OAI211_X1 U15941 ( .C1(n12750), .C2(n15813), .A(n12749), .B(n12748), .ZN(
        n12751) );
  OAI21_X1 U15942 ( .B1(n13886), .B2(n19947), .A(n12751), .ZN(n12752) );
  OAI21_X1 U15943 ( .B1(n13346), .B2(n13586), .A(n12752), .ZN(n12773) );
  NAND2_X1 U15944 ( .A1(n12775), .A2(n12773), .ZN(n12756) );
  NAND2_X1 U15945 ( .A1(n12756), .A2(n12755), .ZN(n12757) );
  AND2_X1 U15946 ( .A1(n13095), .A2(n12757), .ZN(n19832) );
  INV_X1 U15947 ( .A(n19832), .ZN(n12769) );
  OAI222_X1 U15948 ( .A1(n12769), .A2(n14197), .B1(n14193), .B2(n20039), .C1(
        n14191), .C2(n12740), .ZN(P1_U2899) );
  INV_X1 U15949 ( .A(P1_EBX_REG_5__SCAN_IN), .ZN(n12768) );
  INV_X1 U15950 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n19878) );
  NAND2_X1 U15951 ( .A1(n13940), .A2(n19878), .ZN(n12760) );
  NAND2_X1 U15952 ( .A1(n9724), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12758) );
  OAI211_X1 U15953 ( .C1(n13950), .C2(P1_EBX_REG_4__SCAN_IN), .A(n13944), .B(
        n12758), .ZN(n12759) );
  AND2_X1 U15954 ( .A1(n12760), .A2(n12759), .ZN(n19840) );
  NAND2_X1 U15955 ( .A1(n13931), .A2(n12768), .ZN(n12765) );
  NAND2_X1 U15956 ( .A1(n9724), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12762) );
  NAND2_X1 U15957 ( .A1(n13944), .A2(n12762), .ZN(n12763) );
  OAI21_X1 U15958 ( .B1(n13950), .B2(P1_EBX_REG_5__SCAN_IN), .A(n12763), .ZN(
        n12764) );
  AND2_X1 U15959 ( .A1(n19842), .A2(n12766), .ZN(n12767) );
  NOR2_X2 U15960 ( .A1(n19842), .A2(n12766), .ZN(n15789) );
  OR2_X1 U15961 ( .A1(n12767), .A2(n15789), .ZN(n19835) );
  OAI222_X1 U15962 ( .A1(n12769), .A2(n15631), .B1(n19879), .B2(n12768), .C1(
        n14120), .C2(n19835), .ZN(P1_U2867) );
  INV_X1 U15963 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n14190) );
  INV_X1 U15964 ( .A(DATAI_15_), .ZN(n12771) );
  INV_X1 U15965 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n12770) );
  MUX2_X1 U15966 ( .A(n12771), .B(n12770), .S(n20006), .Z(n14192) );
  INV_X1 U15967 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n19881) );
  OAI222_X1 U15968 ( .A1(n13149), .A2(n14190), .B1(n12772), .B2(n14192), .C1(
        n13150), .C2(n19881), .ZN(P1_U2967) );
  INV_X1 U15969 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n19899) );
  INV_X1 U15970 ( .A(n12773), .ZN(n12774) );
  XNOR2_X1 U15971 ( .A(n12775), .B(n12774), .ZN(n19943) );
  INV_X1 U15972 ( .A(n19943), .ZN(n12776) );
  OAI222_X1 U15973 ( .A1(n14191), .A2(n19899), .B1(n14193), .B2(n20035), .C1(
        n14197), .C2(n12776), .ZN(P1_U2900) );
  NAND2_X1 U15974 ( .A1(n20269), .A2(n14513), .ZN(n12796) );
  INV_X1 U15975 ( .A(n12781), .ZN(n12777) );
  OAI21_X1 U15976 ( .B1(n14515), .B2(n12778), .A(n12777), .ZN(n12779) );
  NOR2_X1 U15977 ( .A1(n12779), .A2(n13867), .ZN(n14525) );
  NOR2_X1 U15978 ( .A1(n12780), .A2(n14525), .ZN(n12793) );
  AOI21_X1 U15979 ( .B1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n12782), .A(
        n12781), .ZN(n12791) );
  MUX2_X1 U15980 ( .A(n12783), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n14515), .Z(n12785) );
  NOR2_X1 U15981 ( .A1(n12785), .A2(n12784), .ZN(n12786) );
  NAND2_X1 U15982 ( .A1(n12787), .A2(n12786), .ZN(n12789) );
  NAND2_X1 U15983 ( .A1(n14512), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12788) );
  OAI211_X1 U15984 ( .C1(n12791), .C2(n12790), .A(n12789), .B(n12788), .ZN(
        n12792) );
  AOI21_X1 U15985 ( .B1(n12794), .B2(n12793), .A(n12792), .ZN(n12795) );
  NAND2_X1 U15986 ( .A1(n12796), .A2(n12795), .ZN(n14523) );
  MUX2_X1 U15987 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n14523), .S(
        n12806), .Z(n15442) );
  NAND2_X1 U15988 ( .A1(n15442), .A2(n20898), .ZN(n12798) );
  INV_X1 U15989 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n19765) );
  NAND2_X1 U15990 ( .A1(n19765), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n12801) );
  INV_X1 U15991 ( .A(n12801), .ZN(n12807) );
  NAND2_X1 U15992 ( .A1(n12807), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12797) );
  NAND2_X1 U15993 ( .A1(n12798), .A2(n12797), .ZN(n12803) );
  NAND2_X1 U15994 ( .A1(n15430), .A2(n9900), .ZN(n12799) );
  OAI21_X1 U15995 ( .B1(n12800), .B2(n15430), .A(n12799), .ZN(n15435) );
  OAI22_X1 U15996 ( .A1(n15435), .A2(P1_STATE2_REG_1__SCAN_IN), .B1(n12801), 
        .B2(n9900), .ZN(n12802) );
  NAND2_X1 U15997 ( .A1(n12803), .A2(n12802), .ZN(n15449) );
  INV_X1 U15998 ( .A(n20156), .ZN(n20405) );
  NOR2_X1 U15999 ( .A1(n12804), .A2(n20405), .ZN(n12805) );
  XNOR2_X1 U16000 ( .A(n12805), .B(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n19847) );
  OAI21_X1 U16001 ( .B1(n19847), .B2(n12503), .A(n12806), .ZN(n12809) );
  AOI21_X1 U16002 ( .B1(n15430), .B2(n15813), .A(P1_STATE2_REG_1__SCAN_IN), 
        .ZN(n12808) );
  AOI22_X1 U16003 ( .A1(n12809), .A2(n12808), .B1(
        P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n12807), .ZN(n15448) );
  OAI21_X1 U16004 ( .B1(n15449), .B2(n14516), .A(n15448), .ZN(n12818) );
  OAI21_X1 U16005 ( .B1(n12818), .B2(P1_FLUSH_REG_SCAN_IN), .A(n12810), .ZN(
        n12812) );
  NOR2_X1 U16006 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20670) );
  INV_X1 U16007 ( .A(n20670), .ZN(n15820) );
  NAND2_X1 U16008 ( .A1(n12812), .A2(n20057), .ZN(n20002) );
  NAND2_X1 U16009 ( .A1(n9751), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n12814) );
  NAND2_X1 U16010 ( .A1(n12814), .A2(n20524), .ZN(n20517) );
  NOR2_X1 U16011 ( .A1(n9751), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n12815) );
  AND2_X1 U16012 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n20275), .ZN(n14509) );
  OAI22_X1 U16013 ( .A1(n20517), .A2(n12815), .B1(n20406), .B2(n14509), .ZN(
        n12816) );
  NAND2_X1 U16014 ( .A1(n20002), .A2(n12816), .ZN(n12817) );
  OAI21_X1 U16015 ( .B1(n20002), .B2(n20757), .A(n12817), .ZN(P1_U3477) );
  NOR2_X1 U16016 ( .A1(n12818), .A2(n15824), .ZN(n15457) );
  OAI22_X1 U16017 ( .A1(n20083), .A2(n20518), .B1(n12819), .B2(n14509), .ZN(
        n12820) );
  OAI21_X1 U16018 ( .B1(n15457), .B2(n12820), .A(n20002), .ZN(n12821) );
  OAI21_X1 U16019 ( .B1(n20002), .B2(n20435), .A(n12821), .ZN(P1_U3478) );
  XNOR2_X1 U16020 ( .A(n12823), .B(n12822), .ZN(n19038) );
  XNOR2_X1 U16021 ( .A(n12824), .B(n16147), .ZN(n12825) );
  XNOR2_X1 U16022 ( .A(n12826), .B(n12825), .ZN(n19034) );
  NOR2_X1 U16023 ( .A1(n12926), .A2(n12927), .ZN(n16145) );
  INV_X1 U16024 ( .A(n12929), .ZN(n12827) );
  OAI21_X1 U16025 ( .B1(n16163), .B2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        n12827), .ZN(n16141) );
  NOR2_X1 U16026 ( .A1(n11551), .A2(n18846), .ZN(n12828) );
  AOI221_X1 U16027 ( .B1(n16145), .B2(n16147), .C1(n16141), .C2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A(n12828), .ZN(n12830) );
  NAND2_X1 U16028 ( .A1(n19040), .A2(n16154), .ZN(n12829) );
  OAI211_X1 U16029 ( .C1(n16131), .C2(n18897), .A(n12830), .B(n12829), .ZN(
        n12831) );
  AOI21_X1 U16030 ( .B1(n19034), .B2(n16157), .A(n12831), .ZN(n12832) );
  OAI21_X1 U16031 ( .B1(n19038), .B2(n16139), .A(n12832), .ZN(P2_U3042) );
  NAND2_X1 U16032 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n20670), .ZN(n15463) );
  NAND2_X1 U16033 ( .A1(n13880), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n12833) );
  MUX2_X1 U16034 ( .A(n15463), .B(n12833), .S(n15822), .Z(n12834) );
  NAND2_X1 U16035 ( .A1(n12834), .A2(n19845), .ZN(n12835) );
  INV_X1 U16036 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n12838) );
  INV_X1 U16037 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n15568) );
  INV_X1 U16038 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n12839) );
  INV_X1 U16039 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n12840) );
  INV_X1 U16040 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n13777) );
  INV_X1 U16041 ( .A(n13817), .ZN(n12841) );
  INV_X1 U16042 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n13989) );
  INV_X1 U16043 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n13976) );
  NOR2_X1 U16044 ( .A1(n13861), .A2(n13976), .ZN(n12842) );
  XNOR2_X1 U16045 ( .A(n12842), .B(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14227) );
  NOR2_X1 U16046 ( .A1(n14227), .A2(n20898), .ZN(n12843) );
  NAND2_X1 U16047 ( .A1(n20664), .A2(n12844), .ZN(n12845) );
  NAND2_X1 U16048 ( .A1(n15589), .A2(n12845), .ZN(n19866) );
  INV_X1 U16049 ( .A(n19866), .ZN(n12947) );
  NAND2_X1 U16050 ( .A1(n20664), .A2(n12846), .ZN(n19864) );
  INV_X1 U16051 ( .A(n19864), .ZN(n12939) );
  INV_X1 U16052 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n14069) );
  NOR2_X1 U16053 ( .A1(n13950), .A2(n14069), .ZN(n12855) );
  NAND2_X1 U16054 ( .A1(n20666), .A2(n20439), .ZN(n12847) );
  AND2_X1 U16055 ( .A1(n12855), .A2(n12847), .ZN(n12848) );
  INV_X1 U16056 ( .A(n12849), .ZN(n19992) );
  AOI22_X1 U16057 ( .A1(n12939), .A2(n12394), .B1(n19856), .B2(n19992), .ZN(
        n12861) );
  NAND2_X1 U16058 ( .A1(n13438), .A2(n20666), .ZN(n12851) );
  NAND2_X1 U16059 ( .A1(n12851), .A2(n12850), .ZN(n13414) );
  NAND2_X1 U16060 ( .A1(n13414), .A2(n20439), .ZN(n12853) );
  NOR2_X1 U16061 ( .A1(n12853), .A2(n20010), .ZN(n12852) );
  NAND2_X1 U16062 ( .A1(n19838), .A2(n15545), .ZN(n19826) );
  NAND2_X1 U16063 ( .A1(n19826), .A2(P1_REIP_REG_0__SCAN_IN), .ZN(n12860) );
  INV_X1 U16064 ( .A(n12853), .ZN(n12854) );
  NOR3_X1 U16065 ( .A1(n12855), .A2(n12854), .A3(n20010), .ZN(n12856) );
  NAND2_X1 U16066 ( .A1(n19850), .A2(P1_EBX_REG_0__SCAN_IN), .ZN(n12859) );
  AND2_X1 U16067 ( .A1(n14227), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n12857) );
  OAI21_X1 U16068 ( .B1(n19861), .B2(n19860), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n12858) );
  AND4_X1 U16069 ( .A1(n12861), .A2(n12860), .A3(n12859), .A4(n12858), .ZN(
        n12862) );
  OAI21_X1 U16070 ( .B1(n12947), .B2(n12863), .A(n12862), .ZN(P1_U2840) );
  INV_X1 U16071 ( .A(n20008), .ZN(n12865) );
  OR2_X1 U16072 ( .A1(n20462), .A2(n9751), .ZN(n20401) );
  OAI211_X1 U16073 ( .C1(P1_STATEBS16_REG_SCAN_IN), .C2(n12864), .A(n20377), 
        .B(n20401), .ZN(n12870) );
  INV_X1 U16074 ( .A(n20269), .ZN(n12882) );
  NOR2_X1 U16075 ( .A1(n12882), .A2(n14509), .ZN(n12869) );
  INV_X1 U16076 ( .A(n12866), .ZN(n12867) );
  NAND2_X1 U16077 ( .A1(n9751), .A2(n12868), .ZN(n14507) );
  NOR2_X1 U16078 ( .A1(n20239), .A2(n14507), .ZN(n20243) );
  AOI211_X1 U16079 ( .C1(n20524), .C2(n12870), .A(n12869), .B(n20243), .ZN(
        n12873) );
  INV_X1 U16080 ( .A(n20002), .ZN(n12872) );
  NAND2_X1 U16081 ( .A1(n12872), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n12871) );
  OAI21_X1 U16082 ( .B1(n12873), .B2(n12872), .A(n12871), .ZN(P1_U3475) );
  NAND2_X1 U16083 ( .A1(n13249), .A2(n19866), .ZN(n12881) );
  INV_X1 U16084 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n12917) );
  NAND2_X1 U16085 ( .A1(n19857), .A2(n12917), .ZN(n12941) );
  NAND2_X1 U16086 ( .A1(n12941), .A2(n15545), .ZN(n19855) );
  NAND2_X1 U16087 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(P1_REIP_REG_2__SCAN_IN), 
        .ZN(n12874) );
  OAI211_X1 U16088 ( .C1(P1_REIP_REG_3__SCAN_IN), .C2(P1_REIP_REG_2__SCAN_IN), 
        .A(n12874), .B(P1_REIP_REG_1__SCAN_IN), .ZN(n12878) );
  AOI22_X1 U16089 ( .A1(n19856), .A2(n19954), .B1(n19850), .B2(
        P1_EBX_REG_3__SCAN_IN), .ZN(n12877) );
  INV_X1 U16090 ( .A(n13247), .ZN(n12875) );
  AOI22_X1 U16091 ( .A1(n12875), .A2(n19860), .B1(n19861), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n12876) );
  OAI211_X1 U16092 ( .C1(n19838), .C2(n12878), .A(n12877), .B(n12876), .ZN(
        n12879) );
  AOI21_X1 U16093 ( .B1(P1_REIP_REG_3__SCAN_IN), .B2(n19855), .A(n12879), .ZN(
        n12880) );
  OAI211_X1 U16094 ( .C1(n12882), .C2(n19864), .A(n12881), .B(n12880), .ZN(
        P1_U2837) );
  INV_X1 U16095 ( .A(n15015), .ZN(n12883) );
  OR2_X1 U16096 ( .A1(n12884), .A2(n12883), .ZN(n12886) );
  INV_X1 U16097 ( .A(n13110), .ZN(n12885) );
  AND2_X1 U16098 ( .A1(n12886), .A2(n12885), .ZN(n18773) );
  INV_X1 U16099 ( .A(n18773), .ZN(n12889) );
  OAI222_X1 U16100 ( .A1(n12890), .A2(n18948), .B1(n12889), .B2(n18937), .C1(
        n12888), .C2(n12887), .ZN(P2_U2904) );
  AND2_X1 U16101 ( .A1(n12516), .A2(n12898), .ZN(n12892) );
  OAI211_X1 U16102 ( .C1(n12892), .C2(n12891), .A(n14601), .B(n13040), .ZN(
        n12896) );
  INV_X1 U16103 ( .A(n12901), .ZN(n12894) );
  AOI21_X1 U16104 ( .B1(n10194), .B2(n12894), .A(n9768), .ZN(n18784) );
  NAND2_X1 U16105 ( .A1(n18784), .A2(n14621), .ZN(n12895) );
  OAI211_X1 U16106 ( .C1(n14621), .C2(n12897), .A(n12896), .B(n12895), .ZN(
        P2_U2873) );
  XNOR2_X1 U16107 ( .A(n12516), .B(n12898), .ZN(n12905) );
  AND2_X1 U16108 ( .A1(n12900), .A2(n12899), .ZN(n12902) );
  OR2_X1 U16109 ( .A1(n12902), .A2(n12901), .ZN(n18797) );
  INV_X1 U16110 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n12903) );
  MUX2_X1 U16111 ( .A(n18797), .B(n12903), .S(n14602), .Z(n12904) );
  OAI21_X1 U16112 ( .B1(n12905), .B2(n14630), .A(n12904), .ZN(P2_U2874) );
  NAND2_X1 U16113 ( .A1(n12906), .A2(n13438), .ZN(n12913) );
  NAND2_X1 U16114 ( .A1(n12907), .A2(n12908), .ZN(n13239) );
  OAI21_X1 U16115 ( .B1(n12908), .B2(n12907), .A(n13239), .ZN(n12910) );
  OAI211_X1 U16116 ( .C1(n12910), .C2(n20669), .A(n12118), .B(n12121), .ZN(
        n12911) );
  INV_X1 U16117 ( .A(n12911), .ZN(n12912) );
  XNOR2_X1 U16118 ( .A(n13013), .B(n13011), .ZN(n12914) );
  NAND2_X1 U16119 ( .A1(n12914), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13015) );
  OAI21_X1 U16120 ( .B1(n12914), .B2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n13015), .ZN(n12915) );
  INV_X1 U16121 ( .A(n12915), .ZN(n19986) );
  NOR2_X1 U16122 ( .A1(n19845), .A2(n12917), .ZN(n19982) );
  AOI21_X1 U16123 ( .B1(n19938), .B2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n19982), .ZN(n12918) );
  OAI21_X1 U16124 ( .B1(n15701), .B2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n12918), .ZN(n12919) );
  AOI21_X1 U16125 ( .B1(n19986), .B2(n19944), .A(n12919), .ZN(n12920) );
  OAI21_X1 U16126 ( .B1(n20005), .B2(n12948), .A(n12920), .ZN(P1_U2998) );
  NAND2_X1 U16127 ( .A1(n12922), .A2(n12921), .ZN(n12923) );
  XOR2_X1 U16128 ( .A(n12924), .B(n12923), .Z(n16061) );
  INV_X1 U16129 ( .A(n16061), .ZN(n12937) );
  OAI22_X1 U16130 ( .A1(n16131), .A2(n12925), .B1(n11002), .B2(n18846), .ZN(
        n12931) );
  INV_X1 U16131 ( .A(n12926), .ZN(n12928) );
  MUX2_X1 U16132 ( .A(n12929), .B(n12928), .S(n12927), .Z(n12930) );
  AOI211_X1 U16133 ( .C1(n16154), .C2(n15103), .A(n12931), .B(n12930), .ZN(
        n12936) );
  OR2_X1 U16134 ( .A1(n12933), .A2(n12932), .ZN(n16056) );
  NAND3_X1 U16135 ( .A1(n16056), .A2(n16157), .A3(n12934), .ZN(n12935) );
  OAI211_X1 U16136 ( .C1(n12937), .C2(n16139), .A(n12936), .B(n12935), .ZN(
        P2_U3043) );
  INV_X1 U16137 ( .A(n20406), .ZN(n20465) );
  AOI22_X1 U16138 ( .A1(n12939), .A2(n20465), .B1(n19856), .B2(n12938), .ZN(
        n12946) );
  INV_X1 U16139 ( .A(n15545), .ZN(n19828) );
  AOI22_X1 U16140 ( .A1(P1_EBX_REG_1__SCAN_IN), .A2(n19850), .B1(n19828), .B2(
        P1_REIP_REG_1__SCAN_IN), .ZN(n12940) );
  OAI21_X1 U16141 ( .B1(n19823), .B2(n12944), .A(n12940), .ZN(n12943) );
  INV_X1 U16142 ( .A(n12941), .ZN(n12942) );
  AOI211_X1 U16143 ( .C1(n19860), .C2(n12944), .A(n12943), .B(n12942), .ZN(
        n12945) );
  OAI211_X1 U16144 ( .C1(n12948), .C2(n12947), .A(n12946), .B(n12945), .ZN(
        P1_U2839) );
  INV_X1 U16145 ( .A(n18913), .ZN(n12974) );
  AOI21_X1 U16146 ( .B1(n16065), .B2(n11957), .A(n15403), .ZN(n16053) );
  OAI22_X1 U16147 ( .A1(n18954), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(P2_STATE2_REG_0__SCAN_IN), .ZN(
        n13194) );
  OAI22_X1 U16148 ( .A1(n18954), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(
        n13174), .B2(P2_STATE2_REG_0__SCAN_IN), .ZN(n13181) );
  AND2_X1 U16149 ( .A1(n13194), .A2(n13181), .ZN(n13032) );
  NAND2_X1 U16150 ( .A1(n13032), .A2(n13034), .ZN(n15401) );
  NAND2_X1 U16151 ( .A1(n18863), .A2(n15401), .ZN(n12952) );
  XNOR2_X1 U16152 ( .A(n16053), .B(n12952), .ZN(n12953) );
  NOR4_X1 U16153 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(P2_STATEBS16_REG_SCAN_IN), .A4(n13196), .ZN(n18794) );
  INV_X1 U16154 ( .A(n18794), .ZN(n19614) );
  NAND2_X1 U16155 ( .A1(n12953), .A2(n10036), .ZN(n12973) );
  NAND2_X1 U16156 ( .A1(n12954), .A2(n19736), .ZN(n12955) );
  NAND2_X1 U16157 ( .A1(n12956), .A2(n12955), .ZN(n12967) );
  INV_X1 U16158 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n15830) );
  NAND2_X1 U16159 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19744), .ZN(n19100) );
  NOR2_X1 U16160 ( .A1(n12957), .A2(n19100), .ZN(n16194) );
  OR2_X1 U16161 ( .A1(n19033), .A2(n18794), .ZN(n12958) );
  OR2_X1 U16162 ( .A1(n16194), .A2(n12958), .ZN(n12959) );
  NOR2_X1 U16163 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n12960), .ZN(n12966) );
  NAND2_X1 U16164 ( .A1(n11164), .A2(n12966), .ZN(n12961) );
  NOR2_X1 U16165 ( .A1(n10425), .A2(n12961), .ZN(n16198) );
  INV_X1 U16166 ( .A(n12962), .ZN(n12963) );
  AOI22_X1 U16167 ( .A1(n18918), .A2(P2_REIP_REG_3__SCAN_IN), .B1(n18917), 
        .B2(n19692), .ZN(n12964) );
  OAI21_X1 U16168 ( .B1(n12965), .B2(n18923), .A(n12964), .ZN(n12971) );
  OR2_X1 U16169 ( .A1(n18951), .A2(n12966), .ZN(n15829) );
  OR2_X1 U16170 ( .A1(n12967), .A2(P2_EBX_REG_31__SCAN_IN), .ZN(n12968) );
  NAND2_X1 U16171 ( .A1(n15829), .A2(n12968), .ZN(n18919) );
  INV_X1 U16172 ( .A(n18919), .ZN(n18810) );
  NOR2_X2 U16173 ( .A1(n18918), .A2(n19714), .ZN(n18882) );
  OAI22_X1 U16174 ( .A1(n18810), .A2(n12969), .B1(n16065), .B2(n18911), .ZN(
        n12970) );
  AOI211_X1 U16175 ( .C1(n18925), .C2(n15103), .A(n12971), .B(n12970), .ZN(
        n12972) );
  OAI211_X1 U16176 ( .C1(n12974), .C2(n15105), .A(n12973), .B(n12972), .ZN(
        P2_U2852) );
  AND2_X1 U16177 ( .A1(n12985), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n12975) );
  NAND2_X1 U16178 ( .A1(n11214), .A2(n12975), .ZN(n12982) );
  AND2_X1 U16179 ( .A1(n19226), .A2(n19553), .ZN(n19684) );
  NOR2_X1 U16180 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n19746) );
  AOI221_X4 U16181 ( .B1(n19746), .B2(n15104), .C1(n19719), .C2(n15104), .A(
        P2_STATE2_REG_0__SCAN_IN), .ZN(n19549) );
  OAI21_X1 U16182 ( .B1(n12981), .B2(n19684), .A(n19549), .ZN(n12977) );
  AOI21_X1 U16183 ( .B1(n12985), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n12977), 
        .ZN(n12978) );
  NAND2_X1 U16184 ( .A1(n12982), .A2(n12978), .ZN(n19292) );
  INV_X1 U16185 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n16308) );
  INV_X1 U16186 ( .A(BUF2_REG_21__SCAN_IN), .ZN(n18042) );
  INV_X1 U16187 ( .A(n19553), .ZN(n13214) );
  AOI22_X1 U16188 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n19090), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n19089), .ZN(n19498) );
  INV_X1 U16189 ( .A(n19498), .ZN(n19585) );
  AOI22_X1 U16190 ( .A1(n19329), .A2(n19529), .B1(n19297), .B2(n19585), .ZN(
        n12988) );
  INV_X1 U16191 ( .A(n12981), .ZN(n19255) );
  INV_X1 U16192 ( .A(n19100), .ZN(n19257) );
  INV_X1 U16193 ( .A(n12982), .ZN(n12983) );
  AOI211_X2 U16194 ( .C1(n19255), .C2(n19744), .A(n19257), .B(n12983), .ZN(
        n19296) );
  NOR2_X2 U16195 ( .A1(n12984), .A2(n19426), .ZN(n19584) );
  INV_X1 U16196 ( .A(n12985), .ZN(n19307) );
  NAND2_X1 U16197 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19549), .ZN(n19084) );
  NOR2_X2 U16198 ( .A1(n12986), .A2(n19084), .ZN(n19583) );
  AOI22_X1 U16199 ( .A1(n19296), .A2(n19584), .B1(n19307), .B2(n19583), .ZN(
        n12987) );
  OAI211_X1 U16200 ( .C1(n19301), .C2(n12989), .A(n12988), .B(n12987), .ZN(
        P2_U3109) );
  INV_X1 U16201 ( .A(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12994) );
  INV_X1 U16202 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n16315) );
  INV_X1 U16203 ( .A(BUF2_REG_16__SCAN_IN), .ZN(n18018) );
  AOI22_X1 U16204 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n19089), .B1(
        BUF1_REG_24__SCAN_IN), .B2(n19090), .ZN(n19468) );
  INV_X1 U16205 ( .A(n19468), .ZN(n19555) );
  AOI22_X1 U16206 ( .A1(n19329), .A2(n19465), .B1(n19297), .B2(n19555), .ZN(
        n12993) );
  AND2_X1 U16207 ( .A1(n19740), .A2(n19076), .ZN(n19547) );
  AOI22_X1 U16208 ( .A1(n19296), .A2(n12991), .B1(n19307), .B2(n19547), .ZN(
        n12992) );
  OAI211_X1 U16209 ( .C1(n19301), .C2(n12994), .A(n12993), .B(n12992), .ZN(
        P2_U3104) );
  NOR2_X1 U16210 ( .A1(n15105), .A2(n12954), .ZN(n19552) );
  NAND2_X1 U16211 ( .A1(n19552), .A2(n19162), .ZN(n12995) );
  NOR2_X1 U16212 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n19697), .ZN(
        n19335) );
  NAND2_X1 U16213 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19335), .ZN(
        n13003) );
  NAND2_X1 U16214 ( .A1(n12995), .A2(n13003), .ZN(n13002) );
  INV_X1 U16215 ( .A(n19163), .ZN(n12996) );
  NAND2_X1 U16216 ( .A1(n19335), .A2(n12996), .ZN(n12997) );
  INV_X1 U16217 ( .A(n12997), .ZN(n19413) );
  AND2_X1 U16218 ( .A1(n12997), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n12998) );
  NAND2_X1 U16219 ( .A1(n12999), .A2(n12998), .ZN(n13005) );
  OAI211_X1 U16220 ( .C1(n19714), .C2(n19413), .A(n19549), .B(n13005), .ZN(
        n13000) );
  INV_X1 U16221 ( .A(n13000), .ZN(n13001) );
  NAND2_X1 U16222 ( .A1(n13002), .A2(n13001), .ZN(n19415) );
  INV_X1 U16223 ( .A(n19415), .ZN(n19412) );
  INV_X1 U16224 ( .A(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n13008) );
  INV_X1 U16225 ( .A(n19450), .ZN(n19425) );
  NOR2_X2 U16226 ( .A1(n19424), .A2(n19686), .ZN(n19409) );
  AOI22_X1 U16227 ( .A1(n19425), .A2(n19465), .B1(n19409), .B2(n19555), .ZN(
        n13007) );
  OAI21_X1 U16228 ( .B1(n13003), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n19744), 
        .ZN(n13004) );
  AOI22_X1 U16229 ( .A1(n19414), .A2(n12991), .B1(n19413), .B2(n19547), .ZN(
        n13006) );
  OAI211_X1 U16230 ( .C1(n19412), .C2(n13008), .A(n13007), .B(n13006), .ZN(
        P2_U3136) );
  AOI22_X1 U16231 ( .A1(n19938), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B1(
        n13009), .B2(P1_REIP_REG_2__SCAN_IN), .ZN(n13010) );
  OAI21_X1 U16232 ( .B1(n15701), .B2(n19858), .A(n13010), .ZN(n13025) );
  INV_X1 U16233 ( .A(n13011), .ZN(n13012) );
  OR2_X1 U16234 ( .A1(n13013), .A2(n13012), .ZN(n13014) );
  INV_X1 U16235 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n20722) );
  XNOR2_X1 U16236 ( .A(n13239), .B(n13238), .ZN(n13018) );
  INV_X1 U16237 ( .A(n13016), .ZN(n13017) );
  AOI21_X1 U16238 ( .B1(n13018), .B2(n13383), .A(n13017), .ZN(n13019) );
  NAND2_X1 U16239 ( .A1(n13020), .A2(n13019), .ZN(n13021) );
  NOR2_X1 U16240 ( .A1(n13022), .A2(n13021), .ZN(n19965) );
  INV_X1 U16241 ( .A(n13236), .ZN(n13023) );
  NOR3_X1 U16242 ( .A1(n19965), .A2(n13023), .A3(n19764), .ZN(n13024) );
  AOI211_X1 U16243 ( .C1(n9727), .C2(n19867), .A(n13025), .B(n13024), .ZN(
        n13026) );
  INV_X1 U16244 ( .A(n13026), .ZN(P1_U2997) );
  INV_X1 U16245 ( .A(n18925), .ZN(n18894) );
  NAND2_X1 U16246 ( .A1(n18918), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n13028) );
  AOI22_X1 U16247 ( .A1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n18882), .B1(
        P2_EBX_REG_2__SCAN_IN), .B2(n18919), .ZN(n13027) );
  OAI211_X1 U16248 ( .C1(n18923), .C2(n13029), .A(n13028), .B(n13027), .ZN(
        n13030) );
  AOI21_X1 U16249 ( .B1(n19702), .B2(n18917), .A(n13030), .ZN(n13031) );
  OAI21_X1 U16250 ( .B1(n11148), .B2(n18894), .A(n13031), .ZN(n13037) );
  INV_X1 U16251 ( .A(n13034), .ZN(n13035) );
  NOR2_X1 U16252 ( .A1(n18903), .A2(n13032), .ZN(n13180) );
  INV_X1 U16253 ( .A(n13180), .ZN(n13033) );
  AOI221_X1 U16254 ( .B1(n13035), .B2(n13180), .C1(n13034), .C2(n13033), .A(
        n19614), .ZN(n13036) );
  AOI211_X1 U16255 ( .C1(n13215), .C2(n18913), .A(n13037), .B(n13036), .ZN(
        n13038) );
  INV_X1 U16256 ( .A(n13038), .ZN(P2_U2853) );
  XNOR2_X1 U16257 ( .A(n13040), .B(n13039), .ZN(n13045) );
  INV_X1 U16258 ( .A(n13041), .ZN(n13042) );
  OAI21_X1 U16259 ( .B1(n9768), .B2(n13042), .A(n9842), .ZN(n18776) );
  MUX2_X1 U16260 ( .A(n13043), .B(n18776), .S(n14582), .Z(n13044) );
  OAI21_X1 U16261 ( .B1(n13045), .B2(n14630), .A(n13044), .ZN(P2_U2872) );
  INV_X1 U16262 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n19896) );
  INV_X1 U16263 ( .A(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n13046) );
  OR2_X1 U16264 ( .A1(n13089), .A2(n13046), .ZN(n13058) );
  AOI22_X1 U16265 ( .A1(n12709), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n9732), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n13050) );
  AOI22_X1 U16266 ( .A1(n9741), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12619), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n13049) );
  INV_X1 U16267 ( .A(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n20841) );
  AOI22_X1 U16268 ( .A1(n13803), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n9755), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n13048) );
  AOI22_X1 U16269 ( .A1(n13707), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n13825), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n13047) );
  NAND4_X1 U16270 ( .A1(n13050), .A2(n13049), .A3(n13048), .A4(n13047), .ZN(
        n13056) );
  AOI22_X1 U16271 ( .A1(n13868), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n13867), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n13054) );
  AOI22_X1 U16272 ( .A1(n12367), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n13769), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n13053) );
  AOI22_X1 U16273 ( .A1(n13848), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n9722), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n13052) );
  NAND4_X1 U16274 ( .A1(n13054), .A2(n13053), .A3(n13052), .A4(n13051), .ZN(
        n13055) );
  NAND2_X1 U16275 ( .A1(n13086), .A2(n13371), .ZN(n13057) );
  NAND2_X1 U16276 ( .A1(n13058), .A2(n13057), .ZN(n13060) );
  INV_X1 U16277 ( .A(n13060), .ZN(n13061) );
  NAND2_X1 U16278 ( .A1(n13062), .A2(n13061), .ZN(n13063) );
  INV_X1 U16279 ( .A(n13091), .ZN(n13067) );
  INV_X1 U16280 ( .A(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n13065) );
  NAND2_X1 U16281 ( .A1(n13065), .A2(n13064), .ZN(n13066) );
  NAND2_X1 U16282 ( .A1(n13067), .A2(n13066), .ZN(n19813) );
  AOI22_X1 U16283 ( .A1(n19813), .A2(n13880), .B1(n13887), .B2(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n13068) );
  OAI21_X1 U16284 ( .B1(n13753), .B2(n19896), .A(n13068), .ZN(n13069) );
  XOR2_X1 U16285 ( .A(n13095), .B(n13096), .Z(n19872) );
  INV_X1 U16286 ( .A(n19872), .ZN(n13070) );
  OAI222_X1 U16287 ( .A1(n14191), .A2(n19896), .B1(n14193), .B2(n20043), .C1(
        n14197), .C2(n13070), .ZN(P1_U2898) );
  NOR2_X1 U16288 ( .A1(n19337), .A2(n19131), .ZN(n13071) );
  NOR2_X1 U16289 ( .A1(n19337), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19303) );
  AOI21_X1 U16290 ( .B1(n19604), .B2(n13071), .A(n19303), .ZN(n13077) );
  NOR2_X1 U16291 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19096) );
  NAND2_X1 U16292 ( .A1(n19096), .A2(n10862), .ZN(n19104) );
  NOR2_X1 U16293 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19104), .ZN(
        n19086) );
  INV_X1 U16294 ( .A(n13072), .ZN(n13073) );
  AND2_X1 U16295 ( .A1(n13073), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19595) );
  NOR2_X1 U16296 ( .A1(n19086), .A2(n19595), .ZN(n13081) );
  OAI21_X1 U16297 ( .B1(n13074), .B2(n19086), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n13075) );
  OAI21_X1 U16298 ( .B1(n13077), .B2(n13081), .A(n13075), .ZN(n19091) );
  INV_X1 U16299 ( .A(n19091), .ZN(n13213) );
  NOR2_X2 U16300 ( .A1(n13076), .A2(n19426), .ZN(n19560) );
  INV_X1 U16301 ( .A(n19560), .ZN(n19470) );
  INV_X1 U16302 ( .A(n13077), .ZN(n13082) );
  AOI21_X1 U16303 ( .B1(n13078), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n13079) );
  OAI21_X1 U16304 ( .B1(n19086), .B2(n13079), .A(n19549), .ZN(n13080) );
  INV_X1 U16305 ( .A(n19095), .ZN(n13211) );
  INV_X1 U16306 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n20967) );
  INV_X1 U16307 ( .A(BUF2_REG_25__SCAN_IN), .ZN(n20723) );
  OAI22_X2 U16308 ( .A1(n20967), .A2(n19080), .B1(n20723), .B2(n19079), .ZN(
        n19561) );
  INV_X1 U16309 ( .A(n19561), .ZN(n19474) );
  AOI22_X1 U16310 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n19090), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n19089), .ZN(n19564) );
  INV_X1 U16311 ( .A(n19564), .ZN(n19515) );
  AOI22_X1 U16312 ( .A1(n19515), .A2(n19131), .B1(n19086), .B2(n19559), .ZN(
        n13083) );
  OAI21_X1 U16313 ( .B1(n19474), .B2(n19604), .A(n13083), .ZN(n13084) );
  AOI21_X1 U16314 ( .B1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B2(n13211), .A(
        n13084), .ZN(n13085) );
  OAI21_X1 U16315 ( .B1(n13213), .B2(n19470), .A(n13085), .ZN(P2_U3049) );
  INV_X1 U16316 ( .A(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13088) );
  NAND2_X1 U16317 ( .A1(n13086), .A2(n13382), .ZN(n13087) );
  OAI21_X1 U16318 ( .B1(n13089), .B2(n13088), .A(n13087), .ZN(n13090) );
  INV_X1 U16319 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n13093) );
  OAI21_X1 U16320 ( .B1(n13091), .B2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .A(
        n13129), .ZN(n19807) );
  AOI22_X1 U16321 ( .A1(n19807), .A2(n13880), .B1(n13887), .B2(
        P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n13092) );
  OAI21_X1 U16322 ( .B1(n13753), .B2(n13093), .A(n13092), .ZN(n13094) );
  AOI21_X1 U16323 ( .B1(n13098), .B2(n13097), .A(n13133), .ZN(n19809) );
  INV_X1 U16324 ( .A(n19809), .ZN(n13107) );
  INV_X1 U16325 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n13106) );
  INV_X1 U16326 ( .A(P1_EBX_REG_6__SCAN_IN), .ZN(n19874) );
  NAND2_X1 U16327 ( .A1(n13940), .A2(n19874), .ZN(n13101) );
  NAND2_X1 U16328 ( .A1(n9724), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13099) );
  OAI211_X1 U16329 ( .C1(n13950), .C2(P1_EBX_REG_6__SCAN_IN), .A(n13944), .B(
        n13099), .ZN(n13100) );
  NAND2_X1 U16330 ( .A1(n13931), .A2(n13106), .ZN(n13105) );
  NAND2_X1 U16331 ( .A1(n9724), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n13102) );
  NAND2_X1 U16332 ( .A1(n13944), .A2(n13102), .ZN(n13103) );
  OAI21_X1 U16333 ( .B1(n13950), .B2(P1_EBX_REG_7__SCAN_IN), .A(n13103), .ZN(
        n13104) );
  OAI21_X1 U16334 ( .B1(n9848), .B2(n9877), .A(n13145), .ZN(n19812) );
  OAI222_X1 U16335 ( .A1(n13107), .A2(n15631), .B1(n19879), .B2(n13106), .C1(
        n19812), .C2(n14120), .ZN(P1_U2865) );
  OAI222_X1 U16336 ( .A1(n13107), .A2(n14197), .B1(n14193), .B2(n20050), .C1(
        n14191), .C2(n13093), .ZN(P1_U2897) );
  AOI21_X1 U16337 ( .B1(n13109), .B2(n13108), .A(n13289), .ZN(n13229) );
  INV_X1 U16338 ( .A(n13229), .ZN(n13117) );
  OR2_X1 U16339 ( .A1(n13111), .A2(n13110), .ZN(n13112) );
  NAND2_X1 U16340 ( .A1(n13112), .A2(n13290), .ZN(n18764) );
  INV_X1 U16341 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n18988) );
  OAI22_X1 U16342 ( .A1(n14709), .A2(n18764), .B1(n18988), .B2(n18948), .ZN(
        n13113) );
  AOI21_X1 U16343 ( .B1(n15927), .B2(n13114), .A(n13113), .ZN(n13116) );
  AOI22_X1 U16344 ( .A1(n18929), .A2(BUF2_REG_16__SCAN_IN), .B1(n18931), .B2(
        BUF1_REG_16__SCAN_IN), .ZN(n13115) );
  OAI211_X1 U16345 ( .C1(n13117), .C2(n14714), .A(n13116), .B(n13115), .ZN(
        P2_U2903) );
  INV_X1 U16346 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n13138) );
  AOI22_X1 U16347 ( .A1(n13707), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n9732), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n13121) );
  AOI22_X1 U16348 ( .A1(n13867), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12619), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n13120) );
  AOI22_X1 U16349 ( .A1(n13803), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n9756), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n13119) );
  AOI22_X1 U16350 ( .A1(n13848), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n9722), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13118) );
  NAND4_X1 U16351 ( .A1(n13121), .A2(n13120), .A3(n13119), .A4(n13118), .ZN(
        n13127) );
  AOI22_X1 U16352 ( .A1(n13464), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n13868), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n13125) );
  AOI22_X1 U16353 ( .A1(n9738), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12367), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n13124) );
  AOI22_X1 U16354 ( .A1(n12709), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n13825), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n13123) );
  NAND4_X1 U16355 ( .A1(n13125), .A2(n13124), .A3(n13123), .A4(n13122), .ZN(
        n13126) );
  OR2_X1 U16356 ( .A1(n13127), .A2(n13126), .ZN(n13128) );
  NAND2_X1 U16357 ( .A1(n13505), .A2(n13128), .ZN(n13131) );
  XNOR2_X1 U16358 ( .A(n13129), .B(n19793), .ZN(n19796) );
  AOI22_X1 U16359 ( .A1(n19796), .A2(n13880), .B1(n13887), .B2(
        P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n13130) );
  OAI211_X1 U16360 ( .C1(n13753), .C2(n13138), .A(n13131), .B(n13130), .ZN(
        n13132) );
  INV_X1 U16361 ( .A(n13132), .ZN(n13135) );
  INV_X1 U16362 ( .A(n13133), .ZN(n13134) );
  AOI21_X1 U16363 ( .B1(n13135), .B2(n13134), .A(n13265), .ZN(n19798) );
  INV_X1 U16364 ( .A(n19798), .ZN(n13140) );
  INV_X1 U16365 ( .A(DATAI_8_), .ZN(n13137) );
  NAND2_X1 U16366 ( .A1(n20006), .A2(BUF1_REG_8__SCAN_IN), .ZN(n13136) );
  OAI21_X1 U16367 ( .B1(n20006), .B2(n13137), .A(n13136), .ZN(n19907) );
  INV_X1 U16368 ( .A(n19907), .ZN(n13139) );
  OAI222_X1 U16369 ( .A1(n13140), .A2(n14197), .B1(n14193), .B2(n13139), .C1(
        n13138), .C2(n14191), .ZN(P1_U2896) );
  INV_X1 U16370 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n19792) );
  NAND2_X1 U16371 ( .A1(n19798), .A2(n19876), .ZN(n13148) );
  NAND2_X1 U16372 ( .A1(n13940), .A2(n19792), .ZN(n13143) );
  NAND2_X1 U16373 ( .A1(n9724), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13141) );
  OAI211_X1 U16374 ( .C1(n13950), .C2(P1_EBX_REG_8__SCAN_IN), .A(n13944), .B(
        n13141), .ZN(n13142) );
  NAND2_X1 U16375 ( .A1(n13143), .A2(n13142), .ZN(n13144) );
  AND2_X1 U16376 ( .A1(n13145), .A2(n13144), .ZN(n13146) );
  NOR2_X1 U16377 ( .A1(n9847), .A2(n13146), .ZN(n19795) );
  NAND2_X1 U16378 ( .A1(n19795), .A2(n19875), .ZN(n13147) );
  OAI211_X1 U16379 ( .C1(n19792), .C2(n19879), .A(n13148), .B(n13147), .ZN(
        P1_U2864) );
  AOI22_X1 U16380 ( .A1(n19935), .A2(P1_EAX_REG_21__SCAN_IN), .B1(
        P1_UWORD_REG_5__SCAN_IN), .B2(n19912), .ZN(n13152) );
  NAND2_X1 U16381 ( .A1(n13152), .A2(n13151), .ZN(P1_U2942) );
  AOI22_X1 U16382 ( .A1(n19935), .A2(P1_EAX_REG_0__SCAN_IN), .B1(
        P1_LWORD_REG_0__SCAN_IN), .B2(n19932), .ZN(n13154) );
  INV_X1 U16383 ( .A(n20017), .ZN(n13153) );
  NAND2_X1 U16384 ( .A1(n19920), .A2(n13153), .ZN(n13163) );
  NAND2_X1 U16385 ( .A1(n13154), .A2(n13163), .ZN(P1_U2952) );
  AOI22_X1 U16386 ( .A1(n19935), .A2(P1_EAX_REG_19__SCAN_IN), .B1(
        P1_UWORD_REG_3__SCAN_IN), .B2(n19912), .ZN(n13156) );
  NAND2_X1 U16387 ( .A1(n13156), .A2(n13155), .ZN(P1_U2940) );
  AOI22_X1 U16388 ( .A1(n19935), .A2(P1_EAX_REG_22__SCAN_IN), .B1(
        P1_UWORD_REG_6__SCAN_IN), .B2(n19912), .ZN(n13158) );
  NAND2_X1 U16389 ( .A1(n13158), .A2(n13157), .ZN(P1_U2943) );
  AOI22_X1 U16390 ( .A1(n19935), .A2(P1_EAX_REG_23__SCAN_IN), .B1(
        P1_UWORD_REG_7__SCAN_IN), .B2(n19932), .ZN(n13160) );
  NAND2_X1 U16391 ( .A1(n13160), .A2(n13159), .ZN(P1_U2944) );
  AOI22_X1 U16392 ( .A1(n19935), .A2(P1_EAX_REG_18__SCAN_IN), .B1(
        P1_UWORD_REG_2__SCAN_IN), .B2(n19932), .ZN(n13162) );
  NAND2_X1 U16393 ( .A1(n13162), .A2(n13161), .ZN(P1_U2939) );
  AOI22_X1 U16394 ( .A1(n19935), .A2(P1_EAX_REG_16__SCAN_IN), .B1(
        P1_UWORD_REG_0__SCAN_IN), .B2(n19932), .ZN(n13164) );
  NAND2_X1 U16395 ( .A1(n13164), .A2(n13163), .ZN(P1_U2937) );
  AOI22_X1 U16396 ( .A1(n19935), .A2(P1_EAX_REG_17__SCAN_IN), .B1(
        P1_UWORD_REG_1__SCAN_IN), .B2(n19932), .ZN(n13165) );
  INV_X1 U16397 ( .A(n20023), .ZN(n14180) );
  NAND2_X1 U16398 ( .A1(n19920), .A2(n14180), .ZN(n13166) );
  NAND2_X1 U16399 ( .A1(n13165), .A2(n13166), .ZN(P1_U2938) );
  AOI22_X1 U16400 ( .A1(n19935), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_LWORD_REG_1__SCAN_IN), .B2(n19932), .ZN(n13167) );
  NAND2_X1 U16401 ( .A1(n13167), .A2(n13166), .ZN(P1_U2953) );
  AOI22_X1 U16402 ( .A1(n19935), .A2(P1_EAX_REG_20__SCAN_IN), .B1(
        P1_UWORD_REG_4__SCAN_IN), .B2(n19932), .ZN(n13169) );
  NAND2_X1 U16403 ( .A1(n13169), .A2(n13168), .ZN(P1_U2941) );
  AOI22_X1 U16404 ( .A1(n19935), .A2(P1_EAX_REG_26__SCAN_IN), .B1(
        P1_UWORD_REG_10__SCAN_IN), .B2(n19932), .ZN(n13172) );
  INV_X1 U16405 ( .A(DATAI_10_), .ZN(n13171) );
  NAND2_X1 U16406 ( .A1(n20006), .A2(BUF1_REG_10__SCAN_IN), .ZN(n13170) );
  OAI21_X1 U16407 ( .B1(n20006), .B2(n13171), .A(n13170), .ZN(n14140) );
  NAND2_X1 U16408 ( .A1(n19920), .A2(n14140), .ZN(n19926) );
  NAND2_X1 U16409 ( .A1(n13172), .A2(n19926), .ZN(P1_U2947) );
  NOR2_X1 U16410 ( .A1(n18923), .A2(n13173), .ZN(n13177) );
  OAI22_X1 U16411 ( .A1(n18848), .A2(n13175), .B1(n13174), .B2(n18911), .ZN(
        n13176) );
  AOI211_X1 U16412 ( .C1(P2_EBX_REG_1__SCAN_IN), .C2(n18919), .A(n13177), .B(
        n13176), .ZN(n13179) );
  NAND2_X1 U16413 ( .A1(n19712), .A2(n18917), .ZN(n13178) );
  OAI211_X1 U16414 ( .C1(n11154), .C2(n18894), .A(n13179), .B(n13178), .ZN(
        n13183) );
  OAI21_X1 U16415 ( .B1(n13194), .B2(n13181), .A(n13180), .ZN(n13193) );
  AOI221_X1 U16416 ( .B1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n13193), .C1(
        n12951), .C2(n13193), .A(n19614), .ZN(n13182) );
  AOI211_X1 U16417 ( .C1(n19710), .C2(n18913), .A(n13183), .B(n13182), .ZN(
        n13184) );
  INV_X1 U16418 ( .A(n13184), .ZN(P2_U2854) );
  INV_X1 U16419 ( .A(n13185), .ZN(n13186) );
  INV_X1 U16420 ( .A(n11447), .ZN(n15090) );
  NAND3_X1 U16421 ( .A1(n15091), .A2(n13186), .A3(n15090), .ZN(n13192) );
  OR2_X1 U16422 ( .A1(n16169), .A2(n13187), .ZN(n15089) );
  NOR2_X1 U16423 ( .A1(n10507), .A2(n16164), .ZN(n15094) );
  NOR2_X1 U16424 ( .A1(n15094), .A2(n9743), .ZN(n13190) );
  NAND3_X1 U16425 ( .A1(n15093), .A2(n15092), .A3(n13190), .ZN(n13189) );
  OAI21_X1 U16426 ( .B1(n15089), .B2(n13190), .A(n13189), .ZN(n13191) );
  OAI211_X1 U16427 ( .C1(n11148), .C2(n15072), .A(n13192), .B(n13191), .ZN(
        n16183) );
  OAI21_X1 U16428 ( .B1(n18863), .B2(n9972), .A(n13193), .ZN(n15085) );
  OAI22_X1 U16429 ( .A1(n18863), .A2(n13195), .B1(n13194), .B2(n18903), .ZN(
        n15076) );
  INV_X1 U16430 ( .A(n15076), .ZN(n13197) );
  NOR2_X1 U16431 ( .A1(n13197), .A2(n13196), .ZN(n15079) );
  AOI222_X1 U16432 ( .A1(n16183), .A2(n19606), .B1(n16199), .B2(n13215), .C1(
        n15085), .C2(n15079), .ZN(n13200) );
  NAND2_X1 U16433 ( .A1(n13199), .A2(n16164), .ZN(n13198) );
  OAI21_X1 U16434 ( .B1(n13200), .B2(n13199), .A(n13198), .ZN(P2_U3599) );
  NOR2_X2 U16435 ( .A1(n13201), .A2(n19426), .ZN(n19597) );
  INV_X1 U16436 ( .A(n19597), .ZN(n19507) );
  INV_X1 U16437 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n16291) );
  INV_X1 U16438 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n18058) );
  INV_X1 U16439 ( .A(n19599), .ZN(n19514) );
  AOI22_X1 U16440 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n19090), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n19089), .ZN(n19605) );
  INV_X1 U16441 ( .A(n19605), .ZN(n19536) );
  AND2_X1 U16442 ( .A1(n10390), .A2(n19076), .ZN(n19596) );
  AOI22_X1 U16443 ( .A1(n19536), .A2(n19131), .B1(n19086), .B2(n19596), .ZN(
        n13202) );
  OAI21_X1 U16444 ( .B1(n19514), .B2(n19604), .A(n13202), .ZN(n13203) );
  AOI21_X1 U16445 ( .B1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B2(n13211), .A(
        n13203), .ZN(n13204) );
  OAI21_X1 U16446 ( .B1(n13213), .B2(n19507), .A(n13204), .ZN(P2_U3055) );
  INV_X1 U16447 ( .A(n19584), .ZN(n19494) );
  INV_X1 U16448 ( .A(n19529), .ZN(n19588) );
  INV_X1 U16449 ( .A(n19131), .ZN(n13209) );
  INV_X1 U16450 ( .A(n19604), .ZN(n19087) );
  AOI22_X1 U16451 ( .A1(n19585), .A2(n19087), .B1(n19583), .B2(n19086), .ZN(
        n13205) );
  OAI21_X1 U16452 ( .B1(n19588), .B2(n13209), .A(n13205), .ZN(n13206) );
  AOI21_X1 U16453 ( .B1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B2(n13211), .A(
        n13206), .ZN(n13207) );
  OAI21_X1 U16454 ( .B1(n13213), .B2(n19494), .A(n13207), .ZN(P2_U3053) );
  INV_X1 U16455 ( .A(n12991), .ZN(n19457) );
  INV_X1 U16456 ( .A(n19465), .ZN(n19558) );
  AOI22_X1 U16457 ( .A1(n19555), .A2(n19087), .B1(n19547), .B2(n19086), .ZN(
        n13208) );
  OAI21_X1 U16458 ( .B1(n19558), .B2(n13209), .A(n13208), .ZN(n13210) );
  AOI21_X1 U16459 ( .B1(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B2(n13211), .A(
        n13210), .ZN(n13212) );
  OAI21_X1 U16460 ( .B1(n13213), .B2(n19457), .A(n13212), .ZN(P2_U3048) );
  NAND2_X1 U16461 ( .A1(n13215), .A2(n19707), .ZN(n19423) );
  NOR3_X1 U16462 ( .A1(n19600), .A2(n19537), .A3(n19337), .ZN(n13216) );
  NOR2_X1 U16463 ( .A1(n13216), .A2(n19303), .ZN(n13218) );
  NOR3_X2 U16464 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19697), .A3(
        n19544), .ZN(n19535) );
  NAND3_X1 U16465 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n10862), .ZN(n19461) );
  NOR2_X1 U16466 ( .A1(n19722), .A2(n19461), .ZN(n19464) );
  NOR2_X1 U16467 ( .A1(n19535), .A2(n19464), .ZN(n13221) );
  INV_X1 U16468 ( .A(n11199), .ZN(n13219) );
  OAI21_X1 U16469 ( .B1(n13219), .B2(n19535), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n13217) );
  OAI21_X1 U16470 ( .B1(n13218), .B2(n13221), .A(n13217), .ZN(n19538) );
  INV_X1 U16471 ( .A(n19538), .ZN(n13228) );
  INV_X1 U16472 ( .A(n13218), .ZN(n13222) );
  AOI211_X1 U16473 ( .C1(n13219), .C2(n19714), .A(n19685), .B(n19535), .ZN(
        n13220) );
  AOI211_X2 U16474 ( .C1(n13222), .C2(n13221), .A(n13220), .B(n19426), .ZN(
        n19542) );
  INV_X1 U16475 ( .A(n19542), .ZN(n13226) );
  AOI22_X1 U16476 ( .A1(n19555), .A2(n19537), .B1(n19547), .B2(n19535), .ZN(
        n13223) );
  OAI21_X1 U16477 ( .B1(n19558), .B2(n13224), .A(n13223), .ZN(n13225) );
  AOI21_X1 U16478 ( .B1(n13226), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .A(
        n13225), .ZN(n13227) );
  OAI21_X1 U16479 ( .B1(n13228), .B2(n19457), .A(n13227), .ZN(P2_U3160) );
  NAND2_X1 U16480 ( .A1(n13229), .A2(n14601), .ZN(n13233) );
  AND2_X1 U16481 ( .A1(n9842), .A2(n13230), .ZN(n13231) );
  OR2_X1 U16482 ( .A1(n13231), .A2(n13297), .ZN(n15006) );
  NAND2_X1 U16483 ( .A1(n18761), .A2(n14621), .ZN(n13232) );
  OAI211_X1 U16484 ( .C1(n14621), .C2(n11351), .A(n13233), .B(n13232), .ZN(
        P2_U2871) );
  NAND2_X1 U16485 ( .A1(n13234), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13235) );
  OR2_X1 U16486 ( .A1(n12864), .A2(n13345), .ZN(n13243) );
  NAND2_X1 U16487 ( .A1(n13239), .A2(n13238), .ZN(n13354) );
  INV_X1 U16488 ( .A(n13352), .ZN(n13240) );
  XNOR2_X1 U16489 ( .A(n13354), .B(n13240), .ZN(n13241) );
  NAND2_X1 U16490 ( .A1(n13241), .A2(n13383), .ZN(n13242) );
  NAND2_X1 U16491 ( .A1(n13243), .A2(n13242), .ZN(n13244) );
  OAI21_X1 U16492 ( .B1(n13245), .B2(n13244), .A(n13341), .ZN(n19955) );
  AOI22_X1 U16493 ( .A1(n19938), .A2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B1(
        n13009), .B2(P1_REIP_REG_3__SCAN_IN), .ZN(n13246) );
  OAI21_X1 U16494 ( .B1(n15701), .B2(n13247), .A(n13246), .ZN(n13248) );
  AOI21_X1 U16495 ( .B1(n13249), .B2(n9727), .A(n13248), .ZN(n13250) );
  OAI21_X1 U16496 ( .B1(n19955), .B2(n19764), .A(n13250), .ZN(P1_U2996) );
  XNOR2_X1 U16497 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B(n13251), .ZN(
        n19787) );
  AOI22_X1 U16498 ( .A1(n12709), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n9755), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n13255) );
  AOI22_X1 U16499 ( .A1(n12619), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12367), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n13254) );
  AOI22_X1 U16500 ( .A1(n13867), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n13848), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n13253) );
  NAND4_X1 U16501 ( .A1(n13255), .A2(n13254), .A3(n13253), .A4(n13252), .ZN(
        n13261) );
  AOI22_X1 U16502 ( .A1(n13803), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n9732), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n13259) );
  AOI22_X1 U16503 ( .A1(n13707), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n13825), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n13258) );
  AOI22_X1 U16504 ( .A1(n13868), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n9722), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n13257) );
  AOI22_X1 U16505 ( .A1(n9738), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n13769), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n13256) );
  NAND4_X1 U16506 ( .A1(n13259), .A2(n13258), .A3(n13257), .A4(n13256), .ZN(
        n13260) );
  OR2_X1 U16507 ( .A1(n13261), .A2(n13260), .ZN(n13262) );
  AOI22_X1 U16508 ( .A1(n13505), .A2(n13262), .B1(n13887), .B2(
        P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n13264) );
  NAND2_X1 U16509 ( .A1(n13888), .A2(P1_EAX_REG_9__SCAN_IN), .ZN(n13263) );
  OAI211_X1 U16510 ( .C1(n19787), .C2(n13886), .A(n13264), .B(n13263), .ZN(
        n13266) );
  NOR2_X1 U16511 ( .A1(n13265), .A2(n13266), .ZN(n13267) );
  OR2_X1 U16512 ( .A1(n13320), .A2(n13267), .ZN(n19786) );
  INV_X1 U16513 ( .A(DATAI_9_), .ZN(n13269) );
  NAND2_X1 U16514 ( .A1(n20006), .A2(BUF1_REG_9__SCAN_IN), .ZN(n13268) );
  OAI21_X1 U16515 ( .B1(n20006), .B2(n13269), .A(n13268), .ZN(n19910) );
  AOI22_X1 U16516 ( .A1(n14195), .A2(n19910), .B1(P1_EAX_REG_9__SCAN_IN), .B2(
        n14194), .ZN(n13270) );
  OAI21_X1 U16517 ( .B1(n19786), .B2(n14197), .A(n13270), .ZN(P1_U2895) );
  XNOR2_X1 U16518 ( .A(n13271), .B(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n16040) );
  XNOR2_X1 U16519 ( .A(n13272), .B(n13273), .ZN(n16039) );
  INV_X1 U16520 ( .A(n15065), .ZN(n15053) );
  NOR2_X1 U16521 ( .A1(n11564), .A2(n18846), .ZN(n13274) );
  AOI221_X1 U16522 ( .B1(n13275), .B2(n20739), .C1(n15053), .C2(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(n13274), .ZN(n13278) );
  INV_X1 U16523 ( .A(n18881), .ZN(n13276) );
  AOI22_X1 U16524 ( .A1(n18877), .A2(n16154), .B1(n19059), .B2(n13276), .ZN(
        n13277) );
  OAI211_X1 U16525 ( .C1(n16039), .C2(n16139), .A(n13278), .B(n13277), .ZN(
        n13279) );
  INV_X1 U16526 ( .A(n13279), .ZN(n13280) );
  OAI21_X1 U16527 ( .B1(n16040), .B2(n19056), .A(n13280), .ZN(P2_U3040) );
  INV_X1 U16528 ( .A(P1_EBX_REG_9__SCAN_IN), .ZN(n13287) );
  NAND2_X1 U16529 ( .A1(n13931), .A2(n13287), .ZN(n13284) );
  NAND2_X1 U16530 ( .A1(n9724), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n13281) );
  NAND2_X1 U16531 ( .A1(n13944), .A2(n13281), .ZN(n13282) );
  OAI21_X1 U16532 ( .B1(n13950), .B2(P1_EBX_REG_9__SCAN_IN), .A(n13282), .ZN(
        n13283) );
  NAND2_X1 U16533 ( .A1(n13284), .A2(n13283), .ZN(n13286) );
  INV_X1 U16534 ( .A(n13327), .ZN(n13285) );
  OAI21_X1 U16535 ( .B1(n9847), .B2(n13286), .A(n13285), .ZN(n19784) );
  OAI222_X1 U16536 ( .A1(n19786), .A2(n15631), .B1(n19879), .B2(n13287), .C1(
        n14120), .C2(n19784), .ZN(P1_U2863) );
  OAI21_X1 U16537 ( .B1(n13289), .B2(n13288), .A(n10186), .ZN(n13301) );
  AOI21_X1 U16538 ( .B1(n13291), .B2(n13290), .A(n13332), .ZN(n18749) );
  INV_X1 U16539 ( .A(n18749), .ZN(n13292) );
  INV_X1 U16540 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n18985) );
  OAI22_X1 U16541 ( .A1(n14709), .A2(n13292), .B1(n18985), .B2(n18948), .ZN(
        n13293) );
  AOI21_X1 U16542 ( .B1(n15927), .B2(n13294), .A(n13293), .ZN(n13296) );
  AOI22_X1 U16543 ( .A1(n18929), .A2(BUF2_REG_17__SCAN_IN), .B1(n18931), .B2(
        BUF1_REG_17__SCAN_IN), .ZN(n13295) );
  OAI211_X1 U16544 ( .C1(n13301), .C2(n14714), .A(n13296), .B(n13295), .ZN(
        P2_U2902) );
  XOR2_X1 U16545 ( .A(n13298), .B(n13297), .Z(n18748) );
  NAND2_X1 U16546 ( .A1(n18748), .A2(n14582), .ZN(n13300) );
  NAND2_X1 U16547 ( .A1(n14602), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n13299) );
  OAI211_X1 U16548 ( .C1(n13301), .C2(n14630), .A(n13300), .B(n13299), .ZN(
        P2_U2870) );
  XNOR2_X1 U16549 ( .A(n13302), .B(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n15623) );
  NAND2_X1 U16550 ( .A1(n15623), .A2(n13880), .ZN(n13318) );
  AOI22_X1 U16551 ( .A1(n13707), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n12709), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n13306) );
  AOI22_X1 U16552 ( .A1(n9741), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n13803), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n13305) );
  AOI22_X1 U16553 ( .A1(n13464), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12367), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n13304) );
  AOI22_X1 U16554 ( .A1(n13867), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n9722), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n13303) );
  NAND4_X1 U16555 ( .A1(n13306), .A2(n13305), .A3(n13304), .A4(n13303), .ZN(
        n13312) );
  AOI22_X1 U16556 ( .A1(n12619), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n9757), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n13310) );
  AOI22_X1 U16557 ( .A1(n13868), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n13848), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n13309) );
  AOI22_X1 U16558 ( .A1(n9732), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n13825), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n13308) );
  NAND4_X1 U16559 ( .A1(n13310), .A2(n13309), .A3(n13308), .A4(n13307), .ZN(
        n13311) );
  NOR2_X1 U16560 ( .A1(n13312), .A2(n13311), .ZN(n13315) );
  NAND2_X1 U16561 ( .A1(n13888), .A2(P1_EAX_REG_10__SCAN_IN), .ZN(n13314) );
  NAND2_X1 U16562 ( .A1(n13887), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n13313) );
  OAI211_X1 U16563 ( .C1(n13586), .C2(n13315), .A(n13314), .B(n13313), .ZN(
        n13316) );
  INV_X1 U16564 ( .A(n13316), .ZN(n13317) );
  NAND2_X1 U16565 ( .A1(n13318), .A2(n13317), .ZN(n13319) );
  INV_X1 U16566 ( .A(n13319), .ZN(n13322) );
  INV_X1 U16567 ( .A(n13320), .ZN(n13321) );
  INV_X1 U16568 ( .A(n13458), .ZN(n13512) );
  AOI21_X1 U16569 ( .B1(n13322), .B2(n13321), .A(n13512), .ZN(n15625) );
  INV_X1 U16570 ( .A(n15625), .ZN(n13329) );
  AOI22_X1 U16571 ( .A1(n14195), .A2(n14140), .B1(P1_EAX_REG_10__SCAN_IN), 
        .B2(n14194), .ZN(n13323) );
  OAI21_X1 U16572 ( .B1(n13329), .B2(n14197), .A(n13323), .ZN(P1_U2894) );
  INV_X1 U16573 ( .A(P1_EBX_REG_10__SCAN_IN), .ZN(n13328) );
  MUX2_X1 U16574 ( .A(n13940), .B(n13971), .S(P1_EBX_REG_10__SCAN_IN), .Z(
        n13325) );
  NOR2_X1 U16575 ( .A1(n13951), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n13324) );
  NOR2_X1 U16576 ( .A1(n13325), .A2(n13324), .ZN(n13326) );
  OAI21_X1 U16577 ( .B1(n13327), .B2(n13326), .A(n13536), .ZN(n15620) );
  OAI222_X1 U16578 ( .A1(n13329), .A2(n15631), .B1(n19879), .B2(n13328), .C1(
        n14120), .C2(n15620), .ZN(P1_U2862) );
  OAI21_X1 U16579 ( .B1(n13331), .B2(n13330), .A(n13391), .ZN(n14629) );
  OR2_X1 U16580 ( .A1(n13333), .A2(n13332), .ZN(n13334) );
  NAND2_X1 U16581 ( .A1(n13334), .A2(n14707), .ZN(n18740) );
  INV_X1 U16582 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n18983) );
  OAI22_X1 U16583 ( .A1(n14709), .A2(n18740), .B1(n18983), .B2(n18948), .ZN(
        n13335) );
  AOI21_X1 U16584 ( .B1(n15927), .B2(n13336), .A(n13335), .ZN(n13338) );
  AOI22_X1 U16585 ( .A1(n18929), .A2(BUF2_REG_18__SCAN_IN), .B1(n18931), .B2(
        BUF1_REG_18__SCAN_IN), .ZN(n13337) );
  OAI211_X1 U16586 ( .C1(n14629), .C2(n14714), .A(n13338), .B(n13337), .ZN(
        P2_U2901) );
  NAND2_X1 U16587 ( .A1(n13339), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13340) );
  NAND2_X1 U16588 ( .A1(n13341), .A2(n13340), .ZN(n19941) );
  NAND2_X1 U16589 ( .A1(n13354), .A2(n13352), .ZN(n13342) );
  XNOR2_X1 U16590 ( .A(n13342), .B(n13351), .ZN(n13343) );
  NAND2_X1 U16591 ( .A1(n13343), .A2(n13383), .ZN(n13344) );
  OAI21_X1 U16592 ( .B1(n13346), .B2(n13345), .A(n13344), .ZN(n13348) );
  INV_X1 U16593 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n13347) );
  XNOR2_X1 U16594 ( .A(n13348), .B(n13347), .ZN(n19940) );
  NAND2_X1 U16595 ( .A1(n19941), .A2(n19940), .ZN(n19939) );
  NAND2_X1 U16596 ( .A1(n13348), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13349) );
  NAND2_X1 U16597 ( .A1(n19939), .A2(n13349), .ZN(n15697) );
  NAND2_X1 U16598 ( .A1(n13350), .A2(n13377), .ZN(n13357) );
  AND2_X1 U16599 ( .A1(n13352), .A2(n13351), .ZN(n13353) );
  NAND2_X1 U16600 ( .A1(n13354), .A2(n13353), .ZN(n13361) );
  XNOR2_X1 U16601 ( .A(n13361), .B(n13362), .ZN(n13355) );
  NAND2_X1 U16602 ( .A1(n13355), .A2(n13383), .ZN(n13356) );
  NAND2_X1 U16603 ( .A1(n13357), .A2(n13356), .ZN(n13358) );
  INV_X1 U16604 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n15801) );
  XNOR2_X1 U16605 ( .A(n13358), .B(n15801), .ZN(n15696) );
  NAND2_X1 U16606 ( .A1(n15697), .A2(n15696), .ZN(n15695) );
  NAND2_X1 U16607 ( .A1(n13358), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n13359) );
  NAND2_X1 U16608 ( .A1(n15695), .A2(n13359), .ZN(n15692) );
  NAND2_X1 U16609 ( .A1(n13360), .A2(n13377), .ZN(n13366) );
  INV_X1 U16610 ( .A(n13361), .ZN(n13363) );
  NAND2_X1 U16611 ( .A1(n13363), .A2(n13362), .ZN(n13370) );
  XNOR2_X1 U16612 ( .A(n13370), .B(n13371), .ZN(n13364) );
  NAND2_X1 U16613 ( .A1(n13364), .A2(n13383), .ZN(n13365) );
  NAND2_X1 U16614 ( .A1(n13366), .A2(n13365), .ZN(n15690) );
  OR2_X1 U16615 ( .A1(n15690), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13367) );
  NAND2_X1 U16616 ( .A1(n15690), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13368) );
  NAND2_X1 U16617 ( .A1(n13369), .A2(n13377), .ZN(n13375) );
  INV_X1 U16618 ( .A(n13370), .ZN(n13372) );
  NAND2_X1 U16619 ( .A1(n13372), .A2(n13371), .ZN(n13381) );
  XNOR2_X1 U16620 ( .A(n13381), .B(n13382), .ZN(n13373) );
  NAND2_X1 U16621 ( .A1(n13373), .A2(n13383), .ZN(n13374) );
  NAND2_X1 U16622 ( .A1(n13375), .A2(n13374), .ZN(n15685) );
  AND2_X1 U16623 ( .A1(n15685), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n13376) );
  AND2_X1 U16624 ( .A1(n13378), .A2(n13377), .ZN(n13379) );
  INV_X1 U16625 ( .A(n13381), .ZN(n13384) );
  NAND3_X1 U16626 ( .A1(n13384), .A2(n13383), .A3(n13382), .ZN(n13385) );
  NAND2_X1 U16627 ( .A1(n9750), .A2(n13385), .ZN(n13399) );
  XOR2_X1 U16628 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B(n13399), .Z(
        n13386) );
  XNOR2_X1 U16629 ( .A(n13398), .B(n13386), .ZN(n15777) );
  INV_X1 U16630 ( .A(n15777), .ZN(n13390) );
  AOI22_X1 U16631 ( .A1(n19938), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(
        n13009), .B2(P1_REIP_REG_8__SCAN_IN), .ZN(n13387) );
  OAI21_X1 U16632 ( .B1(n15701), .B2(n19796), .A(n13387), .ZN(n13388) );
  AOI21_X1 U16633 ( .B1(n19798), .B2(n9727), .A(n13388), .ZN(n13389) );
  OAI21_X1 U16634 ( .B1(n13390), .B2(n19764), .A(n13389), .ZN(P1_U2991) );
  INV_X1 U16635 ( .A(n13391), .ZN(n13392) );
  OAI21_X1 U16636 ( .B1(n13392), .B2(n9878), .A(n14613), .ZN(n14715) );
  OR2_X1 U16637 ( .A1(n14626), .A2(n13393), .ZN(n13395) );
  AND2_X1 U16638 ( .A1(n13395), .A2(n13394), .ZN(n18722) );
  NAND2_X1 U16639 ( .A1(n18722), .A2(n14582), .ZN(n13397) );
  NAND2_X1 U16640 ( .A1(n14602), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n13396) );
  OAI211_X1 U16641 ( .C1(n14715), .C2(n14630), .A(n13397), .B(n13396), .ZN(
        P2_U2868) );
  NAND2_X1 U16642 ( .A1(n13399), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13400) );
  NAND2_X1 U16643 ( .A1(n13401), .A2(n13400), .ZN(n14200) );
  INV_X1 U16644 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n13403) );
  NOR2_X1 U16645 ( .A1(n9750), .A2(n13403), .ZN(n14199) );
  NAND2_X1 U16646 ( .A1(n9750), .A2(n13403), .ZN(n14201) );
  INV_X1 U16647 ( .A(n14201), .ZN(n13404) );
  NOR2_X1 U16648 ( .A1(n14199), .A2(n13404), .ZN(n13405) );
  XNOR2_X1 U16649 ( .A(n14200), .B(n13405), .ZN(n13443) );
  AOI22_X1 U16650 ( .A1(n19938), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B1(
        n13009), .B2(P1_REIP_REG_9__SCAN_IN), .ZN(n13407) );
  INV_X1 U16651 ( .A(n15701), .ZN(n15672) );
  NAND2_X1 U16652 ( .A1(n15672), .A2(n19787), .ZN(n13406) );
  OAI211_X1 U16653 ( .C1(n19786), .C2(n20005), .A(n13407), .B(n13406), .ZN(
        n13408) );
  INV_X1 U16654 ( .A(n13408), .ZN(n13409) );
  OAI21_X1 U16655 ( .B1(n13443), .B2(n19764), .A(n13409), .ZN(P1_U2990) );
  NAND2_X1 U16656 ( .A1(n13438), .A2(n15490), .ZN(n13410) );
  NAND2_X1 U16657 ( .A1(n13410), .A2(n20666), .ZN(n13411) );
  OR2_X1 U16658 ( .A1(n13412), .A2(n13411), .ZN(n13417) );
  NAND2_X1 U16659 ( .A1(n9725), .A2(n13891), .ZN(n13413) );
  AOI21_X1 U16660 ( .B1(n13415), .B2(n13414), .A(n13413), .ZN(n13416) );
  NAND3_X1 U16661 ( .A1(n13420), .A2(n13419), .A3(n13418), .ZN(n13422) );
  OAI21_X1 U16662 ( .B1(n20034), .B2(n13436), .A(n13423), .ZN(n13424) );
  OR2_X1 U16663 ( .A1(n12425), .A2(n13424), .ZN(n13425) );
  AOI21_X1 U16664 ( .B1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n15797) );
  NAND2_X1 U16665 ( .A1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n19948) );
  NOR3_X1 U16666 ( .A1(n15797), .A2(n19948), .A3(n15801), .ZN(n14494) );
  NAND3_X1 U16667 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n14369) );
  MUX2_X1 U16668 ( .A(n13427), .B(n20026), .S(n9725), .Z(n13429) );
  NAND2_X1 U16669 ( .A1(n13429), .A2(n13428), .ZN(n13430) );
  OR2_X1 U16670 ( .A1(n13431), .A2(n13430), .ZN(n13432) );
  INV_X1 U16671 ( .A(n19963), .ZN(n14491) );
  NOR2_X1 U16672 ( .A1(n20722), .A2(n12449), .ZN(n13435) );
  INV_X1 U16673 ( .A(n19962), .ZN(n19984) );
  INV_X1 U16674 ( .A(n19985), .ZN(n19971) );
  NAND2_X1 U16675 ( .A1(n19971), .A2(n15797), .ZN(n19975) );
  OAI211_X1 U16676 ( .C1(n14491), .C2(n13435), .A(n19984), .B(n19975), .ZN(
        n19956) );
  NOR2_X1 U16677 ( .A1(n14369), .A2(n19956), .ZN(n13434) );
  NAND2_X1 U16678 ( .A1(n19985), .A2(n15472), .ZN(n19996) );
  INV_X1 U16679 ( .A(n15751), .ZN(n19998) );
  NOR2_X1 U16680 ( .A1(n19988), .A2(n19962), .ZN(n14373) );
  AOI21_X1 U16681 ( .B1(n14494), .B2(n13434), .A(n14373), .ZN(n15768) );
  INV_X1 U16682 ( .A(n13435), .ZN(n19969) );
  NAND2_X1 U16683 ( .A1(n19968), .A2(n15751), .ZN(n19987) );
  NAND2_X1 U16684 ( .A1(n19963), .A2(n19987), .ZN(n14496) );
  OAI21_X1 U16685 ( .B1(n19969), .B2(n14496), .A(n19985), .ZN(n15798) );
  NAND2_X1 U16686 ( .A1(n14494), .A2(n15798), .ZN(n15796) );
  NOR2_X1 U16687 ( .A1(n14369), .A2(n15796), .ZN(n15770) );
  INV_X1 U16688 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n20612) );
  OAI22_X1 U16689 ( .A1(n12340), .A2(n13438), .B1(n13437), .B2(n13436), .ZN(
        n13439) );
  OAI22_X1 U16690 ( .A1(n19845), .A2(n20612), .B1(n15807), .B2(n19784), .ZN(
        n13441) );
  AOI221_X1 U16691 ( .B1(n15768), .B2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .C1(
        n15770), .C2(n13403), .A(n13441), .ZN(n13442) );
  OAI21_X1 U16692 ( .B1(n13443), .B2(n19964), .A(n13442), .ZN(P1_U3022) );
  INV_X1 U16693 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n13543) );
  OAI21_X1 U16694 ( .B1(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n13444), .A(
        n13489), .ZN(n15684) );
  AOI22_X1 U16695 ( .A1(n13880), .A2(n15684), .B1(n13887), .B2(
        P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n13445) );
  OAI21_X1 U16696 ( .B1(n13753), .B2(n13543), .A(n13445), .ZN(n13511) );
  INV_X1 U16697 ( .A(n13511), .ZN(n13446) );
  AOI22_X1 U16698 ( .A1(n12709), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n13803), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n13450) );
  AOI22_X1 U16699 ( .A1(n9739), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12619), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n13449) );
  AOI22_X1 U16700 ( .A1(n12367), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n13848), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13448) );
  AOI22_X1 U16701 ( .A1(n13707), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n13825), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n13447) );
  NAND4_X1 U16702 ( .A1(n13450), .A2(n13449), .A3(n13448), .A4(n13447), .ZN(
        n13456) );
  AOI22_X1 U16703 ( .A1(n13464), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n13867), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n13454) );
  AOI22_X1 U16704 ( .A1(n9732), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n9757), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13453) );
  AOI22_X1 U16705 ( .A1(n13868), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n9722), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n13452) );
  NAND4_X1 U16706 ( .A1(n13454), .A2(n13453), .A3(n13452), .A4(n13451), .ZN(
        n13455) );
  OR2_X1 U16707 ( .A1(n13456), .A2(n13455), .ZN(n13457) );
  NAND2_X1 U16708 ( .A1(n13505), .A2(n13457), .ZN(n13534) );
  XNOR2_X1 U16709 ( .A(n13459), .B(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n14359) );
  NAND2_X1 U16710 ( .A1(n14359), .A2(n13880), .ZN(n13476) );
  AOI22_X1 U16711 ( .A1(n12709), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n13803), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n13463) );
  AOI22_X1 U16712 ( .A1(n9740), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12619), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n13462) );
  AOI22_X1 U16713 ( .A1(n12367), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n13769), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n13461) );
  NAND4_X1 U16714 ( .A1(n13463), .A2(n13462), .A3(n13461), .A4(n13460), .ZN(
        n13470) );
  AOI22_X1 U16715 ( .A1(n13464), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n13868), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n13468) );
  AOI22_X1 U16716 ( .A1(n9732), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n9756), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n13467) );
  AOI22_X1 U16717 ( .A1(n13848), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n9722), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n13466) );
  AOI22_X1 U16718 ( .A1(n13707), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n13825), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n13465) );
  NAND4_X1 U16719 ( .A1(n13468), .A2(n13467), .A3(n13466), .A4(n13465), .ZN(
        n13469) );
  NOR2_X1 U16720 ( .A1(n13470), .A2(n13469), .ZN(n13473) );
  NAND2_X1 U16721 ( .A1(n13888), .A2(P1_EAX_REG_13__SCAN_IN), .ZN(n13472) );
  NAND2_X1 U16722 ( .A1(n13887), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n13471) );
  OAI211_X1 U16723 ( .C1(n13586), .C2(n13473), .A(n13472), .B(n13471), .ZN(
        n13474) );
  INV_X1 U16724 ( .A(n13474), .ZN(n13475) );
  NAND2_X1 U16725 ( .A1(n13476), .A2(n13475), .ZN(n14054) );
  INV_X1 U16726 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n13518) );
  AOI22_X1 U16727 ( .A1(n13707), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n12709), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n13481) );
  AOI22_X1 U16728 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n13868), .B1(
        n13848), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n13480) );
  AOI22_X1 U16729 ( .A1(n12619), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n13769), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n13479) );
  NAND4_X1 U16730 ( .A1(n13481), .A2(n13480), .A3(n13479), .A4(n13478), .ZN(
        n13487) );
  AOI22_X1 U16731 ( .A1(n13803), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n9755), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n13485) );
  AOI22_X1 U16732 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n9741), .B1(
        n12367), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n13484) );
  AOI22_X1 U16733 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n13867), .B1(
        n9722), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n13483) );
  AOI22_X1 U16734 ( .A1(n9732), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n13825), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n13482) );
  NAND4_X1 U16735 ( .A1(n13485), .A2(n13484), .A3(n13483), .A4(n13482), .ZN(
        n13486) );
  OR2_X1 U16736 ( .A1(n13487), .A2(n13486), .ZN(n13488) );
  NAND2_X1 U16737 ( .A1(n13505), .A2(n13488), .ZN(n13492) );
  XNOR2_X1 U16738 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B(n13489), .ZN(
        n15671) );
  INV_X1 U16739 ( .A(n13887), .ZN(n13617) );
  OAI22_X1 U16740 ( .A1(n15671), .A2(n13886), .B1(n13617), .B2(n15605), .ZN(
        n13490) );
  INV_X1 U16741 ( .A(n13490), .ZN(n13491) );
  OAI211_X1 U16742 ( .C1(n13518), .C2(n13753), .A(n13492), .B(n13491), .ZN(
        n13514) );
  XOR2_X1 U16743 ( .A(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B(n13493), .Z(
        n15665) );
  AOI22_X1 U16744 ( .A1(n13707), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n12709), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n13497) );
  AOI22_X1 U16745 ( .A1(n12619), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n9757), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13496) );
  AOI22_X1 U16746 ( .A1(n13464), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12367), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n13495) );
  AOI22_X1 U16747 ( .A1(n13867), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n13848), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13494) );
  NAND4_X1 U16748 ( .A1(n13497), .A2(n13496), .A3(n13495), .A4(n13494), .ZN(
        n13503) );
  AOI22_X1 U16749 ( .A1(n9739), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n13803), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n13501) );
  AOI22_X1 U16750 ( .A1(n9732), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n13825), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n13500) );
  AOI22_X1 U16751 ( .A1(n13868), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n9722), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n13499) );
  NAND4_X1 U16752 ( .A1(n13501), .A2(n13500), .A3(n13499), .A4(n13498), .ZN(
        n13502) );
  OR2_X1 U16753 ( .A1(n13503), .A2(n13502), .ZN(n13504) );
  AOI22_X1 U16754 ( .A1(n13505), .A2(n13504), .B1(n13887), .B2(
        P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n13507) );
  NAND2_X1 U16755 ( .A1(n13888), .A2(P1_EAX_REG_14__SCAN_IN), .ZN(n13506) );
  OAI211_X1 U16756 ( .C1(n15665), .C2(n13886), .A(n13507), .B(n13506), .ZN(
        n13508) );
  OAI21_X1 U16757 ( .B1(n9799), .B2(n13508), .A(n13588), .ZN(n15596) );
  INV_X1 U16758 ( .A(DATAI_14_), .ZN(n20942) );
  NAND2_X1 U16759 ( .A1(n20006), .A2(BUF1_REG_14__SCAN_IN), .ZN(n13509) );
  OAI21_X1 U16760 ( .B1(n20006), .B2(n20942), .A(n13509), .ZN(n19919) );
  AOI22_X1 U16761 ( .A1(n14195), .A2(n19919), .B1(P1_EAX_REG_14__SCAN_IN), 
        .B2(n14194), .ZN(n13510) );
  OAI21_X1 U16762 ( .B1(n15596), .B2(n14197), .A(n13510), .ZN(P1_U2890) );
  OAI21_X1 U16763 ( .B1(n13512), .B2(n13511), .A(n13513), .ZN(n13533) );
  OAI21_X1 U16764 ( .B1(n13533), .B2(n13534), .A(n13513), .ZN(n13515) );
  NAND2_X1 U16765 ( .A1(n13515), .A2(n13514), .ZN(n14056) );
  OAI21_X1 U16766 ( .B1(n13515), .B2(n13514), .A(n14056), .ZN(n15607) );
  INV_X1 U16767 ( .A(DATAI_12_), .ZN(n13517) );
  NAND2_X1 U16768 ( .A1(n20006), .A2(BUF1_REG_12__SCAN_IN), .ZN(n13516) );
  OAI21_X1 U16769 ( .B1(n20006), .B2(n13517), .A(n13516), .ZN(n19915) );
  INV_X1 U16770 ( .A(n19915), .ZN(n13519) );
  OAI222_X1 U16771 ( .A1(n15607), .A2(n14197), .B1(n14193), .B2(n13519), .C1(
        n13518), .C2(n14191), .ZN(P1_U2892) );
  INV_X1 U16772 ( .A(P1_EBX_REG_14__SCAN_IN), .ZN(n13532) );
  INV_X1 U16773 ( .A(P1_EBX_REG_11__SCAN_IN), .ZN(n13538) );
  NAND2_X1 U16774 ( .A1(n13931), .A2(n13538), .ZN(n13522) );
  INV_X1 U16775 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n14210) );
  NAND2_X1 U16776 ( .A1(n13944), .A2(n14210), .ZN(n13520) );
  OAI211_X1 U16777 ( .C1(n13950), .C2(P1_EBX_REG_11__SCAN_IN), .A(n13520), .B(
        n9724), .ZN(n13521) );
  INV_X1 U16778 ( .A(P1_EBX_REG_12__SCAN_IN), .ZN(n15643) );
  NAND2_X1 U16779 ( .A1(n13940), .A2(n15643), .ZN(n13525) );
  NAND2_X1 U16780 ( .A1(n9724), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n13523) );
  OAI211_X1 U16781 ( .C1(n13950), .C2(P1_EBX_REG_12__SCAN_IN), .A(n13944), .B(
        n13523), .ZN(n13524) );
  NAND2_X1 U16782 ( .A1(n13525), .A2(n13524), .ZN(n14500) );
  INV_X1 U16783 ( .A(P1_EBX_REG_13__SCAN_IN), .ZN(n14123) );
  NAND2_X1 U16784 ( .A1(n13931), .A2(n14123), .ZN(n13528) );
  INV_X1 U16785 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n20819) );
  NAND2_X1 U16786 ( .A1(n13944), .A2(n20819), .ZN(n13526) );
  OAI211_X1 U16787 ( .C1(n13950), .C2(P1_EBX_REG_13__SCAN_IN), .A(n13526), .B(
        n9724), .ZN(n13527) );
  MUX2_X1 U16788 ( .A(n13940), .B(n13971), .S(P1_EBX_REG_14__SCAN_IN), .Z(
        n13530) );
  NOR2_X1 U16789 ( .A1(n13951), .A2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n13529) );
  NOR2_X1 U16790 ( .A1(n13530), .A2(n13529), .ZN(n13531) );
  OAI21_X1 U16791 ( .B1(n14058), .B2(n13531), .A(n14116), .ZN(n15594) );
  OAI222_X1 U16792 ( .A1(n15596), .A2(n15631), .B1(n19879), .B2(n13532), .C1(
        n15594), .C2(n14120), .ZN(P1_U2858) );
  XOR2_X1 U16793 ( .A(n13534), .B(n13533), .Z(n15681) );
  NAND2_X1 U16794 ( .A1(n13536), .A2(n13535), .ZN(n13537) );
  NAND2_X1 U16795 ( .A1(n14501), .A2(n13537), .ZN(n15766) );
  OAI22_X1 U16796 ( .A1(n15766), .A2(n14120), .B1(n13538), .B2(n19879), .ZN(
        n13539) );
  AOI21_X1 U16797 ( .B1(n15681), .B2(n19876), .A(n13539), .ZN(n13540) );
  INV_X1 U16798 ( .A(n13540), .ZN(P1_U2861) );
  INV_X1 U16799 ( .A(n15681), .ZN(n13545) );
  INV_X1 U16800 ( .A(DATAI_11_), .ZN(n13542) );
  NAND2_X1 U16801 ( .A1(n20006), .A2(BUF1_REG_11__SCAN_IN), .ZN(n13541) );
  OAI21_X1 U16802 ( .B1(n20006), .B2(n13542), .A(n13541), .ZN(n19913) );
  INV_X1 U16803 ( .A(n19913), .ZN(n13544) );
  OAI222_X1 U16804 ( .A1(n13545), .A2(n14197), .B1(n14193), .B2(n13544), .C1(
        n13543), .C2(n14191), .ZN(P1_U2893) );
  AOI22_X1 U16805 ( .A1(n15162), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n16991), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n13555) );
  AOI22_X1 U16806 ( .A1(n16992), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11806), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13554) );
  AOI22_X1 U16807 ( .A1(n9729), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n16954), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n13546) );
  OAI21_X1 U16808 ( .B1(n16767), .B2(n20836), .A(n13546), .ZN(n13552) );
  AOI22_X1 U16809 ( .A1(n16993), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n16986), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n13550) );
  AOI22_X1 U16810 ( .A1(n11754), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n16974), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n13549) );
  AOI22_X1 U16811 ( .A1(n17000), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n16968), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n13548) );
  AOI22_X1 U16812 ( .A1(n9726), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n16969), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n13547) );
  NAND4_X1 U16813 ( .A1(n13550), .A2(n13549), .A3(n13548), .A4(n13547), .ZN(
        n13551) );
  AOI211_X1 U16814 ( .C1(n16975), .C2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A(
        n13552), .B(n13551), .ZN(n13553) );
  NAND3_X1 U16815 ( .A1(n13555), .A2(n13554), .A3(n13553), .ZN(n17132) );
  INV_X1 U16816 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n15195) );
  AOI211_X1 U16817 ( .C1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .C2(n18630), .A(
        n13558), .B(n13557), .ZN(n15227) );
  INV_X1 U16818 ( .A(n15227), .ZN(n13561) );
  NOR2_X1 U16819 ( .A1(n15229), .A2(n18046), .ZN(n18454) );
  NOR2_X1 U16820 ( .A1(n13564), .A2(n18027), .ZN(n15234) );
  NAND3_X1 U16821 ( .A1(n15219), .A2(n18454), .A3(n15234), .ZN(n15217) );
  NAND2_X1 U16822 ( .A1(n18648), .A2(n18023), .ZN(n16208) );
  NAND2_X1 U16823 ( .A1(P3_EBX_REG_3__SCAN_IN), .A2(n17023), .ZN(n17019) );
  NAND2_X1 U16824 ( .A1(P3_EBX_REG_7__SCAN_IN), .A2(P3_EBX_REG_6__SCAN_IN), 
        .ZN(n17007) );
  INV_X1 U16825 ( .A(n17007), .ZN(n16985) );
  NOR2_X1 U16826 ( .A1(n18052), .A2(n15196), .ZN(n16901) );
  AOI21_X1 U16827 ( .B1(P3_EBX_REG_13__SCAN_IN), .B2(n16901), .A(
        P3_EBX_REG_14__SCAN_IN), .ZN(n13566) );
  NOR2_X1 U16828 ( .A1(n9763), .A2(n13566), .ZN(n13567) );
  INV_X2 U16829 ( .A(n17024), .ZN(n17039) );
  MUX2_X1 U16830 ( .A(n17132), .B(n13567), .S(n17039), .Z(P3_U2689) );
  NAND3_X1 U16831 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_0__SCAN_IN), .A3(P3_STATE2_REG_2__SCAN_IN), .ZN(n18598)
         );
  OAI21_X1 U16832 ( .B1(n13568), .B2(n18624), .A(n16695), .ZN(n15215) );
  NOR2_X1 U16833 ( .A1(n15318), .A2(n15215), .ZN(n18001) );
  INV_X1 U16834 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n16382) );
  NOR2_X1 U16835 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18658) );
  AOI21_X1 U16836 ( .B1(P3_STATE2_REG_2__SCAN_IN), .B2(
        P3_STATE2_REG_1__SCAN_IN), .A(n18658), .ZN(n18510) );
  NOR2_X1 U16837 ( .A1(n18626), .A2(n18510), .ZN(n18011) );
  OAI221_X1 U16838 ( .B1(n18598), .B2(n18001), .C1(n18598), .C2(n16382), .A(
        n18054), .ZN(n18008) );
  INV_X1 U16839 ( .A(n18008), .ZN(n18004) );
  INV_X1 U16840 ( .A(n18667), .ZN(n18602) );
  NAND2_X1 U16841 ( .A1(n18666), .A2(n18599), .ZN(n16377) );
  NAND2_X1 U16842 ( .A1(n18602), .A2(n16377), .ZN(n18002) );
  INV_X1 U16843 ( .A(n18002), .ZN(n18647) );
  NOR2_X1 U16844 ( .A1(n18610), .A2(n18653), .ZN(n17629) );
  NOR2_X1 U16845 ( .A1(n18647), .A2(n17629), .ZN(n15199) );
  AOI21_X1 U16846 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n15199), .ZN(n15200) );
  NOR2_X1 U16847 ( .A1(n18004), .A2(n15200), .ZN(n13570) );
  NOR3_X1 U16848 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .A3(n18653), .ZN(n18083) );
  INV_X1 U16849 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18309) );
  NAND2_X1 U16850 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n18309), .ZN(n18063) );
  NAND2_X1 U16851 ( .A1(n18063), .A2(n18008), .ZN(n15198) );
  OR2_X1 U16852 ( .A1(n18083), .A2(n15198), .ZN(n13569) );
  MUX2_X1 U16853 ( .A(n13570), .B(n13569), .S(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .Z(P3_U2864) );
  NOR2_X1 U16854 ( .A1(n13891), .A2(n20004), .ZN(n13571) );
  NAND2_X1 U16855 ( .A1(n14191), .A2(n13571), .ZN(n14184) );
  XNOR2_X1 U16856 ( .A(n13572), .B(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15592) );
  INV_X1 U16857 ( .A(n15592), .ZN(n14345) );
  AOI22_X1 U16858 ( .A1(n13707), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n9732), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n13576) );
  AOI22_X1 U16859 ( .A1(n13464), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n13867), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n13575) );
  AOI22_X1 U16860 ( .A1(n12619), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n9755), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n13574) );
  AOI22_X1 U16861 ( .A1(n13868), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n13848), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n13573) );
  NAND4_X1 U16862 ( .A1(n13576), .A2(n13575), .A3(n13574), .A4(n13573), .ZN(
        n13582) );
  AOI22_X1 U16863 ( .A1(n9739), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n13803), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n13580) );
  AOI22_X1 U16864 ( .A1(n12709), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n13825), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n13579) );
  AOI22_X1 U16865 ( .A1(n12367), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n13769), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n13578) );
  AOI22_X1 U16866 ( .A1(n9722), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n10197), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n13577) );
  NAND4_X1 U16867 ( .A1(n13580), .A2(n13579), .A3(n13578), .A4(n13577), .ZN(
        n13581) );
  NOR2_X1 U16868 ( .A1(n13582), .A2(n13581), .ZN(n13585) );
  NAND2_X1 U16869 ( .A1(n13888), .A2(P1_EAX_REG_15__SCAN_IN), .ZN(n13584) );
  NAND2_X1 U16870 ( .A1(n13887), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n13583) );
  OAI211_X1 U16871 ( .C1(n13586), .C2(n13585), .A(n13584), .B(n13583), .ZN(
        n13587) );
  AOI21_X1 U16872 ( .B1(n14345), .B2(n13880), .A(n13587), .ZN(n14114) );
  OR2_X1 U16873 ( .A1(n13589), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n13590) );
  NAND2_X1 U16874 ( .A1(n13590), .A2(n13616), .ZN(n15664) );
  AOI22_X1 U16875 ( .A1(n9738), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n13477), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n13594) );
  AOI22_X1 U16876 ( .A1(n13868), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n13867), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n13593) );
  AOI22_X1 U16877 ( .A1(n12126), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n13825), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n13592) );
  AOI22_X1 U16878 ( .A1(n13848), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n9721), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n13591) );
  NAND4_X1 U16879 ( .A1(n13594), .A2(n13593), .A3(n13592), .A4(n13591), .ZN(
        n13600) );
  AOI22_X1 U16880 ( .A1(n13707), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n12709), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n13598) );
  AOI22_X1 U16881 ( .A1(n9732), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n9757), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n13597) );
  AOI22_X1 U16882 ( .A1(n12374), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12367), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n13596) );
  AOI22_X1 U16883 ( .A1(n13769), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10197), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13595) );
  NAND4_X1 U16884 ( .A1(n13598), .A2(n13597), .A3(n13596), .A4(n13595), .ZN(
        n13599) );
  NOR2_X1 U16885 ( .A1(n13600), .A2(n13599), .ZN(n13601) );
  NOR2_X1 U16886 ( .A1(n13883), .A2(n13601), .ZN(n13604) );
  NAND2_X1 U16887 ( .A1(n12396), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n13602) );
  OAI211_X1 U16888 ( .C1(n13753), .C2(n12324), .A(n13886), .B(n13602), .ZN(
        n13603) );
  OAI22_X1 U16889 ( .A1(n15664), .A2(n13886), .B1(n13604), .B2(n13603), .ZN(
        n14107) );
  INV_X1 U16890 ( .A(n14107), .ZN(n13605) );
  AOI22_X1 U16891 ( .A1(n9732), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n9756), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n13609) );
  AOI22_X1 U16892 ( .A1(n9741), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12374), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n13608) );
  AOI22_X1 U16893 ( .A1(n13867), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n13848), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n13607) );
  AOI22_X1 U16894 ( .A1(n12709), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n13825), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n13606) );
  NAND4_X1 U16895 ( .A1(n13609), .A2(n13608), .A3(n13607), .A4(n13606), .ZN(
        n13615) );
  AOI22_X1 U16896 ( .A1(n13707), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n12619), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n13613) );
  AOI22_X1 U16897 ( .A1(n13868), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n9722), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n13612) );
  AOI22_X1 U16898 ( .A1(n12367), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n13769), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n13611) );
  AOI22_X1 U16899 ( .A1(n13464), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n10197), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n13610) );
  NAND4_X1 U16900 ( .A1(n13613), .A2(n13612), .A3(n13611), .A4(n13610), .ZN(
        n13614) );
  NOR2_X1 U16901 ( .A1(n13615), .A2(n13614), .ZN(n13620) );
  XNOR2_X1 U16902 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B(n13616), .ZN(
        n15570) );
  OAI22_X1 U16903 ( .A1(n15570), .A2(n13886), .B1(n13617), .B2(n15568), .ZN(
        n13618) );
  AOI21_X1 U16904 ( .B1(n13888), .B2(P1_EAX_REG_17__SCAN_IN), .A(n13618), .ZN(
        n13619) );
  OAI21_X1 U16905 ( .B1(n13883), .B2(n13620), .A(n13619), .ZN(n14098) );
  OR2_X1 U16906 ( .A1(n13621), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n13622) );
  NAND2_X1 U16907 ( .A1(n13622), .A2(n13685), .ZN(n15566) );
  INV_X1 U16908 ( .A(n15566), .ZN(n13637) );
  AOI22_X1 U16909 ( .A1(n13707), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n12709), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n13626) );
  AOI22_X1 U16910 ( .A1(n12126), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n9732), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n13625) );
  AOI22_X1 U16911 ( .A1(n13868), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n9722), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n13624) );
  AOI22_X1 U16912 ( .A1(n13464), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n10197), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n13623) );
  NAND4_X1 U16913 ( .A1(n13626), .A2(n13625), .A3(n13624), .A4(n13623), .ZN(
        n13632) );
  AOI22_X1 U16914 ( .A1(n9740), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n13803), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n13630) );
  AOI22_X1 U16915 ( .A1(n13867), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n13848), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13629) );
  AOI22_X1 U16916 ( .A1(n9756), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n13825), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n13628) );
  AOI22_X1 U16917 ( .A1(n12367), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n13769), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n13627) );
  NAND4_X1 U16918 ( .A1(n13630), .A2(n13629), .A3(n13628), .A4(n13627), .ZN(
        n13631) );
  OR2_X1 U16919 ( .A1(n13632), .A2(n13631), .ZN(n13635) );
  NAND2_X1 U16920 ( .A1(n12396), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n13633) );
  OAI211_X1 U16921 ( .C1(n13753), .C2(n20934), .A(n13886), .B(n13633), .ZN(
        n13634) );
  AOI21_X1 U16922 ( .B1(n13855), .B2(n13635), .A(n13634), .ZN(n13636) );
  AOI21_X1 U16923 ( .B1(n13637), .B2(n13880), .A(n13636), .ZN(n14091) );
  AOI22_X1 U16924 ( .A1(n12709), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12374), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n13641) );
  AOI22_X1 U16925 ( .A1(n13868), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n13867), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n13640) );
  AOI22_X1 U16926 ( .A1(n9739), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12367), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n13639) );
  AOI22_X1 U16927 ( .A1(n13769), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10197), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n13638) );
  NAND4_X1 U16928 ( .A1(n13641), .A2(n13640), .A3(n13639), .A4(n13638), .ZN(
        n13647) );
  AOI22_X1 U16929 ( .A1(n13464), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12619), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n13645) );
  AOI22_X1 U16930 ( .A1(n9732), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n9755), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13644) );
  AOI22_X1 U16931 ( .A1(n13848), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n9721), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n13643) );
  AOI22_X1 U16932 ( .A1(n13707), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n13825), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n13642) );
  NAND4_X1 U16933 ( .A1(n13645), .A2(n13644), .A3(n13643), .A4(n13642), .ZN(
        n13646) );
  NOR2_X1 U16934 ( .A1(n13647), .A2(n13646), .ZN(n13651) );
  NAND2_X1 U16935 ( .A1(n12396), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n13648) );
  OAI211_X1 U16936 ( .C1(n13753), .C2(n12591), .A(n13886), .B(n13648), .ZN(
        n13649) );
  INV_X1 U16937 ( .A(n13649), .ZN(n13650) );
  OAI21_X1 U16938 ( .B1(n13883), .B2(n13651), .A(n13650), .ZN(n13653) );
  XNOR2_X1 U16939 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B(n13655), .ZN(
        n14307) );
  NAND2_X1 U16940 ( .A1(n13880), .A2(n14307), .ZN(n13652) );
  NAND2_X1 U16941 ( .A1(n13653), .A2(n13652), .ZN(n14078) );
  OR2_X1 U16942 ( .A1(n13654), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n13656) );
  NAND2_X1 U16943 ( .A1(n13656), .A2(n13655), .ZN(n15655) );
  AOI22_X1 U16944 ( .A1(n12709), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n9732), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n13660) );
  AOI22_X1 U16945 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n13803), .B1(
        n9755), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n13659) );
  AOI22_X1 U16946 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n13867), .B1(
        n13848), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13658) );
  AOI22_X1 U16947 ( .A1(n13769), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n10197), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n13657) );
  NAND4_X1 U16948 ( .A1(n13660), .A2(n13659), .A3(n13658), .A4(n13657), .ZN(
        n13666) );
  AOI22_X1 U16949 ( .A1(n9739), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12126), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n13664) );
  AOI22_X1 U16950 ( .A1(n13464), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n12367), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n13663) );
  AOI22_X1 U16951 ( .A1(n13868), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n9722), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n13662) );
  AOI22_X1 U16952 ( .A1(n13707), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n13825), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n13661) );
  NAND4_X1 U16953 ( .A1(n13664), .A2(n13663), .A3(n13662), .A4(n13661), .ZN(
        n13665) );
  NOR2_X1 U16954 ( .A1(n13666), .A2(n13665), .ZN(n13667) );
  NOR2_X1 U16955 ( .A1(n13883), .A2(n13667), .ZN(n13670) );
  NAND2_X1 U16956 ( .A1(n12396), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n13668) );
  OAI211_X1 U16957 ( .C1(n13753), .C2(n12589), .A(n13886), .B(n13668), .ZN(
        n13669) );
  OAI22_X1 U16958 ( .A1(n15655), .A2(n13886), .B1(n13670), .B2(n13669), .ZN(
        n14166) );
  AOI22_X1 U16959 ( .A1(n13707), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n12709), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n13674) );
  AOI22_X1 U16960 ( .A1(n9732), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n9756), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n13673) );
  AOI22_X1 U16961 ( .A1(n9738), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12367), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n13672) );
  AOI22_X1 U16962 ( .A1(n13868), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n13848), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13671) );
  NAND4_X1 U16963 ( .A1(n13674), .A2(n13673), .A3(n13672), .A4(n13671), .ZN(
        n13680) );
  AOI22_X1 U16964 ( .A1(n13803), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n13825), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13678) );
  AOI22_X1 U16965 ( .A1(n13867), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n9722), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13677) );
  AOI22_X1 U16966 ( .A1(n12619), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n13769), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n13676) );
  AOI22_X1 U16967 ( .A1(n13464), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n10197), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n13675) );
  NAND4_X1 U16968 ( .A1(n13678), .A2(n13677), .A3(n13676), .A4(n13675), .ZN(
        n13679) );
  NOR2_X1 U16969 ( .A1(n13680), .A2(n13679), .ZN(n13684) );
  NAND2_X1 U16970 ( .A1(n12396), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n13681) );
  OAI211_X1 U16971 ( .C1(n13753), .C2(n12313), .A(n13886), .B(n13681), .ZN(
        n13682) );
  INV_X1 U16972 ( .A(n13682), .ZN(n13683) );
  OAI21_X1 U16973 ( .B1(n13883), .B2(n13684), .A(n13683), .ZN(n13687) );
  XNOR2_X1 U16974 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B(n13685), .ZN(
        n15556) );
  NAND2_X1 U16975 ( .A1(n15556), .A2(n13880), .ZN(n13686) );
  NAND2_X1 U16976 ( .A1(n13687), .A2(n13686), .ZN(n14086) );
  OR2_X1 U16977 ( .A1(n13689), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n13691) );
  NAND2_X1 U16978 ( .A1(n13691), .A2(n13690), .ZN(n15650) );
  INV_X1 U16979 ( .A(n15650), .ZN(n13706) );
  AOI22_X1 U16980 ( .A1(n13477), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n13867), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n13695) );
  AOI22_X1 U16981 ( .A1(n13707), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n9755), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n13694) );
  AOI22_X1 U16982 ( .A1(n13868), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n9721), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13693) );
  AOI22_X1 U16983 ( .A1(n12374), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n13769), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n13692) );
  NAND4_X1 U16984 ( .A1(n13695), .A2(n13694), .A3(n13693), .A4(n13692), .ZN(
        n13701) );
  AOI22_X1 U16985 ( .A1(n12126), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n9732), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n13699) );
  AOI22_X1 U16986 ( .A1(n9741), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12367), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n13698) );
  AOI22_X1 U16987 ( .A1(n12709), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n13825), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13697) );
  NAND4_X1 U16988 ( .A1(n13699), .A2(n13698), .A3(n13697), .A4(n13696), .ZN(
        n13700) );
  OR2_X1 U16989 ( .A1(n13701), .A2(n13700), .ZN(n13704) );
  NAND2_X1 U16990 ( .A1(n12396), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n13702) );
  OAI211_X1 U16991 ( .C1(n13753), .C2(n12585), .A(n13886), .B(n13702), .ZN(
        n13703) );
  AOI21_X1 U16992 ( .B1(n13855), .B2(n13704), .A(n13703), .ZN(n13705) );
  AOI21_X1 U16993 ( .B1(n13706), .B2(n13880), .A(n13705), .ZN(n14156) );
  AOI22_X1 U16994 ( .A1(n12709), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n9732), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n13711) );
  AOI22_X1 U16995 ( .A1(n9741), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12619), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n13710) );
  AOI22_X1 U16996 ( .A1(n13803), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n9757), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n13709) );
  AOI22_X1 U16997 ( .A1(n13707), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n13825), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n13708) );
  NAND4_X1 U16998 ( .A1(n13711), .A2(n13710), .A3(n13709), .A4(n13708), .ZN(
        n13717) );
  AOI22_X1 U16999 ( .A1(n13868), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n13867), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n13715) );
  AOI22_X1 U17000 ( .A1(n12367), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n13769), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n13714) );
  AOI22_X1 U17001 ( .A1(n13848), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n9722), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n13713) );
  AOI22_X1 U17002 ( .A1(n13464), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n10197), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n13712) );
  NAND4_X1 U17003 ( .A1(n13715), .A2(n13714), .A3(n13713), .A4(n13712), .ZN(
        n13716) );
  NOR2_X1 U17004 ( .A1(n13717), .A2(n13716), .ZN(n13740) );
  AOI22_X1 U17005 ( .A1(n13862), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n12709), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n13722) );
  AOI22_X1 U17006 ( .A1(n13803), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n9756), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n13721) );
  AOI22_X1 U17007 ( .A1(n13843), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n9722), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n13720) );
  AOI22_X1 U17008 ( .A1(n9740), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n13769), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n13719) );
  NAND4_X1 U17009 ( .A1(n13722), .A2(n13721), .A3(n13720), .A4(n13719), .ZN(
        n13728) );
  AOI22_X1 U17010 ( .A1(n12619), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12367), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n13726) );
  AOI22_X1 U17011 ( .A1(n13867), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n13848), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n13725) );
  AOI22_X1 U17012 ( .A1(n9732), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n13825), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n13724) );
  NAND4_X1 U17013 ( .A1(n13726), .A2(n13725), .A3(n13724), .A4(n13723), .ZN(
        n13727) );
  NOR2_X1 U17014 ( .A1(n13728), .A2(n13727), .ZN(n13739) );
  XOR2_X1 U17015 ( .A(n13740), .B(n13739), .Z(n13729) );
  NAND2_X1 U17016 ( .A1(n13729), .A2(n13855), .ZN(n13733) );
  OAI21_X1 U17017 ( .B1(n20439), .B2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n12396), .ZN(n13730) );
  OAI21_X1 U17018 ( .B1(n13753), .B2(n20835), .A(n13730), .ZN(n13731) );
  INV_X1 U17019 ( .A(n13731), .ZN(n13732) );
  NAND2_X1 U17020 ( .A1(n13733), .A2(n13732), .ZN(n13737) );
  NOR2_X1 U17021 ( .A1(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n13734), .ZN(
        n13735) );
  NOR2_X1 U17022 ( .A1(n13756), .A2(n13735), .ZN(n14050) );
  NAND2_X1 U17023 ( .A1(n14050), .A2(n13880), .ZN(n13736) );
  NAND2_X1 U17024 ( .A1(n13737), .A2(n13736), .ZN(n14046) );
  INV_X1 U17025 ( .A(n13738), .ZN(n14044) );
  NOR2_X1 U17026 ( .A1(n13740), .A2(n13739), .ZN(n13763) );
  AOI22_X1 U17027 ( .A1(n12709), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n9732), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n13744) );
  AOI22_X1 U17028 ( .A1(n9738), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12126), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n13743) );
  AOI22_X1 U17029 ( .A1(n13803), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n9757), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n13742) );
  AOI22_X1 U17030 ( .A1(n13862), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n13825), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n13741) );
  NAND4_X1 U17031 ( .A1(n13744), .A2(n13743), .A3(n13742), .A4(n13741), .ZN(
        n13750) );
  AOI22_X1 U17032 ( .A1(n13868), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n13867), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n13748) );
  AOI22_X1 U17033 ( .A1(n12367), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n13769), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n13747) );
  AOI22_X1 U17034 ( .A1(n13848), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n9722), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n13746) );
  NAND4_X1 U17035 ( .A1(n13748), .A2(n13747), .A3(n13746), .A4(n13745), .ZN(
        n13749) );
  OR2_X1 U17036 ( .A1(n13750), .A2(n13749), .ZN(n13762) );
  INV_X1 U17037 ( .A(n13762), .ZN(n13751) );
  XNOR2_X1 U17038 ( .A(n13763), .B(n13751), .ZN(n13755) );
  NAND2_X1 U17039 ( .A1(n12396), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n13752) );
  OAI211_X1 U17040 ( .C1(n13753), .C2(n12319), .A(n13886), .B(n13752), .ZN(
        n13754) );
  AOI21_X1 U17041 ( .B1(n13755), .B2(n13855), .A(n13754), .ZN(n13761) );
  INV_X1 U17042 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n13758) );
  INV_X1 U17043 ( .A(n13756), .ZN(n13757) );
  NAND2_X1 U17044 ( .A1(n13758), .A2(n13757), .ZN(n13759) );
  NAND2_X1 U17045 ( .A1(n13779), .A2(n13759), .ZN(n15520) );
  NOR2_X1 U17046 ( .A1(n15520), .A2(n13886), .ZN(n13760) );
  NAND2_X1 U17047 ( .A1(n13763), .A2(n13762), .ZN(n13785) );
  AOI22_X1 U17048 ( .A1(n13862), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n12709), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n13768) );
  AOI22_X1 U17049 ( .A1(n9740), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n13477), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n13767) );
  AOI22_X1 U17050 ( .A1(n13803), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12126), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n13766) );
  AOI22_X1 U17051 ( .A1(n13848), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n9722), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n13765) );
  NAND4_X1 U17052 ( .A1(n13768), .A2(n13767), .A3(n13766), .A4(n13765), .ZN(
        n13775) );
  AOI22_X1 U17053 ( .A1(n13868), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n13867), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n13773) );
  AOI22_X1 U17054 ( .A1(n9755), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12367), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n13772) );
  AOI22_X1 U17055 ( .A1(n9732), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n13825), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13771) );
  NAND4_X1 U17056 ( .A1(n13773), .A2(n13772), .A3(n13771), .A4(n13770), .ZN(
        n13774) );
  NOR2_X1 U17057 ( .A1(n13775), .A2(n13774), .ZN(n13786) );
  XOR2_X1 U17058 ( .A(n13785), .B(n13786), .Z(n13776) );
  NAND2_X1 U17059 ( .A1(n13776), .A2(n13855), .ZN(n13781) );
  NOR2_X1 U17060 ( .A1(n13777), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13778) );
  AOI211_X1 U17061 ( .C1(n13888), .C2(P1_EAX_REG_25__SCAN_IN), .A(n13880), .B(
        n13778), .ZN(n13780) );
  XNOR2_X1 U17062 ( .A(n13779), .B(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14283) );
  AOI22_X1 U17063 ( .A1(n13781), .A2(n13780), .B1(n13880), .B2(n14283), .ZN(
        n14032) );
  INV_X1 U17064 ( .A(n13782), .ZN(n13783) );
  INV_X1 U17065 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n14024) );
  NAND2_X1 U17066 ( .A1(n13783), .A2(n14024), .ZN(n13784) );
  NAND2_X1 U17067 ( .A1(n13817), .A2(n13784), .ZN(n14275) );
  NOR2_X1 U17068 ( .A1(n13786), .A2(n13785), .ZN(n13802) );
  AOI22_X1 U17069 ( .A1(n12709), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n9732), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n13790) );
  AOI22_X1 U17070 ( .A1(n9738), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12619), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n13789) );
  AOI22_X1 U17071 ( .A1(n12374), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n9757), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n13788) );
  AOI22_X1 U17072 ( .A1(n13862), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n13825), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13787) );
  NAND4_X1 U17073 ( .A1(n13790), .A2(n13789), .A3(n13788), .A4(n13787), .ZN(
        n13796) );
  AOI22_X1 U17074 ( .A1(n13843), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n13867), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n13794) );
  AOI22_X1 U17075 ( .A1(n12367), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n13769), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n13793) );
  AOI22_X1 U17076 ( .A1(n13848), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n9721), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n13792) );
  NAND4_X1 U17077 ( .A1(n13794), .A2(n13793), .A3(n13792), .A4(n13791), .ZN(
        n13795) );
  OR2_X1 U17078 ( .A1(n13796), .A2(n13795), .ZN(n13801) );
  XNOR2_X1 U17079 ( .A(n13802), .B(n13801), .ZN(n13799) );
  OAI21_X1 U17080 ( .B1(n20439), .B2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n12396), .ZN(n13798) );
  NAND2_X1 U17081 ( .A1(n13888), .A2(P1_EAX_REG_26__SCAN_IN), .ZN(n13797) );
  OAI211_X1 U17082 ( .C1(n13799), .C2(n13883), .A(n13798), .B(n13797), .ZN(
        n13800) );
  NAND2_X1 U17083 ( .A1(n13802), .A2(n13801), .ZN(n13823) );
  AOI22_X1 U17084 ( .A1(n13862), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n9732), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n13807) );
  AOI22_X1 U17085 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n13848), .B1(
        n9721), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n13806) );
  AOI22_X1 U17086 ( .A1(n13803), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n13769), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n13805) );
  NAND4_X1 U17087 ( .A1(n13807), .A2(n13806), .A3(n13805), .A4(n13804), .ZN(
        n13813) );
  AOI22_X1 U17088 ( .A1(n12619), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n9756), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n13811) );
  AOI22_X1 U17089 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n13464), .B1(
        n13867), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n13810) );
  AOI22_X1 U17090 ( .A1(n9740), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12367), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n13809) );
  AOI22_X1 U17091 ( .A1(n12709), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n13825), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13808) );
  NAND4_X1 U17092 ( .A1(n13811), .A2(n13810), .A3(n13809), .A4(n13808), .ZN(
        n13812) );
  NOR2_X1 U17093 ( .A1(n13813), .A2(n13812), .ZN(n13824) );
  XOR2_X1 U17094 ( .A(n13823), .B(n13824), .Z(n13814) );
  NAND2_X1 U17095 ( .A1(n13814), .A2(n13855), .ZN(n13819) );
  INV_X1 U17096 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n13815) );
  NOR2_X1 U17097 ( .A1(n13815), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13816) );
  AOI211_X1 U17098 ( .C1(n13888), .C2(P1_EAX_REG_27__SCAN_IN), .A(n13880), .B(
        n13816), .ZN(n13818) );
  XNOR2_X1 U17099 ( .A(n13817), .B(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14265) );
  AOI22_X1 U17100 ( .A1(n13819), .A2(n13818), .B1(n13880), .B2(n14265), .ZN(
        n14012) );
  INV_X1 U17101 ( .A(n13820), .ZN(n13821) );
  INV_X1 U17102 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n14000) );
  NAND2_X1 U17103 ( .A1(n13821), .A2(n14000), .ZN(n13822) );
  NAND2_X1 U17104 ( .A1(n13858), .A2(n13822), .ZN(n14258) );
  NOR2_X1 U17105 ( .A1(n13824), .A2(n13823), .ZN(n13842) );
  INV_X1 U17106 ( .A(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n20818) );
  AOI22_X1 U17107 ( .A1(n12709), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n9732), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n13829) );
  AOI22_X1 U17108 ( .A1(n9739), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12619), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n13828) );
  AOI22_X1 U17109 ( .A1(n12374), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n9756), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n13827) );
  AOI22_X1 U17110 ( .A1(n13862), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n13825), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13826) );
  NAND4_X1 U17111 ( .A1(n13829), .A2(n13828), .A3(n13827), .A4(n13826), .ZN(
        n13835) );
  AOI22_X1 U17112 ( .A1(n13843), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n13867), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n13833) );
  AOI22_X1 U17113 ( .A1(n12367), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n13769), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n13832) );
  AOI22_X1 U17114 ( .A1(n13848), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n12067), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13831) );
  NAND4_X1 U17115 ( .A1(n13833), .A2(n13832), .A3(n13831), .A4(n13830), .ZN(
        n13834) );
  OR2_X1 U17116 ( .A1(n13835), .A2(n13834), .ZN(n13841) );
  XNOR2_X1 U17117 ( .A(n13842), .B(n13841), .ZN(n13839) );
  AOI21_X1 U17118 ( .B1(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n12396), .A(
        n13880), .ZN(n13838) );
  NAND2_X1 U17119 ( .A1(n13888), .A2(P1_EAX_REG_28__SCAN_IN), .ZN(n13837) );
  OAI211_X1 U17120 ( .C1(n13839), .C2(n13883), .A(n13838), .B(n13837), .ZN(
        n13840) );
  OAI21_X1 U17121 ( .B1(n13886), .B2(n14258), .A(n13840), .ZN(n13998) );
  NAND2_X1 U17122 ( .A1(n13842), .A2(n13841), .ZN(n13876) );
  AOI22_X1 U17123 ( .A1(n13862), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n12709), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n13847) );
  AOI22_X1 U17124 ( .A1(n9732), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n13769), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n13846) );
  AOI22_X1 U17125 ( .A1(n13843), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12067), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n13845) );
  NAND4_X1 U17126 ( .A1(n13847), .A2(n13846), .A3(n13845), .A4(n13844), .ZN(
        n13854) );
  AOI22_X1 U17127 ( .A1(n12374), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12619), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n13852) );
  AOI22_X1 U17128 ( .A1(n9740), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12658), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13851) );
  AOI22_X1 U17129 ( .A1(n13477), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n13848), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n13850) );
  AOI22_X1 U17130 ( .A1(n9757), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n13825), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n13849) );
  NAND4_X1 U17131 ( .A1(n13852), .A2(n13851), .A3(n13850), .A4(n13849), .ZN(
        n13853) );
  NOR2_X1 U17132 ( .A1(n13854), .A2(n13853), .ZN(n13877) );
  XOR2_X1 U17133 ( .A(n13876), .B(n13877), .Z(n13856) );
  NAND2_X1 U17134 ( .A1(n13856), .A2(n13855), .ZN(n13860) );
  AOI21_X1 U17135 ( .B1(n13989), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n13857) );
  AOI21_X1 U17136 ( .B1(n13888), .B2(P1_EAX_REG_29__SCAN_IN), .A(n13857), .ZN(
        n13859) );
  XNOR2_X1 U17137 ( .A(n13858), .B(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n13988) );
  AOI22_X1 U17138 ( .A1(n13860), .A2(n13859), .B1(n13880), .B2(n13988), .ZN(
        n13987) );
  XNOR2_X1 U17139 ( .A(n13861), .B(n13976), .ZN(n14238) );
  AOI22_X1 U17140 ( .A1(n13862), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n12709), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n13866) );
  AOI22_X1 U17141 ( .A1(n12374), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12619), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n13865) );
  AOI22_X1 U17142 ( .A1(n13477), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n13769), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n13864) );
  AOI22_X1 U17143 ( .A1(n13848), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n9722), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n13863) );
  NAND4_X1 U17144 ( .A1(n13866), .A2(n13865), .A3(n13864), .A4(n13863), .ZN(
        n13875) );
  AOI22_X1 U17145 ( .A1(n13868), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n13867), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n13873) );
  AOI22_X1 U17146 ( .A1(n9741), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n9755), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n13872) );
  AOI22_X1 U17147 ( .A1(n9732), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n13825), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13871) );
  NAND4_X1 U17148 ( .A1(n13873), .A2(n13872), .A3(n13871), .A4(n13870), .ZN(
        n13874) );
  NOR2_X1 U17149 ( .A1(n13875), .A2(n13874), .ZN(n13879) );
  NOR2_X1 U17150 ( .A1(n13877), .A2(n13876), .ZN(n13878) );
  XOR2_X1 U17151 ( .A(n13879), .B(n13878), .Z(n13884) );
  AOI21_X1 U17152 ( .B1(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n12396), .A(
        n13880), .ZN(n13882) );
  NAND2_X1 U17153 ( .A1(n13888), .A2(P1_EAX_REG_30__SCAN_IN), .ZN(n13881) );
  OAI211_X1 U17154 ( .C1(n13884), .C2(n13883), .A(n13882), .B(n13881), .ZN(
        n13885) );
  OAI21_X1 U17155 ( .B1(n13886), .B2(n14238), .A(n13885), .ZN(n13975) );
  AOI22_X1 U17156 ( .A1(n13888), .A2(P1_EAX_REG_31__SCAN_IN), .B1(n13887), 
        .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n13889) );
  AND2_X1 U17157 ( .A1(n14191), .A2(n20047), .ZN(n13890) );
  NAND2_X1 U17158 ( .A1(n14229), .A2(n13890), .ZN(n13894) );
  NOR3_X1 U17159 ( .A1(n14194), .A2(n20006), .A3(n13891), .ZN(n13892) );
  AOI22_X1 U17160 ( .A1(n14188), .A2(DATAI_31_), .B1(P1_EAX_REG_31__SCAN_IN), 
        .B2(n14194), .ZN(n13893) );
  OAI211_X1 U17161 ( .C1(n14184), .C2(n16291), .A(n13894), .B(n13893), .ZN(
        P1_U2873) );
  AOI22_X1 U17162 ( .A1(n19049), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(
        n16157), .B2(n13895), .ZN(n13901) );
  AOI21_X1 U17163 ( .B1(n19059), .B2(n19712), .A(n13896), .ZN(n13900) );
  NAND2_X1 U17164 ( .A1(n19065), .A2(n13897), .ZN(n13899) );
  OAI211_X1 U17165 ( .C1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(n14998), .B(n19046), .ZN(n13898) );
  AND4_X1 U17166 ( .A1(n13901), .A2(n13900), .A3(n13899), .A4(n13898), .ZN(
        n13902) );
  OAI21_X1 U17167 ( .B1(n11154), .B2(n19061), .A(n13902), .ZN(P2_U3045) );
  NAND2_X1 U17168 ( .A1(n13903), .A2(P1_MEMORYFETCH_REG_SCAN_IN), .ZN(n13905)
         );
  NAND3_X1 U17169 ( .A1(n13905), .A2(n13904), .A3(n19760), .ZN(P1_U2801) );
  AOI22_X1 U17170 ( .A1(n13951), .A2(P1_EBX_REG_31__SCAN_IN), .B1(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n13950), .ZN(n13906) );
  AOI22_X1 U17171 ( .A1(n13951), .A2(P1_EBX_REG_30__SCAN_IN), .B1(
        P1_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n13950), .ZN(n13972) );
  XNOR2_X1 U17172 ( .A(n13906), .B(n13972), .ZN(n13953) );
  OR2_X1 U17173 ( .A1(n13906), .A2(n13971), .ZN(n13952) );
  INV_X1 U17174 ( .A(P1_EBX_REG_15__SCAN_IN), .ZN(n14119) );
  NAND2_X1 U17175 ( .A1(n13931), .A2(n14119), .ZN(n13909) );
  INV_X1 U17176 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15744) );
  NAND2_X1 U17177 ( .A1(n13944), .A2(n15744), .ZN(n13907) );
  OAI211_X1 U17178 ( .C1(n13950), .C2(P1_EBX_REG_15__SCAN_IN), .A(n13907), .B(
        n9724), .ZN(n13908) );
  MUX2_X1 U17179 ( .A(n13948), .B(n9724), .S(P1_EBX_REG_16__SCAN_IN), .Z(
        n13910) );
  OAI21_X1 U17180 ( .B1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n13951), .A(
        n13910), .ZN(n14110) );
  INV_X1 U17181 ( .A(P1_EBX_REG_17__SCAN_IN), .ZN(n15567) );
  NAND2_X1 U17182 ( .A1(n13931), .A2(n15567), .ZN(n13914) );
  INV_X1 U17183 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n13911) );
  NAND2_X1 U17184 ( .A1(n13944), .A2(n13911), .ZN(n13912) );
  OAI211_X1 U17185 ( .C1(n13950), .C2(P1_EBX_REG_17__SCAN_IN), .A(n13912), .B(
        n9724), .ZN(n13913) );
  NAND2_X1 U17186 ( .A1(n13914), .A2(n13913), .ZN(n14101) );
  NAND2_X1 U17187 ( .A1(n14109), .A2(n14101), .ZN(n14103) );
  MUX2_X1 U17188 ( .A(n13948), .B(n13936), .S(P1_EBX_REG_18__SCAN_IN), .Z(
        n13916) );
  INV_X1 U17189 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n14312) );
  NAND2_X1 U17190 ( .A1(n12450), .A2(n14312), .ZN(n13915) );
  NAND2_X1 U17191 ( .A1(n13916), .A2(n13915), .ZN(n14093) );
  INV_X1 U17192 ( .A(P1_EBX_REG_19__SCAN_IN), .ZN(n15552) );
  NAND2_X1 U17193 ( .A1(n13931), .A2(n15552), .ZN(n13919) );
  NAND2_X1 U17194 ( .A1(n13944), .A2(n15721), .ZN(n13917) );
  OAI211_X1 U17195 ( .C1(n13950), .C2(P1_EBX_REG_19__SCAN_IN), .A(n13917), .B(
        n9724), .ZN(n13918) );
  INV_X1 U17196 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n15640) );
  NAND2_X1 U17197 ( .A1(n13940), .A2(n15640), .ZN(n13922) );
  NAND2_X1 U17198 ( .A1(n9724), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n13920) );
  OAI211_X1 U17199 ( .C1(n13950), .C2(P1_EBX_REG_20__SCAN_IN), .A(n13944), .B(
        n13920), .ZN(n13921) );
  INV_X1 U17200 ( .A(P1_EBX_REG_21__SCAN_IN), .ZN(n20795) );
  NAND2_X1 U17201 ( .A1(n13931), .A2(n20795), .ZN(n13925) );
  INV_X1 U17202 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n14305) );
  NAND2_X1 U17203 ( .A1(n13944), .A2(n14305), .ZN(n13923) );
  OAI211_X1 U17204 ( .C1(n13950), .C2(P1_EBX_REG_21__SCAN_IN), .A(n13923), .B(
        n13936), .ZN(n13924) );
  NAND2_X1 U17205 ( .A1(n13925), .A2(n13924), .ZN(n14081) );
  MUX2_X1 U17206 ( .A(n13948), .B(n9724), .S(P1_EBX_REG_22__SCAN_IN), .Z(
        n13926) );
  OAI21_X1 U17207 ( .B1(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n13951), .A(
        n13926), .ZN(n15526) );
  INV_X1 U17208 ( .A(P1_EBX_REG_24__SCAN_IN), .ZN(n15635) );
  NAND2_X1 U17209 ( .A1(n13940), .A2(n15635), .ZN(n13929) );
  NAND2_X1 U17210 ( .A1(n9724), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n13927) );
  OAI211_X1 U17211 ( .C1(n13950), .C2(P1_EBX_REG_24__SCAN_IN), .A(n13944), .B(
        n13927), .ZN(n13928) );
  AND2_X1 U17212 ( .A1(n13929), .A2(n13928), .ZN(n14452) );
  INV_X1 U17213 ( .A(P1_EBX_REG_23__SCAN_IN), .ZN(n13930) );
  NAND2_X1 U17214 ( .A1(n13931), .A2(n13930), .ZN(n13934) );
  INV_X1 U17215 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15709) );
  NAND2_X1 U17216 ( .A1(n13944), .A2(n15709), .ZN(n13932) );
  OAI211_X1 U17217 ( .C1(n13950), .C2(P1_EBX_REG_23__SCAN_IN), .A(n13932), .B(
        n9724), .ZN(n13933) );
  NAND2_X1 U17218 ( .A1(n13934), .A2(n13933), .ZN(n14453) );
  NAND2_X1 U17219 ( .A1(n14452), .A2(n14453), .ZN(n13935) );
  INV_X1 U17220 ( .A(P1_EBX_REG_25__SCAN_IN), .ZN(n14074) );
  NAND2_X1 U17221 ( .A1(n13931), .A2(n14074), .ZN(n13939) );
  INV_X1 U17222 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n14435) );
  NAND2_X1 U17223 ( .A1(n13944), .A2(n14435), .ZN(n13937) );
  OAI211_X1 U17224 ( .C1(n13950), .C2(P1_EBX_REG_25__SCAN_IN), .A(n13937), .B(
        n13936), .ZN(n13938) );
  NAND2_X1 U17225 ( .A1(n13939), .A2(n13938), .ZN(n14037) );
  INV_X1 U17226 ( .A(P1_EBX_REG_26__SCAN_IN), .ZN(n14073) );
  NAND2_X1 U17227 ( .A1(n13940), .A2(n14073), .ZN(n13943) );
  NAND2_X1 U17228 ( .A1(n9724), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n13941) );
  OAI211_X1 U17229 ( .C1(n13950), .C2(P1_EBX_REG_26__SCAN_IN), .A(n13944), .B(
        n13941), .ZN(n13942) );
  AND2_X1 U17230 ( .A1(n13943), .A2(n13942), .ZN(n14019) );
  INV_X1 U17231 ( .A(P1_EBX_REG_27__SCAN_IN), .ZN(n14072) );
  NAND2_X1 U17232 ( .A1(n13931), .A2(n14072), .ZN(n13947) );
  INV_X1 U17233 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14422) );
  NAND2_X1 U17234 ( .A1(n13944), .A2(n14422), .ZN(n13945) );
  OAI211_X1 U17235 ( .C1(n13950), .C2(P1_EBX_REG_27__SCAN_IN), .A(n13945), .B(
        n9724), .ZN(n13946) );
  AND2_X1 U17236 ( .A1(n13947), .A2(n13946), .ZN(n14007) );
  MUX2_X1 U17237 ( .A(n13948), .B(n9724), .S(P1_EBX_REG_28__SCAN_IN), .Z(
        n13949) );
  OAI21_X1 U17238 ( .B1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n13951), .A(
        n13949), .ZN(n13999) );
  OAI22_X1 U17239 ( .A1(n13951), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .B1(
        P1_EBX_REG_29__SCAN_IN), .B2(n13950), .ZN(n13969) );
  OAI22_X1 U17240 ( .A1(n13969), .A2(n13971), .B1(P1_EBX_REG_29__SCAN_IN), 
        .B2(n9724), .ZN(n13984) );
  MUX2_X1 U17241 ( .A(n13953), .B(n13952), .S(n13983), .Z(n14382) );
  NAND2_X1 U17242 ( .A1(n14229), .A2(n19816), .ZN(n13968) );
  INV_X1 U17243 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n20631) );
  INV_X1 U17244 ( .A(P1_REIP_REG_19__SCAN_IN), .ZN(n20629) );
  INV_X1 U17245 ( .A(P1_REIP_REG_18__SCAN_IN), .ZN(n20627) );
  INV_X1 U17246 ( .A(P1_REIP_REG_12__SCAN_IN), .ZN(n20617) );
  INV_X1 U17247 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n20615) );
  INV_X1 U17248 ( .A(P1_REIP_REG_7__SCAN_IN), .ZN(n20609) );
  INV_X1 U17249 ( .A(P1_REIP_REG_5__SCAN_IN), .ZN(n20606) );
  NAND4_X1 U17250 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(P1_REIP_REG_1__SCAN_IN), 
        .A3(P1_REIP_REG_3__SCAN_IN), .A4(P1_REIP_REG_2__SCAN_IN), .ZN(n19827)
         );
  NOR2_X1 U17251 ( .A1(n20606), .A2(n19827), .ZN(n19817) );
  NAND2_X1 U17252 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(n19817), .ZN(n19806) );
  NOR2_X1 U17253 ( .A1(n20609), .A2(n19806), .ZN(n19791) );
  NAND2_X1 U17254 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(n19791), .ZN(n19781) );
  NOR2_X1 U17255 ( .A1(n20612), .A2(n19781), .ZN(n15619) );
  NAND2_X1 U17256 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(n15619), .ZN(n15614) );
  NOR3_X1 U17257 ( .A1(n20617), .A2(n20615), .A3(n15614), .ZN(n14063) );
  NAND3_X1 U17258 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(P1_REIP_REG_13__SCAN_IN), 
        .A3(n14063), .ZN(n15544) );
  NAND3_X1 U17259 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(P1_REIP_REG_16__SCAN_IN), 
        .A3(P1_REIP_REG_15__SCAN_IN), .ZN(n15548) );
  NOR4_X1 U17260 ( .A1(n20629), .A2(n20627), .A3(n15544), .A4(n15548), .ZN(
        n15538) );
  NAND2_X1 U17261 ( .A1(P1_REIP_REG_20__SCAN_IN), .A2(n15538), .ZN(n15529) );
  NOR2_X1 U17262 ( .A1(n20631), .A2(n15529), .ZN(n14047) );
  NAND3_X1 U17263 ( .A1(P1_REIP_REG_23__SCAN_IN), .A2(P1_REIP_REG_22__SCAN_IN), 
        .A3(n14047), .ZN(n13961) );
  INV_X1 U17264 ( .A(n13961), .ZN(n13954) );
  NAND2_X1 U17265 ( .A1(n15545), .A2(n13954), .ZN(n13955) );
  NAND2_X1 U17266 ( .A1(n19826), .A2(n13955), .ZN(n14048) );
  INV_X1 U17267 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n20637) );
  INV_X1 U17268 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n20636) );
  NOR2_X1 U17269 ( .A1(n20637), .A2(n20636), .ZN(n14033) );
  NAND2_X1 U17270 ( .A1(P1_REIP_REG_26__SCAN_IN), .A2(n14033), .ZN(n13956) );
  NAND2_X1 U17271 ( .A1(n19826), .A2(n13956), .ZN(n13957) );
  AND2_X1 U17272 ( .A1(n14048), .A2(n13957), .ZN(n14025) );
  NAND2_X1 U17273 ( .A1(P1_REIP_REG_28__SCAN_IN), .A2(P1_REIP_REG_27__SCAN_IN), 
        .ZN(n13962) );
  NAND2_X1 U17274 ( .A1(n19826), .A2(n13962), .ZN(n13958) );
  NAND2_X1 U17275 ( .A1(P1_REIP_REG_30__SCAN_IN), .A2(P1_REIP_REG_29__SCAN_IN), 
        .ZN(n13964) );
  NAND2_X1 U17276 ( .A1(n19826), .A2(n13964), .ZN(n13959) );
  NAND2_X1 U17277 ( .A1(n14004), .A2(n13959), .ZN(n13979) );
  INV_X1 U17278 ( .A(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n13960) );
  OAI22_X1 U17279 ( .A1(n19870), .A2(n14069), .B1(n13960), .B2(n19823), .ZN(
        n13966) );
  NOR2_X1 U17280 ( .A1(n19838), .A2(n13961), .ZN(n15515) );
  NAND2_X1 U17281 ( .A1(n15515), .A2(n14033), .ZN(n14026) );
  INV_X1 U17282 ( .A(P1_REIP_REG_26__SCAN_IN), .ZN(n20642) );
  NOR2_X1 U17283 ( .A1(n14026), .A2(n20642), .ZN(n14016) );
  INV_X1 U17284 ( .A(n13962), .ZN(n13963) );
  NAND2_X1 U17285 ( .A1(n14016), .A2(n13963), .ZN(n13992) );
  NOR3_X1 U17286 ( .A1(n13992), .A2(P1_REIP_REG_31__SCAN_IN), .A3(n13964), 
        .ZN(n13965) );
  AOI211_X1 U17287 ( .C1(P1_REIP_REG_31__SCAN_IN), .C2(n13979), .A(n13966), 
        .B(n13965), .ZN(n13967) );
  OAI211_X1 U17288 ( .C1(n14382), .C2(n19836), .A(n13968), .B(n13967), .ZN(
        P1_U2809) );
  INV_X1 U17289 ( .A(n13969), .ZN(n13970) );
  AOI22_X1 U17290 ( .A1(n13983), .A2(n13971), .B1(n13970), .B2(n9786), .ZN(
        n13973) );
  AOI21_X2 U17291 ( .B1(n13975), .B2(n13986), .A(n13974), .ZN(n14240) );
  NAND2_X1 U17292 ( .A1(n14240), .A2(n19816), .ZN(n13982) );
  INV_X1 U17293 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n14244) );
  INV_X1 U17294 ( .A(P1_REIP_REG_30__SCAN_IN), .ZN(n14236) );
  OAI21_X1 U17295 ( .B1(n13992), .B2(n14244), .A(n14236), .ZN(n13980) );
  INV_X1 U17296 ( .A(P1_EBX_REG_30__SCAN_IN), .ZN(n14070) );
  NOR2_X1 U17297 ( .A1(n19870), .A2(n14070), .ZN(n13978) );
  OAI22_X1 U17298 ( .A1(n13976), .A2(n19823), .B1(n19829), .B2(n14238), .ZN(
        n13977) );
  AOI211_X1 U17299 ( .C1(n13980), .C2(n13979), .A(n13978), .B(n13977), .ZN(
        n13981) );
  OAI211_X1 U17300 ( .C1(n19836), .C2(n14398), .A(n13982), .B(n13981), .ZN(
        P1_U2810) );
  OAI21_X1 U17301 ( .B1(n9786), .B2(n13984), .A(n13983), .ZN(n14407) );
  OAI21_X1 U17302 ( .B1(n13985), .B2(n13987), .A(n13986), .ZN(n14133) );
  INV_X1 U17303 ( .A(n14133), .ZN(n14248) );
  NAND2_X1 U17304 ( .A1(n14248), .A2(n19816), .ZN(n13996) );
  INV_X1 U17305 ( .A(n14004), .ZN(n13994) );
  INV_X1 U17306 ( .A(n13988), .ZN(n14246) );
  OAI22_X1 U17307 ( .A1(n13989), .A2(n19823), .B1(n19829), .B2(n14246), .ZN(
        n13990) );
  AOI21_X1 U17308 ( .B1(n19850), .B2(P1_EBX_REG_29__SCAN_IN), .A(n13990), .ZN(
        n13991) );
  OAI21_X1 U17309 ( .B1(n13992), .B2(P1_REIP_REG_29__SCAN_IN), .A(n13991), 
        .ZN(n13993) );
  AOI21_X1 U17310 ( .B1(P1_REIP_REG_29__SCAN_IN), .B2(n13994), .A(n13993), 
        .ZN(n13995) );
  OAI211_X1 U17311 ( .C1(n19836), .C2(n14407), .A(n13996), .B(n13995), .ZN(
        P1_U2811) );
  AOI21_X1 U17312 ( .B1(n13998), .B2(n14011), .A(n13985), .ZN(n14260) );
  INV_X1 U17313 ( .A(n14260), .ZN(n14136) );
  AOI21_X1 U17314 ( .B1(n13999), .B2(n14009), .A(n9786), .ZN(n14413) );
  INV_X1 U17315 ( .A(P1_REIP_REG_28__SCAN_IN), .ZN(n14256) );
  NAND3_X1 U17316 ( .A1(n14016), .A2(P1_REIP_REG_27__SCAN_IN), .A3(n14256), 
        .ZN(n14003) );
  OAI22_X1 U17317 ( .A1(n14000), .A2(n19823), .B1(n19829), .B2(n14258), .ZN(
        n14001) );
  AOI21_X1 U17318 ( .B1(n19850), .B2(P1_EBX_REG_28__SCAN_IN), .A(n14001), .ZN(
        n14002) );
  OAI211_X1 U17319 ( .C1(n14004), .C2(n14256), .A(n14003), .B(n14002), .ZN(
        n14005) );
  AOI21_X1 U17320 ( .B1(n14413), .B2(n19856), .A(n14005), .ZN(n14006) );
  OAI21_X1 U17321 ( .B1(n14136), .B2(n15589), .A(n14006), .ZN(P1_U2812) );
  NAND2_X1 U17322 ( .A1(n14021), .A2(n14007), .ZN(n14008) );
  NAND2_X1 U17323 ( .A1(n14009), .A2(n14008), .ZN(n14425) );
  OAI21_X1 U17324 ( .B1(n14010), .B2(n14012), .A(n14011), .ZN(n14139) );
  INV_X1 U17325 ( .A(n14139), .ZN(n14269) );
  NAND2_X1 U17326 ( .A1(n14269), .A2(n19816), .ZN(n14018) );
  INV_X1 U17327 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n20640) );
  AOI22_X1 U17328 ( .A1(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n19861), .B1(
        n19860), .B2(n14265), .ZN(n14013) );
  OAI21_X1 U17329 ( .B1(n19870), .B2(n14072), .A(n14013), .ZN(n14015) );
  NOR2_X1 U17330 ( .A1(n14025), .A2(n20640), .ZN(n14014) );
  AOI211_X1 U17331 ( .C1(n14016), .C2(n20640), .A(n14015), .B(n14014), .ZN(
        n14017) );
  OAI211_X1 U17332 ( .C1(n19836), .C2(n14425), .A(n14018), .B(n14017), .ZN(
        P1_U2813) );
  OR2_X1 U17333 ( .A1(n14039), .A2(n14019), .ZN(n14020) );
  NAND2_X1 U17334 ( .A1(n14021), .A2(n14020), .ZN(n14434) );
  AOI21_X1 U17335 ( .B1(n14023), .B2(n14022), .A(n14010), .ZN(n14277) );
  NAND2_X1 U17336 ( .A1(n14277), .A2(n19816), .ZN(n14030) );
  OAI22_X1 U17337 ( .A1(n14024), .A2(n19823), .B1(n19829), .B2(n14275), .ZN(
        n14028) );
  AOI21_X1 U17338 ( .B1(n20642), .B2(n14026), .A(n14025), .ZN(n14027) );
  AOI211_X1 U17339 ( .C1(P1_EBX_REG_26__SCAN_IN), .C2(n19850), .A(n14028), .B(
        n14027), .ZN(n14029) );
  OAI211_X1 U17340 ( .C1(n19836), .C2(n14434), .A(n14030), .B(n14029), .ZN(
        P1_U2814) );
  OAI21_X1 U17341 ( .B1(n14031), .B2(n14032), .A(n14022), .ZN(n14282) );
  INV_X1 U17342 ( .A(n14048), .ZN(n15516) );
  INV_X1 U17343 ( .A(n14033), .ZN(n14034) );
  OAI211_X1 U17344 ( .C1(P1_REIP_REG_24__SCAN_IN), .C2(P1_REIP_REG_25__SCAN_IN), .A(n15515), .B(n14034), .ZN(n14036) );
  AOI22_X1 U17345 ( .A1(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n19861), .B1(
        n19860), .B2(n14283), .ZN(n14035) );
  OAI211_X1 U17346 ( .C1(n14074), .C2(n19870), .A(n14036), .B(n14035), .ZN(
        n14041) );
  NOR2_X1 U17347 ( .A1(n14454), .A2(n14037), .ZN(n14038) );
  OR2_X1 U17348 ( .A1(n14039), .A2(n14038), .ZN(n14447) );
  NOR2_X1 U17349 ( .A1(n14447), .A2(n19836), .ZN(n14040) );
  AOI211_X1 U17350 ( .C1(n15516), .C2(P1_REIP_REG_25__SCAN_IN), .A(n14041), 
        .B(n14040), .ZN(n14042) );
  OAI21_X1 U17351 ( .B1(n14282), .B2(n15589), .A(n14042), .ZN(P1_U2815) );
  INV_X1 U17352 ( .A(n14044), .ZN(n14045) );
  AOI21_X1 U17353 ( .B1(n14046), .B2(n14043), .A(n14045), .ZN(n14301) );
  INV_X1 U17354 ( .A(n14301), .ZN(n14155) );
  XNOR2_X1 U17355 ( .A(n14451), .B(n14453), .ZN(n15705) );
  AND2_X1 U17356 ( .A1(n19857), .A2(n14047), .ZN(n15524) );
  AOI21_X1 U17357 ( .B1(P1_REIP_REG_22__SCAN_IN), .B2(n15524), .A(
        P1_REIP_REG_23__SCAN_IN), .ZN(n14049) );
  INV_X1 U17358 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n20901) );
  OAI22_X1 U17359 ( .A1(n14049), .A2(n14048), .B1(n20901), .B2(n19823), .ZN(
        n14052) );
  INV_X1 U17360 ( .A(n14050), .ZN(n14299) );
  OAI22_X1 U17361 ( .A1(n19870), .A2(n13930), .B1(n14299), .B2(n19829), .ZN(
        n14051) );
  AOI211_X1 U17362 ( .C1(n15705), .C2(n19856), .A(n14052), .B(n14051), .ZN(
        n14053) );
  OAI21_X1 U17363 ( .B1(n14155), .B2(n15589), .A(n14053), .ZN(P1_U2817) );
  INV_X1 U17364 ( .A(n14054), .ZN(n14055) );
  AOI21_X1 U17365 ( .B1(n14056), .B2(n14055), .A(n9799), .ZN(n14361) );
  NAND2_X1 U17366 ( .A1(n14361), .A2(n19816), .ZN(n14068) );
  INV_X1 U17367 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n14057) );
  NOR2_X1 U17368 ( .A1(n19823), .A2(n14057), .ZN(n14066) );
  INV_X1 U17369 ( .A(n14058), .ZN(n14061) );
  NAND2_X1 U17370 ( .A1(n14503), .A2(n14059), .ZN(n14060) );
  NAND2_X1 U17371 ( .A1(n14061), .A2(n14060), .ZN(n15759) );
  INV_X1 U17372 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n20619) );
  INV_X1 U17373 ( .A(n14063), .ZN(n14062) );
  OAI21_X1 U17374 ( .B1(n19828), .B2(n14062), .A(n19826), .ZN(n15610) );
  OAI22_X1 U17375 ( .A1(n19836), .A2(n15759), .B1(n20619), .B2(n15610), .ZN(
        n14065) );
  NAND2_X1 U17376 ( .A1(n19857), .A2(n14063), .ZN(n15597) );
  OAI22_X1 U17377 ( .A1(P1_REIP_REG_13__SCAN_IN), .A2(n15597), .B1(n14123), 
        .B2(n19870), .ZN(n14064) );
  NOR4_X1 U17378 ( .A1(n14066), .A2(n14065), .A3(n13009), .A4(n14064), .ZN(
        n14067) );
  OAI211_X1 U17379 ( .C1(n19829), .C2(n14359), .A(n14068), .B(n14067), .ZN(
        P1_U2827) );
  OAI22_X1 U17380 ( .A1(n14382), .A2(n14120), .B1(n14069), .B2(n19879), .ZN(
        P1_U2841) );
  INV_X1 U17381 ( .A(n14240), .ZN(n14128) );
  OAI222_X1 U17382 ( .A1(n15631), .A2(n14128), .B1(n19879), .B2(n14070), .C1(
        n14398), .C2(n14120), .ZN(P1_U2842) );
  INV_X1 U17383 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n20732) );
  OAI222_X1 U17384 ( .A1(n20732), .A2(n19879), .B1(n14120), .B2(n14407), .C1(
        n14133), .C2(n15631), .ZN(P1_U2843) );
  AOI22_X1 U17385 ( .A1(n14413), .A2(n19875), .B1(n14111), .B2(
        P1_EBX_REG_28__SCAN_IN), .ZN(n14071) );
  OAI21_X1 U17386 ( .B1(n14136), .B2(n15631), .A(n14071), .ZN(P1_U2844) );
  OAI222_X1 U17387 ( .A1(n14072), .A2(n19879), .B1(n14120), .B2(n14425), .C1(
        n14139), .C2(n15631), .ZN(P1_U2845) );
  INV_X1 U17388 ( .A(n14277), .ZN(n14143) );
  OAI222_X1 U17389 ( .A1(n14073), .A2(n19879), .B1(n14120), .B2(n14434), .C1(
        n14143), .C2(n15631), .ZN(P1_U2846) );
  OAI222_X1 U17390 ( .A1(n14074), .A2(n19879), .B1(n14120), .B2(n14447), .C1(
        n14282), .C2(n15631), .ZN(P1_U2847) );
  AOI22_X1 U17391 ( .A1(n15705), .A2(n19875), .B1(n14111), .B2(
        P1_EBX_REG_23__SCAN_IN), .ZN(n14075) );
  OAI21_X1 U17392 ( .B1(n14155), .B2(n15631), .A(n14075), .ZN(P1_U2849) );
  AND2_X1 U17393 ( .A1(n14163), .A2(n14078), .ZN(n14080) );
  OR2_X1 U17394 ( .A1(n14080), .A2(n14079), .ZN(n15533) );
  INV_X1 U17395 ( .A(n15533), .ZN(n14310) );
  OR2_X1 U17396 ( .A1(n15502), .A2(n14081), .ZN(n14082) );
  NAND2_X1 U17397 ( .A1(n9764), .A2(n14082), .ZN(n15537) );
  OAI22_X1 U17398 ( .A1(n15537), .A2(n14120), .B1(n20795), .B2(n19879), .ZN(
        n14083) );
  AOI21_X1 U17399 ( .B1(n14310), .B2(n19876), .A(n14083), .ZN(n14084) );
  INV_X1 U17400 ( .A(n14084), .ZN(P1_U2851) );
  INV_X1 U17401 ( .A(n14165), .ZN(n14085) );
  AOI21_X1 U17402 ( .B1(n14086), .B2(n14076), .A(n14085), .ZN(n14318) );
  AND2_X1 U17403 ( .A1(n14095), .A2(n14087), .ZN(n14088) );
  OR2_X1 U17404 ( .A1(n14088), .A2(n15501), .ZN(n15725) );
  OAI22_X1 U17405 ( .A1(n15725), .A2(n14120), .B1(n15552), .B2(n19879), .ZN(
        n14089) );
  AOI21_X1 U17406 ( .B1(n14318), .B2(n19876), .A(n14089), .ZN(n14090) );
  INV_X1 U17407 ( .A(n14090), .ZN(P1_U2853) );
  OR2_X1 U17408 ( .A1(n14100), .A2(n14091), .ZN(n14092) );
  AND2_X1 U17409 ( .A1(n14076), .A2(n14092), .ZN(n15563) );
  INV_X1 U17410 ( .A(n15563), .ZN(n14178) );
  INV_X1 U17411 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n14096) );
  NAND2_X1 U17412 ( .A1(n14103), .A2(n14093), .ZN(n14094) );
  NAND2_X1 U17413 ( .A1(n14095), .A2(n14094), .ZN(n15561) );
  OAI222_X1 U17414 ( .A1(n14178), .A2(n15631), .B1(n19879), .B2(n14096), .C1(
        n15561), .C2(n14120), .ZN(P1_U2854) );
  NOR2_X1 U17415 ( .A1(n14097), .A2(n14098), .ZN(n14099) );
  OR2_X1 U17416 ( .A1(n14100), .A2(n14099), .ZN(n15571) );
  OR2_X1 U17417 ( .A1(n14109), .A2(n14101), .ZN(n14102) );
  NAND2_X1 U17418 ( .A1(n14103), .A2(n14102), .ZN(n15732) );
  OAI22_X1 U17419 ( .A1(n15732), .A2(n14120), .B1(n15567), .B2(n19879), .ZN(
        n14104) );
  INV_X1 U17420 ( .A(n14104), .ZN(n14105) );
  OAI21_X1 U17421 ( .B1(n15571), .B2(n15631), .A(n14105), .ZN(P1_U2855) );
  AND2_X1 U17422 ( .A1(n14113), .A2(n14107), .ZN(n14108) );
  OR2_X1 U17423 ( .A1(n14108), .A2(n14097), .ZN(n15578) );
  AOI21_X1 U17424 ( .B1(n14110), .B2(n14118), .A(n14109), .ZN(n15737) );
  AOI22_X1 U17425 ( .A1(n15737), .A2(n19875), .B1(P1_EBX_REG_16__SCAN_IN), 
        .B2(n14111), .ZN(n14112) );
  OAI21_X1 U17426 ( .B1(n15578), .B2(n15631), .A(n14112), .ZN(P1_U2856) );
  AOI21_X1 U17427 ( .B1(n14114), .B2(n13588), .A(n14106), .ZN(n14347) );
  NAND2_X1 U17428 ( .A1(n14116), .A2(n14115), .ZN(n14117) );
  NAND2_X1 U17429 ( .A1(n14118), .A2(n14117), .ZN(n15749) );
  OAI22_X1 U17430 ( .A1(n15749), .A2(n14120), .B1(n14119), .B2(n19879), .ZN(
        n14121) );
  AOI21_X1 U17431 ( .B1(n14347), .B2(n19876), .A(n14121), .ZN(n14122) );
  INV_X1 U17432 ( .A(n14122), .ZN(P1_U2857) );
  OAI22_X1 U17433 ( .A1(n15759), .A2(n14120), .B1(n14123), .B2(n19879), .ZN(
        n14124) );
  AOI21_X1 U17434 ( .B1(n14361), .B2(n19876), .A(n14124), .ZN(n14125) );
  INV_X1 U17435 ( .A(n14125), .ZN(P1_U2859) );
  AOI22_X1 U17436 ( .A1(n14179), .A2(BUF1_REG_30__SCAN_IN), .B1(
        P1_EAX_REG_30__SCAN_IN), .B2(n14194), .ZN(n14127) );
  NOR3_X2 U17437 ( .A1(n14194), .A2(n20047), .A3(n12121), .ZN(n14181) );
  AOI22_X1 U17438 ( .A1(n14181), .A2(n19919), .B1(n14188), .B2(DATAI_30_), 
        .ZN(n14126) );
  OAI211_X1 U17439 ( .C1(n14128), .C2(n14197), .A(n14127), .B(n14126), .ZN(
        P1_U2874) );
  AOI22_X1 U17440 ( .A1(n14179), .A2(BUF1_REG_29__SCAN_IN), .B1(
        P1_EAX_REG_29__SCAN_IN), .B2(n14194), .ZN(n14132) );
  INV_X1 U17441 ( .A(DATAI_13_), .ZN(n14130) );
  NAND2_X1 U17442 ( .A1(n20006), .A2(BUF1_REG_13__SCAN_IN), .ZN(n14129) );
  OAI21_X1 U17443 ( .B1(n20006), .B2(n14130), .A(n14129), .ZN(n19917) );
  AOI22_X1 U17444 ( .A1(n14181), .A2(n19917), .B1(n14188), .B2(DATAI_29_), 
        .ZN(n14131) );
  OAI211_X1 U17445 ( .C1(n14133), .C2(n14197), .A(n14132), .B(n14131), .ZN(
        P1_U2875) );
  AOI22_X1 U17446 ( .A1(n14179), .A2(BUF1_REG_28__SCAN_IN), .B1(
        P1_EAX_REG_28__SCAN_IN), .B2(n14194), .ZN(n14135) );
  AOI22_X1 U17447 ( .A1(n14181), .A2(n19915), .B1(n14188), .B2(DATAI_28_), 
        .ZN(n14134) );
  OAI211_X1 U17448 ( .C1(n14136), .C2(n14197), .A(n14135), .B(n14134), .ZN(
        P1_U2876) );
  AOI22_X1 U17449 ( .A1(n14179), .A2(BUF1_REG_27__SCAN_IN), .B1(
        P1_EAX_REG_27__SCAN_IN), .B2(n14194), .ZN(n14138) );
  AOI22_X1 U17450 ( .A1(n14181), .A2(n19913), .B1(n14188), .B2(DATAI_27_), 
        .ZN(n14137) );
  OAI211_X1 U17451 ( .C1(n14139), .C2(n14197), .A(n14138), .B(n14137), .ZN(
        P1_U2877) );
  AOI22_X1 U17452 ( .A1(n14179), .A2(BUF1_REG_26__SCAN_IN), .B1(
        P1_EAX_REG_26__SCAN_IN), .B2(n14194), .ZN(n14142) );
  AOI22_X1 U17453 ( .A1(n14181), .A2(n14140), .B1(n14188), .B2(DATAI_26_), 
        .ZN(n14141) );
  OAI211_X1 U17454 ( .C1(n14143), .C2(n14197), .A(n14142), .B(n14141), .ZN(
        P1_U2878) );
  AOI22_X1 U17455 ( .A1(n14179), .A2(BUF1_REG_25__SCAN_IN), .B1(
        P1_EAX_REG_25__SCAN_IN), .B2(n14194), .ZN(n14145) );
  AOI22_X1 U17456 ( .A1(n14181), .A2(n19910), .B1(n14188), .B2(DATAI_25_), 
        .ZN(n14144) );
  OAI211_X1 U17457 ( .C1(n14282), .C2(n14197), .A(n14145), .B(n14144), .ZN(
        P1_U2879) );
  AND2_X1 U17458 ( .A1(n14044), .A2(n14146), .ZN(n14147) );
  OR2_X1 U17459 ( .A1(n14147), .A2(n14031), .ZN(n15632) );
  INV_X1 U17460 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n16303) );
  OAI22_X1 U17461 ( .A1(n14184), .A2(n16303), .B1(n12319), .B2(n14191), .ZN(
        n14148) );
  INV_X1 U17462 ( .A(n14148), .ZN(n14150) );
  AOI22_X1 U17463 ( .A1(n14181), .A2(n19907), .B1(n14188), .B2(DATAI_24_), 
        .ZN(n14149) );
  OAI211_X1 U17464 ( .C1(n15632), .C2(n14197), .A(n14150), .B(n14149), .ZN(
        P1_U2880) );
  INV_X1 U17465 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n14151) );
  OAI22_X1 U17466 ( .A1(n14184), .A2(n14151), .B1(n20835), .B2(n14191), .ZN(
        n14153) );
  INV_X1 U17467 ( .A(n14181), .ZN(n14185) );
  NOR2_X1 U17468 ( .A1(n14185), .A2(n20050), .ZN(n14152) );
  AOI211_X1 U17469 ( .C1(n14188), .C2(DATAI_23_), .A(n14153), .B(n14152), .ZN(
        n14154) );
  OAI21_X1 U17470 ( .B1(n14155), .B2(n14197), .A(n14154), .ZN(P1_U2881) );
  OAI21_X1 U17471 ( .B1(n14079), .B2(n14156), .A(n14043), .ZN(n15525) );
  INV_X1 U17472 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n16306) );
  OAI22_X1 U17473 ( .A1(n14184), .A2(n16306), .B1(n12585), .B2(n14191), .ZN(
        n14158) );
  NOR2_X1 U17474 ( .A1(n14185), .A2(n20043), .ZN(n14157) );
  AOI211_X1 U17475 ( .C1(n14188), .C2(DATAI_22_), .A(n14158), .B(n14157), .ZN(
        n14159) );
  OAI21_X1 U17476 ( .B1(n15525), .B2(n14197), .A(n14159), .ZN(P1_U2882) );
  AOI22_X1 U17477 ( .A1(n14179), .A2(BUF1_REG_21__SCAN_IN), .B1(
        P1_EAX_REG_21__SCAN_IN), .B2(n14194), .ZN(n14162) );
  AOI22_X1 U17478 ( .A1(n14181), .A2(n14160), .B1(n14188), .B2(DATAI_21_), 
        .ZN(n14161) );
  OAI211_X1 U17479 ( .C1(n15533), .C2(n14197), .A(n14162), .B(n14161), .ZN(
        P1_U2883) );
  INV_X1 U17480 ( .A(n14163), .ZN(n14164) );
  INV_X1 U17481 ( .A(n15652), .ZN(n14170) );
  INV_X1 U17482 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n19081) );
  OAI22_X1 U17483 ( .A1(n14184), .A2(n19081), .B1(n12589), .B2(n14191), .ZN(
        n14168) );
  NOR2_X1 U17484 ( .A1(n14185), .A2(n20035), .ZN(n14167) );
  AOI211_X1 U17485 ( .C1(n14188), .C2(DATAI_20_), .A(n14168), .B(n14167), .ZN(
        n14169) );
  OAI21_X1 U17486 ( .B1(n14170), .B2(n14197), .A(n14169), .ZN(P1_U2884) );
  INV_X1 U17487 ( .A(n14318), .ZN(n15553) );
  AOI22_X1 U17488 ( .A1(n14179), .A2(BUF1_REG_19__SCAN_IN), .B1(
        P1_EAX_REG_19__SCAN_IN), .B2(n14194), .ZN(n14173) );
  AOI22_X1 U17489 ( .A1(n14181), .A2(n14171), .B1(n14188), .B2(DATAI_19_), 
        .ZN(n14172) );
  OAI211_X1 U17490 ( .C1(n15553), .C2(n14197), .A(n14173), .B(n14172), .ZN(
        P1_U2885) );
  INV_X1 U17491 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n14174) );
  OAI22_X1 U17492 ( .A1(n14184), .A2(n14174), .B1(n20934), .B2(n14191), .ZN(
        n14176) );
  NOR2_X1 U17493 ( .A1(n14185), .A2(n20027), .ZN(n14175) );
  AOI211_X1 U17494 ( .C1(n14188), .C2(DATAI_18_), .A(n14176), .B(n14175), .ZN(
        n14177) );
  OAI21_X1 U17495 ( .B1(n14178), .B2(n14197), .A(n14177), .ZN(P1_U2886) );
  AOI22_X1 U17496 ( .A1(n14179), .A2(BUF1_REG_17__SCAN_IN), .B1(
        P1_EAX_REG_17__SCAN_IN), .B2(n14194), .ZN(n14183) );
  AOI22_X1 U17497 ( .A1(n14181), .A2(n14180), .B1(n14188), .B2(DATAI_17_), 
        .ZN(n14182) );
  OAI211_X1 U17498 ( .C1(n15571), .C2(n14197), .A(n14183), .B(n14182), .ZN(
        P1_U2887) );
  OAI22_X1 U17499 ( .A1(n14184), .A2(n16315), .B1(n12324), .B2(n14191), .ZN(
        n14187) );
  NOR2_X1 U17500 ( .A1(n14185), .A2(n20017), .ZN(n14186) );
  AOI211_X1 U17501 ( .C1(n14188), .C2(DATAI_16_), .A(n14187), .B(n14186), .ZN(
        n14189) );
  OAI21_X1 U17502 ( .B1(n15578), .B2(n14197), .A(n14189), .ZN(P1_U2888) );
  INV_X1 U17503 ( .A(n14347), .ZN(n15590) );
  OAI222_X1 U17504 ( .A1(n15590), .A2(n14197), .B1(n14193), .B2(n14192), .C1(
        n14191), .C2(n14190), .ZN(P1_U2889) );
  INV_X1 U17505 ( .A(n14361), .ZN(n14198) );
  AOI22_X1 U17506 ( .A1(n14195), .A2(n19917), .B1(P1_EAX_REG_13__SCAN_IN), 
        .B2(n14194), .ZN(n14196) );
  OAI21_X1 U17507 ( .B1(n14198), .B2(n14197), .A(n14196), .ZN(P1_U2891) );
  OR2_X1 U17508 ( .A1(n13402), .A2(n20819), .ZN(n14477) );
  NAND2_X1 U17509 ( .A1(n9750), .A2(n20819), .ZN(n14202) );
  NAND2_X1 U17510 ( .A1(n14477), .A2(n14202), .ZN(n14357) );
  INV_X1 U17511 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n14203) );
  NAND2_X1 U17512 ( .A1(n9749), .A2(n14203), .ZN(n14355) );
  NAND2_X1 U17513 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n14204) );
  NAND2_X1 U17514 ( .A1(n9750), .A2(n14204), .ZN(n14351) );
  NAND2_X1 U17515 ( .A1(n14355), .A2(n14351), .ZN(n14205) );
  NOR2_X1 U17516 ( .A1(n14357), .A2(n14205), .ZN(n14476) );
  INV_X1 U17517 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n15734) );
  NAND2_X1 U17518 ( .A1(n9750), .A2(n15734), .ZN(n14206) );
  NAND2_X1 U17519 ( .A1(n14476), .A2(n14206), .ZN(n14338) );
  NOR2_X1 U17520 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n14207) );
  OR2_X1 U17521 ( .A1(n9749), .A2(n14207), .ZN(n14208) );
  AND2_X1 U17522 ( .A1(n14341), .A2(n14208), .ZN(n14329) );
  NAND2_X1 U17523 ( .A1(n9749), .A2(n15744), .ZN(n15656) );
  INV_X1 U17524 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n14209) );
  NAND2_X1 U17525 ( .A1(n14210), .A2(n14209), .ZN(n14350) );
  NAND3_X1 U17526 ( .A1(n20819), .A2(n15734), .A3(n14203), .ZN(n14211) );
  NOR2_X1 U17527 ( .A1(n14350), .A2(n14211), .ZN(n14212) );
  OR2_X1 U17528 ( .A1(n9749), .A2(n14212), .ZN(n14339) );
  NAND2_X1 U17529 ( .A1(n14341), .A2(n14339), .ZN(n15657) );
  NOR2_X1 U17530 ( .A1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n14213) );
  NOR2_X1 U17531 ( .A1(n9749), .A2(n14213), .ZN(n14214) );
  XNOR2_X1 U17532 ( .A(n9749), .B(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14322) );
  NAND2_X1 U17533 ( .A1(n14216), .A2(n9749), .ZN(n15644) );
  INV_X1 U17534 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15497) );
  NAND2_X1 U17535 ( .A1(n14305), .A2(n15497), .ZN(n14218) );
  NOR2_X1 U17536 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14250) );
  NAND2_X1 U17537 ( .A1(n14250), .A2(n15709), .ZN(n14219) );
  NAND2_X1 U17538 ( .A1(n14232), .A2(n14354), .ZN(n14220) );
  AND2_X1 U17539 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14436) );
  NAND2_X1 U17540 ( .A1(n14436), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14430) );
  AND2_X1 U17541 ( .A1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14389) );
  NAND2_X1 U17542 ( .A1(n14263), .A2(n14389), .ZN(n14231) );
  NAND2_X1 U17543 ( .A1(n14220), .A2(n14231), .ZN(n14243) );
  INV_X1 U17544 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14397) );
  MUX2_X1 U17545 ( .A(n14221), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .S(
        n9750), .Z(n14222) );
  OAI211_X1 U17546 ( .C1(n14243), .C2(n14397), .A(n14223), .B(n14222), .ZN(
        n14224) );
  XNOR2_X1 U17547 ( .A(n14224), .B(n12562), .ZN(n14395) );
  INV_X1 U17548 ( .A(P1_REIP_REG_31__SCAN_IN), .ZN(n14225) );
  NOR2_X1 U17549 ( .A1(n19845), .A2(n14225), .ZN(n14391) );
  AOI21_X1 U17550 ( .B1(n19938), .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n14391), .ZN(n14226) );
  OAI21_X1 U17551 ( .B1(n15701), .B2(n14227), .A(n14226), .ZN(n14228) );
  OAI21_X1 U17552 ( .B1(n14395), .B2(n19764), .A(n14230), .ZN(P1_U2968) );
  NOR2_X1 U17553 ( .A1(n14231), .A2(n14221), .ZN(n14234) );
  NOR2_X1 U17554 ( .A1(n14232), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14233) );
  MUX2_X1 U17555 ( .A(n14234), .B(n14233), .S(n14354), .Z(n14235) );
  XNOR2_X1 U17556 ( .A(n14235), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14402) );
  NOR2_X1 U17557 ( .A1(n19845), .A2(n14236), .ZN(n14399) );
  AOI21_X1 U17558 ( .B1(n19938), .B2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n14399), .ZN(n14237) );
  OAI21_X1 U17559 ( .B1(n15701), .B2(n14238), .A(n14237), .ZN(n14239) );
  AOI21_X1 U17560 ( .B1(n14240), .B2(n9727), .A(n14239), .ZN(n14241) );
  OAI21_X1 U17561 ( .B1(n19764), .B2(n14402), .A(n14241), .ZN(P1_U2969) );
  XNOR2_X1 U17562 ( .A(n9750), .B(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14242) );
  XNOR2_X1 U17563 ( .A(n14243), .B(n14242), .ZN(n14411) );
  NOR2_X1 U17564 ( .A1(n19845), .A2(n14244), .ZN(n14404) );
  AOI21_X1 U17565 ( .B1(n19938), .B2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n14404), .ZN(n14245) );
  OAI21_X1 U17566 ( .B1(n15701), .B2(n14246), .A(n14245), .ZN(n14247) );
  AOI21_X1 U17567 ( .B1(n14248), .B2(n9727), .A(n14247), .ZN(n14249) );
  OAI21_X1 U17568 ( .B1(n14411), .B2(n19764), .A(n14249), .ZN(P1_U2970) );
  NAND2_X1 U17569 ( .A1(n9749), .A2(n14430), .ZN(n14271) );
  NAND2_X1 U17570 ( .A1(n14297), .A2(n14271), .ZN(n14254) );
  INV_X1 U17571 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14438) );
  NAND3_X1 U17572 ( .A1(n14250), .A2(n15709), .A3(n14438), .ZN(n14251) );
  NAND2_X1 U17573 ( .A1(n14254), .A2(n14251), .ZN(n14253) );
  MUX2_X1 U17574 ( .A(n14422), .B(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .S(
        n9750), .Z(n14252) );
  OAI211_X1 U17575 ( .C1(n14254), .C2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n14253), .B(n14252), .ZN(n14255) );
  XOR2_X1 U17576 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .B(n14255), .Z(
        n14420) );
  NOR2_X1 U17577 ( .A1(n19845), .A2(n14256), .ZN(n14414) );
  AOI21_X1 U17578 ( .B1(n19938), .B2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n14414), .ZN(n14257) );
  OAI21_X1 U17579 ( .B1(n15701), .B2(n14258), .A(n14257), .ZN(n14259) );
  AOI21_X1 U17580 ( .B1(n14260), .B2(n9727), .A(n14259), .ZN(n14261) );
  OAI21_X1 U17581 ( .B1(n19764), .B2(n14420), .A(n14261), .ZN(P1_U2971) );
  MUX2_X1 U17582 ( .A(n14263), .B(n14262), .S(n14354), .Z(n14264) );
  XNOR2_X1 U17583 ( .A(n14264), .B(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14429) );
  INV_X1 U17584 ( .A(n14265), .ZN(n14267) );
  NOR2_X1 U17585 ( .A1(n19845), .A2(n20640), .ZN(n14421) );
  AOI21_X1 U17586 ( .B1(n19938), .B2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n14421), .ZN(n14266) );
  OAI21_X1 U17587 ( .B1(n15701), .B2(n14267), .A(n14266), .ZN(n14268) );
  AOI21_X1 U17588 ( .B1(n14269), .B2(n9727), .A(n14268), .ZN(n14270) );
  OAI21_X1 U17589 ( .B1(n19764), .B2(n14429), .A(n14270), .ZN(P1_U2972) );
  OAI211_X1 U17590 ( .C1(n14272), .C2(n9749), .A(n14279), .B(n14271), .ZN(
        n14273) );
  XNOR2_X1 U17591 ( .A(n14273), .B(n14438), .ZN(n14443) );
  NOR2_X1 U17592 ( .A1(n19845), .A2(n20642), .ZN(n14431) );
  AOI21_X1 U17593 ( .B1(n19938), .B2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n14431), .ZN(n14274) );
  OAI21_X1 U17594 ( .B1(n15701), .B2(n14275), .A(n14274), .ZN(n14276) );
  AOI21_X1 U17595 ( .B1(n14277), .B2(n9727), .A(n14276), .ZN(n14278) );
  OAI21_X1 U17596 ( .B1(n19764), .B2(n14443), .A(n14278), .ZN(P1_U2973) );
  INV_X1 U17597 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14376) );
  XNOR2_X1 U17598 ( .A(n9750), .B(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14296) );
  OAI211_X1 U17599 ( .C1(n14376), .C2(n9749), .A(n14279), .B(n14296), .ZN(
        n14280) );
  INV_X1 U17600 ( .A(n14282), .ZN(n14287) );
  INV_X1 U17601 ( .A(n14283), .ZN(n14285) );
  NOR2_X1 U17602 ( .A1(n19845), .A2(n20637), .ZN(n14444) );
  AOI21_X1 U17603 ( .B1(n19938), .B2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n14444), .ZN(n14284) );
  OAI21_X1 U17604 ( .B1(n15701), .B2(n14285), .A(n14284), .ZN(n14286) );
  AOI21_X1 U17605 ( .B1(n14287), .B2(n9727), .A(n14286), .ZN(n14288) );
  OAI21_X1 U17606 ( .B1(n19764), .B2(n14448), .A(n14288), .ZN(P1_U2974) );
  NOR2_X1 U17607 ( .A1(n9749), .A2(n15709), .ZN(n14289) );
  OAI22_X1 U17608 ( .A1(n14297), .A2(n14289), .B1(n14354), .B2(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n14291) );
  XNOR2_X1 U17609 ( .A(n9750), .B(n14376), .ZN(n14290) );
  XNOR2_X1 U17610 ( .A(n14291), .B(n14290), .ZN(n14465) );
  INV_X1 U17611 ( .A(n15632), .ZN(n14294) );
  NOR2_X1 U17612 ( .A1(n19845), .A2(n20636), .ZN(n14458) );
  AOI21_X1 U17613 ( .B1(n19938), .B2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n14458), .ZN(n14292) );
  OAI21_X1 U17614 ( .B1(n15701), .B2(n15520), .A(n14292), .ZN(n14293) );
  AOI21_X1 U17615 ( .B1(n14294), .B2(n9727), .A(n14293), .ZN(n14295) );
  OAI21_X1 U17616 ( .B1(n19764), .B2(n14465), .A(n14295), .ZN(P1_U2975) );
  XNOR2_X1 U17617 ( .A(n14297), .B(n14296), .ZN(n15704) );
  AOI22_X1 U17618 ( .A1(n19938), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .B1(
        n13009), .B2(P1_REIP_REG_23__SCAN_IN), .ZN(n14298) );
  OAI21_X1 U17619 ( .B1(n15701), .B2(n14299), .A(n14298), .ZN(n14300) );
  AOI21_X1 U17620 ( .B1(n14301), .B2(n9727), .A(n14300), .ZN(n14302) );
  OAI21_X1 U17621 ( .B1(n15704), .B2(n19764), .A(n14302), .ZN(P1_U2976) );
  INV_X1 U17622 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15721) );
  NOR3_X1 U17623 ( .A1(n14321), .A2(n14354), .A3(n15721), .ZN(n15500) );
  INV_X1 U17624 ( .A(n14303), .ZN(n14304) );
  NAND2_X1 U17625 ( .A1(n14304), .A2(n14354), .ZN(n15495) );
  NOR2_X1 U17626 ( .A1(n15495), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15496) );
  AOI21_X1 U17627 ( .B1(n15500), .B2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n15496), .ZN(n14306) );
  XNOR2_X1 U17628 ( .A(n14306), .B(n14305), .ZN(n15467) );
  INV_X1 U17629 ( .A(n14307), .ZN(n15532) );
  AOI22_X1 U17630 ( .A1(n19938), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B1(
        n13009), .B2(P1_REIP_REG_21__SCAN_IN), .ZN(n14308) );
  OAI21_X1 U17631 ( .B1(n15701), .B2(n15532), .A(n14308), .ZN(n14309) );
  AOI21_X1 U17632 ( .B1(n14310), .B2(n9727), .A(n14309), .ZN(n14311) );
  OAI21_X1 U17633 ( .B1(n15467), .B2(n19764), .A(n14311), .ZN(P1_U2978) );
  NAND2_X1 U17634 ( .A1(n14321), .A2(n14312), .ZN(n14313) );
  MUX2_X1 U17635 ( .A(n14321), .B(n14313), .S(n14354), .Z(n14314) );
  XOR2_X1 U17636 ( .A(n15721), .B(n14314), .Z(n15722) );
  INV_X1 U17637 ( .A(n15722), .ZN(n14320) );
  INV_X1 U17638 ( .A(n15556), .ZN(n14316) );
  AOI22_X1 U17639 ( .A1(n19938), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B1(
        n13009), .B2(P1_REIP_REG_19__SCAN_IN), .ZN(n14315) );
  OAI21_X1 U17640 ( .B1(n15701), .B2(n14316), .A(n14315), .ZN(n14317) );
  AOI21_X1 U17641 ( .B1(n14318), .B2(n9727), .A(n14317), .ZN(n14319) );
  OAI21_X1 U17642 ( .B1(n14320), .B2(n19764), .A(n14319), .ZN(P1_U2980) );
  OAI21_X1 U17643 ( .B1(n14323), .B2(n14322), .A(n14321), .ZN(n14475) );
  NOR2_X1 U17644 ( .A1(n19845), .A2(n20627), .ZN(n14469) );
  AOI21_X1 U17645 ( .B1(n19938), .B2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n14469), .ZN(n14324) );
  OAI21_X1 U17646 ( .B1(n15701), .B2(n15566), .A(n14324), .ZN(n14325) );
  AOI21_X1 U17647 ( .B1(n15563), .B2(n9727), .A(n14325), .ZN(n14326) );
  OAI21_X1 U17648 ( .B1(n19764), .B2(n14475), .A(n14326), .ZN(P1_U2981) );
  INV_X1 U17649 ( .A(n15677), .ZN(n14352) );
  INV_X1 U17650 ( .A(n14350), .ZN(n14327) );
  AOI21_X1 U17651 ( .B1(n14327), .B2(n14203), .A(n9749), .ZN(n14328) );
  NOR2_X1 U17652 ( .A1(n14352), .A2(n14328), .ZN(n14479) );
  AOI21_X1 U17653 ( .B1(n14479), .B2(n14329), .A(n9808), .ZN(n14331) );
  NOR2_X1 U17654 ( .A1(n14331), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n14330) );
  MUX2_X1 U17655 ( .A(n14331), .B(n14330), .S(n14354), .Z(n14332) );
  XNOR2_X1 U17656 ( .A(n14332), .B(n13911), .ZN(n15729) );
  NAND2_X1 U17657 ( .A1(n15729), .A2(n19944), .ZN(n14337) );
  INV_X1 U17658 ( .A(P1_REIP_REG_17__SCAN_IN), .ZN(n14333) );
  OAI22_X1 U17659 ( .A1(n14334), .A2(n15568), .B1(n19845), .B2(n14333), .ZN(
        n14335) );
  AOI21_X1 U17660 ( .B1(n15672), .B2(n15570), .A(n14335), .ZN(n14336) );
  OAI211_X1 U17661 ( .C1(n20005), .C2(n15571), .A(n14337), .B(n14336), .ZN(
        P1_U2982) );
  NOR2_X1 U17662 ( .A1(n15677), .A2(n14338), .ZN(n15658) );
  INV_X1 U17663 ( .A(n15658), .ZN(n14340) );
  NAND2_X1 U17664 ( .A1(n14340), .A2(n14339), .ZN(n14343) );
  NAND2_X1 U17665 ( .A1(n14341), .A2(n15656), .ZN(n14342) );
  XNOR2_X1 U17666 ( .A(n14343), .B(n14342), .ZN(n15747) );
  INV_X1 U17667 ( .A(n15747), .ZN(n14349) );
  AOI22_X1 U17668 ( .A1(n19938), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B1(
        n13009), .B2(P1_REIP_REG_15__SCAN_IN), .ZN(n14344) );
  OAI21_X1 U17669 ( .B1(n15701), .B2(n14345), .A(n14344), .ZN(n14346) );
  AOI21_X1 U17670 ( .B1(n14347), .B2(n9727), .A(n14346), .ZN(n14348) );
  OAI21_X1 U17671 ( .B1(n14349), .B2(n19764), .A(n14348), .ZN(P1_U2984) );
  AOI22_X1 U17672 ( .A1(n14352), .A2(n14351), .B1(n14354), .B2(n14350), .ZN(
        n14489) );
  INV_X1 U17673 ( .A(n14355), .ZN(n14353) );
  AOI21_X1 U17674 ( .B1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n14354), .A(
        n14353), .ZN(n14488) );
  NAND2_X1 U17675 ( .A1(n14489), .A2(n14488), .ZN(n14487) );
  NAND2_X1 U17676 ( .A1(n14487), .A2(n14355), .ZN(n14356) );
  XOR2_X1 U17677 ( .A(n14357), .B(n14356), .Z(n15754) );
  INV_X1 U17678 ( .A(n15754), .ZN(n14363) );
  AOI22_X1 U17679 ( .A1(n19938), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .B1(
        n13009), .B2(P1_REIP_REG_13__SCAN_IN), .ZN(n14358) );
  OAI21_X1 U17680 ( .B1(n15701), .B2(n14359), .A(n14358), .ZN(n14360) );
  AOI21_X1 U17681 ( .B1(n14361), .B2(n9727), .A(n14360), .ZN(n14362) );
  OAI21_X1 U17682 ( .B1(n14363), .B2(n19764), .A(n14362), .ZN(P1_U2986) );
  MUX2_X1 U17683 ( .A(n15676), .B(n15677), .S(n9749), .Z(n14364) );
  XNOR2_X1 U17684 ( .A(n14364), .B(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n15769) );
  INV_X1 U17685 ( .A(n15769), .ZN(n14368) );
  AOI22_X1 U17686 ( .A1(n19938), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .B1(
        n13009), .B2(P1_REIP_REG_10__SCAN_IN), .ZN(n14365) );
  OAI21_X1 U17687 ( .B1(n15701), .B2(n15623), .A(n14365), .ZN(n14366) );
  AOI21_X1 U17688 ( .B1(n15625), .B2(n9727), .A(n14366), .ZN(n14367) );
  OAI21_X1 U17689 ( .B1(n14368), .B2(n19764), .A(n14367), .ZN(P1_U2989) );
  INV_X1 U17690 ( .A(n19988), .ZN(n14468) );
  NOR2_X1 U17691 ( .A1(n15497), .A2(n15721), .ZN(n14374) );
  NOR3_X1 U17692 ( .A1(n15801), .A2(n19969), .A3(n19948), .ZN(n14493) );
  NOR3_X1 U17693 ( .A1(n14209), .A2(n13403), .A3(n14369), .ZN(n14492) );
  NAND2_X1 U17694 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n14492), .ZN(
        n14497) );
  NOR2_X1 U17695 ( .A1(n14203), .A2(n14497), .ZN(n14371) );
  NAND2_X1 U17696 ( .A1(n14493), .A2(n14371), .ZN(n15750) );
  INV_X1 U17697 ( .A(n15750), .ZN(n15468) );
  NAND2_X1 U17698 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15735) );
  NOR3_X1 U17699 ( .A1(n15734), .A2(n13911), .A3(n15735), .ZN(n14471) );
  NAND2_X1 U17700 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n14471), .ZN(
        n14370) );
  NOR2_X1 U17701 ( .A1(n20819), .A2(n14370), .ZN(n15473) );
  NAND2_X1 U17702 ( .A1(n15468), .A2(n15473), .ZN(n15474) );
  INV_X1 U17703 ( .A(n14370), .ZN(n14386) );
  NAND2_X1 U17704 ( .A1(n14371), .A2(n14494), .ZN(n14384) );
  NOR2_X1 U17705 ( .A1(n20819), .A2(n14384), .ZN(n14482) );
  AOI21_X1 U17706 ( .B1(n14386), .B2(n14482), .A(n19985), .ZN(n14372) );
  NAND2_X1 U17707 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15714) );
  NOR2_X1 U17708 ( .A1(n19985), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14375) );
  NOR2_X1 U17709 ( .A1(n15702), .A2(n14375), .ZN(n14460) );
  NAND2_X1 U17710 ( .A1(n19996), .A2(n14376), .ZN(n14378) );
  NAND2_X1 U17711 ( .A1(n19998), .A2(n14430), .ZN(n14377) );
  OAI211_X1 U17712 ( .C1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n15472), .A(
        n14378), .B(n14377), .ZN(n14379) );
  INV_X1 U17713 ( .A(n14379), .ZN(n14380) );
  INV_X1 U17714 ( .A(n14450), .ZN(n14439) );
  NAND2_X1 U17715 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14381) );
  AOI211_X1 U17716 ( .C1(n14468), .C2(n14439), .A(n12562), .B(n14396), .ZN(
        n14393) );
  NOR2_X1 U17717 ( .A1(n14382), .A2(n15807), .ZN(n14392) );
  INV_X1 U17718 ( .A(n14496), .ZN(n19961) );
  NAND2_X1 U17719 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n15468), .ZN(
        n14467) );
  INV_X1 U17720 ( .A(n14467), .ZN(n14383) );
  NAND2_X1 U17721 ( .A1(n19961), .A2(n14383), .ZN(n14461) );
  NOR2_X1 U17722 ( .A1(n19985), .A2(n14384), .ZN(n15469) );
  NAND2_X1 U17723 ( .A1(n15469), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n14385) );
  AND2_X1 U17724 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n14386), .ZN(
        n14387) );
  NAND4_X1 U17725 ( .A1(n14387), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A4(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n14388) );
  INV_X1 U17726 ( .A(n15703), .ZN(n14456) );
  NOR3_X1 U17727 ( .A1(n14456), .A2(n14430), .A3(n14438), .ZN(n14423) );
  NAND2_X1 U17728 ( .A1(n14423), .A2(n14389), .ZN(n14403) );
  NOR4_X1 U17729 ( .A1(n14403), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n14397), .A4(n14221), .ZN(n14390) );
  NOR4_X1 U17730 ( .A1(n14393), .A2(n14392), .A3(n14391), .A4(n14390), .ZN(
        n14394) );
  OAI21_X1 U17731 ( .B1(n14395), .B2(n19964), .A(n14394), .ZN(P1_U3000) );
  INV_X1 U17732 ( .A(n14396), .ZN(n14401) );
  OAI21_X1 U17733 ( .B1(n14403), .B2(n14221), .A(n14397), .ZN(n14400) );
  INV_X1 U17734 ( .A(n14403), .ZN(n14405) );
  AOI21_X1 U17735 ( .B1(n14405), .B2(n14221), .A(n14404), .ZN(n14406) );
  OAI21_X1 U17736 ( .B1(n14407), .B2(n15807), .A(n14406), .ZN(n14408) );
  AOI21_X1 U17737 ( .B1(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n14409), .A(
        n14408), .ZN(n14410) );
  OAI21_X1 U17738 ( .B1(n14411), .B2(n19964), .A(n14410), .ZN(P1_U3002) );
  INV_X1 U17739 ( .A(n14412), .ZN(n14427) );
  INV_X1 U17740 ( .A(n14413), .ZN(n14417) );
  XNOR2_X1 U17741 ( .A(n14422), .B(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14415) );
  AOI21_X1 U17742 ( .B1(n14423), .B2(n14415), .A(n14414), .ZN(n14416) );
  OAI21_X1 U17743 ( .B1(n14417), .B2(n15807), .A(n14416), .ZN(n14418) );
  AOI21_X1 U17744 ( .B1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n14427), .A(
        n14418), .ZN(n14419) );
  OAI21_X1 U17745 ( .B1(n14420), .B2(n19964), .A(n14419), .ZN(P1_U3003) );
  AOI21_X1 U17746 ( .B1(n14423), .B2(n14422), .A(n14421), .ZN(n14424) );
  OAI21_X1 U17747 ( .B1(n14425), .B2(n15807), .A(n14424), .ZN(n14426) );
  AOI21_X1 U17748 ( .B1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n14427), .A(
        n14426), .ZN(n14428) );
  OAI21_X1 U17749 ( .B1(n14429), .B2(n19964), .A(n14428), .ZN(P1_U3004) );
  NOR2_X1 U17750 ( .A1(n14430), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14432) );
  AOI21_X1 U17751 ( .B1(n15703), .B2(n14432), .A(n14431), .ZN(n14433) );
  OAI21_X1 U17752 ( .B1(n14434), .B2(n15807), .A(n14433), .ZN(n14441) );
  AND2_X1 U17753 ( .A1(n14436), .A2(n14435), .ZN(n14437) );
  NAND2_X1 U17754 ( .A1(n15703), .A2(n14437), .ZN(n14446) );
  AOI21_X1 U17755 ( .B1(n14439), .B2(n14446), .A(n14438), .ZN(n14440) );
  NOR2_X1 U17756 ( .A1(n14441), .A2(n14440), .ZN(n14442) );
  OAI21_X1 U17757 ( .B1(n14443), .B2(n19964), .A(n14442), .ZN(P1_U3005) );
  INV_X1 U17758 ( .A(n14444), .ZN(n14445) );
  OAI211_X1 U17759 ( .C1(n14447), .C2(n15807), .A(n14446), .B(n14445), .ZN(
        n14449) );
  AOI21_X1 U17760 ( .B1(n10107), .B2(n14453), .A(n14452), .ZN(n14455) );
  OR2_X1 U17761 ( .A1(n14455), .A2(n14454), .ZN(n15630) );
  INV_X1 U17762 ( .A(n15630), .ZN(n14459) );
  NOR3_X1 U17763 ( .A1(n14456), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(
        n15709), .ZN(n14457) );
  AOI211_X1 U17764 ( .C1(n14459), .C2(n19993), .A(n14458), .B(n14457), .ZN(
        n14464) );
  OAI21_X1 U17765 ( .B1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n14461), .A(
        n14460), .ZN(n14462) );
  NAND2_X1 U17766 ( .A1(n14462), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14463) );
  OAI211_X1 U17767 ( .C1(n14465), .C2(n19964), .A(n14464), .B(n14463), .ZN(
        P1_U3007) );
  OAI21_X1 U17768 ( .B1(n14482), .B2(n19985), .A(n19984), .ZN(n14466) );
  AOI21_X1 U17769 ( .B1(n19963), .B2(n14467), .A(n14466), .ZN(n15733) );
  OAI21_X1 U17770 ( .B1(n14468), .B2(n14471), .A(n15733), .ZN(n15727) );
  NOR2_X1 U17771 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n15726), .ZN(
        n14470) );
  AOI21_X1 U17772 ( .B1(n14471), .B2(n14470), .A(n14469), .ZN(n14472) );
  OAI21_X1 U17773 ( .B1(n15561), .B2(n15807), .A(n14472), .ZN(n14473) );
  AOI21_X1 U17774 ( .B1(n15727), .B2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n14473), .ZN(n14474) );
  OAI21_X1 U17775 ( .B1(n14475), .B2(n19964), .A(n14474), .ZN(P1_U3013) );
  INV_X1 U17776 ( .A(n14476), .ZN(n14478) );
  OAI21_X1 U17777 ( .B1(n14479), .B2(n14478), .A(n14477), .ZN(n14481) );
  XNOR2_X1 U17778 ( .A(n9749), .B(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n14480) );
  XNOR2_X1 U17779 ( .A(n14481), .B(n14480), .ZN(n15669) );
  INV_X1 U17780 ( .A(P1_REIP_REG_14__SCAN_IN), .ZN(n20824) );
  OAI22_X1 U17781 ( .A1(n15733), .A2(n15734), .B1(n19845), .B2(n20824), .ZN(
        n14485) );
  NAND3_X1 U17782 ( .A1(n14482), .A2(n15734), .A3(n15798), .ZN(n14483) );
  OAI21_X1 U17783 ( .B1(n15807), .B2(n15594), .A(n14483), .ZN(n14484) );
  NOR2_X1 U17784 ( .A1(n14485), .A2(n14484), .ZN(n14486) );
  OAI21_X1 U17785 ( .B1(n15669), .B2(n19964), .A(n14486), .ZN(P1_U3017) );
  OAI21_X1 U17786 ( .B1(n14489), .B2(n14488), .A(n14487), .ZN(n14490) );
  INV_X1 U17787 ( .A(n14490), .ZN(n15675) );
  NAND2_X1 U17788 ( .A1(n14492), .A2(n14210), .ZN(n15760) );
  AOI21_X1 U17789 ( .B1(n14493), .B2(n14492), .A(n14491), .ZN(n14495) );
  OAI21_X1 U17790 ( .B1(n14494), .B2(n19985), .A(n19984), .ZN(n15774) );
  AOI211_X1 U17791 ( .C1(n19971), .C2(n14497), .A(n14495), .B(n15774), .ZN(
        n15761) );
  OAI21_X1 U17792 ( .B1(n14496), .B2(n15760), .A(n15761), .ZN(n14499) );
  OAI21_X1 U17793 ( .B1(n14497), .B2(n15796), .A(n14203), .ZN(n14498) );
  OAI21_X1 U17794 ( .B1(n14203), .B2(n14499), .A(n14498), .ZN(n14506) );
  NAND2_X1 U17795 ( .A1(n14501), .A2(n14500), .ZN(n14502) );
  NAND2_X1 U17796 ( .A1(n14503), .A2(n14502), .ZN(n15604) );
  OAI22_X1 U17797 ( .A1(n15604), .A2(n15807), .B1(n19845), .B2(n20617), .ZN(
        n14504) );
  INV_X1 U17798 ( .A(n14504), .ZN(n14505) );
  OAI211_X1 U17799 ( .C1(n15675), .C2(n19964), .A(n14506), .B(n14505), .ZN(
        P1_U3019) );
  MUX2_X1 U17800 ( .A(n20517), .B(n14507), .S(n20008), .Z(n14508) );
  OAI21_X1 U17801 ( .B1(n14509), .B2(n9754), .A(n14508), .ZN(n14510) );
  MUX2_X1 U17802 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n14510), .S(
        n20002), .Z(P1_U3476) );
  NOR3_X1 U17803 ( .A1(n12341), .A2(n14516), .A3(n14515), .ZN(n14511) );
  AOI211_X1 U17804 ( .C1(n20465), .C2(n14513), .A(n14512), .B(n14511), .ZN(
        n15431) );
  INV_X1 U17805 ( .A(n14514), .ZN(n14519) );
  NOR3_X1 U17806 ( .A1(n14516), .A2(n14515), .A3(n14524), .ZN(n14517) );
  AOI21_X1 U17807 ( .B1(n14519), .B2(n14518), .A(n14517), .ZN(n14520) );
  OAI21_X1 U17808 ( .B1(n15431), .B2(n14526), .A(n14520), .ZN(n14522) );
  INV_X1 U17809 ( .A(n14521), .ZN(n15814) );
  MUX2_X1 U17810 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n14522), .S(
        n15814), .Z(P1_U3473) );
  INV_X1 U17811 ( .A(n14523), .ZN(n14527) );
  OAI22_X1 U17812 ( .A1(n14527), .A2(n14526), .B1(n14525), .B2(n14524), .ZN(
        n14528) );
  MUX2_X1 U17813 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n14528), .S(
        n15814), .Z(P1_U3469) );
  INV_X1 U17814 ( .A(n15841), .ZN(n14529) );
  NAND2_X1 U17815 ( .A1(n14529), .A2(n14582), .ZN(n14530) );
  OAI21_X1 U17816 ( .B1(n14621), .B2(n15830), .A(n14530), .ZN(P2_U2856) );
  OAI21_X1 U17817 ( .B1(n14545), .B2(n14532), .A(n14531), .ZN(n15862) );
  OR2_X1 U17818 ( .A1(n14534), .A2(n14533), .ZN(n14631) );
  NAND3_X1 U17819 ( .A1(n14631), .A2(n14535), .A3(n14601), .ZN(n14537) );
  NAND2_X1 U17820 ( .A1(n14602), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n14536) );
  OAI211_X1 U17821 ( .C1(n14602), .C2(n15862), .A(n14537), .B(n14536), .ZN(
        P2_U2858) );
  NOR2_X1 U17822 ( .A1(n14539), .A2(n14538), .ZN(n14541) );
  XNOR2_X1 U17823 ( .A(n14541), .B(n14540), .ZN(n14647) );
  NAND2_X1 U17824 ( .A1(n14602), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n14547) );
  NOR2_X1 U17825 ( .A1(n14543), .A2(n14542), .ZN(n14544) );
  NOR2_X1 U17826 ( .A1(n14545), .A2(n14544), .ZN(n15865) );
  NAND2_X1 U17827 ( .A1(n15865), .A2(n14582), .ZN(n14546) );
  OAI211_X1 U17828 ( .C1(n14647), .C2(n14630), .A(n14547), .B(n14546), .ZN(
        P2_U2859) );
  OAI21_X1 U17829 ( .B1(n14550), .B2(n14549), .A(n14548), .ZN(n14655) );
  XNOR2_X1 U17830 ( .A(n14560), .B(n14551), .ZN(n15884) );
  NOR2_X1 U17831 ( .A1(n15884), .A2(n14602), .ZN(n14552) );
  AOI21_X1 U17832 ( .B1(P2_EBX_REG_27__SCAN_IN), .B2(n14602), .A(n14552), .ZN(
        n14553) );
  OAI21_X1 U17833 ( .B1(n14655), .B2(n14630), .A(n14553), .ZN(P2_U2860) );
  OAI21_X1 U17834 ( .B1(n14556), .B2(n14555), .A(n14554), .ZN(n14663) );
  NAND2_X1 U17835 ( .A1(n14602), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n14562) );
  NOR2_X1 U17836 ( .A1(n14557), .A2(n14558), .ZN(n14559) );
  NOR2_X1 U17837 ( .A1(n14560), .A2(n14559), .ZN(n15889) );
  NAND2_X1 U17838 ( .A1(n15889), .A2(n14582), .ZN(n14561) );
  OAI211_X1 U17839 ( .C1(n14663), .C2(n14630), .A(n14562), .B(n14561), .ZN(
        P2_U2861) );
  OAI21_X1 U17840 ( .B1(n14565), .B2(n14564), .A(n14563), .ZN(n14669) );
  INV_X1 U17841 ( .A(n14557), .ZN(n14570) );
  INV_X1 U17842 ( .A(n14580), .ZN(n14568) );
  INV_X1 U17843 ( .A(n14566), .ZN(n14567) );
  NAND2_X1 U17844 ( .A1(n14568), .A2(n14567), .ZN(n14569) );
  NAND2_X1 U17845 ( .A1(n14570), .A2(n14569), .ZN(n15934) );
  MUX2_X1 U17846 ( .A(n14571), .B(n15934), .S(n14582), .Z(n14572) );
  OAI21_X1 U17847 ( .B1(n14669), .B2(n14630), .A(n14572), .ZN(P2_U2862) );
  AOI21_X1 U17848 ( .B1(n14575), .B2(n14574), .A(n14573), .ZN(n14576) );
  XOR2_X1 U17849 ( .A(n14577), .B(n14576), .Z(n14677) );
  NAND2_X1 U17850 ( .A1(n14602), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n14584) );
  INV_X1 U17851 ( .A(n14578), .ZN(n14581) );
  INV_X1 U17852 ( .A(n14579), .ZN(n14586) );
  AOI21_X1 U17853 ( .B1(n14581), .B2(n14586), .A(n14580), .ZN(n15945) );
  NAND2_X1 U17854 ( .A1(n15945), .A2(n14582), .ZN(n14583) );
  OAI211_X1 U17855 ( .C1(n14677), .C2(n14630), .A(n14584), .B(n14583), .ZN(
        P2_U2863) );
  OAI21_X1 U17856 ( .B1(n14585), .B2(n14587), .A(n14586), .ZN(n16068) );
  AOI21_X1 U17857 ( .B1(n14590), .B2(n14589), .A(n14588), .ZN(n15929) );
  NAND2_X1 U17858 ( .A1(n15929), .A2(n14601), .ZN(n14592) );
  NAND2_X1 U17859 ( .A1(n14602), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n14591) );
  OAI211_X1 U17860 ( .C1(n16068), .C2(n14602), .A(n14592), .B(n14591), .ZN(
        P2_U2864) );
  INV_X1 U17861 ( .A(n14585), .ZN(n14597) );
  INV_X1 U17862 ( .A(n14593), .ZN(n14610) );
  INV_X1 U17863 ( .A(n14594), .ZN(n14595) );
  NAND2_X1 U17864 ( .A1(n14610), .A2(n14595), .ZN(n14596) );
  NAND2_X1 U17865 ( .A1(n14597), .A2(n14596), .ZN(n15966) );
  AOI21_X1 U17866 ( .B1(n14600), .B2(n14598), .A(n14599), .ZN(n14678) );
  NAND2_X1 U17867 ( .A1(n14678), .A2(n14601), .ZN(n14604) );
  NAND2_X1 U17868 ( .A1(n14602), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n14603) );
  OAI211_X1 U17869 ( .C1(n15966), .C2(n14602), .A(n14604), .B(n14603), .ZN(
        P2_U2865) );
  OAI21_X1 U17870 ( .B1(n14612), .B2(n14605), .A(n14598), .ZN(n14695) );
  INV_X1 U17871 ( .A(n14619), .ZN(n14608) );
  INV_X1 U17872 ( .A(n14606), .ZN(n14607) );
  NAND2_X1 U17873 ( .A1(n14608), .A2(n14607), .ZN(n14609) );
  NAND2_X1 U17874 ( .A1(n14610), .A2(n14609), .ZN(n18706) );
  MUX2_X1 U17875 ( .A(n11346), .B(n18706), .S(n14582), .Z(n14611) );
  OAI21_X1 U17876 ( .B1(n14695), .B2(n14630), .A(n14611), .ZN(P2_U2866) );
  AOI21_X1 U17877 ( .B1(n14614), .B2(n14613), .A(n14612), .ZN(n14615) );
  INV_X1 U17878 ( .A(n14615), .ZN(n14703) );
  NOR2_X1 U17879 ( .A1(n14617), .A2(n14616), .ZN(n14618) );
  NOR2_X1 U17880 ( .A1(n14619), .A2(n14618), .ZN(n18710) );
  NOR2_X1 U17881 ( .A1(n14582), .A2(n11345), .ZN(n14620) );
  AOI21_X1 U17882 ( .B1(n18710), .B2(n14621), .A(n14620), .ZN(n14622) );
  OAI21_X1 U17883 ( .B1(n14703), .B2(n14630), .A(n14622), .ZN(P2_U2867) );
  NOR2_X1 U17884 ( .A1(n14624), .A2(n14623), .ZN(n14625) );
  NOR2_X1 U17885 ( .A1(n14626), .A2(n14625), .ZN(n18734) );
  INV_X1 U17886 ( .A(n18734), .ZN(n14816) );
  MUX2_X1 U17887 ( .A(n14627), .B(n14816), .S(n14582), .Z(n14628) );
  OAI21_X1 U17888 ( .B1(n14630), .B2(n14629), .A(n14628), .ZN(P2_U2869) );
  NAND3_X1 U17889 ( .A1(n14631), .A2(n14535), .A3(n15928), .ZN(n14638) );
  AOI21_X1 U17890 ( .B1(n14633), .B2(n14639), .A(n14632), .ZN(n15856) );
  AOI22_X1 U17891 ( .A1(n15856), .A2(n18930), .B1(n18934), .B2(
        P2_EAX_REG_29__SCAN_IN), .ZN(n14637) );
  AOI22_X1 U17892 ( .A1(n18929), .A2(BUF2_REG_29__SCAN_IN), .B1(n18931), .B2(
        BUF1_REG_29__SCAN_IN), .ZN(n14636) );
  MUX2_X1 U17893 ( .A(BUF1_REG_13__SCAN_IN), .B(BUF2_REG_13__SCAN_IN), .S(
        n14634), .Z(n19021) );
  NAND2_X1 U17894 ( .A1(n15927), .A2(n19021), .ZN(n14635) );
  NAND4_X1 U17895 ( .A1(n14638), .A2(n14637), .A3(n14636), .A4(n14635), .ZN(
        P2_U2890) );
  INV_X1 U17896 ( .A(n14639), .ZN(n14640) );
  AOI21_X1 U17897 ( .B1(n14641), .B2(n14648), .A(n14640), .ZN(n15864) );
  INV_X1 U17898 ( .A(n15864), .ZN(n14642) );
  INV_X1 U17899 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n18964) );
  OAI22_X1 U17900 ( .A1(n14642), .A2(n14709), .B1(n18948), .B2(n18964), .ZN(
        n14643) );
  AOI21_X1 U17901 ( .B1(n15927), .B2(n14644), .A(n14643), .ZN(n14646) );
  AOI22_X1 U17902 ( .A1(n18929), .A2(BUF2_REG_28__SCAN_IN), .B1(n18931), .B2(
        BUF1_REG_28__SCAN_IN), .ZN(n14645) );
  OAI211_X1 U17903 ( .C1(n14647), .C2(n14714), .A(n14646), .B(n14645), .ZN(
        P2_U2891) );
  INV_X1 U17904 ( .A(n14648), .ZN(n14649) );
  AOI21_X1 U17905 ( .B1(n14650), .B2(n14658), .A(n14649), .ZN(n15878) );
  INV_X1 U17906 ( .A(n15878), .ZN(n14651) );
  OAI22_X1 U17907 ( .A1(n14651), .A2(n14709), .B1(n18948), .B2(n18966), .ZN(
        n14652) );
  AOI21_X1 U17908 ( .B1(n15927), .B2(n18941), .A(n14652), .ZN(n14654) );
  AOI22_X1 U17909 ( .A1(n18929), .A2(BUF2_REG_27__SCAN_IN), .B1(n18931), .B2(
        BUF1_REG_27__SCAN_IN), .ZN(n14653) );
  OAI211_X1 U17910 ( .C1(n14655), .C2(n14714), .A(n14654), .B(n14653), .ZN(
        P2_U2892) );
  OR2_X1 U17911 ( .A1(n9795), .A2(n14656), .ZN(n14657) );
  NAND2_X1 U17912 ( .A1(n14658), .A2(n14657), .ZN(n15895) );
  INV_X1 U17913 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n18968) );
  OAI22_X1 U17914 ( .A1(n14709), .A2(n15895), .B1(n18948), .B2(n18968), .ZN(
        n14659) );
  AOI21_X1 U17915 ( .B1(n15927), .B2(n14660), .A(n14659), .ZN(n14662) );
  AOI22_X1 U17916 ( .A1(n18929), .A2(BUF2_REG_26__SCAN_IN), .B1(n18931), .B2(
        BUF1_REG_26__SCAN_IN), .ZN(n14661) );
  OAI211_X1 U17917 ( .C1(n14663), .C2(n14714), .A(n14662), .B(n14661), .ZN(
        P2_U2893) );
  AND2_X1 U17918 ( .A1(n14672), .A2(n14664), .ZN(n14665) );
  NOR2_X1 U17919 ( .A1(n9795), .A2(n14665), .ZN(n15899) );
  INV_X1 U17920 ( .A(n15899), .ZN(n14932) );
  OAI22_X1 U17921 ( .A1(n14709), .A2(n14932), .B1(n18948), .B2(n18970), .ZN(
        n14666) );
  AOI21_X1 U17922 ( .B1(n15927), .B2(n18945), .A(n14666), .ZN(n14668) );
  AOI22_X1 U17923 ( .A1(n18929), .A2(BUF2_REG_25__SCAN_IN), .B1(n18931), .B2(
        BUF1_REG_25__SCAN_IN), .ZN(n14667) );
  OAI211_X1 U17924 ( .C1(n14669), .C2(n14714), .A(n14668), .B(n14667), .ZN(
        P2_U2894) );
  NAND2_X1 U17925 ( .A1(n15915), .A2(n14670), .ZN(n14671) );
  NAND2_X1 U17926 ( .A1(n14672), .A2(n14671), .ZN(n15913) );
  INV_X1 U17927 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n18972) );
  OAI22_X1 U17928 ( .A1(n14709), .A2(n15913), .B1(n18948), .B2(n18972), .ZN(
        n14673) );
  AOI21_X1 U17929 ( .B1(n15927), .B2(n14674), .A(n14673), .ZN(n14676) );
  AOI22_X1 U17930 ( .A1(n18929), .A2(BUF2_REG_24__SCAN_IN), .B1(n18931), .B2(
        BUF1_REG_24__SCAN_IN), .ZN(n14675) );
  OAI211_X1 U17931 ( .C1(n14677), .C2(n14714), .A(n14676), .B(n14675), .ZN(
        P2_U2895) );
  INV_X1 U17932 ( .A(n14678), .ZN(n14687) );
  NOR2_X1 U17933 ( .A1(n14681), .A2(n14680), .ZN(n14682) );
  OR2_X1 U17934 ( .A1(n14679), .A2(n14682), .ZN(n15392) );
  INV_X1 U17935 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n18975) );
  OAI22_X1 U17936 ( .A1(n14709), .A2(n15392), .B1(n18975), .B2(n18948), .ZN(
        n14683) );
  AOI21_X1 U17937 ( .B1(n15927), .B2(n14684), .A(n14683), .ZN(n14686) );
  AOI22_X1 U17938 ( .A1(n18929), .A2(BUF2_REG_22__SCAN_IN), .B1(n18931), .B2(
        BUF1_REG_22__SCAN_IN), .ZN(n14685) );
  OAI211_X1 U17939 ( .C1(n14687), .C2(n14714), .A(n14686), .B(n14685), .ZN(
        P2_U2897) );
  INV_X1 U17940 ( .A(n14688), .ZN(n14689) );
  XNOR2_X1 U17941 ( .A(n14698), .B(n14689), .ZN(n18700) );
  INV_X1 U17942 ( .A(n18700), .ZN(n14690) );
  INV_X1 U17943 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n18977) );
  OAI22_X1 U17944 ( .A1(n14709), .A2(n14690), .B1(n18977), .B2(n18948), .ZN(
        n14691) );
  AOI21_X1 U17945 ( .B1(n15927), .B2(n14692), .A(n14691), .ZN(n14694) );
  AOI22_X1 U17946 ( .A1(n18929), .A2(BUF2_REG_21__SCAN_IN), .B1(n18931), .B2(
        BUF1_REG_21__SCAN_IN), .ZN(n14693) );
  OAI211_X1 U17947 ( .C1(n14695), .C2(n14714), .A(n14694), .B(n14693), .ZN(
        P2_U2898) );
  NAND2_X1 U17948 ( .A1(n14705), .A2(n14696), .ZN(n14697) );
  NAND2_X1 U17949 ( .A1(n14698), .A2(n14697), .ZN(n18708) );
  INV_X1 U17950 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n18979) );
  OAI22_X1 U17951 ( .A1(n14709), .A2(n18708), .B1(n18979), .B2(n18948), .ZN(
        n14699) );
  AOI21_X1 U17952 ( .B1(n15927), .B2(n14700), .A(n14699), .ZN(n14702) );
  AOI22_X1 U17953 ( .A1(n18929), .A2(BUF2_REG_20__SCAN_IN), .B1(n18931), .B2(
        BUF1_REG_20__SCAN_IN), .ZN(n14701) );
  OAI211_X1 U17954 ( .C1(n14703), .C2(n14714), .A(n14702), .B(n14701), .ZN(
        P2_U2899) );
  INV_X1 U17955 ( .A(n14705), .ZN(n14706) );
  AOI21_X1 U17956 ( .B1(n10148), .B2(n14707), .A(n14706), .ZN(n18721) );
  INV_X1 U17957 ( .A(n18721), .ZN(n14708) );
  INV_X1 U17958 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n18981) );
  OAI22_X1 U17959 ( .A1(n14709), .A2(n14708), .B1(n18981), .B2(n18948), .ZN(
        n14710) );
  AOI21_X1 U17960 ( .B1(n15927), .B2(n14711), .A(n14710), .ZN(n14713) );
  AOI22_X1 U17961 ( .A1(n18929), .A2(BUF2_REG_19__SCAN_IN), .B1(n18931), .B2(
        BUF1_REG_19__SCAN_IN), .ZN(n14712) );
  OAI211_X1 U17962 ( .C1(n14715), .C2(n14714), .A(n14713), .B(n14712), .ZN(
        P2_U2900) );
  XNOR2_X1 U17963 ( .A(n14716), .B(n14717), .ZN(n14878) );
  INV_X1 U17964 ( .A(n14718), .ZN(n14720) );
  NAND2_X1 U17965 ( .A1(n14720), .A2(n14719), .ZN(n14721) );
  XNOR2_X1 U17966 ( .A(n14722), .B(n14721), .ZN(n14876) );
  NOR2_X1 U17967 ( .A1(n18846), .A2(n19670), .ZN(n14869) );
  XNOR2_X1 U17968 ( .A(n14734), .B(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15846) );
  NOR2_X1 U17969 ( .A1(n19045), .A2(n15846), .ZN(n14723) );
  AOI211_X1 U17970 ( .C1(n19032), .C2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n14869), .B(n14723), .ZN(n14724) );
  OAI21_X1 U17971 ( .B1(n14874), .B2(n16058), .A(n14724), .ZN(n14725) );
  AOI21_X1 U17972 ( .B1(n14876), .B2(n16060), .A(n14725), .ZN(n14726) );
  OAI21_X1 U17973 ( .B1(n19035), .B2(n14878), .A(n14726), .ZN(P2_U2984) );
  OAI21_X1 U17974 ( .B1(n14727), .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n14716), .ZN(n14890) );
  INV_X1 U17975 ( .A(n14728), .ZN(n14729) );
  NOR2_X1 U17976 ( .A1(n14730), .A2(n14729), .ZN(n14731) );
  XNOR2_X1 U17977 ( .A(n14732), .B(n14731), .ZN(n14888) );
  INV_X1 U17978 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n14733) );
  NOR2_X1 U17979 ( .A1(n18846), .A2(n14733), .ZN(n14880) );
  AOI21_X1 U17980 ( .B1(n19032), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n14880), .ZN(n14736) );
  AOI21_X1 U17981 ( .B1(n14752), .B2(n11697), .A(n14734), .ZN(n15838) );
  NAND2_X1 U17982 ( .A1(n16054), .A2(n15838), .ZN(n14735) );
  OAI211_X1 U17983 ( .C1(n15862), .C2(n16058), .A(n14736), .B(n14735), .ZN(
        n14737) );
  AOI21_X1 U17984 ( .B1(n14888), .B2(n16060), .A(n14737), .ZN(n14738) );
  OAI21_X1 U17985 ( .B1(n19035), .B2(n14890), .A(n14738), .ZN(P2_U2985) );
  INV_X1 U17986 ( .A(n14740), .ZN(n14742) );
  NAND2_X1 U17987 ( .A1(n14742), .A2(n14741), .ZN(n14743) );
  NAND2_X1 U17988 ( .A1(n14744), .A2(n14743), .ZN(n15873) );
  NOR2_X1 U17989 ( .A1(n15873), .A2(n11235), .ZN(n14747) );
  INV_X1 U17990 ( .A(n14745), .ZN(n14746) );
  AOI22_X1 U17991 ( .A1(n14757), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B1(
        n14747), .B2(n14746), .ZN(n14750) );
  XOR2_X1 U17992 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .B(n14748), .Z(
        n14749) );
  XNOR2_X1 U17993 ( .A(n14750), .B(n14749), .ZN(n14900) );
  AOI21_X1 U17994 ( .B1(n14895), .B2(n14751), .A(n14727), .ZN(n14898) );
  OAI21_X1 U17995 ( .B1(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n14758), .A(
        n14752), .ZN(n15868) );
  NAND2_X1 U17996 ( .A1(n15865), .A2(n19041), .ZN(n14754) );
  NOR2_X1 U17997 ( .A1(n18846), .A2(n19664), .ZN(n14892) );
  AOI21_X1 U17998 ( .B1(n19032), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n14892), .ZN(n14753) );
  OAI211_X1 U17999 ( .C1(n15868), .C2(n19045), .A(n14754), .B(n14753), .ZN(
        n14755) );
  AOI21_X1 U18000 ( .B1(n14898), .B2(n16055), .A(n14755), .ZN(n14756) );
  OAI21_X1 U18001 ( .B1(n14900), .B2(n19037), .A(n14756), .ZN(P2_U2986) );
  AOI21_X1 U18002 ( .B1(n14768), .B2(n15874), .A(n14758), .ZN(n15837) );
  NOR2_X1 U18003 ( .A1(n18846), .A2(n14759), .ZN(n14901) );
  AOI21_X1 U18004 ( .B1(n19032), .B2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n14901), .ZN(n14760) );
  OAI21_X1 U18005 ( .B1(n15884), .B2(n16058), .A(n14760), .ZN(n14763) );
  NOR2_X1 U18006 ( .A1(n14906), .A2(n19035), .ZN(n14762) );
  OAI21_X1 U18007 ( .B1(n14909), .B2(n19037), .A(n14764), .ZN(P2_U2987) );
  OAI21_X1 U18008 ( .B1(n14925), .B2(n14923), .A(n14921), .ZN(n14766) );
  XNOR2_X1 U18009 ( .A(n14766), .B(n14765), .ZN(n14919) );
  NOR2_X1 U18010 ( .A1(n14926), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14767) );
  OR2_X1 U18011 ( .A1(n14761), .A2(n14767), .ZN(n14910) );
  AOI22_X1 U18012 ( .A1(n15889), .A2(n19041), .B1(
        P2_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n19032), .ZN(n14771) );
  OAI21_X1 U18013 ( .B1(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n9850), .A(
        n14768), .ZN(n15892) );
  OAI22_X1 U18014 ( .A1(n20880), .A2(n18823), .B1(n19045), .B2(n15892), .ZN(
        n14769) );
  INV_X1 U18015 ( .A(n14769), .ZN(n14770) );
  OAI211_X1 U18016 ( .C1(n14910), .C2(n19035), .A(n14771), .B(n14770), .ZN(
        n14772) );
  AOI21_X1 U18017 ( .B1(n14919), .B2(n16060), .A(n14772), .ZN(n14773) );
  INV_X1 U18018 ( .A(n14773), .ZN(P2_U2988) );
  INV_X1 U18019 ( .A(n14774), .ZN(n15998) );
  NOR2_X1 U18020 ( .A1(n14775), .A2(n15998), .ZN(n14776) );
  NAND2_X1 U18021 ( .A1(n14777), .A2(n14833), .ZN(n15990) );
  INV_X1 U18022 ( .A(n15987), .ZN(n14778) );
  INV_X1 U18023 ( .A(n14779), .ZN(n15988) );
  INV_X1 U18024 ( .A(n14782), .ZN(n14783) );
  OR2_X1 U18025 ( .A1(n14783), .A2(n14784), .ZN(n15418) );
  INV_X1 U18026 ( .A(n14784), .ZN(n14785) );
  INV_X1 U18027 ( .A(n14786), .ZN(n14813) );
  NAND2_X1 U18028 ( .A1(n14815), .A2(n14813), .ZN(n15969) );
  INV_X1 U18029 ( .A(n14787), .ZN(n14788) );
  OAI21_X1 U18030 ( .B1(n15969), .B2(n15971), .A(n14788), .ZN(n14806) );
  INV_X1 U18031 ( .A(n14791), .ZN(n14790) );
  NOR2_X1 U18032 ( .A1(n14790), .A2(n14789), .ZN(n14805) );
  NAND2_X1 U18033 ( .A1(n14806), .A2(n14805), .ZN(n14804) );
  NAND2_X1 U18034 ( .A1(n14804), .A2(n14791), .ZN(n14795) );
  NAND2_X1 U18035 ( .A1(n14793), .A2(n14792), .ZN(n14794) );
  XNOR2_X1 U18036 ( .A(n14795), .B(n14794), .ZN(n14973) );
  AOI21_X1 U18037 ( .B1(n14808), .B2(n18695), .A(n15394), .ZN(n15412) );
  NAND2_X1 U18038 ( .A1(n19033), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n14964) );
  NAND2_X1 U18039 ( .A1(n19032), .A2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n14796) );
  OAI211_X1 U18040 ( .C1(n18706), .C2(n16058), .A(n14964), .B(n14796), .ZN(
        n14800) );
  NAND2_X1 U18041 ( .A1(n14797), .A2(n14966), .ZN(n14798) );
  NAND2_X1 U18042 ( .A1(n14952), .A2(n14798), .ZN(n14970) );
  NOR2_X1 U18043 ( .A1(n14970), .A2(n19035), .ZN(n14799) );
  AOI211_X1 U18044 ( .C1(n16054), .C2(n15412), .A(n14800), .B(n14799), .ZN(
        n14801) );
  OAI21_X1 U18045 ( .B1(n14973), .B2(n19037), .A(n14801), .ZN(P2_U2993) );
  OR2_X1 U18046 ( .A1(n14802), .A2(n11625), .ZN(n15976) );
  INV_X1 U18047 ( .A(n15976), .ZN(n14803) );
  OAI21_X1 U18048 ( .B1(n14803), .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n14797), .ZN(n14983) );
  OAI21_X1 U18049 ( .B1(n14806), .B2(n14805), .A(n14804), .ZN(n14974) );
  NAND2_X1 U18050 ( .A1(n14974), .A2(n16060), .ZN(n14812) );
  NOR2_X1 U18051 ( .A1(n20777), .A2(n18846), .ZN(n14976) );
  AOI21_X1 U18052 ( .B1(n19032), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n14976), .ZN(n14807) );
  INV_X1 U18053 ( .A(n14807), .ZN(n14810) );
  OAI21_X1 U18054 ( .B1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n15410), .A(
        n14808), .ZN(n18713) );
  NOR2_X1 U18055 ( .A1(n19045), .A2(n18713), .ZN(n14809) );
  AOI211_X1 U18056 ( .C1(n19041), .C2(n18710), .A(n14810), .B(n14809), .ZN(
        n14811) );
  OAI211_X1 U18057 ( .C1(n19035), .C2(n14983), .A(n14812), .B(n14811), .ZN(
        P2_U2994) );
  NAND2_X1 U18058 ( .A1(n14813), .A2(n15968), .ZN(n14814) );
  XNOR2_X1 U18059 ( .A(n14815), .B(n14814), .ZN(n14994) );
  OAI21_X1 U18060 ( .B1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n9849), .A(
        n15411), .ZN(n18737) );
  OAI22_X1 U18061 ( .A1(n19650), .A2(n18846), .B1(n19045), .B2(n18737), .ZN(
        n14818) );
  NOR2_X1 U18062 ( .A1(n14816), .A2(n16058), .ZN(n14817) );
  AOI211_X1 U18063 ( .C1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(n19032), .A(
        n14818), .B(n14817), .ZN(n14824) );
  NAND2_X1 U18064 ( .A1(n14819), .A2(n14996), .ZN(n15992) );
  OAI21_X1 U18065 ( .B1(n15981), .B2(n14821), .A(n14989), .ZN(n14822) );
  NAND2_X1 U18066 ( .A1(n14822), .A2(n14802), .ZN(n14990) );
  OR2_X1 U18067 ( .A1(n14990), .A2(n19035), .ZN(n14823) );
  OAI211_X1 U18068 ( .C1(n14994), .C2(n19037), .A(n14824), .B(n14823), .ZN(
        P2_U2996) );
  XNOR2_X1 U18069 ( .A(n14826), .B(n14825), .ZN(n15003) );
  INV_X1 U18070 ( .A(n15003), .ZN(n14831) );
  NOR2_X1 U18071 ( .A1(n19647), .A2(n18823), .ZN(n14828) );
  OAI21_X1 U18072 ( .B1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n15395), .A(
        n15408), .ZN(n18758) );
  OAI22_X1 U18073 ( .A1(n10045), .A2(n16064), .B1(n19045), .B2(n18758), .ZN(
        n14827) );
  AOI211_X1 U18074 ( .C1(n18761), .C2(n19041), .A(n14828), .B(n14827), .ZN(
        n14830) );
  INV_X1 U18075 ( .A(n15005), .ZN(n15991) );
  OAI211_X1 U18076 ( .C1(n15991), .C2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n16055), .B(n15981), .ZN(n14829) );
  OAI211_X1 U18077 ( .C1(n14831), .C2(n19037), .A(n14830), .B(n14829), .ZN(
        P2_U2998) );
  INV_X1 U18078 ( .A(n14832), .ZN(n14834) );
  NAND2_X1 U18079 ( .A1(n14834), .A2(n14833), .ZN(n14835) );
  XNOR2_X1 U18080 ( .A(n14836), .B(n14835), .ZN(n15024) );
  INV_X1 U18081 ( .A(n16015), .ZN(n14837) );
  NAND2_X1 U18082 ( .A1(n14837), .A2(n16103), .ZN(n16001) );
  INV_X1 U18083 ( .A(n15992), .ZN(n14838) );
  AOI21_X1 U18084 ( .B1(n16001), .B2(n14839), .A(n14838), .ZN(n15011) );
  NAND2_X1 U18085 ( .A1(n15011), .A2(n16055), .ZN(n14843) );
  OAI21_X1 U18086 ( .B1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n15397), .A(
        n15396), .ZN(n18781) );
  OAI22_X1 U18087 ( .A1(n11608), .A2(n18823), .B1(n19045), .B2(n18781), .ZN(
        n14841) );
  INV_X1 U18088 ( .A(n18784), .ZN(n15020) );
  NOR2_X1 U18089 ( .A1(n15020), .A2(n16058), .ZN(n14840) );
  AOI211_X1 U18090 ( .C1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .C2(n19032), .A(
        n14841), .B(n14840), .ZN(n14842) );
  OAI211_X1 U18091 ( .C1(n19037), .C2(n15024), .A(n14843), .B(n14842), .ZN(
        P2_U3000) );
  NAND2_X1 U18092 ( .A1(n14845), .A2(n14844), .ZN(n14850) );
  INV_X1 U18093 ( .A(n14846), .ZN(n14848) );
  NAND2_X1 U18094 ( .A1(n14848), .A2(n14847), .ZN(n14849) );
  XOR2_X1 U18095 ( .A(n14850), .B(n14849), .Z(n16115) );
  OAI21_X1 U18096 ( .B1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n9823), .A(
        n15398), .ZN(n18802) );
  OAI22_X1 U18097 ( .A1(n11594), .A2(n18846), .B1(n19045), .B2(n18802), .ZN(
        n14853) );
  NOR2_X1 U18098 ( .A1(n14851), .A2(n16058), .ZN(n14852) );
  AOI211_X1 U18099 ( .C1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .C2(n19032), .A(
        n14853), .B(n14852), .ZN(n14855) );
  NOR2_X1 U18100 ( .A1(n11335), .A2(n16015), .ZN(n16002) );
  AOI21_X1 U18101 ( .B1(n16015), .B2(n11335), .A(n16002), .ZN(n16112) );
  NAND2_X1 U18102 ( .A1(n16112), .A2(n16055), .ZN(n14854) );
  OAI211_X1 U18103 ( .C1(n16115), .C2(n19037), .A(n14855), .B(n14854), .ZN(
        P2_U3002) );
  INV_X1 U18104 ( .A(n14856), .ZN(n15026) );
  NOR2_X1 U18105 ( .A1(n14857), .A2(n15026), .ZN(n14861) );
  NAND2_X1 U18106 ( .A1(n14859), .A2(n14858), .ZN(n14860) );
  XNOR2_X1 U18107 ( .A(n14861), .B(n14860), .ZN(n16140) );
  INV_X1 U18108 ( .A(n16014), .ZN(n14862) );
  AOI21_X1 U18109 ( .B1(n16134), .B2(n15025), .A(n14862), .ZN(n16136) );
  NAND2_X1 U18110 ( .A1(n16136), .A2(n16055), .ZN(n14867) );
  OAI21_X1 U18111 ( .B1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n15400), .A(
        n15399), .ZN(n18827) );
  OAI22_X1 U18112 ( .A1(n11585), .A2(n18846), .B1(n19045), .B2(n18827), .ZN(
        n14865) );
  INV_X1 U18113 ( .A(n18830), .ZN(n14863) );
  NOR2_X1 U18114 ( .A1(n14863), .A2(n16058), .ZN(n14864) );
  AOI211_X1 U18115 ( .C1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .C2(n19032), .A(
        n14865), .B(n14864), .ZN(n14866) );
  OAI211_X1 U18116 ( .C1(n16140), .C2(n19037), .A(n14867), .B(n14866), .ZN(
        P2_U3004) );
  NOR2_X1 U18117 ( .A1(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n14868), .ZN(
        n14870) );
  NAND2_X1 U18118 ( .A1(n14871), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14872) );
  OAI211_X1 U18119 ( .C1(n14874), .C2(n19061), .A(n14873), .B(n14872), .ZN(
        n14875) );
  AOI21_X1 U18120 ( .B1(n14876), .B2(n19065), .A(n14875), .ZN(n14877) );
  OAI21_X1 U18121 ( .B1(n19056), .B2(n14878), .A(n14877), .ZN(P2_U3016) );
  INV_X1 U18122 ( .A(n14883), .ZN(n14881) );
  NOR3_X1 U18123 ( .A1(n9881), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n14881), .ZN(n14879) );
  AOI211_X1 U18124 ( .C1(n15856), .C2(n19059), .A(n14880), .B(n14879), .ZN(
        n14886) );
  INV_X1 U18125 ( .A(n14905), .ZN(n14882) );
  NOR2_X1 U18126 ( .A1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n14881), .ZN(
        n14902) );
  NOR2_X1 U18127 ( .A1(n14882), .A2(n14902), .ZN(n14896) );
  INV_X1 U18128 ( .A(n14896), .ZN(n14884) );
  AND3_X1 U18129 ( .A1(n14895), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A3(
        n14883), .ZN(n14891) );
  OAI21_X1 U18130 ( .B1(n14884), .B2(n14891), .A(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14885) );
  OAI211_X1 U18131 ( .C1(n15862), .C2(n19061), .A(n14886), .B(n14885), .ZN(
        n14887) );
  AOI21_X1 U18132 ( .B1(n14888), .B2(n19065), .A(n14887), .ZN(n14889) );
  OAI21_X1 U18133 ( .B1(n19056), .B2(n14890), .A(n14889), .ZN(P2_U3017) );
  NAND2_X1 U18134 ( .A1(n15865), .A2(n16154), .ZN(n14894) );
  AOI211_X1 U18135 ( .C1(n15864), .C2(n19059), .A(n14892), .B(n14891), .ZN(
        n14893) );
  OAI211_X1 U18136 ( .C1(n14896), .C2(n14895), .A(n14894), .B(n14893), .ZN(
        n14897) );
  AOI21_X1 U18137 ( .B1(n14898), .B2(n16157), .A(n14897), .ZN(n14899) );
  OAI21_X1 U18138 ( .B1(n14900), .B2(n16139), .A(n14899), .ZN(P2_U3018) );
  INV_X1 U18139 ( .A(n15884), .ZN(n14908) );
  AOI211_X1 U18140 ( .C1(n15878), .C2(n19059), .A(n14902), .B(n14901), .ZN(
        n14903) );
  OAI21_X1 U18141 ( .B1(n14905), .B2(n14904), .A(n14903), .ZN(n14907) );
  NOR2_X1 U18142 ( .A1(n14910), .A2(n19056), .ZN(n14918) );
  NAND2_X1 U18143 ( .A1(n15889), .A2(n16154), .ZN(n14916) );
  OAI21_X1 U18144 ( .B1(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(n14911), .ZN(n14913) );
  OR2_X1 U18145 ( .A1(n20880), .A2(n18823), .ZN(n14912) );
  OAI21_X1 U18146 ( .B1(n14931), .B2(n14913), .A(n14912), .ZN(n14914) );
  AOI21_X1 U18147 ( .B1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n14927), .A(
        n14914), .ZN(n14915) );
  OAI211_X1 U18148 ( .C1(n15895), .C2(n16131), .A(n14916), .B(n14915), .ZN(
        n14917) );
  AOI211_X1 U18149 ( .C1(n14919), .C2(n19065), .A(n14918), .B(n14917), .ZN(
        n14920) );
  INV_X1 U18150 ( .A(n14920), .ZN(P2_U3020) );
  INV_X1 U18151 ( .A(n14921), .ZN(n14922) );
  NOR2_X1 U18152 ( .A1(n14923), .A2(n14922), .ZN(n14924) );
  XNOR2_X1 U18153 ( .A(n14925), .B(n14924), .ZN(n15937) );
  INV_X1 U18154 ( .A(n15937), .ZN(n14936) );
  AOI21_X1 U18155 ( .B1(n14930), .B2(n14937), .A(n14926), .ZN(n15936) );
  INV_X1 U18156 ( .A(n14927), .ZN(n14929) );
  NAND2_X1 U18157 ( .A1(P2_REIP_REG_25__SCAN_IN), .A2(n19033), .ZN(n14928) );
  OAI221_X1 U18158 ( .B1(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n14931), 
        .C1(n14930), .C2(n14929), .A(n14928), .ZN(n14934) );
  OAI22_X1 U18159 ( .A1(n15934), .A2(n19061), .B1(n16131), .B2(n14932), .ZN(
        n14933) );
  AOI211_X1 U18160 ( .C1(n15936), .C2(n16157), .A(n14934), .B(n14933), .ZN(
        n14935) );
  OAI21_X1 U18161 ( .B1(n14936), .B2(n16139), .A(n14935), .ZN(P2_U3021) );
  OAI21_X1 U18162 ( .B1(n9790), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n14937), .ZN(n15942) );
  INV_X1 U18163 ( .A(n14939), .ZN(n14941) );
  NAND2_X1 U18164 ( .A1(n14941), .A2(n14940), .ZN(n14942) );
  XNOR2_X1 U18165 ( .A(n14938), .B(n14942), .ZN(n15941) );
  NOR2_X1 U18166 ( .A1(n14943), .A2(n14946), .ZN(n14950) );
  NAND2_X1 U18167 ( .A1(n15945), .A2(n16154), .ZN(n14948) );
  NOR2_X1 U18168 ( .A1(n19659), .A2(n18846), .ZN(n14944) );
  AOI21_X1 U18169 ( .B1(n14946), .B2(n14945), .A(n14944), .ZN(n14947) );
  OAI211_X1 U18170 ( .C1(n15913), .C2(n16131), .A(n14948), .B(n14947), .ZN(
        n14949) );
  AOI211_X1 U18171 ( .C1(n15941), .C2(n19065), .A(n14950), .B(n14949), .ZN(
        n14951) );
  OAI21_X1 U18172 ( .B1(n19056), .B2(n15942), .A(n14951), .ZN(P2_U3022) );
  AOI21_X1 U18173 ( .B1(n14956), .B2(n14952), .A(n15950), .ZN(n15962) );
  INV_X1 U18174 ( .A(n15962), .ZN(n14962) );
  XNOR2_X1 U18175 ( .A(n14954), .B(n14953), .ZN(n15963) );
  NAND2_X1 U18176 ( .A1(n15963), .A2(n19065), .ZN(n14961) );
  NOR2_X1 U18177 ( .A1(n15966), .A2(n19061), .ZN(n14959) );
  INV_X1 U18178 ( .A(n14955), .ZN(n16073) );
  AOI22_X1 U18179 ( .A1(n19033), .A2(P2_REIP_REG_22__SCAN_IN), .B1(n14956), 
        .B2(n16073), .ZN(n14957) );
  OAI21_X1 U18180 ( .B1(n16131), .B2(n15392), .A(n14957), .ZN(n14958) );
  AOI211_X1 U18181 ( .C1(n16067), .C2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n14959), .B(n14958), .ZN(n14960) );
  OAI211_X1 U18182 ( .C1(n14962), .C2(n19056), .A(n14961), .B(n14960), .ZN(
        P2_U3024) );
  NAND2_X1 U18183 ( .A1(n19059), .A2(n18700), .ZN(n14963) );
  OAI211_X1 U18184 ( .C1(n18706), .C2(n19061), .A(n14964), .B(n14963), .ZN(
        n14965) );
  AOI21_X1 U18185 ( .B1(n14967), .B2(n14966), .A(n14965), .ZN(n14969) );
  NAND2_X1 U18186 ( .A1(n16067), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n14968) );
  OAI211_X1 U18187 ( .C1(n14970), .C2(n19056), .A(n14969), .B(n14968), .ZN(
        n14971) );
  INV_X1 U18188 ( .A(n14971), .ZN(n14972) );
  OAI21_X1 U18189 ( .B1(n14973), .B2(n16139), .A(n14972), .ZN(P2_U3025) );
  NAND2_X1 U18190 ( .A1(n14974), .A2(n19065), .ZN(n14982) );
  INV_X1 U18191 ( .A(n16079), .ZN(n14980) );
  XNOR2_X1 U18192 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .B(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n14978) );
  NOR2_X1 U18193 ( .A1(n16131), .A2(n18708), .ZN(n14975) );
  AOI211_X1 U18194 ( .C1(n18710), .C2(n16154), .A(n14976), .B(n14975), .ZN(
        n14977) );
  OAI21_X1 U18195 ( .B1(n16080), .B2(n14978), .A(n14977), .ZN(n14979) );
  AOI21_X1 U18196 ( .B1(n14980), .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n14979), .ZN(n14981) );
  OAI211_X1 U18197 ( .C1(n14983), .C2(n19056), .A(n14982), .B(n14981), .ZN(
        P2_U3026) );
  INV_X1 U18198 ( .A(n14984), .ZN(n16120) );
  NOR4_X1 U18199 ( .A1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n15004), .A3(
        n14985), .A4(n16120), .ZN(n14987) );
  NOR2_X1 U18200 ( .A1(n16131), .A2(n18740), .ZN(n14986) );
  AOI211_X1 U18201 ( .C1(P2_REIP_REG_18__SCAN_IN), .C2(n19033), .A(n14987), 
        .B(n14986), .ZN(n14988) );
  OAI21_X1 U18202 ( .B1(n16079), .B2(n14989), .A(n14988), .ZN(n14992) );
  NOR2_X1 U18203 ( .A1(n14990), .A2(n19056), .ZN(n14991) );
  AOI211_X1 U18204 ( .C1(n18734), .C2(n16154), .A(n14992), .B(n14991), .ZN(
        n14993) );
  OAI21_X1 U18205 ( .B1(n14994), .B2(n16139), .A(n14993), .ZN(P2_U3028) );
  OR2_X1 U18206 ( .A1(n16157), .A2(n14995), .ZN(n15002) );
  INV_X1 U18207 ( .A(n14996), .ZN(n14997) );
  NAND2_X1 U18208 ( .A1(n14998), .A2(n14997), .ZN(n14999) );
  NAND2_X1 U18209 ( .A1(n16119), .A2(n14999), .ZN(n16086) );
  NOR2_X1 U18210 ( .A1(n19048), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15000) );
  OR2_X1 U18211 ( .A1(n16086), .A2(n15000), .ZN(n15001) );
  AOI21_X1 U18212 ( .B1(n15981), .B2(n15002), .A(n15001), .ZN(n15422) );
  NAND2_X1 U18213 ( .A1(n15003), .A2(n19065), .ZN(n15010) );
  OAI22_X1 U18214 ( .A1(n15005), .A2(n19056), .B1(n16120), .B2(n15004), .ZN(
        n15424) );
  NOR2_X1 U18215 ( .A1(n15006), .A2(n19061), .ZN(n15008) );
  OAI22_X1 U18216 ( .A1(n16131), .A2(n18764), .B1(n18846), .B2(n19647), .ZN(
        n15007) );
  AOI211_X1 U18217 ( .C1(n15424), .C2(n20745), .A(n15008), .B(n15007), .ZN(
        n15009) );
  OAI211_X1 U18218 ( .C1(n15422), .C2(n20745), .A(n15010), .B(n15009), .ZN(
        P2_U3030) );
  NAND2_X1 U18219 ( .A1(n15011), .A2(n16157), .ZN(n15023) );
  OAI21_X1 U18220 ( .B1(n16163), .B2(n15012), .A(n16119), .ZN(n16110) );
  NOR2_X1 U18221 ( .A1(n15013), .A2(n16120), .ZN(n16111) );
  OAI211_X1 U18222 ( .C1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n16103), .A(
        n16111), .B(n16091), .ZN(n15019) );
  OR2_X1 U18223 ( .A1(n15014), .A2(n16097), .ZN(n15016) );
  NAND2_X1 U18224 ( .A1(n15016), .A2(n15015), .ZN(n18936) );
  INV_X1 U18225 ( .A(n18936), .ZN(n15017) );
  AOI22_X1 U18226 ( .A1(n19059), .A2(n15017), .B1(n19033), .B2(
        P2_REIP_REG_14__SCAN_IN), .ZN(n15018) );
  OAI211_X1 U18227 ( .C1(n15020), .C2(n19061), .A(n15019), .B(n15018), .ZN(
        n15021) );
  AOI21_X1 U18228 ( .B1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n16110), .A(
        n15021), .ZN(n15022) );
  OAI211_X1 U18229 ( .C1(n15024), .C2(n16139), .A(n15023), .B(n15022), .ZN(
        P2_U3032) );
  OAI21_X1 U18230 ( .B1(n14819), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n15025), .ZN(n16022) );
  NOR2_X1 U18231 ( .A1(n15027), .A2(n15026), .ZN(n15028) );
  XNOR2_X1 U18232 ( .A(n15029), .B(n15028), .ZN(n16024) );
  NAND2_X1 U18233 ( .A1(P2_REIP_REG_9__SCAN_IN), .A2(n19033), .ZN(n15030) );
  OAI221_X1 U18234 ( .B1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n16120), .C1(
        n16121), .C2(n16119), .A(n15030), .ZN(n15038) );
  OR2_X1 U18235 ( .A1(n15032), .A2(n10153), .ZN(n15035) );
  INV_X1 U18236 ( .A(n15033), .ZN(n15034) );
  AND2_X1 U18237 ( .A1(n15035), .A2(n15034), .ZN(n18943) );
  INV_X1 U18238 ( .A(n18943), .ZN(n15036) );
  OAI22_X1 U18239 ( .A1(n18844), .A2(n19061), .B1(n16131), .B2(n15036), .ZN(
        n15037) );
  AOI211_X1 U18240 ( .C1(n16024), .C2(n19065), .A(n15038), .B(n15037), .ZN(
        n15039) );
  OAI21_X1 U18241 ( .B1(n16022), .B2(n19056), .A(n15039), .ZN(P2_U3037) );
  XNOR2_X1 U18242 ( .A(n15040), .B(n15041), .ZN(n16029) );
  NAND2_X1 U18243 ( .A1(n15043), .A2(n15061), .ZN(n15044) );
  NAND2_X1 U18244 ( .A1(n15044), .A2(n15062), .ZN(n15048) );
  AND2_X1 U18245 ( .A1(n15046), .A2(n15045), .ZN(n15047) );
  XNOR2_X1 U18246 ( .A(n15048), .B(n15047), .ZN(n16028) );
  NOR2_X1 U18247 ( .A1(n11576), .A2(n18846), .ZN(n15052) );
  INV_X1 U18248 ( .A(n15049), .ZN(n15050) );
  AOI211_X1 U18249 ( .C1(n15066), .C2(n20738), .A(n15050), .B(n15067), .ZN(
        n15051) );
  AOI211_X1 U18250 ( .C1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .C2(n15053), .A(
        n15052), .B(n15051), .ZN(n15056) );
  INV_X1 U18251 ( .A(n18857), .ZN(n15054) );
  AOI22_X1 U18252 ( .A1(n18853), .A2(n16154), .B1(n19059), .B2(n15054), .ZN(
        n15055) );
  OAI211_X1 U18253 ( .C1(n16028), .C2(n16139), .A(n15056), .B(n15055), .ZN(
        n15057) );
  INV_X1 U18254 ( .A(n15057), .ZN(n15058) );
  OAI21_X1 U18255 ( .B1(n16029), .B2(n19056), .A(n15058), .ZN(P2_U3038) );
  XNOR2_X1 U18256 ( .A(n15060), .B(n15059), .ZN(n16033) );
  NAND2_X1 U18257 ( .A1(n15062), .A2(n15061), .ZN(n15063) );
  XNOR2_X1 U18258 ( .A(n15043), .B(n15063), .ZN(n16036) );
  NAND2_X1 U18259 ( .A1(P2_REIP_REG_7__SCAN_IN), .A2(n19033), .ZN(n15064) );
  OAI221_X1 U18260 ( .B1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n15067), .C1(
        n15066), .C2(n15065), .A(n15064), .ZN(n15070) );
  OAI22_X1 U18261 ( .A1(n18870), .A2(n19061), .B1(n16131), .B2(n15068), .ZN(
        n15069) );
  AOI211_X1 U18262 ( .C1(n16036), .C2(n19065), .A(n15070), .B(n15069), .ZN(
        n15071) );
  OAI21_X1 U18263 ( .B1(n16033), .B2(n19056), .A(n15071), .ZN(P2_U3039) );
  INV_X1 U18264 ( .A(n15072), .ZN(n15102) );
  NAND2_X1 U18265 ( .A1(n15074), .A2(n15073), .ZN(n15080) );
  MUX2_X1 U18266 ( .A(n15080), .B(n15091), .S(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Z(n15075) );
  AOI21_X1 U18267 ( .B1(n18926), .B2(n15102), .A(n15075), .ZN(n16181) );
  OAI222_X1 U18268 ( .A1(n15104), .A2(n15077), .B1(n19687), .B2(n16181), .C1(
        n13196), .C2(n15076), .ZN(n15078) );
  MUX2_X1 U18269 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B(n15078), .S(
        n15106), .Z(P2_U3601) );
  INV_X1 U18270 ( .A(n15079), .ZN(n15086) );
  NAND2_X1 U18271 ( .A1(n15091), .A2(n10280), .ZN(n15082) );
  OAI21_X1 U18272 ( .B1(n10510), .B2(n10509), .A(n15080), .ZN(n15081) );
  NAND2_X1 U18273 ( .A1(n15082), .A2(n15081), .ZN(n15083) );
  AOI21_X1 U18274 ( .B1(n15084), .B2(n15102), .A(n15083), .ZN(n16186) );
  OAI222_X1 U18275 ( .A1(n15104), .A2(n19707), .B1(n15086), .B2(n15085), .C1(
        n19687), .C2(n16186), .ZN(n15087) );
  MUX2_X1 U18276 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n15087), .S(
        n15106), .Z(P2_U3600) );
  INV_X1 U18277 ( .A(n15094), .ZN(n15088) );
  AOI22_X1 U18278 ( .A1(n15089), .A2(n15088), .B1(n11447), .B2(n15091), .ZN(
        n15099) );
  NAND2_X1 U18279 ( .A1(n15091), .A2(n15090), .ZN(n15097) );
  NAND2_X1 U18280 ( .A1(n15093), .A2(n15092), .ZN(n15095) );
  AOI21_X1 U18281 ( .B1(n15095), .B2(n10286), .A(n15094), .ZN(n15096) );
  AND2_X1 U18282 ( .A1(n15097), .A2(n15096), .ZN(n15098) );
  MUX2_X1 U18283 ( .A(n15099), .B(n15098), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n15100) );
  NAND2_X1 U18284 ( .A1(n15100), .A2(n10267), .ZN(n15101) );
  AOI21_X1 U18285 ( .B1(n15103), .B2(n15102), .A(n15101), .ZN(n16166) );
  OAI22_X1 U18286 ( .A1(n15105), .A2(n15104), .B1(n16166), .B2(n19687), .ZN(
        n15107) );
  MUX2_X1 U18287 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n15107), .S(
        n15106), .Z(P2_U3596) );
  AOI22_X1 U18288 ( .A1(n15162), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n16777), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n15111) );
  AOI22_X1 U18289 ( .A1(n16968), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n15279), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n15110) );
  AOI22_X1 U18290 ( .A1(n16993), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n16974), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n15109) );
  AOI22_X1 U18291 ( .A1(n15294), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n16969), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n15108) );
  NAND4_X1 U18292 ( .A1(n15111), .A2(n15110), .A3(n15109), .A4(n15108), .ZN(
        n15117) );
  AOI22_X1 U18293 ( .A1(n9726), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n16987), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n15115) );
  AOI22_X1 U18294 ( .A1(n9729), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n15254), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n15114) );
  AOI22_X1 U18295 ( .A1(n16988), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n15318), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n15113) );
  AOI22_X1 U18296 ( .A1(n11754), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n15286), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n15112) );
  NAND4_X1 U18297 ( .A1(n15115), .A2(n15114), .A3(n15113), .A4(n15112), .ZN(
        n15116) );
  NOR2_X1 U18298 ( .A1(n15117), .A2(n15116), .ZN(n16792) );
  AOI22_X1 U18299 ( .A1(n16992), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n15279), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n15122) );
  AOI22_X1 U18300 ( .A1(n15162), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n15318), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n15121) );
  AOI22_X1 U18301 ( .A1(n15118), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n15286), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n15120) );
  AOI22_X1 U18302 ( .A1(n16954), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n16969), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n15119) );
  NAND4_X1 U18303 ( .A1(n15122), .A2(n15121), .A3(n15120), .A4(n15119), .ZN(
        n15128) );
  AOI22_X1 U18304 ( .A1(n16993), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n16974), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n15126) );
  AOI22_X1 U18305 ( .A1(n9729), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11754), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n15125) );
  AOI22_X1 U18306 ( .A1(n16968), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n15254), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n15124) );
  AOI22_X1 U18307 ( .A1(n15294), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n16988), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n15123) );
  NAND4_X1 U18308 ( .A1(n15126), .A2(n15125), .A3(n15124), .A4(n15123), .ZN(
        n15127) );
  NOR2_X1 U18309 ( .A1(n15128), .A2(n15127), .ZN(n16802) );
  AOI22_X1 U18310 ( .A1(n16993), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_7__1__SCAN_IN), .B2(n16974), .ZN(n15132) );
  AOI22_X1 U18311 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n16959), .B1(
        P3_INSTQUEUE_REG_12__1__SCAN_IN), .B2(n16991), .ZN(n15131) );
  AOI22_X1 U18312 ( .A1(n15162), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n15318), .ZN(n15130) );
  AOI22_X1 U18313 ( .A1(n16968), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n16969), .ZN(n15129) );
  NAND4_X1 U18314 ( .A1(n15132), .A2(n15131), .A3(n15130), .A4(n15129), .ZN(
        n15138) );
  AOI22_X1 U18315 ( .A1(n15118), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_4__1__SCAN_IN), .B2(n11754), .ZN(n15136) );
  AOI22_X1 U18316 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n16954), .B1(
        P3_INSTQUEUE_REG_0__1__SCAN_IN), .B2(n15279), .ZN(n15135) );
  AOI22_X1 U18317 ( .A1(n15294), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n16777), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n15134) );
  AOI22_X1 U18318 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n9729), .B1(
        n16988), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n15133) );
  NAND4_X1 U18319 ( .A1(n15136), .A2(n15135), .A3(n15134), .A4(n15133), .ZN(
        n15137) );
  NOR2_X1 U18320 ( .A1(n15138), .A2(n15137), .ZN(n16813) );
  AOI22_X1 U18321 ( .A1(n16993), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n16987), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n15148) );
  AOI22_X1 U18322 ( .A1(n15162), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n16777), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n15147) );
  INV_X1 U18323 ( .A(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n20930) );
  AOI22_X1 U18324 ( .A1(n15118), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n9729), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n15139) );
  OAI21_X1 U18325 ( .B1(n16767), .B2(n20930), .A(n15139), .ZN(n15145) );
  AOI22_X1 U18326 ( .A1(n16968), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n15286), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n15143) );
  AOI22_X1 U18327 ( .A1(n11754), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n16974), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n15142) );
  AOI22_X1 U18328 ( .A1(n15318), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n15254), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n15141) );
  AOI22_X1 U18329 ( .A1(n16988), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n16969), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n15140) );
  NAND4_X1 U18330 ( .A1(n15143), .A2(n15142), .A3(n15141), .A4(n15140), .ZN(
        n15144) );
  AOI211_X1 U18331 ( .C1(n17000), .C2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A(
        n15145), .B(n15144), .ZN(n15146) );
  NAND3_X1 U18332 ( .A1(n15148), .A2(n15147), .A3(n15146), .ZN(n16818) );
  AOI22_X1 U18333 ( .A1(n15149), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n15254), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n15160) );
  AOI22_X1 U18334 ( .A1(n15162), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n16988), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n15159) );
  INV_X1 U18335 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n17009) );
  AOI22_X1 U18336 ( .A1(n11754), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n16974), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n15150) );
  OAI21_X1 U18337 ( .B1(n9785), .B2(n17009), .A(n15150), .ZN(n15157) );
  AOI22_X1 U18338 ( .A1(n16968), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n15279), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n15155) );
  AOI22_X1 U18339 ( .A1(n16959), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n16777), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n15154) );
  AOI22_X1 U18340 ( .A1(n9729), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n16987), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n15153) );
  AOI22_X1 U18341 ( .A1(n16993), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n16969), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n15152) );
  NAND4_X1 U18342 ( .A1(n15155), .A2(n15154), .A3(n15153), .A4(n15152), .ZN(
        n15156) );
  AOI211_X1 U18343 ( .C1(n9726), .C2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A(
        n15157), .B(n15156), .ZN(n15158) );
  NAND3_X1 U18344 ( .A1(n15160), .A2(n15159), .A3(n15158), .ZN(n16819) );
  NAND2_X1 U18345 ( .A1(n16818), .A2(n16819), .ZN(n16817) );
  NOR2_X1 U18346 ( .A1(n16813), .A2(n16817), .ZN(n16809) );
  AOI22_X1 U18347 ( .A1(n9729), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n16987), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n15171) );
  AOI22_X1 U18348 ( .A1(n16992), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n15279), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n15170) );
  AOI22_X1 U18349 ( .A1(n15118), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n15318), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n15161) );
  OAI21_X1 U18350 ( .B1(n10274), .B2(n20798), .A(n15161), .ZN(n15168) );
  AOI22_X1 U18351 ( .A1(n15162), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n15254), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n15166) );
  AOI22_X1 U18352 ( .A1(n11754), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n15286), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n15165) );
  AOI22_X1 U18353 ( .A1(n16993), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n16975), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n15164) );
  AOI22_X1 U18354 ( .A1(n16968), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n16969), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n15163) );
  NAND4_X1 U18355 ( .A1(n15166), .A2(n15165), .A3(n15164), .A4(n15163), .ZN(
        n15167) );
  AOI211_X1 U18356 ( .C1(n17000), .C2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A(
        n15168), .B(n15167), .ZN(n15169) );
  NAND3_X1 U18357 ( .A1(n15171), .A2(n15170), .A3(n15169), .ZN(n16808) );
  NAND2_X1 U18358 ( .A1(n16809), .A2(n16808), .ZN(n16807) );
  NOR2_X1 U18359 ( .A1(n16802), .A2(n16807), .ZN(n17067) );
  AOI22_X1 U18360 ( .A1(n9726), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n15286), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n15181) );
  AOI22_X1 U18361 ( .A1(n16975), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n15279), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n15180) );
  INV_X1 U18362 ( .A(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n20832) );
  AOI22_X1 U18363 ( .A1(n16954), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n16974), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n15172) );
  OAI21_X1 U18364 ( .B1(n9787), .B2(n20832), .A(n15172), .ZN(n15178) );
  AOI22_X1 U18365 ( .A1(n15162), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n9729), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n15176) );
  AOI22_X1 U18366 ( .A1(n15294), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n16777), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n15175) );
  AOI22_X1 U18367 ( .A1(n15318), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n15254), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n15174) );
  AOI22_X1 U18368 ( .A1(n11754), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n16969), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n15173) );
  NAND4_X1 U18369 ( .A1(n15176), .A2(n15175), .A3(n15174), .A4(n15173), .ZN(
        n15177) );
  AOI211_X1 U18370 ( .C1(n16993), .C2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A(
        n15178), .B(n15177), .ZN(n15179) );
  NAND3_X1 U18371 ( .A1(n15181), .A2(n15180), .A3(n15179), .ZN(n17066) );
  NAND2_X1 U18372 ( .A1(n17067), .A2(n17066), .ZN(n17065) );
  XNOR2_X1 U18373 ( .A(n16792), .B(n17065), .ZN(n17064) );
  INV_X1 U18374 ( .A(P3_EBX_REG_26__SCAN_IN), .ZN(n16805) );
  INV_X1 U18375 ( .A(P3_EBX_REG_24__SCAN_IN), .ZN(n16758) );
  INV_X1 U18376 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n16497) );
  NAND2_X1 U18377 ( .A1(n17047), .A2(n16835), .ZN(n16848) );
  INV_X1 U18378 ( .A(P3_EBX_REG_28__SCAN_IN), .ZN(n16440) );
  INV_X1 U18379 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n16800) );
  NOR2_X1 U18380 ( .A1(n16440), .A2(n16800), .ZN(n16796) );
  NAND2_X1 U18381 ( .A1(n17047), .A2(n17034), .ZN(n17037) );
  NAND2_X1 U18382 ( .A1(n17039), .A2(n16801), .ZN(n16804) );
  OAI21_X1 U18383 ( .B1(n16796), .B2(n17037), .A(n16804), .ZN(n16797) );
  OAI221_X1 U18384 ( .B1(P3_EBX_REG_28__SCAN_IN), .B2(n15183), .C1(
        P3_EBX_REG_28__SCAN_IN), .C2(P3_EBX_REG_27__SCAN_IN), .A(n16797), .ZN(
        n15184) );
  OAI21_X1 U18385 ( .B1(n17039), .B2(n17064), .A(n15184), .ZN(P3_U2675) );
  AOI22_X1 U18386 ( .A1(n15151), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n15318), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n15188) );
  AOI22_X1 U18387 ( .A1(n16988), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n16777), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n15187) );
  AOI22_X1 U18388 ( .A1(n15149), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n16974), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n15186) );
  AOI22_X1 U18389 ( .A1(n11754), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n16969), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n15185) );
  NAND4_X1 U18390 ( .A1(n15188), .A2(n15187), .A3(n15186), .A4(n15185), .ZN(
        n15194) );
  AOI22_X1 U18391 ( .A1(n16968), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n15286), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n15192) );
  AOI22_X1 U18392 ( .A1(n16954), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n15254), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n15191) );
  AOI22_X1 U18393 ( .A1(n15162), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n16993), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n15190) );
  AOI22_X1 U18394 ( .A1(n9726), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n15279), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n15189) );
  NAND4_X1 U18395 ( .A1(n15192), .A2(n15191), .A3(n15190), .A4(n15189), .ZN(
        n15193) );
  NOR2_X1 U18396 ( .A1(n15194), .A2(n15193), .ZN(n17137) );
  OAI221_X1 U18397 ( .B1(n16901), .B2(P3_EBX_REG_13__SCAN_IN), .C1(n15196), 
        .C2(n15195), .A(n17039), .ZN(n15197) );
  OAI21_X1 U18398 ( .B1(n17137), .B2(n17039), .A(n15197), .ZN(P3_U2690) );
  NAND2_X1 U18399 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n18240) );
  AOI221_X1 U18400 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n18240), .C1(n15199), 
        .C2(n18240), .A(n15198), .ZN(n18007) );
  NOR2_X1 U18401 ( .A1(n15200), .A2(n18288), .ZN(n15201) );
  OAI21_X1 U18402 ( .B1(n15201), .B2(n18083), .A(n18008), .ZN(n18005) );
  AOI22_X1 U18403 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18007), .B1(
        n18005), .B2(n18013), .ZN(P3_U2865) );
  INV_X1 U18404 ( .A(n18648), .ZN(n18495) );
  NOR4_X1 U18405 ( .A1(n18650), .A2(n15233), .A3(n17200), .A4(n18652), .ZN(
        n15211) );
  INV_X1 U18406 ( .A(n15203), .ZN(n15205) );
  NOR2_X1 U18407 ( .A1(n15205), .A2(n15204), .ZN(n15206) );
  OAI211_X1 U18408 ( .C1(n15229), .C2(n17048), .A(n15219), .B(n15206), .ZN(
        n15241) );
  OAI21_X1 U18409 ( .B1(n15241), .B2(n15208), .A(n15207), .ZN(n15210) );
  NAND2_X1 U18410 ( .A1(n15210), .A2(n15209), .ZN(n15235) );
  NOR4_X2 U18411 ( .A1(n15511), .A2(n15212), .A3(n15211), .A4(n15235), .ZN(
        n18483) );
  NAND2_X1 U18412 ( .A1(n18596), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n18010) );
  OR2_X1 U18413 ( .A1(n16382), .A2(n18598), .ZN(n15213) );
  OAI211_X1 U18414 ( .C1(n18495), .C2(n18483), .A(n18010), .B(n15213), .ZN(
        n18628) );
  INV_X1 U18415 ( .A(n15214), .ZN(n18475) );
  AND2_X1 U18416 ( .A1(n15215), .A2(n18475), .ZN(n18451) );
  NAND3_X1 U18417 ( .A1(n18628), .A2(n18667), .A3(n18451), .ZN(n15216) );
  OAI21_X1 U18418 ( .B1(n18628), .B2(n16695), .A(n15216), .ZN(P3_U3284) );
  NAND2_X2 U18419 ( .A1(n18458), .A2(n15218), .ZN(n18469) );
  NAND3_X1 U18420 ( .A1(n13563), .A2(n18023), .A3(n17200), .ZN(n15221) );
  NAND2_X1 U18421 ( .A1(n15222), .A2(n15221), .ZN(n18452) );
  NAND2_X2 U18422 ( .A1(n17887), .A2(n18465), .ZN(n17903) );
  NAND2_X1 U18423 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n17679) );
  NAND2_X1 U18424 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17682) );
  NOR2_X1 U18425 ( .A1(n17679), .A2(n17682), .ZN(n17320) );
  NAND3_X1 U18426 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A3(n17320), .ZN(n16280) );
  INV_X1 U18427 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n17405) );
  INV_X1 U18428 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n17773) );
  INV_X1 U18429 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n17739) );
  NOR2_X1 U18430 ( .A1(n17773), .A2(n17739), .ZN(n17753) );
  INV_X1 U18431 ( .A(n17753), .ZN(n17413) );
  NOR2_X1 U18432 ( .A1(n17405), .A2(n17413), .ZN(n15224) );
  NAND2_X1 U18433 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n17778) );
  INV_X1 U18434 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n17452) );
  NOR2_X1 U18435 ( .A1(n17778), .A2(n17452), .ZN(n15223) );
  INV_X1 U18436 ( .A(n15223), .ZN(n17736) );
  INV_X1 U18437 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n17831) );
  NAND2_X1 U18438 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n17875) );
  INV_X1 U18439 ( .A(n17875), .ZN(n17844) );
  NAND2_X1 U18440 ( .A1(n17844), .A2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n17858) );
  INV_X1 U18441 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n17864) );
  NOR2_X1 U18442 ( .A1(n17858), .A2(n17864), .ZN(n17854) );
  NAND2_X1 U18443 ( .A1(n17854), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n17829) );
  NOR2_X1 U18444 ( .A1(n17831), .A2(n17829), .ZN(n17800) );
  NAND2_X1 U18445 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n17800), .ZN(
        n16238) );
  INV_X1 U18446 ( .A(n16238), .ZN(n15225) );
  INV_X1 U18447 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n20755) );
  NAND2_X1 U18448 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n17783) );
  INV_X1 U18449 ( .A(n17783), .ZN(n17945) );
  INV_X1 U18450 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n17936) );
  INV_X1 U18451 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n17955) );
  INV_X1 U18452 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n17948) );
  NOR3_X1 U18453 ( .A1(n17936), .A2(n17955), .A3(n17948), .ZN(n17784) );
  AND2_X1 U18454 ( .A1(n17945), .A2(n17784), .ZN(n17901) );
  INV_X1 U18455 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n17902) );
  INV_X1 U18456 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n17930) );
  INV_X1 U18457 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n17907) );
  NOR3_X1 U18458 ( .A1(n17902), .A2(n17930), .A3(n17907), .ZN(n17840) );
  NAND2_X1 U18459 ( .A1(n17901), .A2(n17840), .ZN(n17885) );
  NOR2_X1 U18460 ( .A1(n20755), .A2(n17885), .ZN(n17869) );
  NAND2_X1 U18461 ( .A1(n15225), .A2(n17869), .ZN(n17798) );
  NOR2_X1 U18462 ( .A1(n17736), .A2(n17798), .ZN(n17750) );
  AOI21_X1 U18463 ( .B1(n15224), .B2(n17750), .A(n18465), .ZN(n17732) );
  NAND2_X1 U18464 ( .A1(n15223), .A2(n15224), .ZN(n17740) );
  INV_X1 U18465 ( .A(n17740), .ZN(n17737) );
  NAND2_X1 U18466 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n17737), .ZN(
        n16239) );
  NOR2_X1 U18467 ( .A1(n16238), .A2(n17885), .ZN(n17776) );
  INV_X1 U18468 ( .A(n17776), .ZN(n15383) );
  OAI21_X1 U18469 ( .B1(n16239), .B2(n15383), .A(n18469), .ZN(n17680) );
  INV_X1 U18470 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n20826) );
  NAND2_X1 U18471 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n15224), .ZN(
        n17397) );
  NOR2_X1 U18472 ( .A1(n20826), .A2(n17397), .ZN(n15379) );
  INV_X1 U18473 ( .A(n17840), .ZN(n17785) );
  INV_X1 U18474 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18612) );
  INV_X1 U18475 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n20894) );
  OAI21_X1 U18476 ( .B1(n20755), .B2(n18612), .A(n20894), .ZN(n17973) );
  NAND2_X1 U18477 ( .A1(n17784), .A2(n17973), .ZN(n17899) );
  NOR2_X1 U18478 ( .A1(n17785), .A2(n17899), .ZN(n17797) );
  NAND2_X1 U18479 ( .A1(n15225), .A2(n17797), .ZN(n17735) );
  NOR2_X1 U18480 ( .A1(n17778), .A2(n17735), .ZN(n17780) );
  NAND2_X1 U18481 ( .A1(n15379), .A2(n17780), .ZN(n17683) );
  NAND2_X1 U18482 ( .A1(n18449), .A2(n17683), .ZN(n17720) );
  NAND2_X1 U18483 ( .A1(n17680), .A2(n17720), .ZN(n15226) );
  AOI211_X1 U18484 ( .C1(n17903), .C2(n16280), .A(n17732), .B(n15226), .ZN(
        n15482) );
  AOI21_X1 U18485 ( .B1(n15228), .B2(n15227), .A(n15233), .ZN(n18445) );
  INV_X1 U18486 ( .A(n18445), .ZN(n15240) );
  INV_X1 U18487 ( .A(n18448), .ZN(n16207) );
  OAI21_X1 U18488 ( .B1(n18027), .B2(n15230), .A(n15229), .ZN(n15237) );
  NOR2_X1 U18489 ( .A1(n18654), .A2(n18027), .ZN(n15238) );
  OAI21_X1 U18490 ( .B1(n15231), .B2(n18023), .A(n18652), .ZN(n15232) );
  OAI21_X1 U18491 ( .B1(n15238), .B2(n15232), .A(n18655), .ZN(n16379) );
  NOR3_X1 U18492 ( .A1(n15234), .A2(n15233), .A3(n16379), .ZN(n15236) );
  AOI211_X1 U18493 ( .C1(n16207), .C2(n15237), .A(n15236), .B(n15235), .ZN(
        n15239) );
  NAND2_X1 U18494 ( .A1(n15238), .A2(n18046), .ZN(n15242) );
  AOI221_X4 U18495 ( .B1(n15240), .B2(n15239), .C1(n15242), .C2(n15239), .A(
        n18495), .ZN(n17989) );
  NAND2_X1 U18496 ( .A1(n15482), .A2(n17980), .ZN(n16277) );
  NAND2_X1 U18497 ( .A1(n17989), .A2(n17903), .ZN(n17987) );
  AOI22_X1 U18498 ( .A1(n16954), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n16777), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n15252) );
  AOI22_X1 U18499 ( .A1(n16975), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n15279), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n15251) );
  AOI22_X1 U18500 ( .A1(n16993), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n15318), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n15243) );
  OAI21_X1 U18501 ( .B1(n9787), .B2(n17009), .A(n15243), .ZN(n15249) );
  AOI22_X1 U18502 ( .A1(n15162), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n9726), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n15247) );
  AOI22_X1 U18503 ( .A1(n9729), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n15286), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n15246) );
  AOI22_X1 U18504 ( .A1(n11754), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n16974), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n15245) );
  AOI22_X1 U18505 ( .A1(n16969), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n15254), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n15244) );
  NAND4_X1 U18506 ( .A1(n15247), .A2(n15246), .A3(n15245), .A4(n15244), .ZN(
        n15248) );
  AOI211_X1 U18507 ( .C1(n17000), .C2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A(
        n15249), .B(n15248), .ZN(n15250) );
  INV_X1 U18508 ( .A(n16273), .ZN(n17166) );
  NAND2_X1 U18509 ( .A1(n17919), .A2(n17166), .ZN(n17873) );
  NOR2_X1 U18510 ( .A1(n17928), .A2(n17873), .ZN(n17911) );
  INV_X1 U18511 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n20733) );
  INV_X1 U18512 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n17306) );
  NOR2_X1 U18513 ( .A1(n20733), .A2(n17306), .ZN(n15385) );
  AND2_X1 U18514 ( .A1(n15385), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15483) );
  INV_X1 U18515 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17367) );
  INV_X1 U18516 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n17719) );
  NOR2_X1 U18517 ( .A1(n17719), .A2(n16239), .ZN(n17366) );
  INV_X1 U18518 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n17822) );
  AOI22_X1 U18519 ( .A1(n16993), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n16777), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n15263) );
  AOI22_X1 U18520 ( .A1(n15149), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n16975), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n15262) );
  AOI22_X1 U18521 ( .A1(n16968), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n15286), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n15253) );
  OAI21_X1 U18522 ( .B1(n9785), .B2(n20836), .A(n15253), .ZN(n15260) );
  AOI22_X1 U18523 ( .A1(n16954), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n15254), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n15258) );
  AOI22_X1 U18524 ( .A1(n11754), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n16974), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n15257) );
  AOI22_X1 U18525 ( .A1(n9729), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n15279), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n15256) );
  AOI22_X1 U18526 ( .A1(n15162), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n16969), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n15255) );
  NAND4_X1 U18527 ( .A1(n15258), .A2(n15257), .A3(n15256), .A4(n15255), .ZN(
        n15259) );
  AOI211_X1 U18528 ( .C1(n9726), .C2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A(
        n15260), .B(n15259), .ZN(n15261) );
  NAND3_X1 U18529 ( .A1(n15263), .A2(n15262), .A3(n15261), .ZN(n15343) );
  AOI22_X1 U18530 ( .A1(n15279), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n16991), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n15268) );
  AOI22_X1 U18531 ( .A1(n16993), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n16777), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n15267) );
  AOI22_X1 U18532 ( .A1(n11754), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n16969), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n15266) );
  AOI22_X1 U18533 ( .A1(n9726), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n16974), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n15265) );
  NAND4_X1 U18534 ( .A1(n15268), .A2(n15267), .A3(n15266), .A4(n15265), .ZN(
        n15274) );
  AOI22_X1 U18535 ( .A1(n15162), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n15286), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n15272) );
  AOI22_X1 U18536 ( .A1(n17000), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n16968), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n15271) );
  AOI22_X1 U18537 ( .A1(n16954), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n15318), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n15270) );
  AOI22_X1 U18538 ( .A1(n16975), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n9729), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n15269) );
  NAND4_X1 U18539 ( .A1(n15272), .A2(n15271), .A3(n15270), .A4(n15269), .ZN(
        n15273) );
  AOI22_X1 U18540 ( .A1(n11806), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n16991), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n15278) );
  AOI22_X1 U18541 ( .A1(n16993), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n15286), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n15277) );
  AOI22_X1 U18542 ( .A1(n17000), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n16975), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n15276) );
  AOI22_X1 U18543 ( .A1(n16968), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n16969), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n15275) );
  NAND4_X1 U18544 ( .A1(n15278), .A2(n15277), .A3(n15276), .A4(n15275), .ZN(
        n15285) );
  AOI22_X1 U18545 ( .A1(n9726), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n16974), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n15283) );
  AOI22_X1 U18546 ( .A1(n15162), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n15279), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n15282) );
  AOI22_X1 U18547 ( .A1(n16987), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n16777), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n15281) );
  AOI22_X1 U18548 ( .A1(n9729), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n11754), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n15280) );
  NAND4_X1 U18549 ( .A1(n15283), .A2(n15282), .A3(n15281), .A4(n15280), .ZN(
        n15284) );
  AOI22_X1 U18550 ( .A1(n16992), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n15318), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n15297) );
  AOI22_X1 U18551 ( .A1(n15162), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n15286), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n15296) );
  INV_X1 U18552 ( .A(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n20778) );
  AOI22_X1 U18553 ( .A1(n9729), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n16968), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n15287) );
  OAI21_X1 U18554 ( .B1(n9793), .B2(n20778), .A(n15287), .ZN(n15293) );
  AOI22_X1 U18555 ( .A1(n15279), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n16991), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n15291) );
  AOI22_X1 U18556 ( .A1(n9726), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11754), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n15290) );
  AOI22_X1 U18557 ( .A1(n16993), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n16987), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n15289) );
  AOI22_X1 U18558 ( .A1(n16969), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n16974), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n15288) );
  NAND4_X1 U18559 ( .A1(n15291), .A2(n15290), .A3(n15289), .A4(n15288), .ZN(
        n15292) );
  AOI211_X1 U18560 ( .C1(n15294), .C2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A(
        n15293), .B(n15292), .ZN(n15295) );
  AOI22_X1 U18561 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n16777), .B1(
        P3_INSTQUEUE_REG_14__1__SCAN_IN), .B2(n11806), .ZN(n15305) );
  AOI22_X1 U18562 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n9729), .B1(
        P3_INSTQUEUE_REG_5__1__SCAN_IN), .B2(n16988), .ZN(n15304) );
  AOI22_X1 U18563 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n16974), .B1(
        n16987), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n15298) );
  OAI21_X1 U18564 ( .B1(n20912), .B2(n16990), .A(n15298), .ZN(n15303) );
  AOI22_X1 U18565 ( .A1(n15294), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n16993), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n15302) );
  AOI22_X1 U18566 ( .A1(n15162), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n15279), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n15301) );
  AOI22_X1 U18567 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n16968), .B1(
        n16986), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n15300) );
  AOI22_X1 U18568 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n11754), .B1(
        P3_INSTQUEUE_REG_9__1__SCAN_IN), .B2(n16991), .ZN(n15299) );
  AOI22_X1 U18569 ( .A1(n16959), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n16991), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n15315) );
  AOI22_X1 U18570 ( .A1(n16777), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n15318), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n15314) );
  AOI22_X1 U18571 ( .A1(n16975), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n16968), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n15306) );
  OAI21_X1 U18572 ( .B1(n16837), .B2(n20832), .A(n15306), .ZN(n15312) );
  AOI22_X1 U18573 ( .A1(n15279), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n16974), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n15310) );
  AOI22_X1 U18574 ( .A1(n17000), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n16993), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n15309) );
  AOI22_X1 U18575 ( .A1(n9726), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n11754), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n15308) );
  AOI22_X1 U18576 ( .A1(n9729), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n16969), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n15307) );
  NAND4_X1 U18577 ( .A1(n15310), .A2(n15309), .A3(n15308), .A4(n15307), .ZN(
        n15311) );
  AOI211_X1 U18578 ( .C1(n15162), .C2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A(
        n15312), .B(n15311), .ZN(n15313) );
  NAND3_X1 U18579 ( .A1(n15315), .A2(n15314), .A3(n15313), .ZN(n15342) );
  NAND2_X1 U18580 ( .A1(n15316), .A2(n15342), .ZN(n15334) );
  XNOR2_X1 U18581 ( .A(n17171), .B(n15337), .ZN(n15335) );
  INV_X1 U18582 ( .A(n15342), .ZN(n17176) );
  NOR2_X1 U18583 ( .A1(n20894), .A2(n15328), .ZN(n15329) );
  NOR2_X1 U18584 ( .A1(n15356), .A2(n18612), .ZN(n15327) );
  AOI22_X1 U18585 ( .A1(n15279), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n16974), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n15326) );
  AOI22_X1 U18586 ( .A1(n16975), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n9729), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n15325) );
  AOI22_X1 U18587 ( .A1(n9726), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n16987), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n15317) );
  OAI21_X1 U18588 ( .B1(n9787), .B2(n20930), .A(n15317), .ZN(n15324) );
  AOI22_X1 U18589 ( .A1(n15162), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n16986), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n15322) );
  AOI22_X1 U18590 ( .A1(n17000), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n15318), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n15321) );
  AOI22_X1 U18591 ( .A1(n16777), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n16991), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n15320) );
  AOI22_X1 U18592 ( .A1(n11754), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n16969), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n15319) );
  NAND4_X1 U18593 ( .A1(n15322), .A2(n15321), .A3(n15320), .A4(n15319), .ZN(
        n15323) );
  NAND2_X1 U18594 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n17673), .ZN(
        n17672) );
  NOR2_X1 U18595 ( .A1(n17665), .A2(n17672), .ZN(n17663) );
  NOR2_X1 U18596 ( .A1(n15327), .A2(n17663), .ZN(n17654) );
  XOR2_X1 U18597 ( .A(n17181), .B(n15330), .Z(n15331) );
  XNOR2_X1 U18598 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B(n15331), .ZN(
        n17643) );
  AND2_X1 U18599 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n15331), .ZN(
        n15332) );
  XNOR2_X1 U18600 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B(n15333), .ZN(
        n17628) );
  INV_X1 U18601 ( .A(n15346), .ZN(n17172) );
  XOR2_X1 U18602 ( .A(n17172), .B(n15334), .Z(n17618) );
  XNOR2_X1 U18603 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B(n15335), .ZN(
        n17604) );
  NAND2_X1 U18604 ( .A1(n15337), .A2(n15343), .ZN(n16281) );
  OAI21_X1 U18605 ( .B1(n15338), .B2(n16273), .A(n17551), .ZN(n15340) );
  NAND2_X1 U18606 ( .A1(n17874), .A2(n17800), .ZN(n17501) );
  NAND2_X1 U18607 ( .A1(n17366), .A2(n17808), .ZN(n17715) );
  NAND2_X1 U18608 ( .A1(n15483), .A2(n17686), .ZN(n16230) );
  NOR2_X4 U18609 ( .A1(n18023), .A2(n17903), .ZN(n18447) );
  INV_X1 U18610 ( .A(n18447), .ZN(n17972) );
  INV_X1 U18611 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n20821) );
  NOR2_X1 U18612 ( .A1(n15350), .A2(n17181), .ZN(n15349) );
  NAND2_X1 U18613 ( .A1(n15349), .A2(n15342), .ZN(n15347) );
  NOR2_X1 U18614 ( .A1(n15346), .A2(n15347), .ZN(n15345) );
  NAND2_X1 U18615 ( .A1(n15345), .A2(n15343), .ZN(n15344) );
  NOR2_X1 U18616 ( .A1(n17166), .A2(n15344), .ZN(n15370) );
  XNOR2_X1 U18617 ( .A(n15344), .B(n16273), .ZN(n17596) );
  XNOR2_X1 U18618 ( .A(n15345), .B(n17171), .ZN(n15363) );
  XOR2_X1 U18619 ( .A(n15347), .B(n15346), .Z(n15348) );
  NAND2_X1 U18620 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n15348), .ZN(
        n15362) );
  XNOR2_X1 U18621 ( .A(n17936), .B(n15348), .ZN(n17615) );
  XNOR2_X1 U18622 ( .A(n15349), .B(n17176), .ZN(n15360) );
  XOR2_X1 U18623 ( .A(n17181), .B(n15350), .Z(n15351) );
  NAND2_X1 U18624 ( .A1(n15351), .A2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n15358) );
  XNOR2_X1 U18625 ( .A(n17955), .B(n15351), .ZN(n17641) );
  XOR2_X1 U18626 ( .A(n17187), .B(n15352), .Z(n15353) );
  OR2_X1 U18627 ( .A1(n20894), .A2(n15353), .ZN(n15357) );
  XNOR2_X1 U18628 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n15353), .ZN(
        n17657) );
  AOI21_X1 U18629 ( .B1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n15356), .A(
        n17673), .ZN(n15355) );
  NOR2_X1 U18630 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n15356), .ZN(
        n15354) );
  AOI221_X1 U18631 ( .B1(n17673), .B2(n15356), .C1(n15355), .C2(n20755), .A(
        n15354), .ZN(n17656) );
  NAND2_X1 U18632 ( .A1(n17657), .A2(n17656), .ZN(n17655) );
  NAND2_X1 U18633 ( .A1(n15357), .A2(n17655), .ZN(n17640) );
  NAND2_X1 U18634 ( .A1(n17641), .A2(n17640), .ZN(n17639) );
  NAND2_X1 U18635 ( .A1(n15360), .A2(n15359), .ZN(n15361) );
  NAND2_X1 U18636 ( .A1(n17615), .A2(n17614), .ZN(n17613) );
  NAND2_X1 U18637 ( .A1(n15363), .A2(n15364), .ZN(n15365) );
  NAND2_X1 U18638 ( .A1(n15370), .A2(n15366), .ZN(n15371) );
  INV_X1 U18639 ( .A(n15366), .ZN(n15369) );
  NAND2_X1 U18640 ( .A1(n17596), .A2(n17595), .ZN(n15368) );
  NAND2_X1 U18641 ( .A1(n15370), .A2(n15369), .ZN(n15367) );
  OAI211_X1 U18642 ( .C1(n15370), .C2(n15369), .A(n15368), .B(n15367), .ZN(
        n17576) );
  NAND2_X1 U18643 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n17576), .ZN(
        n17575) );
  INV_X1 U18644 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n17517) );
  NOR2_X2 U18645 ( .A1(n17494), .A2(n17822), .ZN(n17807) );
  NAND2_X1 U18646 ( .A1(n17690), .A2(n15483), .ZN(n16229) );
  AOI22_X1 U18647 ( .A1(n17911), .A2(n16230), .B1(n17982), .B2(n16229), .ZN(
        n15485) );
  OAI21_X1 U18648 ( .B1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n17987), .A(
        n15485), .ZN(n15372) );
  AOI21_X1 U18649 ( .B1(n17993), .B2(n16277), .A(n15372), .ZN(n15388) );
  INV_X1 U18650 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16248) );
  NAND3_X1 U18651 ( .A1(n17919), .A2(n17989), .A3(n16273), .ZN(n17815) );
  INV_X1 U18652 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n17704) );
  INV_X1 U18653 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n17802) );
  NOR2_X1 U18654 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n17557) );
  INV_X1 U18655 ( .A(n17557), .ZN(n17558) );
  NOR4_X1 U18656 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A4(n17558), .ZN(n15374) );
  INV_X1 U18657 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n17782) );
  NAND2_X1 U18658 ( .A1(n15375), .A2(n17366), .ZN(n15377) );
  NAND2_X1 U18659 ( .A1(n17447), .A2(n17773), .ZN(n15376) );
  NOR2_X1 U18660 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n15376), .ZN(
        n17404) );
  NAND2_X1 U18661 ( .A1(n17404), .A2(n17405), .ZN(n17398) );
  NAND2_X1 U18662 ( .A1(n17419), .A2(n17403), .ZN(n17448) );
  NAND2_X1 U18663 ( .A1(n15379), .A2(n17448), .ZN(n17370) );
  OR2_X1 U18664 ( .A1(n17585), .A2(n17357), .ZN(n17348) );
  OAI221_X1 U18665 ( .B1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n17551), 
        .C1(n17704), .C2(n17349), .A(n17348), .ZN(n17332) );
  NOR2_X1 U18666 ( .A1(n17349), .A2(n17551), .ZN(n15380) );
  NAND2_X1 U18667 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17585), .ZN(
        n16271) );
  NAND2_X1 U18668 ( .A1(n17306), .A2(n17551), .ZN(n16272) );
  OAI21_X1 U18669 ( .B1(n17321), .B2(n16271), .A(n15479), .ZN(n15382) );
  XNOR2_X1 U18670 ( .A(n15382), .B(n16248), .ZN(n16251) );
  NAND2_X1 U18671 ( .A1(n17690), .A2(n15385), .ZN(n16278) );
  INV_X1 U18672 ( .A(n18449), .ZN(n18481) );
  INV_X1 U18673 ( .A(n18465), .ZN(n17877) );
  AOI21_X1 U18674 ( .B1(n17877), .B2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n18469), .ZN(n17965) );
  OAI22_X1 U18675 ( .A1(n18481), .A2(n17735), .B1(n15383), .B2(n17965), .ZN(
        n15384) );
  INV_X1 U18676 ( .A(n15384), .ZN(n16279) );
  NOR2_X1 U18677 ( .A1(n16279), .A2(n16239), .ZN(n17702) );
  AND2_X1 U18678 ( .A1(n15385), .A2(n17320), .ZN(n16241) );
  NAND3_X1 U18679 ( .A1(n17989), .A2(n17702), .A3(n16241), .ZN(n16261) );
  NAND2_X1 U18680 ( .A1(n15385), .A2(n17686), .ZN(n16247) );
  INV_X1 U18681 ( .A(n16247), .ZN(n16275) );
  NAND2_X1 U18682 ( .A1(n17911), .A2(n16275), .ZN(n15386) );
  OAI211_X1 U18683 ( .C1(n17999), .C2(n16278), .A(n16261), .B(n15386), .ZN(
        n15487) );
  AOI22_X1 U18684 ( .A1(n17910), .A2(n16251), .B1(n16248), .B2(n15487), .ZN(
        n15387) );
  NAND2_X1 U18685 ( .A1(n17995), .A2(P3_REIP_REG_29__SCAN_IN), .ZN(n16258) );
  OAI211_X1 U18686 ( .C1(n15388), .C2(n16248), .A(n15387), .B(n16258), .ZN(
        P3_U2833) );
  AOI22_X1 U18687 ( .A1(P2_REIP_REG_22__SCAN_IN), .A2(n18918), .B1(
        P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n18882), .ZN(n15417) );
  INV_X1 U18688 ( .A(P2_EBX_REG_22__SCAN_IN), .ZN(n15389) );
  OAI22_X1 U18689 ( .A1(n15390), .A2(n18923), .B1(n18810), .B2(n15389), .ZN(
        n15391) );
  INV_X1 U18690 ( .A(n15391), .ZN(n15416) );
  OAI22_X1 U18691 ( .A1(n15966), .A2(n18894), .B1(n15392), .B2(n18898), .ZN(
        n15393) );
  INV_X1 U18692 ( .A(n15393), .ZN(n15415) );
  OAI21_X1 U18693 ( .B1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n15394), .A(
        n15834), .ZN(n15960) );
  INV_X2 U18694 ( .A(n18903), .ZN(n18863) );
  AOI21_X1 U18695 ( .B1(n15996), .B2(n15396), .A(n15395), .ZN(n18771) );
  AOI21_X1 U18696 ( .B1(n16006), .B2(n15398), .A(n15397), .ZN(n18792) );
  AOI21_X1 U18697 ( .B1(n16021), .B2(n15399), .A(n9823), .ZN(n18816) );
  AOI21_X1 U18698 ( .B1(n18836), .B2(n15406), .A(n15400), .ZN(n18840) );
  AOI21_X1 U18699 ( .B1(n18860), .B2(n15404), .A(n15407), .ZN(n18865) );
  AOI21_X1 U18700 ( .B1(n16052), .B2(n15402), .A(n15405), .ZN(n18888) );
  NOR2_X1 U18701 ( .A1(n16053), .A2(n15401), .ZN(n18902) );
  OAI21_X1 U18702 ( .B1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n15403), .A(
        n15402), .ZN(n19044) );
  NAND2_X1 U18703 ( .A1(n18902), .A2(n19044), .ZN(n18886) );
  NOR2_X1 U18704 ( .A1(n18888), .A2(n18886), .ZN(n18874) );
  OAI21_X1 U18705 ( .B1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n15405), .A(
        n15404), .ZN(n18875) );
  NAND2_X1 U18706 ( .A1(n18874), .A2(n18875), .ZN(n18862) );
  NOR2_X1 U18707 ( .A1(n18865), .A2(n18862), .ZN(n18850) );
  OAI21_X1 U18708 ( .B1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n15407), .A(
        n15406), .ZN(n18851) );
  NAND2_X1 U18709 ( .A1(n18850), .A2(n18851), .ZN(n18838) );
  NOR2_X1 U18710 ( .A1(n18840), .A2(n18838), .ZN(n18826) );
  NAND2_X1 U18711 ( .A1(n18826), .A2(n18827), .ZN(n18814) );
  NOR2_X1 U18712 ( .A1(n18816), .A2(n18814), .ZN(n18801) );
  NAND2_X1 U18713 ( .A1(n18801), .A2(n18802), .ZN(n18790) );
  NOR2_X1 U18714 ( .A1(n18792), .A2(n18790), .ZN(n18780) );
  NAND2_X1 U18715 ( .A1(n18780), .A2(n18781), .ZN(n18769) );
  NOR2_X1 U18716 ( .A1(n18771), .A2(n18769), .ZN(n18757) );
  NAND2_X1 U18717 ( .A1(n18757), .A2(n18758), .ZN(n18741) );
  AOI21_X1 U18718 ( .B1(n15409), .B2(n15408), .A(n9849), .ZN(n18743) );
  AOI21_X1 U18719 ( .B1(n15979), .B2(n15411), .A(n15410), .ZN(n15967) );
  INV_X1 U18720 ( .A(n15967), .ZN(n18725) );
  NAND2_X1 U18721 ( .A1(n18723), .A2(n12951), .ZN(n18712) );
  NAND2_X1 U18722 ( .A1(n18713), .A2(n18712), .ZN(n18711) );
  NAND2_X1 U18723 ( .A1(n18711), .A2(n12951), .ZN(n18702) );
  INV_X1 U18724 ( .A(n15412), .ZN(n18703) );
  OAI211_X1 U18725 ( .C1(n15960), .C2(n15413), .A(n10036), .B(n15833), .ZN(
        n15414) );
  NAND4_X1 U18726 ( .A1(n15417), .A2(n15416), .A3(n15415), .A4(n15414), .ZN(
        P2_U2833) );
  AOI22_X1 U18727 ( .A1(n18748), .A2(n16154), .B1(n19059), .B2(n18749), .ZN(
        n15427) );
  NAND2_X1 U18728 ( .A1(n15419), .A2(n15418), .ZN(n15420) );
  NAND2_X1 U18729 ( .A1(n15421), .A2(n15420), .ZN(n15980) );
  OAI21_X1 U18730 ( .B1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n16163), .A(
        n15422), .ZN(n15423) );
  AOI22_X1 U18731 ( .A1(n15980), .A2(n19065), .B1(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n15423), .ZN(n15426) );
  NAND3_X1 U18732 ( .A1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n14821), .A3(
        n15424), .ZN(n15425) );
  NAND2_X1 U18733 ( .A1(P2_REIP_REG_17__SCAN_IN), .A2(n19033), .ZN(n15984) );
  NAND4_X1 U18734 ( .A1(n15427), .A2(n15426), .A3(n15425), .A4(n15984), .ZN(
        P2_U3029) );
  NOR3_X1 U18735 ( .A1(n15429), .A2(n15428), .A3(n20435), .ZN(n15434) );
  AOI211_X1 U18736 ( .C1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .C2(n15434), .A(
        n15431), .B(n15430), .ZN(n15432) );
  INV_X1 U18737 ( .A(n15432), .ZN(n15433) );
  OAI21_X1 U18738 ( .B1(n15434), .B2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(
        n15433), .ZN(n15438) );
  INV_X1 U18739 ( .A(n15438), .ZN(n15436) );
  OAI21_X1 U18740 ( .B1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n15436), .A(
        n15435), .ZN(n15437) );
  OAI21_X1 U18741 ( .B1(n15438), .B2(n20321), .A(n15437), .ZN(n15439) );
  INV_X1 U18742 ( .A(n15439), .ZN(n15443) );
  INV_X1 U18743 ( .A(n15442), .ZN(n15440) );
  AOI21_X1 U18744 ( .B1(n15440), .B2(n15439), .A(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n15441) );
  AOI21_X1 U18745 ( .B1(n15443), .B2(n15442), .A(n15441), .ZN(n15451) );
  OAI21_X1 U18746 ( .B1(P1_FLUSH_REG_SCAN_IN), .B2(P1_MORE_REG_SCAN_IN), .A(
        n15444), .ZN(n15446) );
  AND4_X1 U18747 ( .A1(n15448), .A2(n15447), .A3(n15446), .A4(n15445), .ZN(
        n15450) );
  OAI211_X1 U18748 ( .C1(n15451), .C2(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A(
        n15450), .B(n15449), .ZN(n15458) );
  NAND4_X1 U18749 ( .A1(n15453), .A2(n12180), .A3(n15452), .A4(n20439), .ZN(
        n15456) );
  OAI21_X1 U18750 ( .B1(n15454), .B2(n20666), .A(n20578), .ZN(n15455) );
  NAND2_X1 U18751 ( .A1(n15456), .A2(n15455), .ZN(n15817) );
  AOI21_X1 U18752 ( .B1(n15459), .B2(n15458), .A(n15457), .ZN(n15460) );
  OAI211_X1 U18753 ( .C1(P1_STATE2_REG_2__SCAN_IN), .C2(n20666), .A(n15460), 
        .B(n15463), .ZN(n15461) );
  NOR2_X1 U18754 ( .A1(n15823), .A2(n15461), .ZN(n15466) );
  OR2_X1 U18755 ( .A1(n15463), .A2(n15462), .ZN(n15464) );
  NAND2_X1 U18756 ( .A1(n15822), .A2(n15464), .ZN(n15465) );
  OAI22_X1 U18757 ( .A1(n15466), .A2(n15822), .B1(n15823), .B2(n15465), .ZN(
        P1_U3161) );
  AOI22_X1 U18758 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n15711), .B1(
        n13009), .B2(P1_REIP_REG_21__SCAN_IN), .ZN(n15477) );
  INV_X1 U18759 ( .A(n15467), .ZN(n15475) );
  NAND2_X1 U18760 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n15468), .ZN(
        n15471) );
  INV_X1 U18761 ( .A(n15469), .ZN(n15470) );
  OAI21_X1 U18762 ( .B1(n15472), .B2(n15471), .A(n15470), .ZN(n15756) );
  NAND2_X1 U18763 ( .A1(n15473), .A2(n15756), .ZN(n15493) );
  OAI21_X1 U18764 ( .B1(n15474), .B2(n15751), .A(n15493), .ZN(n15720) );
  NAND2_X1 U18765 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n15720), .ZN(
        n15506) );
  NOR2_X1 U18766 ( .A1(n15497), .A2(n15506), .ZN(n15715) );
  AOI22_X1 U18767 ( .A1(n15475), .A2(n19994), .B1(n14305), .B2(n15715), .ZN(
        n15476) );
  OAI211_X1 U18768 ( .C1(n15807), .C2(n15537), .A(n15477), .B(n15476), .ZN(
        P1_U3010) );
  NOR2_X1 U18769 ( .A1(n17321), .A2(n16271), .ZN(n15478) );
  NAND2_X1 U18770 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n15478), .ZN(
        n16211) );
  INV_X1 U18771 ( .A(n16211), .ZN(n15480) );
  NOR2_X1 U18772 ( .A1(n15480), .A2(n16209), .ZN(n15481) );
  INV_X1 U18773 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n16231) );
  XNOR2_X1 U18774 ( .A(n15481), .B(n16231), .ZN(n16244) );
  NOR2_X1 U18775 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16248), .ZN(
        n16240) );
  OAI22_X1 U18776 ( .A1(n15483), .A2(n17987), .B1(n15482), .B2(n17928), .ZN(
        n15484) );
  NOR2_X1 U18777 ( .A1(n17918), .A2(n15484), .ZN(n16260) );
  AOI21_X1 U18778 ( .B1(n16260), .B2(n15485), .A(n16231), .ZN(n15486) );
  AOI21_X1 U18779 ( .B1(n16240), .B2(n15487), .A(n15486), .ZN(n15488) );
  NAND2_X1 U18780 ( .A1(n17979), .A2(P3_REIP_REG_30__SCAN_IN), .ZN(n16232) );
  OAI211_X1 U18781 ( .C1(n16244), .C2(n17815), .A(n15488), .B(n16232), .ZN(
        P3_U2832) );
  INV_X1 U18782 ( .A(P1_STATE_REG_1__SCAN_IN), .ZN(n19755) );
  INV_X1 U18783 ( .A(HOLD), .ZN(n20581) );
  INV_X1 U18784 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n20597) );
  NAND2_X1 U18785 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(
        P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n20596) );
  OAI21_X1 U18786 ( .B1(n20581), .B2(n19755), .A(n20596), .ZN(n15489) );
  OAI21_X1 U18787 ( .B1(n20581), .B2(n20597), .A(n15489), .ZN(n15491) );
  OAI211_X1 U18788 ( .C1(n20666), .C2(n19755), .A(n15491), .B(n15490), .ZN(
        P1_U3195) );
  AND2_X1 U18789 ( .A1(n15492), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(P1_U2905)
         );
  OAI221_X1 U18790 ( .B1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n15751), 
        .C1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n15493), .A(n15719), .ZN(
        n15494) );
  AOI22_X1 U18791 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n15494), .B1(
        n13009), .B2(P1_REIP_REG_20__SCAN_IN), .ZN(n15505) );
  NAND2_X1 U18792 ( .A1(n15495), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15499) );
  AOI21_X1 U18793 ( .B1(n15500), .B2(n15497), .A(n15496), .ZN(n15498) );
  OAI21_X1 U18794 ( .B1(n15500), .B2(n15499), .A(n15498), .ZN(n15651) );
  INV_X1 U18795 ( .A(n15501), .ZN(n15503) );
  AOI21_X1 U18796 ( .B1(n9874), .B2(n15503), .A(n15502), .ZN(n15638) );
  AOI22_X1 U18797 ( .A1(n15651), .A2(n19994), .B1(n19993), .B2(n15638), .ZN(
        n15504) );
  OAI211_X1 U18798 ( .C1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .C2(n15506), .A(
        n15505), .B(n15504), .ZN(P1_U3011) );
  NOR3_X1 U18799 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(P2_STATEBS16_REG_SCAN_IN), .ZN(n15507) );
  NAND2_X1 U18800 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19744), .ZN(n19610) );
  NOR2_X1 U18801 ( .A1(n19736), .A2(n19610), .ZN(n16195) );
  NOR4_X1 U18802 ( .A1(n15507), .A2(n19746), .A3(n16195), .A4(n16196), .ZN(
        P2_U3178) );
  AOI221_X1 U18803 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(n16196), .C1(n19729), .C2(
        n16196), .A(n19549), .ZN(n19723) );
  INV_X1 U18804 ( .A(n19723), .ZN(n19720) );
  NOR2_X1 U18805 ( .A1(n15508), .A2(n19720), .ZN(P2_U3047) );
  INV_X2 U18806 ( .A(n17192), .ZN(n17043) );
  NAND2_X1 U18807 ( .A1(n17047), .A2(n17043), .ZN(n17186) );
  INV_X1 U18808 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n17272) );
  NOR2_X1 U18809 ( .A1(n15512), .A2(n17192), .ZN(n17193) );
  AOI22_X1 U18810 ( .A1(n17193), .A2(BUF2_REG_0__SCAN_IN), .B1(n17188), .B2(
        n17673), .ZN(n15513) );
  OAI221_X1 U18811 ( .B1(P3_EAX_REG_0__SCAN_IN), .B2(n17186), .C1(n17272), 
        .C2(n17043), .A(n15513), .ZN(P3_U2735) );
  OAI22_X1 U18812 ( .A1(n13758), .A2(n19823), .B1(n15635), .B2(n19870), .ZN(
        n15514) );
  AOI221_X1 U18813 ( .B1(n15516), .B2(P1_REIP_REG_24__SCAN_IN), .C1(n15515), 
        .C2(n20636), .A(n15514), .ZN(n15519) );
  OAI22_X1 U18814 ( .A1(n15632), .A2(n15589), .B1(n15630), .B2(n19836), .ZN(
        n15517) );
  INV_X1 U18815 ( .A(n15517), .ZN(n15518) );
  OAI211_X1 U18816 ( .C1(n15520), .C2(n19829), .A(n15519), .B(n15518), .ZN(
        P1_U2816) );
  INV_X1 U18817 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n20633) );
  OAI21_X1 U18818 ( .B1(n19828), .B2(n15529), .A(n19826), .ZN(n15540) );
  OAI21_X1 U18819 ( .B1(P1_REIP_REG_21__SCAN_IN), .B2(n19838), .A(n15540), 
        .ZN(n15523) );
  INV_X1 U18820 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n15521) );
  INV_X1 U18821 ( .A(P1_EBX_REG_22__SCAN_IN), .ZN(n15637) );
  OAI22_X1 U18822 ( .A1(n15521), .A2(n19823), .B1(n15637), .B2(n19870), .ZN(
        n15522) );
  AOI221_X1 U18823 ( .B1(n15524), .B2(n20633), .C1(n15523), .C2(
        P1_REIP_REG_22__SCAN_IN), .A(n15522), .ZN(n15528) );
  INV_X1 U18824 ( .A(n15525), .ZN(n15647) );
  AOI21_X1 U18825 ( .B1(n15526), .B2(n9764), .A(n10107), .ZN(n15712) );
  AOI22_X1 U18826 ( .A1(n15647), .A2(n19816), .B1(n19856), .B2(n15712), .ZN(
        n15527) );
  OAI211_X1 U18827 ( .C1(n15650), .C2(n19829), .A(n15528), .B(n15527), .ZN(
        P1_U2818) );
  NOR3_X1 U18828 ( .A1(n19838), .A2(P1_REIP_REG_21__SCAN_IN), .A3(n15529), 
        .ZN(n15531) );
  OAI22_X1 U18829 ( .A1(n15540), .A2(n20631), .B1(n20795), .B2(n19870), .ZN(
        n15530) );
  AOI211_X1 U18830 ( .C1(n19861), .C2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        n15531), .B(n15530), .ZN(n15536) );
  OAI22_X1 U18831 ( .A1(n15533), .A2(n15589), .B1(n15532), .B2(n19829), .ZN(
        n15534) );
  INV_X1 U18832 ( .A(n15534), .ZN(n15535) );
  OAI211_X1 U18833 ( .C1(n19836), .C2(n15537), .A(n15536), .B(n15535), .ZN(
        P1_U2819) );
  AOI21_X1 U18834 ( .B1(n19857), .B2(n15538), .A(P1_REIP_REG_20__SCAN_IN), 
        .ZN(n15539) );
  OAI22_X1 U18835 ( .A1(n15540), .A2(n15539), .B1(n15640), .B2(n19870), .ZN(
        n15541) );
  AOI21_X1 U18836 ( .B1(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n19861), .A(
        n15541), .ZN(n15543) );
  AOI22_X1 U18837 ( .A1(n15652), .A2(n19816), .B1(n19856), .B2(n15638), .ZN(
        n15542) );
  OAI211_X1 U18838 ( .C1(n15655), .C2(n19829), .A(n15543), .B(n15542), .ZN(
        P1_U2820) );
  INV_X1 U18839 ( .A(n15544), .ZN(n15546) );
  OAI21_X1 U18840 ( .B1(n19838), .B2(n15546), .A(n15545), .ZN(n15598) );
  AOI21_X1 U18841 ( .B1(n19826), .B2(n15548), .A(n15598), .ZN(n15576) );
  INV_X1 U18842 ( .A(n15597), .ZN(n15547) );
  NAND3_X1 U18843 ( .A1(n15547), .A2(P1_REIP_REG_13__SCAN_IN), .A3(
        P1_REIP_REG_14__SCAN_IN), .ZN(n15580) );
  NOR2_X1 U18844 ( .A1(n15548), .A2(n15580), .ZN(n15549) );
  NAND2_X1 U18845 ( .A1(n15549), .A2(n20627), .ZN(n15558) );
  AOI21_X1 U18846 ( .B1(n19861), .B2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n13009), .ZN(n15551) );
  NAND3_X1 U18847 ( .A1(P1_REIP_REG_18__SCAN_IN), .A2(n15549), .A3(n20629), 
        .ZN(n15550) );
  OAI211_X1 U18848 ( .C1(n19870), .C2(n15552), .A(n15551), .B(n15550), .ZN(
        n15555) );
  OAI22_X1 U18849 ( .A1(n15553), .A2(n15589), .B1(n19836), .B2(n15725), .ZN(
        n15554) );
  AOI211_X1 U18850 ( .C1(n15556), .C2(n19860), .A(n15555), .B(n15554), .ZN(
        n15557) );
  OAI221_X1 U18851 ( .B1(n20629), .B2(n15576), .C1(n20629), .C2(n15558), .A(
        n15557), .ZN(P1_U2821) );
  AOI21_X1 U18852 ( .B1(n19861), .B2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n13009), .ZN(n15559) );
  OAI211_X1 U18853 ( .C1(n15576), .C2(n20627), .A(n15559), .B(n15558), .ZN(
        n15560) );
  AOI21_X1 U18854 ( .B1(P1_EBX_REG_18__SCAN_IN), .B2(n19850), .A(n15560), .ZN(
        n15565) );
  NOR2_X1 U18855 ( .A1(n15561), .A2(n19836), .ZN(n15562) );
  AOI21_X1 U18856 ( .B1(n15563), .B2(n19816), .A(n15562), .ZN(n15564) );
  OAI211_X1 U18857 ( .C1(n15566), .C2(n19829), .A(n15565), .B(n15564), .ZN(
        P1_U2822) );
  INV_X1 U18858 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n20622) );
  NOR2_X1 U18859 ( .A1(n20622), .A2(n15580), .ZN(n15577) );
  AOI21_X1 U18860 ( .B1(P1_REIP_REG_16__SCAN_IN), .B2(n15577), .A(
        P1_REIP_REG_17__SCAN_IN), .ZN(n15575) );
  OAI22_X1 U18861 ( .A1(n15568), .A2(n19823), .B1(n15567), .B2(n19870), .ZN(
        n15569) );
  AOI211_X1 U18862 ( .C1(n19860), .C2(n15570), .A(n13009), .B(n15569), .ZN(
        n15574) );
  OAI22_X1 U18863 ( .A1(n15571), .A2(n15589), .B1(n19836), .B2(n15732), .ZN(
        n15572) );
  INV_X1 U18864 ( .A(n15572), .ZN(n15573) );
  OAI211_X1 U18865 ( .C1(n15576), .C2(n15575), .A(n15574), .B(n15573), .ZN(
        P1_U2823) );
  INV_X1 U18866 ( .A(P1_REIP_REG_16__SCAN_IN), .ZN(n20624) );
  AOI22_X1 U18867 ( .A1(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n19861), .B1(
        n15577), .B2(n20624), .ZN(n15584) );
  AOI21_X1 U18868 ( .B1(n19850), .B2(P1_EBX_REG_16__SCAN_IN), .A(n13009), .ZN(
        n15583) );
  INV_X1 U18869 ( .A(n15578), .ZN(n15661) );
  INV_X1 U18870 ( .A(n15664), .ZN(n15579) );
  AOI222_X1 U18871 ( .A1(n15661), .A2(n19816), .B1(n15579), .B2(n19860), .C1(
        n19856), .C2(n15737), .ZN(n15582) );
  NOR2_X1 U18872 ( .A1(P1_REIP_REG_15__SCAN_IN), .A2(n15580), .ZN(n15585) );
  OAI21_X1 U18873 ( .B1(n15598), .B2(n15585), .A(P1_REIP_REG_16__SCAN_IN), 
        .ZN(n15581) );
  NAND4_X1 U18874 ( .A1(n15584), .A2(n15583), .A3(n15582), .A4(n15581), .ZN(
        P1_U2824) );
  AOI211_X1 U18875 ( .C1(n19861), .C2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .A(
        n13009), .B(n15585), .ZN(n15586) );
  OAI21_X1 U18876 ( .B1(n19870), .B2(n14119), .A(n15586), .ZN(n15587) );
  AOI21_X1 U18877 ( .B1(P1_REIP_REG_15__SCAN_IN), .B2(n15598), .A(n15587), 
        .ZN(n15588) );
  OAI21_X1 U18878 ( .B1(n15590), .B2(n15589), .A(n15588), .ZN(n15591) );
  AOI21_X1 U18879 ( .B1(n15592), .B2(n19860), .A(n15591), .ZN(n15593) );
  OAI21_X1 U18880 ( .B1(n19836), .B2(n15749), .A(n15593), .ZN(P1_U2825) );
  AOI22_X1 U18881 ( .A1(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n19861), .B1(
        P1_EBX_REG_14__SCAN_IN), .B2(n19850), .ZN(n15603) );
  INV_X1 U18882 ( .A(n15594), .ZN(n15595) );
  AOI21_X1 U18883 ( .B1(n15595), .B2(n19856), .A(n13009), .ZN(n15602) );
  INV_X1 U18884 ( .A(n15596), .ZN(n15666) );
  AOI22_X1 U18885 ( .A1(n15666), .A2(n19816), .B1(n19860), .B2(n15665), .ZN(
        n15601) );
  NOR2_X1 U18886 ( .A1(n20619), .A2(n15597), .ZN(n15599) );
  OAI21_X1 U18887 ( .B1(P1_REIP_REG_14__SCAN_IN), .B2(n15599), .A(n15598), 
        .ZN(n15600) );
  NAND4_X1 U18888 ( .A1(n15603), .A2(n15602), .A3(n15601), .A4(n15600), .ZN(
        P1_U2826) );
  NOR2_X1 U18889 ( .A1(n19838), .A2(n15614), .ZN(n15612) );
  AOI21_X1 U18890 ( .B1(P1_REIP_REG_11__SCAN_IN), .B2(n15612), .A(
        P1_REIP_REG_12__SCAN_IN), .ZN(n15611) );
  INV_X1 U18891 ( .A(n15604), .ZN(n15641) );
  OAI22_X1 U18892 ( .A1(n15605), .A2(n19823), .B1(n15643), .B2(n19870), .ZN(
        n15606) );
  AOI211_X1 U18893 ( .C1(n15641), .C2(n19856), .A(n13009), .B(n15606), .ZN(
        n15609) );
  INV_X1 U18894 ( .A(n15607), .ZN(n15670) );
  AOI22_X1 U18895 ( .A1(n15671), .A2(n19860), .B1(n19816), .B2(n15670), .ZN(
        n15608) );
  OAI211_X1 U18896 ( .C1(n15611), .C2(n15610), .A(n15609), .B(n15608), .ZN(
        P1_U2828) );
  AOI22_X1 U18897 ( .A1(P1_EBX_REG_11__SCAN_IN), .A2(n19850), .B1(n15612), 
        .B2(n20615), .ZN(n15618) );
  INV_X1 U18898 ( .A(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n15613) );
  OAI22_X1 U18899 ( .A1(n15613), .A2(n19823), .B1(n19836), .B2(n15766), .ZN(
        n15616) );
  OAI21_X1 U18900 ( .B1(n19828), .B2(n15614), .A(n19826), .ZN(n15629) );
  OAI21_X1 U18901 ( .B1(n15629), .B2(n20615), .A(n19845), .ZN(n15615) );
  AOI211_X1 U18902 ( .C1(n19816), .C2(n15681), .A(n15616), .B(n15615), .ZN(
        n15617) );
  OAI211_X1 U18903 ( .C1(n15684), .C2(n19829), .A(n15618), .B(n15617), .ZN(
        P1_U2829) );
  AOI21_X1 U18904 ( .B1(n19857), .B2(n15619), .A(P1_REIP_REG_10__SCAN_IN), 
        .ZN(n15628) );
  INV_X1 U18905 ( .A(n15620), .ZN(n15767) );
  AOI22_X1 U18906 ( .A1(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n19861), .B1(
        n19856), .B2(n15767), .ZN(n15621) );
  INV_X1 U18907 ( .A(n15621), .ZN(n15622) );
  AOI211_X1 U18908 ( .C1(n19850), .C2(P1_EBX_REG_10__SCAN_IN), .A(n13009), .B(
        n15622), .ZN(n15627) );
  INV_X1 U18909 ( .A(n15623), .ZN(n15624) );
  AOI22_X1 U18910 ( .A1(n15625), .A2(n19816), .B1(n15624), .B2(n19860), .ZN(
        n15626) );
  OAI211_X1 U18911 ( .C1(n15629), .C2(n15628), .A(n15627), .B(n15626), .ZN(
        P1_U2830) );
  OAI22_X1 U18912 ( .A1(n15632), .A2(n15631), .B1(n15630), .B2(n14120), .ZN(
        n15633) );
  INV_X1 U18913 ( .A(n15633), .ZN(n15634) );
  OAI21_X1 U18914 ( .B1(n19879), .B2(n15635), .A(n15634), .ZN(P1_U2848) );
  AOI22_X1 U18915 ( .A1(n15647), .A2(n19876), .B1(n15712), .B2(n19875), .ZN(
        n15636) );
  OAI21_X1 U18916 ( .B1(n19879), .B2(n15637), .A(n15636), .ZN(P1_U2850) );
  AOI22_X1 U18917 ( .A1(n15652), .A2(n19876), .B1(n19875), .B2(n15638), .ZN(
        n15639) );
  OAI21_X1 U18918 ( .B1(n19879), .B2(n15640), .A(n15639), .ZN(P1_U2852) );
  AOI22_X1 U18919 ( .A1(n15670), .A2(n19876), .B1(n19875), .B2(n15641), .ZN(
        n15642) );
  OAI21_X1 U18920 ( .B1(n19879), .B2(n15643), .A(n15642), .ZN(P1_U2860) );
  AOI22_X1 U18921 ( .A1(n19938), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B1(
        n13009), .B2(P1_REIP_REG_22__SCAN_IN), .ZN(n15649) );
  NAND2_X1 U18922 ( .A1(n15645), .A2(n15644), .ZN(n15646) );
  XNOR2_X1 U18923 ( .A(n15646), .B(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15713) );
  AOI22_X1 U18924 ( .A1(n15647), .A2(n9727), .B1(n19944), .B2(n15713), .ZN(
        n15648) );
  OAI211_X1 U18925 ( .C1(n15701), .C2(n15650), .A(n15649), .B(n15648), .ZN(
        P1_U2977) );
  AOI22_X1 U18926 ( .A1(n19938), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B1(
        n13009), .B2(P1_REIP_REG_20__SCAN_IN), .ZN(n15654) );
  AOI22_X1 U18927 ( .A1(n15652), .A2(n9727), .B1(n15651), .B2(n19944), .ZN(
        n15653) );
  OAI211_X1 U18928 ( .C1(n15701), .C2(n15655), .A(n15654), .B(n15653), .ZN(
        P1_U2979) );
  AOI22_X1 U18929 ( .A1(n19938), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B1(
        n13009), .B2(P1_REIP_REG_16__SCAN_IN), .ZN(n15663) );
  OAI21_X1 U18930 ( .B1(n15658), .B2(n15657), .A(n15656), .ZN(n15660) );
  XNOR2_X1 U18931 ( .A(n15660), .B(n15659), .ZN(n15738) );
  AOI22_X1 U18932 ( .A1(n15738), .A2(n19944), .B1(n9727), .B2(n15661), .ZN(
        n15662) );
  OAI211_X1 U18933 ( .C1(n15701), .C2(n15664), .A(n15663), .B(n15662), .ZN(
        P1_U2983) );
  AOI22_X1 U18934 ( .A1(n19938), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        n13009), .B2(P1_REIP_REG_14__SCAN_IN), .ZN(n15668) );
  AOI22_X1 U18935 ( .A1(n15666), .A2(n9727), .B1(n15672), .B2(n15665), .ZN(
        n15667) );
  OAI211_X1 U18936 ( .C1(n15669), .C2(n19764), .A(n15668), .B(n15667), .ZN(
        P1_U2985) );
  AOI22_X1 U18937 ( .A1(n19938), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        n13009), .B2(P1_REIP_REG_12__SCAN_IN), .ZN(n15674) );
  AOI22_X1 U18938 ( .A1(n15672), .A2(n15671), .B1(n9727), .B2(n15670), .ZN(
        n15673) );
  OAI211_X1 U18939 ( .C1(n15675), .C2(n19764), .A(n15674), .B(n15673), .ZN(
        P1_U2987) );
  AOI22_X1 U18940 ( .A1(n19938), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B1(
        n13009), .B2(P1_REIP_REG_11__SCAN_IN), .ZN(n15683) );
  NOR2_X1 U18941 ( .A1(n15676), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n15679) );
  NOR2_X1 U18942 ( .A1(n15677), .A2(n14209), .ZN(n15678) );
  MUX2_X1 U18943 ( .A(n15679), .B(n15678), .S(n9750), .Z(n15680) );
  XNOR2_X1 U18944 ( .A(n15680), .B(n14210), .ZN(n15763) );
  AOI22_X1 U18945 ( .A1(n19944), .A2(n15763), .B1(n9727), .B2(n15681), .ZN(
        n15682) );
  OAI211_X1 U18946 ( .C1(n15701), .C2(n15684), .A(n15683), .B(n15682), .ZN(
        P1_U2988) );
  AOI22_X1 U18947 ( .A1(n19938), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B1(
        n13009), .B2(P1_REIP_REG_7__SCAN_IN), .ZN(n15689) );
  XNOR2_X1 U18948 ( .A(n15685), .B(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15686) );
  XNOR2_X1 U18949 ( .A(n15687), .B(n15686), .ZN(n15783) );
  AOI22_X1 U18950 ( .A1(n15783), .A2(n19944), .B1(n9727), .B2(n19809), .ZN(
        n15688) );
  OAI211_X1 U18951 ( .C1(n15701), .C2(n19807), .A(n15689), .B(n15688), .ZN(
        P1_U2992) );
  AOI22_X1 U18952 ( .A1(n19938), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B1(
        n13009), .B2(P1_REIP_REG_6__SCAN_IN), .ZN(n15694) );
  XNOR2_X1 U18953 ( .A(n15690), .B(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n15691) );
  XNOR2_X1 U18954 ( .A(n15692), .B(n15691), .ZN(n15793) );
  AOI22_X1 U18955 ( .A1(n15793), .A2(n19944), .B1(n9727), .B2(n19872), .ZN(
        n15693) );
  OAI211_X1 U18956 ( .C1(n15701), .C2(n19813), .A(n15694), .B(n15693), .ZN(
        P1_U2993) );
  AOI22_X1 U18957 ( .A1(n19938), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .B1(
        n13009), .B2(P1_REIP_REG_5__SCAN_IN), .ZN(n15700) );
  OAI21_X1 U18958 ( .B1(n15697), .B2(n15696), .A(n15695), .ZN(n15698) );
  INV_X1 U18959 ( .A(n15698), .ZN(n15804) );
  AOI22_X1 U18960 ( .A1(n15804), .A2(n19944), .B1(n9727), .B2(n19832), .ZN(
        n15699) );
  OAI211_X1 U18961 ( .C1(n15701), .C2(n19830), .A(n15700), .B(n15699), .ZN(
        P1_U2994) );
  INV_X1 U18962 ( .A(n15702), .ZN(n15710) );
  AOI22_X1 U18963 ( .A1(P1_REIP_REG_23__SCAN_IN), .A2(n13009), .B1(n15703), 
        .B2(n15709), .ZN(n15708) );
  INV_X1 U18964 ( .A(n15704), .ZN(n15706) );
  AOI22_X1 U18965 ( .A1(n15706), .A2(n19994), .B1(n19993), .B2(n15705), .ZN(
        n15707) );
  OAI211_X1 U18966 ( .C1(n15710), .C2(n15709), .A(n15708), .B(n15707), .ZN(
        P1_U3008) );
  AOI22_X1 U18967 ( .A1(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n15711), .B1(
        n13009), .B2(P1_REIP_REG_22__SCAN_IN), .ZN(n15718) );
  AOI22_X1 U18968 ( .A1(n15713), .A2(n19994), .B1(n19993), .B2(n15712), .ZN(
        n15717) );
  OAI211_X1 U18969 ( .C1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A(n15715), .B(n15714), .ZN(
        n15716) );
  NAND3_X1 U18970 ( .A1(n15718), .A2(n15717), .A3(n15716), .ZN(P1_U3009) );
  AOI22_X1 U18971 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n9908), .B1(
        n13009), .B2(P1_REIP_REG_19__SCAN_IN), .ZN(n15724) );
  AOI22_X1 U18972 ( .A1(n15722), .A2(n19994), .B1(n15721), .B2(n15720), .ZN(
        n15723) );
  OAI211_X1 U18973 ( .C1(n15807), .C2(n15725), .A(n15724), .B(n15723), .ZN(
        P1_U3012) );
  OAI21_X1 U18974 ( .B1(n15735), .B2(n15745), .A(n13911), .ZN(n15728) );
  AOI22_X1 U18975 ( .A1(n15729), .A2(n19994), .B1(n15728), .B2(n15727), .ZN(
        n15731) );
  NAND2_X1 U18976 ( .A1(n13009), .A2(P1_REIP_REG_17__SCAN_IN), .ZN(n15730) );
  OAI211_X1 U18977 ( .C1(n15807), .C2(n15732), .A(n15731), .B(n15730), .ZN(
        P1_U3014) );
  INV_X1 U18978 ( .A(n15733), .ZN(n15755) );
  AOI21_X1 U18979 ( .B1(n15734), .B2(n19988), .A(n15755), .ZN(n15743) );
  INV_X1 U18980 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15741) );
  AOI21_X1 U18981 ( .B1(n15744), .B2(n15741), .A(n15745), .ZN(n15736) );
  AOI22_X1 U18982 ( .A1(n13009), .A2(P1_REIP_REG_16__SCAN_IN), .B1(n15736), 
        .B2(n15735), .ZN(n15740) );
  AOI22_X1 U18983 ( .A1(n15738), .A2(n19994), .B1(n19993), .B2(n15737), .ZN(
        n15739) );
  OAI211_X1 U18984 ( .C1(n15743), .C2(n15741), .A(n15740), .B(n15739), .ZN(
        P1_U3015) );
  NAND2_X1 U18985 ( .A1(n13009), .A2(P1_REIP_REG_15__SCAN_IN), .ZN(n15742) );
  OAI221_X1 U18986 ( .B1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n15745), 
        .C1(n15744), .C2(n15743), .A(n15742), .ZN(n15746) );
  AOI21_X1 U18987 ( .B1(n15747), .B2(n19994), .A(n15746), .ZN(n15748) );
  OAI21_X1 U18988 ( .B1(n15807), .B2(n15749), .A(n15748), .ZN(P1_U3016) );
  NOR3_X1 U18989 ( .A1(n15751), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A3(
        n15750), .ZN(n15753) );
  NOR2_X1 U18990 ( .A1(n19845), .A2(n20619), .ZN(n15752) );
  AOI211_X1 U18991 ( .C1(n15754), .C2(n19994), .A(n15753), .B(n15752), .ZN(
        n15758) );
  OAI21_X1 U18992 ( .B1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n15756), .A(
        n15755), .ZN(n15757) );
  OAI211_X1 U18993 ( .C1(n15759), .C2(n15807), .A(n15758), .B(n15757), .ZN(
        P1_U3018) );
  OAI22_X1 U18994 ( .A1(n15761), .A2(n14210), .B1(n15796), .B2(n15760), .ZN(
        n15762) );
  AOI21_X1 U18995 ( .B1(n15763), .B2(n19994), .A(n15762), .ZN(n15765) );
  NAND2_X1 U18996 ( .A1(n13009), .A2(P1_REIP_REG_11__SCAN_IN), .ZN(n15764) );
  OAI211_X1 U18997 ( .C1(n15807), .C2(n15766), .A(n15765), .B(n15764), .ZN(
        P1_U3020) );
  AOI22_X1 U18998 ( .A1(n13009), .A2(P1_REIP_REG_10__SCAN_IN), .B1(n19993), 
        .B2(n15767), .ZN(n15773) );
  AOI22_X1 U18999 ( .A1(n15769), .A2(n19994), .B1(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n15768), .ZN(n15772) );
  OAI221_X1 U19000 ( .B1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .C1(n14209), .C2(n13403), .A(
        n15770), .ZN(n15771) );
  NAND3_X1 U19001 ( .A1(n15773), .A2(n15772), .A3(n15771), .ZN(P1_U3021) );
  INV_X1 U19002 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n15781) );
  OR2_X1 U19003 ( .A1(n19948), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n15800) );
  AOI221_X1 U19004 ( .B1(n19969), .B2(n19963), .C1(n19948), .C2(n19963), .A(
        n15774), .ZN(n15802) );
  OAI21_X1 U19005 ( .B1(n14496), .B2(n15800), .A(n15802), .ZN(n15792) );
  AOI21_X1 U19006 ( .B1(n15781), .B2(n19988), .A(n15792), .ZN(n15785) );
  INV_X1 U19007 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n15780) );
  AOI22_X1 U19008 ( .A1(n13009), .A2(P1_REIP_REG_8__SCAN_IN), .B1(n19993), 
        .B2(n19795), .ZN(n15779) );
  NAND2_X1 U19009 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n15776) );
  INV_X1 U19010 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n15786) );
  AOI211_X1 U19011 ( .C1(n15780), .C2(n15786), .A(n15781), .B(n15796), .ZN(
        n15775) );
  AOI22_X1 U19012 ( .A1(n15777), .A2(n19994), .B1(n15776), .B2(n15775), .ZN(
        n15778) );
  OAI211_X1 U19013 ( .C1(n15785), .C2(n15780), .A(n15779), .B(n15778), .ZN(
        P1_U3023) );
  OR2_X1 U19014 ( .A1(n15781), .A2(n15796), .ZN(n15787) );
  OAI22_X1 U19015 ( .A1(n15807), .A2(n19812), .B1(n20609), .B2(n19845), .ZN(
        n15782) );
  AOI21_X1 U19016 ( .B1(n15783), .B2(n19994), .A(n15782), .ZN(n15784) );
  OAI221_X1 U19017 ( .B1(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n15787), .C1(
        n15786), .C2(n15785), .A(n15784), .ZN(P1_U3024) );
  INV_X1 U19018 ( .A(n15788), .ZN(n15791) );
  INV_X1 U19019 ( .A(n15789), .ZN(n15790) );
  AOI21_X1 U19020 ( .B1(n15791), .B2(n15790), .A(n9848), .ZN(n19871) );
  AOI22_X1 U19021 ( .A1(n13009), .A2(P1_REIP_REG_6__SCAN_IN), .B1(n19993), 
        .B2(n19871), .ZN(n15795) );
  AOI22_X1 U19022 ( .A1(n15793), .A2(n19994), .B1(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n15792), .ZN(n15794) );
  OAI211_X1 U19023 ( .C1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .C2(n15796), .A(
        n15795), .B(n15794), .ZN(P1_U3025) );
  INV_X1 U19024 ( .A(n15797), .ZN(n15799) );
  NAND2_X1 U19025 ( .A1(n15799), .A2(n15798), .ZN(n19960) );
  OAI22_X1 U19026 ( .A1(n15802), .A2(n15801), .B1(n15800), .B2(n19960), .ZN(
        n15803) );
  AOI21_X1 U19027 ( .B1(n15804), .B2(n19994), .A(n15803), .ZN(n15806) );
  NAND2_X1 U19028 ( .A1(n13009), .A2(P1_REIP_REG_5__SCAN_IN), .ZN(n15805) );
  OAI211_X1 U19029 ( .C1(n15807), .C2(n19835), .A(n15806), .B(n15805), .ZN(
        P1_U3026) );
  INV_X1 U19030 ( .A(n19847), .ZN(n15811) );
  NAND4_X1 U19031 ( .A1(n15811), .A2(n15810), .A3(n15809), .A4(n15808), .ZN(
        n15812) );
  OAI21_X1 U19032 ( .B1(n15814), .B2(n15813), .A(n15812), .ZN(P1_U3468) );
  NAND4_X1 U19033 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(
        P1_STATE2_REG_0__SCAN_IN), .A3(n12396), .A4(n20666), .ZN(n15815) );
  OAI21_X1 U19034 ( .B1(n15816), .B2(n20439), .A(n15815), .ZN(n20577) );
  OAI21_X1 U19035 ( .B1(n15818), .B2(n20577), .A(n15817), .ZN(n15819) );
  OAI221_X1 U19036 ( .B1(n15820), .B2(n20275), .C1(n15820), .C2(n20666), .A(
        n15819), .ZN(n15821) );
  AOI221_X1 U19037 ( .B1(n15823), .B2(n20898), .C1(n15822), .C2(n20898), .A(
        n15821), .ZN(P1_U3162) );
  NOR2_X1 U19038 ( .A1(n15823), .A2(n15822), .ZN(n15825) );
  OAI22_X1 U19039 ( .A1(n20275), .A2(n15825), .B1(n15824), .B2(n15822), .ZN(
        P1_U3466) );
  INV_X1 U19040 ( .A(n15827), .ZN(n15828) );
  OAI22_X1 U19041 ( .A1(n15828), .A2(n18923), .B1(n19672), .B2(n18848), .ZN(
        n15832) );
  OAI22_X1 U19042 ( .A1(n15830), .A2(n15829), .B1(n11698), .B2(n18911), .ZN(
        n15831) );
  AOI211_X1 U19043 ( .C1(n18917), .C2(n15826), .A(n15832), .B(n15831), .ZN(
        n15840) );
  AOI21_X1 U19044 ( .B1(n15959), .B2(n15834), .A(n15835), .ZN(n15949) );
  INV_X1 U19045 ( .A(n15949), .ZN(n15921) );
  OAI21_X1 U19046 ( .B1(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n15835), .A(
        n15836), .ZN(n15948) );
  AOI21_X1 U19047 ( .B1(n15940), .B2(n15836), .A(n9850), .ZN(n15933) );
  INV_X1 U19048 ( .A(n15933), .ZN(n15902) );
  INV_X1 U19049 ( .A(n15837), .ZN(n15881) );
  INV_X1 U19050 ( .A(n15838), .ZN(n15859) );
  NAND4_X1 U19051 ( .A1(n18794), .A2(n15846), .A3(n18863), .A4(n15845), .ZN(
        n15839) );
  OAI211_X1 U19052 ( .C1(n15841), .C2(n18894), .A(n15840), .B(n15839), .ZN(
        P2_U2824) );
  INV_X1 U19053 ( .A(n18923), .ZN(n18895) );
  AOI22_X1 U19054 ( .A1(n15842), .A2(n18895), .B1(P2_REIP_REG_30__SCAN_IN), 
        .B2(n18918), .ZN(n15850) );
  AOI22_X1 U19055 ( .A1(P2_EBX_REG_30__SCAN_IN), .A2(n18919), .B1(
        P2_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n18882), .ZN(n15849) );
  AOI22_X1 U19056 ( .A1(n15844), .A2(n18925), .B1(n15843), .B2(n18917), .ZN(
        n15848) );
  NAND4_X1 U19057 ( .A1(n15850), .A2(n15849), .A3(n15848), .A4(n15847), .ZN(
        P2_U2825) );
  INV_X1 U19058 ( .A(n15851), .ZN(n15852) );
  OAI22_X1 U19059 ( .A1(n15852), .A2(n18923), .B1(n11697), .B2(n18911), .ZN(
        n15855) );
  INV_X1 U19060 ( .A(P2_EBX_REG_29__SCAN_IN), .ZN(n15853) );
  OAI22_X1 U19061 ( .A1(n18810), .A2(n15853), .B1(n14733), .B2(n18848), .ZN(
        n15854) );
  AOI211_X1 U19062 ( .C1(n15856), .C2(n18917), .A(n15855), .B(n15854), .ZN(
        n15861) );
  OAI211_X1 U19063 ( .C1(n15859), .C2(n15858), .A(n10036), .B(n15857), .ZN(
        n15860) );
  OAI211_X1 U19064 ( .C1(n18894), .C2(n15862), .A(n15861), .B(n15860), .ZN(
        P2_U2826) );
  AOI22_X1 U19065 ( .A1(n15863), .A2(n18895), .B1(P2_REIP_REG_28__SCAN_IN), 
        .B2(n18918), .ZN(n15872) );
  AOI22_X1 U19066 ( .A1(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n18882), .B1(
        P2_EBX_REG_28__SCAN_IN), .B2(n18919), .ZN(n15871) );
  AOI22_X1 U19067 ( .A1(n15865), .A2(n18925), .B1(n15864), .B2(n18917), .ZN(
        n15870) );
  OAI211_X1 U19068 ( .C1(n15868), .C2(n15867), .A(n10036), .B(n15866), .ZN(
        n15869) );
  NAND4_X1 U19069 ( .A1(n15872), .A2(n15871), .A3(n15870), .A4(n15869), .ZN(
        P2_U2827) );
  OAI22_X1 U19070 ( .A1(n15873), .A2(n18923), .B1(n14759), .B2(n18848), .ZN(
        n15877) );
  INV_X1 U19071 ( .A(P2_EBX_REG_27__SCAN_IN), .ZN(n15875) );
  OAI22_X1 U19072 ( .A1(n18810), .A2(n15875), .B1(n15874), .B2(n18911), .ZN(
        n15876) );
  AOI211_X1 U19073 ( .C1(n15878), .C2(n18917), .A(n15877), .B(n15876), .ZN(
        n15883) );
  OAI211_X1 U19074 ( .C1(n15881), .C2(n15880), .A(n10036), .B(n15879), .ZN(
        n15882) );
  OAI211_X1 U19075 ( .C1(n18894), .C2(n15884), .A(n15883), .B(n15882), .ZN(
        P2_U2828) );
  OAI22_X1 U19076 ( .A1(n15885), .A2(n18923), .B1(n20880), .B2(n18848), .ZN(
        n15888) );
  OAI22_X1 U19077 ( .A1(n18810), .A2(n15886), .B1(n10049), .B2(n18911), .ZN(
        n15887) );
  AOI211_X1 U19078 ( .C1(n15889), .C2(n18925), .A(n15888), .B(n15887), .ZN(
        n15894) );
  OAI211_X1 U19079 ( .C1(n15892), .C2(n15891), .A(n10036), .B(n15890), .ZN(
        n15893) );
  OAI211_X1 U19080 ( .C1(n18898), .C2(n15895), .A(n15894), .B(n15893), .ZN(
        P2_U2829) );
  OAI22_X1 U19081 ( .A1(n15896), .A2(n18923), .B1(n11646), .B2(n18848), .ZN(
        n15898) );
  OAI22_X1 U19082 ( .A1(n18810), .A2(n14571), .B1(n15940), .B2(n18911), .ZN(
        n15897) );
  AOI211_X1 U19083 ( .C1(n15899), .C2(n18917), .A(n15898), .B(n15897), .ZN(
        n15904) );
  OAI211_X1 U19084 ( .C1(n15902), .C2(n15901), .A(n10036), .B(n15900), .ZN(
        n15903) );
  OAI211_X1 U19085 ( .C1(n18894), .C2(n15934), .A(n15904), .B(n15903), .ZN(
        P2_U2830) );
  OAI22_X1 U19086 ( .A1(n15905), .A2(n18923), .B1(n10048), .B2(n18911), .ZN(
        n15908) );
  INV_X1 U19087 ( .A(P2_EBX_REG_24__SCAN_IN), .ZN(n15906) );
  OAI22_X1 U19088 ( .A1(n18810), .A2(n15906), .B1(n19659), .B2(n18848), .ZN(
        n15907) );
  AOI211_X1 U19089 ( .C1(n15945), .C2(n18925), .A(n15908), .B(n15907), .ZN(
        n15912) );
  OAI211_X1 U19090 ( .C1(n15948), .C2(n15910), .A(n10036), .B(n15909), .ZN(
        n15911) );
  OAI211_X1 U19091 ( .C1(n18898), .C2(n15913), .A(n15912), .B(n15911), .ZN(
        P2_U2831) );
  AOI22_X1 U19092 ( .A1(P2_REIP_REG_23__SCAN_IN), .A2(n18918), .B1(
        P2_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n18882), .ZN(n15925) );
  AOI22_X1 U19093 ( .A1(n15914), .A2(n18895), .B1(P2_EBX_REG_23__SCAN_IN), 
        .B2(n18919), .ZN(n15924) );
  INV_X1 U19094 ( .A(n16068), .ZN(n15918) );
  OAI21_X1 U19095 ( .B1(n14679), .B2(n15916), .A(n15915), .ZN(n15917) );
  INV_X1 U19096 ( .A(n15917), .ZN(n16066) );
  AOI22_X1 U19097 ( .A1(n15918), .A2(n18925), .B1(n16066), .B2(n18917), .ZN(
        n15923) );
  OAI211_X1 U19098 ( .C1(n15921), .C2(n15920), .A(n10036), .B(n15919), .ZN(
        n15922) );
  NAND4_X1 U19099 ( .A1(n15925), .A2(n15924), .A3(n15923), .A4(n15922), .ZN(
        P2_U2832) );
  AOI22_X1 U19100 ( .A1(n15927), .A2(n15926), .B1(n18934), .B2(
        P2_EAX_REG_23__SCAN_IN), .ZN(n15932) );
  AOI22_X1 U19101 ( .A1(n18929), .A2(BUF2_REG_23__SCAN_IN), .B1(n18931), .B2(
        BUF1_REG_23__SCAN_IN), .ZN(n15931) );
  AOI22_X1 U19102 ( .A1(n15929), .A2(n15928), .B1(n18930), .B2(n16066), .ZN(
        n15930) );
  NAND3_X1 U19103 ( .A1(n15932), .A2(n15931), .A3(n15930), .ZN(P2_U2896) );
  AOI22_X1 U19104 ( .A1(P2_REIP_REG_25__SCAN_IN), .A2(n19033), .B1(n16054), 
        .B2(n15933), .ZN(n15939) );
  INV_X1 U19105 ( .A(n15934), .ZN(n15935) );
  AOI222_X1 U19106 ( .A1(n15937), .A2(n16060), .B1(n16055), .B2(n15936), .C1(
        n19041), .C2(n15935), .ZN(n15938) );
  OAI211_X1 U19107 ( .C1(n15940), .C2(n16064), .A(n15939), .B(n15938), .ZN(
        P2_U2989) );
  AOI22_X1 U19108 ( .A1(P2_REIP_REG_24__SCAN_IN), .A2(n19033), .B1(
        P2_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n19032), .ZN(n15947) );
  INV_X1 U19109 ( .A(n15941), .ZN(n15943) );
  OAI22_X1 U19110 ( .A1(n15943), .A2(n19037), .B1(n19035), .B2(n15942), .ZN(
        n15944) );
  AOI21_X1 U19111 ( .B1(n19041), .B2(n15945), .A(n15944), .ZN(n15946) );
  OAI211_X1 U19112 ( .C1(n19045), .C2(n15948), .A(n15947), .B(n15946), .ZN(
        P2_U2990) );
  AOI22_X1 U19113 ( .A1(P2_REIP_REG_23__SCAN_IN), .A2(n19033), .B1(n16054), 
        .B2(n15949), .ZN(n15958) );
  INV_X1 U19114 ( .A(n15950), .ZN(n15951) );
  AOI21_X1 U19115 ( .B1(n15952), .B2(n15951), .A(n9790), .ZN(n16071) );
  OAI21_X1 U19116 ( .B1(n15955), .B2(n15954), .A(n15953), .ZN(n16069) );
  OAI22_X1 U19117 ( .A1(n16069), .A2(n19037), .B1(n16058), .B2(n16068), .ZN(
        n15956) );
  AOI21_X1 U19118 ( .B1(n16055), .B2(n16071), .A(n15956), .ZN(n15957) );
  OAI211_X1 U19119 ( .C1(n15959), .C2(n16064), .A(n15958), .B(n15957), .ZN(
        P2_U2991) );
  OAI22_X1 U19120 ( .A1(n19656), .A2(n18846), .B1(n19045), .B2(n15960), .ZN(
        n15961) );
  AOI21_X1 U19121 ( .B1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n19032), .A(
        n15961), .ZN(n15965) );
  AOI22_X1 U19122 ( .A1(n15963), .A2(n16060), .B1(n16055), .B2(n15962), .ZN(
        n15964) );
  OAI211_X1 U19123 ( .C1(n16058), .C2(n15966), .A(n15965), .B(n15964), .ZN(
        P2_U2992) );
  AOI22_X1 U19124 ( .A1(P2_REIP_REG_19__SCAN_IN), .A2(n19033), .B1(n16054), 
        .B2(n15967), .ZN(n15978) );
  NAND2_X1 U19125 ( .A1(n15969), .A2(n15968), .ZN(n15974) );
  INV_X1 U19126 ( .A(n15970), .ZN(n15972) );
  OR2_X1 U19127 ( .A1(n15972), .A2(n15971), .ZN(n15973) );
  NAND2_X1 U19128 ( .A1(n14802), .A2(n11625), .ZN(n15975) );
  AND2_X1 U19129 ( .A1(n15976), .A2(n15975), .ZN(n16082) );
  AOI22_X1 U19130 ( .A1(n16082), .A2(n16055), .B1(n19041), .B2(n18722), .ZN(
        n15977) );
  AOI22_X1 U19131 ( .A1(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n19032), .B1(
        n16054), .B2(n18743), .ZN(n15986) );
  AOI22_X1 U19132 ( .A1(n15980), .A2(n16060), .B1(n19041), .B2(n18748), .ZN(
        n15985) );
  MUX2_X1 U19133 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .B(n14821), .S(
        n15981), .Z(n15982) );
  OR2_X1 U19134 ( .A1(n15982), .A2(n19035), .ZN(n15983) );
  NAND4_X1 U19135 ( .A1(n15986), .A2(n15985), .A3(n15984), .A4(n15983), .ZN(
        P2_U2997) );
  AOI22_X1 U19136 ( .A1(P2_REIP_REG_15__SCAN_IN), .A2(n19033), .B1(n16054), 
        .B2(n18771), .ZN(n15995) );
  NAND2_X1 U19137 ( .A1(n15988), .A2(n15987), .ZN(n15989) );
  XNOR2_X1 U19138 ( .A(n15990), .B(n15989), .ZN(n16087) );
  INV_X1 U19139 ( .A(n18776), .ZN(n15993) );
  AOI21_X1 U19140 ( .B1(n14820), .B2(n15992), .A(n15991), .ZN(n16090) );
  AOI222_X1 U19141 ( .A1(n16087), .A2(n16060), .B1(n19041), .B2(n15993), .C1(
        n16055), .C2(n16090), .ZN(n15994) );
  OAI211_X1 U19142 ( .C1(n15996), .C2(n16064), .A(n15995), .B(n15994), .ZN(
        P2_U2999) );
  AOI22_X1 U19143 ( .A1(P2_REIP_REG_13__SCAN_IN), .A2(n19033), .B1(n16054), 
        .B2(n18792), .ZN(n16005) );
  NOR2_X1 U19144 ( .A1(n15998), .A2(n15997), .ZN(n15999) );
  XNOR2_X1 U19145 ( .A(n16000), .B(n15999), .ZN(n16102) );
  OAI21_X1 U19146 ( .B1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n16002), .A(
        n16001), .ZN(n16100) );
  OAI22_X1 U19147 ( .A1(n18797), .A2(n16058), .B1(n16100), .B2(n19035), .ZN(
        n16003) );
  AOI21_X1 U19148 ( .B1(n16102), .B2(n16060), .A(n16003), .ZN(n16004) );
  OAI211_X1 U19149 ( .C1(n16006), .C2(n16064), .A(n16005), .B(n16004), .ZN(
        P2_U3001) );
  AOI22_X1 U19150 ( .A1(P2_REIP_REG_11__SCAN_IN), .A2(n19033), .B1(n16054), 
        .B2(n18816), .ZN(n16020) );
  OR2_X1 U19151 ( .A1(n9976), .A2(n16008), .ZN(n16012) );
  NAND2_X1 U19152 ( .A1(n16010), .A2(n16009), .ZN(n16011) );
  XNOR2_X1 U19153 ( .A(n16012), .B(n16011), .ZN(n16127) );
  INV_X1 U19154 ( .A(n18820), .ZN(n16018) );
  NAND2_X1 U19155 ( .A1(n16014), .A2(n16013), .ZN(n16016) );
  NAND2_X1 U19156 ( .A1(n16016), .A2(n16015), .ZN(n16130) );
  INV_X1 U19157 ( .A(n16130), .ZN(n16017) );
  AOI222_X1 U19158 ( .A1(n16127), .A2(n16060), .B1(n19041), .B2(n16018), .C1(
        n16055), .C2(n16017), .ZN(n16019) );
  OAI211_X1 U19159 ( .C1(n16021), .C2(n16064), .A(n16020), .B(n16019), .ZN(
        P2_U3003) );
  AOI22_X1 U19160 ( .A1(P2_REIP_REG_9__SCAN_IN), .A2(n19033), .B1(n16054), 
        .B2(n18840), .ZN(n16027) );
  INV_X1 U19161 ( .A(n16022), .ZN(n16025) );
  INV_X1 U19162 ( .A(n18844), .ZN(n16023) );
  AOI222_X1 U19163 ( .A1(n16025), .A2(n16055), .B1(n16060), .B2(n16024), .C1(
        n19041), .C2(n16023), .ZN(n16026) );
  OAI211_X1 U19164 ( .C1(n18836), .C2(n16064), .A(n16027), .B(n16026), .ZN(
        P2_U3005) );
  AOI22_X1 U19165 ( .A1(P2_REIP_REG_8__SCAN_IN), .A2(n19033), .B1(
        P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n19032), .ZN(n16032) );
  OAI22_X1 U19166 ( .A1(n16029), .A2(n19035), .B1(n16028), .B2(n19037), .ZN(
        n16030) );
  AOI21_X1 U19167 ( .B1(n19041), .B2(n18853), .A(n16030), .ZN(n16031) );
  OAI211_X1 U19168 ( .C1(n19045), .C2(n18851), .A(n16032), .B(n16031), .ZN(
        P2_U3006) );
  AOI22_X1 U19169 ( .A1(P2_REIP_REG_7__SCAN_IN), .A2(n19033), .B1(n16054), 
        .B2(n18865), .ZN(n16038) );
  INV_X1 U19170 ( .A(n16033), .ZN(n16034) );
  AOI222_X1 U19171 ( .A1(n16036), .A2(n16060), .B1(n19041), .B2(n16035), .C1(
        n16055), .C2(n16034), .ZN(n16037) );
  OAI211_X1 U19172 ( .C1(n18860), .C2(n16064), .A(n16038), .B(n16037), .ZN(
        P2_U3007) );
  AOI22_X1 U19173 ( .A1(P2_REIP_REG_6__SCAN_IN), .A2(n19033), .B1(
        P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n19032), .ZN(n16043) );
  OAI22_X1 U19174 ( .A1(n16040), .A2(n19035), .B1(n16039), .B2(n19037), .ZN(
        n16041) );
  AOI21_X1 U19175 ( .B1(n19041), .B2(n18877), .A(n16041), .ZN(n16042) );
  OAI211_X1 U19176 ( .C1(n19045), .C2(n18875), .A(n16043), .B(n16042), .ZN(
        P2_U3008) );
  AOI22_X1 U19177 ( .A1(P2_REIP_REG_5__SCAN_IN), .A2(n19033), .B1(n16054), 
        .B2(n18888), .ZN(n16051) );
  XOR2_X1 U19178 ( .A(n16044), .B(n16045), .Z(n16144) );
  NAND2_X1 U19179 ( .A1(n16047), .A2(n16046), .ZN(n16048) );
  XNOR2_X1 U19180 ( .A(n16049), .B(n16048), .ZN(n16143) );
  INV_X1 U19181 ( .A(n18893), .ZN(n16142) );
  AOI222_X1 U19182 ( .A1(n16144), .A2(n16060), .B1(n16055), .B2(n16143), .C1(
        n19041), .C2(n16142), .ZN(n16050) );
  OAI211_X1 U19183 ( .C1(n16052), .C2(n16064), .A(n16051), .B(n16050), .ZN(
        P2_U3009) );
  AOI22_X1 U19184 ( .A1(P2_REIP_REG_3__SCAN_IN), .A2(n19033), .B1(n16054), 
        .B2(n16053), .ZN(n16063) );
  NAND3_X1 U19185 ( .A1(n16056), .A2(n16055), .A3(n12934), .ZN(n16057) );
  OAI21_X1 U19186 ( .B1(n16058), .B2(n11119), .A(n16057), .ZN(n16059) );
  AOI21_X1 U19187 ( .B1(n16061), .B2(n16060), .A(n16059), .ZN(n16062) );
  OAI211_X1 U19188 ( .C1(n16065), .C2(n16064), .A(n16063), .B(n16062), .ZN(
        P2_U3011) );
  AOI22_X1 U19189 ( .A1(n16067), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .B1(
        n19059), .B2(n16066), .ZN(n16077) );
  OAI22_X1 U19190 ( .A1(n16069), .A2(n16139), .B1(n19061), .B2(n16068), .ZN(
        n16070) );
  AOI21_X1 U19191 ( .B1(n16157), .B2(n16071), .A(n16070), .ZN(n16076) );
  NAND2_X1 U19192 ( .A1(P2_REIP_REG_23__SCAN_IN), .A2(n19033), .ZN(n16075) );
  OAI211_X1 U19193 ( .C1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(n16073), .B(n16072), .ZN(
        n16074) );
  NAND4_X1 U19194 ( .A1(n16077), .A2(n16076), .A3(n16075), .A4(n16074), .ZN(
        P2_U3023) );
  NAND2_X1 U19195 ( .A1(P2_REIP_REG_19__SCAN_IN), .A2(n19033), .ZN(n16078) );
  OAI221_X1 U19196 ( .B1(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n16080), 
        .C1(n11625), .C2(n16079), .A(n16078), .ZN(n16081) );
  AOI21_X1 U19197 ( .B1(n18721), .B2(n19059), .A(n16081), .ZN(n16084) );
  AOI22_X1 U19198 ( .A1(n16082), .A2(n16157), .B1(n16154), .B2(n18722), .ZN(
        n16083) );
  OAI211_X1 U19199 ( .C1(n16139), .C2(n16085), .A(n16084), .B(n16083), .ZN(
        P2_U3027) );
  AOI22_X1 U19200 ( .A1(n16086), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .B1(
        n19059), .B2(n18773), .ZN(n16096) );
  INV_X1 U19201 ( .A(n16087), .ZN(n16088) );
  OAI22_X1 U19202 ( .A1(n16088), .A2(n16139), .B1(n19061), .B2(n18776), .ZN(
        n16089) );
  AOI21_X1 U19203 ( .B1(n16157), .B2(n16090), .A(n16089), .ZN(n16095) );
  NAND2_X1 U19204 ( .A1(P2_REIP_REG_15__SCAN_IN), .A2(n19033), .ZN(n16094) );
  INV_X1 U19205 ( .A(n16091), .ZN(n16092) );
  NAND3_X1 U19206 ( .A1(n16092), .A2(n16111), .A3(n14820), .ZN(n16093) );
  NAND4_X1 U19207 ( .A1(n16096), .A2(n16095), .A3(n16094), .A4(n16093), .ZN(
        P2_U3031) );
  AOI21_X1 U19208 ( .B1(n16099), .B2(n16098), .A(n16097), .ZN(n18938) );
  AOI22_X1 U19209 ( .A1(n16110), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .B1(
        n19059), .B2(n18938), .ZN(n16108) );
  OAI22_X1 U19210 ( .A1(n18797), .A2(n19061), .B1(n16100), .B2(n19056), .ZN(
        n16101) );
  AOI21_X1 U19211 ( .B1(n16102), .B2(n19065), .A(n16101), .ZN(n16107) );
  NAND2_X1 U19212 ( .A1(P2_REIP_REG_13__SCAN_IN), .A2(n19033), .ZN(n16106) );
  INV_X1 U19213 ( .A(n16103), .ZN(n16104) );
  OAI211_X1 U19214 ( .C1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A(n16111), .B(n16104), .ZN(
        n16105) );
  NAND4_X1 U19215 ( .A1(n16108), .A2(n16107), .A3(n16106), .A4(n16105), .ZN(
        P2_U3033) );
  OAI22_X1 U19216 ( .A1(n16131), .A2(n18808), .B1(n11594), .B2(n18846), .ZN(
        n16109) );
  AOI221_X1 U19217 ( .B1(n16111), .B2(n11335), .C1(n16110), .C2(
        P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A(n16109), .ZN(n16114) );
  AOI22_X1 U19218 ( .A1(n16112), .A2(n16157), .B1(n16154), .B2(n18805), .ZN(
        n16113) );
  OAI211_X1 U19219 ( .C1(n16115), .C2(n16139), .A(n16114), .B(n16113), .ZN(
        P2_U3034) );
  AOI21_X1 U19220 ( .B1(n16118), .B2(n16117), .A(n16116), .ZN(n18940) );
  NOR2_X1 U19221 ( .A1(n18846), .A2(n11591), .ZN(n16125) );
  OAI21_X1 U19222 ( .B1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n16163), .A(
        n16119), .ZN(n16133) );
  NOR2_X1 U19223 ( .A1(n16121), .A2(n16120), .ZN(n16135) );
  AOI22_X1 U19224 ( .A1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n16133), .B1(
        n16135), .B2(n16122), .ZN(n16123) );
  AOI21_X1 U19225 ( .B1(n16134), .B2(n16013), .A(n16123), .ZN(n16124) );
  AOI211_X1 U19226 ( .C1(n19059), .C2(n18940), .A(n16125), .B(n16124), .ZN(
        n16129) );
  NOR2_X1 U19227 ( .A1(n18820), .A2(n19061), .ZN(n16126) );
  AOI21_X1 U19228 ( .B1(n16127), .B2(n19065), .A(n16126), .ZN(n16128) );
  OAI211_X1 U19229 ( .C1(n19056), .C2(n16130), .A(n16129), .B(n16128), .ZN(
        P2_U3035) );
  OAI22_X1 U19230 ( .A1(n16131), .A2(n18833), .B1(n11585), .B2(n18846), .ZN(
        n16132) );
  AOI221_X1 U19231 ( .B1(n16135), .B2(n16134), .C1(n16133), .C2(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A(n16132), .ZN(n16138) );
  AOI22_X1 U19232 ( .A1(n16136), .A2(n16157), .B1(n16154), .B2(n18830), .ZN(
        n16137) );
  OAI211_X1 U19233 ( .C1(n16140), .C2(n16139), .A(n16138), .B(n16137), .ZN(
        P2_U3036) );
  AOI22_X1 U19234 ( .A1(n16141), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .B1(
        n19059), .B2(n18890), .ZN(n16151) );
  AOI222_X1 U19235 ( .A1(n16144), .A2(n19065), .B1(n16157), .B2(n16143), .C1(
        n16154), .C2(n16142), .ZN(n16150) );
  NAND2_X1 U19236 ( .A1(P2_REIP_REG_5__SCAN_IN), .A2(n19033), .ZN(n16149) );
  OAI221_X1 U19237 ( .B1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .C1(n16147), .C2(n16146), .A(
        n16145), .ZN(n16148) );
  NAND4_X1 U19238 ( .A1(n16151), .A2(n16150), .A3(n16149), .A4(n16148), .ZN(
        P2_U3041) );
  AOI22_X1 U19239 ( .A1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n19049), .B1(
        n19065), .B2(n16152), .ZN(n16162) );
  AOI21_X1 U19240 ( .B1(n19059), .B2(n18916), .A(n16153), .ZN(n16160) );
  NAND2_X1 U19241 ( .A1(n18926), .A2(n16154), .ZN(n16159) );
  INV_X1 U19242 ( .A(n16155), .ZN(n16156) );
  NAND2_X1 U19243 ( .A1(n16157), .A2(n16156), .ZN(n16158) );
  AND3_X1 U19244 ( .A1(n16160), .A2(n16159), .A3(n16158), .ZN(n16161) );
  OAI211_X1 U19245 ( .C1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(n16163), .A(
        n16162), .B(n16161), .ZN(P2_U3046) );
  MUX2_X1 U19246 ( .A(n16164), .B(n16183), .S(n16180), .Z(n16193) );
  NOR2_X1 U19247 ( .A1(n16180), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n16165) );
  AOI21_X1 U19248 ( .B1(n16166), .B2(n16180), .A(n16165), .ZN(n16192) );
  AOI22_X1 U19249 ( .A1(n16172), .A2(n16169), .B1(n16168), .B2(n16167), .ZN(
        n16170) );
  OAI21_X1 U19250 ( .B1(n16172), .B2(n16171), .A(n16170), .ZN(n19727) );
  OAI21_X1 U19251 ( .B1(P2_MORE_REG_SCAN_IN), .B2(P2_FLUSH_REG_SCAN_IN), .A(
        n16173), .ZN(n16175) );
  OAI211_X1 U19252 ( .C1(n16176), .C2(n11451), .A(n16175), .B(n16174), .ZN(
        n16177) );
  NOR2_X1 U19253 ( .A1(n19727), .A2(n16177), .ZN(n16178) );
  OAI21_X1 U19254 ( .B1(n16180), .B2(n16179), .A(n16178), .ZN(n16191) );
  INV_X1 U19255 ( .A(n16180), .ZN(n16185) );
  OAI211_X1 U19256 ( .C1(n16186), .C2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B(n16181), .ZN(n16182) );
  OAI21_X1 U19257 ( .B1(n16183), .B2(n19704), .A(n16182), .ZN(n16184) );
  AOI211_X1 U19258 ( .C1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .C2(n16186), .A(
        n16185), .B(n16184), .ZN(n16187) );
  OAI21_X1 U19259 ( .B1(n16192), .B2(n19697), .A(n16187), .ZN(n16189) );
  AOI22_X1 U19260 ( .A1(n16192), .A2(n19697), .B1(n16193), .B2(n19096), .ZN(
        n16188) );
  AOI21_X1 U19261 ( .B1(n16189), .B2(n16188), .A(
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n16190) );
  AOI211_X1 U19262 ( .C1(n16193), .C2(n16192), .A(n16191), .B(n16190), .ZN(
        n16205) );
  INV_X1 U19263 ( .A(n19729), .ZN(n16197) );
  AOI211_X1 U19264 ( .C1(n16197), .C2(n16196), .A(n16195), .B(n16194), .ZN(
        n16204) );
  NOR3_X1 U19265 ( .A1(n16198), .A2(n19734), .A3(n19744), .ZN(n16200) );
  OAI221_X1 U19266 ( .B1(n18954), .B2(n16205), .C1(n18954), .C2(n13196), .A(
        n16200), .ZN(n19613) );
  INV_X1 U19267 ( .A(n19613), .ZN(n16202) );
  INV_X1 U19268 ( .A(n19736), .ZN(n19745) );
  AOI22_X1 U19269 ( .A1(n19745), .A2(n16200), .B1(n19746), .B2(n16199), .ZN(
        n16201) );
  AOI22_X1 U19270 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n16202), .B1(n16201), 
        .B2(n18954), .ZN(n16203) );
  OAI211_X1 U19271 ( .C1(n16205), .C2(n19607), .A(n16204), .B(n16203), .ZN(
        P2_U3176) );
  OAI21_X1 U19272 ( .B1(n19714), .B2(n19613), .A(n16206), .ZN(P2_U3593) );
  NOR2_X1 U19273 ( .A1(n17585), .A2(n16209), .ZN(n16217) );
  OAI21_X1 U19274 ( .B1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n17585), .A(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n16210) );
  OAI221_X1 U19275 ( .B1(n16231), .B2(n16211), .C1(n17585), .C2(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A(n16210), .ZN(n16216) );
  OAI21_X1 U19276 ( .B1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n16231), .A(
        n16211), .ZN(n16214) );
  NAND2_X1 U19277 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n17585), .ZN(
        n16212) );
  OAI22_X1 U19278 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n17585), .B1(
        n16212), .B2(n16231), .ZN(n16213) );
  OAI21_X1 U19279 ( .B1(n16217), .B2(n16214), .A(n16213), .ZN(n16215) );
  OAI21_X1 U19280 ( .B1(n16217), .B2(n16216), .A(n16215), .ZN(n16270) );
  INV_X1 U19281 ( .A(n16218), .ZN(n18450) );
  INV_X1 U19282 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n18583) );
  NOR2_X1 U19283 ( .A1(n18583), .A2(n17993), .ZN(n16264) );
  NAND2_X1 U19284 ( .A1(n9867), .A2(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16220) );
  NOR2_X1 U19285 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18666), .ZN(n17387) );
  OR2_X1 U19286 ( .A1(n16220), .A2(n17471), .ZN(n16235) );
  INV_X1 U19287 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n16222) );
  XOR2_X1 U19288 ( .A(n16222), .B(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .Z(
        n16223) );
  NOR2_X1 U19289 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n17424), .ZN(
        n16254) );
  INV_X1 U19290 ( .A(n16253), .ZN(n16399) );
  INV_X1 U19291 ( .A(n17387), .ZN(n18514) );
  NAND2_X1 U19292 ( .A1(n18390), .A2(n16220), .ZN(n16221) );
  OAI211_X1 U19293 ( .C1(n16399), .C2(n18514), .A(n16221), .B(n17674), .ZN(
        n16255) );
  NOR2_X1 U19294 ( .A1(n16254), .A2(n16255), .ZN(n16233) );
  OAI22_X1 U19295 ( .A1(n16235), .A2(n16223), .B1(n16233), .B2(n16222), .ZN(
        n16224) );
  AOI211_X1 U19296 ( .C1(n17470), .C2(n9742), .A(n16264), .B(n16224), .ZN(
        n16228) );
  NOR2_X1 U19297 ( .A1(n18023), .A2(n16381), .ZN(n17667) );
  INV_X1 U19298 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n18611) );
  NAND3_X1 U19299 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(n18611), .ZN(n16262) );
  OAI21_X1 U19300 ( .B1(n16229), .B2(n16231), .A(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n16225) );
  OAI21_X1 U19301 ( .B1(n16278), .B2(n16262), .A(n16225), .ZN(n16266) );
  INV_X1 U19302 ( .A(n17664), .ZN(n17677) );
  NOR2_X2 U19303 ( .A1(n16273), .A2(n17677), .ZN(n17587) );
  OR2_X1 U19304 ( .A1(n16231), .A2(n16230), .ZN(n16226) );
  XNOR2_X1 U19305 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n16226), .ZN(
        n16267) );
  AOI22_X1 U19306 ( .A1(n17667), .A2(n16266), .B1(n17587), .B2(n16267), .ZN(
        n16227) );
  OAI211_X1 U19307 ( .C1(n17493), .C2(n16270), .A(n16228), .B(n16227), .ZN(
        P3_U2799) );
  XOR2_X1 U19308 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B(n16252), .Z(
        n16417) );
  NAND2_X1 U19309 ( .A1(n17667), .A2(n16229), .ZN(n16245) );
  NAND2_X1 U19310 ( .A1(n17587), .A2(n16230), .ZN(n16246) );
  AOI21_X1 U19311 ( .B1(n16245), .B2(n16246), .A(n16231), .ZN(n16237) );
  INV_X1 U19312 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n16234) );
  OAI221_X1 U19313 ( .B1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n16235), .C1(
        n16234), .C2(n16233), .A(n16232), .ZN(n16236) );
  AOI211_X1 U19314 ( .C1(n17470), .C2(n16417), .A(n16237), .B(n16236), .ZN(
        n16243) );
  INV_X1 U19315 ( .A(n17460), .ZN(n17479) );
  NOR2_X1 U19316 ( .A1(n16239), .A2(n17479), .ZN(n17382) );
  NAND3_X1 U19317 ( .A1(n16241), .A2(n16240), .A3(n17382), .ZN(n16242) );
  OAI211_X1 U19318 ( .C1(n16244), .C2(n17493), .A(n16243), .B(n16242), .ZN(
        P3_U2800) );
  AOI21_X1 U19319 ( .B1(n16248), .B2(n16278), .A(n16245), .ZN(n16250) );
  AOI21_X1 U19320 ( .B1(n16248), .B2(n16247), .A(n16246), .ZN(n16249) );
  AOI211_X1 U19321 ( .C1(n17586), .C2(n16251), .A(n16250), .B(n16249), .ZN(
        n16259) );
  AOI21_X1 U19322 ( .B1(n16430), .B2(n16253), .A(n16252), .ZN(n16426) );
  OAI21_X1 U19323 ( .B1(n16254), .B2(n17470), .A(n16426), .ZN(n16257) );
  OAI221_X1 U19324 ( .B1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n9867), .C1(
        P3_PHYADDRPOINTER_REG_29__SCAN_IN), .C2(n18390), .A(n16255), .ZN(
        n16256) );
  NAND4_X1 U19325 ( .A1(n16259), .A2(n16258), .A3(n16257), .A4(n16256), .ZN(
        P3_U2801) );
  OAI21_X1 U19326 ( .B1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n17987), .A(
        n16260), .ZN(n16265) );
  NOR2_X1 U19327 ( .A1(n16262), .A2(n16261), .ZN(n16263) );
  AOI211_X1 U19328 ( .C1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .C2(n16265), .A(
        n16264), .B(n16263), .ZN(n16269) );
  AOI22_X1 U19329 ( .A1(n17911), .A2(n16267), .B1(n17982), .B2(n16266), .ZN(
        n16268) );
  OAI211_X1 U19330 ( .C1(n16270), .C2(n17815), .A(n16269), .B(n16268), .ZN(
        P3_U2831) );
  NAND2_X1 U19331 ( .A1(n16272), .A2(n16271), .ZN(n17308) );
  OAI211_X1 U19332 ( .C1(n16281), .C2(n17321), .A(n17919), .B(n16273), .ZN(
        n16274) );
  OAI22_X1 U19333 ( .A1(n16275), .A2(n17873), .B1(n17307), .B2(n16274), .ZN(
        n16276) );
  AOI211_X1 U19334 ( .C1(n18447), .C2(n16278), .A(n16277), .B(n16276), .ZN(
        n16287) );
  NAND2_X1 U19335 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17993), .ZN(
        n16286) );
  INV_X1 U19336 ( .A(n17873), .ZN(n17733) );
  AOI22_X1 U19337 ( .A1(n18447), .A2(n17807), .B1(n17808), .B2(n17733), .ZN(
        n17786) );
  NOR3_X1 U19338 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17740), .A3(
        n16280), .ZN(n17312) );
  AOI22_X1 U19339 ( .A1(n17979), .A2(P3_REIP_REG_28__SCAN_IN), .B1(n17769), 
        .B2(n17312), .ZN(n16285) );
  OAI221_X1 U19340 ( .B1(n16283), .B2(n16282), .C1(n16283), .C2(n17308), .A(
        n17910), .ZN(n16284) );
  OAI211_X1 U19341 ( .C1(n16287), .C2(n16286), .A(n16285), .B(n16284), .ZN(
        P3_U2834) );
  NOR3_X1 U19342 ( .A1(P3_BE_N_REG_2__SCAN_IN), .A2(P3_W_R_N_REG_SCAN_IN), 
        .A3(P3_BE_N_REG_0__SCAN_IN), .ZN(n16289) );
  NOR4_X1 U19343 ( .A1(P3_BE_N_REG_1__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_D_C_N_REG_SCAN_IN), .A4(P3_ADS_N_REG_SCAN_IN), .ZN(n16288) );
  NAND4_X1 U19344 ( .A1(P3_M_IO_N_REG_SCAN_IN), .A2(n16289), .A3(n16288), .A4(
        U215), .ZN(U213) );
  INV_X1 U19345 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n16292) );
  INV_X2 U19346 ( .A(U214), .ZN(n16338) );
  NOR2_X2 U19347 ( .A1(n16338), .A2(n16290), .ZN(n16339) );
  INV_X1 U19348 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n18955) );
  OAI222_X1 U19349 ( .A1(U214), .A2(n16292), .B1(n16329), .B2(n16291), .C1(
        U212), .C2(n18955), .ZN(U216) );
  AOI222_X1 U19350 ( .A1(n16338), .A2(P1_DATAO_REG_30__SCAN_IN), .B1(n16339), 
        .B2(BUF1_REG_30__SCAN_IN), .C1(n16332), .C2(P2_DATAO_REG_30__SCAN_IN), 
        .ZN(n16293) );
  INV_X1 U19351 ( .A(n16293), .ZN(U217) );
  INV_X1 U19352 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n18961) );
  AOI22_X1 U19353 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n16339), .B1(
        P1_DATAO_REG_29__SCAN_IN), .B2(n16338), .ZN(n16294) );
  OAI21_X1 U19354 ( .B1(n18961), .B2(U212), .A(n16294), .ZN(U218) );
  INV_X1 U19355 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n16296) );
  AOI22_X1 U19356 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(n16332), .B1(
        P1_DATAO_REG_28__SCAN_IN), .B2(n16338), .ZN(n16295) );
  OAI21_X1 U19357 ( .B1(n16296), .B2(n16329), .A(n16295), .ZN(U219) );
  INV_X1 U19358 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n16298) );
  AOI22_X1 U19359 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(n16332), .B1(
        P1_DATAO_REG_27__SCAN_IN), .B2(n16338), .ZN(n16297) );
  OAI21_X1 U19360 ( .B1(n16298), .B2(n16329), .A(n16297), .ZN(U220) );
  INV_X1 U19361 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n16300) );
  AOI22_X1 U19362 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(n16332), .B1(
        P1_DATAO_REG_26__SCAN_IN), .B2(n16338), .ZN(n16299) );
  OAI21_X1 U19363 ( .B1(n16300), .B2(n16329), .A(n16299), .ZN(U221) );
  AOI22_X1 U19364 ( .A1(P2_DATAO_REG_25__SCAN_IN), .A2(n16332), .B1(
        P1_DATAO_REG_25__SCAN_IN), .B2(n16338), .ZN(n16301) );
  OAI21_X1 U19365 ( .B1(n20967), .B2(n16329), .A(n16301), .ZN(U222) );
  AOI22_X1 U19366 ( .A1(P2_DATAO_REG_24__SCAN_IN), .A2(n16332), .B1(
        P1_DATAO_REG_24__SCAN_IN), .B2(n16338), .ZN(n16302) );
  OAI21_X1 U19367 ( .B1(n16303), .B2(n16329), .A(n16302), .ZN(U223) );
  AOI22_X1 U19368 ( .A1(P2_DATAO_REG_23__SCAN_IN), .A2(n16332), .B1(
        P1_DATAO_REG_23__SCAN_IN), .B2(n16338), .ZN(n16304) );
  OAI21_X1 U19369 ( .B1(n14151), .B2(n16329), .A(n16304), .ZN(U224) );
  AOI22_X1 U19370 ( .A1(P2_DATAO_REG_22__SCAN_IN), .A2(n16332), .B1(
        P1_DATAO_REG_22__SCAN_IN), .B2(n16338), .ZN(n16305) );
  OAI21_X1 U19371 ( .B1(n16306), .B2(n16329), .A(n16305), .ZN(U225) );
  AOI22_X1 U19372 ( .A1(P2_DATAO_REG_21__SCAN_IN), .A2(n16332), .B1(
        P1_DATAO_REG_21__SCAN_IN), .B2(n16338), .ZN(n16307) );
  OAI21_X1 U19373 ( .B1(n16308), .B2(n16329), .A(n16307), .ZN(U226) );
  AOI22_X1 U19374 ( .A1(P2_DATAO_REG_20__SCAN_IN), .A2(n16332), .B1(
        P1_DATAO_REG_20__SCAN_IN), .B2(n16338), .ZN(n16309) );
  OAI21_X1 U19375 ( .B1(n19081), .B2(n16329), .A(n16309), .ZN(U227) );
  INV_X1 U19376 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n20944) );
  INV_X1 U19377 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n16310) );
  INV_X1 U19378 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n20963) );
  OAI222_X1 U19379 ( .A1(U214), .A2(n20944), .B1(n16329), .B2(n16310), .C1(
        U212), .C2(n20963), .ZN(U228) );
  AOI22_X1 U19380 ( .A1(P2_DATAO_REG_18__SCAN_IN), .A2(n16332), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(n16338), .ZN(n16311) );
  OAI21_X1 U19381 ( .B1(n14174), .B2(n16329), .A(n16311), .ZN(U229) );
  INV_X1 U19382 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n16313) );
  AOI22_X1 U19383 ( .A1(P2_DATAO_REG_17__SCAN_IN), .A2(n16332), .B1(
        P1_DATAO_REG_17__SCAN_IN), .B2(n16338), .ZN(n16312) );
  OAI21_X1 U19384 ( .B1(n16313), .B2(n16329), .A(n16312), .ZN(U230) );
  AOI22_X1 U19385 ( .A1(P2_DATAO_REG_16__SCAN_IN), .A2(n16332), .B1(
        P1_DATAO_REG_16__SCAN_IN), .B2(n16338), .ZN(n16314) );
  OAI21_X1 U19386 ( .B1(n16315), .B2(n16329), .A(n16314), .ZN(U231) );
  INV_X1 U19387 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n16357) );
  AOI22_X1 U19388 ( .A1(BUF1_REG_15__SCAN_IN), .A2(n16339), .B1(
        P1_DATAO_REG_15__SCAN_IN), .B2(n16338), .ZN(n16316) );
  OAI21_X1 U19389 ( .B1(n16357), .B2(U212), .A(n16316), .ZN(U232) );
  INV_X1 U19390 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n16318) );
  AOI22_X1 U19391 ( .A1(P2_DATAO_REG_14__SCAN_IN), .A2(n16332), .B1(
        P1_DATAO_REG_14__SCAN_IN), .B2(n16338), .ZN(n16317) );
  OAI21_X1 U19392 ( .B1(n16318), .B2(n16329), .A(n16317), .ZN(U233) );
  INV_X1 U19393 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n16320) );
  AOI22_X1 U19394 ( .A1(P2_DATAO_REG_13__SCAN_IN), .A2(n16332), .B1(
        P1_DATAO_REG_13__SCAN_IN), .B2(n16338), .ZN(n16319) );
  OAI21_X1 U19395 ( .B1(n16320), .B2(n16329), .A(n16319), .ZN(U234) );
  INV_X1 U19396 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n16353) );
  AOI22_X1 U19397 ( .A1(BUF1_REG_12__SCAN_IN), .A2(n16339), .B1(
        P1_DATAO_REG_12__SCAN_IN), .B2(n16338), .ZN(n16321) );
  OAI21_X1 U19398 ( .B1(n16353), .B2(U212), .A(n16321), .ZN(U235) );
  INV_X1 U19399 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n16323) );
  AOI22_X1 U19400 ( .A1(P2_DATAO_REG_11__SCAN_IN), .A2(n16332), .B1(
        P1_DATAO_REG_11__SCAN_IN), .B2(n16338), .ZN(n16322) );
  OAI21_X1 U19401 ( .B1(n16323), .B2(n16329), .A(n16322), .ZN(U236) );
  INV_X1 U19402 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n16351) );
  AOI22_X1 U19403 ( .A1(BUF1_REG_10__SCAN_IN), .A2(n16339), .B1(
        P1_DATAO_REG_10__SCAN_IN), .B2(n16338), .ZN(n16324) );
  OAI21_X1 U19404 ( .B1(n16351), .B2(U212), .A(n16324), .ZN(U237) );
  AOI22_X1 U19405 ( .A1(P2_DATAO_REG_9__SCAN_IN), .A2(n16332), .B1(
        P1_DATAO_REG_9__SCAN_IN), .B2(n16338), .ZN(n16325) );
  OAI21_X1 U19406 ( .B1(n16326), .B2(n16329), .A(n16325), .ZN(U238) );
  AOI22_X1 U19407 ( .A1(P2_DATAO_REG_8__SCAN_IN), .A2(n16332), .B1(
        P1_DATAO_REG_8__SCAN_IN), .B2(n16338), .ZN(n16327) );
  OAI21_X1 U19408 ( .B1(n11896), .B2(n16329), .A(n16327), .ZN(U239) );
  INV_X1 U19409 ( .A(BUF1_REG_7__SCAN_IN), .ZN(n16330) );
  AOI22_X1 U19410 ( .A1(P2_DATAO_REG_7__SCAN_IN), .A2(n16332), .B1(
        P1_DATAO_REG_7__SCAN_IN), .B2(n16338), .ZN(n16328) );
  OAI21_X1 U19411 ( .B1(n16330), .B2(n16329), .A(n16328), .ZN(U240) );
  INV_X1 U19412 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n16346) );
  AOI22_X1 U19413 ( .A1(BUF1_REG_6__SCAN_IN), .A2(n16339), .B1(
        P1_DATAO_REG_6__SCAN_IN), .B2(n16338), .ZN(n16331) );
  OAI21_X1 U19414 ( .B1(n16346), .B2(U212), .A(n16331), .ZN(U241) );
  INV_X1 U19415 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n20856) );
  AOI22_X1 U19416 ( .A1(BUF1_REG_5__SCAN_IN), .A2(n16339), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n16332), .ZN(n16333) );
  OAI21_X1 U19417 ( .B1(n20856), .B2(U214), .A(n16333), .ZN(U242) );
  INV_X1 U19418 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n16344) );
  AOI22_X1 U19419 ( .A1(BUF1_REG_4__SCAN_IN), .A2(n16339), .B1(
        P1_DATAO_REG_4__SCAN_IN), .B2(n16338), .ZN(n16334) );
  OAI21_X1 U19420 ( .B1(n16344), .B2(U212), .A(n16334), .ZN(U243) );
  INV_X1 U19421 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n16343) );
  AOI22_X1 U19422 ( .A1(BUF1_REG_3__SCAN_IN), .A2(n16339), .B1(
        P1_DATAO_REG_3__SCAN_IN), .B2(n16338), .ZN(n16335) );
  OAI21_X1 U19423 ( .B1(n16343), .B2(U212), .A(n16335), .ZN(U244) );
  INV_X1 U19424 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n16342) );
  AOI22_X1 U19425 ( .A1(BUF1_REG_2__SCAN_IN), .A2(n16339), .B1(
        P1_DATAO_REG_2__SCAN_IN), .B2(n16338), .ZN(n16336) );
  OAI21_X1 U19426 ( .B1(n16342), .B2(U212), .A(n16336), .ZN(U245) );
  INV_X1 U19427 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n20754) );
  AOI22_X1 U19428 ( .A1(BUF1_REG_1__SCAN_IN), .A2(n16339), .B1(
        P1_DATAO_REG_1__SCAN_IN), .B2(n16338), .ZN(n16337) );
  OAI21_X1 U19429 ( .B1(n20754), .B2(U212), .A(n16337), .ZN(U246) );
  INV_X1 U19430 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n16341) );
  AOI22_X1 U19431 ( .A1(BUF1_REG_0__SCAN_IN), .A2(n16339), .B1(
        P1_DATAO_REG_0__SCAN_IN), .B2(n16338), .ZN(n16340) );
  OAI21_X1 U19432 ( .B1(n16341), .B2(U212), .A(n16340), .ZN(U247) );
  INV_X1 U19433 ( .A(BUF2_REG_0__SCAN_IN), .ZN(n18014) );
  AOI22_X1 U19434 ( .A1(n16371), .A2(n16341), .B1(n18014), .B2(U215), .ZN(U251) );
  INV_X1 U19435 ( .A(BUF2_REG_1__SCAN_IN), .ZN(n18024) );
  AOI22_X1 U19436 ( .A1(n16371), .A2(n20754), .B1(n18024), .B2(U215), .ZN(U252) );
  INV_X1 U19437 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n18028) );
  AOI22_X1 U19438 ( .A1(n16371), .A2(n16342), .B1(n18028), .B2(U215), .ZN(U253) );
  INV_X1 U19439 ( .A(BUF2_REG_3__SCAN_IN), .ZN(n18033) );
  AOI22_X1 U19440 ( .A1(n16371), .A2(n16343), .B1(n18033), .B2(U215), .ZN(U254) );
  INV_X1 U19441 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n18038) );
  AOI22_X1 U19442 ( .A1(n16371), .A2(n16344), .B1(n18038), .B2(U215), .ZN(U255) );
  OAI22_X1 U19443 ( .A1(U215), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n16367), .ZN(n16345) );
  INV_X1 U19444 ( .A(n16345), .ZN(U256) );
  INV_X1 U19445 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n18048) );
  AOI22_X1 U19446 ( .A1(n16371), .A2(n16346), .B1(n18048), .B2(U215), .ZN(U257) );
  INV_X1 U19447 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n16347) );
  INV_X1 U19448 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n18055) );
  AOI22_X1 U19449 ( .A1(n16371), .A2(n16347), .B1(n18055), .B2(U215), .ZN(U258) );
  OAI22_X1 U19450 ( .A1(U215), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n16367), .ZN(n16348) );
  INV_X1 U19451 ( .A(n16348), .ZN(U259) );
  INV_X1 U19452 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n16349) );
  INV_X1 U19453 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n17159) );
  AOI22_X1 U19454 ( .A1(n16371), .A2(n16349), .B1(n17159), .B2(U215), .ZN(U260) );
  INV_X1 U19455 ( .A(BUF2_REG_10__SCAN_IN), .ZN(n16350) );
  AOI22_X1 U19456 ( .A1(n16367), .A2(n16351), .B1(n16350), .B2(U215), .ZN(U261) );
  INV_X1 U19457 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n16352) );
  INV_X1 U19458 ( .A(BUF2_REG_11__SCAN_IN), .ZN(n17149) );
  AOI22_X1 U19459 ( .A1(n16371), .A2(n16352), .B1(n17149), .B2(U215), .ZN(U262) );
  INV_X1 U19460 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n17145) );
  AOI22_X1 U19461 ( .A1(n16367), .A2(n16353), .B1(n17145), .B2(U215), .ZN(U263) );
  INV_X1 U19462 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n16354) );
  INV_X1 U19463 ( .A(BUF2_REG_13__SCAN_IN), .ZN(n17140) );
  AOI22_X1 U19464 ( .A1(n16371), .A2(n16354), .B1(n17140), .B2(U215), .ZN(U264) );
  OAI22_X1 U19465 ( .A1(U215), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n16371), .ZN(n16355) );
  INV_X1 U19466 ( .A(n16355), .ZN(U265) );
  INV_X1 U19467 ( .A(BUF2_REG_15__SCAN_IN), .ZN(n16356) );
  AOI22_X1 U19468 ( .A1(n16371), .A2(n16357), .B1(n16356), .B2(U215), .ZN(U266) );
  INV_X1 U19469 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n16358) );
  AOI22_X1 U19470 ( .A1(n16371), .A2(n16358), .B1(n18018), .B2(U215), .ZN(U267) );
  OAI22_X1 U19471 ( .A1(U215), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n16367), .ZN(n16359) );
  INV_X1 U19472 ( .A(n16359), .ZN(U268) );
  INV_X1 U19473 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n16360) );
  INV_X1 U19474 ( .A(BUF2_REG_18__SCAN_IN), .ZN(n19070) );
  AOI22_X1 U19475 ( .A1(n16367), .A2(n16360), .B1(n19070), .B2(U215), .ZN(U269) );
  INV_X1 U19476 ( .A(BUF2_REG_19__SCAN_IN), .ZN(n18034) );
  AOI22_X1 U19477 ( .A1(n16371), .A2(n20963), .B1(n18034), .B2(U215), .ZN(U270) );
  INV_X1 U19478 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n16361) );
  INV_X1 U19479 ( .A(BUF2_REG_20__SCAN_IN), .ZN(n20770) );
  AOI22_X1 U19480 ( .A1(n16367), .A2(n16361), .B1(n20770), .B2(U215), .ZN(U271) );
  INV_X1 U19481 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n16362) );
  AOI22_X1 U19482 ( .A1(n16371), .A2(n16362), .B1(n18042), .B2(U215), .ZN(U272) );
  INV_X1 U19483 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n16363) );
  INV_X1 U19484 ( .A(BUF2_REG_22__SCAN_IN), .ZN(n18047) );
  AOI22_X1 U19485 ( .A1(n16367), .A2(n16363), .B1(n18047), .B2(U215), .ZN(U273) );
  OAI22_X1 U19486 ( .A1(U215), .A2(P2_DATAO_REG_23__SCAN_IN), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n16371), .ZN(n16364) );
  INV_X1 U19487 ( .A(n16364), .ZN(U274) );
  OAI22_X1 U19488 ( .A1(U215), .A2(P2_DATAO_REG_24__SCAN_IN), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n16367), .ZN(n16365) );
  INV_X1 U19489 ( .A(n16365), .ZN(U275) );
  INV_X1 U19490 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n16366) );
  AOI22_X1 U19491 ( .A1(n16367), .A2(n16366), .B1(n20723), .B2(U215), .ZN(U276) );
  INV_X1 U19492 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n16368) );
  INV_X1 U19493 ( .A(BUF2_REG_26__SCAN_IN), .ZN(n18029) );
  AOI22_X1 U19494 ( .A1(n16371), .A2(n16368), .B1(n18029), .B2(U215), .ZN(U277) );
  OAI22_X1 U19495 ( .A1(U215), .A2(P2_DATAO_REG_27__SCAN_IN), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n16371), .ZN(n16369) );
  INV_X1 U19496 ( .A(n16369), .ZN(U278) );
  OAI22_X1 U19497 ( .A1(U215), .A2(P2_DATAO_REG_28__SCAN_IN), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n16371), .ZN(n16370) );
  INV_X1 U19498 ( .A(n16370), .ZN(U279) );
  INV_X1 U19499 ( .A(BUF2_REG_29__SCAN_IN), .ZN(n18043) );
  AOI22_X1 U19500 ( .A1(n16371), .A2(n18961), .B1(n18043), .B2(U215), .ZN(U280) );
  INV_X1 U19501 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n18958) );
  INV_X1 U19502 ( .A(BUF2_REG_30__SCAN_IN), .ZN(n18049) );
  AOI22_X1 U19503 ( .A1(n16371), .A2(n18958), .B1(n18049), .B2(U215), .ZN(U281) );
  AOI22_X1 U19504 ( .A1(n16371), .A2(n18955), .B1(n18058), .B2(U215), .ZN(U282) );
  INV_X1 U19505 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n16372) );
  INV_X1 U19506 ( .A(P3_DATAO_REG_30__SCAN_IN), .ZN(n20772) );
  OAI222_X1 U19507 ( .A1(P2_DATAO_REG_31__SCAN_IN), .A2(n18958), .B1(
        P1_DATAO_REG_31__SCAN_IN), .B2(n16372), .C1(P3_DATAO_REG_31__SCAN_IN), 
        .C2(n20772), .ZN(n16373) );
  INV_X2 U19508 ( .A(n20676), .ZN(n20677) );
  INV_X1 U19509 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n20869) );
  INV_X1 U19510 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n19642) );
  AOI22_X1 U19511 ( .A1(n20677), .A2(n20869), .B1(n19642), .B2(n20676), .ZN(
        U347) );
  INV_X1 U19512 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n20948) );
  INV_X1 U19513 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n19641) );
  AOI22_X1 U19514 ( .A1(n20677), .A2(n20948), .B1(n19641), .B2(n20676), .ZN(
        U348) );
  INV_X1 U19515 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n18541) );
  INV_X1 U19516 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n19640) );
  AOI22_X1 U19517 ( .A1(n20677), .A2(n18541), .B1(n19640), .B2(n20676), .ZN(
        U349) );
  INV_X1 U19518 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n18540) );
  INV_X1 U19519 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n20804) );
  AOI22_X1 U19520 ( .A1(n20677), .A2(n18540), .B1(n20804), .B2(n20676), .ZN(
        U350) );
  INV_X1 U19521 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n18538) );
  INV_X1 U19522 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n19639) );
  AOI22_X1 U19523 ( .A1(n20677), .A2(n18538), .B1(n19639), .B2(n20676), .ZN(
        U351) );
  INV_X1 U19524 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n18536) );
  INV_X1 U19525 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n19638) );
  AOI22_X1 U19526 ( .A1(n20677), .A2(n18536), .B1(n19638), .B2(n20676), .ZN(
        U352) );
  INV_X1 U19527 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n20803) );
  INV_X1 U19528 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n19637) );
  AOI22_X1 U19529 ( .A1(n20677), .A2(n20803), .B1(n19637), .B2(n20676), .ZN(
        U353) );
  INV_X1 U19530 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n18533) );
  AOI22_X1 U19531 ( .A1(n20677), .A2(n18533), .B1(n19636), .B2(n20676), .ZN(
        U354) );
  INV_X1 U19532 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n18581) );
  INV_X1 U19533 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n19667) );
  AOI22_X1 U19534 ( .A1(n20677), .A2(n18581), .B1(n19667), .B2(n16373), .ZN(
        U356) );
  INV_X1 U19535 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n18577) );
  INV_X1 U19536 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n19666) );
  AOI22_X1 U19537 ( .A1(n20677), .A2(n18577), .B1(n19666), .B2(n16373), .ZN(
        U357) );
  INV_X1 U19538 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n18576) );
  INV_X1 U19539 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n19663) );
  AOI22_X1 U19540 ( .A1(n20677), .A2(n18576), .B1(n19663), .B2(n20676), .ZN(
        U358) );
  INV_X1 U19541 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n18574) );
  INV_X1 U19542 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n19662) );
  AOI22_X1 U19543 ( .A1(n20677), .A2(n18574), .B1(n19662), .B2(n20676), .ZN(
        U359) );
  INV_X1 U19544 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n18572) );
  INV_X1 U19545 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n19661) );
  AOI22_X1 U19546 ( .A1(n20677), .A2(n18572), .B1(n19661), .B2(n20676), .ZN(
        U360) );
  INV_X1 U19547 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n20797) );
  INV_X1 U19548 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n19660) );
  AOI22_X1 U19549 ( .A1(n20677), .A2(n20797), .B1(n19660), .B2(n20676), .ZN(
        U361) );
  INV_X1 U19550 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n18569) );
  INV_X1 U19551 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n19658) );
  AOI22_X1 U19552 ( .A1(n20677), .A2(n18569), .B1(n19658), .B2(n20676), .ZN(
        U362) );
  INV_X1 U19553 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n18568) );
  INV_X1 U19554 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n19657) );
  AOI22_X1 U19555 ( .A1(n20677), .A2(n18568), .B1(n19657), .B2(n20676), .ZN(
        U363) );
  INV_X1 U19556 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n18566) );
  INV_X1 U19557 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n19655) );
  AOI22_X1 U19558 ( .A1(n20677), .A2(n18566), .B1(n19655), .B2(n20676), .ZN(
        U364) );
  INV_X1 U19559 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n18531) );
  INV_X1 U19560 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n19635) );
  AOI22_X1 U19561 ( .A1(n20677), .A2(n18531), .B1(n19635), .B2(n20676), .ZN(
        U365) );
  INV_X1 U19562 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n18563) );
  INV_X1 U19563 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n19653) );
  AOI22_X1 U19564 ( .A1(n20677), .A2(n18563), .B1(n19653), .B2(n16373), .ZN(
        U366) );
  INV_X1 U19565 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n18562) );
  INV_X1 U19566 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n19652) );
  AOI22_X1 U19567 ( .A1(n20677), .A2(n18562), .B1(n19652), .B2(n16373), .ZN(
        U367) );
  INV_X1 U19568 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n18560) );
  INV_X1 U19569 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n19651) );
  AOI22_X1 U19570 ( .A1(n20677), .A2(n18560), .B1(n19651), .B2(n16373), .ZN(
        U368) );
  INV_X1 U19571 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n18557) );
  INV_X1 U19572 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n19649) );
  AOI22_X1 U19573 ( .A1(n20677), .A2(n18557), .B1(n19649), .B2(n16373), .ZN(
        U369) );
  INV_X1 U19574 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n18556) );
  INV_X1 U19575 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n19648) );
  AOI22_X1 U19576 ( .A1(n20677), .A2(n18556), .B1(n19648), .B2(n16373), .ZN(
        U370) );
  INV_X1 U19577 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n18554) );
  INV_X1 U19578 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n19646) );
  AOI22_X1 U19579 ( .A1(n20677), .A2(n18554), .B1(n19646), .B2(n16373), .ZN(
        U371) );
  INV_X1 U19580 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n18551) );
  INV_X1 U19581 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n19645) );
  AOI22_X1 U19582 ( .A1(n20677), .A2(n18551), .B1(n19645), .B2(n20676), .ZN(
        U372) );
  INV_X1 U19583 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n18550) );
  INV_X1 U19584 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n19644) );
  AOI22_X1 U19585 ( .A1(n20677), .A2(n18550), .B1(n19644), .B2(n20676), .ZN(
        U373) );
  INV_X1 U19586 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n18548) );
  INV_X1 U19587 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n19643) );
  AOI22_X1 U19588 ( .A1(n20677), .A2(n18548), .B1(n19643), .B2(n20676), .ZN(
        U374) );
  INV_X1 U19589 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n18546) );
  INV_X1 U19590 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n20729) );
  AOI22_X1 U19591 ( .A1(n20677), .A2(n18546), .B1(n20729), .B2(n20676), .ZN(
        U375) );
  INV_X1 U19592 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n18530) );
  INV_X1 U19593 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n19634) );
  AOI22_X1 U19594 ( .A1(n20677), .A2(n18530), .B1(n19634), .B2(n20676), .ZN(
        U376) );
  INV_X1 U19595 ( .A(P3_ADS_N_REG_SCAN_IN), .ZN(n16374) );
  NOR2_X1 U19596 ( .A1(P3_STATE_REG_2__SCAN_IN), .A2(n20812), .ZN(n20688) );
  OAI21_X1 U19597 ( .B1(n18519), .B2(n20688), .A(n18663), .ZN(n18515) );
  INV_X1 U19598 ( .A(n18515), .ZN(n18595) );
  OAI21_X1 U19599 ( .B1(n16374), .B2(n18519), .A(n18516), .ZN(P3_U2633) );
  INV_X1 U19600 ( .A(n16380), .ZN(n16375) );
  OAI21_X1 U19601 ( .B1(n16375), .B2(n17238), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n16376) );
  OAI21_X1 U19602 ( .B1(n16377), .B2(n18504), .A(n16376), .ZN(P3_U2634) );
  INV_X1 U19603 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n20947) );
  AOI21_X1 U19604 ( .B1(n18519), .B2(n20947), .A(P3_D_C_N_REG_SCAN_IN), .ZN(
        n16378) );
  AOI22_X1 U19605 ( .A1(n18665), .A2(P3_CODEFETCH_REG_SCAN_IN), .B1(n16378), 
        .B2(n18663), .ZN(P3_U2635) );
  NOR2_X1 U19606 ( .A1(P3_STATE_REG_2__SCAN_IN), .A2(P3_STATE_REG_1__SCAN_IN), 
        .ZN(n18517) );
  OAI21_X1 U19607 ( .B1(n18517), .B2(BS16), .A(n18595), .ZN(n18594) );
  OAI21_X1 U19608 ( .B1(n18595), .B2(n18653), .A(n18594), .ZN(P3_U2636) );
  AND3_X1 U19609 ( .A1(n18443), .A2(n16380), .A3(n16379), .ZN(n18491) );
  NOR2_X1 U19610 ( .A1(n18491), .A2(n18495), .ZN(n18643) );
  OAI21_X1 U19611 ( .B1(n18643), .B2(n16382), .A(n16381), .ZN(P3_U2637) );
  NOR4_X1 U19612 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_10__SCAN_IN), .A3(P3_DATAWIDTH_REG_11__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_12__SCAN_IN), .ZN(n16392) );
  NOR4_X1 U19613 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_6__SCAN_IN), .A3(P3_DATAWIDTH_REG_7__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_8__SCAN_IN), .ZN(n16391) );
  NOR2_X1 U19614 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_31__SCAN_IN), .ZN(n20687) );
  AOI211_X1 U19615 ( .C1(P3_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A(P3_DATAWIDTH_REG_3__SCAN_IN), .B(
        P3_DATAWIDTH_REG_4__SCAN_IN), .ZN(n16383) );
  NAND2_X1 U19616 ( .A1(n20687), .A2(n16383), .ZN(n16389) );
  NOR4_X1 U19617 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_19__SCAN_IN), .A3(P3_DATAWIDTH_REG_20__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_21__SCAN_IN), .ZN(n16387) );
  NOR4_X1 U19618 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_13__SCAN_IN), .A3(P3_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_17__SCAN_IN), .ZN(n16386) );
  NOR4_X1 U19619 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_27__SCAN_IN), .A3(P3_DATAWIDTH_REG_28__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_29__SCAN_IN), .ZN(n16385) );
  NOR4_X1 U19620 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_23__SCAN_IN), .A3(P3_DATAWIDTH_REG_25__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_30__SCAN_IN), .ZN(n16384) );
  NAND4_X1 U19621 ( .A1(n16387), .A2(n16386), .A3(n16385), .A4(n16384), .ZN(
        n16388) );
  NOR4_X1 U19622 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_2__SCAN_IN), .A3(n16389), .A4(n16388), .ZN(n16390) );
  NAND3_X1 U19623 ( .A1(n16392), .A2(n16391), .A3(n16390), .ZN(n18635) );
  NOR2_X1 U19624 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n18635), .ZN(n18632) );
  INV_X1 U19625 ( .A(n18635), .ZN(n18640) );
  INV_X1 U19626 ( .A(P3_REIP_REG_0__SCAN_IN), .ZN(n18633) );
  INV_X1 U19627 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20950) );
  INV_X1 U19628 ( .A(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(n18637) );
  NAND4_X1 U19629 ( .A1(n18640), .A2(n18633), .A3(n20950), .A4(n18637), .ZN(
        n16393) );
  INV_X1 U19630 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n18592) );
  AOI22_X1 U19631 ( .A1(n18632), .A2(n16393), .B1(n18635), .B2(n18592), .ZN(
        P3_U2638) );
  INV_X1 U19632 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .ZN(n18589) );
  NAND2_X1 U19633 ( .A1(n18632), .A2(n20950), .ZN(n18638) );
  OAI211_X1 U19634 ( .C1(n18640), .C2(n18589), .A(n16393), .B(n18638), .ZN(
        P3_U2639) );
  AOI22_X1 U19635 ( .A1(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .A2(n16709), .B1(
        P3_EBX_REG_31__SCAN_IN), .B2(n16750), .ZN(n16413) );
  NOR2_X1 U19636 ( .A1(P3_EBX_REG_30__SCAN_IN), .A2(n16711), .ZN(n16409) );
  NAND2_X1 U19637 ( .A1(n16478), .A2(n16758), .ZN(n16477) );
  NOR2_X1 U19638 ( .A1(P3_EBX_REG_25__SCAN_IN), .A2(n16477), .ZN(n16462) );
  NAND2_X1 U19639 ( .A1(n16462), .A2(n16805), .ZN(n16456) );
  NOR2_X1 U19640 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(n16456), .ZN(n16446) );
  NAND2_X1 U19641 ( .A1(n16446), .A2(n16440), .ZN(n16439) );
  NOR2_X1 U19642 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n16439), .ZN(n16423) );
  INV_X1 U19643 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n18580) );
  NAND2_X1 U19644 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .ZN(n16433) );
  NOR2_X1 U19645 ( .A1(n18580), .A2(n16433), .ZN(n16397) );
  NAND2_X1 U19646 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n16394), .ZN(n16396) );
  NAND2_X1 U19647 ( .A1(P3_REIP_REG_26__SCAN_IN), .A2(P3_REIP_REG_25__SCAN_IN), 
        .ZN(n16395) );
  AOI221_X1 U19648 ( .B1(n16396), .B2(n16739), .C1(n16395), .C2(n16739), .A(
        n16737), .ZN(n16460) );
  OAI21_X1 U19649 ( .B1(n16397), .B2(n16710), .A(n16460), .ZN(n16428) );
  INV_X1 U19650 ( .A(n16428), .ZN(n16398) );
  NOR2_X1 U19651 ( .A1(n16710), .A2(n16396), .ZN(n16461) );
  NAND3_X1 U19652 ( .A1(P3_REIP_REG_26__SCAN_IN), .A2(n16461), .A3(
        P3_REIP_REG_25__SCAN_IN), .ZN(n16435) );
  INV_X1 U19653 ( .A(n16435), .ZN(n16449) );
  AND2_X1 U19654 ( .A1(n16449), .A2(n16397), .ZN(n16410) );
  INV_X1 U19655 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n18586) );
  NAND2_X1 U19656 ( .A1(n16410), .A2(n18586), .ZN(n16418) );
  AOI21_X1 U19657 ( .B1(n16398), .B2(n16418), .A(n18583), .ZN(n16408) );
  INV_X1 U19658 ( .A(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n16436) );
  NOR2_X1 U19659 ( .A1(n17670), .A2(n17313), .ZN(n16401) );
  NAND2_X1 U19660 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n16401), .ZN(
        n16400) );
  AOI21_X1 U19661 ( .B1(n16436), .B2(n16400), .A(n16399), .ZN(n17305) );
  OAI21_X1 U19662 ( .B1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n16401), .A(
        n16400), .ZN(n17330) );
  INV_X1 U19663 ( .A(n17330), .ZN(n16445) );
  NAND2_X1 U19664 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17333), .ZN(
        n16402) );
  AOI21_X1 U19665 ( .B1(n10073), .B2(n16402), .A(n16401), .ZN(n17334) );
  INV_X1 U19666 ( .A(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n16470) );
  NAND2_X1 U19667 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n16405), .ZN(
        n16404) );
  INV_X1 U19668 ( .A(n16402), .ZN(n16403) );
  AOI21_X1 U19669 ( .B1(n16470), .B2(n16404), .A(n16403), .ZN(n17344) );
  XOR2_X1 U19670 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .B(n16405), .Z(
        n17359) );
  NOR2_X1 U19671 ( .A1(n16406), .A2(n16667), .ZN(n16472) );
  NOR2_X1 U19672 ( .A1(n17359), .A2(n16472), .ZN(n16471) );
  NOR2_X1 U19673 ( .A1(n16471), .A2(n16667), .ZN(n16464) );
  NOR2_X1 U19674 ( .A1(n16463), .A2(n16667), .ZN(n16453) );
  NOR2_X1 U19675 ( .A1(n17334), .A2(n16453), .ZN(n16452) );
  NOR2_X1 U19676 ( .A1(n16452), .A2(n16667), .ZN(n16444) );
  NOR2_X1 U19677 ( .A1(n16443), .A2(n16667), .ZN(n16432) );
  NOR2_X1 U19678 ( .A1(n17305), .A2(n16432), .ZN(n16431) );
  NOR2_X1 U19679 ( .A1(n16431), .A2(n16667), .ZN(n16425) );
  NOR2_X1 U19680 ( .A1(n16424), .A2(n16667), .ZN(n16416) );
  NAND2_X1 U19681 ( .A1(n9742), .A2(n9882), .ZN(n16741) );
  NOR3_X1 U19682 ( .A1(n16417), .A2(n16416), .A3(n16741), .ZN(n16407) );
  AOI211_X1 U19683 ( .C1(n16409), .C2(n16423), .A(n16408), .B(n16407), .ZN(
        n16412) );
  NAND3_X1 U19684 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n16410), .A3(n18583), 
        .ZN(n16411) );
  NAND3_X1 U19685 ( .A1(n16413), .A2(n16412), .A3(n16411), .ZN(P3_U2640) );
  AOI22_X1 U19686 ( .A1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n16709), .B1(
        P3_REIP_REG_30__SCAN_IN), .B2(n16428), .ZN(n16421) );
  XNOR2_X1 U19687 ( .A(P3_EBX_REG_30__SCAN_IN), .B(n16423), .ZN(n16414) );
  AOI22_X1 U19688 ( .A1(P3_EBX_REG_30__SCAN_IN), .A2(n16750), .B1(n16751), 
        .B2(n16414), .ZN(n16420) );
  AOI21_X1 U19689 ( .B1(n16417), .B2(n16416), .A(n9780), .ZN(n16415) );
  OAI21_X1 U19690 ( .B1(n16417), .B2(n16416), .A(n16415), .ZN(n16419) );
  NAND4_X1 U19691 ( .A1(n16421), .A2(n16420), .A3(n16419), .A4(n16418), .ZN(
        P3_U2641) );
  NOR3_X1 U19692 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n16435), .A3(n16433), 
        .ZN(n16422) );
  AOI21_X1 U19693 ( .B1(P3_EBX_REG_29__SCAN_IN), .B2(n16750), .A(n16422), .ZN(
        n16429) );
  AOI211_X1 U19694 ( .C1(P3_EBX_REG_29__SCAN_IN), .C2(n16439), .A(n16423), .B(
        n16711), .ZN(n16427) );
  INV_X1 U19695 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n18578) );
  AOI211_X1 U19696 ( .C1(n17305), .C2(n16432), .A(n16431), .B(n9780), .ZN(
        n16438) );
  OAI21_X1 U19697 ( .B1(P3_REIP_REG_28__SCAN_IN), .B2(P3_REIP_REG_27__SCAN_IN), 
        .A(n16433), .ZN(n16434) );
  OAI22_X1 U19698 ( .A1(n16436), .A2(n16740), .B1(n16435), .B2(n16434), .ZN(
        n16437) );
  AOI211_X1 U19699 ( .C1(P3_EBX_REG_28__SCAN_IN), .C2(n16750), .A(n16438), .B(
        n16437), .ZN(n16442) );
  OAI211_X1 U19700 ( .C1(n16446), .C2(n16440), .A(n16751), .B(n16439), .ZN(
        n16441) );
  OAI211_X1 U19701 ( .C1(n16460), .C2(n18578), .A(n16442), .B(n16441), .ZN(
        P3_U2643) );
  INV_X1 U19702 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n18575) );
  AOI22_X1 U19703 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n16709), .B1(
        n16750), .B2(P3_EBX_REG_27__SCAN_IN), .ZN(n16451) );
  AOI211_X1 U19704 ( .C1(n16445), .C2(n16444), .A(n16443), .B(n9780), .ZN(
        n16448) );
  AOI211_X1 U19705 ( .C1(P3_EBX_REG_27__SCAN_IN), .C2(n16456), .A(n16446), .B(
        n16711), .ZN(n16447) );
  AOI211_X1 U19706 ( .C1(n16449), .C2(n18575), .A(n16448), .B(n16447), .ZN(
        n16450) );
  OAI211_X1 U19707 ( .C1(n16460), .C2(n18575), .A(n16451), .B(n16450), .ZN(
        P3_U2644) );
  AOI21_X1 U19708 ( .B1(n16461), .B2(P3_REIP_REG_25__SCAN_IN), .A(
        P3_REIP_REG_26__SCAN_IN), .ZN(n16459) );
  AOI211_X1 U19709 ( .C1(n17334), .C2(n16453), .A(n16452), .B(n9780), .ZN(
        n16455) );
  NOR2_X1 U19710 ( .A1(n10073), .A2(n16740), .ZN(n16454) );
  AOI211_X1 U19711 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n16750), .A(n16455), .B(
        n16454), .ZN(n16458) );
  OAI211_X1 U19712 ( .C1(n16462), .C2(n16805), .A(n16751), .B(n16456), .ZN(
        n16457) );
  OAI211_X1 U19713 ( .C1(n16460), .C2(n16459), .A(n16458), .B(n16457), .ZN(
        P3_U2645) );
  INV_X1 U19714 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n20927) );
  AOI22_X1 U19715 ( .A1(n16750), .A2(P3_EBX_REG_25__SCAN_IN), .B1(n16461), 
        .B2(n20927), .ZN(n16469) );
  OAI21_X1 U19716 ( .B1(P3_REIP_REG_24__SCAN_IN), .B2(n16710), .A(n16481), 
        .ZN(n16467) );
  AOI211_X1 U19717 ( .C1(P3_EBX_REG_25__SCAN_IN), .C2(n16477), .A(n16462), .B(
        n16711), .ZN(n16466) );
  AOI211_X1 U19718 ( .C1(n17344), .C2(n16464), .A(n16463), .B(n9780), .ZN(
        n16465) );
  AOI211_X1 U19719 ( .C1(P3_REIP_REG_25__SCAN_IN), .C2(n16467), .A(n16466), 
        .B(n16465), .ZN(n16468) );
  OAI211_X1 U19720 ( .C1(n16470), .C2(n16740), .A(n16469), .B(n16468), .ZN(
        P3_U2646) );
  INV_X1 U19721 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n18571) );
  AOI211_X1 U19722 ( .C1(n17359), .C2(n16472), .A(n16471), .B(n9780), .ZN(
        n16476) );
  INV_X1 U19723 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n17363) );
  NAND2_X1 U19724 ( .A1(n16739), .A2(n18571), .ZN(n16473) );
  OAI22_X1 U19725 ( .A1(n17363), .A2(n16740), .B1(n16474), .B2(n16473), .ZN(
        n16475) );
  AOI211_X1 U19726 ( .C1(P3_EBX_REG_24__SCAN_IN), .C2(n16750), .A(n16476), .B(
        n16475), .ZN(n16480) );
  OAI211_X1 U19727 ( .C1(n16478), .C2(n16758), .A(n16751), .B(n16477), .ZN(
        n16479) );
  OAI211_X1 U19728 ( .C1(n16481), .C2(n18571), .A(n16480), .B(n16479), .ZN(
        P3_U2647) );
  AOI21_X1 U19729 ( .B1(n16739), .B2(n16482), .A(n16737), .ZN(n16513) );
  INV_X1 U19730 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n18567) );
  AOI211_X1 U19731 ( .C1(n17394), .C2(n16484), .A(n16483), .B(n9780), .ZN(
        n16489) );
  OAI211_X1 U19732 ( .C1(n16496), .C2(n16487), .A(n16751), .B(n16485), .ZN(
        n16486) );
  OAI21_X1 U19733 ( .B1(n16487), .B2(n16743), .A(n16486), .ZN(n16488) );
  AOI211_X1 U19734 ( .C1(n16709), .C2(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n16489), .B(n16488), .ZN(n16493) );
  INV_X1 U19735 ( .A(n16502), .ZN(n16491) );
  OAI211_X1 U19736 ( .C1(P3_REIP_REG_22__SCAN_IN), .C2(P3_REIP_REG_21__SCAN_IN), .A(n16491), .B(n16490), .ZN(n16492) );
  OAI211_X1 U19737 ( .C1(n16513), .C2(n18567), .A(n16493), .B(n16492), .ZN(
        P3_U2649) );
  INV_X1 U19738 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n18565) );
  AOI211_X1 U19739 ( .C1(n17412), .C2(n16495), .A(n16494), .B(n9780), .ZN(
        n16500) );
  AOI211_X1 U19740 ( .C1(P3_EBX_REG_21__SCAN_IN), .C2(n16504), .A(n16496), .B(
        n16711), .ZN(n16499) );
  OAI22_X1 U19741 ( .A1(n17409), .A2(n16740), .B1(n16743), .B2(n16497), .ZN(
        n16498) );
  NOR3_X1 U19742 ( .A1(n16500), .A2(n16499), .A3(n16498), .ZN(n16501) );
  OAI221_X1 U19743 ( .B1(P3_REIP_REG_21__SCAN_IN), .B2(n16502), .C1(n18565), 
        .C2(n16513), .A(n16501), .ZN(P3_U2650) );
  INV_X1 U19744 ( .A(n16520), .ZN(n16503) );
  AOI21_X1 U19745 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(n16503), .A(n16711), .ZN(
        n16505) );
  AOI22_X1 U19746 ( .A1(n16750), .A2(P3_EBX_REG_20__SCAN_IN), .B1(n16505), 
        .B2(n16504), .ZN(n16512) );
  AOI211_X1 U19747 ( .C1(n17425), .C2(n16507), .A(n16506), .B(n9780), .ZN(
        n16510) );
  NOR3_X1 U19748 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(n16508), .A3(n16566), 
        .ZN(n16509) );
  AOI211_X1 U19749 ( .C1(n16709), .C2(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n16510), .B(n16509), .ZN(n16511) );
  OAI211_X1 U19750 ( .C1(n18564), .C2(n16513), .A(n16512), .B(n16511), .ZN(
        P3_U2651) );
  INV_X1 U19751 ( .A(n16519), .ZN(n16514) );
  INV_X1 U19752 ( .A(n16737), .ZN(n16753) );
  NAND2_X1 U19753 ( .A1(n16710), .A2(n16753), .ZN(n16752) );
  OAI21_X1 U19754 ( .B1(n16572), .B2(n16710), .A(n16753), .ZN(n16546) );
  AOI21_X1 U19755 ( .B1(n16514), .B2(n16752), .A(n16546), .ZN(n16545) );
  INV_X1 U19756 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n18561) );
  INV_X1 U19757 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n17445) );
  NOR2_X1 U19758 ( .A1(n17445), .A2(n16536), .ZN(n16515) );
  OAI21_X1 U19759 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n16515), .A(
        n17386), .ZN(n17433) );
  INV_X1 U19760 ( .A(n16515), .ZN(n16525) );
  OAI21_X1 U19761 ( .B1(n16549), .B2(n16525), .A(n9742), .ZN(n16517) );
  OAI21_X1 U19762 ( .B1(n17433), .B2(n16517), .A(n9882), .ZN(n16516) );
  AOI21_X1 U19763 ( .B1(n17433), .B2(n16517), .A(n16516), .ZN(n16518) );
  AOI211_X1 U19764 ( .C1(n16750), .C2(P3_EBX_REG_19__SCAN_IN), .A(n17979), .B(
        n16518), .ZN(n16524) );
  INV_X1 U19765 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n18559) );
  NAND2_X1 U19766 ( .A1(n16519), .A2(n16548), .ZN(n16534) );
  AOI221_X1 U19767 ( .B1(P3_REIP_REG_19__SCAN_IN), .B2(P3_REIP_REG_18__SCAN_IN), .C1(n18561), .C2(n18559), .A(n16534), .ZN(n16522) );
  AOI211_X1 U19768 ( .C1(P3_EBX_REG_19__SCAN_IN), .C2(n16529), .A(n16520), .B(
        n16711), .ZN(n16521) );
  AOI211_X1 U19769 ( .C1(n16709), .C2(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n16522), .B(n16521), .ZN(n16523) );
  OAI211_X1 U19770 ( .C1(n16545), .C2(n18561), .A(n16524), .B(n16523), .ZN(
        P3_U2652) );
  AOI22_X1 U19771 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n16709), .B1(
        n16750), .B2(P3_EBX_REG_18__SCAN_IN), .ZN(n16532) );
  INV_X1 U19772 ( .A(n16526), .ZN(n16528) );
  INV_X1 U19773 ( .A(n16536), .ZN(n17429) );
  OAI21_X1 U19774 ( .B1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n17429), .A(
        n16525), .ZN(n17442) );
  INV_X1 U19775 ( .A(n17442), .ZN(n16527) );
  OAI221_X1 U19776 ( .B1(n16528), .B2(n16527), .C1(n16526), .C2(n17442), .A(
        n9882), .ZN(n16531) );
  OAI211_X1 U19777 ( .C1(n16540), .C2(n16887), .A(n16751), .B(n16529), .ZN(
        n16530) );
  AND4_X1 U19778 ( .A1(n16532), .A2(n17993), .A3(n16531), .A4(n16530), .ZN(
        n16533) );
  OAI221_X1 U19779 ( .B1(P3_REIP_REG_18__SCAN_IN), .B2(n16534), .C1(n18559), 
        .C2(n16545), .A(n16533), .ZN(P3_U2653) );
  NOR3_X1 U19780 ( .A1(P3_REIP_REG_17__SCAN_IN), .A2(n16547), .A3(n16566), 
        .ZN(n16535) );
  AOI211_X1 U19781 ( .C1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .C2(n16709), .A(
        n17979), .B(n16535), .ZN(n16544) );
  OAI21_X1 U19782 ( .B1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n16537), .A(
        n16536), .ZN(n17454) );
  INV_X1 U19783 ( .A(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n16559) );
  NAND2_X1 U19784 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n17468), .ZN(
        n16561) );
  AOI21_X1 U19785 ( .B1(n16559), .B2(n16561), .A(n16537), .ZN(n17469) );
  OAI21_X1 U19786 ( .B1(n17469), .B2(n16549), .A(n9742), .ZN(n16539) );
  OAI21_X1 U19787 ( .B1(n17454), .B2(n16539), .A(n9882), .ZN(n16538) );
  AOI21_X1 U19788 ( .B1(n17454), .B2(n16539), .A(n16538), .ZN(n16542) );
  AOI211_X1 U19789 ( .C1(P3_EBX_REG_17__SCAN_IN), .C2(n16556), .A(n16540), .B(
        n16711), .ZN(n16541) );
  AOI211_X1 U19790 ( .C1(P3_EBX_REG_17__SCAN_IN), .C2(n16750), .A(n16542), .B(
        n16541), .ZN(n16543) );
  OAI211_X1 U19791 ( .C1(n16545), .C2(n18558), .A(n16544), .B(n16543), .ZN(
        P3_U2654) );
  INV_X1 U19792 ( .A(n16546), .ZN(n16575) );
  INV_X1 U19793 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n18555) );
  OAI211_X1 U19794 ( .C1(P3_REIP_REG_16__SCAN_IN), .C2(P3_REIP_REG_15__SCAN_IN), .A(n16548), .B(n16547), .ZN(n16554) );
  INV_X1 U19795 ( .A(n17469), .ZN(n16552) );
  NAND2_X1 U19796 ( .A1(n9742), .A2(n16549), .ZN(n16551) );
  NAND2_X1 U19797 ( .A1(n16552), .A2(n16551), .ZN(n16550) );
  OAI211_X1 U19798 ( .C1(n16552), .C2(n16551), .A(n9882), .B(n16550), .ZN(
        n16553) );
  OAI211_X1 U19799 ( .C1(n16575), .C2(n18555), .A(n16554), .B(n16553), .ZN(
        n16555) );
  AOI211_X1 U19800 ( .C1(n16750), .C2(P3_EBX_REG_16__SCAN_IN), .A(n17979), .B(
        n16555), .ZN(n16558) );
  OAI211_X1 U19801 ( .C1(n16560), .C2(n16914), .A(n16751), .B(n16556), .ZN(
        n16557) );
  OAI211_X1 U19802 ( .C1(n16740), .C2(n16559), .A(n16558), .B(n16557), .ZN(
        P3_U2655) );
  INV_X1 U19803 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n16570) );
  AOI211_X1 U19804 ( .C1(P3_EBX_REG_15__SCAN_IN), .C2(n16578), .A(n16560), .B(
        n16711), .ZN(n16568) );
  INV_X1 U19805 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n18553) );
  OAI21_X1 U19806 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n17468), .A(
        n16561), .ZN(n17484) );
  OR2_X1 U19807 ( .A1(n16562), .A2(n16667), .ZN(n16564) );
  AOI21_X1 U19808 ( .B1(n17484), .B2(n16564), .A(n9780), .ZN(n16563) );
  OAI21_X1 U19809 ( .B1(n17484), .B2(n16564), .A(n16563), .ZN(n16565) );
  OAI221_X1 U19810 ( .B1(P3_REIP_REG_15__SCAN_IN), .B2(n16566), .C1(n18553), 
        .C2(n16575), .A(n16565), .ZN(n16567) );
  AOI211_X1 U19811 ( .C1(n16709), .C2(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A(
        n16568), .B(n16567), .ZN(n16569) );
  OAI211_X1 U19812 ( .C1(n16743), .C2(n16570), .A(n16569), .B(n17993), .ZN(
        P3_U2656) );
  NOR2_X1 U19813 ( .A1(n17670), .A2(n17506), .ZN(n17508) );
  INV_X1 U19814 ( .A(n17508), .ZN(n16582) );
  OR2_X1 U19815 ( .A1(n17509), .A2(n16582), .ZN(n16583) );
  AOI21_X1 U19816 ( .B1(n17498), .B2(n16583), .A(n17468), .ZN(n17500) );
  OAI21_X1 U19817 ( .B1(n17509), .B2(n16597), .A(n9742), .ZN(n16571) );
  XNOR2_X1 U19818 ( .A(n17500), .B(n16571), .ZN(n16577) );
  NOR3_X1 U19819 ( .A1(n16710), .A2(n16572), .A3(n16586), .ZN(n16573) );
  AOI22_X1 U19820 ( .A1(n16750), .A2(P3_EBX_REG_14__SCAN_IN), .B1(
        P3_REIP_REG_13__SCAN_IN), .B2(n16573), .ZN(n16574) );
  OAI211_X1 U19821 ( .C1(n18552), .C2(n16575), .A(n16574), .B(n17993), .ZN(
        n16576) );
  AOI21_X1 U19822 ( .B1(n16577), .B2(n9882), .A(n16576), .ZN(n16581) );
  OAI211_X1 U19823 ( .C1(n16590), .C2(n16579), .A(n16751), .B(n16578), .ZN(
        n16580) );
  OAI211_X1 U19824 ( .C1(n16740), .C2(n17498), .A(n16581), .B(n16580), .ZN(
        P3_U2657) );
  AOI22_X1 U19825 ( .A1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n16709), .B1(
        n16750), .B2(P3_EBX_REG_13__SCAN_IN), .ZN(n16595) );
  INV_X1 U19826 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n16605) );
  NOR2_X1 U19827 ( .A1(n16605), .A2(n16582), .ZN(n16584) );
  OAI21_X1 U19828 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n16584), .A(
        n16583), .ZN(n17511) );
  INV_X1 U19829 ( .A(n16584), .ZN(n16596) );
  OAI21_X1 U19830 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16596), .A(
        n9742), .ZN(n16585) );
  XOR2_X1 U19831 ( .A(n17511), .B(n16585), .Z(n16588) );
  NOR2_X1 U19832 ( .A1(n16710), .A2(n16586), .ZN(n16587) );
  AOI22_X1 U19833 ( .A1(n9882), .A2(n16588), .B1(n16587), .B2(n18549), .ZN(
        n16594) );
  INV_X1 U19834 ( .A(n16600), .ZN(n16589) );
  AOI21_X1 U19835 ( .B1(n16739), .B2(n16589), .A(n16737), .ZN(n16609) );
  OAI21_X1 U19836 ( .B1(P3_REIP_REG_12__SCAN_IN), .B2(n16710), .A(n16609), 
        .ZN(n16592) );
  AOI211_X1 U19837 ( .C1(P3_EBX_REG_13__SCAN_IN), .C2(n16602), .A(n16590), .B(
        n16711), .ZN(n16591) );
  AOI211_X1 U19838 ( .C1(P3_REIP_REG_13__SCAN_IN), .C2(n16592), .A(n17979), 
        .B(n16591), .ZN(n16593) );
  NAND3_X1 U19839 ( .A1(n16595), .A2(n16594), .A3(n16593), .ZN(P3_U2658) );
  INV_X1 U19840 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n18547) );
  OAI21_X1 U19841 ( .B1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n17508), .A(
        n16596), .ZN(n17522) );
  NAND2_X1 U19842 ( .A1(n9742), .A2(n16597), .ZN(n16598) );
  XOR2_X1 U19843 ( .A(n17522), .B(n16598), .Z(n16601) );
  NOR2_X1 U19844 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n16710), .ZN(n16599) );
  AOI22_X1 U19845 ( .A1(n9882), .A2(n16601), .B1(n16600), .B2(n16599), .ZN(
        n16604) );
  OAI211_X1 U19846 ( .C1(n16611), .C2(n16938), .A(n16751), .B(n16602), .ZN(
        n16603) );
  OAI211_X1 U19847 ( .C1(n16740), .C2(n16605), .A(n16604), .B(n16603), .ZN(
        n16606) );
  AOI211_X1 U19848 ( .C1(n16750), .C2(P3_EBX_REG_12__SCAN_IN), .A(n17979), .B(
        n16606), .ZN(n16607) );
  OAI21_X1 U19849 ( .B1(n18547), .B2(n16609), .A(n16607), .ZN(P3_U2659) );
  OR2_X1 U19850 ( .A1(n17544), .A2(n16666), .ZN(n16619) );
  AOI21_X1 U19851 ( .B1(n17534), .B2(n16619), .A(n17508), .ZN(n17537) );
  NOR2_X1 U19852 ( .A1(n16608), .A2(n16667), .ZN(n16621) );
  XNOR2_X1 U19853 ( .A(n17537), .B(n16621), .ZN(n16616) );
  AOI21_X1 U19854 ( .B1(n16681), .B2(P3_EBX_REG_11__SCAN_IN), .A(n17979), .ZN(
        n16615) );
  NAND3_X1 U19855 ( .A1(n16739), .A2(P3_REIP_REG_8__SCAN_IN), .A3(n16642), 
        .ZN(n16641) );
  AOI221_X1 U19856 ( .B1(n16610), .B2(n18545), .C1(n16641), .C2(n18545), .A(
        n16609), .ZN(n16613) );
  AOI211_X1 U19857 ( .C1(P3_EBX_REG_11__SCAN_IN), .C2(n16628), .A(n16611), .B(
        n16711), .ZN(n16612) );
  AOI211_X1 U19858 ( .C1(n16709), .C2(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n16613), .B(n16612), .ZN(n16614) );
  OAI211_X1 U19859 ( .C1(n9780), .C2(n16616), .A(n16615), .B(n16614), .ZN(
        P3_U2660) );
  INV_X1 U19860 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n18543) );
  NOR2_X1 U19861 ( .A1(n18543), .A2(n16641), .ZN(n16627) );
  INV_X1 U19862 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n18544) );
  AOI21_X1 U19863 ( .B1(n16739), .B2(n16617), .A(n16737), .ZN(n16647) );
  OAI21_X1 U19864 ( .B1(P3_REIP_REG_9__SCAN_IN), .B2(n16641), .A(n16647), .ZN(
        n16626) );
  INV_X1 U19865 ( .A(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n16624) );
  NAND3_X1 U19866 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n16618) );
  NOR2_X1 U19867 ( .A1(n16618), .A2(n16666), .ZN(n16620) );
  OAI21_X1 U19868 ( .B1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n16620), .A(
        n16619), .ZN(n17546) );
  INV_X1 U19869 ( .A(n17546), .ZN(n16622) );
  INV_X1 U19870 ( .A(n16620), .ZN(n16632) );
  OAI21_X1 U19871 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16632), .A(
        n9742), .ZN(n16634) );
  OAI221_X1 U19872 ( .B1(n16622), .B2(n16621), .C1(n17546), .C2(n16634), .A(
        n9882), .ZN(n16623) );
  OAI211_X1 U19873 ( .C1(n16624), .C2(n16740), .A(n17993), .B(n16623), .ZN(
        n16625) );
  AOI221_X1 U19874 ( .B1(n16627), .B2(n18544), .C1(n16626), .C2(
        P3_REIP_REG_10__SCAN_IN), .A(n16625), .ZN(n16630) );
  OAI211_X1 U19875 ( .C1(n16631), .C2(n20809), .A(n16751), .B(n16628), .ZN(
        n16629) );
  OAI211_X1 U19876 ( .C1(n20809), .C2(n16743), .A(n16630), .B(n16629), .ZN(
        P3_U2661) );
  AOI211_X1 U19877 ( .C1(P3_EBX_REG_9__SCAN_IN), .C2(n16649), .A(n16631), .B(
        n16711), .ZN(n16639) );
  INV_X1 U19878 ( .A(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n17581) );
  INV_X1 U19879 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n17590) );
  NOR2_X1 U19880 ( .A1(n17577), .A2(n17590), .ZN(n17579) );
  NAND2_X1 U19881 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17579), .ZN(
        n16654) );
  NOR2_X1 U19882 ( .A1(n17581), .A2(n16654), .ZN(n16643) );
  OAI21_X1 U19883 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n16643), .A(
        n16632), .ZN(n17568) );
  NAND2_X1 U19884 ( .A1(n9882), .A2(n16667), .ZN(n16728) );
  INV_X1 U19885 ( .A(n17568), .ZN(n16635) );
  INV_X1 U19886 ( .A(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n17545) );
  NAND2_X1 U19887 ( .A1(n16643), .A2(n17545), .ZN(n16633) );
  OAI22_X1 U19888 ( .A1(n16635), .A2(n16634), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16633), .ZN(n16636) );
  AOI22_X1 U19889 ( .A1(n16750), .A2(P3_EBX_REG_9__SCAN_IN), .B1(n9882), .B2(
        n16636), .ZN(n16637) );
  OAI211_X1 U19890 ( .C1(n17568), .C2(n16728), .A(n16637), .B(n17993), .ZN(
        n16638) );
  AOI211_X1 U19891 ( .C1(n16709), .C2(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A(
        n16639), .B(n16638), .ZN(n16640) );
  OAI221_X1 U19892 ( .B1(P3_REIP_REG_9__SCAN_IN), .B2(n16641), .C1(n18543), 
        .C2(n16647), .A(n16640), .ZN(P3_U2662) );
  AOI21_X1 U19893 ( .B1(n16739), .B2(n16642), .A(P3_REIP_REG_8__SCAN_IN), .ZN(
        n16646) );
  AOI21_X1 U19894 ( .B1(n17581), .B2(n16654), .A(n16643), .ZN(n17583) );
  OAI21_X1 U19895 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16666), .A(
        n9742), .ZN(n16665) );
  OAI21_X1 U19896 ( .B1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n16667), .A(
        n16665), .ZN(n16644) );
  XNOR2_X1 U19897 ( .A(n17583), .B(n16644), .ZN(n16645) );
  OAI22_X1 U19898 ( .A1(n16647), .A2(n16646), .B1(n9780), .B2(n16645), .ZN(
        n16648) );
  AOI211_X1 U19899 ( .C1(n16750), .C2(P3_EBX_REG_8__SCAN_IN), .A(n17979), .B(
        n16648), .ZN(n16652) );
  OAI211_X1 U19900 ( .C1(n16658), .C2(n16650), .A(n16751), .B(n16649), .ZN(
        n16651) );
  OAI211_X1 U19901 ( .C1(n16740), .C2(n17581), .A(n16652), .B(n16651), .ZN(
        P3_U2663) );
  INV_X1 U19902 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n18537) );
  OAI21_X1 U19903 ( .B1(n16672), .B2(n16710), .A(n16753), .ZN(n16682) );
  AOI21_X1 U19904 ( .B1(n16739), .B2(n18537), .A(n16682), .ZN(n16664) );
  AOI22_X1 U19905 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n16709), .B1(
        n16750), .B2(P3_EBX_REG_7__SCAN_IN), .ZN(n16663) );
  NOR3_X1 U19906 ( .A1(P3_REIP_REG_7__SCAN_IN), .A2(n16710), .A3(n16653), .ZN(
        n16661) );
  INV_X1 U19907 ( .A(n16666), .ZN(n16655) );
  OAI21_X1 U19908 ( .B1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n16655), .A(
        n16654), .ZN(n17602) );
  INV_X1 U19909 ( .A(n17602), .ZN(n16657) );
  INV_X1 U19910 ( .A(n16665), .ZN(n16656) );
  AOI221_X1 U19911 ( .B1(n16657), .B2(n16656), .C1(n17602), .C2(n16665), .A(
        n9780), .ZN(n16660) );
  AOI211_X1 U19912 ( .C1(P3_EBX_REG_7__SCAN_IN), .C2(n16673), .A(n16658), .B(
        n16711), .ZN(n16659) );
  NOR4_X1 U19913 ( .A1(n17995), .A2(n16661), .A3(n16660), .A4(n16659), .ZN(
        n16662) );
  OAI211_X1 U19914 ( .C1(n16664), .C2(n18539), .A(n16663), .B(n16662), .ZN(
        P3_U2664) );
  AOI22_X1 U19915 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n16709), .B1(
        n16750), .B2(P3_EBX_REG_6__SCAN_IN), .ZN(n16678) );
  NOR2_X1 U19916 ( .A1(n9780), .A2(n16665), .ZN(n16670) );
  OAI21_X1 U19917 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n16680), .A(
        n16666), .ZN(n17609) );
  INV_X1 U19918 ( .A(n16680), .ZN(n16668) );
  INV_X1 U19919 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n16742) );
  OAI21_X1 U19920 ( .B1(n16667), .B2(n16742), .A(n9882), .ZN(n16744) );
  AOI211_X1 U19921 ( .C1(n9742), .C2(n16668), .A(n17609), .B(n16744), .ZN(
        n16669) );
  AOI211_X1 U19922 ( .C1(n16670), .C2(n17609), .A(n17979), .B(n16669), .ZN(
        n16677) );
  NOR2_X1 U19923 ( .A1(P3_REIP_REG_6__SCAN_IN), .A2(n16710), .ZN(n16671) );
  AOI22_X1 U19924 ( .A1(P3_REIP_REG_6__SCAN_IN), .A2(n16682), .B1(n16672), 
        .B2(n16671), .ZN(n16676) );
  OAI211_X1 U19925 ( .C1(n16685), .C2(n16674), .A(n16751), .B(n16673), .ZN(
        n16675) );
  NAND4_X1 U19926 ( .A1(n16678), .A2(n16677), .A3(n16676), .A4(n16675), .ZN(
        P3_U2665) );
  INV_X1 U19927 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n17620) );
  NAND2_X1 U19928 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n16679), .ZN(
        n16691) );
  AOI21_X1 U19929 ( .B1(n17620), .B2(n16691), .A(n16680), .ZN(n17622) );
  OAI21_X1 U19930 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16691), .A(
        n9742), .ZN(n16692) );
  XOR2_X1 U19931 ( .A(n17622), .B(n16692), .Z(n16690) );
  AOI21_X1 U19932 ( .B1(n16681), .B2(P3_EBX_REG_5__SCAN_IN), .A(n17979), .ZN(
        n16689) );
  INV_X1 U19933 ( .A(n16682), .ZN(n16683) );
  AOI221_X1 U19934 ( .B1(n16710), .B2(n18535), .C1(n16684), .C2(n18535), .A(
        n16683), .ZN(n16687) );
  AOI211_X1 U19935 ( .C1(P3_EBX_REG_5__SCAN_IN), .C2(n16700), .A(n16685), .B(
        n16711), .ZN(n16686) );
  AOI211_X1 U19936 ( .C1(n16709), .C2(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .A(
        n16687), .B(n16686), .ZN(n16688) );
  OAI211_X1 U19937 ( .C1(n9780), .C2(n16690), .A(n16689), .B(n16688), .ZN(
        P3_U2666) );
  AND2_X1 U19938 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17631), .ZN(
        n16707) );
  OAI21_X1 U19939 ( .B1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n16707), .A(
        n16691), .ZN(n17634) );
  INV_X1 U19940 ( .A(n17634), .ZN(n16693) );
  NAND2_X1 U19941 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n16742), .ZN(
        n16723) );
  INV_X1 U19942 ( .A(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n16698) );
  NAND2_X1 U19943 ( .A1(n17631), .A2(n16698), .ZN(n17638) );
  OAI22_X1 U19944 ( .A1(n16693), .A2(n16692), .B1(n16723), .B2(n17638), .ZN(
        n16697) );
  NAND2_X1 U19945 ( .A1(n16694), .A2(n18669), .ZN(n16720) );
  AOI21_X1 U19946 ( .B1(n9787), .B2(n16695), .A(n16720), .ZN(n16696) );
  AOI211_X1 U19947 ( .C1(n9882), .C2(n16697), .A(n17979), .B(n16696), .ZN(
        n16706) );
  OAI21_X1 U19948 ( .B1(n16699), .B2(n16710), .A(n16753), .ZN(n16716) );
  OAI22_X1 U19949 ( .A1(n16698), .A2(n16740), .B1(n16743), .B2(n17020), .ZN(
        n16704) );
  NAND2_X1 U19950 ( .A1(n16739), .A2(n16699), .ZN(n16702) );
  OAI211_X1 U19951 ( .C1(n16712), .C2(n17020), .A(n16751), .B(n16700), .ZN(
        n16701) );
  OAI21_X1 U19952 ( .B1(P3_REIP_REG_4__SCAN_IN), .B2(n16702), .A(n16701), .ZN(
        n16703) );
  AOI211_X1 U19953 ( .C1(P3_REIP_REG_4__SCAN_IN), .C2(n16716), .A(n16704), .B(
        n16703), .ZN(n16705) );
  OAI211_X1 U19954 ( .C1(n17634), .C2(n16728), .A(n16706), .B(n16705), .ZN(
        P3_U2667) );
  NAND2_X1 U19955 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n16721) );
  AOI21_X1 U19956 ( .B1(n17645), .B2(n16721), .A(n16707), .ZN(n17649) );
  OAI21_X1 U19957 ( .B1(n17662), .B2(n16723), .A(n9742), .ZN(n16708) );
  XOR2_X1 U19958 ( .A(n17649), .B(n16708), .Z(n16719) );
  AOI22_X1 U19959 ( .A1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n16709), .B1(
        n16750), .B2(P3_EBX_REG_3__SCAN_IN), .ZN(n16718) );
  OAI21_X1 U19960 ( .B1(n16710), .B2(n16732), .A(n18532), .ZN(n16715) );
  AOI211_X1 U19961 ( .C1(P3_EBX_REG_3__SCAN_IN), .C2(n16725), .A(n16712), .B(
        n16711), .ZN(n16714) );
  NAND2_X1 U19962 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n18460) );
  NOR2_X1 U19963 ( .A1(n18630), .A2(n18460), .ZN(n18457) );
  OAI21_X1 U19964 ( .B1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n18457), .A(
        n9787), .ZN(n18601) );
  NOR2_X1 U19965 ( .A1(n16720), .A2(n18601), .ZN(n16713) );
  AOI211_X1 U19966 ( .C1(n16716), .C2(n16715), .A(n16714), .B(n16713), .ZN(
        n16717) );
  OAI211_X1 U19967 ( .C1(n9780), .C2(n16719), .A(n16718), .B(n16717), .ZN(
        P3_U2668) );
  NAND2_X1 U19968 ( .A1(n18617), .A2(n18478), .ZN(n18455) );
  INV_X1 U19969 ( .A(n18455), .ZN(n18461) );
  NOR2_X1 U19970 ( .A1(n18461), .A2(n18457), .ZN(n18613) );
  INV_X1 U19971 ( .A(n16720), .ZN(n18671) );
  AOI22_X1 U19972 ( .A1(P3_REIP_REG_2__SCAN_IN), .A2(n16737), .B1(n18613), 
        .B2(n18671), .ZN(n16735) );
  OAI21_X1 U19973 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n16721), .ZN(n17658) );
  INV_X1 U19974 ( .A(n17658), .ZN(n16724) );
  NOR2_X1 U19975 ( .A1(n17662), .A2(n16723), .ZN(n16722) );
  AOI211_X1 U19976 ( .C1(n16724), .C2(n16723), .A(n16722), .B(n16741), .ZN(
        n16731) );
  OAI22_X1 U19977 ( .A1(n17662), .A2(n16740), .B1(n16743), .B2(n16726), .ZN(
        n16730) );
  OAI211_X1 U19978 ( .C1(n16738), .C2(n16726), .A(n16751), .B(n16725), .ZN(
        n16727) );
  OAI21_X1 U19979 ( .B1(n16728), .B2(n17658), .A(n16727), .ZN(n16729) );
  NOR3_X1 U19980 ( .A1(n16731), .A2(n16730), .A3(n16729), .ZN(n16734) );
  OAI211_X1 U19981 ( .C1(P3_REIP_REG_2__SCAN_IN), .C2(P3_REIP_REG_1__SCAN_IN), 
        .A(n16739), .B(n16732), .ZN(n16733) );
  NAND3_X1 U19982 ( .A1(n16735), .A2(n16734), .A3(n16733), .ZN(P3_U2669) );
  AND2_X1 U19983 ( .A1(n18478), .A2(n16736), .ZN(n18621) );
  AOI22_X1 U19984 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n16737), .B1(n18621), 
        .B2(n18671), .ZN(n16749) );
  AOI21_X1 U19985 ( .B1(P3_EBX_REG_1__SCAN_IN), .B2(P3_EBX_REG_0__SCAN_IN), 
        .A(n16738), .ZN(n17032) );
  INV_X1 U19986 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n18529) );
  AOI22_X1 U19987 ( .A1(n16751), .A2(n17032), .B1(n16739), .B2(n18529), .ZN(
        n16748) );
  OAI21_X1 U19988 ( .B1(n16742), .B2(n16741), .A(n16740), .ZN(n16746) );
  INV_X1 U19989 ( .A(P3_EBX_REG_1__SCAN_IN), .ZN(n17035) );
  OAI22_X1 U19990 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n16744), .B1(
        n17035), .B2(n16743), .ZN(n16745) );
  AOI21_X1 U19991 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n16746), .A(
        n16745), .ZN(n16747) );
  NAND3_X1 U19992 ( .A1(n16749), .A2(n16748), .A3(n16747), .ZN(P3_U2670) );
  NOR2_X1 U19993 ( .A1(n16751), .A2(n16750), .ZN(n16756) );
  INV_X1 U19994 ( .A(P3_EBX_REG_0__SCAN_IN), .ZN(n17038) );
  AOI22_X1 U19995 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(n16752), .B1(n18671), 
        .B2(n18630), .ZN(n16755) );
  NAND3_X1 U19996 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n18602), .A3(
        n16753), .ZN(n16754) );
  OAI211_X1 U19997 ( .C1(n16756), .C2(n17038), .A(n16755), .B(n16754), .ZN(
        P3_U2671) );
  INV_X1 U19998 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n16764) );
  INV_X1 U19999 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n16759) );
  NAND4_X1 U20000 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(P3_EBX_REG_21__SCAN_IN), 
        .A3(n16835), .A4(n16796), .ZN(n16757) );
  NOR4_X1 U20001 ( .A1(n16759), .A2(n16758), .A3(n16812), .A4(n16757), .ZN(
        n16760) );
  NAND3_X1 U20002 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(P3_EBX_REG_25__SCAN_IN), 
        .A3(n16760), .ZN(n16763) );
  NAND2_X1 U20003 ( .A1(n17039), .A2(P3_EBX_REG_31__SCAN_IN), .ZN(n16762) );
  NAND2_X1 U20004 ( .A1(n16791), .A2(n17047), .ZN(n16761) );
  OAI22_X1 U20005 ( .A1(n16791), .A2(n16762), .B1(P3_EBX_REG_31__SCAN_IN), 
        .B2(n16761), .ZN(P3_U2672) );
  NAND2_X1 U20006 ( .A1(n16764), .A2(n16763), .ZN(n16765) );
  NAND2_X1 U20007 ( .A1(n16765), .A2(n17039), .ZN(n16790) );
  AOI22_X1 U20008 ( .A1(n16993), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n16975), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n16776) );
  AOI22_X1 U20009 ( .A1(n15162), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n9729), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n16775) );
  AOI22_X1 U20010 ( .A1(n15318), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n16974), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n16766) );
  OAI21_X1 U20011 ( .B1(n16767), .B2(n17009), .A(n16766), .ZN(n16773) );
  AOI22_X1 U20012 ( .A1(n16954), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n16777), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n16771) );
  AOI22_X1 U20013 ( .A1(n15149), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n9726), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n16770) );
  AOI22_X1 U20014 ( .A1(n16968), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n16986), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n16769) );
  AOI22_X1 U20015 ( .A1(n16969), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n16991), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n16768) );
  NAND4_X1 U20016 ( .A1(n16771), .A2(n16770), .A3(n16769), .A4(n16768), .ZN(
        n16772) );
  AOI211_X1 U20017 ( .C1(n11754), .C2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A(
        n16773), .B(n16772), .ZN(n16774) );
  NAND3_X1 U20018 ( .A1(n16776), .A2(n16775), .A3(n16774), .ZN(n16789) );
  AOI22_X1 U20019 ( .A1(n16975), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n16991), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n16781) );
  AOI22_X1 U20020 ( .A1(n15162), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11754), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n16780) );
  AOI22_X1 U20021 ( .A1(n16969), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n11806), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n16779) );
  AOI22_X1 U20022 ( .A1(n16993), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n16777), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n16778) );
  NAND4_X1 U20023 ( .A1(n16781), .A2(n16780), .A3(n16779), .A4(n16778), .ZN(
        n16787) );
  AOI22_X1 U20024 ( .A1(n16968), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n15279), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n16785) );
  AOI22_X1 U20025 ( .A1(n9729), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n16987), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n16784) );
  AOI22_X1 U20026 ( .A1(n9726), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n16974), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n16783) );
  AOI22_X1 U20027 ( .A1(n15149), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n16986), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n16782) );
  NAND4_X1 U20028 ( .A1(n16785), .A2(n16784), .A3(n16783), .A4(n16782), .ZN(
        n16786) );
  NOR2_X1 U20029 ( .A1(n16787), .A2(n16786), .ZN(n16794) );
  NOR3_X1 U20030 ( .A1(n16794), .A2(n16792), .A3(n17065), .ZN(n16788) );
  XNOR2_X1 U20031 ( .A(n16789), .B(n16788), .ZN(n17055) );
  OAI22_X1 U20032 ( .A1(n16791), .A2(n16790), .B1(n17055), .B2(n17039), .ZN(
        P3_U2673) );
  NOR2_X1 U20033 ( .A1(n16792), .A2(n17065), .ZN(n16793) );
  XOR2_X1 U20034 ( .A(n16794), .B(n16793), .Z(n17059) );
  NOR2_X1 U20035 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n16801), .ZN(n16795) );
  AOI22_X1 U20036 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n16797), .B1(n16796), 
        .B2(n16795), .ZN(n16798) );
  OAI21_X1 U20037 ( .B1(n17039), .B2(n17059), .A(n16798), .ZN(P3_U2674) );
  OAI211_X1 U20038 ( .C1(n17067), .C2(n17066), .A(n17024), .B(n17065), .ZN(
        n16799) );
  OAI221_X1 U20039 ( .B1(P3_EBX_REG_27__SCAN_IN), .B2(n16801), .C1(n16800), 
        .C2(n16804), .A(n16799), .ZN(P3_U2676) );
  AOI21_X1 U20040 ( .B1(n16802), .B2(n16807), .A(n17067), .ZN(n17072) );
  NAND2_X1 U20041 ( .A1(n17024), .A2(n17072), .ZN(n16803) );
  OAI221_X1 U20042 ( .B1(P3_EBX_REG_26__SCAN_IN), .B2(n16806), .C1(n16805), 
        .C2(n16804), .A(n16803), .ZN(P3_U2677) );
  INV_X1 U20043 ( .A(n16806), .ZN(n16811) );
  AOI21_X1 U20044 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n17039), .A(n16815), .ZN(
        n16810) );
  OAI21_X1 U20045 ( .B1(n16809), .B2(n16808), .A(n16807), .ZN(n17081) );
  OAI22_X1 U20046 ( .A1(n16811), .A2(n16810), .B1(n17039), .B2(n17081), .ZN(
        P3_U2678) );
  NOR2_X1 U20047 ( .A1(n16812), .A2(n16816), .ZN(n16821) );
  AOI21_X1 U20048 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n17039), .A(n16821), .ZN(
        n16814) );
  XNOR2_X1 U20049 ( .A(n16813), .B(n16817), .ZN(n17086) );
  OAI22_X1 U20050 ( .A1(n16815), .A2(n16814), .B1(n17039), .B2(n17086), .ZN(
        P3_U2679) );
  INV_X1 U20051 ( .A(n16816), .ZN(n16834) );
  AOI21_X1 U20052 ( .B1(P3_EBX_REG_23__SCAN_IN), .B2(n17039), .A(n16834), .ZN(
        n16820) );
  OAI21_X1 U20053 ( .B1(n16819), .B2(n16818), .A(n16817), .ZN(n17091) );
  OAI22_X1 U20054 ( .A1(n16821), .A2(n16820), .B1(n17039), .B2(n17091), .ZN(
        P3_U2680) );
  AOI21_X1 U20055 ( .B1(P3_EBX_REG_22__SCAN_IN), .B2(n17039), .A(n16822), .ZN(
        n16833) );
  AOI22_X1 U20056 ( .A1(n15149), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n16987), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n16826) );
  AOI22_X1 U20057 ( .A1(n15162), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11754), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n16825) );
  AOI22_X1 U20058 ( .A1(n16993), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n16969), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n16824) );
  AOI22_X1 U20059 ( .A1(n16959), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n16974), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n16823) );
  NAND4_X1 U20060 ( .A1(n16826), .A2(n16825), .A3(n16824), .A4(n16823), .ZN(
        n16832) );
  AOI22_X1 U20061 ( .A1(n9726), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11806), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n16830) );
  AOI22_X1 U20062 ( .A1(n15279), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n16991), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n16829) );
  AOI22_X1 U20063 ( .A1(n9729), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n16968), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n16828) );
  AOI22_X1 U20064 ( .A1(n16988), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n16992), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n16827) );
  NAND4_X1 U20065 ( .A1(n16830), .A2(n16829), .A3(n16828), .A4(n16827), .ZN(
        n16831) );
  NOR2_X1 U20066 ( .A1(n16832), .A2(n16831), .ZN(n17093) );
  OAI22_X1 U20067 ( .A1(n16834), .A2(n16833), .B1(n17093), .B2(n17039), .ZN(
        P3_U2681) );
  NOR2_X1 U20068 ( .A1(n17024), .A2(n16835), .ZN(n16859) );
  AOI22_X1 U20069 ( .A1(n15162), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n16968), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n16846) );
  AOI22_X1 U20070 ( .A1(n16993), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11788), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n16845) );
  INV_X1 U20071 ( .A(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n20872) );
  AOI22_X1 U20072 ( .A1(n15318), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n16974), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n16836) );
  OAI21_X1 U20073 ( .B1(n16837), .B2(n20872), .A(n16836), .ZN(n16843) );
  AOI22_X1 U20074 ( .A1(n9726), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11754), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n16841) );
  AOI22_X1 U20075 ( .A1(n16975), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n9729), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n16840) );
  AOI22_X1 U20076 ( .A1(n17000), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n16991), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n16839) );
  AOI22_X1 U20077 ( .A1(n15279), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n16969), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n16838) );
  NAND4_X1 U20078 ( .A1(n16841), .A2(n16840), .A3(n16839), .A4(n16838), .ZN(
        n16842) );
  AOI211_X1 U20079 ( .C1(n16959), .C2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A(
        n16843), .B(n16842), .ZN(n16844) );
  NAND3_X1 U20080 ( .A1(n16846), .A2(n16845), .A3(n16844), .ZN(n17097) );
  AOI22_X1 U20081 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n16859), .B1(n17024), 
        .B2(n17097), .ZN(n16847) );
  OAI21_X1 U20082 ( .B1(P3_EBX_REG_21__SCAN_IN), .B2(n16848), .A(n16847), .ZN(
        P3_U2682) );
  AOI22_X1 U20083 ( .A1(n15151), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n15279), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n16852) );
  AOI22_X1 U20084 ( .A1(n16954), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n16986), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n16851) );
  AOI22_X1 U20085 ( .A1(n17000), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n16968), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n16850) );
  AOI22_X1 U20086 ( .A1(n11754), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n16969), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n16849) );
  NAND4_X1 U20087 ( .A1(n16852), .A2(n16851), .A3(n16850), .A4(n16849), .ZN(
        n16858) );
  AOI22_X1 U20088 ( .A1(n15162), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n9726), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n16856) );
  AOI22_X1 U20089 ( .A1(n16992), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n16974), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n16855) );
  AOI22_X1 U20090 ( .A1(n16988), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n11806), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n16854) );
  AOI22_X1 U20091 ( .A1(n16993), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n16991), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n16853) );
  NAND4_X1 U20092 ( .A1(n16856), .A2(n16855), .A3(n16854), .A4(n16853), .ZN(
        n16857) );
  NOR2_X1 U20093 ( .A1(n16858), .A2(n16857), .ZN(n17105) );
  INV_X1 U20094 ( .A(n16872), .ZN(n16860) );
  OAI21_X1 U20095 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(n16860), .A(n16859), .ZN(
        n16861) );
  OAI21_X1 U20096 ( .B1(n17105), .B2(n17039), .A(n16861), .ZN(P3_U2683) );
  AOI22_X1 U20097 ( .A1(n15151), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n16986), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n16865) );
  AOI22_X1 U20098 ( .A1(n15162), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n16968), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n16864) );
  AOI22_X1 U20099 ( .A1(n11754), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n16969), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n16863) );
  AOI22_X1 U20100 ( .A1(n16975), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n11806), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n16862) );
  NAND4_X1 U20101 ( .A1(n16865), .A2(n16864), .A3(n16863), .A4(n16862), .ZN(
        n16871) );
  AOI22_X1 U20102 ( .A1(n16993), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n15279), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n16869) );
  AOI22_X1 U20103 ( .A1(n15149), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n16991), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n16868) );
  AOI22_X1 U20104 ( .A1(n9726), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n16974), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n16867) );
  AOI22_X1 U20105 ( .A1(n16954), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11788), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n16866) );
  NAND4_X1 U20106 ( .A1(n16869), .A2(n16868), .A3(n16867), .A4(n16866), .ZN(
        n16870) );
  NOR2_X1 U20107 ( .A1(n16871), .A2(n16870), .ZN(n17110) );
  OAI21_X1 U20108 ( .B1(P3_EBX_REG_19__SCAN_IN), .B2(n9833), .A(n16872), .ZN(
        n16873) );
  AOI22_X1 U20109 ( .A1(n17024), .A2(n17110), .B1(n16873), .B2(n17039), .ZN(
        P3_U2684) );
  NAND2_X1 U20110 ( .A1(n17039), .A2(n16884), .ZN(n16899) );
  AOI22_X1 U20111 ( .A1(n16968), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n16986), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n16883) );
  AOI22_X1 U20112 ( .A1(n16992), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n16974), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n16882) );
  AOI22_X1 U20113 ( .A1(n15279), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n16991), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n16874) );
  OAI21_X1 U20114 ( .B1(n9793), .B2(n20798), .A(n16874), .ZN(n16880) );
  AOI22_X1 U20115 ( .A1(n9726), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11806), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n16878) );
  AOI22_X1 U20116 ( .A1(n16993), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n16954), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n16877) );
  AOI22_X1 U20117 ( .A1(n15162), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n11754), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n16876) );
  AOI22_X1 U20118 ( .A1(n17000), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n16969), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n16875) );
  NAND4_X1 U20119 ( .A1(n16878), .A2(n16877), .A3(n16876), .A4(n16875), .ZN(
        n16879) );
  AOI211_X1 U20120 ( .C1(n9729), .C2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A(
        n16880), .B(n16879), .ZN(n16881) );
  NAND3_X1 U20121 ( .A1(n16883), .A2(n16882), .A3(n16881), .ZN(n17111) );
  NOR3_X1 U20122 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n18052), .A3(n16884), .ZN(
        n16885) );
  AOI21_X1 U20123 ( .B1(n17024), .B2(n17111), .A(n16885), .ZN(n16886) );
  OAI21_X1 U20124 ( .B1(n16887), .B2(n16899), .A(n16886), .ZN(P3_U2685) );
  NOR2_X1 U20125 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n16888), .ZN(n16900) );
  AOI22_X1 U20126 ( .A1(n16968), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n11788), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n16892) );
  AOI22_X1 U20127 ( .A1(n11754), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n16986), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n16891) );
  AOI22_X1 U20128 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n16988), .B1(
        P3_INSTQUEUE_REG_11__1__SCAN_IN), .B2(n16991), .ZN(n16890) );
  AOI22_X1 U20129 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n16969), .B1(
        n9726), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n16889) );
  NAND4_X1 U20130 ( .A1(n16892), .A2(n16891), .A3(n16890), .A4(n16889), .ZN(
        n16898) );
  AOI22_X1 U20131 ( .A1(n17000), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_15__1__SCAN_IN), .B2(n15279), .ZN(n16896) );
  AOI22_X1 U20132 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n16993), .B1(
        n15162), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n16895) );
  AOI22_X1 U20133 ( .A1(n9729), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_0__1__SCAN_IN), .B2(n15318), .ZN(n16894) );
  AOI22_X1 U20134 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n16954), .B1(
        P3_INSTQUEUE_REG_6__1__SCAN_IN), .B2(n16974), .ZN(n16893) );
  NAND4_X1 U20135 ( .A1(n16896), .A2(n16895), .A3(n16894), .A4(n16893), .ZN(
        n16897) );
  NOR2_X1 U20136 ( .A1(n16898), .A2(n16897), .ZN(n17121) );
  OAI22_X1 U20137 ( .A1(n16900), .A2(n16899), .B1(n17121), .B2(n17039), .ZN(
        P3_U2686) );
  NAND4_X1 U20138 ( .A1(P3_EBX_REG_15__SCAN_IN), .A2(P3_EBX_REG_14__SCAN_IN), 
        .A3(P3_EBX_REG_13__SCAN_IN), .A4(n16901), .ZN(n16915) );
  NAND2_X1 U20139 ( .A1(n17039), .A2(n16902), .ZN(n16926) );
  AOI22_X1 U20140 ( .A1(n9726), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11788), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n16912) );
  AOI22_X1 U20141 ( .A1(n16968), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n16974), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n16911) );
  AOI22_X1 U20142 ( .A1(n11754), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n15279), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n16903) );
  OAI21_X1 U20143 ( .B1(n9785), .B2(n20930), .A(n16903), .ZN(n16909) );
  AOI22_X1 U20144 ( .A1(n16993), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n16991), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n16907) );
  AOI22_X1 U20145 ( .A1(n15162), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n16975), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n16906) );
  AOI22_X1 U20146 ( .A1(n17000), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n16987), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n16905) );
  AOI22_X1 U20147 ( .A1(n16959), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n16969), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n16904) );
  NAND4_X1 U20148 ( .A1(n16907), .A2(n16906), .A3(n16905), .A4(n16904), .ZN(
        n16908) );
  AOI211_X1 U20149 ( .C1(n9729), .C2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A(
        n16909), .B(n16908), .ZN(n16910) );
  NAND3_X1 U20150 ( .A1(n16912), .A2(n16911), .A3(n16910), .ZN(n17122) );
  NAND2_X1 U20151 ( .A1(n17024), .A2(n17122), .ZN(n16913) );
  OAI221_X1 U20152 ( .B1(P3_EBX_REG_16__SCAN_IN), .B2(n16915), .C1(n16914), 
        .C2(n16926), .A(n16913), .ZN(P3_U2687) );
  NOR2_X1 U20153 ( .A1(P3_EBX_REG_15__SCAN_IN), .A2(n9763), .ZN(n16927) );
  AOI22_X1 U20154 ( .A1(n9726), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n16986), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n16919) );
  AOI22_X1 U20155 ( .A1(n15162), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n16974), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n16918) );
  AOI22_X1 U20156 ( .A1(n9729), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n16969), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n16917) );
  AOI22_X1 U20157 ( .A1(n16992), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n15279), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n16916) );
  NAND4_X1 U20158 ( .A1(n16919), .A2(n16918), .A3(n16917), .A4(n16916), .ZN(
        n16925) );
  AOI22_X1 U20159 ( .A1(n16968), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n16991), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n16923) );
  AOI22_X1 U20160 ( .A1(n17000), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n16987), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n16922) );
  AOI22_X1 U20161 ( .A1(n11754), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n11806), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n16921) );
  AOI22_X1 U20162 ( .A1(n16993), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n16975), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n16920) );
  NAND4_X1 U20163 ( .A1(n16923), .A2(n16922), .A3(n16921), .A4(n16920), .ZN(
        n16924) );
  NOR2_X1 U20164 ( .A1(n16925), .A2(n16924), .ZN(n17131) );
  OAI22_X1 U20165 ( .A1(n16927), .A2(n16926), .B1(n17131), .B2(n17039), .ZN(
        P3_U2688) );
  AOI22_X1 U20166 ( .A1(n9726), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n16991), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n16931) );
  AOI22_X1 U20167 ( .A1(n15162), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n16975), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n16930) );
  AOI22_X1 U20168 ( .A1(n16992), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11806), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n16929) );
  AOI22_X1 U20169 ( .A1(n16969), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n16974), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n16928) );
  NAND4_X1 U20170 ( .A1(n16931), .A2(n16930), .A3(n16929), .A4(n16928), .ZN(
        n16937) );
  AOI22_X1 U20171 ( .A1(n9729), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n15279), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n16935) );
  AOI22_X1 U20172 ( .A1(n16968), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n16954), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n16934) );
  AOI22_X1 U20173 ( .A1(n16993), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n16959), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n16933) );
  AOI22_X1 U20174 ( .A1(n17000), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11754), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n16932) );
  NAND4_X1 U20175 ( .A1(n16935), .A2(n16934), .A3(n16933), .A4(n16932), .ZN(
        n16936) );
  NOR2_X1 U20176 ( .A1(n16937), .A2(n16936), .ZN(n17142) );
  NOR2_X1 U20177 ( .A1(n17024), .A2(n16939), .ZN(n16951) );
  OAI222_X1 U20178 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n17047), .B1(
        P3_EBX_REG_12__SCAN_IN), .B2(n16939), .C1(n16951), .C2(n16938), .ZN(
        n16940) );
  OAI21_X1 U20179 ( .B1(n17142), .B2(n17039), .A(n16940), .ZN(P3_U2691) );
  AOI22_X1 U20180 ( .A1(n16975), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11806), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n16944) );
  AOI22_X1 U20181 ( .A1(n16992), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n16991), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n16943) );
  AOI22_X1 U20182 ( .A1(n9729), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n16954), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n16942) );
  AOI22_X1 U20183 ( .A1(n15279), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n16969), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n16941) );
  NAND4_X1 U20184 ( .A1(n16944), .A2(n16943), .A3(n16942), .A4(n16941), .ZN(
        n16950) );
  AOI22_X1 U20185 ( .A1(n17000), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n16993), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n16948) );
  AOI22_X1 U20186 ( .A1(n15162), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n16968), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n16947) );
  AOI22_X1 U20187 ( .A1(n11754), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n16974), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n16946) );
  AOI22_X1 U20188 ( .A1(n9726), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n16959), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n16945) );
  NAND4_X1 U20189 ( .A1(n16948), .A2(n16947), .A3(n16946), .A4(n16945), .ZN(
        n16949) );
  NOR2_X1 U20190 ( .A1(n16950), .A2(n16949), .ZN(n17146) );
  OAI21_X1 U20191 ( .B1(P3_EBX_REG_11__SCAN_IN), .B2(n16952), .A(n16951), .ZN(
        n16953) );
  OAI21_X1 U20192 ( .B1(n17146), .B2(n17039), .A(n16953), .ZN(P3_U2692) );
  AOI22_X1 U20193 ( .A1(n16954), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n16991), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n16958) );
  AOI22_X1 U20194 ( .A1(n17000), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n15162), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n16957) );
  AOI22_X1 U20195 ( .A1(n16993), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n16975), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n16956) );
  AOI22_X1 U20196 ( .A1(n15279), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n16969), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n16955) );
  NAND4_X1 U20197 ( .A1(n16958), .A2(n16957), .A3(n16956), .A4(n16955), .ZN(
        n16965) );
  AOI22_X1 U20198 ( .A1(n9729), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n16974), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n16963) );
  AOI22_X1 U20199 ( .A1(n16968), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n16959), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n16962) );
  AOI22_X1 U20200 ( .A1(n11754), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n11806), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n16961) );
  AOI22_X1 U20201 ( .A1(n9726), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11788), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n16960) );
  NAND4_X1 U20202 ( .A1(n16963), .A2(n16962), .A3(n16961), .A4(n16960), .ZN(
        n16964) );
  NOR2_X1 U20203 ( .A1(n16965), .A2(n16964), .ZN(n17153) );
  OAI22_X1 U20204 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n18052), .B1(n17024), 
        .B2(n16982), .ZN(n16966) );
  OAI21_X1 U20205 ( .B1(P3_EBX_REG_10__SCAN_IN), .B2(n16982), .A(n16966), .ZN(
        n16967) );
  OAI21_X1 U20206 ( .B1(n17153), .B2(n17039), .A(n16967), .ZN(P3_U2693) );
  AOI22_X1 U20207 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n16987), .B1(
        n11754), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n16973) );
  AOI22_X1 U20208 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n16968), .B1(
        n15279), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n16972) );
  AOI22_X1 U20209 ( .A1(n17000), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_15__1__SCAN_IN), .B2(n11806), .ZN(n16971) );
  AOI22_X1 U20210 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n16969), .B1(
        P3_INSTQUEUE_REG_11__1__SCAN_IN), .B2(n16777), .ZN(n16970) );
  NAND4_X1 U20211 ( .A1(n16973), .A2(n16972), .A3(n16971), .A4(n16970), .ZN(
        n16981) );
  AOI22_X1 U20212 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n16991), .B1(
        P3_INSTQUEUE_REG_5__1__SCAN_IN), .B2(n16974), .ZN(n16979) );
  AOI22_X1 U20213 ( .A1(n16993), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_7__1__SCAN_IN), .B2(n9726), .ZN(n16978) );
  AOI22_X1 U20214 ( .A1(n9729), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n16986), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n16977) );
  AOI22_X1 U20215 ( .A1(n15162), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n16975), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n16976) );
  NAND4_X1 U20216 ( .A1(n16979), .A2(n16978), .A3(n16977), .A4(n16976), .ZN(
        n16980) );
  NOR2_X1 U20217 ( .A1(n16981), .A2(n16980), .ZN(n17156) );
  NOR2_X1 U20218 ( .A1(n17024), .A2(n16982), .ZN(n16983) );
  OAI21_X1 U20219 ( .B1(P3_EBX_REG_9__SCAN_IN), .B2(n17006), .A(n16983), .ZN(
        n16984) );
  OAI21_X1 U20220 ( .B1(n17156), .B2(n17039), .A(n16984), .ZN(P3_U2694) );
  AND2_X1 U20221 ( .A1(n17047), .A2(n17015), .ZN(n17018) );
  NAND2_X1 U20222 ( .A1(P3_EBX_REG_5__SCAN_IN), .A2(n17018), .ZN(n17014) );
  INV_X1 U20223 ( .A(n17014), .ZN(n17008) );
  AOI22_X1 U20224 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n17039), .B1(n16985), .B2(
        n17008), .ZN(n17005) );
  AOI22_X1 U20225 ( .A1(n15118), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n11754), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n17003) );
  AOI22_X1 U20226 ( .A1(n15162), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n16986), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n17002) );
  AOI22_X1 U20227 ( .A1(n16988), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n16987), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n16989) );
  OAI21_X1 U20228 ( .B1(n16990), .B2(n20930), .A(n16989), .ZN(n16999) );
  AOI22_X1 U20229 ( .A1(n16992), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n16991), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n16997) );
  AOI22_X1 U20230 ( .A1(n16968), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n16974), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n16996) );
  AOI22_X1 U20231 ( .A1(n15279), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11806), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n16995) );
  AOI22_X1 U20232 ( .A1(n16993), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n9729), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n16994) );
  NAND4_X1 U20233 ( .A1(n16997), .A2(n16996), .A3(n16995), .A4(n16994), .ZN(
        n16998) );
  AOI211_X1 U20234 ( .C1(n17000), .C2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A(
        n16999), .B(n16998), .ZN(n17001) );
  NAND3_X1 U20235 ( .A1(n17003), .A2(n17002), .A3(n17001), .ZN(n17161) );
  INV_X1 U20236 ( .A(n17161), .ZN(n17004) );
  OAI22_X1 U20237 ( .A1(n17006), .A2(n17005), .B1(n17004), .B2(n17039), .ZN(
        P3_U2695) );
  NOR2_X1 U20238 ( .A1(n17007), .A2(n17014), .ZN(n17011) );
  AOI22_X1 U20239 ( .A1(P3_EBX_REG_7__SCAN_IN), .A2(n17039), .B1(
        P3_EBX_REG_6__SCAN_IN), .B2(n17008), .ZN(n17010) );
  OAI22_X1 U20240 ( .A1(n17011), .A2(n17010), .B1(n17009), .B2(n17039), .ZN(
        P3_U2696) );
  INV_X1 U20241 ( .A(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17013) );
  NAND3_X1 U20242 ( .A1(n17014), .A2(P3_EBX_REG_6__SCAN_IN), .A3(n17039), .ZN(
        n17012) );
  OAI221_X1 U20243 ( .B1(n17014), .B2(P3_EBX_REG_6__SCAN_IN), .C1(n17039), 
        .C2(n17013), .A(n17012), .ZN(P3_U2697) );
  INV_X1 U20244 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n17017) );
  OAI211_X1 U20245 ( .C1(P3_EBX_REG_5__SCAN_IN), .C2(n17015), .A(n17014), .B(
        n17039), .ZN(n17016) );
  OAI21_X1 U20246 ( .B1(n17039), .B2(n17017), .A(n17016), .ZN(P3_U2698) );
  AOI21_X1 U20247 ( .B1(n17020), .B2(n17019), .A(n17018), .ZN(n17021) );
  OAI22_X1 U20248 ( .A1(n17039), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n17021), .B2(n17024), .ZN(n17022) );
  INV_X1 U20249 ( .A(n17022), .ZN(P3_U2699) );
  NAND2_X1 U20250 ( .A1(n17047), .A2(n17023), .ZN(n17026) );
  NOR2_X1 U20251 ( .A1(n17024), .A2(n17023), .ZN(n17028) );
  AOI22_X1 U20252 ( .A1(P3_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n17024), .B1(
        P3_EBX_REG_3__SCAN_IN), .B2(n17028), .ZN(n17025) );
  OAI21_X1 U20253 ( .B1(P3_EBX_REG_3__SCAN_IN), .B2(n17026), .A(n17025), .ZN(
        P3_U2700) );
  INV_X1 U20254 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17031) );
  INV_X1 U20255 ( .A(n17027), .ZN(n17029) );
  OAI21_X1 U20256 ( .B1(P3_EBX_REG_2__SCAN_IN), .B2(n17029), .A(n17028), .ZN(
        n17030) );
  OAI21_X1 U20257 ( .B1(n17039), .B2(n17031), .A(n17030), .ZN(P3_U2701) );
  INV_X1 U20258 ( .A(n17032), .ZN(n17036) );
  INV_X1 U20259 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17033) );
  OAI222_X1 U20260 ( .A1(n17036), .A2(n17037), .B1(n17035), .B2(n17034), .C1(
        n17033), .C2(n17039), .ZN(P3_U2702) );
  AND2_X1 U20261 ( .A1(n17038), .A2(n17037), .ZN(n17040) );
  OAI22_X1 U20262 ( .A1(n17041), .A2(n17040), .B1(n20930), .B2(n17039), .ZN(
        P3_U2703) );
  INV_X1 U20263 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n17266) );
  INV_X1 U20264 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n20918) );
  INV_X1 U20265 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n17303) );
  INV_X1 U20266 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n17284) );
  NAND2_X1 U20267 ( .A1(P3_EAX_REG_1__SCAN_IN), .A2(P3_EAX_REG_0__SCAN_IN), 
        .ZN(n17194) );
  NAND4_X1 U20268 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(P3_EAX_REG_2__SCAN_IN), 
        .A3(P3_EAX_REG_5__SCAN_IN), .A4(P3_EAX_REG_4__SCAN_IN), .ZN(n17042) );
  NOR2_X1 U20269 ( .A1(n17194), .A2(n17042), .ZN(n17174) );
  NAND4_X1 U20270 ( .A1(P3_EAX_REG_14__SCAN_IN), .A2(P3_EAX_REG_13__SCAN_IN), 
        .A3(P3_EAX_REG_11__SCAN_IN), .A4(P3_EAX_REG_10__SCAN_IN), .ZN(n17044)
         );
  NAND4_X1 U20271 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(P3_EAX_REG_8__SCAN_IN), 
        .A3(P3_EAX_REG_9__SCAN_IN), .A4(n17045), .ZN(n17133) );
  NOR2_X2 U20272 ( .A1(n17303), .A2(n17133), .ZN(n17128) );
  NAND2_X1 U20273 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(P3_EAX_REG_18__SCAN_IN), 
        .ZN(n17092) );
  NAND4_X1 U20274 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(P3_EAX_REG_21__SCAN_IN), 
        .A3(P3_EAX_REG_20__SCAN_IN), .A4(P3_EAX_REG_17__SCAN_IN), .ZN(n17046)
         );
  NOR3_X2 U20275 ( .A1(n17124), .A2(n17092), .A3(n17046), .ZN(n17088) );
  NAND2_X1 U20276 ( .A1(P3_EAX_REG_23__SCAN_IN), .A2(n17088), .ZN(n17087) );
  NAND2_X1 U20277 ( .A1(P3_EAX_REG_24__SCAN_IN), .A2(n17083), .ZN(n17082) );
  NAND2_X1 U20278 ( .A1(P3_EAX_REG_29__SCAN_IN), .A2(n17060), .ZN(n17056) );
  NAND2_X1 U20279 ( .A1(P3_EAX_REG_30__SCAN_IN), .A2(n17052), .ZN(n17051) );
  NAND2_X1 U20280 ( .A1(n17051), .A2(P3_EAX_REG_31__SCAN_IN), .ZN(n17050) );
  NOR2_X2 U20281 ( .A1(n17048), .A2(n17180), .ZN(n17116) );
  NAND2_X1 U20282 ( .A1(BUF2_REG_31__SCAN_IN), .A2(n17116), .ZN(n17049) );
  OAI221_X1 U20283 ( .B1(n17051), .B2(P3_EAX_REG_31__SCAN_IN), .C1(n17050), 
        .C2(n17185), .A(n17049), .ZN(P3_U2704) );
  NOR2_X2 U20284 ( .A1(n18041), .A2(n17180), .ZN(n17123) );
  AOI22_X1 U20285 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17123), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n17116), .ZN(n17054) );
  OAI211_X1 U20286 ( .C1(n17052), .C2(P3_EAX_REG_30__SCAN_IN), .A(n17180), .B(
        n17051), .ZN(n17053) );
  OAI211_X1 U20287 ( .C1(n17055), .C2(n17198), .A(n17054), .B(n17053), .ZN(
        P3_U2705) );
  AOI22_X1 U20288 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17123), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n17116), .ZN(n17058) );
  OAI211_X1 U20289 ( .C1(n17060), .C2(P3_EAX_REG_29__SCAN_IN), .A(n17180), .B(
        n17056), .ZN(n17057) );
  OAI211_X1 U20290 ( .C1(n17198), .C2(n17059), .A(n17058), .B(n17057), .ZN(
        P3_U2706) );
  AOI22_X1 U20291 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17123), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n17116), .ZN(n17063) );
  AOI211_X1 U20292 ( .C1(n17266), .C2(n17068), .A(n17060), .B(n17185), .ZN(
        n17061) );
  INV_X1 U20293 ( .A(n17061), .ZN(n17062) );
  OAI211_X1 U20294 ( .C1(n17198), .C2(n17064), .A(n17063), .B(n17062), .ZN(
        P3_U2707) );
  OAI21_X1 U20295 ( .B1(n17067), .B2(n17066), .A(n17065), .ZN(n17071) );
  AOI22_X1 U20296 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17123), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n17116), .ZN(n17070) );
  OAI211_X1 U20297 ( .C1(n17073), .C2(P3_EAX_REG_27__SCAN_IN), .A(n17180), .B(
        n17068), .ZN(n17069) );
  OAI211_X1 U20298 ( .C1(n17198), .C2(n17071), .A(n17070), .B(n17069), .ZN(
        P3_U2708) );
  INV_X1 U20299 ( .A(n17116), .ZN(n17127) );
  AOI22_X1 U20300 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17123), .B1(n17072), .B2(
        n17188), .ZN(n17076) );
  AOI211_X1 U20301 ( .C1(n20918), .C2(n17077), .A(n17073), .B(n17185), .ZN(
        n17074) );
  INV_X1 U20302 ( .A(n17074), .ZN(n17075) );
  OAI211_X1 U20303 ( .C1(n17127), .C2(n18029), .A(n17076), .B(n17075), .ZN(
        P3_U2709) );
  AOI22_X1 U20304 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17123), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n17116), .ZN(n17080) );
  OAI211_X1 U20305 ( .C1(n17078), .C2(P3_EAX_REG_25__SCAN_IN), .A(n17180), .B(
        n17077), .ZN(n17079) );
  OAI211_X1 U20306 ( .C1(n17198), .C2(n17081), .A(n17080), .B(n17079), .ZN(
        P3_U2710) );
  AOI22_X1 U20307 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17123), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n17116), .ZN(n17085) );
  OAI211_X1 U20308 ( .C1(n17083), .C2(P3_EAX_REG_24__SCAN_IN), .A(n17180), .B(
        n17082), .ZN(n17084) );
  OAI211_X1 U20309 ( .C1(n17198), .C2(n17086), .A(n17085), .B(n17084), .ZN(
        P3_U2711) );
  AOI22_X1 U20310 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17123), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n17116), .ZN(n17090) );
  OAI211_X1 U20311 ( .C1(P3_EAX_REG_23__SCAN_IN), .C2(n17088), .A(n17180), .B(
        n17087), .ZN(n17089) );
  OAI211_X1 U20312 ( .C1(n17198), .C2(n17091), .A(n17090), .B(n17089), .ZN(
        P3_U2712) );
  INV_X1 U20313 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n17245) );
  INV_X1 U20314 ( .A(n17113), .ZN(n17117) );
  NAND2_X1 U20315 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n17106), .ZN(n17102) );
  NAND2_X1 U20316 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(n17099), .ZN(n17098) );
  NAND2_X1 U20317 ( .A1(n17098), .A2(P3_EAX_REG_22__SCAN_IN), .ZN(n17096) );
  OAI22_X1 U20318 ( .A1(n17093), .A2(n17198), .B1(n18047), .B2(n17127), .ZN(
        n17094) );
  AOI21_X1 U20319 ( .B1(BUF2_REG_6__SCAN_IN), .B2(n17123), .A(n17094), .ZN(
        n17095) );
  OAI221_X1 U20320 ( .B1(n17098), .B2(P3_EAX_REG_22__SCAN_IN), .C1(n17096), 
        .C2(n17185), .A(n17095), .ZN(P3_U2713) );
  AOI22_X1 U20321 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17123), .B1(n17188), .B2(
        n17097), .ZN(n17101) );
  OAI211_X1 U20322 ( .C1(n17099), .C2(P3_EAX_REG_21__SCAN_IN), .A(n17180), .B(
        n17098), .ZN(n17100) );
  OAI211_X1 U20323 ( .C1(n17127), .C2(n18042), .A(n17101), .B(n17100), .ZN(
        P3_U2714) );
  AOI22_X1 U20324 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17123), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n17116), .ZN(n17104) );
  OAI211_X1 U20325 ( .C1(n17106), .C2(P3_EAX_REG_20__SCAN_IN), .A(n17180), .B(
        n17102), .ZN(n17103) );
  OAI211_X1 U20326 ( .C1(n17105), .C2(n17198), .A(n17104), .B(n17103), .ZN(
        P3_U2715) );
  AOI22_X1 U20327 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17123), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n17116), .ZN(n17109) );
  INV_X1 U20328 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n17249) );
  NAND2_X1 U20329 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n17113), .ZN(n17112) );
  AOI211_X1 U20330 ( .C1(n17249), .C2(n17112), .A(n17106), .B(n17185), .ZN(
        n17107) );
  INV_X1 U20331 ( .A(n17107), .ZN(n17108) );
  OAI211_X1 U20332 ( .C1(n17110), .C2(n17198), .A(n17109), .B(n17108), .ZN(
        P3_U2716) );
  AOI22_X1 U20333 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17123), .B1(n17188), .B2(
        n17111), .ZN(n17115) );
  OAI211_X1 U20334 ( .C1(n17113), .C2(P3_EAX_REG_18__SCAN_IN), .A(n17180), .B(
        n17112), .ZN(n17114) );
  OAI211_X1 U20335 ( .C1(n17127), .C2(n19070), .A(n17115), .B(n17114), .ZN(
        P3_U2717) );
  AOI22_X1 U20336 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17123), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n17116), .ZN(n17120) );
  INV_X1 U20337 ( .A(n17124), .ZN(n17118) );
  OAI211_X1 U20338 ( .C1(n17118), .C2(P3_EAX_REG_17__SCAN_IN), .A(n17180), .B(
        n17117), .ZN(n17119) );
  OAI211_X1 U20339 ( .C1(n17121), .C2(n17198), .A(n17120), .B(n17119), .ZN(
        P3_U2718) );
  AOI22_X1 U20340 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17123), .B1(n17188), .B2(
        n17122), .ZN(n17126) );
  OAI211_X1 U20341 ( .C1(P3_EAX_REG_16__SCAN_IN), .C2(n17128), .A(n17180), .B(
        n17124), .ZN(n17125) );
  OAI211_X1 U20342 ( .C1(n17127), .C2(n18018), .A(n17126), .B(n17125), .ZN(
        P3_U2719) );
  AOI211_X1 U20343 ( .C1(n17303), .C2(n17133), .A(n17185), .B(n17128), .ZN(
        n17129) );
  AOI21_X1 U20344 ( .B1(n17193), .B2(BUF2_REG_15__SCAN_IN), .A(n17129), .ZN(
        n17130) );
  OAI21_X1 U20345 ( .B1(n17131), .B2(n17198), .A(n17130), .ZN(P3_U2720) );
  INV_X1 U20346 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n20936) );
  INV_X1 U20347 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n17290) );
  INV_X1 U20348 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n20741) );
  NOR3_X1 U20349 ( .A1(n18052), .A2(n17160), .A3(n20741), .ZN(n17155) );
  NAND2_X1 U20350 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(n17155), .ZN(n17154) );
  NOR2_X1 U20351 ( .A1(n17290), .A2(n17154), .ZN(n17150) );
  NAND2_X1 U20352 ( .A1(P3_EAX_REG_11__SCAN_IN), .A2(n17150), .ZN(n17141) );
  NOR2_X1 U20353 ( .A1(n20936), .A2(n17141), .ZN(n17144) );
  NAND2_X1 U20354 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n17144), .ZN(n17136) );
  AOI22_X1 U20355 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17193), .B1(n17188), .B2(
        n17132), .ZN(n17135) );
  NAND3_X1 U20356 ( .A1(P3_EAX_REG_14__SCAN_IN), .A2(n17180), .A3(n17133), 
        .ZN(n17134) );
  OAI211_X1 U20357 ( .C1(P3_EAX_REG_14__SCAN_IN), .C2(n17136), .A(n17135), .B(
        n17134), .ZN(P3_U2721) );
  INV_X1 U20358 ( .A(n17193), .ZN(n17184) );
  INV_X1 U20359 ( .A(n17136), .ZN(n17139) );
  AOI21_X1 U20360 ( .B1(P3_EAX_REG_13__SCAN_IN), .B2(n17180), .A(n17144), .ZN(
        n17138) );
  OAI222_X1 U20361 ( .A1(n17184), .A2(n17140), .B1(n17139), .B2(n17138), .C1(
        n17198), .C2(n17137), .ZN(P3_U2722) );
  INV_X1 U20362 ( .A(n17141), .ZN(n17148) );
  AOI21_X1 U20363 ( .B1(P3_EAX_REG_12__SCAN_IN), .B2(n17180), .A(n17148), .ZN(
        n17143) );
  OAI222_X1 U20364 ( .A1(n17184), .A2(n17145), .B1(n17144), .B2(n17143), .C1(
        n17198), .C2(n17142), .ZN(P3_U2723) );
  AOI21_X1 U20365 ( .B1(P3_EAX_REG_11__SCAN_IN), .B2(n17180), .A(n17150), .ZN(
        n17147) );
  OAI222_X1 U20366 ( .A1(n17184), .A2(n17149), .B1(n17148), .B2(n17147), .C1(
        n17198), .C2(n17146), .ZN(P3_U2724) );
  AOI211_X1 U20367 ( .C1(n17290), .C2(n17154), .A(n17185), .B(n17150), .ZN(
        n17151) );
  AOI21_X1 U20368 ( .B1(n17193), .B2(BUF2_REG_10__SCAN_IN), .A(n17151), .ZN(
        n17152) );
  OAI21_X1 U20369 ( .B1(n17153), .B2(n17198), .A(n17152), .ZN(P3_U2725) );
  INV_X1 U20370 ( .A(n17154), .ZN(n17158) );
  AOI21_X1 U20371 ( .B1(P3_EAX_REG_9__SCAN_IN), .B2(n17180), .A(n17155), .ZN(
        n17157) );
  OAI222_X1 U20372 ( .A1(n17184), .A2(n17159), .B1(n17158), .B2(n17157), .C1(
        n17198), .C2(n17156), .ZN(P3_U2726) );
  OR2_X1 U20373 ( .A1(n18052), .A2(n17160), .ZN(n17163) );
  NAND2_X1 U20374 ( .A1(n17180), .A2(n17160), .ZN(n17165) );
  AOI22_X1 U20375 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17193), .B1(n17188), .B2(
        n17161), .ZN(n17162) );
  OAI221_X1 U20376 ( .B1(P3_EAX_REG_8__SCAN_IN), .B2(n17163), .C1(n20741), 
        .C2(n17165), .A(n17162), .ZN(P3_U2727) );
  NOR2_X1 U20377 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(n17167), .ZN(n17164) );
  OAI222_X1 U20378 ( .A1(n17184), .A2(n18055), .B1(n17198), .B2(n17166), .C1(
        n17165), .C2(n17164), .ZN(P3_U2728) );
  AOI211_X1 U20379 ( .C1(n17284), .C2(n17168), .A(n17185), .B(n17167), .ZN(
        n17169) );
  AOI21_X1 U20380 ( .B1(n17193), .B2(BUF2_REG_6__SCAN_IN), .A(n17169), .ZN(
        n17170) );
  OAI21_X1 U20381 ( .B1(n17171), .B2(n17198), .A(n17170), .ZN(P3_U2729) );
  INV_X1 U20382 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n17278) );
  INV_X1 U20383 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n17276) );
  NOR3_X1 U20384 ( .A1(n17276), .A2(n17194), .A3(n17186), .ZN(n17179) );
  INV_X1 U20385 ( .A(n17179), .ZN(n17190) );
  NOR2_X1 U20386 ( .A1(n17278), .A2(n17190), .ZN(n17182) );
  AND2_X1 U20387 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(n17182), .ZN(n17177) );
  AOI21_X1 U20388 ( .B1(P3_EAX_REG_5__SCAN_IN), .B2(n17180), .A(n17177), .ZN(
        n17175) );
  INV_X1 U20389 ( .A(n17186), .ZN(n17195) );
  AOI22_X1 U20390 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17193), .B1(n17188), .B2(
        n17172), .ZN(n17173) );
  OAI221_X1 U20391 ( .B1(n17175), .B2(n17174), .C1(n17175), .C2(n17195), .A(
        n17173), .ZN(P3_U2730) );
  AOI21_X1 U20392 ( .B1(P3_EAX_REG_4__SCAN_IN), .B2(n17180), .A(n17182), .ZN(
        n17178) );
  OAI222_X1 U20393 ( .A1(n17184), .A2(n18038), .B1(n17178), .B2(n17177), .C1(
        n17198), .C2(n17176), .ZN(P3_U2731) );
  AOI21_X1 U20394 ( .B1(P3_EAX_REG_3__SCAN_IN), .B2(n17180), .A(n17179), .ZN(
        n17183) );
  OAI222_X1 U20395 ( .A1(n17184), .A2(n18033), .B1(n17183), .B2(n17182), .C1(
        n17198), .C2(n17181), .ZN(P3_U2732) );
  OAI22_X1 U20396 ( .A1(n17186), .A2(n17194), .B1(n17276), .B2(n17185), .ZN(
        n17189) );
  AOI222_X1 U20397 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17193), .B1(n17190), .B2(
        n17189), .C1(n17188), .C2(n17187), .ZN(n17191) );
  INV_X1 U20398 ( .A(n17191), .ZN(P3_U2733) );
  AOI22_X1 U20399 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17193), .B1(
        P3_EAX_REG_1__SCAN_IN), .B2(n17192), .ZN(n17197) );
  OAI211_X1 U20400 ( .C1(P3_EAX_REG_1__SCAN_IN), .C2(P3_EAX_REG_0__SCAN_IN), 
        .A(n17195), .B(n17194), .ZN(n17196) );
  OAI211_X1 U20401 ( .C1(n17199), .C2(n17198), .A(n17197), .B(n17196), .ZN(
        P3_U2734) );
  NAND2_X1 U20402 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n17387), .ZN(n18649) );
  INV_X2 U20403 ( .A(n18649), .ZN(n17235) );
  AND2_X1 U20404 ( .A1(n17215), .A2(P3_DATAO_REG_31__SCAN_IN), .ZN(P3_U2736)
         );
  INV_X1 U20405 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n17270) );
  NAND2_X1 U20406 ( .A1(n17218), .A2(n18012), .ZN(n17217) );
  AOI22_X1 U20407 ( .A1(n17235), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(
        P3_DATAO_REG_30__SCAN_IN), .B2(n17234), .ZN(n17201) );
  OAI21_X1 U20408 ( .B1(n17270), .B2(n17217), .A(n17201), .ZN(P3_U2737) );
  INV_X1 U20409 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n17268) );
  AOI22_X1 U20410 ( .A1(n17235), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n17234), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n17202) );
  OAI21_X1 U20411 ( .B1(n17268), .B2(n17217), .A(n17202), .ZN(P3_U2738) );
  AOI22_X1 U20412 ( .A1(n17235), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n17234), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n17203) );
  OAI21_X1 U20413 ( .B1(n17266), .B2(n17217), .A(n17203), .ZN(P3_U2739) );
  INV_X1 U20414 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n17264) );
  AOI22_X1 U20415 ( .A1(n17235), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n17215), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n17204) );
  OAI21_X1 U20416 ( .B1(n17264), .B2(n17217), .A(n17204), .ZN(P3_U2740) );
  AOI22_X1 U20417 ( .A1(n17235), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n17215), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n17205) );
  OAI21_X1 U20418 ( .B1(n20918), .B2(n17217), .A(n17205), .ZN(P3_U2741) );
  INV_X1 U20419 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n17261) );
  AOI22_X1 U20420 ( .A1(n17235), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n17234), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n17206) );
  OAI21_X1 U20421 ( .B1(n17261), .B2(n17217), .A(n17206), .ZN(P3_U2742) );
  INV_X1 U20422 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n17259) );
  AOI22_X1 U20423 ( .A1(n17235), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n17215), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n17207) );
  OAI21_X1 U20424 ( .B1(n17259), .B2(n17217), .A(n17207), .ZN(P3_U2743) );
  INV_X1 U20425 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n17257) );
  AOI22_X1 U20426 ( .A1(n17235), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n17234), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n17208) );
  OAI21_X1 U20427 ( .B1(n17257), .B2(n17217), .A(n17208), .ZN(P3_U2744) );
  INV_X1 U20428 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n17255) );
  AOI22_X1 U20429 ( .A1(n17235), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n17215), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n17209) );
  OAI21_X1 U20430 ( .B1(n17255), .B2(n17217), .A(n17209), .ZN(P3_U2745) );
  INV_X1 U20431 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n17253) );
  AOI22_X1 U20432 ( .A1(n17235), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n17215), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n17210) );
  OAI21_X1 U20433 ( .B1(n17253), .B2(n17217), .A(n17210), .ZN(P3_U2746) );
  INV_X1 U20434 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n17251) );
  AOI22_X1 U20435 ( .A1(n17235), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n17215), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n17211) );
  OAI21_X1 U20436 ( .B1(n17251), .B2(n17217), .A(n17211), .ZN(P3_U2747) );
  AOI22_X1 U20437 ( .A1(n17235), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n17215), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n17212) );
  OAI21_X1 U20438 ( .B1(n17249), .B2(n17217), .A(n17212), .ZN(P3_U2748) );
  INV_X1 U20439 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n17247) );
  AOI22_X1 U20440 ( .A1(n17235), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n17215), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n17213) );
  OAI21_X1 U20441 ( .B1(n17247), .B2(n17217), .A(n17213), .ZN(P3_U2749) );
  AOI22_X1 U20442 ( .A1(n17235), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n17215), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n17214) );
  OAI21_X1 U20443 ( .B1(n17245), .B2(n17217), .A(n17214), .ZN(P3_U2750) );
  INV_X1 U20444 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n17243) );
  AOI22_X1 U20445 ( .A1(n17235), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n17215), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n17216) );
  OAI21_X1 U20446 ( .B1(n17243), .B2(n17217), .A(n17216), .ZN(P3_U2751) );
  AOI22_X1 U20447 ( .A1(n17235), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n17234), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n17219) );
  OAI21_X1 U20448 ( .B1(n17303), .B2(n17237), .A(n17219), .ZN(P3_U2752) );
  INV_X1 U20449 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n17299) );
  AOI22_X1 U20450 ( .A1(n17235), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n17234), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n17220) );
  OAI21_X1 U20451 ( .B1(n17299), .B2(n17237), .A(n17220), .ZN(P3_U2753) );
  INV_X1 U20452 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n17297) );
  AOI22_X1 U20453 ( .A1(n17235), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n17234), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n17221) );
  OAI21_X1 U20454 ( .B1(n17297), .B2(n17237), .A(n17221), .ZN(P3_U2754) );
  AOI22_X1 U20455 ( .A1(n17235), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n17234), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n17222) );
  OAI21_X1 U20456 ( .B1(n20936), .B2(n17237), .A(n17222), .ZN(P3_U2755) );
  INV_X1 U20457 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n17292) );
  AOI22_X1 U20458 ( .A1(n17235), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n17234), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n17223) );
  OAI21_X1 U20459 ( .B1(n17292), .B2(n17237), .A(n17223), .ZN(P3_U2756) );
  AOI22_X1 U20460 ( .A1(n17235), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n17234), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n17224) );
  OAI21_X1 U20461 ( .B1(n17290), .B2(n17237), .A(n17224), .ZN(P3_U2757) );
  INV_X1 U20462 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n17288) );
  AOI22_X1 U20463 ( .A1(n17235), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n17234), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n17225) );
  OAI21_X1 U20464 ( .B1(n17288), .B2(n17237), .A(n17225), .ZN(P3_U2758) );
  AOI22_X1 U20465 ( .A1(n17235), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n17234), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n17226) );
  OAI21_X1 U20466 ( .B1(n20741), .B2(n17237), .A(n17226), .ZN(P3_U2759) );
  INV_X1 U20467 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n20896) );
  AOI22_X1 U20468 ( .A1(n17235), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n17234), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n17227) );
  OAI21_X1 U20469 ( .B1(n20896), .B2(n17237), .A(n17227), .ZN(P3_U2760) );
  AOI22_X1 U20470 ( .A1(n17235), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n17234), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n17228) );
  OAI21_X1 U20471 ( .B1(n17284), .B2(n17237), .A(n17228), .ZN(P3_U2761) );
  INV_X1 U20472 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n17282) );
  AOI22_X1 U20473 ( .A1(n17235), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n17234), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n17229) );
  OAI21_X1 U20474 ( .B1(n17282), .B2(n17237), .A(n17229), .ZN(P3_U2762) );
  INV_X1 U20475 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n17280) );
  AOI22_X1 U20476 ( .A1(n17235), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n17234), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n17230) );
  OAI21_X1 U20477 ( .B1(n17280), .B2(n17237), .A(n17230), .ZN(P3_U2763) );
  AOI22_X1 U20478 ( .A1(n17235), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n17234), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n17231) );
  OAI21_X1 U20479 ( .B1(n17278), .B2(n17237), .A(n17231), .ZN(P3_U2764) );
  AOI22_X1 U20480 ( .A1(n17235), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n17234), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n17232) );
  OAI21_X1 U20481 ( .B1(n17276), .B2(n17237), .A(n17232), .ZN(P3_U2765) );
  INV_X1 U20482 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n17274) );
  AOI22_X1 U20483 ( .A1(n17235), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n17234), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n17233) );
  OAI21_X1 U20484 ( .B1(n17274), .B2(n17237), .A(n17233), .ZN(P3_U2766) );
  AOI22_X1 U20485 ( .A1(n17235), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n17234), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n17236) );
  OAI21_X1 U20486 ( .B1(n17272), .B2(n17237), .A(n17236), .ZN(P3_U2767) );
  INV_X1 U20487 ( .A(n17238), .ZN(n17240) );
  NOR2_X1 U20488 ( .A1(n18023), .A2(n17239), .ZN(n18496) );
  NAND2_X2 U20489 ( .A1(n17240), .A2(n18496), .ZN(n17302) );
  AOI22_X1 U20490 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17294), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n17293), .ZN(n17242) );
  OAI21_X1 U20491 ( .B1(n17243), .B2(n17302), .A(n17242), .ZN(P3_U2768) );
  AOI22_X1 U20492 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17294), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n17293), .ZN(n17244) );
  OAI21_X1 U20493 ( .B1(n17245), .B2(n17302), .A(n17244), .ZN(P3_U2769) );
  AOI22_X1 U20494 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17294), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n17293), .ZN(n17246) );
  OAI21_X1 U20495 ( .B1(n17247), .B2(n17302), .A(n17246), .ZN(P3_U2770) );
  AOI22_X1 U20496 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n9758), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n17293), .ZN(n17248) );
  OAI21_X1 U20497 ( .B1(n17249), .B2(n17302), .A(n17248), .ZN(P3_U2771) );
  AOI22_X1 U20498 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n9758), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n17293), .ZN(n17250) );
  OAI21_X1 U20499 ( .B1(n17251), .B2(n17302), .A(n17250), .ZN(P3_U2772) );
  AOI22_X1 U20500 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n9758), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n17293), .ZN(n17252) );
  OAI21_X1 U20501 ( .B1(n17253), .B2(n17302), .A(n17252), .ZN(P3_U2773) );
  AOI22_X1 U20502 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n9758), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n17293), .ZN(n17254) );
  OAI21_X1 U20503 ( .B1(n17255), .B2(n17302), .A(n17254), .ZN(P3_U2774) );
  AOI22_X1 U20504 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n9758), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n17293), .ZN(n17256) );
  OAI21_X1 U20505 ( .B1(n17257), .B2(n17302), .A(n17256), .ZN(P3_U2775) );
  AOI22_X1 U20506 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n9758), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n17293), .ZN(n17258) );
  OAI21_X1 U20507 ( .B1(n17259), .B2(n17302), .A(n17258), .ZN(P3_U2776) );
  AOI22_X1 U20508 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n9758), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n17293), .ZN(n17260) );
  OAI21_X1 U20509 ( .B1(n17261), .B2(n17302), .A(n17260), .ZN(P3_U2777) );
  AOI22_X1 U20510 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n9758), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n17293), .ZN(n17262) );
  OAI21_X1 U20511 ( .B1(n20918), .B2(n17302), .A(n17262), .ZN(P3_U2778) );
  AOI22_X1 U20512 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n9758), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n17293), .ZN(n17263) );
  OAI21_X1 U20513 ( .B1(n17264), .B2(n17302), .A(n17263), .ZN(P3_U2779) );
  AOI22_X1 U20514 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17294), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n17293), .ZN(n17265) );
  OAI21_X1 U20515 ( .B1(n17266), .B2(n17302), .A(n17265), .ZN(P3_U2780) );
  AOI22_X1 U20516 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17294), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n17293), .ZN(n17267) );
  OAI21_X1 U20517 ( .B1(n17268), .B2(n17302), .A(n17267), .ZN(P3_U2781) );
  AOI22_X1 U20518 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17294), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n17293), .ZN(n17269) );
  OAI21_X1 U20519 ( .B1(n17270), .B2(n17302), .A(n17269), .ZN(P3_U2782) );
  AOI22_X1 U20520 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17294), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n17293), .ZN(n17271) );
  OAI21_X1 U20521 ( .B1(n17272), .B2(n17302), .A(n17271), .ZN(P3_U2783) );
  AOI22_X1 U20522 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17294), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n17293), .ZN(n17273) );
  OAI21_X1 U20523 ( .B1(n17274), .B2(n17302), .A(n17273), .ZN(P3_U2784) );
  AOI22_X1 U20524 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17294), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n17293), .ZN(n17275) );
  OAI21_X1 U20525 ( .B1(n17276), .B2(n17302), .A(n17275), .ZN(P3_U2785) );
  AOI22_X1 U20526 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17294), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n17293), .ZN(n17277) );
  OAI21_X1 U20527 ( .B1(n17278), .B2(n17302), .A(n17277), .ZN(P3_U2786) );
  AOI22_X1 U20528 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17294), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n17300), .ZN(n17279) );
  OAI21_X1 U20529 ( .B1(n17280), .B2(n17302), .A(n17279), .ZN(P3_U2787) );
  AOI22_X1 U20530 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17294), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n17300), .ZN(n17281) );
  OAI21_X1 U20531 ( .B1(n17282), .B2(n17302), .A(n17281), .ZN(P3_U2788) );
  AOI22_X1 U20532 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17294), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n17300), .ZN(n17283) );
  OAI21_X1 U20533 ( .B1(n17284), .B2(n17302), .A(n17283), .ZN(P3_U2789) );
  AOI22_X1 U20534 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17294), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n17300), .ZN(n17285) );
  OAI21_X1 U20535 ( .B1(n20896), .B2(n17302), .A(n17285), .ZN(P3_U2790) );
  AOI22_X1 U20536 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17294), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n17300), .ZN(n17286) );
  OAI21_X1 U20537 ( .B1(n20741), .B2(n17302), .A(n17286), .ZN(P3_U2791) );
  AOI22_X1 U20538 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17294), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n17300), .ZN(n17287) );
  OAI21_X1 U20539 ( .B1(n17288), .B2(n17302), .A(n17287), .ZN(P3_U2792) );
  AOI22_X1 U20540 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n9758), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n17293), .ZN(n17289) );
  OAI21_X1 U20541 ( .B1(n17290), .B2(n17302), .A(n17289), .ZN(P3_U2793) );
  AOI22_X1 U20542 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17294), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n17300), .ZN(n17291) );
  OAI21_X1 U20543 ( .B1(n17292), .B2(n17302), .A(n17291), .ZN(P3_U2794) );
  AOI22_X1 U20544 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n9758), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n17293), .ZN(n17295) );
  OAI21_X1 U20545 ( .B1(n20936), .B2(n17302), .A(n17295), .ZN(P3_U2795) );
  AOI22_X1 U20546 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17294), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n17300), .ZN(n17296) );
  OAI21_X1 U20547 ( .B1(n17297), .B2(n17302), .A(n17296), .ZN(P3_U2796) );
  AOI22_X1 U20548 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17294), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n17300), .ZN(n17298) );
  OAI21_X1 U20549 ( .B1(n17299), .B2(n17302), .A(n17298), .ZN(P3_U2797) );
  AOI22_X1 U20550 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n17294), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n17300), .ZN(n17301) );
  OAI21_X1 U20551 ( .B1(n17303), .B2(n17302), .A(n17301), .ZN(P3_U2798) );
  AOI21_X1 U20552 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n17333), .A(
        n18514), .ZN(n17304) );
  AOI211_X1 U20553 ( .C1(n17629), .C2(n17313), .A(n17646), .B(n17304), .ZN(
        n17338) );
  OAI21_X1 U20554 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n17424), .A(
        n17338), .ZN(n17319) );
  AOI22_X1 U20555 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n17319), .B1(
        n17470), .B2(n17305), .ZN(n17318) );
  NOR2_X1 U20556 ( .A1(n17667), .A2(n17587), .ZN(n17417) );
  INV_X1 U20557 ( .A(n17587), .ZN(n17540) );
  OAI22_X1 U20558 ( .A1(n17690), .A2(n17678), .B1(n17686), .B2(n17540), .ZN(
        n17340) );
  NOR2_X1 U20559 ( .A1(n20733), .A2(n17340), .ZN(n17324) );
  NOR3_X1 U20560 ( .A1(n17417), .A2(n17324), .A3(n17306), .ZN(n17311) );
  AOI211_X1 U20561 ( .C1(n17309), .C2(n17308), .A(n17307), .B(n17493), .ZN(
        n17310) );
  AOI211_X1 U20562 ( .C1(n17460), .C2(n17312), .A(n17311), .B(n17310), .ZN(
        n17317) );
  NAND2_X1 U20563 ( .A1(n17995), .A2(P3_REIP_REG_28__SCAN_IN), .ZN(n17316) );
  NOR2_X1 U20564 ( .A1(n17471), .A2(n17313), .ZN(n17327) );
  OAI211_X1 U20565 ( .C1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A(n17327), .B(n17314), .ZN(n17315) );
  NAND4_X1 U20566 ( .A1(n17318), .A2(n17317), .A3(n17316), .A4(n17315), .ZN(
        P3_U2802) );
  AOI22_X1 U20567 ( .A1(n17979), .A2(P3_REIP_REG_27__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n17319), .ZN(n17329) );
  INV_X1 U20568 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n17326) );
  AOI21_X1 U20569 ( .B1(n17320), .B2(n17382), .A(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n17323) );
  NAND2_X1 U20570 ( .A1(n9893), .A2(n17321), .ZN(n17322) );
  XNOR2_X1 U20571 ( .A(n17585), .B(n17322), .ZN(n17694) );
  OAI22_X1 U20572 ( .A1(n17324), .A2(n17323), .B1(n17694), .B2(n17493), .ZN(
        n17325) );
  AOI21_X1 U20573 ( .B1(n17327), .B2(n17326), .A(n17325), .ZN(n17328) );
  OAI211_X1 U20574 ( .C1(n17521), .C2(n17330), .A(n17329), .B(n17328), .ZN(
        P3_U2803) );
  AOI21_X1 U20575 ( .B1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n17332), .A(
        n17331), .ZN(n17700) );
  AOI21_X1 U20576 ( .B1(n17333), .B2(n18390), .A(
        P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n17337) );
  OAI21_X1 U20577 ( .B1(n17470), .B2(n17390), .A(n17334), .ZN(n17336) );
  NAND2_X1 U20578 ( .A1(n17995), .A2(P3_REIP_REG_26__SCAN_IN), .ZN(n17335) );
  OAI211_X1 U20579 ( .C1(n17338), .C2(n17337), .A(n17336), .B(n17335), .ZN(
        n17339) );
  AOI21_X1 U20580 ( .B1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n17340), .A(
        n17339), .ZN(n17342) );
  INV_X1 U20581 ( .A(n17682), .ZN(n17701) );
  NAND4_X1 U20582 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n17701), .A3(
        n17382), .A4(n20821), .ZN(n17341) );
  OAI211_X1 U20583 ( .C1(n17700), .C2(n17493), .A(n17342), .B(n17341), .ZN(
        P3_U2804) );
  AND2_X1 U20584 ( .A1(n17352), .A2(n18390), .ZN(n17375) );
  AOI211_X1 U20585 ( .C1(n17387), .C2(n17343), .A(n17646), .B(n17375), .ZN(
        n17379) );
  OAI21_X1 U20586 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n17424), .A(
        n17379), .ZN(n17362) );
  AOI22_X1 U20587 ( .A1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n17362), .B1(
        n17470), .B2(n17344), .ZN(n17356) );
  XNOR2_X1 U20588 ( .A(n17345), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n17711) );
  OAI21_X1 U20589 ( .B1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n17347), .A(
        n17346), .ZN(n17709) );
  OAI21_X1 U20590 ( .B1(n17551), .B2(n17349), .A(n17348), .ZN(n17350) );
  XNOR2_X1 U20591 ( .A(n17350), .B(n17704), .ZN(n17713) );
  OAI22_X1 U20592 ( .A1(n17678), .A2(n17709), .B1(n17493), .B2(n17713), .ZN(
        n17351) );
  AOI21_X1 U20593 ( .B1(n17587), .B2(n17711), .A(n17351), .ZN(n17355) );
  NAND2_X1 U20594 ( .A1(n17995), .A2(P3_REIP_REG_25__SCAN_IN), .ZN(n17707) );
  NOR2_X1 U20595 ( .A1(n17471), .A2(n17352), .ZN(n17364) );
  OAI211_X1 U20596 ( .C1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A(n17364), .B(n17353), .ZN(n17354) );
  NAND4_X1 U20597 ( .A1(n17356), .A2(n17355), .A3(n17707), .A4(n17354), .ZN(
        P3_U2805) );
  AOI21_X1 U20598 ( .B1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n17358), .A(
        n17357), .ZN(n17725) );
  AOI22_X1 U20599 ( .A1(n17979), .A2(P3_REIP_REG_24__SCAN_IN), .B1(n17470), 
        .B2(n17359), .ZN(n17360) );
  INV_X1 U20600 ( .A(n17360), .ZN(n17361) );
  AOI221_X1 U20601 ( .B1(n17364), .B2(n17363), .C1(n17362), .C2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A(n17361), .ZN(n17369) );
  AOI22_X1 U20602 ( .A1(n17716), .A2(n17667), .B1(n17715), .B2(n17587), .ZN(
        n17365) );
  INV_X1 U20603 ( .A(n17365), .ZN(n17381) );
  AND2_X1 U20604 ( .A1(n17367), .A2(n17366), .ZN(n17714) );
  AOI22_X1 U20605 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17381), .B1(
        n17460), .B2(n17714), .ZN(n17368) );
  OAI211_X1 U20606 ( .C1(n17725), .C2(n17493), .A(n17369), .B(n17368), .ZN(
        P3_U2806) );
  AOI22_X1 U20607 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n17551), .B1(
        n17370), .B2(n17398), .ZN(n17371) );
  NAND2_X1 U20608 ( .A1(n17419), .A2(n17371), .ZN(n17372) );
  XNOR2_X1 U20609 ( .A(n17372), .B(n17719), .ZN(n17730) );
  INV_X1 U20610 ( .A(n17659), .ZN(n17373) );
  AOI22_X1 U20611 ( .A1(n17376), .A2(n17375), .B1(n17374), .B2(n17373), .ZN(
        n17377) );
  NAND2_X1 U20612 ( .A1(n17979), .A2(P3_REIP_REG_23__SCAN_IN), .ZN(n17729) );
  OAI211_X1 U20613 ( .C1(n17379), .C2(n17378), .A(n17377), .B(n17729), .ZN(
        n17380) );
  AOI221_X1 U20614 ( .B1(n17382), .B2(n17719), .C1(n17381), .C2(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A(n17380), .ZN(n17383) );
  OAI21_X1 U20615 ( .B1(n17493), .B2(n17730), .A(n17383), .ZN(P3_U2807) );
  OR2_X1 U20616 ( .A1(n17385), .A2(n17471), .ZN(n17410) );
  AOI211_X1 U20617 ( .C1(n17409), .C2(n17391), .A(n17384), .B(n17410), .ZN(
        n17393) );
  AOI22_X1 U20618 ( .A1(n17387), .A2(n17386), .B1(n17629), .B2(n17385), .ZN(
        n17388) );
  NAND2_X1 U20619 ( .A1(n17388), .A2(n17674), .ZN(n17422) );
  AOI21_X1 U20620 ( .B1(n17390), .B2(n17389), .A(n17422), .ZN(n17408) );
  NAND2_X1 U20621 ( .A1(n17979), .A2(P3_REIP_REG_22__SCAN_IN), .ZN(n17746) );
  OAI21_X1 U20622 ( .B1(n17408), .B2(n17391), .A(n17746), .ZN(n17392) );
  AOI211_X1 U20623 ( .C1(n17394), .C2(n17470), .A(n17393), .B(n17392), .ZN(
        n17402) );
  NOR2_X1 U20624 ( .A1(n17808), .A2(n17540), .ZN(n17490) );
  INV_X1 U20625 ( .A(n17490), .ZN(n17395) );
  OAI21_X1 U20626 ( .B1(n17678), .B2(n17807), .A(n17395), .ZN(n17441) );
  INV_X1 U20627 ( .A(n17441), .ZN(n17478) );
  OAI21_X1 U20628 ( .B1(n17737), .B2(n17417), .A(n17478), .ZN(n17414) );
  INV_X1 U20629 ( .A(n17419), .ZN(n17396) );
  AOI221_X1 U20630 ( .B1(n17403), .B2(n17398), .C1(n17397), .C2(n17398), .A(
        n17396), .ZN(n17399) );
  XNOR2_X1 U20631 ( .A(n17399), .B(n20826), .ZN(n17744) );
  AOI22_X1 U20632 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n17414), .B1(
        n17586), .B2(n17744), .ZN(n17401) );
  NAND3_X1 U20633 ( .A1(n17737), .A2(n17460), .A3(n20826), .ZN(n17400) );
  NAND3_X1 U20634 ( .A1(n17402), .A2(n17401), .A3(n17400), .ZN(P3_U2808) );
  NOR3_X1 U20635 ( .A1(n17452), .A2(n17551), .A3(n17403), .ZN(n17435) );
  INV_X1 U20636 ( .A(n17448), .ZN(n17436) );
  AOI22_X1 U20637 ( .A1(n17753), .A2(n17435), .B1(n17436), .B2(n17404), .ZN(
        n17406) );
  XNOR2_X1 U20638 ( .A(n17406), .B(n17405), .ZN(n17757) );
  NAND2_X1 U20639 ( .A1(n17995), .A2(P3_REIP_REG_21__SCAN_IN), .ZN(n17407) );
  OAI221_X1 U20640 ( .B1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n17410), .C1(
        n17409), .C2(n17408), .A(n17407), .ZN(n17411) );
  AOI21_X1 U20641 ( .B1(n17470), .B2(n17412), .A(n17411), .ZN(n17416) );
  NOR3_X1 U20642 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17736), .A3(
        n17413), .ZN(n17748) );
  AOI22_X1 U20643 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17414), .B1(
        n17460), .B2(n17748), .ZN(n17415) );
  OAI211_X1 U20644 ( .C1(n17757), .C2(n17493), .A(n17416), .B(n17415), .ZN(
        P3_U2809) );
  NOR2_X1 U20645 ( .A1(n17736), .A2(n17773), .ZN(n17759) );
  AND2_X1 U20646 ( .A1(n17739), .A2(n17759), .ZN(n17763) );
  OAI21_X1 U20647 ( .B1(n17417), .B2(n17759), .A(n17478), .ZN(n17418) );
  INV_X1 U20648 ( .A(n17418), .ZN(n17440) );
  OAI221_X1 U20649 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n17447), 
        .C1(n17773), .C2(n17435), .A(n17419), .ZN(n17420) );
  XNOR2_X1 U20650 ( .A(n17739), .B(n17420), .ZN(n17767) );
  OAI22_X1 U20651 ( .A1(n17440), .A2(n17739), .B1(n17493), .B2(n17767), .ZN(
        n17421) );
  AOI21_X1 U20652 ( .B1(n17460), .B2(n17763), .A(n17421), .ZN(n17428) );
  NAND2_X1 U20653 ( .A1(n17995), .A2(P3_REIP_REG_20__SCAN_IN), .ZN(n17765) );
  OAI221_X1 U20654 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n17423), .C1(
        P3_PHYADDRPOINTER_REG_20__SCAN_IN), .C2(n18390), .A(n17422), .ZN(
        n17427) );
  OAI21_X1 U20655 ( .B1(n17470), .B2(n17390), .A(n17425), .ZN(n17426) );
  NAND4_X1 U20656 ( .A1(n17428), .A2(n17765), .A3(n17427), .A4(n17426), .ZN(
        P3_U2810) );
  AOI21_X1 U20657 ( .B1(n17629), .B2(n17430), .A(n17646), .ZN(n17455) );
  OAI21_X1 U20658 ( .B1(n17429), .B2(n18514), .A(n17455), .ZN(n17444) );
  NOR2_X1 U20659 ( .A1(n17471), .A2(n17430), .ZN(n17446) );
  OAI211_X1 U20660 ( .C1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(n17446), .B(n17431), .ZN(n17432) );
  NAND2_X1 U20661 ( .A1(n17995), .A2(P3_REIP_REG_19__SCAN_IN), .ZN(n17771) );
  OAI211_X1 U20662 ( .C1(n17521), .C2(n17433), .A(n17432), .B(n17771), .ZN(
        n17434) );
  AOI21_X1 U20663 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n17444), .A(
        n17434), .ZN(n17439) );
  AOI21_X1 U20664 ( .B1(n17447), .B2(n17436), .A(n17435), .ZN(n17437) );
  XNOR2_X1 U20665 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B(n17437), .ZN(
        n17770) );
  NOR2_X1 U20666 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17736), .ZN(
        n17768) );
  AOI22_X1 U20667 ( .A1(n17586), .A2(n17770), .B1(n17460), .B2(n17768), .ZN(
        n17438) );
  OAI211_X1 U20668 ( .C1(n17440), .C2(n17773), .A(n17439), .B(n17438), .ZN(
        P3_U2811) );
  AOI21_X1 U20669 ( .B1(n17460), .B2(n17778), .A(n17441), .ZN(n17463) );
  OAI22_X1 U20670 ( .A1(n17993), .A2(n18559), .B1(n17521), .B2(n17442), .ZN(
        n17443) );
  AOI221_X1 U20671 ( .B1(n17446), .B2(n17445), .C1(n17444), .C2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(n17443), .ZN(n17451) );
  AOI21_X1 U20672 ( .B1(n17585), .B2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n17447), .ZN(n17449) );
  XNOR2_X1 U20673 ( .A(n17449), .B(n17448), .ZN(n17788) );
  NOR2_X1 U20674 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17778), .ZN(
        n17787) );
  AOI22_X1 U20675 ( .A1(n17586), .A2(n17788), .B1(n17460), .B2(n17787), .ZN(
        n17450) );
  OAI211_X1 U20676 ( .C1(n17463), .C2(n17452), .A(n17451), .B(n17450), .ZN(
        P3_U2812) );
  AOI21_X1 U20677 ( .B1(n18390), .B2(n17453), .A(
        P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n17456) );
  OAI22_X1 U20678 ( .A1(n17456), .A2(n17455), .B1(n17659), .B2(n17454), .ZN(
        n17457) );
  AOI21_X1 U20679 ( .B1(n17995), .B2(P3_REIP_REG_17__SCAN_IN), .A(n17457), 
        .ZN(n17462) );
  OAI21_X1 U20680 ( .B1(n17459), .B2(n17782), .A(n17458), .ZN(n17793) );
  NOR2_X1 U20681 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n17802), .ZN(
        n17792) );
  AOI22_X1 U20682 ( .A1(n17586), .A2(n17793), .B1(n17460), .B2(n17792), .ZN(
        n17461) );
  OAI211_X1 U20683 ( .C1(n17463), .C2(n17782), .A(n17462), .B(n17461), .ZN(
        P3_U2813) );
  AOI21_X1 U20684 ( .B1(n17585), .B2(n17465), .A(n17464), .ZN(n17466) );
  XNOR2_X1 U20685 ( .A(n17466), .B(n17802), .ZN(n17804) );
  AOI21_X1 U20686 ( .B1(n17629), .B2(n17467), .A(n17646), .ZN(n17497) );
  OAI21_X1 U20687 ( .B1(n17468), .B2(n18514), .A(n17497), .ZN(n17486) );
  AOI22_X1 U20688 ( .A1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n17486), .B1(
        n17470), .B2(n17469), .ZN(n17475) );
  OR2_X1 U20689 ( .A1(n17506), .A2(n17471), .ZN(n17523) );
  NOR2_X1 U20690 ( .A1(n17472), .A2(n17523), .ZN(n17488) );
  OAI211_X1 U20691 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(n17488), .B(n17473), .ZN(n17474) );
  OAI211_X1 U20692 ( .C1(n18555), .C2(n17993), .A(n17475), .B(n17474), .ZN(
        n17476) );
  AOI21_X1 U20693 ( .B1(n17586), .B2(n17804), .A(n17476), .ZN(n17477) );
  OAI221_X1 U20694 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n17479), 
        .C1(n17802), .C2(n17478), .A(n17477), .ZN(P3_U2814) );
  NOR3_X1 U20695 ( .A1(n17831), .A2(n17858), .A3(n17480), .ZN(n17481) );
  NAND2_X1 U20696 ( .A1(n17552), .A2(n17551), .ZN(n17563) );
  NOR3_X1 U20697 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n17558), .A3(
        n17563), .ZN(n17526) );
  AOI22_X1 U20698 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n17481), .B1(
        n17526), .B2(n17517), .ZN(n17482) );
  AOI221_X1 U20699 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n17864), 
        .C1(n17551), .C2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A(n17482), .ZN(
        n17483) );
  XNOR2_X1 U20700 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B(n17483), .ZN(
        n17814) );
  INV_X1 U20701 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n17487) );
  OAI22_X1 U20702 ( .A1(n17993), .A2(n18553), .B1(n17521), .B2(n17484), .ZN(
        n17485) );
  AOI221_X1 U20703 ( .B1(n17488), .B2(n17487), .C1(n17486), .C2(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A(n17485), .ZN(n17492) );
  NAND2_X1 U20704 ( .A1(n17822), .A2(n17501), .ZN(n17812) );
  NOR2_X1 U20705 ( .A1(n17807), .A2(n17678), .ZN(n17489) );
  NAND2_X1 U20706 ( .A1(n17494), .A2(n17822), .ZN(n17818) );
  AOI22_X1 U20707 ( .A1(n17490), .A2(n17812), .B1(n17489), .B2(n17818), .ZN(
        n17491) );
  OAI211_X1 U20708 ( .C1(n17493), .C2(n17814), .A(n17492), .B(n17491), .ZN(
        P3_U2815) );
  OAI21_X1 U20709 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n17495), .A(
        n17494), .ZN(n17839) );
  NAND2_X1 U20710 ( .A1(n18390), .A2(n17496), .ZN(n17536) );
  AOI221_X1 U20711 ( .B1(n17509), .B2(n17498), .C1(n17536), .C2(n17498), .A(
        n17497), .ZN(n17499) );
  NOR2_X1 U20712 ( .A1(n17993), .A2(n18552), .ZN(n17832) );
  AOI211_X1 U20713 ( .C1(n17500), .C2(n17373), .A(n17499), .B(n17832), .ZN(
        n17505) );
  INV_X1 U20714 ( .A(n17829), .ZN(n17824) );
  OAI221_X1 U20715 ( .B1(n17874), .B2(P3_INSTADDRPOINTER_REG_14__SCAN_IN), 
        .C1(n17824), .C2(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A(n17501), .ZN(
        n17502) );
  INV_X1 U20716 ( .A(n17502), .ZN(n17836) );
  NAND2_X1 U20717 ( .A1(n17585), .A2(n17874), .ZN(n17564) );
  INV_X1 U20718 ( .A(n17564), .ZN(n17555) );
  NAND2_X1 U20719 ( .A1(n17854), .A2(n17555), .ZN(n17515) );
  NAND2_X1 U20720 ( .A1(n17526), .A2(n17864), .ZN(n17516) );
  AOI22_X1 U20721 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n17515), .B1(
        n17516), .B2(n17517), .ZN(n17503) );
  XNOR2_X1 U20722 ( .A(n17831), .B(n17503), .ZN(n17835) );
  AOI22_X1 U20723 ( .A1(n17587), .A2(n17836), .B1(n17586), .B2(n17835), .ZN(
        n17504) );
  OAI211_X1 U20724 ( .C1(n17678), .C2(n17839), .A(n17505), .B(n17504), .ZN(
        P3_U2816) );
  NAND2_X1 U20725 ( .A1(n17854), .A2(n17517), .ZN(n17853) );
  AOI21_X1 U20726 ( .B1(n17629), .B2(n17506), .A(n17646), .ZN(n17507) );
  OAI21_X1 U20727 ( .B1(n17508), .B2(n18514), .A(n17507), .ZN(n17525) );
  NOR2_X1 U20728 ( .A1(n17993), .A2(n18549), .ZN(n17513) );
  OAI21_X1 U20729 ( .B1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A(n17509), .ZN(n17510) );
  OAI22_X1 U20730 ( .A1(n17521), .A2(n17511), .B1(n17523), .B2(n17510), .ZN(
        n17512) );
  AOI211_X1 U20731 ( .C1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .C2(n17525), .A(
        n17513), .B(n17512), .ZN(n17520) );
  INV_X1 U20732 ( .A(n17848), .ZN(n17514) );
  AND2_X1 U20733 ( .A1(n17854), .A2(n17874), .ZN(n17846) );
  OAI22_X1 U20734 ( .A1(n17514), .A2(n17678), .B1(n17846), .B2(n17540), .ZN(
        n17529) );
  NAND2_X1 U20735 ( .A1(n17516), .A2(n17515), .ZN(n17518) );
  XNOR2_X1 U20736 ( .A(n17518), .B(n17517), .ZN(n17841) );
  AOI22_X1 U20737 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n17529), .B1(
        n17586), .B2(n17841), .ZN(n17519) );
  OAI211_X1 U20738 ( .C1(n17574), .C2(n17853), .A(n17520), .B(n17519), .ZN(
        P3_U2817) );
  OAI22_X1 U20739 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n17523), .B1(
        n17522), .B2(n17521), .ZN(n17524) );
  AOI21_X1 U20740 ( .B1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n17525), .A(
        n17524), .ZN(n17532) );
  INV_X1 U20741 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n17842) );
  NAND2_X1 U20742 ( .A1(n17844), .A2(n17555), .ZN(n17553) );
  INV_X1 U20743 ( .A(n17526), .ZN(n17527) );
  OAI21_X1 U20744 ( .B1(n17842), .B2(n17553), .A(n17527), .ZN(n17528) );
  XNOR2_X1 U20745 ( .A(n17528), .B(n17864), .ZN(n17861) );
  AOI22_X1 U20746 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n17529), .B1(
        n17586), .B2(n17861), .ZN(n17531) );
  NAND2_X1 U20747 ( .A1(n17995), .A2(P3_REIP_REG_12__SCAN_IN), .ZN(n17862) );
  OR3_X1 U20748 ( .A1(n17858), .A2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A3(
        n17574), .ZN(n17530) );
  NAND4_X1 U20749 ( .A1(n17532), .A2(n17531), .A3(n17862), .A4(n17530), .ZN(
        P3_U2818) );
  NOR2_X1 U20750 ( .A1(n18057), .A2(n17533), .ZN(n17606) );
  NAND2_X1 U20751 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n17606), .ZN(
        n17591) );
  OAI22_X1 U20752 ( .A1(n17671), .A2(n17534), .B1(n17544), .B2(n17591), .ZN(
        n17535) );
  AOI22_X1 U20753 ( .A1(n17537), .A2(n17373), .B1(n17536), .B2(n17535), .ZN(
        n17543) );
  OAI21_X1 U20754 ( .B1(n17563), .B2(n17558), .A(n17553), .ZN(n17538) );
  XOR2_X1 U20755 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n17538), .Z(
        n17867) );
  NOR2_X1 U20756 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n17875), .ZN(
        n17866) );
  INV_X1 U20757 ( .A(n17574), .ZN(n17539) );
  AOI22_X1 U20758 ( .A1(n17586), .A2(n17867), .B1(n17866), .B2(n17539), .ZN(
        n17542) );
  NOR2_X1 U20759 ( .A1(n17844), .A2(n17574), .ZN(n17559) );
  OAI22_X1 U20760 ( .A1(n17874), .A2(n17540), .B1(n17678), .B2(n17868), .ZN(
        n17562) );
  OAI21_X1 U20761 ( .B1(n17559), .B2(n17562), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n17541) );
  NAND2_X1 U20762 ( .A1(n17995), .A2(P3_REIP_REG_11__SCAN_IN), .ZN(n17881) );
  NAND4_X1 U20763 ( .A1(n17543), .A2(n17542), .A3(n17541), .A4(n17881), .ZN(
        P3_U2819) );
  NOR2_X1 U20764 ( .A1(n17993), .A2(n18544), .ZN(n17550) );
  NOR2_X1 U20765 ( .A1(n17544), .A2(n17591), .ZN(n17548) );
  NAND2_X1 U20766 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n17578) );
  NOR3_X1 U20767 ( .A1(n17578), .A2(n17545), .A3(n17591), .ZN(n17570) );
  AOI21_X1 U20768 ( .B1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n17567), .A(
        n17570), .ZN(n17547) );
  OAI22_X1 U20769 ( .A1(n17548), .A2(n17547), .B1(n17659), .B2(n17546), .ZN(
        n17549) );
  AOI211_X1 U20770 ( .C1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .C2(n17562), .A(
        n17550), .B(n17549), .ZN(n17561) );
  INV_X1 U20771 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n17892) );
  OR2_X1 U20772 ( .A1(n17892), .A2(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n17891) );
  NAND4_X1 U20773 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n17552), .A3(
        n17892), .A4(n17551), .ZN(n17554) );
  OAI211_X1 U20774 ( .C1(n17555), .C2(n17891), .A(n17554), .B(n17553), .ZN(
        n17556) );
  AOI21_X1 U20775 ( .B1(n17557), .B2(n17563), .A(n17556), .ZN(n17883) );
  AOI22_X1 U20776 ( .A1(n17586), .A2(n17883), .B1(n17559), .B2(n17558), .ZN(
        n17560) );
  NAND2_X1 U20777 ( .A1(n17561), .A2(n17560), .ZN(P3_U2820) );
  INV_X1 U20778 ( .A(n17562), .ZN(n17573) );
  NAND2_X1 U20779 ( .A1(n17564), .A2(n17563), .ZN(n17565) );
  XNOR2_X1 U20780 ( .A(n17565), .B(n17892), .ZN(n17896) );
  NOR2_X1 U20781 ( .A1(n17993), .A2(n18543), .ZN(n17895) );
  NOR2_X1 U20782 ( .A1(n17578), .A2(n17591), .ZN(n17566) );
  AOI21_X1 U20783 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n17567), .A(
        n17566), .ZN(n17569) );
  OAI22_X1 U20784 ( .A1(n17570), .A2(n17569), .B1(n17659), .B2(n17568), .ZN(
        n17571) );
  AOI211_X1 U20785 ( .C1(n17586), .C2(n17896), .A(n17895), .B(n17571), .ZN(
        n17572) );
  OAI221_X1 U20786 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n17574), .C1(
        n17892), .C2(n17573), .A(n17572), .ZN(P3_U2821) );
  OAI21_X1 U20787 ( .B1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n17576), .A(
        n17575), .ZN(n17915) );
  AOI21_X1 U20788 ( .B1(n17629), .B2(n17577), .A(n17646), .ZN(n17592) );
  OAI211_X1 U20789 ( .C1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .C2(n17579), .A(
        n18390), .B(n17578), .ZN(n17580) );
  NAND2_X1 U20790 ( .A1(n17979), .A2(P3_REIP_REG_8__SCAN_IN), .ZN(n17904) );
  OAI211_X1 U20791 ( .C1(n17592), .C2(n17581), .A(n17580), .B(n17904), .ZN(
        n17582) );
  AOI21_X1 U20792 ( .B1(n17583), .B2(n17373), .A(n17582), .ZN(n17589) );
  OAI21_X1 U20793 ( .B1(n17585), .B2(n17912), .A(n17584), .ZN(n17909) );
  AOI22_X1 U20794 ( .A1(n17587), .A2(n17912), .B1(n17586), .B2(n17909), .ZN(
        n17588) );
  OAI211_X1 U20795 ( .C1(n17678), .C2(n17915), .A(n17589), .B(n17588), .ZN(
        P3_U2822) );
  AOI22_X1 U20796 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n17592), .B1(
        n17591), .B2(n17590), .ZN(n17593) );
  AOI21_X1 U20797 ( .B1(n17979), .B2(P3_REIP_REG_7__SCAN_IN), .A(n17593), .ZN(
        n17601) );
  AOI21_X1 U20798 ( .B1(n17596), .B2(n17595), .A(n17594), .ZN(n17597) );
  XNOR2_X1 U20799 ( .A(n17597), .B(n17902), .ZN(n17921) );
  AOI21_X1 U20800 ( .B1(n17902), .B2(n17599), .A(n17598), .ZN(n17920) );
  AOI22_X1 U20801 ( .A1(n17667), .A2(n17921), .B1(n17664), .B2(n17920), .ZN(
        n17600) );
  OAI211_X1 U20802 ( .C1(n17659), .C2(n17602), .A(n17601), .B(n17600), .ZN(
        P3_U2823) );
  AOI21_X1 U20803 ( .B1(n17605), .B2(n17604), .A(n17603), .ZN(n17926) );
  AOI22_X1 U20804 ( .A1(n17664), .A2(n17926), .B1(n17606), .B2(n20957), .ZN(
        n17612) );
  NOR2_X1 U20805 ( .A1(n17671), .A2(n17606), .ZN(n17624) );
  OAI21_X1 U20806 ( .B1(n17608), .B2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n17607), .ZN(n17934) );
  OAI22_X1 U20807 ( .A1(n17659), .A2(n17609), .B1(n17678), .B2(n17934), .ZN(
        n17610) );
  AOI21_X1 U20808 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n17624), .A(
        n17610), .ZN(n17611) );
  OAI211_X1 U20809 ( .C1(n17993), .C2(n18537), .A(n17612), .B(n17611), .ZN(
        P3_U2824) );
  OAI21_X1 U20810 ( .B1(n17615), .B2(n17614), .A(n17613), .ZN(n17941) );
  OAI21_X1 U20811 ( .B1(n17618), .B2(n17617), .A(n17616), .ZN(n17619) );
  XNOR2_X1 U20812 ( .A(n17619), .B(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n17935) );
  AOI22_X1 U20813 ( .A1(n17664), .A2(n17935), .B1(n17995), .B2(
        P3_REIP_REG_5__SCAN_IN), .ZN(n17626) );
  OAI21_X1 U20814 ( .B1(n17646), .B2(n17621), .A(n17620), .ZN(n17623) );
  AOI22_X1 U20815 ( .A1(n17624), .A2(n17623), .B1(n17622), .B2(n17373), .ZN(
        n17625) );
  OAI211_X1 U20816 ( .C1(n17678), .C2(n17941), .A(n17626), .B(n17625), .ZN(
        P3_U2825) );
  AOI21_X1 U20817 ( .B1(n9873), .B2(n17628), .A(n17627), .ZN(n17942) );
  AOI22_X1 U20818 ( .A1(n17664), .A2(n17942), .B1(n17995), .B2(
        P3_REIP_REG_4__SCAN_IN), .ZN(n17637) );
  INV_X1 U20819 ( .A(n17629), .ZN(n17630) );
  OAI21_X1 U20820 ( .B1(n17631), .B2(n17630), .A(n17674), .ZN(n17648) );
  OAI21_X1 U20821 ( .B1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n17633), .A(
        n17632), .ZN(n17953) );
  OAI22_X1 U20822 ( .A1(n17659), .A2(n17634), .B1(n17678), .B2(n17953), .ZN(
        n17635) );
  AOI21_X1 U20823 ( .B1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n17648), .A(
        n17635), .ZN(n17636) );
  OAI211_X1 U20824 ( .C1(n18057), .C2(n17638), .A(n17637), .B(n17636), .ZN(
        P3_U2826) );
  OAI21_X1 U20825 ( .B1(n17641), .B2(n17640), .A(n17639), .ZN(n17962) );
  AOI21_X1 U20826 ( .B1(n17644), .B2(n17643), .A(n17642), .ZN(n17960) );
  AOI22_X1 U20827 ( .A1(n17664), .A2(n17960), .B1(n17995), .B2(
        P3_REIP_REG_3__SCAN_IN), .ZN(n17651) );
  OAI21_X1 U20828 ( .B1(n17646), .B2(n17662), .A(n17645), .ZN(n17647) );
  AOI22_X1 U20829 ( .A1(n17649), .A2(n17373), .B1(n17648), .B2(n17647), .ZN(
        n17650) );
  OAI211_X1 U20830 ( .C1(n17678), .C2(n17962), .A(n17651), .B(n17650), .ZN(
        P3_U2827) );
  AOI21_X1 U20831 ( .B1(n17654), .B2(n17653), .A(n17652), .ZN(n17964) );
  INV_X1 U20832 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n20867) );
  NOR2_X1 U20833 ( .A1(n17993), .A2(n20867), .ZN(n17963) );
  OAI21_X1 U20834 ( .B1(n17657), .B2(n17656), .A(n17655), .ZN(n17971) );
  OAI22_X1 U20835 ( .A1(n17659), .A2(n17658), .B1(n17678), .B2(n17971), .ZN(
        n17660) );
  AOI211_X1 U20836 ( .C1(n17664), .C2(n17964), .A(n17963), .B(n17660), .ZN(
        n17661) );
  OAI221_X1 U20837 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n18057), .C1(
        n17662), .C2(n17674), .A(n17661), .ZN(P3_U2828) );
  AOI21_X1 U20838 ( .B1(n17665), .B2(n17672), .A(n17663), .ZN(n17978) );
  AOI22_X1 U20839 ( .A1(n17664), .A2(n17978), .B1(n17995), .B2(
        P3_REIP_REG_1__SCAN_IN), .ZN(n17669) );
  NOR2_X1 U20840 ( .A1(n17673), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n17666) );
  XNOR2_X1 U20841 ( .A(n17666), .B(n17665), .ZN(n17981) );
  AOI22_X1 U20842 ( .A1(n17667), .A2(n17981), .B1(n17670), .B2(n17373), .ZN(
        n17668) );
  OAI211_X1 U20843 ( .C1(n17671), .C2(n17670), .A(n17669), .B(n17668), .ZN(
        P3_U2829) );
  OAI21_X1 U20844 ( .B1(n17673), .B2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n17672), .ZN(n17998) );
  INV_X1 U20845 ( .A(n17998), .ZN(n18000) );
  NAND3_X1 U20846 ( .A1(n18610), .A2(n18514), .A3(n17674), .ZN(n17675) );
  AOI22_X1 U20847 ( .A1(n17995), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17675), .ZN(n17676) );
  OAI221_X1 U20848 ( .B1(n18000), .B2(n17678), .C1(n17998), .C2(n17677), .A(
        n17676), .ZN(P3_U2830) );
  NOR3_X1 U20849 ( .A1(n17741), .A2(n17740), .A3(n20826), .ZN(n17727) );
  NAND3_X1 U20850 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n17701), .A3(
        n17727), .ZN(n17695) );
  NOR2_X1 U20851 ( .A1(n20821), .A2(n17695), .ZN(n17691) );
  NAND2_X1 U20852 ( .A1(n18465), .A2(n18481), .ZN(n17826) );
  AOI22_X1 U20853 ( .A1(n18469), .A2(n17704), .B1(n17679), .B2(n17826), .ZN(
        n17689) );
  NOR2_X1 U20854 ( .A1(n18469), .A2(n17877), .ZN(n17944) );
  INV_X1 U20855 ( .A(n17944), .ZN(n17781) );
  INV_X1 U20856 ( .A(n17680), .ZN(n17681) );
  AOI211_X1 U20857 ( .C1(n17781), .C2(n20826), .A(n17732), .B(n17681), .ZN(
        n17718) );
  OAI21_X1 U20858 ( .B1(n17683), .B2(n17682), .A(n18449), .ZN(n17684) );
  OAI211_X1 U20859 ( .C1(n17701), .C2(n17944), .A(n17718), .B(n17684), .ZN(
        n17685) );
  INV_X1 U20860 ( .A(n17685), .ZN(n17705) );
  OAI21_X1 U20861 ( .B1(n17873), .B2(n17686), .A(n17705), .ZN(n17687) );
  INV_X1 U20862 ( .A(n17687), .ZN(n17688) );
  OAI211_X1 U20863 ( .C1(n17690), .C2(n17972), .A(n17689), .B(n17688), .ZN(
        n17696) );
  NAND2_X1 U20864 ( .A1(n17995), .A2(P3_REIP_REG_27__SCAN_IN), .ZN(n17692) );
  OAI211_X1 U20865 ( .C1(n17694), .C2(n17815), .A(n17693), .B(n17692), .ZN(
        P3_U2835) );
  AOI22_X1 U20866 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n17918), .B1(
        n17995), .B2(P3_REIP_REG_26__SCAN_IN), .ZN(n17699) );
  INV_X1 U20867 ( .A(n17695), .ZN(n17697) );
  OAI221_X1 U20868 ( .B1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n17697), 
        .C1(n20821), .C2(n17696), .A(n17989), .ZN(n17698) );
  OAI211_X1 U20869 ( .C1(n17700), .C2(n17815), .A(n17699), .B(n17698), .ZN(
        P3_U2836) );
  NAND3_X1 U20870 ( .A1(n17702), .A2(n17701), .A3(n17704), .ZN(n17703) );
  OAI21_X1 U20871 ( .B1(n17705), .B2(n17704), .A(n17703), .ZN(n17706) );
  AOI22_X1 U20872 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n17918), .B1(
        n17989), .B2(n17706), .ZN(n17708) );
  OAI211_X1 U20873 ( .C1(n17709), .C2(n17999), .A(n17708), .B(n17707), .ZN(
        n17710) );
  AOI21_X1 U20874 ( .B1(n17911), .B2(n17711), .A(n17710), .ZN(n17712) );
  OAI21_X1 U20875 ( .B1(n17815), .B2(n17713), .A(n17712), .ZN(P3_U2837) );
  AOI22_X1 U20876 ( .A1(n17979), .A2(P3_REIP_REG_24__SCAN_IN), .B1(n17769), 
        .B2(n17714), .ZN(n17724) );
  AOI22_X1 U20877 ( .A1(n18447), .A2(n17716), .B1(n17733), .B2(n17715), .ZN(
        n17717) );
  NAND3_X1 U20878 ( .A1(n17718), .A2(n17717), .A3(n17980), .ZN(n17722) );
  NOR2_X1 U20879 ( .A1(n17719), .A2(n17722), .ZN(n17721) );
  AOI21_X1 U20880 ( .B1(n17721), .B2(n17720), .A(n17979), .ZN(n17726) );
  OAI211_X1 U20881 ( .C1(n17903), .C2(n17722), .A(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B(n17726), .ZN(n17723) );
  OAI211_X1 U20882 ( .C1(n17725), .C2(n17815), .A(n17724), .B(n17723), .ZN(
        P3_U2838) );
  OAI221_X1 U20883 ( .B1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n17727), 
        .C1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n17980), .A(n17726), .ZN(
        n17728) );
  OAI211_X1 U20884 ( .C1(n17815), .C2(n17730), .A(n17729), .B(n17728), .ZN(
        P3_U2839) );
  OAI22_X1 U20885 ( .A1(n17807), .A2(n17972), .B1(n17808), .B2(n17873), .ZN(
        n17749) );
  OAI22_X1 U20886 ( .A1(n17887), .A2(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .B1(
        n17753), .B2(n18481), .ZN(n17731) );
  NOR4_X1 U20887 ( .A1(n17732), .A2(n20826), .A3(n17749), .A4(n17731), .ZN(
        n17743) );
  NOR2_X1 U20888 ( .A1(n18447), .A2(n17733), .ZN(n17775) );
  INV_X1 U20889 ( .A(n18469), .ZN(n17990) );
  AOI21_X1 U20890 ( .B1(n17776), .B2(n17759), .A(n17990), .ZN(n17734) );
  AOI221_X1 U20891 ( .B1(n17736), .B2(n18449), .C1(n17735), .C2(n18449), .A(
        n17734), .ZN(n17758) );
  OAI21_X1 U20892 ( .B1(n17737), .B2(n17775), .A(n17758), .ZN(n17738) );
  AOI21_X1 U20893 ( .B1(n18469), .B2(n17739), .A(n17738), .ZN(n17751) );
  OR2_X1 U20894 ( .A1(n17741), .A2(n17740), .ZN(n17742) );
  AOI22_X1 U20895 ( .A1(n17743), .A2(n17751), .B1(n20826), .B2(n17742), .ZN(
        n17745) );
  AOI22_X1 U20896 ( .A1(n17989), .A2(n17745), .B1(n17910), .B2(n17744), .ZN(
        n17747) );
  OAI211_X1 U20897 ( .C1(n17980), .C2(n20826), .A(n17747), .B(n17746), .ZN(
        P3_U2840) );
  AOI22_X1 U20898 ( .A1(n17995), .A2(P3_REIP_REG_21__SCAN_IN), .B1(n17769), 
        .B2(n17748), .ZN(n17756) );
  NOR2_X1 U20899 ( .A1(n17928), .A2(n17749), .ZN(n17796) );
  OAI21_X1 U20900 ( .B1(n18465), .B2(n17750), .A(n17796), .ZN(n17760) );
  INV_X1 U20901 ( .A(n17826), .ZN(n17752) );
  OAI21_X1 U20902 ( .B1(n17753), .B2(n17752), .A(n17751), .ZN(n17754) );
  OAI211_X1 U20903 ( .C1(n17760), .C2(n17754), .A(
        P3_INSTADDRPOINTER_REG_21__SCAN_IN), .B(n17993), .ZN(n17755) );
  OAI211_X1 U20904 ( .C1(n17757), .C2(n17815), .A(n17756), .B(n17755), .ZN(
        P3_U2841) );
  NAND3_X1 U20905 ( .A1(n17773), .A2(P3_STATE2_REG_2__SCAN_IN), .A3(n17826), 
        .ZN(n17762) );
  OAI21_X1 U20906 ( .B1(n17759), .B2(n17775), .A(n17758), .ZN(n17761) );
  OAI21_X1 U20907 ( .B1(n17761), .B2(n17760), .A(n17993), .ZN(n17774) );
  NAND2_X1 U20908 ( .A1(n17762), .A2(n17774), .ZN(n17764) );
  AOI22_X1 U20909 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n17764), .B1(
        n17769), .B2(n17763), .ZN(n17766) );
  OAI211_X1 U20910 ( .C1(n17767), .C2(n17815), .A(n17766), .B(n17765), .ZN(
        P3_U2842) );
  AOI22_X1 U20911 ( .A1(n17910), .A2(n17770), .B1(n17769), .B2(n17768), .ZN(
        n17772) );
  OAI211_X1 U20912 ( .C1(n17774), .C2(n17773), .A(n17772), .B(n17771), .ZN(
        P3_U2843) );
  INV_X1 U20913 ( .A(n17775), .ZN(n17876) );
  NAND2_X1 U20914 ( .A1(n17877), .A2(n20755), .ZN(n17943) );
  NAND3_X1 U20915 ( .A1(n17776), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        n17943), .ZN(n17777) );
  AOI22_X1 U20916 ( .A1(n17778), .A2(n17876), .B1(n17781), .B2(n17777), .ZN(
        n17779) );
  OAI211_X1 U20917 ( .C1(n17780), .C2(n18481), .A(n17796), .B(n17779), .ZN(
        n17791) );
  OAI221_X1 U20918 ( .B1(n17791), .B2(n17782), .C1(n17791), .C2(n17781), .A(
        P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n17790) );
  INV_X1 U20919 ( .A(n17973), .ZN(n17946) );
  OAI22_X1 U20920 ( .A1(n17946), .A2(n18481), .B1(n17783), .B2(n17965), .ZN(
        n17954) );
  NAND2_X1 U20921 ( .A1(n17784), .A2(n17954), .ZN(n17916) );
  NOR2_X1 U20922 ( .A1(n17785), .A2(n17916), .ZN(n17823) );
  NAND2_X1 U20923 ( .A1(n17800), .A2(n17823), .ZN(n17809) );
  AOI211_X1 U20924 ( .C1(n17786), .C2(n17809), .A(n17822), .B(n17928), .ZN(
        n17803) );
  AOI22_X1 U20925 ( .A1(n17910), .A2(n17788), .B1(n17803), .B2(n17787), .ZN(
        n17789) );
  OAI221_X1 U20926 ( .B1(n17995), .B2(n17790), .C1(n17993), .C2(n18559), .A(
        n17789), .ZN(P3_U2844) );
  NAND2_X1 U20927 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n17791), .ZN(
        n17795) );
  AOI22_X1 U20928 ( .A1(n17910), .A2(n17793), .B1(n17803), .B2(n17792), .ZN(
        n17794) );
  OAI221_X1 U20929 ( .B1(n17979), .B2(n17795), .C1(n17993), .C2(n18558), .A(
        n17794), .ZN(P3_U2845) );
  INV_X1 U20930 ( .A(n17796), .ZN(n17801) );
  NOR2_X1 U20931 ( .A1(n17797), .A2(n18481), .ZN(n17871) );
  AOI21_X1 U20932 ( .B1(n18469), .B2(n17885), .A(n17871), .ZN(n17827) );
  OAI21_X1 U20933 ( .B1(n17822), .B2(n17877), .A(n17798), .ZN(n17799) );
  OAI211_X1 U20934 ( .C1(n17887), .C2(n17800), .A(n17827), .B(n17799), .ZN(
        n17811) );
  OAI221_X1 U20935 ( .B1(n17801), .B2(n17903), .C1(n17801), .C2(n17811), .A(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n17806) );
  AOI22_X1 U20936 ( .A1(n17804), .A2(n17910), .B1(n17803), .B2(n17802), .ZN(
        n17805) );
  OAI221_X1 U20937 ( .B1(n17995), .B2(n17806), .C1(n17993), .C2(n18555), .A(
        n17805), .ZN(P3_U2846) );
  NOR2_X1 U20938 ( .A1(n17807), .A2(n17999), .ZN(n17819) );
  NOR2_X1 U20939 ( .A1(n17808), .A2(n17873), .ZN(n17813) );
  NAND2_X1 U20940 ( .A1(n17822), .A2(n17809), .ZN(n17810) );
  AOI22_X1 U20941 ( .A1(n17813), .A2(n17812), .B1(n17811), .B2(n17810), .ZN(
        n17816) );
  OAI22_X1 U20942 ( .A1(n17816), .A2(n17928), .B1(n17815), .B2(n17814), .ZN(
        n17817) );
  AOI21_X1 U20943 ( .B1(n17819), .B2(n17818), .A(n17817), .ZN(n17821) );
  NAND2_X1 U20944 ( .A1(n17995), .A2(P3_REIP_REG_15__SCAN_IN), .ZN(n17820) );
  OAI211_X1 U20945 ( .C1(n17980), .C2(n17822), .A(n17821), .B(n17820), .ZN(
        P3_U2847) );
  AOI21_X1 U20946 ( .B1(n17824), .B2(n17823), .A(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n17825) );
  INV_X1 U20947 ( .A(n17825), .ZN(n17834) );
  NAND2_X1 U20948 ( .A1(n17989), .A2(n17826), .ZN(n17991) );
  AOI21_X1 U20949 ( .B1(n17854), .B2(n17869), .A(n18465), .ZN(n17850) );
  OAI211_X1 U20950 ( .C1(n17854), .C2(n18481), .A(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B(n17827), .ZN(n17828) );
  AOI211_X1 U20951 ( .C1(n18469), .C2(n17829), .A(n17850), .B(n17828), .ZN(
        n17830) );
  OAI222_X1 U20952 ( .A1(n17980), .A2(n17831), .B1(n17991), .B2(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .C1(n17928), .C2(n17830), .ZN(
        n17833) );
  AOI21_X1 U20953 ( .B1(n17834), .B2(n17833), .A(n17832), .ZN(n17838) );
  AOI22_X1 U20954 ( .A1(n17911), .A2(n17836), .B1(n17910), .B2(n17835), .ZN(
        n17837) );
  OAI211_X1 U20955 ( .C1(n17999), .C2(n17839), .A(n17838), .B(n17837), .ZN(
        P3_U2848) );
  NAND3_X1 U20956 ( .A1(n17989), .A2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        n17954), .ZN(n17947) );
  NOR3_X1 U20957 ( .A1(n17936), .A2(n17948), .A3(n17947), .ZN(n17931) );
  AOI222_X1 U20958 ( .A1(n17868), .A2(n17982), .B1(n17874), .B2(n17911), .C1(
        n17840), .C2(n17931), .ZN(n17898) );
  AOI22_X1 U20959 ( .A1(n17979), .A2(P3_REIP_REG_13__SCAN_IN), .B1(n17910), 
        .B2(n17841), .ZN(n17852) );
  AOI21_X1 U20960 ( .B1(n18469), .B2(n17842), .A(n17864), .ZN(n17856) );
  INV_X1 U20961 ( .A(n17885), .ZN(n17843) );
  AOI21_X1 U20962 ( .B1(n17844), .B2(n17843), .A(n17990), .ZN(n17845) );
  AOI21_X1 U20963 ( .B1(n18449), .B2(n17858), .A(n17845), .ZN(n17878) );
  OAI21_X1 U20964 ( .B1(n17846), .B2(n17873), .A(n17878), .ZN(n17847) );
  AOI211_X1 U20965 ( .C1(n18447), .C2(n17848), .A(n17871), .B(n17847), .ZN(
        n17855) );
  OAI211_X1 U20966 ( .C1(n17887), .C2(n17856), .A(n17989), .B(n17855), .ZN(
        n17849) );
  OAI211_X1 U20967 ( .C1(n17850), .C2(n17849), .A(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B(n17993), .ZN(n17851) );
  OAI211_X1 U20968 ( .C1(n17898), .C2(n17853), .A(n17852), .B(n17851), .ZN(
        P3_U2849) );
  AND2_X1 U20969 ( .A1(n17854), .A2(n17869), .ZN(n17857) );
  OAI211_X1 U20970 ( .C1(n17857), .C2(n18465), .A(n17856), .B(n17855), .ZN(
        n17860) );
  OAI22_X1 U20971 ( .A1(n17898), .A2(n17858), .B1(n17864), .B2(n17928), .ZN(
        n17859) );
  AOI22_X1 U20972 ( .A1(n17910), .A2(n17861), .B1(n17860), .B2(n17859), .ZN(
        n17863) );
  OAI211_X1 U20973 ( .C1(n17980), .C2(n17864), .A(n17863), .B(n17862), .ZN(
        P3_U2850) );
  INV_X1 U20974 ( .A(n17898), .ZN(n17865) );
  AOI22_X1 U20975 ( .A1(n17910), .A2(n17867), .B1(n17866), .B2(n17865), .ZN(
        n17882) );
  OAI22_X1 U20976 ( .A1(n18465), .A2(n17869), .B1(n17868), .B2(n17972), .ZN(
        n17870) );
  NOR3_X1 U20977 ( .A1(n17871), .A2(n17928), .A3(n17870), .ZN(n17872) );
  OAI21_X1 U20978 ( .B1(n17874), .B2(n17873), .A(n17872), .ZN(n17884) );
  OAI21_X1 U20979 ( .B1(n17877), .B2(n17876), .A(n17875), .ZN(n17886) );
  NAND2_X1 U20980 ( .A1(n17878), .A2(n17886), .ZN(n17879) );
  OAI211_X1 U20981 ( .C1(n17884), .C2(n17879), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n17993), .ZN(n17880) );
  NAND3_X1 U20982 ( .A1(n17882), .A2(n17881), .A3(n17880), .ZN(P3_U2851) );
  AOI22_X1 U20983 ( .A1(n17995), .A2(P3_REIP_REG_10__SCAN_IN), .B1(n17910), 
        .B2(n17883), .ZN(n17890) );
  AOI21_X1 U20984 ( .B1(n18469), .B2(n17885), .A(n17884), .ZN(n17893) );
  OAI211_X1 U20985 ( .C1(n17887), .C2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n17893), .B(n17886), .ZN(n17888) );
  NAND3_X1 U20986 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n17993), .A3(
        n17888), .ZN(n17889) );
  OAI211_X1 U20987 ( .C1(n17898), .C2(n17891), .A(n17890), .B(n17889), .ZN(
        P3_U2852) );
  NOR3_X1 U20988 ( .A1(n17979), .A2(n17893), .A3(n17892), .ZN(n17894) );
  AOI211_X1 U20989 ( .C1(n17910), .C2(n17896), .A(n17895), .B(n17894), .ZN(
        n17897) );
  OAI21_X1 U20990 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n17898), .A(
        n17897), .ZN(P3_U2853) );
  AND3_X1 U20991 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A3(n17931), .ZN(n17908) );
  NAND2_X1 U20992 ( .A1(n18449), .A2(n17899), .ZN(n17900) );
  OAI211_X1 U20993 ( .C1(n17901), .C2(n17944), .A(n17900), .B(n17943), .ZN(
        n17927) );
  AOI211_X1 U20994 ( .C1(n17903), .C2(n17930), .A(n17902), .B(n17927), .ZN(
        n17925) );
  OAI21_X1 U20995 ( .B1(n17925), .B2(n17987), .A(n17980), .ZN(n17906) );
  INV_X1 U20996 ( .A(n17904), .ZN(n17905) );
  AOI221_X1 U20997 ( .B1(n17908), .B2(n17907), .C1(n17906), .C2(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A(n17905), .ZN(n17914) );
  AOI22_X1 U20998 ( .A1(n17912), .A2(n17911), .B1(n17910), .B2(n17909), .ZN(
        n17913) );
  OAI211_X1 U20999 ( .C1(n17999), .C2(n17915), .A(n17914), .B(n17913), .ZN(
        P3_U2854) );
  NOR2_X1 U21000 ( .A1(n17930), .A2(n17916), .ZN(n17917) );
  OAI21_X1 U21001 ( .B1(n17917), .B2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n17989), .ZN(n17924) );
  AOI22_X1 U21002 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n17918), .B1(
        n17995), .B2(P3_REIP_REG_7__SCAN_IN), .ZN(n17923) );
  INV_X1 U21003 ( .A(n17919), .ZN(n18444) );
  NOR2_X1 U21004 ( .A1(n18444), .A2(n17928), .ZN(n17988) );
  AOI22_X1 U21005 ( .A1(n17982), .A2(n17921), .B1(n17920), .B2(n17988), .ZN(
        n17922) );
  OAI211_X1 U21006 ( .C1(n17925), .C2(n17924), .A(n17923), .B(n17922), .ZN(
        P3_U2855) );
  AOI22_X1 U21007 ( .A1(n17995), .A2(P3_REIP_REG_6__SCAN_IN), .B1(n17988), 
        .B2(n17926), .ZN(n17933) );
  INV_X1 U21008 ( .A(n17927), .ZN(n17929) );
  OAI21_X1 U21009 ( .B1(n17929), .B2(n17928), .A(n17980), .ZN(n17937) );
  AOI22_X1 U21010 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n17937), .B1(
        n17931), .B2(n17930), .ZN(n17932) );
  OAI211_X1 U21011 ( .C1(n17999), .C2(n17934), .A(n17933), .B(n17932), .ZN(
        P3_U2856) );
  AOI22_X1 U21012 ( .A1(n17995), .A2(P3_REIP_REG_5__SCAN_IN), .B1(n17988), 
        .B2(n17935), .ZN(n17940) );
  OAI21_X1 U21013 ( .B1(n17948), .B2(n17947), .A(n17936), .ZN(n17938) );
  NAND2_X1 U21014 ( .A1(n17938), .A2(n17937), .ZN(n17939) );
  OAI211_X1 U21015 ( .C1(n17999), .C2(n17941), .A(n17940), .B(n17939), .ZN(
        P3_U2857) );
  AOI22_X1 U21016 ( .A1(n17995), .A2(P3_REIP_REG_4__SCAN_IN), .B1(n17988), 
        .B2(n17942), .ZN(n17952) );
  OAI21_X1 U21017 ( .B1(n17945), .B2(n17944), .A(n17943), .ZN(n17966) );
  AOI211_X1 U21018 ( .C1(n18449), .C2(n17946), .A(n17955), .B(n17966), .ZN(
        n17957) );
  OAI21_X1 U21019 ( .B1(n17957), .B2(n17987), .A(n17980), .ZN(n17950) );
  INV_X1 U21020 ( .A(n17947), .ZN(n17949) );
  AOI22_X1 U21021 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n17950), .B1(
        n17949), .B2(n17948), .ZN(n17951) );
  OAI211_X1 U21022 ( .C1(n17999), .C2(n17953), .A(n17952), .B(n17951), .ZN(
        P3_U2858) );
  NOR2_X1 U21023 ( .A1(n17993), .A2(n18532), .ZN(n17959) );
  OAI21_X1 U21024 ( .B1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n17954), .A(
        n17989), .ZN(n17956) );
  OAI22_X1 U21025 ( .A1(n17957), .A2(n17956), .B1(n17955), .B2(n17980), .ZN(
        n17958) );
  AOI211_X1 U21026 ( .C1(n17988), .C2(n17960), .A(n17959), .B(n17958), .ZN(
        n17961) );
  OAI21_X1 U21027 ( .B1(n17999), .B2(n17962), .A(n17961), .ZN(P3_U2859) );
  AOI21_X1 U21028 ( .B1(n17988), .B2(n17964), .A(n17963), .ZN(n17977) );
  NOR2_X1 U21029 ( .A1(n18612), .A2(n17965), .ZN(n17970) );
  NOR2_X1 U21030 ( .A1(n20755), .A2(n18612), .ZN(n17967) );
  AOI21_X1 U21031 ( .B1(n18449), .B2(n17967), .A(n17966), .ZN(n17968) );
  INV_X1 U21032 ( .A(n17968), .ZN(n17969) );
  MUX2_X1 U21033 ( .A(n17970), .B(n17969), .S(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .Z(n17975) );
  OAI22_X1 U21034 ( .A1(n18481), .A2(n17973), .B1(n17972), .B2(n17971), .ZN(
        n17974) );
  OAI21_X1 U21035 ( .B1(n17975), .B2(n17974), .A(n17989), .ZN(n17976) );
  OAI211_X1 U21036 ( .C1(n17980), .C2(n20894), .A(n17977), .B(n17976), .ZN(
        P3_U2860) );
  OAI21_X1 U21037 ( .B1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n18469), .A(
        n18612), .ZN(n17986) );
  AOI22_X1 U21038 ( .A1(n17979), .A2(P3_REIP_REG_1__SCAN_IN), .B1(n17988), 
        .B2(n17978), .ZN(n17985) );
  OAI21_X1 U21039 ( .B1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n17991), .A(
        n17980), .ZN(n17983) );
  AOI22_X1 U21040 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n17983), .B1(
        n17982), .B2(n17981), .ZN(n17984) );
  OAI211_X1 U21041 ( .C1(n17987), .C2(n17986), .A(n17985), .B(n17984), .ZN(
        P3_U2861) );
  INV_X1 U21042 ( .A(n17988), .ZN(n17997) );
  AOI21_X1 U21043 ( .B1(n17990), .B2(n17989), .A(n20755), .ZN(n17994) );
  NOR2_X1 U21044 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n17991), .ZN(
        n17992) );
  AOI221_X1 U21045 ( .B1(P3_REIP_REG_0__SCAN_IN), .B2(n17995), .C1(n17994), 
        .C2(n17993), .A(n17992), .ZN(n17996) );
  OAI221_X1 U21046 ( .B1(n18000), .B2(n17999), .C1(n17998), .C2(n17997), .A(
        n17996), .ZN(P3_U2862) );
  OAI211_X1 U21047 ( .C1(P3_FLUSH_REG_SCAN_IN), .C2(n18001), .A(
        P3_STATE2_REG_2__SCAN_IN), .B(P3_STATE2_REG_1__SCAN_IN), .ZN(n18502)
         );
  OAI21_X1 U21048 ( .B1(n18004), .B2(n18002), .A(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18003) );
  OAI221_X1 U21049 ( .B1(n18004), .B2(n18502), .C1(n18004), .C2(n18063), .A(
        n18003), .ZN(P3_U2863) );
  NOR2_X1 U21050 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18013), .ZN(
        n18194) );
  INV_X1 U21051 ( .A(n18194), .ZN(n18148) );
  NOR2_X1 U21052 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18487), .ZN(
        n18289) );
  NAND2_X1 U21053 ( .A1(n18083), .A2(n18289), .ZN(n18310) );
  AND2_X1 U21054 ( .A1(n18148), .A2(n18310), .ZN(n18006) );
  OAI22_X1 U21055 ( .A1(n18007), .A2(n18487), .B1(n18006), .B2(n18005), .ZN(
        P3_U2866) );
  NOR2_X1 U21056 ( .A1(n18009), .A2(n18008), .ZN(P3_U2867) );
  NOR2_X1 U21057 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18471) );
  NOR2_X1 U21058 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18105) );
  NAND2_X1 U21059 ( .A1(n18471), .A2(n18105), .ZN(n18062) );
  NOR2_X1 U21060 ( .A1(n18011), .A2(n18010), .ZN(n18053) );
  NAND2_X1 U21061 ( .A1(n18053), .A2(n18012), .ZN(n18394) );
  NOR2_X1 U21062 ( .A1(n18013), .A2(n18487), .ZN(n18015) );
  NAND2_X1 U21063 ( .A1(n18015), .A2(n18288), .ZN(n18334) );
  NOR2_X2 U21064 ( .A1(n18309), .A2(n18334), .ZN(n18436) );
  AND2_X1 U21065 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n18390), .ZN(n18386) );
  NOR2_X2 U21066 ( .A1(n18054), .A2(n18014), .ZN(n18385) );
  INV_X1 U21067 ( .A(n18505), .ZN(n18357) );
  NOR2_X1 U21068 ( .A1(n18288), .A2(n18309), .ZN(n18470) );
  INV_X1 U21069 ( .A(n18470), .ZN(n18016) );
  INV_X1 U21070 ( .A(n18015), .ZN(n18020) );
  NOR2_X2 U21071 ( .A1(n18016), .A2(n18020), .ZN(n18384) );
  INV_X1 U21072 ( .A(n18062), .ZN(n18121) );
  NOR2_X1 U21073 ( .A1(n18384), .A2(n18121), .ZN(n18084) );
  NOR2_X1 U21074 ( .A1(n18357), .A2(n18084), .ZN(n18056) );
  AOI22_X1 U21075 ( .A1(n18436), .A2(n18386), .B1(n18385), .B2(n18056), .ZN(
        n18022) );
  AOI21_X1 U21076 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n18084), .ZN(n18017) );
  NOR2_X1 U21077 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18288), .ZN(
        n18263) );
  NOR2_X1 U21078 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18309), .ZN(
        n18238) );
  NOR2_X1 U21079 ( .A1(n18263), .A2(n18238), .ZN(n18311) );
  NOR2_X1 U21080 ( .A1(n18311), .A2(n18020), .ZN(n18356) );
  AOI22_X1 U21081 ( .A1(n18362), .A2(n18017), .B1(n18390), .B2(n18356), .ZN(
        n18059) );
  NOR2_X2 U21082 ( .A1(n18057), .A2(n18018), .ZN(n18391) );
  INV_X1 U21083 ( .A(n18263), .ZN(n18019) );
  NOR2_X2 U21084 ( .A1(n18020), .A2(n18019), .ZN(n18363) );
  AOI22_X1 U21085 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n18059), .B1(
        n18391), .B2(n18363), .ZN(n18021) );
  OAI211_X1 U21086 ( .C1(n18062), .C2(n18394), .A(n18022), .B(n18021), .ZN(
        P3_U2868) );
  NAND2_X1 U21087 ( .A1(n18053), .A2(n18023), .ZN(n18400) );
  AND2_X1 U21088 ( .A1(n18390), .A2(BUF2_REG_17__SCAN_IN), .ZN(n18397) );
  NOR2_X2 U21089 ( .A1(n18054), .A2(n18024), .ZN(n18395) );
  AOI22_X1 U21090 ( .A1(n18363), .A2(n18397), .B1(n18056), .B2(n18395), .ZN(
        n18026) );
  NOR2_X2 U21091 ( .A1(n20723), .A2(n18057), .ZN(n18396) );
  AOI22_X1 U21092 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n18059), .B1(
        n18436), .B2(n18396), .ZN(n18025) );
  OAI211_X1 U21093 ( .C1(n18062), .C2(n18400), .A(n18026), .B(n18025), .ZN(
        P3_U2869) );
  NAND2_X1 U21094 ( .A1(n18053), .A2(n18027), .ZN(n18406) );
  NOR2_X2 U21095 ( .A1(n18057), .A2(n19070), .ZN(n18403) );
  NOR2_X2 U21096 ( .A1(n18054), .A2(n18028), .ZN(n18401) );
  AOI22_X1 U21097 ( .A1(n18363), .A2(n18403), .B1(n18056), .B2(n18401), .ZN(
        n18031) );
  NOR2_X2 U21098 ( .A1(n18029), .A2(n18057), .ZN(n18402) );
  AOI22_X1 U21099 ( .A1(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n18059), .B1(
        n18436), .B2(n18402), .ZN(n18030) );
  OAI211_X1 U21100 ( .C1(n18062), .C2(n18406), .A(n18031), .B(n18030), .ZN(
        P3_U2870) );
  NAND2_X1 U21101 ( .A1(n18053), .A2(n18032), .ZN(n18412) );
  AND2_X1 U21102 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n18390), .ZN(n18408) );
  NOR2_X2 U21103 ( .A1(n18033), .A2(n18054), .ZN(n18407) );
  AOI22_X1 U21104 ( .A1(n18436), .A2(n18408), .B1(n18056), .B2(n18407), .ZN(
        n18036) );
  NOR2_X2 U21105 ( .A1(n18034), .A2(n18057), .ZN(n18409) );
  AOI22_X1 U21106 ( .A1(P3_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n18059), .B1(
        n18363), .B2(n18409), .ZN(n18035) );
  OAI211_X1 U21107 ( .C1(n18062), .C2(n18412), .A(n18036), .B(n18035), .ZN(
        P3_U2871) );
  NAND2_X1 U21108 ( .A1(n18053), .A2(n18037), .ZN(n18418) );
  NOR2_X2 U21109 ( .A1(n20770), .A2(n18057), .ZN(n18414) );
  NOR2_X2 U21110 ( .A1(n18038), .A2(n18054), .ZN(n18413) );
  AOI22_X1 U21111 ( .A1(n18363), .A2(n18414), .B1(n18056), .B2(n18413), .ZN(
        n18040) );
  AND2_X1 U21112 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n18390), .ZN(n18415) );
  AOI22_X1 U21113 ( .A1(P3_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n18059), .B1(
        n18436), .B2(n18415), .ZN(n18039) );
  OAI211_X1 U21114 ( .C1(n18062), .C2(n18418), .A(n18040), .B(n18039), .ZN(
        P3_U2872) );
  NAND2_X1 U21115 ( .A1(n18053), .A2(n18041), .ZN(n18424) );
  NOR2_X2 U21116 ( .A1(n18042), .A2(n18057), .ZN(n18420) );
  AND2_X1 U21117 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n18362), .ZN(n18419) );
  AOI22_X1 U21118 ( .A1(n18363), .A2(n18420), .B1(n18056), .B2(n18419), .ZN(
        n18045) );
  NOR2_X2 U21119 ( .A1(n18043), .A2(n18057), .ZN(n18421) );
  AOI22_X1 U21120 ( .A1(P3_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n18059), .B1(
        n18436), .B2(n18421), .ZN(n18044) );
  OAI211_X1 U21121 ( .C1(n18062), .C2(n18424), .A(n18045), .B(n18044), .ZN(
        P3_U2873) );
  NAND2_X1 U21122 ( .A1(n18053), .A2(n18046), .ZN(n18430) );
  NOR2_X2 U21123 ( .A1(n18047), .A2(n18057), .ZN(n18426) );
  NOR2_X2 U21124 ( .A1(n18048), .A2(n18054), .ZN(n18425) );
  AOI22_X1 U21125 ( .A1(n18363), .A2(n18426), .B1(n18056), .B2(n18425), .ZN(
        n18051) );
  NOR2_X2 U21126 ( .A1(n18049), .A2(n18057), .ZN(n18427) );
  AOI22_X1 U21127 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n18059), .B1(
        n18436), .B2(n18427), .ZN(n18050) );
  OAI211_X1 U21128 ( .C1(n18062), .C2(n18430), .A(n18051), .B(n18050), .ZN(
        P3_U2874) );
  NAND2_X1 U21129 ( .A1(n18053), .A2(n18052), .ZN(n18440) );
  AND2_X1 U21130 ( .A1(BUF2_REG_23__SCAN_IN), .A2(n18390), .ZN(n18435) );
  NOR2_X2 U21131 ( .A1(n18055), .A2(n18054), .ZN(n18432) );
  AOI22_X1 U21132 ( .A1(n18363), .A2(n18435), .B1(n18056), .B2(n18432), .ZN(
        n18061) );
  NOR2_X2 U21133 ( .A1(n18058), .A2(n18057), .ZN(n18434) );
  AOI22_X1 U21134 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n18059), .B1(
        n18436), .B2(n18434), .ZN(n18060) );
  OAI211_X1 U21135 ( .C1(n18062), .C2(n18440), .A(n18061), .B(n18060), .ZN(
        P3_U2875) );
  NAND2_X1 U21136 ( .A1(n18238), .A2(n18105), .ZN(n18082) );
  INV_X1 U21137 ( .A(n18105), .ZN(n18149) );
  NAND2_X1 U21138 ( .A1(n18288), .A2(n18505), .ZN(n18239) );
  NOR2_X1 U21139 ( .A1(n18149), .A2(n18239), .ZN(n18078) );
  AOI22_X1 U21140 ( .A1(n18363), .A2(n18386), .B1(n18385), .B2(n18078), .ZN(
        n18065) );
  NOR2_X1 U21141 ( .A1(n18487), .A2(n18240), .ZN(n18387) );
  NAND2_X1 U21142 ( .A1(n18362), .A2(n18063), .ZN(n18241) );
  NOR2_X1 U21143 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18241), .ZN(
        n18150) );
  AOI22_X1 U21144 ( .A1(n18390), .A2(n18387), .B1(n18105), .B2(n18150), .ZN(
        n18079) );
  AOI22_X1 U21145 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n18079), .B1(
        n18384), .B2(n18391), .ZN(n18064) );
  OAI211_X1 U21146 ( .C1(n18394), .C2(n18082), .A(n18065), .B(n18064), .ZN(
        P3_U2876) );
  AOI22_X1 U21147 ( .A1(n18363), .A2(n18396), .B1(n18395), .B2(n18078), .ZN(
        n18067) );
  AOI22_X1 U21148 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n18079), .B1(
        n18384), .B2(n18397), .ZN(n18066) );
  OAI211_X1 U21149 ( .C1(n18400), .C2(n18082), .A(n18067), .B(n18066), .ZN(
        P3_U2877) );
  AOI22_X1 U21150 ( .A1(n18384), .A2(n18403), .B1(n18401), .B2(n18078), .ZN(
        n18069) );
  AOI22_X1 U21151 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n18079), .B1(
        n18363), .B2(n18402), .ZN(n18068) );
  OAI211_X1 U21152 ( .C1(n18406), .C2(n18082), .A(n18069), .B(n18068), .ZN(
        P3_U2878) );
  AOI22_X1 U21153 ( .A1(n18384), .A2(n18409), .B1(n18407), .B2(n18078), .ZN(
        n18071) );
  AOI22_X1 U21154 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n18079), .B1(
        n18363), .B2(n18408), .ZN(n18070) );
  OAI211_X1 U21155 ( .C1(n18412), .C2(n18082), .A(n18071), .B(n18070), .ZN(
        P3_U2879) );
  AOI22_X1 U21156 ( .A1(n18363), .A2(n18415), .B1(n18413), .B2(n18078), .ZN(
        n18073) );
  AOI22_X1 U21157 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n18079), .B1(
        n18384), .B2(n18414), .ZN(n18072) );
  OAI211_X1 U21158 ( .C1(n18418), .C2(n18082), .A(n18073), .B(n18072), .ZN(
        P3_U2880) );
  AOI22_X1 U21159 ( .A1(n18384), .A2(n18420), .B1(n18419), .B2(n18078), .ZN(
        n18075) );
  AOI22_X1 U21160 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n18079), .B1(
        n18363), .B2(n18421), .ZN(n18074) );
  OAI211_X1 U21161 ( .C1(n18424), .C2(n18082), .A(n18075), .B(n18074), .ZN(
        P3_U2881) );
  AOI22_X1 U21162 ( .A1(n18363), .A2(n18427), .B1(n18425), .B2(n18078), .ZN(
        n18077) );
  AOI22_X1 U21163 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n18079), .B1(
        n18384), .B2(n18426), .ZN(n18076) );
  OAI211_X1 U21164 ( .C1(n18430), .C2(n18082), .A(n18077), .B(n18076), .ZN(
        P3_U2882) );
  AOI22_X1 U21165 ( .A1(n18384), .A2(n18435), .B1(n18432), .B2(n18078), .ZN(
        n18081) );
  AOI22_X1 U21166 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n18079), .B1(
        n18363), .B2(n18434), .ZN(n18080) );
  OAI211_X1 U21167 ( .C1(n18440), .C2(n18082), .A(n18081), .B(n18080), .ZN(
        P3_U2883) );
  NAND2_X1 U21168 ( .A1(n18263), .A2(n18105), .ZN(n18104) );
  INV_X1 U21169 ( .A(n18082), .ZN(n18144) );
  INV_X1 U21170 ( .A(n18104), .ZN(n18167) );
  NOR2_X1 U21171 ( .A1(n18144), .A2(n18167), .ZN(n18126) );
  NOR2_X1 U21172 ( .A1(n18357), .A2(n18126), .ZN(n18100) );
  AOI22_X1 U21173 ( .A1(n18384), .A2(n18386), .B1(n18385), .B2(n18100), .ZN(
        n18087) );
  INV_X1 U21174 ( .A(n18083), .ZN(n18359) );
  OAI21_X1 U21175 ( .B1(n18084), .B2(n18359), .A(n18126), .ZN(n18085) );
  OAI211_X1 U21176 ( .C1(n18167), .C2(n18599), .A(n18362), .B(n18085), .ZN(
        n18101) );
  AOI22_X1 U21177 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n18101), .B1(
        n18121), .B2(n18391), .ZN(n18086) );
  OAI211_X1 U21178 ( .C1(n18394), .C2(n18104), .A(n18087), .B(n18086), .ZN(
        P3_U2884) );
  AOI22_X1 U21179 ( .A1(n18384), .A2(n18396), .B1(n18395), .B2(n18100), .ZN(
        n18089) );
  AOI22_X1 U21180 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n18101), .B1(
        n18121), .B2(n18397), .ZN(n18088) );
  OAI211_X1 U21181 ( .C1(n18400), .C2(n18104), .A(n18089), .B(n18088), .ZN(
        P3_U2885) );
  AOI22_X1 U21182 ( .A1(n18121), .A2(n18403), .B1(n18401), .B2(n18100), .ZN(
        n18091) );
  AOI22_X1 U21183 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n18101), .B1(
        n18384), .B2(n18402), .ZN(n18090) );
  OAI211_X1 U21184 ( .C1(n18406), .C2(n18104), .A(n18091), .B(n18090), .ZN(
        P3_U2886) );
  AOI22_X1 U21185 ( .A1(n18121), .A2(n18409), .B1(n18407), .B2(n18100), .ZN(
        n18093) );
  AOI22_X1 U21186 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n18101), .B1(
        n18384), .B2(n18408), .ZN(n18092) );
  OAI211_X1 U21187 ( .C1(n18412), .C2(n18104), .A(n18093), .B(n18092), .ZN(
        P3_U2887) );
  AOI22_X1 U21188 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n18101), .B1(
        n18413), .B2(n18100), .ZN(n18095) );
  AOI22_X1 U21189 ( .A1(n18384), .A2(n18415), .B1(n18121), .B2(n18414), .ZN(
        n18094) );
  OAI211_X1 U21190 ( .C1(n18418), .C2(n18104), .A(n18095), .B(n18094), .ZN(
        P3_U2888) );
  AOI22_X1 U21191 ( .A1(n18384), .A2(n18421), .B1(n18419), .B2(n18100), .ZN(
        n18097) );
  AOI22_X1 U21192 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n18101), .B1(
        n18121), .B2(n18420), .ZN(n18096) );
  OAI211_X1 U21193 ( .C1(n18424), .C2(n18104), .A(n18097), .B(n18096), .ZN(
        P3_U2889) );
  AOI22_X1 U21194 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n18101), .B1(
        n18425), .B2(n18100), .ZN(n18099) );
  AOI22_X1 U21195 ( .A1(n18384), .A2(n18427), .B1(n18121), .B2(n18426), .ZN(
        n18098) );
  OAI211_X1 U21196 ( .C1(n18430), .C2(n18104), .A(n18099), .B(n18098), .ZN(
        P3_U2890) );
  AOI22_X1 U21197 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n18101), .B1(
        n18432), .B2(n18100), .ZN(n18103) );
  AOI22_X1 U21198 ( .A1(n18384), .A2(n18434), .B1(n18121), .B2(n18435), .ZN(
        n18102) );
  OAI211_X1 U21199 ( .C1(n18440), .C2(n18104), .A(n18103), .B(n18102), .ZN(
        P3_U2891) );
  NAND2_X1 U21200 ( .A1(n18470), .A2(n18105), .ZN(n18125) );
  AOI22_X1 U21201 ( .A1(n18121), .A2(n18386), .B1(n18385), .B2(n18120), .ZN(
        n18107) );
  AOI21_X1 U21202 ( .B1(n18288), .B2(n18359), .A(n18241), .ZN(n18195) );
  NAND2_X1 U21203 ( .A1(n18105), .A2(n18195), .ZN(n18122) );
  AOI22_X1 U21204 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n18122), .B1(
        n18391), .B2(n18144), .ZN(n18106) );
  OAI211_X1 U21205 ( .C1(n18394), .C2(n18125), .A(n18107), .B(n18106), .ZN(
        P3_U2892) );
  AOI22_X1 U21206 ( .A1(n18121), .A2(n18396), .B1(n18395), .B2(n18120), .ZN(
        n18109) );
  AOI22_X1 U21207 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n18122), .B1(
        n18397), .B2(n18144), .ZN(n18108) );
  OAI211_X1 U21208 ( .C1(n18400), .C2(n18125), .A(n18109), .B(n18108), .ZN(
        P3_U2893) );
  AOI22_X1 U21209 ( .A1(n18121), .A2(n18402), .B1(n18401), .B2(n18120), .ZN(
        n18111) );
  AOI22_X1 U21210 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n18122), .B1(
        n18403), .B2(n18144), .ZN(n18110) );
  OAI211_X1 U21211 ( .C1(n18406), .C2(n18125), .A(n18111), .B(n18110), .ZN(
        P3_U2894) );
  AOI22_X1 U21212 ( .A1(n18409), .A2(n18144), .B1(n18407), .B2(n18120), .ZN(
        n18113) );
  AOI22_X1 U21213 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n18122), .B1(
        n18121), .B2(n18408), .ZN(n18112) );
  OAI211_X1 U21214 ( .C1(n18412), .C2(n18125), .A(n18113), .B(n18112), .ZN(
        P3_U2895) );
  AOI22_X1 U21215 ( .A1(n18414), .A2(n18144), .B1(n18413), .B2(n18120), .ZN(
        n18115) );
  AOI22_X1 U21216 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n18122), .B1(
        n18121), .B2(n18415), .ZN(n18114) );
  OAI211_X1 U21217 ( .C1(n18418), .C2(n18125), .A(n18115), .B(n18114), .ZN(
        P3_U2896) );
  AOI22_X1 U21218 ( .A1(n18121), .A2(n18421), .B1(n18419), .B2(n18120), .ZN(
        n18117) );
  AOI22_X1 U21219 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n18122), .B1(
        n18420), .B2(n18144), .ZN(n18116) );
  OAI211_X1 U21220 ( .C1(n18424), .C2(n18125), .A(n18117), .B(n18116), .ZN(
        P3_U2897) );
  AOI22_X1 U21221 ( .A1(n18121), .A2(n18427), .B1(n18425), .B2(n18120), .ZN(
        n18119) );
  AOI22_X1 U21222 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n18122), .B1(
        n18426), .B2(n18144), .ZN(n18118) );
  OAI211_X1 U21223 ( .C1(n18430), .C2(n18125), .A(n18119), .B(n18118), .ZN(
        P3_U2898) );
  AOI22_X1 U21224 ( .A1(n18435), .A2(n18144), .B1(n18432), .B2(n18120), .ZN(
        n18124) );
  AOI22_X1 U21225 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n18122), .B1(
        n18121), .B2(n18434), .ZN(n18123) );
  OAI211_X1 U21226 ( .C1(n18440), .C2(n18125), .A(n18124), .B(n18123), .ZN(
        P3_U2899) );
  NAND2_X1 U21227 ( .A1(n18471), .A2(n18194), .ZN(n18147) );
  INV_X1 U21228 ( .A(n18125), .ZN(n18190) );
  INV_X1 U21229 ( .A(n18147), .ZN(n18211) );
  NOR2_X1 U21230 ( .A1(n18190), .A2(n18211), .ZN(n18172) );
  NOR2_X1 U21231 ( .A1(n18357), .A2(n18172), .ZN(n18142) );
  AOI22_X1 U21232 ( .A1(n18391), .A2(n18167), .B1(n18385), .B2(n18142), .ZN(
        n18129) );
  OAI21_X1 U21233 ( .B1(n18126), .B2(n18359), .A(n18172), .ZN(n18127) );
  OAI211_X1 U21234 ( .C1(n18211), .C2(n18599), .A(n18362), .B(n18127), .ZN(
        n18143) );
  AOI22_X1 U21235 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n18143), .B1(
        n18386), .B2(n18144), .ZN(n18128) );
  OAI211_X1 U21236 ( .C1(n18394), .C2(n18147), .A(n18129), .B(n18128), .ZN(
        P3_U2900) );
  AOI22_X1 U21237 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n18143), .B1(
        n18395), .B2(n18142), .ZN(n18131) );
  AOI22_X1 U21238 ( .A1(n18396), .A2(n18144), .B1(n18397), .B2(n18167), .ZN(
        n18130) );
  OAI211_X1 U21239 ( .C1(n18400), .C2(n18147), .A(n18131), .B(n18130), .ZN(
        P3_U2901) );
  AOI22_X1 U21240 ( .A1(n18402), .A2(n18144), .B1(n18401), .B2(n18142), .ZN(
        n18133) );
  AOI22_X1 U21241 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n18143), .B1(
        n18403), .B2(n18167), .ZN(n18132) );
  OAI211_X1 U21242 ( .C1(n18406), .C2(n18147), .A(n18133), .B(n18132), .ZN(
        P3_U2902) );
  AOI22_X1 U21243 ( .A1(n18409), .A2(n18167), .B1(n18407), .B2(n18142), .ZN(
        n18135) );
  AOI22_X1 U21244 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n18143), .B1(
        n18408), .B2(n18144), .ZN(n18134) );
  OAI211_X1 U21245 ( .C1(n18412), .C2(n18147), .A(n18135), .B(n18134), .ZN(
        P3_U2903) );
  AOI22_X1 U21246 ( .A1(n18414), .A2(n18167), .B1(n18413), .B2(n18142), .ZN(
        n18137) );
  AOI22_X1 U21247 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n18143), .B1(
        n18415), .B2(n18144), .ZN(n18136) );
  OAI211_X1 U21248 ( .C1(n18418), .C2(n18147), .A(n18137), .B(n18136), .ZN(
        P3_U2904) );
  AOI22_X1 U21249 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n18143), .B1(
        n18419), .B2(n18142), .ZN(n18139) );
  AOI22_X1 U21250 ( .A1(n18421), .A2(n18144), .B1(n18420), .B2(n18167), .ZN(
        n18138) );
  OAI211_X1 U21251 ( .C1(n18424), .C2(n18147), .A(n18139), .B(n18138), .ZN(
        P3_U2905) );
  AOI22_X1 U21252 ( .A1(n18427), .A2(n18144), .B1(n18425), .B2(n18142), .ZN(
        n18141) );
  AOI22_X1 U21253 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n18143), .B1(
        n18426), .B2(n18167), .ZN(n18140) );
  OAI211_X1 U21254 ( .C1(n18430), .C2(n18147), .A(n18141), .B(n18140), .ZN(
        P3_U2906) );
  AOI22_X1 U21255 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n18143), .B1(
        n18432), .B2(n18142), .ZN(n18146) );
  AOI22_X1 U21256 ( .A1(n18434), .A2(n18144), .B1(n18435), .B2(n18167), .ZN(
        n18145) );
  OAI211_X1 U21257 ( .C1(n18440), .C2(n18147), .A(n18146), .B(n18145), .ZN(
        P3_U2907) );
  NAND2_X1 U21258 ( .A1(n18238), .A2(n18194), .ZN(n18171) );
  NOR2_X1 U21259 ( .A1(n18239), .A2(n18148), .ZN(n18166) );
  AOI22_X1 U21260 ( .A1(n18386), .A2(n18167), .B1(n18385), .B2(n18166), .ZN(
        n18153) );
  NOR2_X1 U21261 ( .A1(n18288), .A2(n18149), .ZN(n18151) );
  AOI22_X1 U21262 ( .A1(n18390), .A2(n18151), .B1(n18150), .B2(n18194), .ZN(
        n18168) );
  AOI22_X1 U21263 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n18168), .B1(
        n18391), .B2(n18190), .ZN(n18152) );
  OAI211_X1 U21264 ( .C1(n18394), .C2(n18171), .A(n18153), .B(n18152), .ZN(
        P3_U2908) );
  AOI22_X1 U21265 ( .A1(n18395), .A2(n18166), .B1(n18397), .B2(n18190), .ZN(
        n18155) );
  AOI22_X1 U21266 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n18168), .B1(
        n18396), .B2(n18167), .ZN(n18154) );
  OAI211_X1 U21267 ( .C1(n18400), .C2(n18171), .A(n18155), .B(n18154), .ZN(
        P3_U2909) );
  AOI22_X1 U21268 ( .A1(n18403), .A2(n18190), .B1(n18401), .B2(n18166), .ZN(
        n18157) );
  AOI22_X1 U21269 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n18168), .B1(
        n18402), .B2(n18167), .ZN(n18156) );
  OAI211_X1 U21270 ( .C1(n18406), .C2(n18171), .A(n18157), .B(n18156), .ZN(
        P3_U2910) );
  AOI22_X1 U21271 ( .A1(n18408), .A2(n18167), .B1(n18407), .B2(n18166), .ZN(
        n18159) );
  AOI22_X1 U21272 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n18168), .B1(
        n18409), .B2(n18190), .ZN(n18158) );
  OAI211_X1 U21273 ( .C1(n18412), .C2(n18171), .A(n18159), .B(n18158), .ZN(
        P3_U2911) );
  AOI22_X1 U21274 ( .A1(n18414), .A2(n18190), .B1(n18413), .B2(n18166), .ZN(
        n18161) );
  AOI22_X1 U21275 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n18168), .B1(
        n18415), .B2(n18167), .ZN(n18160) );
  OAI211_X1 U21276 ( .C1(n18418), .C2(n18171), .A(n18161), .B(n18160), .ZN(
        P3_U2912) );
  AOI22_X1 U21277 ( .A1(n18421), .A2(n18167), .B1(n18419), .B2(n18166), .ZN(
        n18163) );
  AOI22_X1 U21278 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n18168), .B1(
        n18420), .B2(n18190), .ZN(n18162) );
  OAI211_X1 U21279 ( .C1(n18424), .C2(n18171), .A(n18163), .B(n18162), .ZN(
        P3_U2913) );
  AOI22_X1 U21280 ( .A1(n18426), .A2(n18190), .B1(n18425), .B2(n18166), .ZN(
        n18165) );
  AOI22_X1 U21281 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n18168), .B1(
        n18427), .B2(n18167), .ZN(n18164) );
  OAI211_X1 U21282 ( .C1(n18430), .C2(n18171), .A(n18165), .B(n18164), .ZN(
        P3_U2914) );
  AOI22_X1 U21283 ( .A1(n18434), .A2(n18167), .B1(n18432), .B2(n18166), .ZN(
        n18170) );
  AOI22_X1 U21284 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n18168), .B1(
        n18435), .B2(n18190), .ZN(n18169) );
  OAI211_X1 U21285 ( .C1(n18440), .C2(n18171), .A(n18170), .B(n18169), .ZN(
        P3_U2915) );
  NAND2_X1 U21286 ( .A1(n18263), .A2(n18194), .ZN(n18193) );
  INV_X1 U21287 ( .A(n18171), .ZN(n18234) );
  INV_X1 U21288 ( .A(n18193), .ZN(n18259) );
  NOR2_X1 U21289 ( .A1(n18234), .A2(n18259), .ZN(n18216) );
  NOR2_X1 U21290 ( .A1(n18357), .A2(n18216), .ZN(n18188) );
  AOI22_X1 U21291 ( .A1(n18386), .A2(n18190), .B1(n18385), .B2(n18188), .ZN(
        n18175) );
  OAI21_X1 U21292 ( .B1(n18172), .B2(n18359), .A(n18216), .ZN(n18173) );
  OAI211_X1 U21293 ( .C1(n18259), .C2(n18599), .A(n18362), .B(n18173), .ZN(
        n18189) );
  AOI22_X1 U21294 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n18189), .B1(
        n18391), .B2(n18211), .ZN(n18174) );
  OAI211_X1 U21295 ( .C1(n18394), .C2(n18193), .A(n18175), .B(n18174), .ZN(
        P3_U2916) );
  AOI22_X1 U21296 ( .A1(n18395), .A2(n18188), .B1(n18397), .B2(n18211), .ZN(
        n18177) );
  AOI22_X1 U21297 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n18189), .B1(
        n18396), .B2(n18190), .ZN(n18176) );
  OAI211_X1 U21298 ( .C1(n18400), .C2(n18193), .A(n18177), .B(n18176), .ZN(
        P3_U2917) );
  AOI22_X1 U21299 ( .A1(n18402), .A2(n18190), .B1(n18401), .B2(n18188), .ZN(
        n18179) );
  AOI22_X1 U21300 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n18189), .B1(
        n18403), .B2(n18211), .ZN(n18178) );
  OAI211_X1 U21301 ( .C1(n18406), .C2(n18193), .A(n18179), .B(n18178), .ZN(
        P3_U2918) );
  AOI22_X1 U21302 ( .A1(n18408), .A2(n18190), .B1(n18407), .B2(n18188), .ZN(
        n18181) );
  AOI22_X1 U21303 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n18189), .B1(
        n18409), .B2(n18211), .ZN(n18180) );
  OAI211_X1 U21304 ( .C1(n18412), .C2(n18193), .A(n18181), .B(n18180), .ZN(
        P3_U2919) );
  AOI22_X1 U21305 ( .A1(n18415), .A2(n18190), .B1(n18413), .B2(n18188), .ZN(
        n18183) );
  AOI22_X1 U21306 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n18189), .B1(
        n18414), .B2(n18211), .ZN(n18182) );
  OAI211_X1 U21307 ( .C1(n18418), .C2(n18193), .A(n18183), .B(n18182), .ZN(
        P3_U2920) );
  AOI22_X1 U21308 ( .A1(n18420), .A2(n18211), .B1(n18419), .B2(n18188), .ZN(
        n18185) );
  AOI22_X1 U21309 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n18189), .B1(
        n18421), .B2(n18190), .ZN(n18184) );
  OAI211_X1 U21310 ( .C1(n18424), .C2(n18193), .A(n18185), .B(n18184), .ZN(
        P3_U2921) );
  AOI22_X1 U21311 ( .A1(n18427), .A2(n18190), .B1(n18425), .B2(n18188), .ZN(
        n18187) );
  AOI22_X1 U21312 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n18189), .B1(
        n18426), .B2(n18211), .ZN(n18186) );
  OAI211_X1 U21313 ( .C1(n18430), .C2(n18193), .A(n18187), .B(n18186), .ZN(
        P3_U2922) );
  AOI22_X1 U21314 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n18189), .B1(
        n18432), .B2(n18188), .ZN(n18192) );
  AOI22_X1 U21315 ( .A1(n18434), .A2(n18190), .B1(n18435), .B2(n18211), .ZN(
        n18191) );
  OAI211_X1 U21316 ( .C1(n18440), .C2(n18193), .A(n18192), .B(n18191), .ZN(
        P3_U2923) );
  NAND2_X1 U21317 ( .A1(n18470), .A2(n18194), .ZN(n18215) );
  AOI22_X1 U21318 ( .A1(n18386), .A2(n18211), .B1(n18385), .B2(n18210), .ZN(
        n18197) );
  NAND2_X1 U21319 ( .A1(n18195), .A2(n18194), .ZN(n18212) );
  AOI22_X1 U21320 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n18212), .B1(
        n18391), .B2(n18234), .ZN(n18196) );
  OAI211_X1 U21321 ( .C1(n18394), .C2(n18215), .A(n18197), .B(n18196), .ZN(
        P3_U2924) );
  AOI22_X1 U21322 ( .A1(n18396), .A2(n18211), .B1(n18395), .B2(n18210), .ZN(
        n18199) );
  AOI22_X1 U21323 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n18212), .B1(
        n18397), .B2(n18234), .ZN(n18198) );
  OAI211_X1 U21324 ( .C1(n18400), .C2(n18215), .A(n18199), .B(n18198), .ZN(
        P3_U2925) );
  AOI22_X1 U21325 ( .A1(n18402), .A2(n18211), .B1(n18401), .B2(n18210), .ZN(
        n18201) );
  AOI22_X1 U21326 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n18212), .B1(
        n18403), .B2(n18234), .ZN(n18200) );
  OAI211_X1 U21327 ( .C1(n18406), .C2(n18215), .A(n18201), .B(n18200), .ZN(
        P3_U2926) );
  AOI22_X1 U21328 ( .A1(n18408), .A2(n18211), .B1(n18407), .B2(n18210), .ZN(
        n18203) );
  AOI22_X1 U21329 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n18212), .B1(
        n18409), .B2(n18234), .ZN(n18202) );
  OAI211_X1 U21330 ( .C1(n18412), .C2(n18215), .A(n18203), .B(n18202), .ZN(
        P3_U2927) );
  AOI22_X1 U21331 ( .A1(n18414), .A2(n18234), .B1(n18413), .B2(n18210), .ZN(
        n18205) );
  AOI22_X1 U21332 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n18212), .B1(
        n18415), .B2(n18211), .ZN(n18204) );
  OAI211_X1 U21333 ( .C1(n18418), .C2(n18215), .A(n18205), .B(n18204), .ZN(
        P3_U2928) );
  AOI22_X1 U21334 ( .A1(n18421), .A2(n18211), .B1(n18419), .B2(n18210), .ZN(
        n18207) );
  AOI22_X1 U21335 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n18212), .B1(
        n18420), .B2(n18234), .ZN(n18206) );
  OAI211_X1 U21336 ( .C1(n18424), .C2(n18215), .A(n18207), .B(n18206), .ZN(
        P3_U2929) );
  AOI22_X1 U21337 ( .A1(n18427), .A2(n18211), .B1(n18425), .B2(n18210), .ZN(
        n18209) );
  AOI22_X1 U21338 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n18212), .B1(
        n18426), .B2(n18234), .ZN(n18208) );
  OAI211_X1 U21339 ( .C1(n18430), .C2(n18215), .A(n18209), .B(n18208), .ZN(
        P3_U2930) );
  AOI22_X1 U21340 ( .A1(n18435), .A2(n18234), .B1(n18432), .B2(n18210), .ZN(
        n18214) );
  AOI22_X1 U21341 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n18212), .B1(
        n18434), .B2(n18211), .ZN(n18213) );
  OAI211_X1 U21342 ( .C1(n18440), .C2(n18215), .A(n18214), .B(n18213), .ZN(
        P3_U2931) );
  NAND2_X1 U21343 ( .A1(n18471), .A2(n18289), .ZN(n18237) );
  INV_X1 U21344 ( .A(n18215), .ZN(n18282) );
  INV_X1 U21345 ( .A(n18237), .ZN(n18305) );
  NOR2_X1 U21346 ( .A1(n18282), .A2(n18305), .ZN(n18264) );
  NOR2_X1 U21347 ( .A1(n18357), .A2(n18264), .ZN(n18232) );
  AOI22_X1 U21348 ( .A1(n18386), .A2(n18234), .B1(n18385), .B2(n18232), .ZN(
        n18219) );
  OAI21_X1 U21349 ( .B1(n18216), .B2(n18359), .A(n18264), .ZN(n18217) );
  OAI211_X1 U21350 ( .C1(n18305), .C2(n18599), .A(n18362), .B(n18217), .ZN(
        n18233) );
  AOI22_X1 U21351 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n18233), .B1(
        n18391), .B2(n18259), .ZN(n18218) );
  OAI211_X1 U21352 ( .C1(n18394), .C2(n18237), .A(n18219), .B(n18218), .ZN(
        P3_U2932) );
  AOI22_X1 U21353 ( .A1(n18395), .A2(n18232), .B1(n18397), .B2(n18259), .ZN(
        n18221) );
  AOI22_X1 U21354 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n18233), .B1(
        n18396), .B2(n18234), .ZN(n18220) );
  OAI211_X1 U21355 ( .C1(n18400), .C2(n18237), .A(n18221), .B(n18220), .ZN(
        P3_U2933) );
  AOI22_X1 U21356 ( .A1(n18402), .A2(n18234), .B1(n18401), .B2(n18232), .ZN(
        n18223) );
  AOI22_X1 U21357 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n18233), .B1(
        n18403), .B2(n18259), .ZN(n18222) );
  OAI211_X1 U21358 ( .C1(n18406), .C2(n18237), .A(n18223), .B(n18222), .ZN(
        P3_U2934) );
  AOI22_X1 U21359 ( .A1(n18408), .A2(n18234), .B1(n18407), .B2(n18232), .ZN(
        n18225) );
  AOI22_X1 U21360 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n18233), .B1(
        n18409), .B2(n18259), .ZN(n18224) );
  OAI211_X1 U21361 ( .C1(n18412), .C2(n18237), .A(n18225), .B(n18224), .ZN(
        P3_U2935) );
  AOI22_X1 U21362 ( .A1(n18414), .A2(n18259), .B1(n18413), .B2(n18232), .ZN(
        n18227) );
  AOI22_X1 U21363 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n18233), .B1(
        n18415), .B2(n18234), .ZN(n18226) );
  OAI211_X1 U21364 ( .C1(n18418), .C2(n18237), .A(n18227), .B(n18226), .ZN(
        P3_U2936) );
  AOI22_X1 U21365 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n18233), .B1(
        n18419), .B2(n18232), .ZN(n18229) );
  AOI22_X1 U21366 ( .A1(n18421), .A2(n18234), .B1(n18420), .B2(n18259), .ZN(
        n18228) );
  OAI211_X1 U21367 ( .C1(n18424), .C2(n18237), .A(n18229), .B(n18228), .ZN(
        P3_U2937) );
  AOI22_X1 U21368 ( .A1(n18426), .A2(n18259), .B1(n18425), .B2(n18232), .ZN(
        n18231) );
  AOI22_X1 U21369 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n18233), .B1(
        n18427), .B2(n18234), .ZN(n18230) );
  OAI211_X1 U21370 ( .C1(n18430), .C2(n18237), .A(n18231), .B(n18230), .ZN(
        P3_U2938) );
  AOI22_X1 U21371 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n18233), .B1(
        n18432), .B2(n18232), .ZN(n18236) );
  AOI22_X1 U21372 ( .A1(n18434), .A2(n18234), .B1(n18435), .B2(n18259), .ZN(
        n18235) );
  OAI211_X1 U21373 ( .C1(n18440), .C2(n18237), .A(n18236), .B(n18235), .ZN(
        P3_U2939) );
  NAND2_X1 U21374 ( .A1(n18238), .A2(n18289), .ZN(n18286) );
  INV_X1 U21375 ( .A(n18289), .ZN(n18287) );
  NOR2_X1 U21376 ( .A1(n18239), .A2(n18287), .ZN(n18258) );
  AOI22_X1 U21377 ( .A1(n18391), .A2(n18282), .B1(n18385), .B2(n18258), .ZN(
        n18245) );
  NOR2_X1 U21378 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18240), .ZN(
        n18243) );
  INV_X1 U21379 ( .A(n18241), .ZN(n18388) );
  NOR2_X1 U21380 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18287), .ZN(
        n18242) );
  AOI22_X1 U21381 ( .A1(n18390), .A2(n18243), .B1(n18388), .B2(n18242), .ZN(
        n18260) );
  AOI22_X1 U21382 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n18260), .B1(
        n18386), .B2(n18259), .ZN(n18244) );
  OAI211_X1 U21383 ( .C1(n18394), .C2(n18286), .A(n18245), .B(n18244), .ZN(
        P3_U2940) );
  AOI22_X1 U21384 ( .A1(n18396), .A2(n18259), .B1(n18395), .B2(n18258), .ZN(
        n18247) );
  AOI22_X1 U21385 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n18260), .B1(
        n18397), .B2(n18282), .ZN(n18246) );
  OAI211_X1 U21386 ( .C1(n18400), .C2(n18286), .A(n18247), .B(n18246), .ZN(
        P3_U2941) );
  AOI22_X1 U21387 ( .A1(n18402), .A2(n18259), .B1(n18401), .B2(n18258), .ZN(
        n18249) );
  AOI22_X1 U21388 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n18260), .B1(
        n18403), .B2(n18282), .ZN(n18248) );
  OAI211_X1 U21389 ( .C1(n18406), .C2(n18286), .A(n18249), .B(n18248), .ZN(
        P3_U2942) );
  AOI22_X1 U21390 ( .A1(n18408), .A2(n18259), .B1(n18407), .B2(n18258), .ZN(
        n18251) );
  AOI22_X1 U21391 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n18260), .B1(
        n18409), .B2(n18282), .ZN(n18250) );
  OAI211_X1 U21392 ( .C1(n18412), .C2(n18286), .A(n18251), .B(n18250), .ZN(
        P3_U2943) );
  AOI22_X1 U21393 ( .A1(n18414), .A2(n18282), .B1(n18413), .B2(n18258), .ZN(
        n18253) );
  AOI22_X1 U21394 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n18260), .B1(
        n18415), .B2(n18259), .ZN(n18252) );
  OAI211_X1 U21395 ( .C1(n18418), .C2(n18286), .A(n18253), .B(n18252), .ZN(
        P3_U2944) );
  AOI22_X1 U21396 ( .A1(n18421), .A2(n18259), .B1(n18419), .B2(n18258), .ZN(
        n18255) );
  AOI22_X1 U21397 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n18260), .B1(
        n18420), .B2(n18282), .ZN(n18254) );
  OAI211_X1 U21398 ( .C1(n18424), .C2(n18286), .A(n18255), .B(n18254), .ZN(
        P3_U2945) );
  AOI22_X1 U21399 ( .A1(n18426), .A2(n18282), .B1(n18425), .B2(n18258), .ZN(
        n18257) );
  AOI22_X1 U21400 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n18260), .B1(
        n18427), .B2(n18259), .ZN(n18256) );
  OAI211_X1 U21401 ( .C1(n18430), .C2(n18286), .A(n18257), .B(n18256), .ZN(
        P3_U2946) );
  AOI22_X1 U21402 ( .A1(n18435), .A2(n18282), .B1(n18432), .B2(n18258), .ZN(
        n18262) );
  AOI22_X1 U21403 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n18260), .B1(
        n18434), .B2(n18259), .ZN(n18261) );
  OAI211_X1 U21404 ( .C1(n18440), .C2(n18286), .A(n18262), .B(n18261), .ZN(
        P3_U2947) );
  NAND2_X1 U21405 ( .A1(n18263), .A2(n18289), .ZN(n18285) );
  AOI21_X1 U21406 ( .B1(n18286), .B2(n18285), .A(n18357), .ZN(n18280) );
  AOI22_X1 U21407 ( .A1(n18386), .A2(n18282), .B1(n18385), .B2(n18280), .ZN(
        n18267) );
  INV_X1 U21408 ( .A(n18285), .ZN(n18351) );
  OAI211_X1 U21409 ( .C1(n18264), .C2(n18359), .A(n18286), .B(n18285), .ZN(
        n18265) );
  OAI211_X1 U21410 ( .C1(n18351), .C2(n18599), .A(n18362), .B(n18265), .ZN(
        n18281) );
  AOI22_X1 U21411 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n18281), .B1(
        n18391), .B2(n18305), .ZN(n18266) );
  OAI211_X1 U21412 ( .C1(n18394), .C2(n18285), .A(n18267), .B(n18266), .ZN(
        P3_U2948) );
  AOI22_X1 U21413 ( .A1(n18396), .A2(n18282), .B1(n18395), .B2(n18280), .ZN(
        n18269) );
  AOI22_X1 U21414 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n18281), .B1(
        n18397), .B2(n18305), .ZN(n18268) );
  OAI211_X1 U21415 ( .C1(n18400), .C2(n18285), .A(n18269), .B(n18268), .ZN(
        P3_U2949) );
  AOI22_X1 U21416 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n18281), .B1(
        n18401), .B2(n18280), .ZN(n18271) );
  AOI22_X1 U21417 ( .A1(n18402), .A2(n18282), .B1(n18403), .B2(n18305), .ZN(
        n18270) );
  OAI211_X1 U21418 ( .C1(n18406), .C2(n18285), .A(n18271), .B(n18270), .ZN(
        P3_U2950) );
  AOI22_X1 U21419 ( .A1(n18409), .A2(n18305), .B1(n18407), .B2(n18280), .ZN(
        n18273) );
  AOI22_X1 U21420 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n18281), .B1(
        n18408), .B2(n18282), .ZN(n18272) );
  OAI211_X1 U21421 ( .C1(n18412), .C2(n18285), .A(n18273), .B(n18272), .ZN(
        P3_U2951) );
  AOI22_X1 U21422 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n18281), .B1(
        n18413), .B2(n18280), .ZN(n18275) );
  AOI22_X1 U21423 ( .A1(n18415), .A2(n18282), .B1(n18414), .B2(n18305), .ZN(
        n18274) );
  OAI211_X1 U21424 ( .C1(n18418), .C2(n18285), .A(n18275), .B(n18274), .ZN(
        P3_U2952) );
  AOI22_X1 U21425 ( .A1(n18420), .A2(n18305), .B1(n18419), .B2(n18280), .ZN(
        n18277) );
  AOI22_X1 U21426 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n18281), .B1(
        n18421), .B2(n18282), .ZN(n18276) );
  OAI211_X1 U21427 ( .C1(n18424), .C2(n18285), .A(n18277), .B(n18276), .ZN(
        P3_U2953) );
  AOI22_X1 U21428 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n18281), .B1(
        n18425), .B2(n18280), .ZN(n18279) );
  AOI22_X1 U21429 ( .A1(n18427), .A2(n18282), .B1(n18426), .B2(n18305), .ZN(
        n18278) );
  OAI211_X1 U21430 ( .C1(n18430), .C2(n18285), .A(n18279), .B(n18278), .ZN(
        P3_U2954) );
  AOI22_X1 U21431 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n18281), .B1(
        n18432), .B2(n18280), .ZN(n18284) );
  AOI22_X1 U21432 ( .A1(n18434), .A2(n18282), .B1(n18435), .B2(n18305), .ZN(
        n18283) );
  OAI211_X1 U21433 ( .C1(n18440), .C2(n18285), .A(n18284), .B(n18283), .ZN(
        P3_U2955) );
  NAND2_X1 U21434 ( .A1(n18470), .A2(n18289), .ZN(n18333) );
  INV_X1 U21435 ( .A(n18286), .ZN(n18328) );
  NOR2_X1 U21436 ( .A1(n18288), .A2(n18287), .ZN(n18335) );
  AND2_X1 U21437 ( .A1(n18505), .A2(n18335), .ZN(n18304) );
  AOI22_X1 U21438 ( .A1(n18391), .A2(n18328), .B1(n18385), .B2(n18304), .ZN(
        n18291) );
  OAI211_X1 U21439 ( .C1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .C2(n18390), .A(
        n18388), .B(n18289), .ZN(n18306) );
  AOI22_X1 U21440 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n18306), .B1(
        n18386), .B2(n18305), .ZN(n18290) );
  OAI211_X1 U21441 ( .C1(n18394), .C2(n18333), .A(n18291), .B(n18290), .ZN(
        P3_U2956) );
  AOI22_X1 U21442 ( .A1(n18395), .A2(n18304), .B1(n18397), .B2(n18328), .ZN(
        n18293) );
  AOI22_X1 U21443 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n18306), .B1(
        n18396), .B2(n18305), .ZN(n18292) );
  OAI211_X1 U21444 ( .C1(n18400), .C2(n18333), .A(n18293), .B(n18292), .ZN(
        P3_U2957) );
  AOI22_X1 U21445 ( .A1(n18402), .A2(n18305), .B1(n18401), .B2(n18304), .ZN(
        n18295) );
  AOI22_X1 U21446 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n18306), .B1(
        n18403), .B2(n18328), .ZN(n18294) );
  OAI211_X1 U21447 ( .C1(n18406), .C2(n18333), .A(n18295), .B(n18294), .ZN(
        P3_U2958) );
  AOI22_X1 U21448 ( .A1(n18408), .A2(n18305), .B1(n18407), .B2(n18304), .ZN(
        n18297) );
  AOI22_X1 U21449 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n18306), .B1(
        n18409), .B2(n18328), .ZN(n18296) );
  OAI211_X1 U21450 ( .C1(n18412), .C2(n18333), .A(n18297), .B(n18296), .ZN(
        P3_U2959) );
  AOI22_X1 U21451 ( .A1(n18415), .A2(n18305), .B1(n18413), .B2(n18304), .ZN(
        n18299) );
  AOI22_X1 U21452 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n18306), .B1(
        n18414), .B2(n18328), .ZN(n18298) );
  OAI211_X1 U21453 ( .C1(n18418), .C2(n18333), .A(n18299), .B(n18298), .ZN(
        P3_U2960) );
  AOI22_X1 U21454 ( .A1(n18420), .A2(n18328), .B1(n18419), .B2(n18304), .ZN(
        n18301) );
  AOI22_X1 U21455 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n18306), .B1(
        n18421), .B2(n18305), .ZN(n18300) );
  OAI211_X1 U21456 ( .C1(n18424), .C2(n18333), .A(n18301), .B(n18300), .ZN(
        P3_U2961) );
  AOI22_X1 U21457 ( .A1(n18427), .A2(n18305), .B1(n18425), .B2(n18304), .ZN(
        n18303) );
  AOI22_X1 U21458 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n18306), .B1(
        n18426), .B2(n18328), .ZN(n18302) );
  OAI211_X1 U21459 ( .C1(n18430), .C2(n18333), .A(n18303), .B(n18302), .ZN(
        P3_U2962) );
  AOI22_X1 U21460 ( .A1(n18434), .A2(n18305), .B1(n18432), .B2(n18304), .ZN(
        n18308) );
  AOI22_X1 U21461 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n18306), .B1(
        n18435), .B2(n18328), .ZN(n18307) );
  OAI211_X1 U21462 ( .C1(n18440), .C2(n18333), .A(n18308), .B(n18307), .ZN(
        P3_U2963) );
  INV_X1 U21463 ( .A(n18334), .ZN(n18389) );
  NAND2_X1 U21464 ( .A1(n18389), .A2(n18309), .ZN(n18332) );
  AOI21_X1 U21465 ( .B1(n18333), .B2(n18332), .A(n18357), .ZN(n18327) );
  AOI22_X1 U21466 ( .A1(n18391), .A2(n18351), .B1(n18385), .B2(n18327), .ZN(
        n18314) );
  INV_X1 U21467 ( .A(n18332), .ZN(n18433) );
  AOI221_X1 U21468 ( .B1(n18311), .B2(n18333), .C1(n18310), .C2(n18333), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n18312) );
  OAI21_X1 U21469 ( .B1(n18433), .B2(n18312), .A(n18362), .ZN(n18329) );
  AOI22_X1 U21470 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n18329), .B1(
        n18386), .B2(n18328), .ZN(n18313) );
  OAI211_X1 U21471 ( .C1(n18394), .C2(n18332), .A(n18314), .B(n18313), .ZN(
        P3_U2964) );
  AOI22_X1 U21472 ( .A1(n18395), .A2(n18327), .B1(n18397), .B2(n18351), .ZN(
        n18316) );
  AOI22_X1 U21473 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n18329), .B1(
        n18396), .B2(n18328), .ZN(n18315) );
  OAI211_X1 U21474 ( .C1(n18400), .C2(n18332), .A(n18316), .B(n18315), .ZN(
        P3_U2965) );
  AOI22_X1 U21475 ( .A1(n18403), .A2(n18351), .B1(n18401), .B2(n18327), .ZN(
        n18318) );
  AOI22_X1 U21476 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n18329), .B1(
        n18402), .B2(n18328), .ZN(n18317) );
  OAI211_X1 U21477 ( .C1(n18406), .C2(n18332), .A(n18318), .B(n18317), .ZN(
        P3_U2966) );
  AOI22_X1 U21478 ( .A1(n18409), .A2(n18351), .B1(n18407), .B2(n18327), .ZN(
        n18320) );
  AOI22_X1 U21479 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n18329), .B1(
        n18408), .B2(n18328), .ZN(n18319) );
  OAI211_X1 U21480 ( .C1(n18412), .C2(n18332), .A(n18320), .B(n18319), .ZN(
        P3_U2967) );
  AOI22_X1 U21481 ( .A1(n18414), .A2(n18351), .B1(n18413), .B2(n18327), .ZN(
        n18322) );
  AOI22_X1 U21482 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n18329), .B1(
        n18415), .B2(n18328), .ZN(n18321) );
  OAI211_X1 U21483 ( .C1(n18418), .C2(n18332), .A(n18322), .B(n18321), .ZN(
        P3_U2968) );
  AOI22_X1 U21484 ( .A1(n18421), .A2(n18328), .B1(n18419), .B2(n18327), .ZN(
        n18324) );
  AOI22_X1 U21485 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n18329), .B1(
        n18420), .B2(n18351), .ZN(n18323) );
  OAI211_X1 U21486 ( .C1(n18424), .C2(n18332), .A(n18324), .B(n18323), .ZN(
        P3_U2969) );
  AOI22_X1 U21487 ( .A1(n18426), .A2(n18351), .B1(n18425), .B2(n18327), .ZN(
        n18326) );
  AOI22_X1 U21488 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n18329), .B1(
        n18427), .B2(n18328), .ZN(n18325) );
  OAI211_X1 U21489 ( .C1(n18430), .C2(n18332), .A(n18326), .B(n18325), .ZN(
        P3_U2970) );
  AOI22_X1 U21490 ( .A1(n18434), .A2(n18328), .B1(n18432), .B2(n18327), .ZN(
        n18331) );
  AOI22_X1 U21491 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n18329), .B1(
        n18435), .B2(n18351), .ZN(n18330) );
  OAI211_X1 U21492 ( .C1(n18440), .C2(n18332), .A(n18331), .B(n18330), .ZN(
        P3_U2971) );
  INV_X1 U21493 ( .A(n18436), .ZN(n18355) );
  INV_X1 U21494 ( .A(n18333), .ZN(n18379) );
  NOR2_X1 U21495 ( .A1(n18357), .A2(n18334), .ZN(n18350) );
  AOI22_X1 U21496 ( .A1(n18391), .A2(n18379), .B1(n18385), .B2(n18350), .ZN(
        n18337) );
  AOI22_X1 U21497 ( .A1(n18390), .A2(n18335), .B1(n18389), .B2(n18388), .ZN(
        n18352) );
  AOI22_X1 U21498 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n18352), .B1(
        n18386), .B2(n18351), .ZN(n18336) );
  OAI211_X1 U21499 ( .C1(n18394), .C2(n18355), .A(n18337), .B(n18336), .ZN(
        P3_U2972) );
  AOI22_X1 U21500 ( .A1(n18395), .A2(n18350), .B1(n18397), .B2(n18379), .ZN(
        n18339) );
  AOI22_X1 U21501 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n18352), .B1(
        n18396), .B2(n18351), .ZN(n18338) );
  OAI211_X1 U21502 ( .C1(n18355), .C2(n18400), .A(n18339), .B(n18338), .ZN(
        P3_U2973) );
  AOI22_X1 U21503 ( .A1(n18403), .A2(n18379), .B1(n18401), .B2(n18350), .ZN(
        n18341) );
  AOI22_X1 U21504 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n18352), .B1(
        n18402), .B2(n18351), .ZN(n18340) );
  OAI211_X1 U21505 ( .C1(n18355), .C2(n18406), .A(n18341), .B(n18340), .ZN(
        P3_U2974) );
  AOI22_X1 U21506 ( .A1(n18408), .A2(n18351), .B1(n18407), .B2(n18350), .ZN(
        n18343) );
  AOI22_X1 U21507 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n18352), .B1(
        n18409), .B2(n18379), .ZN(n18342) );
  OAI211_X1 U21508 ( .C1(n18355), .C2(n18412), .A(n18343), .B(n18342), .ZN(
        P3_U2975) );
  AOI22_X1 U21509 ( .A1(n18415), .A2(n18351), .B1(n18413), .B2(n18350), .ZN(
        n18345) );
  AOI22_X1 U21510 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n18352), .B1(
        n18414), .B2(n18379), .ZN(n18344) );
  OAI211_X1 U21511 ( .C1(n18355), .C2(n18418), .A(n18345), .B(n18344), .ZN(
        P3_U2976) );
  AOI22_X1 U21512 ( .A1(n18420), .A2(n18379), .B1(n18419), .B2(n18350), .ZN(
        n18347) );
  AOI22_X1 U21513 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n18352), .B1(
        n18421), .B2(n18351), .ZN(n18346) );
  OAI211_X1 U21514 ( .C1(n18355), .C2(n18424), .A(n18347), .B(n18346), .ZN(
        P3_U2977) );
  AOI22_X1 U21515 ( .A1(n18427), .A2(n18351), .B1(n18425), .B2(n18350), .ZN(
        n18349) );
  AOI22_X1 U21516 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n18352), .B1(
        n18426), .B2(n18379), .ZN(n18348) );
  OAI211_X1 U21517 ( .C1(n18355), .C2(n18430), .A(n18349), .B(n18348), .ZN(
        P3_U2978) );
  AOI22_X1 U21518 ( .A1(n18434), .A2(n18351), .B1(n18432), .B2(n18350), .ZN(
        n18354) );
  AOI22_X1 U21519 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n18352), .B1(
        n18435), .B2(n18379), .ZN(n18353) );
  OAI211_X1 U21520 ( .C1(n18355), .C2(n18440), .A(n18354), .B(n18353), .ZN(
        P3_U2979) );
  INV_X1 U21521 ( .A(n18363), .ZN(n18383) );
  INV_X1 U21522 ( .A(n18356), .ZN(n18358) );
  NOR2_X1 U21523 ( .A1(n18357), .A2(n18358), .ZN(n18378) );
  AOI22_X1 U21524 ( .A1(n18386), .A2(n18379), .B1(n18385), .B2(n18378), .ZN(
        n18365) );
  NOR2_X1 U21525 ( .A1(n18379), .A2(n18433), .ZN(n18360) );
  OAI21_X1 U21526 ( .B1(n18360), .B2(n18359), .A(n18358), .ZN(n18361) );
  OAI211_X1 U21527 ( .C1(n18363), .C2(n18599), .A(n18362), .B(n18361), .ZN(
        n18380) );
  AOI22_X1 U21528 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n18380), .B1(
        n18391), .B2(n18433), .ZN(n18364) );
  OAI211_X1 U21529 ( .C1(n18383), .C2(n18394), .A(n18365), .B(n18364), .ZN(
        P3_U2980) );
  AOI22_X1 U21530 ( .A1(n18395), .A2(n18378), .B1(n18397), .B2(n18433), .ZN(
        n18367) );
  AOI22_X1 U21531 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n18380), .B1(
        n18396), .B2(n18379), .ZN(n18366) );
  OAI211_X1 U21532 ( .C1(n18383), .C2(n18400), .A(n18367), .B(n18366), .ZN(
        P3_U2981) );
  AOI22_X1 U21533 ( .A1(n18403), .A2(n18433), .B1(n18401), .B2(n18378), .ZN(
        n18369) );
  AOI22_X1 U21534 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n18380), .B1(
        n18402), .B2(n18379), .ZN(n18368) );
  OAI211_X1 U21535 ( .C1(n18383), .C2(n18406), .A(n18369), .B(n18368), .ZN(
        P3_U2982) );
  AOI22_X1 U21536 ( .A1(n18408), .A2(n18379), .B1(n18407), .B2(n18378), .ZN(
        n18371) );
  AOI22_X1 U21537 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n18380), .B1(
        n18409), .B2(n18433), .ZN(n18370) );
  OAI211_X1 U21538 ( .C1(n18383), .C2(n18412), .A(n18371), .B(n18370), .ZN(
        P3_U2983) );
  AOI22_X1 U21539 ( .A1(n18414), .A2(n18433), .B1(n18413), .B2(n18378), .ZN(
        n18373) );
  AOI22_X1 U21540 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n18380), .B1(
        n18415), .B2(n18379), .ZN(n18372) );
  OAI211_X1 U21541 ( .C1(n18383), .C2(n18418), .A(n18373), .B(n18372), .ZN(
        P3_U2984) );
  AOI22_X1 U21542 ( .A1(n18421), .A2(n18379), .B1(n18419), .B2(n18378), .ZN(
        n18375) );
  AOI22_X1 U21543 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n18380), .B1(
        n18420), .B2(n18433), .ZN(n18374) );
  OAI211_X1 U21544 ( .C1(n18383), .C2(n18424), .A(n18375), .B(n18374), .ZN(
        P3_U2985) );
  AOI22_X1 U21545 ( .A1(n18426), .A2(n18433), .B1(n18425), .B2(n18378), .ZN(
        n18377) );
  AOI22_X1 U21546 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n18380), .B1(
        n18427), .B2(n18379), .ZN(n18376) );
  OAI211_X1 U21547 ( .C1(n18383), .C2(n18430), .A(n18377), .B(n18376), .ZN(
        P3_U2986) );
  AOI22_X1 U21548 ( .A1(n18435), .A2(n18433), .B1(n18432), .B2(n18378), .ZN(
        n18382) );
  AOI22_X1 U21549 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n18380), .B1(
        n18434), .B2(n18379), .ZN(n18381) );
  OAI211_X1 U21550 ( .C1(n18383), .C2(n18440), .A(n18382), .B(n18381), .ZN(
        P3_U2987) );
  INV_X1 U21551 ( .A(n18384), .ZN(n18441) );
  AND2_X1 U21552 ( .A1(n18505), .A2(n18387), .ZN(n18431) );
  AOI22_X1 U21553 ( .A1(n18386), .A2(n18433), .B1(n18385), .B2(n18431), .ZN(
        n18393) );
  AOI22_X1 U21554 ( .A1(n18390), .A2(n18389), .B1(n18388), .B2(n18387), .ZN(
        n18437) );
  AOI22_X1 U21555 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n18437), .B1(
        n18391), .B2(n18436), .ZN(n18392) );
  OAI211_X1 U21556 ( .C1(n18441), .C2(n18394), .A(n18393), .B(n18392), .ZN(
        P3_U2988) );
  AOI22_X1 U21557 ( .A1(n18396), .A2(n18433), .B1(n18395), .B2(n18431), .ZN(
        n18399) );
  AOI22_X1 U21558 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n18437), .B1(
        n18436), .B2(n18397), .ZN(n18398) );
  OAI211_X1 U21559 ( .C1(n18441), .C2(n18400), .A(n18399), .B(n18398), .ZN(
        P3_U2989) );
  AOI22_X1 U21560 ( .A1(n18402), .A2(n18433), .B1(n18401), .B2(n18431), .ZN(
        n18405) );
  AOI22_X1 U21561 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n18437), .B1(
        n18436), .B2(n18403), .ZN(n18404) );
  OAI211_X1 U21562 ( .C1(n18441), .C2(n18406), .A(n18405), .B(n18404), .ZN(
        P3_U2990) );
  AOI22_X1 U21563 ( .A1(n18408), .A2(n18433), .B1(n18407), .B2(n18431), .ZN(
        n18411) );
  AOI22_X1 U21564 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n18437), .B1(
        n18436), .B2(n18409), .ZN(n18410) );
  OAI211_X1 U21565 ( .C1(n18441), .C2(n18412), .A(n18411), .B(n18410), .ZN(
        P3_U2991) );
  AOI22_X1 U21566 ( .A1(n18436), .A2(n18414), .B1(n18413), .B2(n18431), .ZN(
        n18417) );
  AOI22_X1 U21567 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n18437), .B1(
        n18415), .B2(n18433), .ZN(n18416) );
  OAI211_X1 U21568 ( .C1(n18441), .C2(n18418), .A(n18417), .B(n18416), .ZN(
        P3_U2992) );
  AOI22_X1 U21569 ( .A1(n18436), .A2(n18420), .B1(n18419), .B2(n18431), .ZN(
        n18423) );
  AOI22_X1 U21570 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n18437), .B1(
        n18421), .B2(n18433), .ZN(n18422) );
  OAI211_X1 U21571 ( .C1(n18441), .C2(n18424), .A(n18423), .B(n18422), .ZN(
        P3_U2993) );
  AOI22_X1 U21572 ( .A1(n18436), .A2(n18426), .B1(n18425), .B2(n18431), .ZN(
        n18429) );
  AOI22_X1 U21573 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n18437), .B1(
        n18427), .B2(n18433), .ZN(n18428) );
  OAI211_X1 U21574 ( .C1(n18441), .C2(n18430), .A(n18429), .B(n18428), .ZN(
        P3_U2994) );
  AOI22_X1 U21575 ( .A1(n18434), .A2(n18433), .B1(n18432), .B2(n18431), .ZN(
        n18439) );
  AOI22_X1 U21576 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n18437), .B1(
        n18436), .B2(n18435), .ZN(n18438) );
  OAI211_X1 U21577 ( .C1(n18441), .C2(n18440), .A(n18439), .B(n18438), .ZN(
        P3_U2995) );
  OAI22_X1 U21578 ( .A1(n18445), .A2(n18444), .B1(n18443), .B2(n18442), .ZN(
        n18446) );
  AOI211_X1 U21579 ( .C1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .C2(n18483), .A(
        n18451), .B(n18450), .ZN(n18494) );
  AOI21_X1 U21580 ( .B1(n18454), .B2(n18453), .A(n18452), .ZN(n18476) );
  NAND2_X1 U21581 ( .A1(n18469), .A2(n18460), .ZN(n18456) );
  OAI211_X1 U21582 ( .C1(n18457), .C2(n18476), .A(n18456), .B(n18455), .ZN(
        n18606) );
  NOR2_X1 U21583 ( .A1(n18483), .A2(n18606), .ZN(n18463) );
  OAI21_X1 U21584 ( .B1(n18465), .B2(n18630), .A(n18458), .ZN(n18474) );
  NOR2_X1 U21585 ( .A1(n18459), .A2(n18474), .ZN(n18466) );
  OAI22_X1 U21586 ( .A1(n18461), .A2(n18481), .B1(n18466), .B2(n18460), .ZN(
        n18603) );
  NAND2_X1 U21587 ( .A1(n18607), .A2(n18603), .ZN(n18462) );
  OAI22_X1 U21588 ( .A1(n18463), .A2(n18607), .B1(n18483), .B2(n18462), .ZN(
        n18490) );
  NAND2_X1 U21589 ( .A1(n18465), .A2(n18464), .ZN(n18468) );
  INV_X1 U21590 ( .A(n18466), .ZN(n18467) );
  AOI22_X1 U21591 ( .A1(n18621), .A2(n18468), .B1(n18624), .B2(n18467), .ZN(
        n18618) );
  AOI22_X1 U21592 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18469), .B1(
        n18468), .B2(n18630), .ZN(n18625) );
  AOI222_X1 U21593 ( .A1(n18618), .A2(n18625), .B1(n18618), .B2(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .C1(n18625), .C2(n18470), .ZN(
        n18472) );
  INV_X1 U21594 ( .A(n18483), .ZN(n18482) );
  AOI21_X1 U21595 ( .B1(n18472), .B2(n18482), .A(n18471), .ZN(n18485) );
  NAND2_X1 U21596 ( .A1(n18624), .A2(n18617), .ZN(n18473) );
  OAI221_X1 U21597 ( .B1(n18624), .B2(n18617), .C1(n18475), .C2(n18474), .A(
        n18473), .ZN(n18480) );
  INV_X1 U21598 ( .A(n18476), .ZN(n18477) );
  NAND3_X1 U21599 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n18478), .A3(
        n18477), .ZN(n18479) );
  OAI211_X1 U21600 ( .C1(n18613), .C2(n18481), .A(n18480), .B(n18479), .ZN(
        n18615) );
  AOI22_X1 U21601 ( .A1(n18483), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n18615), .B2(n18482), .ZN(n18486) );
  OR2_X1 U21602 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18486), .ZN(
        n18484) );
  AOI221_X1 U21603 ( .B1(n18485), .B2(n18484), .C1(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .C2(n18486), .A(
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n18489) );
  OAI21_X1 U21604 ( .B1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(n18486), .ZN(n18488) );
  AOI222_X1 U21605 ( .A1(n18490), .A2(n18489), .B1(n18490), .B2(n18488), .C1(
        n18489), .C2(n18487), .ZN(n18493) );
  OAI21_X1 U21606 ( .B1(P3_MORE_REG_SCAN_IN), .B2(P3_FLUSH_REG_SCAN_IN), .A(
        n18491), .ZN(n18492) );
  NAND4_X1 U21607 ( .A1(n18645), .A2(n18494), .A3(n18493), .A4(n18492), .ZN(
        n18500) );
  AOI211_X1 U21608 ( .C1(n18497), .C2(n18496), .A(n18495), .B(n18500), .ZN(
        n18597) );
  AOI21_X1 U21609 ( .B1(n18650), .B2(n18666), .A(n18597), .ZN(n18506) );
  NOR2_X1 U21610 ( .A1(n18655), .A2(n18649), .ZN(n18503) );
  AOI211_X1 U21611 ( .C1(n18626), .C2(n18658), .A(P3_STATE2_REG_0__SCAN_IN), 
        .B(n18503), .ZN(n18498) );
  AOI211_X1 U21612 ( .C1(n18648), .C2(n18500), .A(n18499), .B(n18498), .ZN(
        n18501) );
  OAI221_X1 U21613 ( .B1(n18596), .B2(n18506), .C1(n18596), .C2(n18502), .A(
        n18501), .ZN(P3_U2996) );
  INV_X1 U21614 ( .A(n18503), .ZN(n18509) );
  NAND4_X1 U21615 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(
        P3_STATE2_REG_1__SCAN_IN), .A3(n18650), .A4(n18666), .ZN(n18511) );
  INV_X1 U21616 ( .A(n18504), .ZN(n18507) );
  NAND3_X1 U21617 ( .A1(n18507), .A2(n18506), .A3(n18505), .ZN(n18508) );
  NAND4_X1 U21618 ( .A1(n9780), .A2(n18509), .A3(n18511), .A4(n18508), .ZN(
        P3_U2997) );
  OAI21_X1 U21619 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(
        P3_STATEBS16_REG_SCAN_IN), .A(n18510), .ZN(n18513) );
  INV_X1 U21620 ( .A(n18511), .ZN(n18512) );
  AOI21_X1 U21621 ( .B1(n18514), .B2(n18513), .A(n18512), .ZN(P3_U2998) );
  INV_X1 U21622 ( .A(P3_DATAWIDTH_REG_31__SCAN_IN), .ZN(n20854) );
  NOR2_X1 U21623 ( .A1(n18595), .A2(n20854), .ZN(P3_U2999) );
  AND2_X1 U21624 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n18516), .ZN(
        P3_U3000) );
  AND2_X1 U21625 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n18516), .ZN(
        P3_U3001) );
  AND2_X1 U21626 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n18516), .ZN(
        P3_U3002) );
  AND2_X1 U21627 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n18516), .ZN(
        P3_U3003) );
  AND2_X1 U21628 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n18516), .ZN(
        P3_U3004) );
  AND2_X1 U21629 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n18516), .ZN(
        P3_U3005) );
  INV_X1 U21630 ( .A(P3_DATAWIDTH_REG_24__SCAN_IN), .ZN(n20915) );
  NOR2_X1 U21631 ( .A1(n18595), .A2(n20915), .ZN(P3_U3006) );
  AND2_X1 U21632 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n18516), .ZN(
        P3_U3007) );
  AND2_X1 U21633 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n18516), .ZN(
        P3_U3008) );
  AND2_X1 U21634 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n18516), .ZN(
        P3_U3009) );
  AND2_X1 U21635 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n18516), .ZN(
        P3_U3010) );
  AND2_X1 U21636 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n18516), .ZN(
        P3_U3011) );
  AND2_X1 U21637 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n18516), .ZN(
        P3_U3012) );
  AND2_X1 U21638 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n18516), .ZN(
        P3_U3013) );
  AND2_X1 U21639 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n18516), .ZN(
        P3_U3014) );
  INV_X1 U21640 ( .A(P3_DATAWIDTH_REG_15__SCAN_IN), .ZN(n20789) );
  NOR2_X1 U21641 ( .A1(n18595), .A2(n20789), .ZN(P3_U3015) );
  AND2_X1 U21642 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n18516), .ZN(
        P3_U3016) );
  AND2_X1 U21643 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n18515), .ZN(
        P3_U3017) );
  AND2_X1 U21644 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n18515), .ZN(
        P3_U3018) );
  AND2_X1 U21645 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n18515), .ZN(
        P3_U3019) );
  AND2_X1 U21646 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n18515), .ZN(
        P3_U3020) );
  AND2_X1 U21647 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n18515), .ZN(P3_U3021) );
  AND2_X1 U21648 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n18515), .ZN(P3_U3022) );
  AND2_X1 U21649 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n18515), .ZN(P3_U3023) );
  AND2_X1 U21650 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n18515), .ZN(P3_U3024) );
  AND2_X1 U21651 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n18515), .ZN(P3_U3025) );
  AND2_X1 U21652 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n18516), .ZN(P3_U3026) );
  AND2_X1 U21653 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n18516), .ZN(P3_U3027) );
  AND2_X1 U21654 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n18516), .ZN(P3_U3028) );
  OAI21_X1 U21655 ( .B1(n20581), .B2(n18517), .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n18518) );
  INV_X1 U21656 ( .A(n18518), .ZN(n18521) );
  NOR2_X1 U21657 ( .A1(n18655), .A2(n20812), .ZN(n18524) );
  NOR2_X1 U21658 ( .A1(n18524), .A2(n18519), .ZN(n18526) );
  INV_X1 U21659 ( .A(NA), .ZN(n20589) );
  OAI21_X1 U21660 ( .B1(P3_STATE_REG_1__SCAN_IN), .B2(n20589), .A(
        P3_STATE_REG_2__SCAN_IN), .ZN(n18525) );
  INV_X1 U21661 ( .A(n18525), .ZN(n18520) );
  OAI22_X1 U21662 ( .A1(n18665), .A2(n18521), .B1(n18526), .B2(n18520), .ZN(
        P3_U3029) );
  OAI22_X1 U21663 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(
        P3_REQUESTPENDING_REG_SCAN_IN), .B1(n20947), .B2(n20581), .ZN(n18523)
         );
  OAI21_X1 U21664 ( .B1(P3_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .A(
        P3_STATE_REG_0__SCAN_IN), .ZN(n18527) );
  INV_X1 U21665 ( .A(n18524), .ZN(n18522) );
  OAI211_X1 U21666 ( .C1(n18523), .C2(n18527), .A(n18652), .B(n18522), .ZN(
        P3_U3030) );
  AOI21_X1 U21667 ( .B1(n18524), .B2(n20589), .A(n18523), .ZN(n18528) );
  OAI22_X1 U21668 ( .A1(n18528), .A2(n18527), .B1(n18526), .B2(n18525), .ZN(
        P3_U3031) );
  OAI222_X1 U21669 ( .A1(n18582), .A2(n20867), .B1(n18530), .B2(n18665), .C1(
        n18529), .C2(n18579), .ZN(P3_U3032) );
  OAI222_X1 U21670 ( .A1(n18582), .A2(n18532), .B1(n18531), .B2(n18665), .C1(
        n20867), .C2(n18579), .ZN(P3_U3033) );
  INV_X1 U21671 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n18534) );
  OAI222_X1 U21672 ( .A1(n18582), .A2(n18534), .B1(n18533), .B2(n18665), .C1(
        n18532), .C2(n18579), .ZN(P3_U3034) );
  OAI222_X1 U21673 ( .A1(n18582), .A2(n18535), .B1(n20803), .B2(n18665), .C1(
        n18534), .C2(n18579), .ZN(P3_U3035) );
  OAI222_X1 U21674 ( .A1(n18582), .A2(n18537), .B1(n18536), .B2(n18584), .C1(
        n18535), .C2(n18579), .ZN(P3_U3036) );
  OAI222_X1 U21675 ( .A1(n18582), .A2(n18539), .B1(n18538), .B2(n18584), .C1(
        n18537), .C2(n18579), .ZN(P3_U3037) );
  INV_X1 U21676 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n18542) );
  OAI222_X1 U21677 ( .A1(n18582), .A2(n18542), .B1(n18540), .B2(n18665), .C1(
        n18539), .C2(n18579), .ZN(P3_U3038) );
  OAI222_X1 U21678 ( .A1(n18542), .A2(n18579), .B1(n18541), .B2(n18584), .C1(
        n18543), .C2(n18582), .ZN(P3_U3039) );
  OAI222_X1 U21679 ( .A1(n18582), .A2(n18544), .B1(n20948), .B2(n18665), .C1(
        n18543), .C2(n18579), .ZN(P3_U3040) );
  OAI222_X1 U21680 ( .A1(n18582), .A2(n18545), .B1(n20869), .B2(n18665), .C1(
        n18544), .C2(n18579), .ZN(P3_U3041) );
  OAI222_X1 U21681 ( .A1(n18582), .A2(n18547), .B1(n18546), .B2(n18665), .C1(
        n18545), .C2(n18587), .ZN(P3_U3042) );
  OAI222_X1 U21682 ( .A1(n18582), .A2(n18549), .B1(n18548), .B2(n18665), .C1(
        n18547), .C2(n18587), .ZN(P3_U3043) );
  OAI222_X1 U21683 ( .A1(n18582), .A2(n18552), .B1(n18550), .B2(n18665), .C1(
        n18549), .C2(n18587), .ZN(P3_U3044) );
  OAI222_X1 U21684 ( .A1(n18552), .A2(n18579), .B1(n18551), .B2(n18665), .C1(
        n18553), .C2(n18582), .ZN(P3_U3045) );
  OAI222_X1 U21685 ( .A1(n18582), .A2(n18555), .B1(n18554), .B2(n18665), .C1(
        n18553), .C2(n18587), .ZN(P3_U3046) );
  OAI222_X1 U21686 ( .A1(n18582), .A2(n18558), .B1(n18556), .B2(n18665), .C1(
        n18555), .C2(n18587), .ZN(P3_U3047) );
  OAI222_X1 U21687 ( .A1(n18558), .A2(n18579), .B1(n18557), .B2(n18665), .C1(
        n18559), .C2(n18582), .ZN(P3_U3048) );
  OAI222_X1 U21688 ( .A1(n18582), .A2(n18561), .B1(n18560), .B2(n18665), .C1(
        n18559), .C2(n18587), .ZN(P3_U3049) );
  OAI222_X1 U21689 ( .A1(n18582), .A2(n18564), .B1(n18562), .B2(n18665), .C1(
        n18561), .C2(n18587), .ZN(P3_U3050) );
  OAI222_X1 U21690 ( .A1(n18564), .A2(n18579), .B1(n18563), .B2(n18665), .C1(
        n18565), .C2(n18582), .ZN(P3_U3051) );
  OAI222_X1 U21691 ( .A1(n18582), .A2(n18567), .B1(n18566), .B2(n18665), .C1(
        n18565), .C2(n18579), .ZN(P3_U3052) );
  OAI222_X1 U21692 ( .A1(n18582), .A2(n18570), .B1(n18568), .B2(n18665), .C1(
        n18567), .C2(n18587), .ZN(P3_U3053) );
  OAI222_X1 U21693 ( .A1(n18570), .A2(n18579), .B1(n18569), .B2(n18665), .C1(
        n18571), .C2(n18582), .ZN(P3_U3054) );
  OAI222_X1 U21694 ( .A1(n18571), .A2(n18579), .B1(n20797), .B2(n18584), .C1(
        n20927), .C2(n18582), .ZN(P3_U3055) );
  INV_X1 U21695 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n18573) );
  OAI222_X1 U21696 ( .A1(n18582), .A2(n18573), .B1(n18572), .B2(n18584), .C1(
        n20927), .C2(n18587), .ZN(P3_U3056) );
  OAI222_X1 U21697 ( .A1(n18582), .A2(n18575), .B1(n18574), .B2(n18584), .C1(
        n18573), .C2(n18579), .ZN(P3_U3057) );
  OAI222_X1 U21698 ( .A1(n18582), .A2(n18578), .B1(n18576), .B2(n18584), .C1(
        n18575), .C2(n18587), .ZN(P3_U3058) );
  OAI222_X1 U21699 ( .A1(n18578), .A2(n18579), .B1(n18577), .B2(n18584), .C1(
        n18580), .C2(n18582), .ZN(P3_U3059) );
  OAI222_X1 U21700 ( .A1(n18582), .A2(n18586), .B1(n18581), .B2(n18584), .C1(
        n18580), .C2(n18579), .ZN(P3_U3060) );
  INV_X1 U21701 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n18585) );
  OAI222_X1 U21702 ( .A1(n18587), .A2(n18586), .B1(n18585), .B2(n18584), .C1(
        n18583), .C2(n18582), .ZN(P3_U3061) );
  INV_X1 U21703 ( .A(P3_BE_N_REG_3__SCAN_IN), .ZN(n18588) );
  AOI22_X1 U21704 ( .A1(n18665), .A2(n18589), .B1(n18588), .B2(n18663), .ZN(
        P3_U3274) );
  INV_X1 U21705 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n18590) );
  INV_X1 U21706 ( .A(P3_BE_N_REG_2__SCAN_IN), .ZN(n20870) );
  AOI22_X1 U21707 ( .A1(n18665), .A2(n18590), .B1(n20870), .B2(n18663), .ZN(
        P3_U3275) );
  INV_X1 U21708 ( .A(P3_BE_N_REG_1__SCAN_IN), .ZN(n18591) );
  AOI22_X1 U21709 ( .A1(n18665), .A2(n18592), .B1(n18591), .B2(n18663), .ZN(
        P3_U3276) );
  MUX2_X1 U21710 ( .A(P3_BE_N_REG_0__SCAN_IN), .B(P3_BYTEENABLE_REG_0__SCAN_IN), .S(n18665), .Z(P3_U3277) );
  OAI21_X1 U21711 ( .B1(P3_DATAWIDTH_REG_0__SCAN_IN), .B2(n18595), .A(n18594), 
        .ZN(n18593) );
  INV_X1 U21712 ( .A(n18593), .ZN(P3_U3280) );
  OAI21_X1 U21713 ( .B1(n18595), .B2(n20950), .A(n18594), .ZN(P3_U3281) );
  NOR2_X1 U21714 ( .A1(n18597), .A2(n18596), .ZN(n18600) );
  OAI21_X1 U21715 ( .B1(n18600), .B2(n18599), .A(n18598), .ZN(P3_U3282) );
  INV_X1 U21716 ( .A(n18628), .ZN(n18631) );
  INV_X1 U21717 ( .A(n18601), .ZN(n18605) );
  NOR2_X1 U21718 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n18602), .ZN(
        n18604) );
  AOI22_X1 U21719 ( .A1(n18626), .A2(n18605), .B1(n18604), .B2(n18603), .ZN(
        n18609) );
  AOI21_X1 U21720 ( .B1(n18667), .B2(n18606), .A(n18631), .ZN(n18608) );
  OAI22_X1 U21721 ( .A1(n18631), .A2(n18609), .B1(n18608), .B2(n18607), .ZN(
        P3_U3285) );
  NOR2_X1 U21722 ( .A1(n18610), .A2(n20755), .ZN(n18619) );
  AOI22_X1 U21723 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n18612), .B1(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n18611), .ZN(n18620) );
  INV_X1 U21724 ( .A(n18620), .ZN(n18614) );
  AOI222_X1 U21725 ( .A1(n18615), .A2(n18667), .B1(n18619), .B2(n18614), .C1(
        n18626), .C2(n18613), .ZN(n18616) );
  AOI22_X1 U21726 ( .A1(n18631), .A2(n18617), .B1(n18616), .B2(n18628), .ZN(
        P3_U3288) );
  INV_X1 U21727 ( .A(n18618), .ZN(n18622) );
  AOI222_X1 U21728 ( .A1(n18622), .A2(n18667), .B1(n18626), .B2(n18621), .C1(
        n18620), .C2(n18619), .ZN(n18623) );
  AOI22_X1 U21729 ( .A1(n18631), .A2(n18624), .B1(n18623), .B2(n18628), .ZN(
        P3_U3289) );
  INV_X1 U21730 ( .A(n18625), .ZN(n18627) );
  AOI222_X1 U21731 ( .A1(n20755), .A2(P3_STATE2_REG_1__SCAN_IN), .B1(n18667), 
        .B2(n18627), .C1(n18630), .C2(n18626), .ZN(n18629) );
  AOI22_X1 U21732 ( .A1(n18631), .A2(n18630), .B1(n18629), .B2(n18628), .ZN(
        P3_U3290) );
  NAND2_X1 U21733 ( .A1(n18632), .A2(n18633), .ZN(n18639) );
  NOR2_X1 U21734 ( .A1(n18635), .A2(n18633), .ZN(n18634) );
  AOI22_X1 U21735 ( .A1(P3_BYTEENABLE_REG_2__SCAN_IN), .A2(n18635), .B1(
        P3_REIP_REG_1__SCAN_IN), .B2(n18634), .ZN(n18636) );
  OAI221_X1 U21736 ( .B1(P3_DATAWIDTH_REG_0__SCAN_IN), .B2(n18638), .C1(n18637), .C2(n18639), .A(n18636), .ZN(P3_U3292) );
  OAI21_X1 U21737 ( .B1(n18640), .B2(P3_BYTEENABLE_REG_0__SCAN_IN), .A(n18639), 
        .ZN(n18641) );
  INV_X1 U21738 ( .A(n18641), .ZN(P3_U3293) );
  INV_X1 U21739 ( .A(P3_W_R_N_REG_SCAN_IN), .ZN(n18642) );
  AOI22_X1 U21740 ( .A1(n18665), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n18642), 
        .B2(n18663), .ZN(P3_U3294) );
  INV_X1 U21741 ( .A(n18643), .ZN(n18646) );
  NAND2_X1 U21742 ( .A1(n18646), .A2(P3_MORE_REG_SCAN_IN), .ZN(n18644) );
  OAI21_X1 U21743 ( .B1(n18646), .B2(n18645), .A(n18644), .ZN(P3_U3295) );
  OAI22_X1 U21744 ( .A1(n18650), .A2(n18649), .B1(n18648), .B2(n18647), .ZN(
        n18651) );
  NOR2_X1 U21745 ( .A1(n18669), .A2(n18651), .ZN(n18662) );
  AOI21_X1 U21746 ( .B1(n18654), .B2(n18653), .A(n18652), .ZN(n18656) );
  OAI211_X1 U21747 ( .C1(n18657), .C2(n18656), .A(P3_STATE2_REG_2__SCAN_IN), 
        .B(n18655), .ZN(n18659) );
  AOI21_X1 U21748 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n18659), .A(n18658), 
        .ZN(n18661) );
  NAND2_X1 U21749 ( .A1(n18662), .A2(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n18660) );
  OAI21_X1 U21750 ( .B1(n18662), .B2(n18661), .A(n18660), .ZN(P3_U3296) );
  INV_X1 U21751 ( .A(P3_MEMORYFETCH_REG_SCAN_IN), .ZN(n18672) );
  INV_X1 U21752 ( .A(P3_M_IO_N_REG_SCAN_IN), .ZN(n18664) );
  AOI22_X1 U21753 ( .A1(n18665), .A2(n18672), .B1(n18664), .B2(n18663), .ZN(
        P3_U3297) );
  AOI21_X1 U21754 ( .B1(n18667), .B2(n18666), .A(n18669), .ZN(n18673) );
  INV_X1 U21755 ( .A(P3_READREQUEST_REG_SCAN_IN), .ZN(n18670) );
  AOI22_X1 U21756 ( .A1(n18673), .A2(n18670), .B1(n18669), .B2(n18668), .ZN(
        P3_U3298) );
  AOI21_X1 U21757 ( .B1(n18673), .B2(n18672), .A(n18671), .ZN(P3_U3299) );
  INV_X1 U21758 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n19617) );
  INV_X1 U21759 ( .A(P2_ADS_N_REG_SCAN_IN), .ZN(n18674) );
  INV_X1 U21760 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n19633) );
  NAND2_X1 U21761 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n19633), .ZN(n19623) );
  AOI22_X1 U21762 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(n19623), .B1(
        P2_STATE_REG_1__SCAN_IN), .B2(n19617), .ZN(n19683) );
  INV_X1 U21763 ( .A(n19683), .ZN(n19616) );
  OAI21_X1 U21764 ( .B1(n19617), .B2(n18674), .A(n19616), .ZN(P2_U2815) );
  INV_X1 U21765 ( .A(P2_CODEFETCH_REG_SCAN_IN), .ZN(n18676) );
  OAI22_X1 U21766 ( .A1(n19735), .A2(n18676), .B1(n18954), .B2(n18675), .ZN(
        P2_U2816) );
  NAND2_X1 U21767 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n19617), .ZN(n19753) );
  AOI22_X1 U21768 ( .A1(P2_D_C_N_REG_SCAN_IN), .A2(n19753), .B1(n19625), .B2(
        n19617), .ZN(n18677) );
  OAI21_X1 U21769 ( .B1(P2_CODEFETCH_REG_SCAN_IN), .B2(n19753), .A(n18677), 
        .ZN(P2_U2817) );
  OAI21_X1 U21770 ( .B1(n19625), .B2(BS16), .A(n19683), .ZN(n19681) );
  OAI21_X1 U21771 ( .B1(n19683), .B2(n12954), .A(n19681), .ZN(P2_U2818) );
  NOR4_X1 U21772 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_21__SCAN_IN), .A3(P2_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_23__SCAN_IN), .ZN(n18681) );
  NOR4_X1 U21773 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_17__SCAN_IN), .A3(P2_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_19__SCAN_IN), .ZN(n18680) );
  NOR4_X1 U21774 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_29__SCAN_IN), .A3(P2_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_31__SCAN_IN), .ZN(n18679) );
  NOR4_X1 U21775 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_25__SCAN_IN), .A3(P2_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_27__SCAN_IN), .ZN(n18678) );
  NAND4_X1 U21776 ( .A1(n18681), .A2(n18680), .A3(n18679), .A4(n18678), .ZN(
        n18687) );
  NOR4_X1 U21777 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_4__SCAN_IN), .A3(P2_DATAWIDTH_REG_5__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_7__SCAN_IN), .ZN(n18685) );
  AOI211_X1 U21778 ( .C1(P2_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_0__SCAN_IN), .A(P2_DATAWIDTH_REG_6__SCAN_IN), .B(
        P2_DATAWIDTH_REG_2__SCAN_IN), .ZN(n18684) );
  NOR4_X1 U21779 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_13__SCAN_IN), .A3(P2_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_15__SCAN_IN), .ZN(n18683) );
  NOR4_X1 U21780 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_9__SCAN_IN), .A3(P2_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_11__SCAN_IN), .ZN(n18682) );
  NAND4_X1 U21781 ( .A1(n18685), .A2(n18684), .A3(n18683), .A4(n18682), .ZN(
        n18686) );
  NOR2_X1 U21782 ( .A1(n18687), .A2(n18686), .ZN(n18694) );
  INV_X1 U21783 ( .A(n18694), .ZN(n18693) );
  NOR2_X1 U21784 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n18693), .ZN(n18688) );
  INV_X1 U21785 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n19679) );
  AOI22_X1 U21786 ( .A1(n18688), .A2(n10947), .B1(n18693), .B2(n19679), .ZN(
        P2_U2820) );
  OR3_X1 U21787 ( .A1(P2_REIP_REG_0__SCAN_IN), .A2(P2_DATAWIDTH_REG_1__SCAN_IN), .A3(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n18692) );
  INV_X1 U21788 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n19677) );
  AOI22_X1 U21789 ( .A1(n18688), .A2(n18692), .B1(n18693), .B2(n19677), .ZN(
        P2_U2821) );
  INV_X1 U21790 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n19682) );
  NAND2_X1 U21791 ( .A1(n18688), .A2(n19682), .ZN(n18691) );
  OAI21_X1 U21792 ( .B1(n10947), .B2(n13175), .A(n18694), .ZN(n18689) );
  OAI21_X1 U21793 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n18694), .A(n18689), 
        .ZN(n18690) );
  OAI221_X1 U21794 ( .B1(n18691), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n18691), .C2(P2_REIP_REG_0__SCAN_IN), .A(n18690), .ZN(P2_U2822) );
  INV_X1 U21795 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n19675) );
  OAI221_X1 U21796 ( .B1(n18694), .B2(n19675), .C1(n18693), .C2(n18692), .A(
        n18691), .ZN(P2_U2823) );
  OAI22_X1 U21797 ( .A1(n18695), .A2(n18911), .B1(n19654), .B2(n18848), .ZN(
        n18699) );
  INV_X1 U21798 ( .A(n18696), .ZN(n18697) );
  OAI22_X1 U21799 ( .A1(n18697), .A2(n18923), .B1(n11346), .B2(n18810), .ZN(
        n18698) );
  AOI211_X1 U21800 ( .C1(n18700), .C2(n18917), .A(n18699), .B(n18698), .ZN(
        n18705) );
  OAI211_X1 U21801 ( .C1(n18703), .C2(n18702), .A(n10036), .B(n18701), .ZN(
        n18704) );
  OAI211_X1 U21802 ( .C1(n18894), .C2(n18706), .A(n18705), .B(n18704), .ZN(
        P2_U2834) );
  AOI22_X1 U21803 ( .A1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n18882), .B1(
        P2_REIP_REG_20__SCAN_IN), .B2(n18918), .ZN(n18717) );
  AOI22_X1 U21804 ( .A1(n18707), .A2(n18895), .B1(P2_EBX_REG_20__SCAN_IN), 
        .B2(n18919), .ZN(n18716) );
  INV_X1 U21805 ( .A(n18708), .ZN(n18709) );
  AOI22_X1 U21806 ( .A1(n18710), .A2(n18925), .B1(n18709), .B2(n18917), .ZN(
        n18715) );
  OAI211_X1 U21807 ( .C1(n18713), .C2(n18712), .A(n10036), .B(n18711), .ZN(
        n18714) );
  NAND4_X1 U21808 ( .A1(n18717), .A2(n18716), .A3(n18715), .A4(n18714), .ZN(
        P2_U2835) );
  AOI22_X1 U21809 ( .A1(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n18882), .B1(
        P2_EBX_REG_19__SCAN_IN), .B2(n18919), .ZN(n18718) );
  OAI21_X1 U21810 ( .B1(n18719), .B2(n18923), .A(n18718), .ZN(n18720) );
  AOI211_X1 U21811 ( .C1(P2_REIP_REG_19__SCAN_IN), .C2(n18918), .A(n19033), 
        .B(n18720), .ZN(n18728) );
  AOI22_X1 U21812 ( .A1(n18722), .A2(n18925), .B1(n18721), .B2(n18917), .ZN(
        n18727) );
  OAI211_X1 U21813 ( .C1(n18725), .C2(n18724), .A(n10036), .B(n18723), .ZN(
        n18726) );
  NAND3_X1 U21814 ( .A1(n18728), .A2(n18727), .A3(n18726), .ZN(P2_U2836) );
  AOI22_X1 U21815 ( .A1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n18882), .B1(
        P2_EBX_REG_18__SCAN_IN), .B2(n18919), .ZN(n18729) );
  OAI211_X1 U21816 ( .C1(n18848), .C2(n19650), .A(n18729), .B(n18846), .ZN(
        n18730) );
  INV_X1 U21817 ( .A(n18730), .ZN(n18731) );
  OAI21_X1 U21818 ( .B1(n18732), .B2(n18923), .A(n18731), .ZN(n18733) );
  AOI21_X1 U21819 ( .B1(n18734), .B2(n18925), .A(n18733), .ZN(n18739) );
  OAI211_X1 U21820 ( .C1(n18737), .C2(n18736), .A(n10036), .B(n18735), .ZN(
        n18738) );
  OAI211_X1 U21821 ( .C1(n18898), .C2(n18740), .A(n18739), .B(n18738), .ZN(
        P2_U2837) );
  NAND2_X1 U21822 ( .A1(n18863), .A2(n18741), .ZN(n18742) );
  XOR2_X1 U21823 ( .A(n18743), .B(n18742), .Z(n18752) );
  INV_X1 U21824 ( .A(n18744), .ZN(n18746) );
  AOI22_X1 U21825 ( .A1(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n18882), .B1(
        P2_EBX_REG_17__SCAN_IN), .B2(n18919), .ZN(n18745) );
  OAI21_X1 U21826 ( .B1(n18746), .B2(n18923), .A(n18745), .ZN(n18747) );
  AOI211_X1 U21827 ( .C1(P2_REIP_REG_17__SCAN_IN), .C2(n18918), .A(n19033), 
        .B(n18747), .ZN(n18751) );
  AOI22_X1 U21828 ( .A1(n18749), .A2(n18917), .B1(n18748), .B2(n18925), .ZN(
        n18750) );
  OAI211_X1 U21829 ( .C1(n19614), .C2(n18752), .A(n18751), .B(n18750), .ZN(
        P2_U2838) );
  OAI21_X1 U21830 ( .B1(n19647), .B2(n18848), .A(n18846), .ZN(n18756) );
  INV_X1 U21831 ( .A(n18753), .ZN(n18754) );
  OAI22_X1 U21832 ( .A1(n18754), .A2(n18923), .B1(n18810), .B2(n11351), .ZN(
        n18755) );
  AOI211_X1 U21833 ( .C1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .C2(n18882), .A(
        n18756), .B(n18755), .ZN(n18763) );
  NOR2_X1 U21834 ( .A1(n18903), .A2(n18757), .ZN(n18759) );
  XNOR2_X1 U21835 ( .A(n18759), .B(n18758), .ZN(n18760) );
  AOI22_X1 U21836 ( .A1(n18761), .A2(n18925), .B1(n10036), .B2(n18760), .ZN(
        n18762) );
  OAI211_X1 U21837 ( .C1(n18764), .C2(n18898), .A(n18763), .B(n18762), .ZN(
        P2_U2839) );
  INV_X1 U21838 ( .A(n18765), .ZN(n18767) );
  AOI22_X1 U21839 ( .A1(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n18882), .B1(
        P2_EBX_REG_15__SCAN_IN), .B2(n18919), .ZN(n18766) );
  OAI21_X1 U21840 ( .B1(n18767), .B2(n18923), .A(n18766), .ZN(n18768) );
  AOI211_X1 U21841 ( .C1(P2_REIP_REG_15__SCAN_IN), .C2(n18918), .A(n19033), 
        .B(n18768), .ZN(n18775) );
  NAND2_X1 U21842 ( .A1(n18863), .A2(n18769), .ZN(n18770) );
  XNOR2_X1 U21843 ( .A(n18771), .B(n18770), .ZN(n18772) );
  AOI22_X1 U21844 ( .A1(n18773), .A2(n18917), .B1(n18794), .B2(n18772), .ZN(
        n18774) );
  OAI211_X1 U21845 ( .C1(n18776), .C2(n18894), .A(n18775), .B(n18774), .ZN(
        P2_U2840) );
  AOI22_X1 U21846 ( .A1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n18882), .B1(
        P2_EBX_REG_14__SCAN_IN), .B2(n18919), .ZN(n18777) );
  OAI21_X1 U21847 ( .B1(n18778), .B2(n18923), .A(n18777), .ZN(n18779) );
  AOI211_X1 U21848 ( .C1(P2_REIP_REG_14__SCAN_IN), .C2(n18918), .A(n19033), 
        .B(n18779), .ZN(n18786) );
  NOR2_X1 U21849 ( .A1(n18903), .A2(n18780), .ZN(n18782) );
  XNOR2_X1 U21850 ( .A(n18782), .B(n18781), .ZN(n18783) );
  AOI22_X1 U21851 ( .A1(n18784), .A2(n18925), .B1(n10036), .B2(n18783), .ZN(
        n18785) );
  OAI211_X1 U21852 ( .C1(n18936), .C2(n18898), .A(n18786), .B(n18785), .ZN(
        P2_U2841) );
  AOI22_X1 U21853 ( .A1(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n18882), .B1(
        P2_EBX_REG_13__SCAN_IN), .B2(n18919), .ZN(n18787) );
  OAI21_X1 U21854 ( .B1(n18788), .B2(n18923), .A(n18787), .ZN(n18789) );
  AOI211_X1 U21855 ( .C1(P2_REIP_REG_13__SCAN_IN), .C2(n18918), .A(n19033), 
        .B(n18789), .ZN(n18796) );
  NAND2_X1 U21856 ( .A1(n18863), .A2(n18790), .ZN(n18791) );
  XNOR2_X1 U21857 ( .A(n18792), .B(n18791), .ZN(n18793) );
  AOI22_X1 U21858 ( .A1(n18938), .A2(n18917), .B1(n18794), .B2(n18793), .ZN(
        n18795) );
  OAI211_X1 U21859 ( .C1(n18797), .C2(n18894), .A(n18796), .B(n18795), .ZN(
        P2_U2842) );
  AOI22_X1 U21860 ( .A1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n18882), .B1(
        P2_EBX_REG_12__SCAN_IN), .B2(n18919), .ZN(n18798) );
  OAI21_X1 U21861 ( .B1(n18799), .B2(n18923), .A(n18798), .ZN(n18800) );
  AOI211_X1 U21862 ( .C1(P2_REIP_REG_12__SCAN_IN), .C2(n18918), .A(n19033), 
        .B(n18800), .ZN(n18807) );
  NOR2_X1 U21863 ( .A1(n18903), .A2(n18801), .ZN(n18803) );
  XNOR2_X1 U21864 ( .A(n18803), .B(n18802), .ZN(n18804) );
  AOI22_X1 U21865 ( .A1(n18805), .A2(n18925), .B1(n10036), .B2(n18804), .ZN(
        n18806) );
  OAI211_X1 U21866 ( .C1(n18808), .C2(n18898), .A(n18807), .B(n18806), .ZN(
        P2_U2843) );
  OAI21_X1 U21867 ( .B1(n11591), .B2(n18848), .A(n18846), .ZN(n18813) );
  OAI22_X1 U21868 ( .A1(n18811), .A2(n18923), .B1(n18810), .B2(n18809), .ZN(
        n18812) );
  AOI211_X1 U21869 ( .C1(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .C2(n18882), .A(
        n18813), .B(n18812), .ZN(n18819) );
  NAND2_X1 U21870 ( .A1(n18863), .A2(n18814), .ZN(n18815) );
  XNOR2_X1 U21871 ( .A(n18816), .B(n18815), .ZN(n18817) );
  AOI22_X1 U21872 ( .A1(n18940), .A2(n18917), .B1(n10036), .B2(n18817), .ZN(
        n18818) );
  OAI211_X1 U21873 ( .C1(n18820), .C2(n18894), .A(n18819), .B(n18818), .ZN(
        P2_U2844) );
  INV_X1 U21874 ( .A(n18821), .ZN(n18822) );
  AOI22_X1 U21875 ( .A1(n18822), .A2(n18895), .B1(P2_EBX_REG_10__SCAN_IN), 
        .B2(n18919), .ZN(n18824) );
  OAI211_X1 U21876 ( .C1(n11585), .C2(n18848), .A(n18824), .B(n18823), .ZN(
        n18825) );
  AOI21_X1 U21877 ( .B1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n18882), .A(
        n18825), .ZN(n18832) );
  NOR2_X1 U21878 ( .A1(n18903), .A2(n18826), .ZN(n18828) );
  XNOR2_X1 U21879 ( .A(n18828), .B(n18827), .ZN(n18829) );
  AOI22_X1 U21880 ( .A1(n18830), .A2(n18925), .B1(n10036), .B2(n18829), .ZN(
        n18831) );
  OAI211_X1 U21881 ( .C1(n18833), .C2(n18898), .A(n18832), .B(n18831), .ZN(
        P2_U2845) );
  AOI22_X1 U21882 ( .A1(n18834), .A2(n18895), .B1(P2_EBX_REG_9__SCAN_IN), .B2(
        n18919), .ZN(n18835) );
  OAI21_X1 U21883 ( .B1(n18836), .B2(n18911), .A(n18835), .ZN(n18837) );
  AOI211_X1 U21884 ( .C1(P2_REIP_REG_9__SCAN_IN), .C2(n18918), .A(n19033), .B(
        n18837), .ZN(n18843) );
  NAND2_X1 U21885 ( .A1(n18863), .A2(n18838), .ZN(n18839) );
  XNOR2_X1 U21886 ( .A(n18840), .B(n18839), .ZN(n18841) );
  AOI22_X1 U21887 ( .A1(n18917), .A2(n18943), .B1(n10036), .B2(n18841), .ZN(
        n18842) );
  OAI211_X1 U21888 ( .C1(n18894), .C2(n18844), .A(n18843), .B(n18842), .ZN(
        P2_U2846) );
  AOI22_X1 U21889 ( .A1(n18845), .A2(n18895), .B1(P2_EBX_REG_8__SCAN_IN), .B2(
        n18919), .ZN(n18847) );
  OAI211_X1 U21890 ( .C1(n11576), .C2(n18848), .A(n18847), .B(n18846), .ZN(
        n18849) );
  AOI21_X1 U21891 ( .B1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n18882), .A(
        n18849), .ZN(n18856) );
  NOR2_X1 U21892 ( .A1(n18903), .A2(n18850), .ZN(n18852) );
  XNOR2_X1 U21893 ( .A(n18852), .B(n18851), .ZN(n18854) );
  AOI22_X1 U21894 ( .A1(n10036), .A2(n18854), .B1(n18925), .B2(n18853), .ZN(
        n18855) );
  OAI211_X1 U21895 ( .C1(n18898), .C2(n18857), .A(n18856), .B(n18855), .ZN(
        P2_U2847) );
  AOI22_X1 U21896 ( .A1(n18858), .A2(n18895), .B1(P2_EBX_REG_7__SCAN_IN), .B2(
        n18919), .ZN(n18859) );
  OAI21_X1 U21897 ( .B1(n18860), .B2(n18911), .A(n18859), .ZN(n18861) );
  AOI211_X1 U21898 ( .C1(P2_REIP_REG_7__SCAN_IN), .C2(n18918), .A(n19033), .B(
        n18861), .ZN(n18869) );
  NAND2_X1 U21899 ( .A1(n18863), .A2(n18862), .ZN(n18864) );
  XNOR2_X1 U21900 ( .A(n18865), .B(n18864), .ZN(n18866) );
  AOI22_X1 U21901 ( .A1(n18917), .A2(n18867), .B1(n10036), .B2(n18866), .ZN(
        n18868) );
  OAI211_X1 U21902 ( .C1(n18894), .C2(n18870), .A(n18869), .B(n18868), .ZN(
        P2_U2848) );
  AOI22_X1 U21903 ( .A1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n18882), .B1(
        P2_EBX_REG_6__SCAN_IN), .B2(n18919), .ZN(n18871) );
  OAI21_X1 U21904 ( .B1(n18872), .B2(n18923), .A(n18871), .ZN(n18873) );
  AOI211_X1 U21905 ( .C1(P2_REIP_REG_6__SCAN_IN), .C2(n18918), .A(n19033), .B(
        n18873), .ZN(n18880) );
  NOR2_X1 U21906 ( .A1(n18903), .A2(n18874), .ZN(n18876) );
  XNOR2_X1 U21907 ( .A(n18876), .B(n18875), .ZN(n18878) );
  AOI22_X1 U21908 ( .A1(n10036), .A2(n18878), .B1(n18925), .B2(n18877), .ZN(
        n18879) );
  OAI211_X1 U21909 ( .C1(n18898), .C2(n18881), .A(n18880), .B(n18879), .ZN(
        P2_U2849) );
  AOI22_X1 U21910 ( .A1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n18882), .B1(
        P2_EBX_REG_5__SCAN_IN), .B2(n18919), .ZN(n18883) );
  OAI21_X1 U21911 ( .B1(n18884), .B2(n18923), .A(n18883), .ZN(n18885) );
  AOI211_X1 U21912 ( .C1(P2_REIP_REG_5__SCAN_IN), .C2(n18918), .A(n19033), .B(
        n18885), .ZN(n18892) );
  NAND2_X1 U21913 ( .A1(n18863), .A2(n18886), .ZN(n18887) );
  XNOR2_X1 U21914 ( .A(n18888), .B(n18887), .ZN(n18889) );
  AOI22_X1 U21915 ( .A1(n18917), .A2(n18890), .B1(n10036), .B2(n18889), .ZN(
        n18891) );
  OAI211_X1 U21916 ( .C1(n18894), .C2(n18893), .A(n18892), .B(n18891), .ZN(
        P2_U2850) );
  AOI22_X1 U21917 ( .A1(n18896), .A2(n18895), .B1(P2_EBX_REG_4__SCAN_IN), .B2(
        n18919), .ZN(n18910) );
  INV_X1 U21918 ( .A(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n18899) );
  OAI22_X1 U21919 ( .A1(n18899), .A2(n18911), .B1(n18898), .B2(n18897), .ZN(
        n18900) );
  AOI211_X1 U21920 ( .C1(P2_REIP_REG_4__SCAN_IN), .C2(n18918), .A(n19033), .B(
        n18900), .ZN(n18909) );
  AOI22_X1 U21921 ( .A1(n18901), .A2(n18913), .B1(n18925), .B2(n19040), .ZN(
        n18908) );
  INV_X1 U21922 ( .A(n19044), .ZN(n18906) );
  NOR2_X1 U21923 ( .A1(n18903), .A2(n18902), .ZN(n18905) );
  AOI21_X1 U21924 ( .B1(n18906), .B2(n18905), .A(n19614), .ZN(n18904) );
  OAI21_X1 U21925 ( .B1(n18906), .B2(n18905), .A(n18904), .ZN(n18907) );
  NAND4_X1 U21926 ( .A1(n18910), .A2(n18909), .A3(n18908), .A4(n18907), .ZN(
        P2_U2851) );
  NAND2_X1 U21927 ( .A1(n18911), .A2(n19614), .ZN(n18914) );
  AOI22_X1 U21928 ( .A1(n18914), .A2(P2_PHYADDRPOINTER_REG_0__SCAN_IN), .B1(
        n18913), .B2(n18912), .ZN(n18928) );
  INV_X1 U21929 ( .A(n18915), .ZN(n18922) );
  AOI22_X1 U21930 ( .A1(n18918), .A2(P2_REIP_REG_0__SCAN_IN), .B1(n18917), 
        .B2(n18916), .ZN(n18921) );
  NAND2_X1 U21931 ( .A1(n18919), .A2(P2_EBX_REG_0__SCAN_IN), .ZN(n18920) );
  OAI211_X1 U21932 ( .C1(n18923), .C2(n18922), .A(n18921), .B(n18920), .ZN(
        n18924) );
  AOI21_X1 U21933 ( .B1(n18926), .B2(n18925), .A(n18924), .ZN(n18927) );
  NAND2_X1 U21934 ( .A1(n18928), .A2(n18927), .ZN(P2_U2855) );
  AOI22_X1 U21935 ( .A1(n15826), .A2(n18930), .B1(n18929), .B2(
        BUF2_REG_31__SCAN_IN), .ZN(n18933) );
  AOI22_X1 U21936 ( .A1(BUF1_REG_31__SCAN_IN), .A2(n18931), .B1(
        P2_EAX_REG_31__SCAN_IN), .B2(n18934), .ZN(n18932) );
  NAND2_X1 U21937 ( .A1(n18933), .A2(n18932), .ZN(P2_U2888) );
  AOI22_X1 U21938 ( .A1(n18946), .A2(n19023), .B1(n18934), .B2(
        P2_EAX_REG_14__SCAN_IN), .ZN(n18935) );
  OAI21_X1 U21939 ( .B1(n18937), .B2(n18936), .A(n18935), .ZN(P2_U2905) );
  INV_X1 U21940 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n18993) );
  AOI22_X1 U21941 ( .A1(n18946), .A2(n19021), .B1(n18944), .B2(n18938), .ZN(
        n18939) );
  OAI21_X1 U21942 ( .B1(n18948), .B2(n18993), .A(n18939), .ZN(P2_U2906) );
  AOI22_X1 U21943 ( .A1(n18946), .A2(n18941), .B1(n18944), .B2(n18940), .ZN(
        n18942) );
  OAI21_X1 U21944 ( .B1(n18948), .B2(n20931), .A(n18942), .ZN(P2_U2908) );
  AOI22_X1 U21945 ( .A1(n18946), .A2(n18945), .B1(n18944), .B2(n18943), .ZN(
        n18947) );
  OAI21_X1 U21946 ( .B1(n18948), .B2(n19000), .A(n18947), .ZN(P2_U2910) );
  NAND2_X1 U21947 ( .A1(n18950), .A2(n18949), .ZN(n18952) );
  NAND2_X1 U21948 ( .A1(n18952), .A2(n18951), .ZN(n18953) );
  NAND2_X1 U21949 ( .A1(n19719), .A2(n18954), .ZN(n18956) );
  NOR2_X1 U21950 ( .A1(n18962), .A2(n18955), .ZN(P2_U2920) );
  OR2_X1 U21951 ( .A1(n19019), .A2(n19739), .ZN(n18987) );
  INV_X1 U21952 ( .A(n18987), .ZN(n18959) );
  AOI22_X1 U21953 ( .A1(P2_EAX_REG_30__SCAN_IN), .A2(n18959), .B1(n19017), 
        .B2(P2_UWORD_REG_14__SCAN_IN), .ZN(n18957) );
  OAI21_X1 U21954 ( .B1(n18958), .B2(n18962), .A(n18957), .ZN(P2_U2921) );
  AOI22_X1 U21955 ( .A1(P2_EAX_REG_29__SCAN_IN), .A2(n18959), .B1(n19017), 
        .B2(P2_UWORD_REG_13__SCAN_IN), .ZN(n18960) );
  OAI21_X1 U21956 ( .B1(n18962), .B2(n18961), .A(n18960), .ZN(P2_U2922) );
  AOI22_X1 U21957 ( .A1(n19017), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(n19006), 
        .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n18963) );
  OAI21_X1 U21958 ( .B1(n18964), .B2(n18987), .A(n18963), .ZN(P2_U2923) );
  AOI22_X1 U21959 ( .A1(n19017), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(n19006), 
        .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n18965) );
  OAI21_X1 U21960 ( .B1(n18966), .B2(n18987), .A(n18965), .ZN(P2_U2924) );
  AOI22_X1 U21961 ( .A1(n19017), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(n19006), 
        .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n18967) );
  OAI21_X1 U21962 ( .B1(n18968), .B2(n18987), .A(n18967), .ZN(P2_U2925) );
  AOI22_X1 U21963 ( .A1(n19017), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(n19006), 
        .B2(P2_DATAO_REG_25__SCAN_IN), .ZN(n18969) );
  OAI21_X1 U21964 ( .B1(n18970), .B2(n18987), .A(n18969), .ZN(P2_U2926) );
  AOI22_X1 U21965 ( .A1(n19017), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n19006), 
        .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n18971) );
  OAI21_X1 U21966 ( .B1(n18972), .B2(n18987), .A(n18971), .ZN(P2_U2927) );
  INV_X1 U21967 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n20851) );
  AOI22_X1 U21968 ( .A1(n19017), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n19006), 
        .B2(P2_DATAO_REG_23__SCAN_IN), .ZN(n18973) );
  OAI21_X1 U21969 ( .B1(n20851), .B2(n18987), .A(n18973), .ZN(P2_U2928) );
  AOI22_X1 U21970 ( .A1(n19017), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(n19006), 
        .B2(P2_DATAO_REG_22__SCAN_IN), .ZN(n18974) );
  OAI21_X1 U21971 ( .B1(n18975), .B2(n18987), .A(n18974), .ZN(P2_U2929) );
  AOI22_X1 U21972 ( .A1(n19017), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n19006), 
        .B2(P2_DATAO_REG_21__SCAN_IN), .ZN(n18976) );
  OAI21_X1 U21973 ( .B1(n18977), .B2(n18987), .A(n18976), .ZN(P2_U2930) );
  AOI22_X1 U21974 ( .A1(n19017), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n19006), 
        .B2(P2_DATAO_REG_20__SCAN_IN), .ZN(n18978) );
  OAI21_X1 U21975 ( .B1(n18979), .B2(n18987), .A(n18978), .ZN(P2_U2931) );
  AOI22_X1 U21976 ( .A1(n19017), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n19006), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n18980) );
  OAI21_X1 U21977 ( .B1(n18981), .B2(n18987), .A(n18980), .ZN(P2_U2932) );
  AOI22_X1 U21978 ( .A1(n19017), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n19006), 
        .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n18982) );
  OAI21_X1 U21979 ( .B1(n18983), .B2(n18987), .A(n18982), .ZN(P2_U2933) );
  AOI22_X1 U21980 ( .A1(n19017), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n19006), 
        .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n18984) );
  OAI21_X1 U21981 ( .B1(n18985), .B2(n18987), .A(n18984), .ZN(P2_U2934) );
  AOI22_X1 U21982 ( .A1(n19017), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(n19006), 
        .B2(P2_DATAO_REG_16__SCAN_IN), .ZN(n18986) );
  OAI21_X1 U21983 ( .B1(n18988), .B2(n18987), .A(n18986), .ZN(P2_U2935) );
  AOI22_X1 U21984 ( .A1(n19017), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n19006), 
        .B2(P2_DATAO_REG_15__SCAN_IN), .ZN(n18989) );
  OAI21_X1 U21985 ( .B1(n12890), .B2(n19019), .A(n18989), .ZN(P2_U2936) );
  INV_X1 U21986 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n18991) );
  AOI22_X1 U21987 ( .A1(n19017), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n19006), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n18990) );
  OAI21_X1 U21988 ( .B1(n18991), .B2(n19019), .A(n18990), .ZN(P2_U2937) );
  AOI22_X1 U21989 ( .A1(n19017), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n19006), 
        .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n18992) );
  OAI21_X1 U21990 ( .B1(n18993), .B2(n19019), .A(n18992), .ZN(P2_U2938) );
  AOI22_X1 U21991 ( .A1(n19017), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(n19006), 
        .B2(P2_DATAO_REG_12__SCAN_IN), .ZN(n18994) );
  OAI21_X1 U21992 ( .B1(n18995), .B2(n19019), .A(n18994), .ZN(P2_U2939) );
  AOI22_X1 U21993 ( .A1(n19017), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n19006), 
        .B2(P2_DATAO_REG_11__SCAN_IN), .ZN(n18996) );
  OAI21_X1 U21994 ( .B1(n20931), .B2(n19019), .A(n18996), .ZN(P2_U2940) );
  AOI22_X1 U21995 ( .A1(n19017), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n19006), 
        .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n18997) );
  OAI21_X1 U21996 ( .B1(n18998), .B2(n19019), .A(n18997), .ZN(P2_U2941) );
  AOI22_X1 U21997 ( .A1(n19017), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n19006), 
        .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n18999) );
  OAI21_X1 U21998 ( .B1(n19000), .B2(n19019), .A(n18999), .ZN(P2_U2942) );
  AOI22_X1 U21999 ( .A1(n19017), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n19006), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n19001) );
  OAI21_X1 U22000 ( .B1(n19002), .B2(n19019), .A(n19001), .ZN(P2_U2943) );
  AOI22_X1 U22001 ( .A1(n19017), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n19006), 
        .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n19003) );
  OAI21_X1 U22002 ( .B1(n11992), .B2(n19019), .A(n19003), .ZN(P2_U2944) );
  AOI22_X1 U22003 ( .A1(n19017), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n19006), 
        .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n19004) );
  OAI21_X1 U22004 ( .B1(n19005), .B2(n19019), .A(n19004), .ZN(P2_U2945) );
  INV_X1 U22005 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n19008) );
  AOI22_X1 U22006 ( .A1(n19017), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n19006), 
        .B2(P2_DATAO_REG_5__SCAN_IN), .ZN(n19007) );
  OAI21_X1 U22007 ( .B1(n19008), .B2(n19019), .A(n19007), .ZN(P2_U2946) );
  INV_X1 U22008 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n19010) );
  AOI22_X1 U22009 ( .A1(n19017), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n19006), 
        .B2(P2_DATAO_REG_4__SCAN_IN), .ZN(n19009) );
  OAI21_X1 U22010 ( .B1(n19010), .B2(n19019), .A(n19009), .ZN(P2_U2947) );
  INV_X1 U22011 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n19012) );
  AOI22_X1 U22012 ( .A1(n19017), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n19006), 
        .B2(P2_DATAO_REG_3__SCAN_IN), .ZN(n19011) );
  OAI21_X1 U22013 ( .B1(n19012), .B2(n19019), .A(n19011), .ZN(P2_U2948) );
  INV_X1 U22014 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n19014) );
  AOI22_X1 U22015 ( .A1(n19017), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n19006), 
        .B2(P2_DATAO_REG_2__SCAN_IN), .ZN(n19013) );
  OAI21_X1 U22016 ( .B1(n19014), .B2(n19019), .A(n19013), .ZN(P2_U2949) );
  INV_X1 U22017 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n19016) );
  AOI22_X1 U22018 ( .A1(n19017), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n19006), 
        .B2(P2_DATAO_REG_1__SCAN_IN), .ZN(n19015) );
  OAI21_X1 U22019 ( .B1(n19016), .B2(n19019), .A(n19015), .ZN(P2_U2950) );
  INV_X1 U22020 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n19020) );
  AOI22_X1 U22021 ( .A1(n19017), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n19006), 
        .B2(P2_DATAO_REG_0__SCAN_IN), .ZN(n19018) );
  OAI21_X1 U22022 ( .B1(n19020), .B2(n19019), .A(n19018), .ZN(P2_U2951) );
  AOI22_X1 U22023 ( .A1(n19029), .A2(P2_EAX_REG_29__SCAN_IN), .B1(n19028), 
        .B2(P2_UWORD_REG_13__SCAN_IN), .ZN(n19022) );
  NAND2_X1 U22024 ( .A1(n19024), .A2(n19021), .ZN(n19026) );
  NAND2_X1 U22025 ( .A1(n19022), .A2(n19026), .ZN(P2_U2965) );
  AOI22_X1 U22026 ( .A1(n19029), .A2(P2_EAX_REG_30__SCAN_IN), .B1(n19028), 
        .B2(P2_UWORD_REG_14__SCAN_IN), .ZN(n19025) );
  NAND2_X1 U22027 ( .A1(n19024), .A2(n19023), .ZN(n19030) );
  NAND2_X1 U22028 ( .A1(n19025), .A2(n19030), .ZN(P2_U2966) );
  AOI22_X1 U22029 ( .A1(n19029), .A2(P2_EAX_REG_13__SCAN_IN), .B1(n19028), 
        .B2(P2_LWORD_REG_13__SCAN_IN), .ZN(n19027) );
  NAND2_X1 U22030 ( .A1(n19027), .A2(n19026), .ZN(P2_U2980) );
  AOI22_X1 U22031 ( .A1(n19029), .A2(P2_EAX_REG_14__SCAN_IN), .B1(n19028), 
        .B2(P2_LWORD_REG_14__SCAN_IN), .ZN(n19031) );
  NAND2_X1 U22032 ( .A1(n19031), .A2(n19030), .ZN(P2_U2981) );
  AOI22_X1 U22033 ( .A1(P2_REIP_REG_4__SCAN_IN), .A2(n19033), .B1(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n19032), .ZN(n19043) );
  INV_X1 U22034 ( .A(n19034), .ZN(n19036) );
  OAI22_X1 U22035 ( .A1(n19038), .A2(n19037), .B1(n19036), .B2(n19035), .ZN(
        n19039) );
  AOI21_X1 U22036 ( .B1(n19041), .B2(n19040), .A(n19039), .ZN(n19042) );
  OAI211_X1 U22037 ( .C1(n19045), .C2(n19044), .A(n19043), .B(n19042), .ZN(
        P2_U3010) );
  NOR2_X1 U22038 ( .A1(n19047), .A2(n19046), .ZN(n19051) );
  NOR2_X1 U22039 ( .A1(n19048), .A2(n19052), .ZN(n19050) );
  NOR3_X1 U22040 ( .A1(n19051), .A2(n19050), .A3(n19049), .ZN(n19068) );
  NAND3_X1 U22041 ( .A1(n19053), .A2(n19052), .A3(n19067), .ZN(n19054) );
  OAI21_X1 U22042 ( .B1(n19056), .B2(n19055), .A(n19054), .ZN(n19057) );
  AOI211_X1 U22043 ( .C1(n19059), .C2(n19702), .A(n19058), .B(n19057), .ZN(
        n19060) );
  OAI21_X1 U22044 ( .B1(n11148), .B2(n19061), .A(n19060), .ZN(n19062) );
  AOI211_X1 U22045 ( .C1(n19065), .C2(n19064), .A(n19063), .B(n19062), .ZN(
        n19066) );
  OAI21_X1 U22046 ( .B1(n19068), .B2(n19067), .A(n19066), .ZN(P2_U3044) );
  AOI22_X1 U22047 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n19090), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n19089), .ZN(n19480) );
  INV_X1 U22048 ( .A(n19480), .ZN(n19567) );
  AOI22_X1 U22049 ( .A1(n19567), .A2(n19087), .B1(n19086), .B2(n19565), .ZN(
        n19072) );
  NOR2_X2 U22050 ( .A1(n19069), .A2(n19426), .ZN(n19566) );
  OAI22_X2 U22051 ( .A1(n14174), .A2(n19080), .B1(n19070), .B2(n19079), .ZN(
        n19518) );
  AOI22_X1 U22052 ( .A1(n19566), .A2(n19091), .B1(n19131), .B2(n19518), .ZN(
        n19071) );
  OAI211_X1 U22053 ( .C1(n19095), .C2(n10477), .A(n19072), .B(n19071), .ZN(
        P2_U3050) );
  AOI22_X1 U22054 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n19090), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n19089), .ZN(n19486) );
  INV_X1 U22055 ( .A(n19486), .ZN(n19573) );
  AOI22_X1 U22056 ( .A1(n19573), .A2(n19087), .B1(n19086), .B2(n19571), .ZN(
        n19075) );
  NOR2_X2 U22057 ( .A1(n19073), .A2(n19426), .ZN(n19572) );
  AOI22_X1 U22058 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n19090), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n19089), .ZN(n19576) );
  AOI22_X1 U22059 ( .A1(n19572), .A2(n19091), .B1(n19131), .B2(n19522), .ZN(
        n19074) );
  OAI211_X1 U22060 ( .C1(n19095), .C2(n11169), .A(n19075), .B(n19074), .ZN(
        P2_U3051) );
  AOI22_X1 U22061 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n19089), .B1(
        BUF1_REG_28__SCAN_IN), .B2(n19090), .ZN(n19492) );
  INV_X1 U22062 ( .A(n19492), .ZN(n19579) );
  AND2_X1 U22063 ( .A1(n19077), .A2(n19076), .ZN(n19577) );
  AOI22_X1 U22064 ( .A1(n19579), .A2(n19087), .B1(n19086), .B2(n19577), .ZN(
        n19083) );
  NOR2_X2 U22065 ( .A1(n19078), .A2(n19426), .ZN(n19578) );
  OAI22_X2 U22066 ( .A1(n19081), .A2(n19080), .B1(n20770), .B2(n19079), .ZN(
        n19525) );
  AOI22_X1 U22067 ( .A1(n19578), .A2(n19091), .B1(n19131), .B2(n19525), .ZN(
        n19082) );
  OAI211_X1 U22068 ( .C1(n19095), .C2(n10773), .A(n19083), .B(n19082), .ZN(
        P2_U3052) );
  AOI22_X1 U22069 ( .A1(BUF2_REG_30__SCAN_IN), .A2(n19089), .B1(
        BUF1_REG_30__SCAN_IN), .B2(n19090), .ZN(n19504) );
  NOR2_X2 U22070 ( .A1(n19085), .A2(n19084), .ZN(n19589) );
  AOI22_X1 U22071 ( .A1(n19591), .A2(n19087), .B1(n19086), .B2(n19589), .ZN(
        n19093) );
  NOR2_X2 U22072 ( .A1(n19088), .A2(n19426), .ZN(n19590) );
  AOI22_X1 U22073 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n19090), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n19089), .ZN(n19594) );
  INV_X1 U22074 ( .A(n19594), .ZN(n19532) );
  AOI22_X1 U22075 ( .A1(n19590), .A2(n19091), .B1(n19131), .B2(n19532), .ZN(
        n19092) );
  OAI211_X1 U22076 ( .C1(n19095), .C2(n19094), .A(n19093), .B(n19092), .ZN(
        P2_U3054) );
  INV_X1 U22077 ( .A(n19096), .ZN(n19165) );
  NOR2_X1 U22078 ( .A1(n19336), .A2(n19165), .ZN(n19107) );
  INV_X1 U22079 ( .A(n19107), .ZN(n19128) );
  AND2_X1 U22080 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19128), .ZN(n19097) );
  AND2_X1 U22081 ( .A1(n19098), .A2(n19097), .ZN(n19103) );
  NAND2_X1 U22082 ( .A1(n19744), .A2(n19104), .ZN(n19099) );
  NAND2_X1 U22083 ( .A1(n19100), .A2(n19099), .ZN(n19101) );
  INV_X1 U22084 ( .A(n19547), .ZN(n19456) );
  OAI22_X1 U22085 ( .A1(n19129), .A2(n19457), .B1(n19456), .B2(n19128), .ZN(
        n19102) );
  INV_X1 U22086 ( .A(n19102), .ZN(n19109) );
  NAND2_X1 U22087 ( .A1(n19226), .A2(n19338), .ZN(n19105) );
  AOI21_X1 U22088 ( .B1(n19105), .B2(n19104), .A(n19103), .ZN(n19106) );
  OAI211_X1 U22089 ( .C1(n19107), .C2(n19714), .A(n19106), .B(n19549), .ZN(
        n19132) );
  AOI22_X1 U22090 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19132), .B1(
        n19131), .B2(n19555), .ZN(n19108) );
  OAI211_X1 U22091 ( .C1(n19558), .C2(n19153), .A(n19109), .B(n19108), .ZN(
        P2_U3056) );
  INV_X1 U22092 ( .A(n19559), .ZN(n19469) );
  OAI22_X1 U22093 ( .A1(n19129), .A2(n19470), .B1(n19469), .B2(n19128), .ZN(
        n19110) );
  INV_X1 U22094 ( .A(n19110), .ZN(n19112) );
  AOI22_X1 U22095 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19132), .B1(
        n19131), .B2(n19561), .ZN(n19111) );
  OAI211_X1 U22096 ( .C1(n19564), .C2(n19153), .A(n19112), .B(n19111), .ZN(
        P2_U3057) );
  INV_X1 U22097 ( .A(n19518), .ZN(n19570) );
  INV_X1 U22098 ( .A(n19566), .ZN(n19476) );
  INV_X1 U22099 ( .A(n19565), .ZN(n19475) );
  OAI22_X1 U22100 ( .A1(n19129), .A2(n19476), .B1(n19475), .B2(n19128), .ZN(
        n19113) );
  INV_X1 U22101 ( .A(n19113), .ZN(n19115) );
  AOI22_X1 U22102 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19132), .B1(
        n19131), .B2(n19567), .ZN(n19114) );
  OAI211_X1 U22103 ( .C1(n19570), .C2(n19153), .A(n19115), .B(n19114), .ZN(
        P2_U3058) );
  INV_X1 U22104 ( .A(n19572), .ZN(n19482) );
  INV_X1 U22105 ( .A(n19571), .ZN(n19481) );
  OAI22_X1 U22106 ( .A1(n19129), .A2(n19482), .B1(n19481), .B2(n19128), .ZN(
        n19116) );
  INV_X1 U22107 ( .A(n19116), .ZN(n19118) );
  AOI22_X1 U22108 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19132), .B1(
        n19131), .B2(n19573), .ZN(n19117) );
  OAI211_X1 U22109 ( .C1(n19576), .C2(n19153), .A(n19118), .B(n19117), .ZN(
        P2_U3059) );
  INV_X1 U22110 ( .A(n19578), .ZN(n19488) );
  INV_X1 U22111 ( .A(n19577), .ZN(n19487) );
  OAI22_X1 U22112 ( .A1(n19129), .A2(n19488), .B1(n19487), .B2(n19128), .ZN(
        n19119) );
  INV_X1 U22113 ( .A(n19119), .ZN(n19121) );
  AOI22_X1 U22114 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19132), .B1(
        n19131), .B2(n19579), .ZN(n19120) );
  OAI211_X1 U22115 ( .C1(n19582), .C2(n19153), .A(n19121), .B(n19120), .ZN(
        P2_U3060) );
  INV_X1 U22116 ( .A(n19583), .ZN(n19493) );
  OAI22_X1 U22117 ( .A1(n19129), .A2(n19494), .B1(n19493), .B2(n19128), .ZN(
        n19122) );
  INV_X1 U22118 ( .A(n19122), .ZN(n19124) );
  AOI22_X1 U22119 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19132), .B1(
        n19131), .B2(n19585), .ZN(n19123) );
  OAI211_X1 U22120 ( .C1(n19588), .C2(n19153), .A(n19124), .B(n19123), .ZN(
        P2_U3061) );
  INV_X1 U22121 ( .A(n19590), .ZN(n19500) );
  INV_X1 U22122 ( .A(n19589), .ZN(n19499) );
  OAI22_X1 U22123 ( .A1(n19129), .A2(n19500), .B1(n19499), .B2(n19128), .ZN(
        n19125) );
  INV_X1 U22124 ( .A(n19125), .ZN(n19127) );
  AOI22_X1 U22125 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19132), .B1(
        n19131), .B2(n19591), .ZN(n19126) );
  OAI211_X1 U22126 ( .C1(n19594), .C2(n19153), .A(n19127), .B(n19126), .ZN(
        P2_U3062) );
  INV_X1 U22127 ( .A(n19596), .ZN(n19506) );
  OAI22_X1 U22128 ( .A1(n19129), .A2(n19507), .B1(n19506), .B2(n19128), .ZN(
        n19130) );
  INV_X1 U22129 ( .A(n19130), .ZN(n19134) );
  AOI22_X1 U22130 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19132), .B1(
        n19131), .B2(n19599), .ZN(n19133) );
  OAI211_X1 U22131 ( .C1(n19605), .C2(n19153), .A(n19134), .B(n19133), .ZN(
        P2_U3063) );
  NOR2_X1 U22132 ( .A1(n19368), .A2(n19165), .ZN(n19156) );
  OAI21_X1 U22133 ( .B1(n19135), .B2(n19156), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19136) );
  OR2_X1 U22134 ( .A1(n19371), .A2(n19165), .ZN(n19137) );
  NAND2_X1 U22135 ( .A1(n19136), .A2(n19137), .ZN(n19157) );
  AOI22_X1 U22136 ( .A1(n19157), .A2(n12991), .B1(n19547), .B2(n19156), .ZN(
        n19142) );
  AOI21_X1 U22137 ( .B1(n11218), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n19140) );
  INV_X1 U22138 ( .A(n19153), .ZN(n19158) );
  OAI21_X1 U22139 ( .B1(n19186), .B2(n19158), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19138) );
  NAND3_X1 U22140 ( .A1(n19138), .A2(n19685), .A3(n19137), .ZN(n19139) );
  OAI211_X1 U22141 ( .C1(n19156), .C2(n19140), .A(n19139), .B(n19549), .ZN(
        n19159) );
  AOI22_X1 U22142 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19159), .B1(
        n19186), .B2(n19465), .ZN(n19141) );
  OAI211_X1 U22143 ( .C1(n19468), .C2(n19153), .A(n19142), .B(n19141), .ZN(
        P2_U3064) );
  AOI22_X1 U22144 ( .A1(n19157), .A2(n19560), .B1(n19559), .B2(n19156), .ZN(
        n19144) );
  AOI22_X1 U22145 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19159), .B1(
        n19158), .B2(n19561), .ZN(n19143) );
  OAI211_X1 U22146 ( .C1(n19564), .C2(n19194), .A(n19144), .B(n19143), .ZN(
        P2_U3065) );
  AOI22_X1 U22147 ( .A1(n19157), .A2(n19566), .B1(n19565), .B2(n19156), .ZN(
        n19146) );
  AOI22_X1 U22148 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19159), .B1(
        n19186), .B2(n19518), .ZN(n19145) );
  OAI211_X1 U22149 ( .C1(n19480), .C2(n19153), .A(n19146), .B(n19145), .ZN(
        P2_U3066) );
  AOI22_X1 U22150 ( .A1(n19157), .A2(n19572), .B1(n19571), .B2(n19156), .ZN(
        n19148) );
  AOI22_X1 U22151 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19159), .B1(
        n19186), .B2(n19522), .ZN(n19147) );
  OAI211_X1 U22152 ( .C1(n19486), .C2(n19153), .A(n19148), .B(n19147), .ZN(
        P2_U3067) );
  AOI22_X1 U22153 ( .A1(n19157), .A2(n19578), .B1(n19577), .B2(n19156), .ZN(
        n19150) );
  AOI22_X1 U22154 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19159), .B1(
        n19186), .B2(n19525), .ZN(n19149) );
  OAI211_X1 U22155 ( .C1(n19492), .C2(n19153), .A(n19150), .B(n19149), .ZN(
        P2_U3068) );
  AOI22_X1 U22156 ( .A1(n19157), .A2(n19584), .B1(n19583), .B2(n19156), .ZN(
        n19152) );
  AOI22_X1 U22157 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19159), .B1(
        n19186), .B2(n19529), .ZN(n19151) );
  OAI211_X1 U22158 ( .C1(n19498), .C2(n19153), .A(n19152), .B(n19151), .ZN(
        P2_U3069) );
  AOI22_X1 U22159 ( .A1(n19157), .A2(n19590), .B1(n19589), .B2(n19156), .ZN(
        n19155) );
  AOI22_X1 U22160 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19159), .B1(
        n19158), .B2(n19591), .ZN(n19154) );
  OAI211_X1 U22161 ( .C1(n19594), .C2(n19194), .A(n19155), .B(n19154), .ZN(
        P2_U3070) );
  AOI22_X1 U22162 ( .A1(n19157), .A2(n19597), .B1(n19596), .B2(n19156), .ZN(
        n19161) );
  AOI22_X1 U22163 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19159), .B1(
        n19158), .B2(n19599), .ZN(n19160) );
  OAI211_X1 U22164 ( .C1(n19605), .C2(n19194), .A(n19161), .B(n19160), .ZN(
        P2_U3071) );
  NOR2_X1 U22165 ( .A1(n19163), .A2(n19165), .ZN(n19189) );
  AOI22_X1 U22166 ( .A1(n19555), .A2(n19186), .B1(n19547), .B2(n19189), .ZN(
        n19175) );
  INV_X1 U22167 ( .A(n19226), .ZN(n19164) );
  OAI21_X1 U22168 ( .B1(n19164), .B2(n19686), .A(n19685), .ZN(n19173) );
  NOR2_X1 U22169 ( .A1(n10862), .A2(n19165), .ZN(n19169) );
  INV_X1 U22170 ( .A(n19189), .ZN(n19166) );
  OAI211_X1 U22171 ( .C1(n19167), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19337), 
        .B(n19166), .ZN(n19168) );
  OAI211_X1 U22172 ( .C1(n19173), .C2(n19169), .A(n19549), .B(n19168), .ZN(
        n19191) );
  INV_X1 U22173 ( .A(n19169), .ZN(n19172) );
  OAI21_X1 U22174 ( .B1(n19170), .B2(n19189), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19171) );
  OAI21_X1 U22175 ( .B1(n19173), .B2(n19172), .A(n19171), .ZN(n19190) );
  AOI22_X1 U22176 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19191), .B1(
        n12991), .B2(n19190), .ZN(n19174) );
  OAI211_X1 U22177 ( .C1(n19558), .C2(n19224), .A(n19175), .B(n19174), .ZN(
        P2_U3072) );
  AOI22_X1 U22178 ( .A1(n19561), .A2(n19186), .B1(n19559), .B2(n19189), .ZN(
        n19177) );
  AOI22_X1 U22179 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19191), .B1(
        n19560), .B2(n19190), .ZN(n19176) );
  OAI211_X1 U22180 ( .C1(n19564), .C2(n19224), .A(n19177), .B(n19176), .ZN(
        P2_U3073) );
  AOI22_X1 U22181 ( .A1(n19518), .A2(n19216), .B1(n19189), .B2(n19565), .ZN(
        n19179) );
  AOI22_X1 U22182 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19191), .B1(
        n19566), .B2(n19190), .ZN(n19178) );
  OAI211_X1 U22183 ( .C1(n19480), .C2(n19194), .A(n19179), .B(n19178), .ZN(
        P2_U3074) );
  AOI22_X1 U22184 ( .A1(n19522), .A2(n19216), .B1(n19189), .B2(n19571), .ZN(
        n19181) );
  AOI22_X1 U22185 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19191), .B1(
        n19572), .B2(n19190), .ZN(n19180) );
  OAI211_X1 U22186 ( .C1(n19486), .C2(n19194), .A(n19181), .B(n19180), .ZN(
        P2_U3075) );
  AOI22_X1 U22187 ( .A1(n19579), .A2(n19186), .B1(n19577), .B2(n19189), .ZN(
        n19183) );
  AOI22_X1 U22188 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19191), .B1(
        n19578), .B2(n19190), .ZN(n19182) );
  OAI211_X1 U22189 ( .C1(n19582), .C2(n19224), .A(n19183), .B(n19182), .ZN(
        P2_U3076) );
  AOI22_X1 U22190 ( .A1(n19585), .A2(n19186), .B1(n19583), .B2(n19189), .ZN(
        n19185) );
  AOI22_X1 U22191 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19191), .B1(
        n19584), .B2(n19190), .ZN(n19184) );
  OAI211_X1 U22192 ( .C1(n19588), .C2(n19224), .A(n19185), .B(n19184), .ZN(
        P2_U3077) );
  AOI22_X1 U22193 ( .A1(n19591), .A2(n19186), .B1(n19189), .B2(n19589), .ZN(
        n19188) );
  AOI22_X1 U22194 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19191), .B1(
        n19590), .B2(n19190), .ZN(n19187) );
  OAI211_X1 U22195 ( .C1(n19594), .C2(n19224), .A(n19188), .B(n19187), .ZN(
        P2_U3078) );
  AOI22_X1 U22196 ( .A1(n19536), .A2(n19216), .B1(n19596), .B2(n19189), .ZN(
        n19193) );
  AOI22_X1 U22197 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19191), .B1(
        n19597), .B2(n19190), .ZN(n19192) );
  OAI211_X1 U22198 ( .C1(n19514), .C2(n19194), .A(n19193), .B(n19192), .ZN(
        P2_U3079) );
  NOR2_X1 U22199 ( .A1(n19196), .A2(n19195), .ZN(n19419) );
  NAND2_X1 U22200 ( .A1(n19419), .A2(n19697), .ZN(n19201) );
  INV_X1 U22201 ( .A(n11221), .ZN(n19197) );
  NAND3_X1 U22202 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n19697), .A3(
        n10862), .ZN(n19233) );
  NOR2_X1 U22203 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19233), .ZN(
        n19219) );
  OAI21_X1 U22204 ( .B1(n19197), .B2(n19219), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19198) );
  OAI21_X1 U22205 ( .B1(n19201), .B2(n19337), .A(n19198), .ZN(n19220) );
  AOI22_X1 U22206 ( .A1(n19220), .A2(n12991), .B1(n19547), .B2(n19219), .ZN(
        n19205) );
  AOI21_X1 U22207 ( .B1(n11221), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n19203) );
  OAI21_X1 U22208 ( .B1(n19216), .B2(n19247), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19200) );
  AOI21_X1 U22209 ( .B1(n19201), .B2(n19200), .A(n19426), .ZN(n19202) );
  AOI22_X1 U22210 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n19221), .B1(
        n19247), .B2(n19465), .ZN(n19204) );
  OAI211_X1 U22211 ( .C1(n19468), .C2(n19224), .A(n19205), .B(n19204), .ZN(
        P2_U3080) );
  AOI22_X1 U22212 ( .A1(n19220), .A2(n19560), .B1(n19559), .B2(n19219), .ZN(
        n19207) );
  AOI22_X1 U22213 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19221), .B1(
        n19216), .B2(n19561), .ZN(n19206) );
  OAI211_X1 U22214 ( .C1(n19564), .C2(n19254), .A(n19207), .B(n19206), .ZN(
        P2_U3081) );
  AOI22_X1 U22215 ( .A1(n19220), .A2(n19566), .B1(n19565), .B2(n19219), .ZN(
        n19209) );
  AOI22_X1 U22216 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19221), .B1(
        n19247), .B2(n19518), .ZN(n19208) );
  OAI211_X1 U22217 ( .C1(n19480), .C2(n19224), .A(n19209), .B(n19208), .ZN(
        P2_U3082) );
  AOI22_X1 U22218 ( .A1(n19220), .A2(n19572), .B1(n19571), .B2(n19219), .ZN(
        n19211) );
  AOI22_X1 U22219 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19221), .B1(
        n19247), .B2(n19522), .ZN(n19210) );
  OAI211_X1 U22220 ( .C1(n19486), .C2(n19224), .A(n19211), .B(n19210), .ZN(
        P2_U3083) );
  AOI22_X1 U22221 ( .A1(n19220), .A2(n19578), .B1(n19577), .B2(n19219), .ZN(
        n19213) );
  AOI22_X1 U22222 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19221), .B1(
        n19216), .B2(n19579), .ZN(n19212) );
  OAI211_X1 U22223 ( .C1(n19582), .C2(n19254), .A(n19213), .B(n19212), .ZN(
        P2_U3084) );
  AOI22_X1 U22224 ( .A1(n19220), .A2(n19584), .B1(n19583), .B2(n19219), .ZN(
        n19215) );
  AOI22_X1 U22225 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19221), .B1(
        n19247), .B2(n19529), .ZN(n19214) );
  OAI211_X1 U22226 ( .C1(n19498), .C2(n19224), .A(n19215), .B(n19214), .ZN(
        P2_U3085) );
  AOI22_X1 U22227 ( .A1(n19220), .A2(n19590), .B1(n19589), .B2(n19219), .ZN(
        n19218) );
  AOI22_X1 U22228 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19221), .B1(
        n19216), .B2(n19591), .ZN(n19217) );
  OAI211_X1 U22229 ( .C1(n19594), .C2(n19254), .A(n19218), .B(n19217), .ZN(
        P2_U3086) );
  AOI22_X1 U22230 ( .A1(n19220), .A2(n19597), .B1(n19596), .B2(n19219), .ZN(
        n19223) );
  AOI22_X1 U22231 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19221), .B1(
        n19247), .B2(n19536), .ZN(n19222) );
  OAI211_X1 U22232 ( .C1(n19514), .C2(n19224), .A(n19223), .B(n19222), .ZN(
        P2_U3087) );
  NOR2_X1 U22233 ( .A1(n19722), .A2(n19233), .ZN(n19260) );
  AOI22_X1 U22234 ( .A1(n19555), .A2(n19247), .B1(n19547), .B2(n19260), .ZN(
        n19236) );
  AOI21_X1 U22235 ( .B1(n19226), .B2(n19459), .A(n19337), .ZN(n19230) );
  INV_X1 U22236 ( .A(n19260), .ZN(n19227) );
  NAND2_X1 U22237 ( .A1(n11211), .A2(n19227), .ZN(n19231) );
  NOR2_X1 U22238 ( .A1(n19231), .A2(n19744), .ZN(n19228) );
  AOI21_X1 U22239 ( .B1(n19230), .B2(n19233), .A(n19228), .ZN(n19229) );
  OAI211_X1 U22240 ( .C1(n19260), .C2(n19714), .A(n19229), .B(n19549), .ZN(
        n19251) );
  INV_X1 U22241 ( .A(n19230), .ZN(n19234) );
  INV_X1 U22242 ( .A(n19231), .ZN(n19232) );
  OAI22_X1 U22243 ( .A1(n19234), .A2(n19233), .B1(n19232), .B2(n19744), .ZN(
        n19250) );
  AOI22_X1 U22244 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n19251), .B1(
        n12991), .B2(n19250), .ZN(n19235) );
  OAI211_X1 U22245 ( .C1(n19558), .C2(n19275), .A(n19236), .B(n19235), .ZN(
        P2_U3088) );
  AOI22_X1 U22246 ( .A1(n19561), .A2(n19247), .B1(n19559), .B2(n19260), .ZN(
        n19238) );
  AOI22_X1 U22247 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19251), .B1(
        n19560), .B2(n19250), .ZN(n19237) );
  OAI211_X1 U22248 ( .C1(n19564), .C2(n19275), .A(n19238), .B(n19237), .ZN(
        P2_U3089) );
  AOI22_X1 U22249 ( .A1(n19518), .A2(n19280), .B1(n19260), .B2(n19565), .ZN(
        n19240) );
  AOI22_X1 U22250 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19251), .B1(
        n19566), .B2(n19250), .ZN(n19239) );
  OAI211_X1 U22251 ( .C1(n19480), .C2(n19254), .A(n19240), .B(n19239), .ZN(
        P2_U3090) );
  AOI22_X1 U22252 ( .A1(n19522), .A2(n19280), .B1(n19260), .B2(n19571), .ZN(
        n19242) );
  AOI22_X1 U22253 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19251), .B1(
        n19572), .B2(n19250), .ZN(n19241) );
  OAI211_X1 U22254 ( .C1(n19486), .C2(n19254), .A(n19242), .B(n19241), .ZN(
        P2_U3091) );
  AOI22_X1 U22255 ( .A1(n19579), .A2(n19247), .B1(n19577), .B2(n19260), .ZN(
        n19244) );
  AOI22_X1 U22256 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19251), .B1(
        n19578), .B2(n19250), .ZN(n19243) );
  OAI211_X1 U22257 ( .C1(n19582), .C2(n19275), .A(n19244), .B(n19243), .ZN(
        P2_U3092) );
  AOI22_X1 U22258 ( .A1(n19585), .A2(n19247), .B1(n19583), .B2(n19260), .ZN(
        n19246) );
  AOI22_X1 U22259 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19251), .B1(
        n19584), .B2(n19250), .ZN(n19245) );
  OAI211_X1 U22260 ( .C1(n19588), .C2(n19275), .A(n19246), .B(n19245), .ZN(
        P2_U3093) );
  AOI22_X1 U22261 ( .A1(n19591), .A2(n19247), .B1(n19260), .B2(n19589), .ZN(
        n19249) );
  AOI22_X1 U22262 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19251), .B1(
        n19590), .B2(n19250), .ZN(n19248) );
  OAI211_X1 U22263 ( .C1(n19594), .C2(n19275), .A(n19249), .B(n19248), .ZN(
        P2_U3094) );
  AOI22_X1 U22264 ( .A1(n19536), .A2(n19280), .B1(n19596), .B2(n19260), .ZN(
        n19253) );
  AOI22_X1 U22265 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19251), .B1(
        n19597), .B2(n19250), .ZN(n19252) );
  OAI211_X1 U22266 ( .C1(n19514), .C2(n19254), .A(n19253), .B(n19252), .ZN(
        P2_U3095) );
  NOR2_X1 U22267 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19255), .ZN(
        n19278) );
  NOR2_X1 U22268 ( .A1(n19260), .A2(n19278), .ZN(n19258) );
  NOR3_X1 U22269 ( .A1(n19256), .A2(n19278), .A3(n19744), .ZN(n19261) );
  AOI211_X2 U22270 ( .C1(n19258), .C2(n19744), .A(n19257), .B(n19261), .ZN(
        n19279) );
  AOI22_X1 U22271 ( .A1(n19279), .A2(n12991), .B1(n19547), .B2(n19278), .ZN(
        n19264) );
  AOI21_X1 U22272 ( .B1(n19275), .B2(n19295), .A(n12954), .ZN(n19259) );
  AOI221_X1 U22273 ( .B1(n19714), .B2(n19260), .C1(n19714), .C2(n19259), .A(
        n19278), .ZN(n19262) );
  AOI22_X1 U22274 ( .A1(P2_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n19281), .B1(
        n19280), .B2(n19555), .ZN(n19263) );
  OAI211_X1 U22275 ( .C1(n19558), .C2(n19295), .A(n19264), .B(n19263), .ZN(
        P2_U3096) );
  AOI22_X1 U22276 ( .A1(n19279), .A2(n19560), .B1(n19559), .B2(n19278), .ZN(
        n19266) );
  AOI22_X1 U22277 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19281), .B1(
        n19280), .B2(n19561), .ZN(n19265) );
  OAI211_X1 U22278 ( .C1(n19564), .C2(n19295), .A(n19266), .B(n19265), .ZN(
        P2_U3097) );
  AOI22_X1 U22279 ( .A1(n19279), .A2(n19566), .B1(n19565), .B2(n19278), .ZN(
        n19268) );
  AOI22_X1 U22280 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19281), .B1(
        n19297), .B2(n19518), .ZN(n19267) );
  OAI211_X1 U22281 ( .C1(n19480), .C2(n19275), .A(n19268), .B(n19267), .ZN(
        P2_U3098) );
  AOI22_X1 U22282 ( .A1(n19279), .A2(n19572), .B1(n19571), .B2(n19278), .ZN(
        n19270) );
  AOI22_X1 U22283 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19281), .B1(
        n19297), .B2(n19522), .ZN(n19269) );
  OAI211_X1 U22284 ( .C1(n19486), .C2(n19275), .A(n19270), .B(n19269), .ZN(
        P2_U3099) );
  AOI22_X1 U22285 ( .A1(n19279), .A2(n19578), .B1(n19577), .B2(n19278), .ZN(
        n19272) );
  AOI22_X1 U22286 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19281), .B1(
        n19297), .B2(n19525), .ZN(n19271) );
  OAI211_X1 U22287 ( .C1(n19492), .C2(n19275), .A(n19272), .B(n19271), .ZN(
        P2_U3100) );
  AOI22_X1 U22288 ( .A1(n19279), .A2(n19584), .B1(n19583), .B2(n19278), .ZN(
        n19274) );
  AOI22_X1 U22289 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19281), .B1(
        n19297), .B2(n19529), .ZN(n19273) );
  OAI211_X1 U22290 ( .C1(n19498), .C2(n19275), .A(n19274), .B(n19273), .ZN(
        P2_U3101) );
  AOI22_X1 U22291 ( .A1(n19279), .A2(n19590), .B1(n19589), .B2(n19278), .ZN(
        n19277) );
  AOI22_X1 U22292 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19281), .B1(
        n19280), .B2(n19591), .ZN(n19276) );
  OAI211_X1 U22293 ( .C1(n19594), .C2(n19295), .A(n19277), .B(n19276), .ZN(
        P2_U3102) );
  AOI22_X1 U22294 ( .A1(n19279), .A2(n19597), .B1(n19596), .B2(n19278), .ZN(
        n19283) );
  AOI22_X1 U22295 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19281), .B1(
        n19280), .B2(n19599), .ZN(n19282) );
  OAI211_X1 U22296 ( .C1(n19605), .C2(n19295), .A(n19283), .B(n19282), .ZN(
        P2_U3103) );
  AOI22_X1 U22297 ( .A1(n19296), .A2(n19560), .B1(n19307), .B2(n19559), .ZN(
        n19285) );
  AOI22_X1 U22298 ( .A1(n19329), .A2(n19515), .B1(n19297), .B2(n19561), .ZN(
        n19284) );
  OAI211_X1 U22299 ( .C1(n19301), .C2(n20859), .A(n19285), .B(n19284), .ZN(
        P2_U3105) );
  AOI22_X1 U22300 ( .A1(n19296), .A2(n19566), .B1(n19307), .B2(n19565), .ZN(
        n19287) );
  AOI22_X1 U22301 ( .A1(n19329), .A2(n19518), .B1(n19297), .B2(n19567), .ZN(
        n19286) );
  OAI211_X1 U22302 ( .C1(n19301), .C2(n20774), .A(n19287), .B(n19286), .ZN(
        P2_U3106) );
  AOI22_X1 U22303 ( .A1(n19296), .A2(n19572), .B1(n19307), .B2(n19571), .ZN(
        n19289) );
  AOI22_X1 U22304 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19292), .B1(
        n19329), .B2(n19522), .ZN(n19288) );
  OAI211_X1 U22305 ( .C1(n19486), .C2(n19295), .A(n19289), .B(n19288), .ZN(
        P2_U3107) );
  AOI22_X1 U22306 ( .A1(n19296), .A2(n19578), .B1(n19307), .B2(n19577), .ZN(
        n19291) );
  AOI22_X1 U22307 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19292), .B1(
        n19329), .B2(n19525), .ZN(n19290) );
  OAI211_X1 U22308 ( .C1(n19492), .C2(n19295), .A(n19291), .B(n19290), .ZN(
        P2_U3108) );
  AOI22_X1 U22309 ( .A1(n19296), .A2(n19590), .B1(n19307), .B2(n19589), .ZN(
        n19294) );
  AOI22_X1 U22310 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19292), .B1(
        n19329), .B2(n19532), .ZN(n19293) );
  OAI211_X1 U22311 ( .C1(n19504), .C2(n19295), .A(n19294), .B(n19293), .ZN(
        P2_U3110) );
  AOI22_X1 U22312 ( .A1(n19296), .A2(n19597), .B1(n19307), .B2(n19596), .ZN(
        n19299) );
  AOI22_X1 U22313 ( .A1(n19329), .A2(n19536), .B1(n19297), .B2(n19599), .ZN(
        n19298) );
  OAI211_X1 U22314 ( .C1(n19301), .C2(n19300), .A(n19299), .B(n19298), .ZN(
        P2_U3111) );
  NAND2_X1 U22315 ( .A1(n19335), .A2(n10862), .ZN(n19346) );
  NOR2_X1 U22316 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19346), .ZN(
        n19328) );
  AOI22_X1 U22317 ( .A1(n19465), .A2(n19363), .B1(n19547), .B2(n19328), .ZN(
        n19314) );
  NOR3_X1 U22318 ( .A1(n19363), .A2(n19329), .A3(n19337), .ZN(n19304) );
  NOR2_X1 U22319 ( .A1(n19304), .A2(n19303), .ZN(n19312) );
  NOR2_X1 U22320 ( .A1(n19312), .A2(n19307), .ZN(n19305) );
  AOI211_X1 U22321 ( .C1(P2_STATE2_REG_2__SCAN_IN), .C2(n19308), .A(
        P2_STATE2_REG_3__SCAN_IN), .B(n19305), .ZN(n19306) );
  OAI21_X1 U22322 ( .B1(n19328), .B2(n19306), .A(n19549), .ZN(n19331) );
  NOR2_X1 U22323 ( .A1(n19307), .A2(n19328), .ZN(n19311) );
  INV_X1 U22324 ( .A(n19308), .ZN(n19309) );
  OAI21_X1 U22325 ( .B1(n19309), .B2(n19328), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19310) );
  AOI22_X1 U22326 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19331), .B1(
        n12991), .B2(n19330), .ZN(n19313) );
  OAI211_X1 U22327 ( .C1(n19468), .C2(n19325), .A(n19314), .B(n19313), .ZN(
        P2_U3112) );
  AOI22_X1 U22328 ( .A1(n19561), .A2(n19329), .B1(n19559), .B2(n19328), .ZN(
        n19316) );
  AOI22_X1 U22329 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19331), .B1(
        n19330), .B2(n19560), .ZN(n19315) );
  OAI211_X1 U22330 ( .C1(n19564), .C2(n19362), .A(n19316), .B(n19315), .ZN(
        P2_U3113) );
  AOI22_X1 U22331 ( .A1(n19518), .A2(n19363), .B1(n19328), .B2(n19565), .ZN(
        n19318) );
  AOI22_X1 U22332 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19331), .B1(
        n19330), .B2(n19566), .ZN(n19317) );
  OAI211_X1 U22333 ( .C1(n19480), .C2(n19325), .A(n19318), .B(n19317), .ZN(
        P2_U3114) );
  AOI22_X1 U22334 ( .A1(n19522), .A2(n19363), .B1(n19328), .B2(n19571), .ZN(
        n19320) );
  AOI22_X1 U22335 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19331), .B1(
        n19330), .B2(n19572), .ZN(n19319) );
  OAI211_X1 U22336 ( .C1(n19486), .C2(n19325), .A(n19320), .B(n19319), .ZN(
        P2_U3115) );
  AOI22_X1 U22337 ( .A1(n19525), .A2(n19363), .B1(n19328), .B2(n19577), .ZN(
        n19322) );
  AOI22_X1 U22338 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19331), .B1(
        n19330), .B2(n19578), .ZN(n19321) );
  OAI211_X1 U22339 ( .C1(n19492), .C2(n19325), .A(n19322), .B(n19321), .ZN(
        P2_U3116) );
  AOI22_X1 U22340 ( .A1(n19529), .A2(n19363), .B1(n19583), .B2(n19328), .ZN(
        n19324) );
  AOI22_X1 U22341 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19331), .B1(
        n19330), .B2(n19584), .ZN(n19323) );
  OAI211_X1 U22342 ( .C1(n19498), .C2(n19325), .A(n19324), .B(n19323), .ZN(
        P2_U3117) );
  AOI22_X1 U22343 ( .A1(n19591), .A2(n19329), .B1(n19328), .B2(n19589), .ZN(
        n19327) );
  AOI22_X1 U22344 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19331), .B1(
        n19330), .B2(n19590), .ZN(n19326) );
  OAI211_X1 U22345 ( .C1(n19594), .C2(n19362), .A(n19327), .B(n19326), .ZN(
        P2_U3118) );
  AOI22_X1 U22346 ( .A1(n19599), .A2(n19329), .B1(n19596), .B2(n19328), .ZN(
        n19333) );
  AOI22_X1 U22347 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19331), .B1(
        n19330), .B2(n19597), .ZN(n19332) );
  OAI211_X1 U22348 ( .C1(n19605), .C2(n19362), .A(n19333), .B(n19332), .ZN(
        P2_U3119) );
  INV_X1 U22349 ( .A(n19335), .ZN(n19372) );
  NOR2_X1 U22350 ( .A1(n19336), .A2(n19372), .ZN(n19373) );
  AOI22_X1 U22351 ( .A1(n19465), .A2(n19395), .B1(n19547), .B2(n19373), .ZN(
        n19349) );
  AOI21_X1 U22352 ( .B1(n19552), .B2(n19338), .A(n19337), .ZN(n19343) );
  INV_X1 U22353 ( .A(n19373), .ZN(n19339) );
  NAND2_X1 U22354 ( .A1(n19340), .A2(n19339), .ZN(n19344) );
  NOR2_X1 U22355 ( .A1(n19344), .A2(n19744), .ZN(n19341) );
  AOI21_X1 U22356 ( .B1(n19343), .B2(n19346), .A(n19341), .ZN(n19342) );
  OAI211_X1 U22357 ( .C1(n19373), .C2(n19714), .A(n19342), .B(n19549), .ZN(
        n19365) );
  INV_X1 U22358 ( .A(n19343), .ZN(n19347) );
  INV_X1 U22359 ( .A(n19344), .ZN(n19345) );
  OAI22_X1 U22360 ( .A1(n19347), .A2(n19346), .B1(n19345), .B2(n19744), .ZN(
        n19364) );
  AOI22_X1 U22361 ( .A1(P2_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n19365), .B1(
        n12991), .B2(n19364), .ZN(n19348) );
  OAI211_X1 U22362 ( .C1(n19468), .C2(n19362), .A(n19349), .B(n19348), .ZN(
        P2_U3120) );
  AOI22_X1 U22363 ( .A1(n19515), .A2(n19395), .B1(n19559), .B2(n19373), .ZN(
        n19351) );
  AOI22_X1 U22364 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19365), .B1(
        n19560), .B2(n19364), .ZN(n19350) );
  OAI211_X1 U22365 ( .C1(n19474), .C2(n19362), .A(n19351), .B(n19350), .ZN(
        P2_U3121) );
  AOI22_X1 U22366 ( .A1(n19567), .A2(n19363), .B1(n19373), .B2(n19565), .ZN(
        n19353) );
  AOI22_X1 U22367 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19365), .B1(
        n19566), .B2(n19364), .ZN(n19352) );
  OAI211_X1 U22368 ( .C1(n19570), .C2(n19390), .A(n19353), .B(n19352), .ZN(
        P2_U3122) );
  AOI22_X1 U22369 ( .A1(n19573), .A2(n19363), .B1(n19373), .B2(n19571), .ZN(
        n19355) );
  AOI22_X1 U22370 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19365), .B1(
        n19572), .B2(n19364), .ZN(n19354) );
  OAI211_X1 U22371 ( .C1(n19576), .C2(n19390), .A(n19355), .B(n19354), .ZN(
        P2_U3123) );
  AOI22_X1 U22372 ( .A1(n19525), .A2(n19395), .B1(n19577), .B2(n19373), .ZN(
        n19357) );
  AOI22_X1 U22373 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19365), .B1(
        n19578), .B2(n19364), .ZN(n19356) );
  OAI211_X1 U22374 ( .C1(n19492), .C2(n19362), .A(n19357), .B(n19356), .ZN(
        P2_U3124) );
  AOI22_X1 U22375 ( .A1(n19585), .A2(n19363), .B1(n19583), .B2(n19373), .ZN(
        n19359) );
  AOI22_X1 U22376 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19365), .B1(
        n19584), .B2(n19364), .ZN(n19358) );
  OAI211_X1 U22377 ( .C1(n19588), .C2(n19390), .A(n19359), .B(n19358), .ZN(
        P2_U3125) );
  AOI22_X1 U22378 ( .A1(n19532), .A2(n19395), .B1(n19373), .B2(n19589), .ZN(
        n19361) );
  AOI22_X1 U22379 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19365), .B1(
        n19590), .B2(n19364), .ZN(n19360) );
  OAI211_X1 U22380 ( .C1(n19504), .C2(n19362), .A(n19361), .B(n19360), .ZN(
        P2_U3126) );
  AOI22_X1 U22381 ( .A1(n19599), .A2(n19363), .B1(n19596), .B2(n19373), .ZN(
        n19367) );
  AOI22_X1 U22382 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19365), .B1(
        n19597), .B2(n19364), .ZN(n19366) );
  OAI211_X1 U22383 ( .C1(n19605), .C2(n19390), .A(n19367), .B(n19366), .ZN(
        P2_U3127) );
  INV_X1 U22384 ( .A(n19374), .ZN(n19369) );
  NOR2_X1 U22385 ( .A1(n19368), .A2(n19372), .ZN(n19393) );
  OAI21_X1 U22386 ( .B1(n19369), .B2(n19393), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19370) );
  OAI21_X1 U22387 ( .B1(n19372), .B2(n19371), .A(n19370), .ZN(n19394) );
  AOI22_X1 U22388 ( .A1(n19394), .A2(n12991), .B1(n19547), .B2(n19393), .ZN(
        n19379) );
  AOI221_X1 U22389 ( .B1(n19409), .B2(P2_STATEBS16_REG_SCAN_IN), .C1(n19395), 
        .C2(P2_STATEBS16_REG_SCAN_IN), .A(n19373), .ZN(n19375) );
  MUX2_X1 U22390 ( .A(n19375), .B(n19374), .S(P2_STATE2_REG_2__SCAN_IN), .Z(
        n19376) );
  NOR2_X1 U22391 ( .A1(n19376), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19377) );
  AOI22_X1 U22392 ( .A1(P2_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19396), .B1(
        n19409), .B2(n19465), .ZN(n19378) );
  OAI211_X1 U22393 ( .C1(n19468), .C2(n19390), .A(n19379), .B(n19378), .ZN(
        P2_U3128) );
  INV_X1 U22394 ( .A(n19409), .ZN(n19418) );
  AOI22_X1 U22395 ( .A1(n19394), .A2(n19560), .B1(n19559), .B2(n19393), .ZN(
        n19381) );
  AOI22_X1 U22396 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19396), .B1(
        n19395), .B2(n19561), .ZN(n19380) );
  OAI211_X1 U22397 ( .C1(n19564), .C2(n19418), .A(n19381), .B(n19380), .ZN(
        P2_U3129) );
  AOI22_X1 U22398 ( .A1(n19394), .A2(n19566), .B1(n19565), .B2(n19393), .ZN(
        n19383) );
  AOI22_X1 U22399 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19396), .B1(
        n19409), .B2(n19518), .ZN(n19382) );
  OAI211_X1 U22400 ( .C1(n19480), .C2(n19390), .A(n19383), .B(n19382), .ZN(
        P2_U3130) );
  AOI22_X1 U22401 ( .A1(n19394), .A2(n19572), .B1(n19571), .B2(n19393), .ZN(
        n19385) );
  AOI22_X1 U22402 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19396), .B1(
        n19409), .B2(n19522), .ZN(n19384) );
  OAI211_X1 U22403 ( .C1(n19486), .C2(n19390), .A(n19385), .B(n19384), .ZN(
        P2_U3131) );
  AOI22_X1 U22404 ( .A1(n19394), .A2(n19578), .B1(n19577), .B2(n19393), .ZN(
        n19387) );
  AOI22_X1 U22405 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19396), .B1(
        n19409), .B2(n19525), .ZN(n19386) );
  OAI211_X1 U22406 ( .C1(n19492), .C2(n19390), .A(n19387), .B(n19386), .ZN(
        P2_U3132) );
  AOI22_X1 U22407 ( .A1(n19394), .A2(n19584), .B1(n19583), .B2(n19393), .ZN(
        n19389) );
  AOI22_X1 U22408 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19396), .B1(
        n19409), .B2(n19529), .ZN(n19388) );
  OAI211_X1 U22409 ( .C1(n19498), .C2(n19390), .A(n19389), .B(n19388), .ZN(
        P2_U3133) );
  AOI22_X1 U22410 ( .A1(n19394), .A2(n19590), .B1(n19589), .B2(n19393), .ZN(
        n19392) );
  AOI22_X1 U22411 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19396), .B1(
        n19395), .B2(n19591), .ZN(n19391) );
  OAI211_X1 U22412 ( .C1(n19594), .C2(n19418), .A(n19392), .B(n19391), .ZN(
        P2_U3134) );
  AOI22_X1 U22413 ( .A1(n19394), .A2(n19597), .B1(n19596), .B2(n19393), .ZN(
        n19398) );
  AOI22_X1 U22414 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19396), .B1(
        n19395), .B2(n19599), .ZN(n19397) );
  OAI211_X1 U22415 ( .C1(n19605), .C2(n19418), .A(n19398), .B(n19397), .ZN(
        P2_U3135) );
  AOI22_X1 U22416 ( .A1(n19414), .A2(n19560), .B1(n19413), .B2(n19559), .ZN(
        n19400) );
  AOI22_X1 U22417 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19415), .B1(
        n19425), .B2(n19515), .ZN(n19399) );
  OAI211_X1 U22418 ( .C1(n19474), .C2(n19418), .A(n19400), .B(n19399), .ZN(
        P2_U3137) );
  AOI22_X1 U22419 ( .A1(n19414), .A2(n19566), .B1(n19413), .B2(n19565), .ZN(
        n19402) );
  AOI22_X1 U22420 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19415), .B1(
        n19409), .B2(n19567), .ZN(n19401) );
  OAI211_X1 U22421 ( .C1(n19570), .C2(n19450), .A(n19402), .B(n19401), .ZN(
        P2_U3138) );
  AOI22_X1 U22422 ( .A1(n19414), .A2(n19572), .B1(n19413), .B2(n19571), .ZN(
        n19404) );
  AOI22_X1 U22423 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19415), .B1(
        n19409), .B2(n19573), .ZN(n19403) );
  OAI211_X1 U22424 ( .C1(n19576), .C2(n19450), .A(n19404), .B(n19403), .ZN(
        P2_U3139) );
  AOI22_X1 U22425 ( .A1(n19414), .A2(n19578), .B1(n19413), .B2(n19577), .ZN(
        n19406) );
  AOI22_X1 U22426 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19415), .B1(
        n19409), .B2(n19579), .ZN(n19405) );
  OAI211_X1 U22427 ( .C1(n19582), .C2(n19450), .A(n19406), .B(n19405), .ZN(
        P2_U3140) );
  AOI22_X1 U22428 ( .A1(n19414), .A2(n19584), .B1(n19413), .B2(n19583), .ZN(
        n19408) );
  AOI22_X1 U22429 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19415), .B1(
        n19409), .B2(n19585), .ZN(n19407) );
  OAI211_X1 U22430 ( .C1(n19588), .C2(n19450), .A(n19408), .B(n19407), .ZN(
        P2_U3141) );
  AOI22_X1 U22431 ( .A1(n19414), .A2(n19590), .B1(n19413), .B2(n19589), .ZN(
        n19411) );
  AOI22_X1 U22432 ( .A1(n19409), .A2(n19591), .B1(n19425), .B2(n19532), .ZN(
        n19410) );
  OAI211_X1 U22433 ( .C1(n19412), .C2(n20775), .A(n19411), .B(n19410), .ZN(
        P2_U3142) );
  AOI22_X1 U22434 ( .A1(n19414), .A2(n19597), .B1(n19413), .B2(n19596), .ZN(
        n19417) );
  AOI22_X1 U22435 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19415), .B1(
        n19425), .B2(n19536), .ZN(n19416) );
  OAI211_X1 U22436 ( .C1(n19514), .C2(n19418), .A(n19417), .B(n19416), .ZN(
        P2_U3143) );
  NAND2_X1 U22437 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19419), .ZN(
        n19428) );
  OR2_X1 U22438 ( .A1(n19428), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19422) );
  INV_X1 U22439 ( .A(n19420), .ZN(n19421) );
  NOR2_X1 U22440 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19461), .ZN(
        n19445) );
  NOR3_X1 U22441 ( .A1(n19421), .A2(n19445), .A3(n19744), .ZN(n19427) );
  AOI21_X1 U22442 ( .B1(n19744), .B2(n19422), .A(n19427), .ZN(n19446) );
  AOI22_X1 U22443 ( .A1(n19446), .A2(n12991), .B1(n19547), .B2(n19445), .ZN(
        n19432) );
  OAI21_X1 U22444 ( .B1(n19425), .B2(n19451), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19429) );
  AOI211_X1 U22445 ( .C1(n19429), .C2(n19428), .A(n19427), .B(n19426), .ZN(
        n19430) );
  AOI22_X1 U22446 ( .A1(P2_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n19447), .B1(
        n19451), .B2(n19465), .ZN(n19431) );
  OAI211_X1 U22447 ( .C1(n19468), .C2(n19450), .A(n19432), .B(n19431), .ZN(
        P2_U3144) );
  AOI22_X1 U22448 ( .A1(n19446), .A2(n19560), .B1(n19559), .B2(n19445), .ZN(
        n19434) );
  AOI22_X1 U22449 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n19447), .B1(
        n19451), .B2(n19515), .ZN(n19433) );
  OAI211_X1 U22450 ( .C1(n19474), .C2(n19450), .A(n19434), .B(n19433), .ZN(
        P2_U3145) );
  AOI22_X1 U22451 ( .A1(n19446), .A2(n19566), .B1(n19565), .B2(n19445), .ZN(
        n19436) );
  AOI22_X1 U22452 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n19447), .B1(
        n19451), .B2(n19518), .ZN(n19435) );
  OAI211_X1 U22453 ( .C1(n19480), .C2(n19450), .A(n19436), .B(n19435), .ZN(
        P2_U3146) );
  AOI22_X1 U22454 ( .A1(n19446), .A2(n19572), .B1(n19571), .B2(n19445), .ZN(
        n19438) );
  AOI22_X1 U22455 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19447), .B1(
        n19451), .B2(n19522), .ZN(n19437) );
  OAI211_X1 U22456 ( .C1(n19486), .C2(n19450), .A(n19438), .B(n19437), .ZN(
        P2_U3147) );
  AOI22_X1 U22457 ( .A1(n19446), .A2(n19578), .B1(n19577), .B2(n19445), .ZN(
        n19440) );
  AOI22_X1 U22458 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n19447), .B1(
        n19451), .B2(n19525), .ZN(n19439) );
  OAI211_X1 U22459 ( .C1(n19492), .C2(n19450), .A(n19440), .B(n19439), .ZN(
        P2_U3148) );
  AOI22_X1 U22460 ( .A1(n19446), .A2(n19584), .B1(n19583), .B2(n19445), .ZN(
        n19442) );
  AOI22_X1 U22461 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19447), .B1(
        n19451), .B2(n19529), .ZN(n19441) );
  OAI211_X1 U22462 ( .C1(n19498), .C2(n19450), .A(n19442), .B(n19441), .ZN(
        P2_U3149) );
  AOI22_X1 U22463 ( .A1(n19446), .A2(n19590), .B1(n19589), .B2(n19445), .ZN(
        n19444) );
  AOI22_X1 U22464 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19447), .B1(
        n19451), .B2(n19532), .ZN(n19443) );
  OAI211_X1 U22465 ( .C1(n19504), .C2(n19450), .A(n19444), .B(n19443), .ZN(
        P2_U3150) );
  AOI22_X1 U22466 ( .A1(n19446), .A2(n19597), .B1(n19596), .B2(n19445), .ZN(
        n19449) );
  AOI22_X1 U22467 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n19447), .B1(
        n19451), .B2(n19536), .ZN(n19448) );
  OAI211_X1 U22468 ( .C1(n19514), .C2(n19450), .A(n19449), .B(n19448), .ZN(
        P2_U3151) );
  INV_X1 U22469 ( .A(n19464), .ZN(n19505) );
  AND2_X1 U22470 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19505), .ZN(n19452) );
  AND2_X1 U22471 ( .A1(n19453), .A2(n19452), .ZN(n19460) );
  INV_X1 U22472 ( .A(n19461), .ZN(n19454) );
  AOI21_X1 U22473 ( .B1(n19714), .B2(n19454), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19455) );
  OAI22_X1 U22474 ( .A1(n19508), .A2(n19457), .B1(n19456), .B2(n19505), .ZN(
        n19458) );
  INV_X1 U22475 ( .A(n19458), .ZN(n19467) );
  NAND2_X1 U22476 ( .A1(n19552), .A2(n19459), .ZN(n19462) );
  AOI21_X1 U22477 ( .B1(n19462), .B2(n19461), .A(n19460), .ZN(n19463) );
  OAI211_X1 U22478 ( .C1(n19464), .C2(n19714), .A(n19463), .B(n19549), .ZN(
        n19510) );
  AOI22_X1 U22479 ( .A1(P2_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n19510), .B1(
        n19537), .B2(n19465), .ZN(n19466) );
  OAI211_X1 U22480 ( .C1(n19468), .C2(n19513), .A(n19467), .B(n19466), .ZN(
        P2_U3152) );
  OAI22_X1 U22481 ( .A1(n19508), .A2(n19470), .B1(n19469), .B2(n19505), .ZN(
        n19471) );
  INV_X1 U22482 ( .A(n19471), .ZN(n19473) );
  AOI22_X1 U22483 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19510), .B1(
        n19537), .B2(n19515), .ZN(n19472) );
  OAI211_X1 U22484 ( .C1(n19474), .C2(n19513), .A(n19473), .B(n19472), .ZN(
        P2_U3153) );
  OAI22_X1 U22485 ( .A1(n19508), .A2(n19476), .B1(n19475), .B2(n19505), .ZN(
        n19477) );
  INV_X1 U22486 ( .A(n19477), .ZN(n19479) );
  AOI22_X1 U22487 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19510), .B1(
        n19537), .B2(n19518), .ZN(n19478) );
  OAI211_X1 U22488 ( .C1(n19480), .C2(n19513), .A(n19479), .B(n19478), .ZN(
        P2_U3154) );
  OAI22_X1 U22489 ( .A1(n19508), .A2(n19482), .B1(n19481), .B2(n19505), .ZN(
        n19483) );
  INV_X1 U22490 ( .A(n19483), .ZN(n19485) );
  AOI22_X1 U22491 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19510), .B1(
        n19537), .B2(n19522), .ZN(n19484) );
  OAI211_X1 U22492 ( .C1(n19486), .C2(n19513), .A(n19485), .B(n19484), .ZN(
        P2_U3155) );
  OAI22_X1 U22493 ( .A1(n19508), .A2(n19488), .B1(n19487), .B2(n19505), .ZN(
        n19489) );
  INV_X1 U22494 ( .A(n19489), .ZN(n19491) );
  AOI22_X1 U22495 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19510), .B1(
        n19537), .B2(n19525), .ZN(n19490) );
  OAI211_X1 U22496 ( .C1(n19492), .C2(n19513), .A(n19491), .B(n19490), .ZN(
        P2_U3156) );
  OAI22_X1 U22497 ( .A1(n19508), .A2(n19494), .B1(n19493), .B2(n19505), .ZN(
        n19495) );
  INV_X1 U22498 ( .A(n19495), .ZN(n19497) );
  AOI22_X1 U22499 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19510), .B1(
        n19537), .B2(n19529), .ZN(n19496) );
  OAI211_X1 U22500 ( .C1(n19498), .C2(n19513), .A(n19497), .B(n19496), .ZN(
        P2_U3157) );
  OAI22_X1 U22501 ( .A1(n19508), .A2(n19500), .B1(n19499), .B2(n19505), .ZN(
        n19501) );
  INV_X1 U22502 ( .A(n19501), .ZN(n19503) );
  AOI22_X1 U22503 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19510), .B1(
        n19537), .B2(n19532), .ZN(n19502) );
  OAI211_X1 U22504 ( .C1(n19504), .C2(n19513), .A(n19503), .B(n19502), .ZN(
        P2_U3158) );
  OAI22_X1 U22505 ( .A1(n19508), .A2(n19507), .B1(n19506), .B2(n19505), .ZN(
        n19509) );
  INV_X1 U22506 ( .A(n19509), .ZN(n19512) );
  AOI22_X1 U22507 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19510), .B1(
        n19537), .B2(n19536), .ZN(n19511) );
  OAI211_X1 U22508 ( .C1(n19514), .C2(n19513), .A(n19512), .B(n19511), .ZN(
        P2_U3159) );
  AOI22_X1 U22509 ( .A1(n19515), .A2(n19600), .B1(n19535), .B2(n19559), .ZN(
        n19517) );
  AOI22_X1 U22510 ( .A1(n19560), .A2(n19538), .B1(n19537), .B2(n19561), .ZN(
        n19516) );
  OAI211_X1 U22511 ( .C1(n19542), .C2(n20884), .A(n19517), .B(n19516), .ZN(
        P2_U3161) );
  INV_X1 U22512 ( .A(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n19521) );
  AOI22_X1 U22513 ( .A1(n19518), .A2(n19600), .B1(n19535), .B2(n19565), .ZN(
        n19520) );
  AOI22_X1 U22514 ( .A1(n19566), .A2(n19538), .B1(n19537), .B2(n19567), .ZN(
        n19519) );
  OAI211_X1 U22515 ( .C1(n19542), .C2(n19521), .A(n19520), .B(n19519), .ZN(
        P2_U3162) );
  AOI22_X1 U22516 ( .A1(n19573), .A2(n19537), .B1(n19535), .B2(n19571), .ZN(
        n19524) );
  AOI22_X1 U22517 ( .A1(n19572), .A2(n19538), .B1(n19600), .B2(n19522), .ZN(
        n19523) );
  OAI211_X1 U22518 ( .C1(n19542), .C2(n11174), .A(n19524), .B(n19523), .ZN(
        P2_U3163) );
  AOI22_X1 U22519 ( .A1(n19579), .A2(n19537), .B1(n19535), .B2(n19577), .ZN(
        n19527) );
  AOI22_X1 U22520 ( .A1(n19578), .A2(n19538), .B1(n19600), .B2(n19525), .ZN(
        n19526) );
  OAI211_X1 U22521 ( .C1(n19542), .C2(n19528), .A(n19527), .B(n19526), .ZN(
        P2_U3164) );
  AOI22_X1 U22522 ( .A1(n19529), .A2(n19600), .B1(n19583), .B2(n19535), .ZN(
        n19531) );
  AOI22_X1 U22523 ( .A1(n19584), .A2(n19538), .B1(n19537), .B2(n19585), .ZN(
        n19530) );
  OAI211_X1 U22524 ( .C1(n19542), .C2(n11201), .A(n19531), .B(n19530), .ZN(
        P2_U3165) );
  AOI22_X1 U22525 ( .A1(n19532), .A2(n19600), .B1(n19535), .B2(n19589), .ZN(
        n19534) );
  AOI22_X1 U22526 ( .A1(n19590), .A2(n19538), .B1(n19537), .B2(n19591), .ZN(
        n19533) );
  OAI211_X1 U22527 ( .C1(n19542), .C2(n11274), .A(n19534), .B(n19533), .ZN(
        P2_U3166) );
  INV_X1 U22528 ( .A(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n19541) );
  AOI22_X1 U22529 ( .A1(n19536), .A2(n19600), .B1(n19535), .B2(n19596), .ZN(
        n19540) );
  AOI22_X1 U22530 ( .A1(n19597), .A2(n19538), .B1(n19537), .B2(n19599), .ZN(
        n19539) );
  OAI211_X1 U22531 ( .C1(n19542), .C2(n19541), .A(n19540), .B(n19539), .ZN(
        P2_U3167) );
  NOR2_X1 U22532 ( .A1(n19595), .A2(n19744), .ZN(n19543) );
  NAND2_X1 U22533 ( .A1(n11204), .A2(n19543), .ZN(n19548) );
  NOR2_X1 U22534 ( .A1(n19697), .A2(n19544), .ZN(n19554) );
  INV_X1 U22535 ( .A(n19554), .ZN(n19545) );
  OAI21_X1 U22536 ( .B1(n19545), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n19744), 
        .ZN(n19546) );
  AND2_X1 U22537 ( .A1(n19548), .A2(n19546), .ZN(n19598) );
  AOI22_X1 U22538 ( .A1(n19598), .A2(n12991), .B1(n19547), .B2(n19595), .ZN(
        n19557) );
  OAI211_X1 U22539 ( .C1(n19595), .C2(n19714), .A(n19549), .B(n19548), .ZN(
        n19550) );
  INV_X1 U22540 ( .A(n19550), .ZN(n19551) );
  OAI221_X1 U22541 ( .B1(n19554), .B2(n19553), .C1(n19554), .C2(n19552), .A(
        n19551), .ZN(n19601) );
  AOI22_X1 U22542 ( .A1(P2_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n19601), .B1(
        n19600), .B2(n19555), .ZN(n19556) );
  OAI211_X1 U22543 ( .C1(n19558), .C2(n19604), .A(n19557), .B(n19556), .ZN(
        P2_U3168) );
  AOI22_X1 U22544 ( .A1(n19598), .A2(n19560), .B1(n19559), .B2(n19595), .ZN(
        n19563) );
  AOI22_X1 U22545 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n19601), .B1(
        n19600), .B2(n19561), .ZN(n19562) );
  OAI211_X1 U22546 ( .C1(n19564), .C2(n19604), .A(n19563), .B(n19562), .ZN(
        P2_U3169) );
  AOI22_X1 U22547 ( .A1(n19598), .A2(n19566), .B1(n19565), .B2(n19595), .ZN(
        n19569) );
  AOI22_X1 U22548 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n19601), .B1(
        n19600), .B2(n19567), .ZN(n19568) );
  OAI211_X1 U22549 ( .C1(n19570), .C2(n19604), .A(n19569), .B(n19568), .ZN(
        P2_U3170) );
  AOI22_X1 U22550 ( .A1(n19598), .A2(n19572), .B1(n19571), .B2(n19595), .ZN(
        n19575) );
  AOI22_X1 U22551 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n19601), .B1(
        n19600), .B2(n19573), .ZN(n19574) );
  OAI211_X1 U22552 ( .C1(n19576), .C2(n19604), .A(n19575), .B(n19574), .ZN(
        P2_U3171) );
  AOI22_X1 U22553 ( .A1(n19598), .A2(n19578), .B1(n19577), .B2(n19595), .ZN(
        n19581) );
  AOI22_X1 U22554 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n19601), .B1(
        n19600), .B2(n19579), .ZN(n19580) );
  OAI211_X1 U22555 ( .C1(n19582), .C2(n19604), .A(n19581), .B(n19580), .ZN(
        P2_U3172) );
  AOI22_X1 U22556 ( .A1(n19598), .A2(n19584), .B1(n19583), .B2(n19595), .ZN(
        n19587) );
  AOI22_X1 U22557 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19601), .B1(
        n19600), .B2(n19585), .ZN(n19586) );
  OAI211_X1 U22558 ( .C1(n19588), .C2(n19604), .A(n19587), .B(n19586), .ZN(
        P2_U3173) );
  AOI22_X1 U22559 ( .A1(n19598), .A2(n19590), .B1(n19589), .B2(n19595), .ZN(
        n19593) );
  AOI22_X1 U22560 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19601), .B1(
        n19600), .B2(n19591), .ZN(n19592) );
  OAI211_X1 U22561 ( .C1(n19594), .C2(n19604), .A(n19593), .B(n19592), .ZN(
        P2_U3174) );
  AOI22_X1 U22562 ( .A1(n19598), .A2(n19597), .B1(n19596), .B2(n19595), .ZN(
        n19603) );
  AOI22_X1 U22563 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n19601), .B1(
        n19600), .B2(n19599), .ZN(n19602) );
  OAI211_X1 U22564 ( .C1(n19605), .C2(n19604), .A(n19603), .B(n19602), .ZN(
        P2_U3175) );
  NAND3_X1 U22565 ( .A1(n19736), .A2(n19606), .A3(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n19608) );
  NAND2_X1 U22566 ( .A1(n19608), .A2(n19607), .ZN(n19612) );
  NAND2_X1 U22567 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n19745), .ZN(n19609) );
  AOI21_X1 U22568 ( .B1(n19610), .B2(n19613), .A(n19609), .ZN(n19611) );
  AOI21_X1 U22569 ( .B1(n19613), .B2(n19612), .A(n19611), .ZN(n19615) );
  NAND2_X1 U22570 ( .A1(n19615), .A2(n19614), .ZN(P2_U3177) );
  AND2_X1 U22571 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n19616), .ZN(
        P2_U3179) );
  AND2_X1 U22572 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n19616), .ZN(
        P2_U3180) );
  AND2_X1 U22573 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n19616), .ZN(
        P2_U3181) );
  AND2_X1 U22574 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n19616), .ZN(
        P2_U3182) );
  AND2_X1 U22575 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n19616), .ZN(
        P2_U3183) );
  AND2_X1 U22576 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n19616), .ZN(
        P2_U3184) );
  AND2_X1 U22577 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n19616), .ZN(
        P2_U3185) );
  AND2_X1 U22578 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n19616), .ZN(
        P2_U3186) );
  AND2_X1 U22579 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n19616), .ZN(
        P2_U3187) );
  AND2_X1 U22580 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n19616), .ZN(
        P2_U3188) );
  AND2_X1 U22581 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n19616), .ZN(
        P2_U3189) );
  AND2_X1 U22582 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n19616), .ZN(
        P2_U3190) );
  AND2_X1 U22583 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n19616), .ZN(
        P2_U3191) );
  AND2_X1 U22584 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n19616), .ZN(
        P2_U3192) );
  AND2_X1 U22585 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n19616), .ZN(
        P2_U3193) );
  AND2_X1 U22586 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n19616), .ZN(
        P2_U3194) );
  AND2_X1 U22587 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n19616), .ZN(
        P2_U3195) );
  AND2_X1 U22588 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n19616), .ZN(
        P2_U3196) );
  AND2_X1 U22589 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n19616), .ZN(
        P2_U3197) );
  AND2_X1 U22590 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n19616), .ZN(
        P2_U3198) );
  AND2_X1 U22591 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n19616), .ZN(
        P2_U3199) );
  AND2_X1 U22592 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n19616), .ZN(
        P2_U3200) );
  AND2_X1 U22593 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n19616), .ZN(P2_U3201) );
  AND2_X1 U22594 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n19616), .ZN(P2_U3202) );
  AND2_X1 U22595 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n19616), .ZN(P2_U3203) );
  INV_X1 U22596 ( .A(P2_DATAWIDTH_REG_6__SCAN_IN), .ZN(n20724) );
  NOR2_X1 U22597 ( .A1(n20724), .A2(n19683), .ZN(P2_U3204) );
  AND2_X1 U22598 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n19616), .ZN(P2_U3205) );
  AND2_X1 U22599 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n19616), .ZN(P2_U3206) );
  AND2_X1 U22600 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n19616), .ZN(P2_U3207) );
  AND2_X1 U22601 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n19616), .ZN(P2_U3208) );
  INV_X1 U22602 ( .A(P2_STATE_REG_1__SCAN_IN), .ZN(n19626) );
  NOR2_X1 U22603 ( .A1(n19736), .A2(n19626), .ZN(n19624) );
  INV_X1 U22604 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n19751) );
  OR3_X1 U22605 ( .A1(n19624), .A2(n19751), .A3(n19617), .ZN(n19619) );
  INV_X2 U22606 ( .A(n19753), .ZN(n19665) );
  AOI211_X1 U22607 ( .C1(n20581), .C2(P2_REQUESTPENDING_REG_SCAN_IN), .A(
        n19625), .B(n19665), .ZN(n19618) );
  NOR3_X1 U22608 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(P2_STATE_REG_1__SCAN_IN), 
        .A3(n20589), .ZN(n19630) );
  AOI211_X1 U22609 ( .C1(n19633), .C2(n19619), .A(n19618), .B(n19630), .ZN(
        n19620) );
  INV_X1 U22610 ( .A(n19620), .ZN(P2_U3209) );
  AOI21_X1 U22611 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(n20581), .A(n19633), 
        .ZN(n19627) );
  NOR3_X1 U22612 ( .A1(n19617), .A2(n19627), .A3(n19751), .ZN(n19621) );
  NOR3_X1 U22613 ( .A1(n19741), .A2(n19624), .A3(n19621), .ZN(n19622) );
  OAI21_X1 U22614 ( .B1(n20581), .B2(n19623), .A(n19622), .ZN(P2_U3210) );
  AOI22_X1 U22615 ( .A1(n19625), .A2(n19751), .B1(n19624), .B2(n20589), .ZN(
        n19632) );
  OAI21_X1 U22616 ( .B1(P2_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .A(
        P2_STATE_REG_0__SCAN_IN), .ZN(n19631) );
  NOR2_X1 U22617 ( .A1(n19626), .A2(n19633), .ZN(n19628) );
  AOI21_X1 U22618 ( .B1(n19628), .B2(n19745), .A(n19627), .ZN(n19629) );
  OAI22_X1 U22619 ( .A1(n19632), .A2(n19631), .B1(n19630), .B2(n19629), .ZN(
        P2_U3211) );
  NAND2_X1 U22620 ( .A1(n19665), .A2(n19633), .ZN(n19673) );
  CLKBUF_X1 U22621 ( .A(n19673), .Z(n19668) );
  OAI222_X1 U22622 ( .A1(n19669), .A2(n13175), .B1(n19634), .B2(n19665), .C1(
        n11958), .C2(n19668), .ZN(P2_U3212) );
  OAI222_X1 U22623 ( .A1(n19669), .A2(n11958), .B1(n19635), .B2(n19665), .C1(
        n11002), .C2(n19668), .ZN(P2_U3213) );
  OAI222_X1 U22624 ( .A1(n19669), .A2(n11002), .B1(n19636), .B2(n19665), .C1(
        n11551), .C2(n19668), .ZN(P2_U3214) );
  OAI222_X1 U22625 ( .A1(n19668), .A2(n11557), .B1(n19637), .B2(n19665), .C1(
        n11551), .C2(n19669), .ZN(P2_U3215) );
  OAI222_X1 U22626 ( .A1(n19673), .A2(n11564), .B1(n19638), .B2(n19665), .C1(
        n11557), .C2(n19669), .ZN(P2_U3216) );
  OAI222_X1 U22627 ( .A1(n19673), .A2(n11570), .B1(n19639), .B2(n19665), .C1(
        n11564), .C2(n19669), .ZN(P2_U3217) );
  OAI222_X1 U22628 ( .A1(n19673), .A2(n11576), .B1(n20804), .B2(n19665), .C1(
        n11570), .C2(n19669), .ZN(P2_U3218) );
  OAI222_X1 U22629 ( .A1(n19673), .A2(n11579), .B1(n19640), .B2(n19665), .C1(
        n11576), .C2(n19669), .ZN(P2_U3219) );
  OAI222_X1 U22630 ( .A1(n19673), .A2(n11585), .B1(n19641), .B2(n19665), .C1(
        n11579), .C2(n19669), .ZN(P2_U3220) );
  OAI222_X1 U22631 ( .A1(n19668), .A2(n11591), .B1(n19642), .B2(n19665), .C1(
        n11585), .C2(n19669), .ZN(P2_U3221) );
  OAI222_X1 U22632 ( .A1(n19668), .A2(n11594), .B1(n20729), .B2(n19665), .C1(
        n11591), .C2(n19669), .ZN(P2_U3222) );
  OAI222_X1 U22633 ( .A1(n19668), .A2(n11602), .B1(n19643), .B2(n19665), .C1(
        n11594), .C2(n19669), .ZN(P2_U3223) );
  OAI222_X1 U22634 ( .A1(n19668), .A2(n11608), .B1(n19644), .B2(n19665), .C1(
        n11602), .C2(n19669), .ZN(P2_U3224) );
  OAI222_X1 U22635 ( .A1(n19668), .A2(n11611), .B1(n19645), .B2(n19665), .C1(
        n11608), .C2(n19669), .ZN(P2_U3225) );
  OAI222_X1 U22636 ( .A1(n19668), .A2(n19647), .B1(n19646), .B2(n19665), .C1(
        n11611), .C2(n19669), .ZN(P2_U3226) );
  OAI222_X1 U22637 ( .A1(n19673), .A2(n11622), .B1(n19648), .B2(n19665), .C1(
        n19647), .C2(n19669), .ZN(P2_U3227) );
  OAI222_X1 U22638 ( .A1(n19673), .A2(n19650), .B1(n19649), .B2(n19665), .C1(
        n11622), .C2(n19669), .ZN(P2_U3228) );
  OAI222_X1 U22639 ( .A1(n19673), .A2(n11628), .B1(n19651), .B2(n19665), .C1(
        n19650), .C2(n19669), .ZN(P2_U3229) );
  OAI222_X1 U22640 ( .A1(n19673), .A2(n20777), .B1(n19652), .B2(n19665), .C1(
        n11628), .C2(n19669), .ZN(P2_U3230) );
  OAI222_X1 U22641 ( .A1(n19673), .A2(n19654), .B1(n19653), .B2(n19665), .C1(
        n20777), .C2(n19669), .ZN(P2_U3231) );
  OAI222_X1 U22642 ( .A1(n19673), .A2(n19656), .B1(n19655), .B2(n19665), .C1(
        n19654), .C2(n19669), .ZN(P2_U3232) );
  OAI222_X1 U22643 ( .A1(n19668), .A2(n11641), .B1(n19657), .B2(n19665), .C1(
        n19656), .C2(n19669), .ZN(P2_U3233) );
  OAI222_X1 U22644 ( .A1(n19668), .A2(n19659), .B1(n19658), .B2(n19665), .C1(
        n11641), .C2(n19669), .ZN(P2_U3234) );
  OAI222_X1 U22645 ( .A1(n19668), .A2(n11646), .B1(n19660), .B2(n19665), .C1(
        n19659), .C2(n19669), .ZN(P2_U3235) );
  OAI222_X1 U22646 ( .A1(n19668), .A2(n20880), .B1(n19661), .B2(n19665), .C1(
        n11646), .C2(n19669), .ZN(P2_U3236) );
  OAI222_X1 U22647 ( .A1(n19668), .A2(n14759), .B1(n19662), .B2(n19665), .C1(
        n20880), .C2(n19669), .ZN(P2_U3237) );
  OAI222_X1 U22648 ( .A1(n19669), .A2(n14759), .B1(n19663), .B2(n19665), .C1(
        n19664), .C2(n19668), .ZN(P2_U3238) );
  OAI222_X1 U22649 ( .A1(n19668), .A2(n14733), .B1(n19666), .B2(n19665), .C1(
        n19664), .C2(n19669), .ZN(P2_U3239) );
  OAI222_X1 U22650 ( .A1(n19668), .A2(n19670), .B1(n19667), .B2(n19665), .C1(
        n14733), .C2(n19669), .ZN(P2_U3240) );
  INV_X1 U22651 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n19671) );
  OAI222_X1 U22652 ( .A1(n19673), .A2(n19672), .B1(n19671), .B2(n19665), .C1(
        n19670), .C2(n19669), .ZN(P2_U3241) );
  INV_X1 U22653 ( .A(P2_BE_N_REG_3__SCAN_IN), .ZN(n19674) );
  AOI22_X1 U22654 ( .A1(n19665), .A2(n19675), .B1(n19674), .B2(n19753), .ZN(
        P2_U3585) );
  MUX2_X1 U22655 ( .A(P2_BE_N_REG_2__SCAN_IN), .B(P2_BYTEENABLE_REG_2__SCAN_IN), .S(n19665), .Z(P2_U3586) );
  INV_X1 U22656 ( .A(P2_BE_N_REG_1__SCAN_IN), .ZN(n19676) );
  AOI22_X1 U22657 ( .A1(n19665), .A2(n19677), .B1(n19676), .B2(n19753), .ZN(
        P2_U3587) );
  INV_X1 U22658 ( .A(P2_BE_N_REG_0__SCAN_IN), .ZN(n19678) );
  AOI22_X1 U22659 ( .A1(n19665), .A2(n19679), .B1(n19678), .B2(n19753), .ZN(
        P2_U3588) );
  OAI21_X1 U22660 ( .B1(n19683), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .A(n19681), 
        .ZN(n19680) );
  INV_X1 U22661 ( .A(n19680), .ZN(P2_U3591) );
  OAI21_X1 U22662 ( .B1(n19683), .B2(n19682), .A(n19681), .ZN(P2_U3592) );
  NAND2_X1 U22663 ( .A1(n19684), .A2(n19685), .ZN(n19695) );
  NAND2_X1 U22664 ( .A1(n19685), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19709) );
  OR2_X1 U22665 ( .A1(n19686), .A2(n19709), .ZN(n19698) );
  NAND2_X1 U22666 ( .A1(n19687), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19688) );
  OR2_X1 U22667 ( .A1(n19707), .A2(n19688), .ZN(n19689) );
  NAND2_X1 U22668 ( .A1(n19689), .A2(n19705), .ZN(n19699) );
  NAND2_X1 U22669 ( .A1(n19698), .A2(n19699), .ZN(n19691) );
  NAND2_X1 U22670 ( .A1(n19691), .A2(n19690), .ZN(n19694) );
  NAND2_X1 U22671 ( .A1(n19692), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19693) );
  AND3_X1 U22672 ( .A1(n19695), .A2(n19694), .A3(n19693), .ZN(n19696) );
  AOI22_X1 U22673 ( .A1(n19723), .A2(n19697), .B1(n19696), .B2(n19720), .ZN(
        P2_U3602) );
  OAI21_X1 U22674 ( .B1(n19700), .B2(n19699), .A(n19698), .ZN(n19701) );
  AOI21_X1 U22675 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19702), .A(n19701), 
        .ZN(n19703) );
  AOI22_X1 U22676 ( .A1(n19723), .A2(n19704), .B1(n19703), .B2(n19720), .ZN(
        P2_U3603) );
  INV_X1 U22677 ( .A(n19705), .ZN(n19715) );
  OR3_X1 U22678 ( .A1(n19707), .A2(n19715), .A3(n19706), .ZN(n19708) );
  OAI21_X1 U22679 ( .B1(n19710), .B2(n19709), .A(n19708), .ZN(n19711) );
  AOI21_X1 U22680 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19712), .A(n19711), 
        .ZN(n19713) );
  AOI22_X1 U22681 ( .A1(n19723), .A2(n10862), .B1(n19713), .B2(n19720), .ZN(
        P2_U3604) );
  OAI22_X1 U22682 ( .A1(n19716), .A2(n19715), .B1(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n19714), .ZN(n19717) );
  AOI21_X1 U22683 ( .B1(n19719), .B2(n19718), .A(n19717), .ZN(n19721) );
  AOI22_X1 U22684 ( .A1(n19723), .A2(n19722), .B1(n19721), .B2(n19720), .ZN(
        P2_U3605) );
  INV_X1 U22685 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n20808) );
  AOI22_X1 U22686 ( .A1(n19665), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n20808), 
        .B2(n19753), .ZN(P2_U3608) );
  INV_X1 U22687 ( .A(n19724), .ZN(n19725) );
  NOR2_X1 U22688 ( .A1(n19726), .A2(n19725), .ZN(n19728) );
  AOI211_X1 U22689 ( .C1(n19730), .C2(n19729), .A(n19728), .B(n19727), .ZN(
        n19732) );
  INV_X1 U22690 ( .A(P2_MORE_REG_SCAN_IN), .ZN(n20933) );
  INV_X1 U22691 ( .A(n19733), .ZN(n19731) );
  AOI22_X1 U22692 ( .A1(n19733), .A2(n19732), .B1(n20933), .B2(n19731), .ZN(
        P2_U3609) );
  NOR2_X1 U22693 ( .A1(n19734), .A2(n19744), .ZN(n19738) );
  AOI21_X1 U22694 ( .B1(n19017), .B2(n19736), .A(n19735), .ZN(n19737) );
  OAI21_X1 U22695 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19738), .A(n19737), 
        .ZN(n19752) );
  AOI21_X1 U22696 ( .B1(n19741), .B2(P2_STATEBS16_REG_SCAN_IN), .A(n19739), 
        .ZN(n19743) );
  NOR3_X1 U22697 ( .A1(n19741), .A2(n19740), .A3(n18954), .ZN(n19742) );
  MUX2_X1 U22698 ( .A(n19743), .B(n19742), .S(n10944), .Z(n19749) );
  OAI22_X1 U22699 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19746), .B1(n19745), 
        .B2(n19744), .ZN(n19747) );
  INV_X1 U22700 ( .A(n19747), .ZN(n19748) );
  OAI21_X1 U22701 ( .B1(n19749), .B2(n19748), .A(n19752), .ZN(n19750) );
  OAI21_X1 U22702 ( .B1(n19752), .B2(n19751), .A(n19750), .ZN(P2_U3610) );
  INV_X1 U22703 ( .A(P2_M_IO_N_REG_SCAN_IN), .ZN(n20928) );
  AOI22_X1 U22704 ( .A1(n19665), .A2(n19754), .B1(n20928), .B2(n19753), .ZN(
        P2_U3611) );
  AOI21_X1 U22705 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n20597), .A(n20585), 
        .ZN(n19762) );
  INV_X1 U22706 ( .A(P1_ADS_N_REG_SCAN_IN), .ZN(n19756) );
  INV_X2 U22707 ( .A(n20662), .ZN(n20675) );
  AOI21_X1 U22708 ( .B1(n19762), .B2(n19756), .A(n20675), .ZN(P1_U2802) );
  OAI21_X1 U22709 ( .B1(n19758), .B2(n19757), .A(P1_CODEFETCH_REG_SCAN_IN), 
        .ZN(n19759) );
  OAI21_X1 U22710 ( .B1(n19760), .B2(n15822), .A(n19759), .ZN(P1_U2803) );
  NOR2_X1 U22711 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(P1_STATE_REG_0__SCAN_IN), 
        .ZN(n19763) );
  OAI21_X1 U22712 ( .B1(n19763), .B2(P1_D_C_N_REG_SCAN_IN), .A(n20662), .ZN(
        n19761) );
  OAI21_X1 U22713 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(n20662), .A(n19761), 
        .ZN(P1_U2804) );
  NOR2_X1 U22714 ( .A1(n20675), .A2(n19762), .ZN(n20654) );
  OAI21_X1 U22715 ( .B1(BS16), .B2(n19763), .A(n20654), .ZN(n20652) );
  OAI21_X1 U22716 ( .B1(n20654), .B2(n20439), .A(n20652), .ZN(P1_U2805) );
  OAI21_X1 U22717 ( .B1(n19766), .B2(n19765), .A(n19764), .ZN(P1_U2806) );
  NOR4_X1 U22718 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_21__SCAN_IN), .A3(P1_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_23__SCAN_IN), .ZN(n19770) );
  NOR4_X1 U22719 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_17__SCAN_IN), .A3(P1_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_19__SCAN_IN), .ZN(n19769) );
  NOR4_X1 U22720 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_29__SCAN_IN), .A3(P1_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_31__SCAN_IN), .ZN(n19768) );
  NOR4_X1 U22721 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_25__SCAN_IN), .A3(P1_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_27__SCAN_IN), .ZN(n19767) );
  NAND4_X1 U22722 ( .A1(n19770), .A2(n19769), .A3(n19768), .A4(n19767), .ZN(
        n19776) );
  NOR4_X1 U22723 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_5__SCAN_IN), .A3(P1_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_7__SCAN_IN), .ZN(n19774) );
  AOI211_X1 U22724 ( .C1(P1_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A(P1_DATAWIDTH_REG_2__SCAN_IN), .B(
        P1_DATAWIDTH_REG_3__SCAN_IN), .ZN(n19773) );
  NOR4_X1 U22725 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_13__SCAN_IN), .A3(P1_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_15__SCAN_IN), .ZN(n19772) );
  NOR4_X1 U22726 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_9__SCAN_IN), .A3(P1_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_11__SCAN_IN), .ZN(n19771) );
  NAND4_X1 U22727 ( .A1(n19774), .A2(n19773), .A3(n19772), .A4(n19771), .ZN(
        n19775) );
  NOR2_X1 U22728 ( .A1(n19776), .A2(n19775), .ZN(n20659) );
  INV_X1 U22729 ( .A(n20659), .ZN(n19779) );
  NAND2_X1 U22730 ( .A1(n20659), .A2(n12475), .ZN(n20656) );
  NOR3_X1 U22731 ( .A1(P1_DATAWIDTH_REG_1__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A3(n20656), .ZN(n19778) );
  AOI21_X1 U22732 ( .B1(P1_BYTEENABLE_REG_1__SCAN_IN), .B2(n19779), .A(n19778), 
        .ZN(n19777) );
  OAI21_X1 U22733 ( .B1(n12917), .B2(n19779), .A(n19777), .ZN(P1_U2807) );
  NAND2_X1 U22734 ( .A1(n20659), .A2(n12917), .ZN(n20660) );
  AOI21_X1 U22735 ( .B1(P1_BYTEENABLE_REG_3__SCAN_IN), .B2(n19779), .A(n19778), 
        .ZN(n19780) );
  OAI21_X1 U22736 ( .B1(P1_DATAWIDTH_REG_1__SCAN_IN), .B2(n20660), .A(n19780), 
        .ZN(P1_U2808) );
  OAI21_X1 U22737 ( .B1(n19828), .B2(n19781), .A(n19826), .ZN(n19802) );
  NOR3_X1 U22738 ( .A1(n19838), .A2(P1_REIP_REG_9__SCAN_IN), .A3(n19781), .ZN(
        n19782) );
  AOI211_X1 U22739 ( .C1(n19861), .C2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .A(
        n13009), .B(n19782), .ZN(n19783) );
  OAI21_X1 U22740 ( .B1(n19836), .B2(n19784), .A(n19783), .ZN(n19785) );
  AOI21_X1 U22741 ( .B1(P1_EBX_REG_9__SCAN_IN), .B2(n19850), .A(n19785), .ZN(
        n19790) );
  INV_X1 U22742 ( .A(n19786), .ZN(n19788) );
  AOI22_X1 U22743 ( .A1(n19788), .A2(n19816), .B1(n19860), .B2(n19787), .ZN(
        n19789) );
  OAI211_X1 U22744 ( .C1(n19802), .C2(n20612), .A(n19790), .B(n19789), .ZN(
        P1_U2831) );
  AOI21_X1 U22745 ( .B1(n19857), .B2(n19791), .A(P1_REIP_REG_8__SCAN_IN), .ZN(
        n19801) );
  OAI22_X1 U22746 ( .A1(n19793), .A2(n19823), .B1(n19792), .B2(n19870), .ZN(
        n19794) );
  AOI211_X1 U22747 ( .C1(n19856), .C2(n19795), .A(n13009), .B(n19794), .ZN(
        n19800) );
  INV_X1 U22748 ( .A(n19796), .ZN(n19797) );
  AOI22_X1 U22749 ( .A1(n19798), .A2(n19816), .B1(n19797), .B2(n19860), .ZN(
        n19799) );
  OAI211_X1 U22750 ( .C1(n19802), .C2(n19801), .A(n19800), .B(n19799), .ZN(
        P1_U2832) );
  NOR3_X1 U22751 ( .A1(n19838), .A2(n19806), .A3(P1_REIP_REG_7__SCAN_IN), .ZN(
        n19805) );
  INV_X1 U22752 ( .A(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n19803) );
  OAI21_X1 U22753 ( .B1(n19823), .B2(n19803), .A(n19845), .ZN(n19804) );
  AOI211_X1 U22754 ( .C1(n19850), .C2(P1_EBX_REG_7__SCAN_IN), .A(n19805), .B(
        n19804), .ZN(n19811) );
  AOI21_X1 U22755 ( .B1(n19857), .B2(n19806), .A(n19828), .ZN(n19814) );
  OAI22_X1 U22756 ( .A1(n19814), .A2(n20609), .B1(n19807), .B2(n19829), .ZN(
        n19808) );
  AOI21_X1 U22757 ( .B1(n19809), .B2(n19816), .A(n19808), .ZN(n19810) );
  OAI211_X1 U22758 ( .C1(n19836), .C2(n19812), .A(n19811), .B(n19810), .ZN(
        P1_U2833) );
  AOI21_X1 U22759 ( .B1(n19861), .B2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n13009), .ZN(n19821) );
  AOI22_X1 U22760 ( .A1(P1_EBX_REG_6__SCAN_IN), .A2(n19850), .B1(n19856), .B2(
        n19871), .ZN(n19820) );
  INV_X1 U22761 ( .A(P1_REIP_REG_6__SCAN_IN), .ZN(n20730) );
  OAI22_X1 U22762 ( .A1(n19814), .A2(n20730), .B1(n19813), .B2(n19829), .ZN(
        n19815) );
  AOI21_X1 U22763 ( .B1(n19872), .B2(n19816), .A(n19815), .ZN(n19819) );
  NAND3_X1 U22764 ( .A1(n19857), .A2(n20730), .A3(n19817), .ZN(n19818) );
  NAND4_X1 U22765 ( .A1(n19821), .A2(n19820), .A3(n19819), .A4(n19818), .ZN(
        P1_U2834) );
  NOR3_X1 U22766 ( .A1(n19838), .A2(n19827), .A3(P1_REIP_REG_5__SCAN_IN), .ZN(
        n19825) );
  OAI21_X1 U22767 ( .B1(n19823), .B2(n19822), .A(n19845), .ZN(n19824) );
  AOI211_X1 U22768 ( .C1(n19850), .C2(P1_EBX_REG_5__SCAN_IN), .A(n19825), .B(
        n19824), .ZN(n19834) );
  OAI21_X1 U22769 ( .B1(n19828), .B2(n19827), .A(n19826), .ZN(n19854) );
  OAI22_X1 U22770 ( .A1(n19854), .A2(n20606), .B1(n19830), .B2(n19829), .ZN(
        n19831) );
  AOI21_X1 U22771 ( .B1(n19832), .B2(n19866), .A(n19831), .ZN(n19833) );
  OAI211_X1 U22772 ( .C1(n19836), .C2(n19835), .A(n19834), .B(n19833), .ZN(
        P1_U2835) );
  INV_X1 U22773 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n20604) );
  NAND3_X1 U22774 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_3__SCAN_IN), 
        .A3(P1_REIP_REG_2__SCAN_IN), .ZN(n19837) );
  NOR3_X1 U22775 ( .A1(n19838), .A2(P1_REIP_REG_4__SCAN_IN), .A3(n19837), .ZN(
        n19849) );
  AOI21_X1 U22776 ( .B1(n12761), .B2(n19841), .A(n19840), .ZN(n19844) );
  INV_X1 U22777 ( .A(n19842), .ZN(n19843) );
  NOR2_X1 U22778 ( .A1(n19844), .A2(n19843), .ZN(n19949) );
  AOI22_X1 U22779 ( .A1(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n19861), .B1(
        n19856), .B2(n19949), .ZN(n19846) );
  OAI211_X1 U22780 ( .C1(n19847), .C2(n19864), .A(n19846), .B(n19845), .ZN(
        n19848) );
  AOI211_X1 U22781 ( .C1(n19850), .C2(P1_EBX_REG_4__SCAN_IN), .A(n19849), .B(
        n19848), .ZN(n19853) );
  INV_X1 U22782 ( .A(n19947), .ZN(n19851) );
  AOI22_X1 U22783 ( .A1(n19943), .A2(n19866), .B1(n19851), .B2(n19860), .ZN(
        n19852) );
  OAI211_X1 U22784 ( .C1(n19854), .C2(n20604), .A(n19853), .B(n19852), .ZN(
        P1_U2836) );
  AOI22_X1 U22785 ( .A1(n19856), .A2(n19967), .B1(P1_REIP_REG_2__SCAN_IN), 
        .B2(n19855), .ZN(n19869) );
  INV_X1 U22786 ( .A(P1_REIP_REG_2__SCAN_IN), .ZN(n20600) );
  NAND3_X1 U22787 ( .A1(n19857), .A2(n20600), .A3(P1_REIP_REG_1__SCAN_IN), 
        .ZN(n19863) );
  INV_X1 U22788 ( .A(n19858), .ZN(n19859) );
  AOI22_X1 U22789 ( .A1(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n19861), .B1(
        n19860), .B2(n19859), .ZN(n19862) );
  OAI211_X1 U22790 ( .C1(n19864), .C2(n9754), .A(n19863), .B(n19862), .ZN(
        n19865) );
  AOI21_X1 U22791 ( .B1(n19867), .B2(n19866), .A(n19865), .ZN(n19868) );
  OAI211_X1 U22792 ( .C1(n20857), .C2(n19870), .A(n19869), .B(n19868), .ZN(
        P1_U2838) );
  AOI22_X1 U22793 ( .A1(n19872), .A2(n19876), .B1(n19875), .B2(n19871), .ZN(
        n19873) );
  OAI21_X1 U22794 ( .B1(n19879), .B2(n19874), .A(n19873), .ZN(P1_U2866) );
  AOI22_X1 U22795 ( .A1(n19943), .A2(n19876), .B1(n19875), .B2(n19949), .ZN(
        n19877) );
  OAI21_X1 U22796 ( .B1(n19879), .B2(n19878), .A(n19877), .ZN(P1_U2868) );
  AOI22_X1 U22797 ( .A1(P1_EAX_REG_15__SCAN_IN), .A2(n19885), .B1(n19903), 
        .B2(P1_DATAO_REG_15__SCAN_IN), .ZN(n19880) );
  OAI21_X1 U22798 ( .B1(n19881), .B2(n19887), .A(n19880), .ZN(P1_U2921) );
  INV_X1 U22799 ( .A(P1_LWORD_REG_14__SCAN_IN), .ZN(n20747) );
  AOI22_X1 U22800 ( .A1(P1_EAX_REG_14__SCAN_IN), .A2(n19885), .B1(n19903), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n19882) );
  OAI21_X1 U22801 ( .B1(n20747), .B2(n19887), .A(n19882), .ZN(P1_U2922) );
  INV_X1 U22802 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n19884) );
  AOI22_X1 U22803 ( .A1(P1_LWORD_REG_13__SCAN_IN), .A2(n20667), .B1(n19903), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n19883) );
  OAI21_X1 U22804 ( .B1(n19884), .B2(n19905), .A(n19883), .ZN(P1_U2923) );
  INV_X1 U22805 ( .A(P1_LWORD_REG_12__SCAN_IN), .ZN(n20833) );
  AOI22_X1 U22806 ( .A1(P1_EAX_REG_12__SCAN_IN), .A2(n19885), .B1(n19903), 
        .B2(P1_DATAO_REG_12__SCAN_IN), .ZN(n19886) );
  OAI21_X1 U22807 ( .B1(n20833), .B2(n19887), .A(n19886), .ZN(P1_U2924) );
  AOI22_X1 U22808 ( .A1(P1_LWORD_REG_11__SCAN_IN), .A2(n20667), .B1(n19903), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n19888) );
  OAI21_X1 U22809 ( .B1(n13543), .B2(n19905), .A(n19888), .ZN(P1_U2925) );
  INV_X1 U22810 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n19890) );
  AOI22_X1 U22811 ( .A1(P1_LWORD_REG_10__SCAN_IN), .A2(n20667), .B1(n19903), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n19889) );
  OAI21_X1 U22812 ( .B1(n19890), .B2(n19905), .A(n19889), .ZN(P1_U2926) );
  INV_X1 U22813 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n19892) );
  AOI22_X1 U22814 ( .A1(P1_LWORD_REG_9__SCAN_IN), .A2(n20667), .B1(n19903), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n19891) );
  OAI21_X1 U22815 ( .B1(n19892), .B2(n19905), .A(n19891), .ZN(P1_U2927) );
  AOI22_X1 U22816 ( .A1(P1_LWORD_REG_8__SCAN_IN), .A2(n20667), .B1(n19903), 
        .B2(P1_DATAO_REG_8__SCAN_IN), .ZN(n19893) );
  OAI21_X1 U22817 ( .B1(n13138), .B2(n19905), .A(n19893), .ZN(P1_U2928) );
  AOI22_X1 U22818 ( .A1(P1_LWORD_REG_7__SCAN_IN), .A2(n20667), .B1(n19903), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n19894) );
  OAI21_X1 U22819 ( .B1(n13093), .B2(n19905), .A(n19894), .ZN(P1_U2929) );
  AOI22_X1 U22820 ( .A1(P1_LWORD_REG_6__SCAN_IN), .A2(n20667), .B1(n19903), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n19895) );
  OAI21_X1 U22821 ( .B1(n19896), .B2(n19905), .A(n19895), .ZN(P1_U2930) );
  AOI22_X1 U22822 ( .A1(P1_LWORD_REG_5__SCAN_IN), .A2(n20667), .B1(n19903), 
        .B2(P1_DATAO_REG_5__SCAN_IN), .ZN(n19897) );
  OAI21_X1 U22823 ( .B1(n12740), .B2(n19905), .A(n19897), .ZN(P1_U2931) );
  AOI22_X1 U22824 ( .A1(P1_LWORD_REG_4__SCAN_IN), .A2(n20667), .B1(n19903), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n19898) );
  OAI21_X1 U22825 ( .B1(n19899), .B2(n19905), .A(n19898), .ZN(P1_U2932) );
  AOI22_X1 U22826 ( .A1(P1_LWORD_REG_3__SCAN_IN), .A2(n20667), .B1(n19903), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n19900) );
  OAI21_X1 U22827 ( .B1(n12675), .B2(n19905), .A(n19900), .ZN(P1_U2933) );
  AOI22_X1 U22828 ( .A1(P1_LWORD_REG_2__SCAN_IN), .A2(n20667), .B1(n19903), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n19901) );
  OAI21_X1 U22829 ( .B1(n12643), .B2(n19905), .A(n19901), .ZN(P1_U2934) );
  AOI22_X1 U22830 ( .A1(P1_LWORD_REG_1__SCAN_IN), .A2(n20667), .B1(n19903), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n19902) );
  OAI21_X1 U22831 ( .B1(n12440), .B2(n19905), .A(n19902), .ZN(P1_U2935) );
  AOI22_X1 U22832 ( .A1(P1_LWORD_REG_0__SCAN_IN), .A2(n20667), .B1(n19903), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n19904) );
  OAI21_X1 U22833 ( .B1(n19906), .B2(n19905), .A(n19904), .ZN(P1_U2936) );
  AOI22_X1 U22834 ( .A1(n19909), .A2(P1_EAX_REG_24__SCAN_IN), .B1(
        P1_UWORD_REG_8__SCAN_IN), .B2(n19912), .ZN(n19908) );
  NAND2_X1 U22835 ( .A1(n19920), .A2(n19907), .ZN(n19922) );
  NAND2_X1 U22836 ( .A1(n19908), .A2(n19922), .ZN(P1_U2945) );
  AOI22_X1 U22837 ( .A1(n19909), .A2(P1_EAX_REG_25__SCAN_IN), .B1(
        P1_UWORD_REG_9__SCAN_IN), .B2(n19912), .ZN(n19911) );
  NAND2_X1 U22838 ( .A1(n19920), .A2(n19910), .ZN(n19924) );
  NAND2_X1 U22839 ( .A1(n19911), .A2(n19924), .ZN(P1_U2946) );
  AOI22_X1 U22840 ( .A1(n19935), .A2(P1_EAX_REG_27__SCAN_IN), .B1(
        P1_UWORD_REG_11__SCAN_IN), .B2(n19912), .ZN(n19914) );
  NAND2_X1 U22841 ( .A1(n19920), .A2(n19913), .ZN(n19928) );
  NAND2_X1 U22842 ( .A1(n19914), .A2(n19928), .ZN(P1_U2948) );
  AOI22_X1 U22843 ( .A1(n19935), .A2(P1_EAX_REG_28__SCAN_IN), .B1(
        P1_UWORD_REG_12__SCAN_IN), .B2(n19932), .ZN(n19916) );
  NAND2_X1 U22844 ( .A1(n19920), .A2(n19915), .ZN(n19930) );
  NAND2_X1 U22845 ( .A1(n19916), .A2(n19930), .ZN(P1_U2949) );
  AOI22_X1 U22846 ( .A1(n19935), .A2(P1_EAX_REG_29__SCAN_IN), .B1(
        P1_UWORD_REG_13__SCAN_IN), .B2(n19932), .ZN(n19918) );
  NAND2_X1 U22847 ( .A1(n19920), .A2(n19917), .ZN(n19933) );
  NAND2_X1 U22848 ( .A1(n19918), .A2(n19933), .ZN(P1_U2950) );
  AOI22_X1 U22849 ( .A1(n19935), .A2(P1_EAX_REG_30__SCAN_IN), .B1(
        P1_UWORD_REG_14__SCAN_IN), .B2(n19932), .ZN(n19921) );
  NAND2_X1 U22850 ( .A1(n19920), .A2(n19919), .ZN(n19936) );
  NAND2_X1 U22851 ( .A1(n19921), .A2(n19936), .ZN(P1_U2951) );
  AOI22_X1 U22852 ( .A1(n19935), .A2(P1_EAX_REG_8__SCAN_IN), .B1(
        P1_LWORD_REG_8__SCAN_IN), .B2(n19932), .ZN(n19923) );
  NAND2_X1 U22853 ( .A1(n19923), .A2(n19922), .ZN(P1_U2960) );
  AOI22_X1 U22854 ( .A1(n19935), .A2(P1_EAX_REG_9__SCAN_IN), .B1(
        P1_LWORD_REG_9__SCAN_IN), .B2(n19932), .ZN(n19925) );
  NAND2_X1 U22855 ( .A1(n19925), .A2(n19924), .ZN(P1_U2961) );
  AOI22_X1 U22856 ( .A1(n19935), .A2(P1_EAX_REG_10__SCAN_IN), .B1(
        P1_LWORD_REG_10__SCAN_IN), .B2(n19932), .ZN(n19927) );
  NAND2_X1 U22857 ( .A1(n19927), .A2(n19926), .ZN(P1_U2962) );
  AOI22_X1 U22858 ( .A1(n19935), .A2(P1_EAX_REG_11__SCAN_IN), .B1(
        P1_LWORD_REG_11__SCAN_IN), .B2(n19932), .ZN(n19929) );
  NAND2_X1 U22859 ( .A1(n19929), .A2(n19928), .ZN(P1_U2963) );
  AOI22_X1 U22860 ( .A1(n19935), .A2(P1_EAX_REG_12__SCAN_IN), .B1(
        P1_LWORD_REG_12__SCAN_IN), .B2(n19932), .ZN(n19931) );
  NAND2_X1 U22861 ( .A1(n19931), .A2(n19930), .ZN(P1_U2964) );
  AOI22_X1 U22862 ( .A1(n19935), .A2(P1_EAX_REG_13__SCAN_IN), .B1(
        P1_LWORD_REG_13__SCAN_IN), .B2(n19932), .ZN(n19934) );
  NAND2_X1 U22863 ( .A1(n19934), .A2(n19933), .ZN(P1_U2965) );
  AOI22_X1 U22864 ( .A1(n19935), .A2(P1_EAX_REG_14__SCAN_IN), .B1(
        P1_LWORD_REG_14__SCAN_IN), .B2(n19932), .ZN(n19937) );
  NAND2_X1 U22865 ( .A1(n19937), .A2(n19936), .ZN(P1_U2966) );
  AOI22_X1 U22866 ( .A1(n19938), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B1(
        n13009), .B2(P1_REIP_REG_4__SCAN_IN), .ZN(n19946) );
  OAI21_X1 U22867 ( .B1(n19941), .B2(n19940), .A(n19939), .ZN(n19942) );
  INV_X1 U22868 ( .A(n19942), .ZN(n19950) );
  AOI22_X1 U22869 ( .A1(n19950), .A2(n19944), .B1(n9727), .B2(n19943), .ZN(
        n19945) );
  OAI211_X1 U22870 ( .C1(n15701), .C2(n19947), .A(n19946), .B(n19945), .ZN(
        P1_U2995) );
  OAI21_X1 U22871 ( .B1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A(n19948), .ZN(n19953) );
  AOI22_X1 U22872 ( .A1(n13009), .A2(P1_REIP_REG_4__SCAN_IN), .B1(n19993), 
        .B2(n19949), .ZN(n19952) );
  AOI22_X1 U22873 ( .A1(n19950), .A2(n19994), .B1(
        P1_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n19956), .ZN(n19951) );
  OAI211_X1 U22874 ( .C1(n19960), .C2(n19953), .A(n19952), .B(n19951), .ZN(
        P1_U3027) );
  AOI22_X1 U22875 ( .A1(n13009), .A2(P1_REIP_REG_3__SCAN_IN), .B1(n19993), 
        .B2(n19954), .ZN(n19959) );
  INV_X1 U22876 ( .A(n19955), .ZN(n19957) );
  AOI22_X1 U22877 ( .A1(n19957), .A2(n19994), .B1(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n19956), .ZN(n19958) );
  OAI211_X1 U22878 ( .C1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .C2(n19960), .A(
        n19959), .B(n19958), .ZN(P1_U3028) );
  NAND2_X1 U22879 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n19961), .ZN(
        n19980) );
  AOI21_X1 U22880 ( .B1(n12449), .B2(n19963), .A(n19962), .ZN(n19979) );
  NOR2_X1 U22881 ( .A1(n19965), .A2(n19964), .ZN(n19977) );
  NAND2_X1 U22882 ( .A1(n13009), .A2(P1_REIP_REG_2__SCAN_IN), .ZN(n19974) );
  NAND2_X1 U22883 ( .A1(n19993), .A2(n19967), .ZN(n19973) );
  NOR2_X1 U22884 ( .A1(n19969), .A2(n19968), .ZN(n19970) );
  NAND2_X1 U22885 ( .A1(n19971), .A2(n19970), .ZN(n19972) );
  NAND4_X1 U22886 ( .A1(n19975), .A2(n19974), .A3(n19973), .A4(n19972), .ZN(
        n19976) );
  AOI21_X1 U22887 ( .B1(n19977), .B2(n13236), .A(n19976), .ZN(n19978) );
  OAI221_X1 U22888 ( .B1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n19980), .C1(
        n20722), .C2(n19979), .A(n19978), .ZN(P1_U3029) );
  INV_X1 U22889 ( .A(n19981), .ZN(n19983) );
  AOI21_X1 U22890 ( .B1(n19993), .B2(n19983), .A(n19982), .ZN(n19991) );
  OAI21_X1 U22891 ( .B1(n19985), .B2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n19984), .ZN(n19997) );
  AOI22_X1 U22892 ( .A1(n19986), .A2(n19994), .B1(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n19997), .ZN(n19990) );
  NAND3_X1 U22893 ( .A1(n12449), .A2(n19988), .A3(n19987), .ZN(n19989) );
  NAND3_X1 U22894 ( .A1(n19991), .A2(n19990), .A3(n19989), .ZN(P1_U3030) );
  AOI22_X1 U22895 ( .A1(n19995), .A2(n19994), .B1(n19993), .B2(n19992), .ZN(
        n20001) );
  OAI22_X1 U22896 ( .A1(n19998), .A2(n19997), .B1(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n19996), .ZN(n19999) );
  NAND3_X1 U22897 ( .A1(n20001), .A2(n20000), .A3(n19999), .ZN(P1_U3031) );
  NOR2_X1 U22898 ( .A1(n20003), .A2(n20002), .ZN(P1_U3032) );
  NOR2_X2 U22899 ( .A1(n20005), .A2(n20004), .ZN(n20046) );
  AOI22_X1 U22900 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n20046), .B1(DATAI_16_), 
        .B2(n20007), .ZN(n20478) );
  AOI22_X1 U22901 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n20046), .B1(DATAI_24_), 
        .B2(n20007), .ZN(n20529) );
  INV_X1 U22902 ( .A(n20529), .ZN(n20475) );
  NOR2_X2 U22903 ( .A1(n20048), .A2(n20010), .ZN(n20515) );
  NAND3_X1 U22904 ( .A1(n20368), .A2(n20321), .A3(n20757), .ZN(n20056) );
  NOR2_X1 U22905 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20056), .ZN(
        n20049) );
  AOI22_X1 U22906 ( .A1(n20571), .A2(n20475), .B1(n20515), .B2(n20049), .ZN(
        n20022) );
  INV_X1 U22907 ( .A(n20018), .ZN(n20011) );
  NOR2_X1 U22908 ( .A1(n20011), .A2(n12396), .ZN(n20155) );
  NOR3_X1 U22909 ( .A1(n20079), .A2(n20571), .A3(n20518), .ZN(n20012) );
  NAND2_X1 U22910 ( .A1(n20524), .A2(n20439), .ZN(n20403) );
  INV_X1 U22911 ( .A(n20403), .ZN(n20186) );
  NOR2_X1 U22912 ( .A1(n20012), .A2(n20186), .ZN(n20020) );
  INV_X1 U22913 ( .A(n20020), .ZN(n20015) );
  INV_X1 U22914 ( .A(n9754), .ZN(n20013) );
  NAND2_X1 U22915 ( .A1(n9821), .A2(n20406), .ZN(n20019) );
  INV_X1 U22916 ( .A(n20270), .ZN(n20014) );
  NAND2_X1 U22917 ( .A1(n20014), .A2(n20326), .ZN(n20158) );
  AOI22_X1 U22918 ( .A1(n20015), .A2(n20019), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n20158), .ZN(n20016) );
  OAI211_X1 U22919 ( .C1(n20049), .C2(n20275), .A(n20328), .B(n20016), .ZN(
        n20052) );
  NOR2_X2 U22920 ( .A1(n20017), .A2(n20057), .ZN(n20516) );
  OR2_X1 U22921 ( .A1(n20018), .A2(n12396), .ZN(n20330) );
  OAI22_X1 U22922 ( .A1(n20020), .A2(n20019), .B1(n20330), .B2(n20158), .ZN(
        n20051) );
  AOI22_X1 U22923 ( .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n20052), .B1(
        n20516), .B2(n20051), .ZN(n20021) );
  OAI211_X1 U22924 ( .C1(n20478), .C2(n20076), .A(n20022), .B(n20021), .ZN(
        P1_U3033) );
  AOI22_X1 U22925 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n20046), .B1(DATAI_25_), 
        .B2(n20007), .ZN(n20535) );
  INV_X1 U22926 ( .A(n20535), .ZN(n20479) );
  NOR2_X2 U22927 ( .A1(n20048), .A2(n12180), .ZN(n20530) );
  AOI22_X1 U22928 ( .A1(n20571), .A2(n20479), .B1(n20530), .B2(n20049), .ZN(
        n20025) );
  NOR2_X2 U22929 ( .A1(n20023), .A2(n20057), .ZN(n20531) );
  AOI22_X1 U22930 ( .A1(P1_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n20052), .B1(
        n20531), .B2(n20051), .ZN(n20024) );
  OAI211_X1 U22931 ( .C1(n20482), .C2(n20076), .A(n20025), .B(n20024), .ZN(
        P1_U3034) );
  AOI22_X1 U22932 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n20046), .B1(DATAI_26_), 
        .B2(n20007), .ZN(n20541) );
  INV_X1 U22933 ( .A(n20541), .ZN(n20483) );
  NOR2_X2 U22934 ( .A1(n20048), .A2(n20026), .ZN(n20536) );
  AOI22_X1 U22935 ( .A1(n20571), .A2(n20483), .B1(n20536), .B2(n20049), .ZN(
        n20029) );
  NOR2_X2 U22936 ( .A1(n20027), .A2(n20057), .ZN(n20537) );
  AOI22_X1 U22937 ( .A1(P1_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n20052), .B1(
        n20537), .B2(n20051), .ZN(n20028) );
  OAI211_X1 U22938 ( .C1(n20486), .C2(n20076), .A(n20029), .B(n20028), .ZN(
        P1_U3035) );
  AOI22_X1 U22939 ( .A1(DATAI_19_), .A2(n20007), .B1(BUF1_REG_19__SCAN_IN), 
        .B2(n20046), .ZN(n20490) );
  AOI22_X1 U22940 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n20046), .B1(DATAI_27_), 
        .B2(n20007), .ZN(n20547) );
  INV_X1 U22941 ( .A(n20547), .ZN(n20487) );
  NOR2_X2 U22942 ( .A1(n20048), .A2(n20030), .ZN(n20542) );
  AOI22_X1 U22943 ( .A1(n20571), .A2(n20487), .B1(n20542), .B2(n20049), .ZN(
        n20033) );
  NOR2_X2 U22944 ( .A1(n20031), .A2(n20057), .ZN(n20543) );
  AOI22_X1 U22945 ( .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n20052), .B1(
        n20543), .B2(n20051), .ZN(n20032) );
  OAI211_X1 U22946 ( .C1(n20490), .C2(n20076), .A(n20033), .B(n20032), .ZN(
        P1_U3036) );
  AOI22_X1 U22947 ( .A1(DATAI_20_), .A2(n20007), .B1(BUF1_REG_20__SCAN_IN), 
        .B2(n20046), .ZN(n20494) );
  INV_X1 U22948 ( .A(n20553), .ZN(n20491) );
  NOR2_X2 U22949 ( .A1(n20048), .A2(n20034), .ZN(n20548) );
  AOI22_X1 U22950 ( .A1(n20571), .A2(n20491), .B1(n20548), .B2(n20049), .ZN(
        n20037) );
  NOR2_X2 U22951 ( .A1(n20035), .A2(n20057), .ZN(n20549) );
  AOI22_X1 U22952 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n20052), .B1(
        n20549), .B2(n20051), .ZN(n20036) );
  OAI211_X1 U22953 ( .C1(n20494), .C2(n20076), .A(n20037), .B(n20036), .ZN(
        P1_U3037) );
  AOI22_X1 U22954 ( .A1(DATAI_21_), .A2(n20007), .B1(BUF1_REG_21__SCAN_IN), 
        .B2(n20046), .ZN(n20498) );
  AOI22_X1 U22955 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n20046), .B1(DATAI_29_), 
        .B2(n20007), .ZN(n20559) );
  INV_X1 U22956 ( .A(n20559), .ZN(n20495) );
  NOR2_X2 U22957 ( .A1(n20048), .A2(n20038), .ZN(n20554) );
  AOI22_X1 U22958 ( .A1(n20571), .A2(n20495), .B1(n20554), .B2(n20049), .ZN(
        n20041) );
  NOR2_X2 U22959 ( .A1(n20039), .A2(n20057), .ZN(n20555) );
  AOI22_X1 U22960 ( .A1(P1_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n20052), .B1(
        n20555), .B2(n20051), .ZN(n20040) );
  OAI211_X1 U22961 ( .C1(n20498), .C2(n20076), .A(n20041), .B(n20040), .ZN(
        P1_U3038) );
  AOI22_X1 U22962 ( .A1(DATAI_22_), .A2(n20007), .B1(BUF1_REG_22__SCAN_IN), 
        .B2(n20046), .ZN(n20502) );
  AOI22_X1 U22963 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n20046), .B1(DATAI_30_), 
        .B2(n20007), .ZN(n20565) );
  INV_X1 U22964 ( .A(n20565), .ZN(n20499) );
  NOR2_X2 U22965 ( .A1(n20048), .A2(n20042), .ZN(n20560) );
  AOI22_X1 U22966 ( .A1(n20571), .A2(n20499), .B1(n20560), .B2(n20049), .ZN(
        n20045) );
  NOR2_X2 U22967 ( .A1(n20043), .A2(n20057), .ZN(n20561) );
  AOI22_X1 U22968 ( .A1(P1_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n20052), .B1(
        n20561), .B2(n20051), .ZN(n20044) );
  OAI211_X1 U22969 ( .C1(n20502), .C2(n20076), .A(n20045), .B(n20044), .ZN(
        P1_U3039) );
  AOI22_X1 U22970 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n20046), .B1(DATAI_23_), 
        .B2(n20007), .ZN(n20510) );
  AOI22_X1 U22971 ( .A1(DATAI_31_), .A2(n20007), .B1(BUF1_REG_31__SCAN_IN), 
        .B2(n20046), .ZN(n20576) );
  INV_X1 U22972 ( .A(n20576), .ZN(n20505) );
  NOR2_X2 U22973 ( .A1(n20048), .A2(n20047), .ZN(n20567) );
  AOI22_X1 U22974 ( .A1(n20571), .A2(n20505), .B1(n20567), .B2(n20049), .ZN(
        n20054) );
  NOR2_X2 U22975 ( .A1(n20050), .A2(n20057), .ZN(n20569) );
  AOI22_X1 U22976 ( .A1(P1_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n20052), .B1(
        n20569), .B2(n20051), .ZN(n20053) );
  OAI211_X1 U22977 ( .C1(n20510), .C2(n20076), .A(n20054), .B(n20053), .ZN(
        P1_U3040) );
  INV_X1 U22978 ( .A(n20055), .ZN(n20436) );
  NOR2_X1 U22979 ( .A1(n20435), .A2(n20056), .ZN(n20077) );
  AOI21_X1 U22980 ( .B1(n9821), .B2(n20436), .A(n20077), .ZN(n20058) );
  OAI22_X1 U22981 ( .A1(n20058), .A2(n20518), .B1(n20056), .B2(n12396), .ZN(
        n20078) );
  AOI22_X1 U22982 ( .A1(n20516), .A2(n20078), .B1(n20515), .B2(n20077), .ZN(
        n20062) );
  INV_X1 U22983 ( .A(n20056), .ZN(n20060) );
  OAI211_X1 U22984 ( .C1(n20122), .C2(n20439), .A(n20524), .B(n20058), .ZN(
        n20059) );
  OAI211_X1 U22985 ( .C1(n20524), .C2(n20060), .A(n20523), .B(n20059), .ZN(
        n20080) );
  INV_X1 U22986 ( .A(n20117), .ZN(n20073) );
  INV_X1 U22987 ( .A(n20478), .ZN(n20526) );
  AOI22_X1 U22988 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n20080), .B1(
        n20073), .B2(n20526), .ZN(n20061) );
  OAI211_X1 U22989 ( .C1(n20529), .C2(n20076), .A(n20062), .B(n20061), .ZN(
        P1_U3041) );
  AOI22_X1 U22990 ( .A1(n20531), .A2(n20078), .B1(n20530), .B2(n20077), .ZN(
        n20064) );
  AOI22_X1 U22991 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n20080), .B1(
        n20079), .B2(n20479), .ZN(n20063) );
  OAI211_X1 U22992 ( .C1(n20482), .C2(n20117), .A(n20064), .B(n20063), .ZN(
        P1_U3042) );
  AOI22_X1 U22993 ( .A1(n20537), .A2(n20078), .B1(n20536), .B2(n20077), .ZN(
        n20066) );
  AOI22_X1 U22994 ( .A1(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n20080), .B1(
        n20079), .B2(n20483), .ZN(n20065) );
  OAI211_X1 U22995 ( .C1(n20486), .C2(n20117), .A(n20066), .B(n20065), .ZN(
        P1_U3043) );
  AOI22_X1 U22996 ( .A1(n20543), .A2(n20078), .B1(n20542), .B2(n20077), .ZN(
        n20068) );
  AOI22_X1 U22997 ( .A1(P1_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n20080), .B1(
        n20079), .B2(n20487), .ZN(n20067) );
  OAI211_X1 U22998 ( .C1(n20490), .C2(n20117), .A(n20068), .B(n20067), .ZN(
        P1_U3044) );
  AOI22_X1 U22999 ( .A1(n20549), .A2(n20078), .B1(n20548), .B2(n20077), .ZN(
        n20070) );
  INV_X1 U23000 ( .A(n20494), .ZN(n20550) );
  AOI22_X1 U23001 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n20080), .B1(
        n20073), .B2(n20550), .ZN(n20069) );
  OAI211_X1 U23002 ( .C1(n20553), .C2(n20076), .A(n20070), .B(n20069), .ZN(
        P1_U3045) );
  AOI22_X1 U23003 ( .A1(n20555), .A2(n20078), .B1(n20554), .B2(n20077), .ZN(
        n20072) );
  AOI22_X1 U23004 ( .A1(P1_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n20080), .B1(
        n20079), .B2(n20495), .ZN(n20071) );
  OAI211_X1 U23005 ( .C1(n20498), .C2(n20117), .A(n20072), .B(n20071), .ZN(
        P1_U3046) );
  AOI22_X1 U23006 ( .A1(n20561), .A2(n20078), .B1(n20560), .B2(n20077), .ZN(
        n20075) );
  INV_X1 U23007 ( .A(n20502), .ZN(n20562) );
  AOI22_X1 U23008 ( .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n20080), .B1(
        n20073), .B2(n20562), .ZN(n20074) );
  OAI211_X1 U23009 ( .C1(n20565), .C2(n20076), .A(n20075), .B(n20074), .ZN(
        P1_U3047) );
  AOI22_X1 U23010 ( .A1(n20569), .A2(n20078), .B1(n20567), .B2(n20077), .ZN(
        n20082) );
  AOI22_X1 U23011 ( .A1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n20080), .B1(
        n20079), .B2(n20505), .ZN(n20081) );
  OAI211_X1 U23012 ( .C1(n20510), .C2(n20117), .A(n20082), .B(n20081), .ZN(
        P1_U3048) );
  NAND2_X1 U23013 ( .A1(n9751), .A2(n20083), .ZN(n20463) );
  INV_X1 U23014 ( .A(n20515), .ZN(n20322) );
  NAND3_X1 U23015 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20368), .A3(
        n20321), .ZN(n20125) );
  OR2_X1 U23016 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20125), .ZN(
        n20111) );
  OAI22_X1 U23017 ( .A1(n20117), .A2(n20529), .B1(n20322), .B2(n20111), .ZN(
        n20084) );
  INV_X1 U23018 ( .A(n20084), .ZN(n20092) );
  NAND2_X1 U23019 ( .A1(n20149), .A2(n20117), .ZN(n20085) );
  AOI21_X1 U23020 ( .B1(n20085), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n20518), 
        .ZN(n20087) );
  NAND2_X1 U23021 ( .A1(n9821), .A2(n20465), .ZN(n20089) );
  AOI22_X1 U23022 ( .A1(n20087), .A2(n20089), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20111), .ZN(n20086) );
  OAI21_X1 U23023 ( .B1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n20326), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n20212) );
  NAND3_X1 U23024 ( .A1(n20328), .A2(n20086), .A3(n20212), .ZN(n20114) );
  INV_X1 U23025 ( .A(n20087), .ZN(n20090) );
  INV_X1 U23026 ( .A(n20326), .ZN(n20088) );
  NAND2_X1 U23027 ( .A1(n20088), .A2(n20368), .ZN(n20215) );
  OAI22_X1 U23028 ( .A1(n20090), .A2(n20089), .B1(n20330), .B2(n20215), .ZN(
        n20113) );
  AOI22_X1 U23029 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n20114), .B1(
        n20516), .B2(n20113), .ZN(n20091) );
  OAI211_X1 U23030 ( .C1(n20478), .C2(n20149), .A(n20092), .B(n20091), .ZN(
        P1_U3049) );
  INV_X1 U23031 ( .A(n20530), .ZN(n20335) );
  OAI22_X1 U23032 ( .A1(n20117), .A2(n20535), .B1(n20335), .B2(n20111), .ZN(
        n20093) );
  INV_X1 U23033 ( .A(n20093), .ZN(n20095) );
  AOI22_X1 U23034 ( .A1(P1_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n20114), .B1(
        n20531), .B2(n20113), .ZN(n20094) );
  OAI211_X1 U23035 ( .C1(n20482), .C2(n20149), .A(n20095), .B(n20094), .ZN(
        P1_U3050) );
  INV_X1 U23036 ( .A(n20536), .ZN(n20339) );
  OAI22_X1 U23037 ( .A1(n20117), .A2(n20541), .B1(n20339), .B2(n20111), .ZN(
        n20096) );
  INV_X1 U23038 ( .A(n20096), .ZN(n20098) );
  AOI22_X1 U23039 ( .A1(P1_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n20114), .B1(
        n20537), .B2(n20113), .ZN(n20097) );
  OAI211_X1 U23040 ( .C1(n20486), .C2(n20149), .A(n20098), .B(n20097), .ZN(
        P1_U3051) );
  INV_X1 U23041 ( .A(n20542), .ZN(n20343) );
  OAI22_X1 U23042 ( .A1(n20117), .A2(n20547), .B1(n20343), .B2(n20111), .ZN(
        n20099) );
  INV_X1 U23043 ( .A(n20099), .ZN(n20101) );
  AOI22_X1 U23044 ( .A1(P1_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n20114), .B1(
        n20543), .B2(n20113), .ZN(n20100) );
  OAI211_X1 U23045 ( .C1(n20490), .C2(n20149), .A(n20101), .B(n20100), .ZN(
        P1_U3052) );
  INV_X1 U23046 ( .A(n20548), .ZN(n20347) );
  OAI22_X1 U23047 ( .A1(n20149), .A2(n20494), .B1(n20347), .B2(n20111), .ZN(
        n20102) );
  INV_X1 U23048 ( .A(n20102), .ZN(n20104) );
  AOI22_X1 U23049 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n20114), .B1(
        n20549), .B2(n20113), .ZN(n20103) );
  OAI211_X1 U23050 ( .C1(n20553), .C2(n20117), .A(n20104), .B(n20103), .ZN(
        P1_U3053) );
  INV_X1 U23051 ( .A(n20554), .ZN(n20351) );
  OAI22_X1 U23052 ( .A1(n20149), .A2(n20498), .B1(n20351), .B2(n20111), .ZN(
        n20105) );
  INV_X1 U23053 ( .A(n20105), .ZN(n20107) );
  AOI22_X1 U23054 ( .A1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n20114), .B1(
        n20555), .B2(n20113), .ZN(n20106) );
  OAI211_X1 U23055 ( .C1(n20559), .C2(n20117), .A(n20107), .B(n20106), .ZN(
        P1_U3054) );
  INV_X1 U23056 ( .A(n20560), .ZN(n20355) );
  OAI22_X1 U23057 ( .A1(n20149), .A2(n20502), .B1(n20355), .B2(n20111), .ZN(
        n20108) );
  INV_X1 U23058 ( .A(n20108), .ZN(n20110) );
  AOI22_X1 U23059 ( .A1(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n20114), .B1(
        n20561), .B2(n20113), .ZN(n20109) );
  OAI211_X1 U23060 ( .C1(n20565), .C2(n20117), .A(n20110), .B(n20109), .ZN(
        P1_U3055) );
  INV_X1 U23061 ( .A(n20567), .ZN(n20360) );
  OAI22_X1 U23062 ( .A1(n20149), .A2(n20510), .B1(n20360), .B2(n20111), .ZN(
        n20112) );
  INV_X1 U23063 ( .A(n20112), .ZN(n20116) );
  AOI22_X1 U23064 ( .A1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n20114), .B1(
        n20569), .B2(n20113), .ZN(n20115) );
  OAI211_X1 U23065 ( .C1(n20576), .C2(n20117), .A(n20116), .B(n20115), .ZN(
        P1_U3056) );
  NOR2_X1 U23066 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n20367), .ZN(
        n20120) );
  INV_X1 U23067 ( .A(n20120), .ZN(n20148) );
  OAI22_X1 U23068 ( .A1(n20149), .A2(n20529), .B1(n20322), .B2(n20148), .ZN(
        n20118) );
  INV_X1 U23069 ( .A(n20118), .ZN(n20129) );
  AND2_X1 U23070 ( .A1(n12394), .A2(n20119), .ZN(n20512) );
  AOI21_X1 U23071 ( .B1(n9821), .B2(n20512), .A(n20120), .ZN(n20126) );
  INV_X1 U23072 ( .A(n20517), .ZN(n20121) );
  AOI21_X1 U23073 ( .B1(n20122), .B2(n20524), .A(n20121), .ZN(n20127) );
  INV_X1 U23074 ( .A(n20127), .ZN(n20123) );
  AOI22_X1 U23075 ( .A1(n20126), .A2(n20123), .B1(n20518), .B2(n20125), .ZN(
        n20124) );
  NAND2_X1 U23076 ( .A1(n20523), .A2(n20124), .ZN(n20152) );
  OAI22_X1 U23077 ( .A1(n20127), .A2(n20126), .B1(n12396), .B2(n20125), .ZN(
        n20151) );
  AOI22_X1 U23078 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n20152), .B1(
        n20516), .B2(n20151), .ZN(n20128) );
  OAI211_X1 U23079 ( .C1(n20478), .C2(n20183), .A(n20129), .B(n20128), .ZN(
        P1_U3057) );
  OAI22_X1 U23080 ( .A1(n20149), .A2(n20535), .B1(n20335), .B2(n20148), .ZN(
        n20130) );
  INV_X1 U23081 ( .A(n20130), .ZN(n20132) );
  AOI22_X1 U23082 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n20152), .B1(
        n20531), .B2(n20151), .ZN(n20131) );
  OAI211_X1 U23083 ( .C1(n20482), .C2(n20183), .A(n20132), .B(n20131), .ZN(
        P1_U3058) );
  OAI22_X1 U23084 ( .A1(n20183), .A2(n20486), .B1(n20339), .B2(n20148), .ZN(
        n20133) );
  INV_X1 U23085 ( .A(n20133), .ZN(n20135) );
  AOI22_X1 U23086 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n20152), .B1(
        n20537), .B2(n20151), .ZN(n20134) );
  OAI211_X1 U23087 ( .C1(n20541), .C2(n20149), .A(n20135), .B(n20134), .ZN(
        P1_U3059) );
  OAI22_X1 U23088 ( .A1(n20149), .A2(n20547), .B1(n20343), .B2(n20148), .ZN(
        n20136) );
  INV_X1 U23089 ( .A(n20136), .ZN(n20138) );
  AOI22_X1 U23090 ( .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20152), .B1(
        n20543), .B2(n20151), .ZN(n20137) );
  OAI211_X1 U23091 ( .C1(n20490), .C2(n20183), .A(n20138), .B(n20137), .ZN(
        P1_U3060) );
  OAI22_X1 U23092 ( .A1(n20149), .A2(n20553), .B1(n20347), .B2(n20148), .ZN(
        n20139) );
  INV_X1 U23093 ( .A(n20139), .ZN(n20141) );
  AOI22_X1 U23094 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n20152), .B1(
        n20549), .B2(n20151), .ZN(n20140) );
  OAI211_X1 U23095 ( .C1(n20494), .C2(n20183), .A(n20141), .B(n20140), .ZN(
        P1_U3061) );
  OAI22_X1 U23096 ( .A1(n20149), .A2(n20559), .B1(n20351), .B2(n20148), .ZN(
        n20142) );
  INV_X1 U23097 ( .A(n20142), .ZN(n20144) );
  AOI22_X1 U23098 ( .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n20152), .B1(
        n20555), .B2(n20151), .ZN(n20143) );
  OAI211_X1 U23099 ( .C1(n20498), .C2(n20183), .A(n20144), .B(n20143), .ZN(
        P1_U3062) );
  OAI22_X1 U23100 ( .A1(n20183), .A2(n20502), .B1(n20355), .B2(n20148), .ZN(
        n20145) );
  INV_X1 U23101 ( .A(n20145), .ZN(n20147) );
  AOI22_X1 U23102 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20152), .B1(
        n20561), .B2(n20151), .ZN(n20146) );
  OAI211_X1 U23103 ( .C1(n20565), .C2(n20149), .A(n20147), .B(n20146), .ZN(
        P1_U3063) );
  OAI22_X1 U23104 ( .A1(n20149), .A2(n20576), .B1(n20360), .B2(n20148), .ZN(
        n20150) );
  INV_X1 U23105 ( .A(n20150), .ZN(n20154) );
  AOI22_X1 U23106 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n20152), .B1(
        n20569), .B2(n20151), .ZN(n20153) );
  OAI211_X1 U23107 ( .C1(n20510), .C2(n20183), .A(n20154), .B(n20153), .ZN(
        P1_U3064) );
  INV_X1 U23108 ( .A(n20155), .ZN(n20466) );
  NOR2_X1 U23109 ( .A1(n9754), .A2(n20156), .ZN(n20240) );
  NAND3_X1 U23110 ( .A1(n20240), .A2(n20524), .A3(n20406), .ZN(n20157) );
  OAI21_X1 U23111 ( .B1(n20158), .B2(n20466), .A(n20157), .ZN(n20179) );
  NAND3_X1 U23112 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n20368), .A3(
        n20757), .ZN(n20184) );
  NOR2_X1 U23113 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20184), .ZN(
        n20178) );
  AOI22_X1 U23114 ( .A1(n20516), .A2(n20179), .B1(n20515), .B2(n20178), .ZN(
        n20164) );
  AOI21_X1 U23115 ( .B1(n20183), .B2(n20203), .A(n20439), .ZN(n20159) );
  AOI21_X1 U23116 ( .B1(n20240), .B2(n20406), .A(n20159), .ZN(n20160) );
  NOR2_X1 U23117 ( .A1(n20160), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20162) );
  INV_X1 U23118 ( .A(n20183), .ZN(n20169) );
  AOI22_X1 U23119 ( .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n20180), .B1(
        n20169), .B2(n20475), .ZN(n20163) );
  OAI211_X1 U23120 ( .C1(n20478), .C2(n20203), .A(n20164), .B(n20163), .ZN(
        P1_U3065) );
  AOI22_X1 U23121 ( .A1(n20531), .A2(n20179), .B1(n20530), .B2(n20178), .ZN(
        n20166) );
  AOI22_X1 U23122 ( .A1(P1_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n20180), .B1(
        n20169), .B2(n20479), .ZN(n20165) );
  OAI211_X1 U23123 ( .C1(n20482), .C2(n20203), .A(n20166), .B(n20165), .ZN(
        P1_U3066) );
  AOI22_X1 U23124 ( .A1(n20537), .A2(n20179), .B1(n20536), .B2(n20178), .ZN(
        n20168) );
  AOI22_X1 U23125 ( .A1(P1_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n20180), .B1(
        n20169), .B2(n20483), .ZN(n20167) );
  OAI211_X1 U23126 ( .C1(n20486), .C2(n20203), .A(n20168), .B(n20167), .ZN(
        P1_U3067) );
  AOI22_X1 U23127 ( .A1(n20543), .A2(n20179), .B1(n20542), .B2(n20178), .ZN(
        n20171) );
  AOI22_X1 U23128 ( .A1(P1_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n20180), .B1(
        n20169), .B2(n20487), .ZN(n20170) );
  OAI211_X1 U23129 ( .C1(n20490), .C2(n20203), .A(n20171), .B(n20170), .ZN(
        P1_U3068) );
  AOI22_X1 U23130 ( .A1(n20549), .A2(n20179), .B1(n20548), .B2(n20178), .ZN(
        n20173) );
  AOI22_X1 U23131 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n20180), .B1(
        n20206), .B2(n20550), .ZN(n20172) );
  OAI211_X1 U23132 ( .C1(n20553), .C2(n20183), .A(n20173), .B(n20172), .ZN(
        P1_U3069) );
  AOI22_X1 U23133 ( .A1(n20555), .A2(n20179), .B1(n20554), .B2(n20178), .ZN(
        n20175) );
  INV_X1 U23134 ( .A(n20498), .ZN(n20556) );
  AOI22_X1 U23135 ( .A1(P1_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n20180), .B1(
        n20206), .B2(n20556), .ZN(n20174) );
  OAI211_X1 U23136 ( .C1(n20559), .C2(n20183), .A(n20175), .B(n20174), .ZN(
        P1_U3070) );
  AOI22_X1 U23137 ( .A1(n20561), .A2(n20179), .B1(n20560), .B2(n20178), .ZN(
        n20177) );
  AOI22_X1 U23138 ( .A1(P1_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n20180), .B1(
        n20206), .B2(n20562), .ZN(n20176) );
  OAI211_X1 U23139 ( .C1(n20565), .C2(n20183), .A(n20177), .B(n20176), .ZN(
        P1_U3071) );
  AOI22_X1 U23140 ( .A1(n20569), .A2(n20179), .B1(n20567), .B2(n20178), .ZN(
        n20182) );
  INV_X1 U23141 ( .A(n20510), .ZN(n20570) );
  AOI22_X1 U23142 ( .A1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n20180), .B1(
        n20206), .B2(n20570), .ZN(n20181) );
  OAI211_X1 U23143 ( .C1(n20576), .C2(n20183), .A(n20182), .B(n20181), .ZN(
        P1_U3072) );
  NOR2_X1 U23144 ( .A1(n20435), .A2(n20184), .ZN(n20204) );
  AOI21_X1 U23145 ( .B1(n20240), .B2(n20436), .A(n20204), .ZN(n20185) );
  OAI22_X1 U23146 ( .A1(n20185), .A2(n20518), .B1(n20184), .B2(n12396), .ZN(
        n20205) );
  AOI22_X1 U23147 ( .A1(n20516), .A2(n20205), .B1(n20515), .B2(n20204), .ZN(
        n20190) );
  INV_X1 U23148 ( .A(n20184), .ZN(n20188) );
  OAI21_X1 U23149 ( .B1(n20239), .B2(n20186), .A(n20185), .ZN(n20187) );
  OAI211_X1 U23150 ( .C1(n20524), .C2(n20188), .A(n20523), .B(n20187), .ZN(
        n20207) );
  AOI22_X1 U23151 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n20207), .B1(
        n20206), .B2(n20475), .ZN(n20189) );
  OAI211_X1 U23152 ( .C1(n20478), .C2(n20238), .A(n20190), .B(n20189), .ZN(
        P1_U3073) );
  AOI22_X1 U23153 ( .A1(n20531), .A2(n20205), .B1(n20530), .B2(n20204), .ZN(
        n20192) );
  AOI22_X1 U23154 ( .A1(P1_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n20207), .B1(
        n20206), .B2(n20479), .ZN(n20191) );
  OAI211_X1 U23155 ( .C1(n20482), .C2(n20238), .A(n20192), .B(n20191), .ZN(
        P1_U3074) );
  AOI22_X1 U23156 ( .A1(n20537), .A2(n20205), .B1(n20536), .B2(n20204), .ZN(
        n20194) );
  INV_X1 U23157 ( .A(n20238), .ZN(n20230) );
  INV_X1 U23158 ( .A(n20486), .ZN(n20538) );
  AOI22_X1 U23159 ( .A1(P1_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n20207), .B1(
        n20230), .B2(n20538), .ZN(n20193) );
  OAI211_X1 U23160 ( .C1(n20541), .C2(n20203), .A(n20194), .B(n20193), .ZN(
        P1_U3075) );
  AOI22_X1 U23161 ( .A1(n20543), .A2(n20205), .B1(n20542), .B2(n20204), .ZN(
        n20196) );
  INV_X1 U23162 ( .A(n20490), .ZN(n20544) );
  AOI22_X1 U23163 ( .A1(P1_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20207), .B1(
        n20230), .B2(n20544), .ZN(n20195) );
  OAI211_X1 U23164 ( .C1(n20547), .C2(n20203), .A(n20196), .B(n20195), .ZN(
        P1_U3076) );
  AOI22_X1 U23165 ( .A1(n20549), .A2(n20205), .B1(n20548), .B2(n20204), .ZN(
        n20198) );
  AOI22_X1 U23166 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n20207), .B1(
        n20206), .B2(n20491), .ZN(n20197) );
  OAI211_X1 U23167 ( .C1(n20494), .C2(n20238), .A(n20198), .B(n20197), .ZN(
        P1_U3077) );
  AOI22_X1 U23168 ( .A1(n20555), .A2(n20205), .B1(n20554), .B2(n20204), .ZN(
        n20200) );
  AOI22_X1 U23169 ( .A1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20207), .B1(
        n20206), .B2(n20495), .ZN(n20199) );
  OAI211_X1 U23170 ( .C1(n20498), .C2(n20238), .A(n20200), .B(n20199), .ZN(
        P1_U3078) );
  AOI22_X1 U23171 ( .A1(n20561), .A2(n20205), .B1(n20560), .B2(n20204), .ZN(
        n20202) );
  AOI22_X1 U23172 ( .A1(P1_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n20207), .B1(
        n20230), .B2(n20562), .ZN(n20201) );
  OAI211_X1 U23173 ( .C1(n20565), .C2(n20203), .A(n20202), .B(n20201), .ZN(
        P1_U3079) );
  AOI22_X1 U23174 ( .A1(n20569), .A2(n20205), .B1(n20567), .B2(n20204), .ZN(
        n20209) );
  AOI22_X1 U23175 ( .A1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n20207), .B1(
        n20206), .B2(n20505), .ZN(n20208) );
  OAI211_X1 U23176 ( .C1(n20510), .C2(n20238), .A(n20209), .B(n20208), .ZN(
        P1_U3080) );
  NOR2_X1 U23177 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20241), .ZN(
        n20233) );
  AOI22_X1 U23178 ( .A1(n20255), .A2(n20526), .B1(n20515), .B2(n20233), .ZN(
        n20219) );
  NAND3_X1 U23179 ( .A1(n20266), .A2(n20238), .A3(n20524), .ZN(n20210) );
  NAND2_X1 U23180 ( .A1(n20210), .A2(n20403), .ZN(n20214) );
  NAND2_X1 U23181 ( .A1(n20240), .A2(n20465), .ZN(n20216) );
  INV_X1 U23182 ( .A(n20233), .ZN(n20211) );
  AOI22_X1 U23183 ( .A1(n20214), .A2(n20216), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20211), .ZN(n20213) );
  NAND3_X1 U23184 ( .A1(n20473), .A2(n20213), .A3(n20212), .ZN(n20235) );
  INV_X1 U23185 ( .A(n20214), .ZN(n20217) );
  OAI22_X1 U23186 ( .A1(n20217), .A2(n20216), .B1(n20215), .B2(n20466), .ZN(
        n20234) );
  AOI22_X1 U23187 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n20235), .B1(
        n20516), .B2(n20234), .ZN(n20218) );
  OAI211_X1 U23188 ( .C1(n20529), .C2(n20238), .A(n20219), .B(n20218), .ZN(
        P1_U3081) );
  INV_X1 U23189 ( .A(n20482), .ZN(n20532) );
  AOI22_X1 U23190 ( .A1(n20255), .A2(n20532), .B1(n20530), .B2(n20233), .ZN(
        n20221) );
  AOI22_X1 U23191 ( .A1(P1_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n20235), .B1(
        n20531), .B2(n20234), .ZN(n20220) );
  OAI211_X1 U23192 ( .C1(n20535), .C2(n20238), .A(n20221), .B(n20220), .ZN(
        P1_U3082) );
  AOI22_X1 U23193 ( .A1(n20230), .A2(n20483), .B1(n20536), .B2(n20233), .ZN(
        n20223) );
  AOI22_X1 U23194 ( .A1(P1_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n20235), .B1(
        n20537), .B2(n20234), .ZN(n20222) );
  OAI211_X1 U23195 ( .C1(n20486), .C2(n20266), .A(n20223), .B(n20222), .ZN(
        P1_U3083) );
  AOI22_X1 U23196 ( .A1(n20255), .A2(n20544), .B1(n20542), .B2(n20233), .ZN(
        n20225) );
  AOI22_X1 U23197 ( .A1(P1_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n20235), .B1(
        n20543), .B2(n20234), .ZN(n20224) );
  OAI211_X1 U23198 ( .C1(n20547), .C2(n20238), .A(n20225), .B(n20224), .ZN(
        P1_U3084) );
  AOI22_X1 U23199 ( .A1(n20255), .A2(n20550), .B1(n20548), .B2(n20233), .ZN(
        n20227) );
  AOI22_X1 U23200 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n20235), .B1(
        n20549), .B2(n20234), .ZN(n20226) );
  OAI211_X1 U23201 ( .C1(n20553), .C2(n20238), .A(n20227), .B(n20226), .ZN(
        P1_U3085) );
  AOI22_X1 U23202 ( .A1(n20255), .A2(n20556), .B1(n20554), .B2(n20233), .ZN(
        n20229) );
  AOI22_X1 U23203 ( .A1(P1_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n20235), .B1(
        n20555), .B2(n20234), .ZN(n20228) );
  OAI211_X1 U23204 ( .C1(n20559), .C2(n20238), .A(n20229), .B(n20228), .ZN(
        P1_U3086) );
  AOI22_X1 U23205 ( .A1(n20230), .A2(n20499), .B1(n20560), .B2(n20233), .ZN(
        n20232) );
  AOI22_X1 U23206 ( .A1(P1_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n20235), .B1(
        n20561), .B2(n20234), .ZN(n20231) );
  OAI211_X1 U23207 ( .C1(n20502), .C2(n20266), .A(n20232), .B(n20231), .ZN(
        P1_U3087) );
  AOI22_X1 U23208 ( .A1(n20255), .A2(n20570), .B1(n20567), .B2(n20233), .ZN(
        n20237) );
  AOI22_X1 U23209 ( .A1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n20235), .B1(
        n20569), .B2(n20234), .ZN(n20236) );
  OAI211_X1 U23210 ( .C1(n20576), .C2(n20238), .A(n20237), .B(n20236), .ZN(
        P1_U3088) );
  AOI21_X1 U23211 ( .B1(n20240), .B2(n20512), .A(n20261), .ZN(n20242) );
  OAI22_X1 U23212 ( .A1(n20242), .A2(n20518), .B1(n20241), .B2(n12396), .ZN(
        n20262) );
  AOI22_X1 U23213 ( .A1(n20516), .A2(n20262), .B1(n20515), .B2(n20261), .ZN(
        n20246) );
  OAI21_X1 U23214 ( .B1(n20244), .B2(n20243), .A(n20523), .ZN(n20263) );
  AOI22_X1 U23215 ( .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n20263), .B1(
        n20255), .B2(n20475), .ZN(n20245) );
  OAI211_X1 U23216 ( .C1(n20478), .C2(n20258), .A(n20246), .B(n20245), .ZN(
        P1_U3089) );
  AOI22_X1 U23217 ( .A1(n20531), .A2(n20262), .B1(n20530), .B2(n20261), .ZN(
        n20248) );
  AOI22_X1 U23218 ( .A1(P1_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n20263), .B1(
        n20255), .B2(n20479), .ZN(n20247) );
  OAI211_X1 U23219 ( .C1(n20482), .C2(n20258), .A(n20248), .B(n20247), .ZN(
        P1_U3090) );
  AOI22_X1 U23220 ( .A1(n20537), .A2(n20262), .B1(n20536), .B2(n20261), .ZN(
        n20250) );
  AOI22_X1 U23221 ( .A1(P1_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n20263), .B1(
        n20255), .B2(n20483), .ZN(n20249) );
  OAI211_X1 U23222 ( .C1(n20486), .C2(n20258), .A(n20250), .B(n20249), .ZN(
        P1_U3091) );
  AOI22_X1 U23223 ( .A1(n20543), .A2(n20262), .B1(n20542), .B2(n20261), .ZN(
        n20252) );
  AOI22_X1 U23224 ( .A1(P1_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n20263), .B1(
        n20255), .B2(n20487), .ZN(n20251) );
  OAI211_X1 U23225 ( .C1(n20490), .C2(n20258), .A(n20252), .B(n20251), .ZN(
        P1_U3092) );
  AOI22_X1 U23226 ( .A1(n20549), .A2(n20262), .B1(n20548), .B2(n20261), .ZN(
        n20254) );
  AOI22_X1 U23227 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n20263), .B1(
        n20292), .B2(n20550), .ZN(n20253) );
  OAI211_X1 U23228 ( .C1(n20553), .C2(n20266), .A(n20254), .B(n20253), .ZN(
        P1_U3093) );
  AOI22_X1 U23229 ( .A1(n20555), .A2(n20262), .B1(n20554), .B2(n20261), .ZN(
        n20257) );
  AOI22_X1 U23230 ( .A1(P1_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n20263), .B1(
        n20255), .B2(n20495), .ZN(n20256) );
  OAI211_X1 U23231 ( .C1(n20498), .C2(n20258), .A(n20257), .B(n20256), .ZN(
        P1_U3094) );
  AOI22_X1 U23232 ( .A1(n20561), .A2(n20262), .B1(n20560), .B2(n20261), .ZN(
        n20260) );
  AOI22_X1 U23233 ( .A1(P1_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n20263), .B1(
        n20292), .B2(n20562), .ZN(n20259) );
  OAI211_X1 U23234 ( .C1(n20565), .C2(n20266), .A(n20260), .B(n20259), .ZN(
        P1_U3095) );
  AOI22_X1 U23235 ( .A1(n20569), .A2(n20262), .B1(n20567), .B2(n20261), .ZN(
        n20265) );
  AOI22_X1 U23236 ( .A1(P1_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n20263), .B1(
        n20292), .B2(n20570), .ZN(n20264) );
  OAI211_X1 U23237 ( .C1(n20576), .C2(n20266), .A(n20265), .B(n20264), .ZN(
        P1_U3096) );
  INV_X1 U23238 ( .A(n20377), .ZN(n20371) );
  INV_X1 U23239 ( .A(n20267), .ZN(n20268) );
  NAND2_X1 U23240 ( .A1(n20269), .A2(n9754), .ZN(n20325) );
  INV_X1 U23241 ( .A(n20325), .ZN(n20369) );
  NAND3_X1 U23242 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n20321), .A3(
        n20757), .ZN(n20296) );
  NOR2_X1 U23243 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20296), .ZN(
        n20290) );
  AOI21_X1 U23244 ( .B1(n20369), .B2(n20406), .A(n20290), .ZN(n20272) );
  AND2_X1 U23245 ( .A1(n20270), .A2(n20326), .ZN(n20409) );
  INV_X1 U23246 ( .A(n20409), .ZN(n20411) );
  OAI22_X1 U23247 ( .A1(n20272), .A2(n20518), .B1(n20330), .B2(n20411), .ZN(
        n20291) );
  AOI22_X1 U23248 ( .A1(n20516), .A2(n20291), .B1(n20515), .B2(n20290), .ZN(
        n20277) );
  INV_X1 U23249 ( .A(n20320), .ZN(n20271) );
  OAI21_X1 U23250 ( .B1(n20271), .B2(n20292), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20273) );
  NAND2_X1 U23251 ( .A1(n20273), .A2(n20272), .ZN(n20274) );
  OAI211_X1 U23252 ( .C1(n20290), .C2(n20275), .A(n20328), .B(n20274), .ZN(
        n20293) );
  AOI22_X1 U23253 ( .A1(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n20293), .B1(
        n20292), .B2(n20475), .ZN(n20276) );
  OAI211_X1 U23254 ( .C1(n20478), .C2(n20320), .A(n20277), .B(n20276), .ZN(
        P1_U3097) );
  AOI22_X1 U23255 ( .A1(n20531), .A2(n20291), .B1(n20530), .B2(n20290), .ZN(
        n20279) );
  AOI22_X1 U23256 ( .A1(P1_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n20293), .B1(
        n20292), .B2(n20479), .ZN(n20278) );
  OAI211_X1 U23257 ( .C1(n20482), .C2(n20320), .A(n20279), .B(n20278), .ZN(
        P1_U3098) );
  AOI22_X1 U23258 ( .A1(n20537), .A2(n20291), .B1(n20536), .B2(n20290), .ZN(
        n20281) );
  AOI22_X1 U23259 ( .A1(P1_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n20293), .B1(
        n20292), .B2(n20483), .ZN(n20280) );
  OAI211_X1 U23260 ( .C1(n20486), .C2(n20320), .A(n20281), .B(n20280), .ZN(
        P1_U3099) );
  AOI22_X1 U23261 ( .A1(n20543), .A2(n20291), .B1(n20542), .B2(n20290), .ZN(
        n20283) );
  AOI22_X1 U23262 ( .A1(P1_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n20293), .B1(
        n20292), .B2(n20487), .ZN(n20282) );
  OAI211_X1 U23263 ( .C1(n20490), .C2(n20320), .A(n20283), .B(n20282), .ZN(
        P1_U3100) );
  AOI22_X1 U23264 ( .A1(n20549), .A2(n20291), .B1(n20548), .B2(n20290), .ZN(
        n20285) );
  AOI22_X1 U23265 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n20293), .B1(
        n20292), .B2(n20491), .ZN(n20284) );
  OAI211_X1 U23266 ( .C1(n20494), .C2(n20320), .A(n20285), .B(n20284), .ZN(
        P1_U3101) );
  AOI22_X1 U23267 ( .A1(n20555), .A2(n20291), .B1(n20554), .B2(n20290), .ZN(
        n20287) );
  AOI22_X1 U23268 ( .A1(P1_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n20293), .B1(
        n20292), .B2(n20495), .ZN(n20286) );
  OAI211_X1 U23269 ( .C1(n20498), .C2(n20320), .A(n20287), .B(n20286), .ZN(
        P1_U3102) );
  AOI22_X1 U23270 ( .A1(n20561), .A2(n20291), .B1(n20560), .B2(n20290), .ZN(
        n20289) );
  AOI22_X1 U23271 ( .A1(P1_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n20293), .B1(
        n20292), .B2(n20499), .ZN(n20288) );
  OAI211_X1 U23272 ( .C1(n20502), .C2(n20320), .A(n20289), .B(n20288), .ZN(
        P1_U3103) );
  AOI22_X1 U23273 ( .A1(n20569), .A2(n20291), .B1(n20567), .B2(n20290), .ZN(
        n20295) );
  AOI22_X1 U23274 ( .A1(P1_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n20293), .B1(
        n20292), .B2(n20505), .ZN(n20294) );
  OAI211_X1 U23275 ( .C1(n20510), .C2(n20320), .A(n20295), .B(n20294), .ZN(
        P1_U3104) );
  NOR2_X1 U23276 ( .A1(n20435), .A2(n20296), .ZN(n20314) );
  AOI21_X1 U23277 ( .B1(n20369), .B2(n20436), .A(n20314), .ZN(n20297) );
  OAI22_X1 U23278 ( .A1(n20297), .A2(n20518), .B1(n20296), .B2(n12396), .ZN(
        n20315) );
  AOI22_X1 U23279 ( .A1(n20516), .A2(n20315), .B1(n20515), .B2(n20314), .ZN(
        n20301) );
  INV_X1 U23280 ( .A(n20296), .ZN(n20299) );
  OAI211_X1 U23281 ( .C1(n20377), .C2(n20439), .A(n20524), .B(n20297), .ZN(
        n20298) );
  OAI211_X1 U23282 ( .C1(n20524), .C2(n20299), .A(n20523), .B(n20298), .ZN(
        n20317) );
  AOI22_X1 U23283 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n20317), .B1(
        n20316), .B2(n20526), .ZN(n20300) );
  OAI211_X1 U23284 ( .C1(n20529), .C2(n20320), .A(n20301), .B(n20300), .ZN(
        P1_U3105) );
  AOI22_X1 U23285 ( .A1(n20531), .A2(n20315), .B1(n20530), .B2(n20314), .ZN(
        n20303) );
  AOI22_X1 U23286 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n20317), .B1(
        n20316), .B2(n20532), .ZN(n20302) );
  OAI211_X1 U23287 ( .C1(n20535), .C2(n20320), .A(n20303), .B(n20302), .ZN(
        P1_U3106) );
  AOI22_X1 U23288 ( .A1(n20537), .A2(n20315), .B1(n20536), .B2(n20314), .ZN(
        n20305) );
  AOI22_X1 U23289 ( .A1(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n20317), .B1(
        n20316), .B2(n20538), .ZN(n20304) );
  OAI211_X1 U23290 ( .C1(n20541), .C2(n20320), .A(n20305), .B(n20304), .ZN(
        P1_U3107) );
  AOI22_X1 U23291 ( .A1(n20543), .A2(n20315), .B1(n20542), .B2(n20314), .ZN(
        n20307) );
  AOI22_X1 U23292 ( .A1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n20317), .B1(
        n20316), .B2(n20544), .ZN(n20306) );
  OAI211_X1 U23293 ( .C1(n20547), .C2(n20320), .A(n20307), .B(n20306), .ZN(
        P1_U3108) );
  AOI22_X1 U23294 ( .A1(n20549), .A2(n20315), .B1(n20548), .B2(n20314), .ZN(
        n20309) );
  AOI22_X1 U23295 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n20317), .B1(
        n20316), .B2(n20550), .ZN(n20308) );
  OAI211_X1 U23296 ( .C1(n20553), .C2(n20320), .A(n20309), .B(n20308), .ZN(
        P1_U3109) );
  AOI22_X1 U23297 ( .A1(n20555), .A2(n20315), .B1(n20554), .B2(n20314), .ZN(
        n20311) );
  AOI22_X1 U23298 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n20317), .B1(
        n20316), .B2(n20556), .ZN(n20310) );
  OAI211_X1 U23299 ( .C1(n20559), .C2(n20320), .A(n20311), .B(n20310), .ZN(
        P1_U3110) );
  AOI22_X1 U23300 ( .A1(n20561), .A2(n20315), .B1(n20560), .B2(n20314), .ZN(
        n20313) );
  AOI22_X1 U23301 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n20317), .B1(
        n20316), .B2(n20562), .ZN(n20312) );
  OAI211_X1 U23302 ( .C1(n20565), .C2(n20320), .A(n20313), .B(n20312), .ZN(
        P1_U3111) );
  AOI22_X1 U23303 ( .A1(n20569), .A2(n20315), .B1(n20567), .B2(n20314), .ZN(
        n20319) );
  AOI22_X1 U23304 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n20317), .B1(
        n20316), .B2(n20570), .ZN(n20318) );
  OAI211_X1 U23305 ( .C1(n20576), .C2(n20320), .A(n20319), .B(n20318), .ZN(
        P1_U3112) );
  NAND3_X1 U23306 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n20321), .ZN(n20370) );
  OR2_X1 U23307 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20370), .ZN(
        n20359) );
  OAI22_X1 U23308 ( .A1(n20366), .A2(n20529), .B1(n20322), .B2(n20359), .ZN(
        n20323) );
  INV_X1 U23309 ( .A(n20323), .ZN(n20334) );
  NAND3_X1 U23310 ( .A1(n20391), .A2(n20366), .A3(n20524), .ZN(n20324) );
  NAND2_X1 U23311 ( .A1(n20324), .A2(n20403), .ZN(n20329) );
  OR2_X1 U23312 ( .A1(n20325), .A2(n20406), .ZN(n20331) );
  AOI22_X1 U23313 ( .A1(n20329), .A2(n20331), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20359), .ZN(n20327) );
  OR2_X1 U23314 ( .A1(n20326), .A2(n20368), .ZN(n20467) );
  NAND2_X1 U23315 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20467), .ZN(n20472) );
  NAND3_X1 U23316 ( .A1(n20328), .A2(n20327), .A3(n20472), .ZN(n20363) );
  INV_X1 U23317 ( .A(n20329), .ZN(n20332) );
  OAI22_X1 U23318 ( .A1(n20332), .A2(n20331), .B1(n20330), .B2(n20467), .ZN(
        n20362) );
  AOI22_X1 U23319 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n20363), .B1(
        n20516), .B2(n20362), .ZN(n20333) );
  OAI211_X1 U23320 ( .C1(n20478), .C2(n20391), .A(n20334), .B(n20333), .ZN(
        P1_U3113) );
  OAI22_X1 U23321 ( .A1(n20391), .A2(n20482), .B1(n20335), .B2(n20359), .ZN(
        n20336) );
  INV_X1 U23322 ( .A(n20336), .ZN(n20338) );
  AOI22_X1 U23323 ( .A1(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n20363), .B1(
        n20531), .B2(n20362), .ZN(n20337) );
  OAI211_X1 U23324 ( .C1(n20535), .C2(n20366), .A(n20338), .B(n20337), .ZN(
        P1_U3114) );
  OAI22_X1 U23325 ( .A1(n20391), .A2(n20486), .B1(n20339), .B2(n20359), .ZN(
        n20340) );
  INV_X1 U23326 ( .A(n20340), .ZN(n20342) );
  AOI22_X1 U23327 ( .A1(P1_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n20363), .B1(
        n20537), .B2(n20362), .ZN(n20341) );
  OAI211_X1 U23328 ( .C1(n20541), .C2(n20366), .A(n20342), .B(n20341), .ZN(
        P1_U3115) );
  OAI22_X1 U23329 ( .A1(n20391), .A2(n20490), .B1(n20343), .B2(n20359), .ZN(
        n20344) );
  INV_X1 U23330 ( .A(n20344), .ZN(n20346) );
  AOI22_X1 U23331 ( .A1(P1_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n20363), .B1(
        n20543), .B2(n20362), .ZN(n20345) );
  OAI211_X1 U23332 ( .C1(n20547), .C2(n20366), .A(n20346), .B(n20345), .ZN(
        P1_U3116) );
  OAI22_X1 U23333 ( .A1(n20391), .A2(n20494), .B1(n20347), .B2(n20359), .ZN(
        n20348) );
  INV_X1 U23334 ( .A(n20348), .ZN(n20350) );
  AOI22_X1 U23335 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n20363), .B1(
        n20549), .B2(n20362), .ZN(n20349) );
  OAI211_X1 U23336 ( .C1(n20553), .C2(n20366), .A(n20350), .B(n20349), .ZN(
        P1_U3117) );
  OAI22_X1 U23337 ( .A1(n20391), .A2(n20498), .B1(n20351), .B2(n20359), .ZN(
        n20352) );
  INV_X1 U23338 ( .A(n20352), .ZN(n20354) );
  AOI22_X1 U23339 ( .A1(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n20363), .B1(
        n20555), .B2(n20362), .ZN(n20353) );
  OAI211_X1 U23340 ( .C1(n20559), .C2(n20366), .A(n20354), .B(n20353), .ZN(
        P1_U3118) );
  OAI22_X1 U23341 ( .A1(n20366), .A2(n20565), .B1(n20355), .B2(n20359), .ZN(
        n20356) );
  INV_X1 U23342 ( .A(n20356), .ZN(n20358) );
  AOI22_X1 U23343 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n20363), .B1(
        n20561), .B2(n20362), .ZN(n20357) );
  OAI211_X1 U23344 ( .C1(n20502), .C2(n20391), .A(n20358), .B(n20357), .ZN(
        P1_U3119) );
  OAI22_X1 U23345 ( .A1(n20391), .A2(n20510), .B1(n20360), .B2(n20359), .ZN(
        n20361) );
  INV_X1 U23346 ( .A(n20361), .ZN(n20365) );
  AOI22_X1 U23347 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n20363), .B1(
        n20569), .B2(n20362), .ZN(n20364) );
  OAI211_X1 U23348 ( .C1(n20576), .C2(n20366), .A(n20365), .B(n20364), .ZN(
        P1_U3120) );
  NOR2_X1 U23349 ( .A1(n20368), .A2(n20367), .ZN(n20394) );
  AOI21_X1 U23350 ( .B1(n20369), .B2(n20512), .A(n20394), .ZN(n20372) );
  OAI22_X1 U23351 ( .A1(n20372), .A2(n20518), .B1(n20370), .B2(n12396), .ZN(
        n20395) );
  AOI22_X1 U23352 ( .A1(n20516), .A2(n20395), .B1(n20515), .B2(n20394), .ZN(
        n20379) );
  INV_X1 U23353 ( .A(n20370), .ZN(n20375) );
  OAI21_X1 U23354 ( .B1(n20371), .B2(n20518), .A(n20517), .ZN(n20373) );
  NAND2_X1 U23355 ( .A1(n20373), .A2(n20372), .ZN(n20374) );
  OAI211_X1 U23356 ( .C1(n20524), .C2(n20375), .A(n20523), .B(n20374), .ZN(
        n20397) );
  INV_X1 U23357 ( .A(n20433), .ZN(n20388) );
  AOI22_X1 U23358 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n20397), .B1(
        n20388), .B2(n20526), .ZN(n20378) );
  OAI211_X1 U23359 ( .C1(n20529), .C2(n20391), .A(n20379), .B(n20378), .ZN(
        P1_U3121) );
  AOI22_X1 U23360 ( .A1(n20531), .A2(n20395), .B1(n20530), .B2(n20394), .ZN(
        n20381) );
  INV_X1 U23361 ( .A(n20391), .ZN(n20396) );
  AOI22_X1 U23362 ( .A1(P1_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n20397), .B1(
        n20396), .B2(n20479), .ZN(n20380) );
  OAI211_X1 U23363 ( .C1(n20482), .C2(n20433), .A(n20381), .B(n20380), .ZN(
        P1_U3122) );
  AOI22_X1 U23364 ( .A1(n20537), .A2(n20395), .B1(n20536), .B2(n20394), .ZN(
        n20383) );
  AOI22_X1 U23365 ( .A1(P1_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n20397), .B1(
        n20388), .B2(n20538), .ZN(n20382) );
  OAI211_X1 U23366 ( .C1(n20541), .C2(n20391), .A(n20383), .B(n20382), .ZN(
        P1_U3123) );
  AOI22_X1 U23367 ( .A1(n20543), .A2(n20395), .B1(n20542), .B2(n20394), .ZN(
        n20385) );
  AOI22_X1 U23368 ( .A1(P1_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n20397), .B1(
        n20388), .B2(n20544), .ZN(n20384) );
  OAI211_X1 U23369 ( .C1(n20547), .C2(n20391), .A(n20385), .B(n20384), .ZN(
        P1_U3124) );
  AOI22_X1 U23370 ( .A1(n20549), .A2(n20395), .B1(n20548), .B2(n20394), .ZN(
        n20387) );
  AOI22_X1 U23371 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n20397), .B1(
        n20388), .B2(n20550), .ZN(n20386) );
  OAI211_X1 U23372 ( .C1(n20553), .C2(n20391), .A(n20387), .B(n20386), .ZN(
        P1_U3125) );
  AOI22_X1 U23373 ( .A1(n20555), .A2(n20395), .B1(n20554), .B2(n20394), .ZN(
        n20390) );
  AOI22_X1 U23374 ( .A1(P1_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n20397), .B1(
        n20388), .B2(n20556), .ZN(n20389) );
  OAI211_X1 U23375 ( .C1(n20559), .C2(n20391), .A(n20390), .B(n20389), .ZN(
        P1_U3126) );
  AOI22_X1 U23376 ( .A1(n20561), .A2(n20395), .B1(n20560), .B2(n20394), .ZN(
        n20393) );
  AOI22_X1 U23377 ( .A1(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n20397), .B1(
        n20396), .B2(n20499), .ZN(n20392) );
  OAI211_X1 U23378 ( .C1(n20502), .C2(n20433), .A(n20393), .B(n20392), .ZN(
        P1_U3127) );
  AOI22_X1 U23379 ( .A1(n20569), .A2(n20395), .B1(n20567), .B2(n20394), .ZN(
        n20399) );
  AOI22_X1 U23380 ( .A1(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n20397), .B1(
        n20396), .B2(n20505), .ZN(n20398) );
  OAI211_X1 U23381 ( .C1(n20510), .C2(n20433), .A(n20399), .B(n20398), .ZN(
        P1_U3128) );
  NAND3_X1 U23382 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n20757), .ZN(n20437) );
  NOR2_X1 U23383 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20437), .ZN(
        n20428) );
  AOI22_X1 U23384 ( .A1(n20458), .A2(n20526), .B1(n20515), .B2(n20428), .ZN(
        n20415) );
  INV_X1 U23385 ( .A(n20458), .ZN(n20402) );
  NAND3_X1 U23386 ( .A1(n20402), .A2(n20524), .A3(n20433), .ZN(n20404) );
  NAND2_X1 U23387 ( .A1(n20404), .A2(n20403), .ZN(n20410) );
  NOR2_X1 U23388 ( .A1(n9754), .A2(n20405), .ZN(n20513) );
  NAND2_X1 U23389 ( .A1(n20513), .A2(n20406), .ZN(n20412) );
  INV_X1 U23390 ( .A(n20428), .ZN(n20407) );
  AOI22_X1 U23391 ( .A1(n20410), .A2(n20412), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20407), .ZN(n20408) );
  INV_X1 U23392 ( .A(n20410), .ZN(n20413) );
  AOI22_X1 U23393 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n20430), .B1(
        n20516), .B2(n20429), .ZN(n20414) );
  OAI211_X1 U23394 ( .C1(n20529), .C2(n20433), .A(n20415), .B(n20414), .ZN(
        P1_U3129) );
  AOI22_X1 U23395 ( .A1(n20458), .A2(n20532), .B1(n20530), .B2(n20428), .ZN(
        n20417) );
  AOI22_X1 U23396 ( .A1(P1_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n20430), .B1(
        n20531), .B2(n20429), .ZN(n20416) );
  OAI211_X1 U23397 ( .C1(n20535), .C2(n20433), .A(n20417), .B(n20416), .ZN(
        P1_U3130) );
  AOI22_X1 U23398 ( .A1(n20458), .A2(n20538), .B1(n20536), .B2(n20428), .ZN(
        n20419) );
  AOI22_X1 U23399 ( .A1(P1_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n20430), .B1(
        n20537), .B2(n20429), .ZN(n20418) );
  OAI211_X1 U23400 ( .C1(n20541), .C2(n20433), .A(n20419), .B(n20418), .ZN(
        P1_U3131) );
  AOI22_X1 U23401 ( .A1(n20458), .A2(n20544), .B1(n20542), .B2(n20428), .ZN(
        n20421) );
  AOI22_X1 U23402 ( .A1(P1_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n20430), .B1(
        n20543), .B2(n20429), .ZN(n20420) );
  OAI211_X1 U23403 ( .C1(n20547), .C2(n20433), .A(n20421), .B(n20420), .ZN(
        P1_U3132) );
  AOI22_X1 U23404 ( .A1(n20458), .A2(n20550), .B1(n20548), .B2(n20428), .ZN(
        n20423) );
  AOI22_X1 U23405 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n20430), .B1(
        n20549), .B2(n20429), .ZN(n20422) );
  OAI211_X1 U23406 ( .C1(n20553), .C2(n20433), .A(n20423), .B(n20422), .ZN(
        P1_U3133) );
  AOI22_X1 U23407 ( .A1(n20458), .A2(n20556), .B1(n20554), .B2(n20428), .ZN(
        n20425) );
  AOI22_X1 U23408 ( .A1(P1_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n20430), .B1(
        n20555), .B2(n20429), .ZN(n20424) );
  OAI211_X1 U23409 ( .C1(n20559), .C2(n20433), .A(n20425), .B(n20424), .ZN(
        P1_U3134) );
  AOI22_X1 U23410 ( .A1(n20458), .A2(n20562), .B1(n20560), .B2(n20428), .ZN(
        n20427) );
  AOI22_X1 U23411 ( .A1(P1_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n20430), .B1(
        n20561), .B2(n20429), .ZN(n20426) );
  OAI211_X1 U23412 ( .C1(n20565), .C2(n20433), .A(n20427), .B(n20426), .ZN(
        P1_U3135) );
  AOI22_X1 U23413 ( .A1(n20458), .A2(n20570), .B1(n20567), .B2(n20428), .ZN(
        n20432) );
  AOI22_X1 U23414 ( .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n20430), .B1(
        n20569), .B2(n20429), .ZN(n20431) );
  OAI211_X1 U23415 ( .C1(n20576), .C2(n20433), .A(n20432), .B(n20431), .ZN(
        P1_U3136) );
  NOR2_X1 U23416 ( .A1(n20435), .A2(n20437), .ZN(n20456) );
  AOI21_X1 U23417 ( .B1(n20513), .B2(n20436), .A(n20456), .ZN(n20438) );
  OAI22_X1 U23418 ( .A1(n20438), .A2(n20518), .B1(n20437), .B2(n12396), .ZN(
        n20457) );
  AOI22_X1 U23419 ( .A1(n20516), .A2(n20457), .B1(n20515), .B2(n20456), .ZN(
        n20443) );
  INV_X1 U23420 ( .A(n20437), .ZN(n20441) );
  OAI211_X1 U23421 ( .C1(n20462), .C2(n20439), .A(n20524), .B(n20438), .ZN(
        n20440) );
  OAI211_X1 U23422 ( .C1(n20524), .C2(n20441), .A(n20523), .B(n20440), .ZN(
        n20459) );
  AOI22_X1 U23423 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n20459), .B1(
        n20458), .B2(n20475), .ZN(n20442) );
  OAI211_X1 U23424 ( .C1(n20478), .C2(n20468), .A(n20443), .B(n20442), .ZN(
        P1_U3137) );
  AOI22_X1 U23425 ( .A1(n20531), .A2(n20457), .B1(n20530), .B2(n20456), .ZN(
        n20445) );
  AOI22_X1 U23426 ( .A1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n20459), .B1(
        n20458), .B2(n20479), .ZN(n20444) );
  OAI211_X1 U23427 ( .C1(n20482), .C2(n20468), .A(n20445), .B(n20444), .ZN(
        P1_U3138) );
  AOI22_X1 U23428 ( .A1(n20537), .A2(n20457), .B1(n20536), .B2(n20456), .ZN(
        n20447) );
  AOI22_X1 U23429 ( .A1(P1_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n20459), .B1(
        n20458), .B2(n20483), .ZN(n20446) );
  OAI211_X1 U23430 ( .C1(n20486), .C2(n20468), .A(n20447), .B(n20446), .ZN(
        P1_U3139) );
  AOI22_X1 U23431 ( .A1(n20543), .A2(n20457), .B1(n20542), .B2(n20456), .ZN(
        n20449) );
  AOI22_X1 U23432 ( .A1(P1_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n20459), .B1(
        n20458), .B2(n20487), .ZN(n20448) );
  OAI211_X1 U23433 ( .C1(n20490), .C2(n20468), .A(n20449), .B(n20448), .ZN(
        P1_U3140) );
  AOI22_X1 U23434 ( .A1(n20549), .A2(n20457), .B1(n20548), .B2(n20456), .ZN(
        n20451) );
  AOI22_X1 U23435 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n20459), .B1(
        n20458), .B2(n20491), .ZN(n20450) );
  OAI211_X1 U23436 ( .C1(n20494), .C2(n20468), .A(n20451), .B(n20450), .ZN(
        P1_U3141) );
  AOI22_X1 U23437 ( .A1(n20555), .A2(n20457), .B1(n20554), .B2(n20456), .ZN(
        n20453) );
  AOI22_X1 U23438 ( .A1(P1_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n20459), .B1(
        n20458), .B2(n20495), .ZN(n20452) );
  OAI211_X1 U23439 ( .C1(n20498), .C2(n20468), .A(n20453), .B(n20452), .ZN(
        P1_U3142) );
  AOI22_X1 U23440 ( .A1(n20561), .A2(n20457), .B1(n20560), .B2(n20456), .ZN(
        n20455) );
  AOI22_X1 U23441 ( .A1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n20459), .B1(
        n20458), .B2(n20499), .ZN(n20454) );
  OAI211_X1 U23442 ( .C1(n20502), .C2(n20468), .A(n20455), .B(n20454), .ZN(
        P1_U3143) );
  AOI22_X1 U23443 ( .A1(n20569), .A2(n20457), .B1(n20567), .B2(n20456), .ZN(
        n20461) );
  AOI22_X1 U23444 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n20459), .B1(
        n20458), .B2(n20505), .ZN(n20460) );
  OAI211_X1 U23445 ( .C1(n20510), .C2(n20468), .A(n20461), .B(n20460), .ZN(
        P1_U3144) );
  INV_X1 U23446 ( .A(n20462), .ZN(n20519) );
  INV_X1 U23447 ( .A(n20463), .ZN(n20464) );
  NAND2_X1 U23448 ( .A1(n20513), .A2(n20465), .ZN(n20470) );
  OAI22_X1 U23449 ( .A1(n20470), .A2(n20518), .B1(n20467), .B2(n20466), .ZN(
        n20504) );
  NOR2_X1 U23450 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20514), .ZN(
        n20503) );
  AOI22_X1 U23451 ( .A1(n20516), .A2(n20504), .B1(n20515), .B2(n20503), .ZN(
        n20477) );
  INV_X1 U23452 ( .A(n20575), .ZN(n20469) );
  OAI21_X1 U23453 ( .B1(n20469), .B2(n20506), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20471) );
  AOI21_X1 U23454 ( .B1(n20471), .B2(n20470), .A(P1_STATE2_REG_3__SCAN_IN), 
        .ZN(n20474) );
  AOI22_X1 U23455 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n20507), .B1(
        n20506), .B2(n20475), .ZN(n20476) );
  OAI211_X1 U23456 ( .C1(n20478), .C2(n20575), .A(n20477), .B(n20476), .ZN(
        P1_U3145) );
  AOI22_X1 U23457 ( .A1(n20531), .A2(n20504), .B1(n20530), .B2(n20503), .ZN(
        n20481) );
  AOI22_X1 U23458 ( .A1(P1_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n20507), .B1(
        n20506), .B2(n20479), .ZN(n20480) );
  OAI211_X1 U23459 ( .C1(n20482), .C2(n20575), .A(n20481), .B(n20480), .ZN(
        P1_U3146) );
  AOI22_X1 U23460 ( .A1(n20537), .A2(n20504), .B1(n20536), .B2(n20503), .ZN(
        n20485) );
  AOI22_X1 U23461 ( .A1(P1_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n20507), .B1(
        n20506), .B2(n20483), .ZN(n20484) );
  OAI211_X1 U23462 ( .C1(n20486), .C2(n20575), .A(n20485), .B(n20484), .ZN(
        P1_U3147) );
  AOI22_X1 U23463 ( .A1(n20543), .A2(n20504), .B1(n20542), .B2(n20503), .ZN(
        n20489) );
  AOI22_X1 U23464 ( .A1(P1_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n20507), .B1(
        n20506), .B2(n20487), .ZN(n20488) );
  OAI211_X1 U23465 ( .C1(n20490), .C2(n20575), .A(n20489), .B(n20488), .ZN(
        P1_U3148) );
  AOI22_X1 U23466 ( .A1(n20549), .A2(n20504), .B1(n20548), .B2(n20503), .ZN(
        n20493) );
  AOI22_X1 U23467 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n20507), .B1(
        n20506), .B2(n20491), .ZN(n20492) );
  OAI211_X1 U23468 ( .C1(n20494), .C2(n20575), .A(n20493), .B(n20492), .ZN(
        P1_U3149) );
  AOI22_X1 U23469 ( .A1(n20555), .A2(n20504), .B1(n20554), .B2(n20503), .ZN(
        n20497) );
  AOI22_X1 U23470 ( .A1(P1_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n20507), .B1(
        n20506), .B2(n20495), .ZN(n20496) );
  OAI211_X1 U23471 ( .C1(n20498), .C2(n20575), .A(n20497), .B(n20496), .ZN(
        P1_U3150) );
  AOI22_X1 U23472 ( .A1(n20561), .A2(n20504), .B1(n20560), .B2(n20503), .ZN(
        n20501) );
  AOI22_X1 U23473 ( .A1(P1_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n20507), .B1(
        n20506), .B2(n20499), .ZN(n20500) );
  OAI211_X1 U23474 ( .C1(n20502), .C2(n20575), .A(n20501), .B(n20500), .ZN(
        P1_U3151) );
  AOI22_X1 U23475 ( .A1(n20569), .A2(n20504), .B1(n20567), .B2(n20503), .ZN(
        n20509) );
  AOI22_X1 U23476 ( .A1(P1_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n20507), .B1(
        n20506), .B2(n20505), .ZN(n20508) );
  OAI211_X1 U23477 ( .C1(n20510), .C2(n20575), .A(n20509), .B(n20508), .ZN(
        P1_U3152) );
  INV_X1 U23478 ( .A(n20511), .ZN(n20566) );
  AOI21_X1 U23479 ( .B1(n20513), .B2(n20512), .A(n20566), .ZN(n20520) );
  OAI22_X1 U23480 ( .A1(n20520), .A2(n20518), .B1(n20514), .B2(n12396), .ZN(
        n20568) );
  AOI22_X1 U23481 ( .A1(n20516), .A2(n20568), .B1(n20515), .B2(n20566), .ZN(
        n20528) );
  OAI21_X1 U23482 ( .B1(n20519), .B2(n20518), .A(n20517), .ZN(n20521) );
  NAND2_X1 U23483 ( .A1(n20521), .A2(n20520), .ZN(n20522) );
  OAI211_X1 U23484 ( .C1(n20525), .C2(n20524), .A(n20523), .B(n20522), .ZN(
        n20572) );
  AOI22_X1 U23485 ( .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n20572), .B1(
        n20571), .B2(n20526), .ZN(n20527) );
  OAI211_X1 U23486 ( .C1(n20529), .C2(n20575), .A(n20528), .B(n20527), .ZN(
        P1_U3153) );
  AOI22_X1 U23487 ( .A1(n20531), .A2(n20568), .B1(n20530), .B2(n20566), .ZN(
        n20534) );
  AOI22_X1 U23488 ( .A1(P1_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n20572), .B1(
        n20571), .B2(n20532), .ZN(n20533) );
  OAI211_X1 U23489 ( .C1(n20535), .C2(n20575), .A(n20534), .B(n20533), .ZN(
        P1_U3154) );
  AOI22_X1 U23490 ( .A1(n20537), .A2(n20568), .B1(n20536), .B2(n20566), .ZN(
        n20540) );
  AOI22_X1 U23491 ( .A1(P1_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n20572), .B1(
        n20571), .B2(n20538), .ZN(n20539) );
  OAI211_X1 U23492 ( .C1(n20541), .C2(n20575), .A(n20540), .B(n20539), .ZN(
        P1_U3155) );
  AOI22_X1 U23493 ( .A1(n20543), .A2(n20568), .B1(n20542), .B2(n20566), .ZN(
        n20546) );
  AOI22_X1 U23494 ( .A1(P1_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n20572), .B1(
        n20571), .B2(n20544), .ZN(n20545) );
  OAI211_X1 U23495 ( .C1(n20547), .C2(n20575), .A(n20546), .B(n20545), .ZN(
        P1_U3156) );
  AOI22_X1 U23496 ( .A1(n20549), .A2(n20568), .B1(n20548), .B2(n20566), .ZN(
        n20552) );
  AOI22_X1 U23497 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n20572), .B1(
        n20571), .B2(n20550), .ZN(n20551) );
  OAI211_X1 U23498 ( .C1(n20553), .C2(n20575), .A(n20552), .B(n20551), .ZN(
        P1_U3157) );
  AOI22_X1 U23499 ( .A1(n20555), .A2(n20568), .B1(n20554), .B2(n20566), .ZN(
        n20558) );
  AOI22_X1 U23500 ( .A1(P1_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n20572), .B1(
        n20571), .B2(n20556), .ZN(n20557) );
  OAI211_X1 U23501 ( .C1(n20559), .C2(n20575), .A(n20558), .B(n20557), .ZN(
        P1_U3158) );
  AOI22_X1 U23502 ( .A1(n20561), .A2(n20568), .B1(n20560), .B2(n20566), .ZN(
        n20564) );
  AOI22_X1 U23503 ( .A1(P1_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n20572), .B1(
        n20571), .B2(n20562), .ZN(n20563) );
  OAI211_X1 U23504 ( .C1(n20565), .C2(n20575), .A(n20564), .B(n20563), .ZN(
        P1_U3159) );
  AOI22_X1 U23505 ( .A1(n20569), .A2(n20568), .B1(n20567), .B2(n20566), .ZN(
        n20574) );
  AOI22_X1 U23506 ( .A1(P1_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n20572), .B1(
        n20571), .B2(n20570), .ZN(n20573) );
  OAI211_X1 U23507 ( .C1(n20576), .C2(n20575), .A(n20574), .B(n20573), .ZN(
        P1_U3160) );
  AOI21_X1 U23508 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n15822), .A(n20577), 
        .ZN(n20579) );
  NAND2_X1 U23509 ( .A1(n20579), .A2(n20578), .ZN(P1_U3163) );
  AND2_X1 U23510 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n20580), .ZN(
        P1_U3164) );
  AND2_X1 U23511 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n20580), .ZN(
        P1_U3165) );
  AND2_X1 U23512 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n20580), .ZN(
        P1_U3166) );
  AND2_X1 U23513 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n20580), .ZN(
        P1_U3167) );
  AND2_X1 U23514 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n20580), .ZN(
        P1_U3168) );
  AND2_X1 U23515 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n20580), .ZN(
        P1_U3169) );
  AND2_X1 U23516 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n20580), .ZN(
        P1_U3170) );
  AND2_X1 U23517 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n20580), .ZN(
        P1_U3171) );
  AND2_X1 U23518 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n20580), .ZN(
        P1_U3172) );
  AND2_X1 U23519 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n20580), .ZN(
        P1_U3173) );
  AND2_X1 U23520 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n20580), .ZN(
        P1_U3174) );
  AND2_X1 U23521 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n20580), .ZN(
        P1_U3175) );
  AND2_X1 U23522 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n20580), .ZN(
        P1_U3176) );
  AND2_X1 U23523 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n20580), .ZN(
        P1_U3177) );
  AND2_X1 U23524 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n20580), .ZN(
        P1_U3178) );
  AND2_X1 U23525 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n20580), .ZN(
        P1_U3179) );
  AND2_X1 U23526 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n20580), .ZN(
        P1_U3180) );
  AND2_X1 U23527 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n20580), .ZN(
        P1_U3181) );
  AND2_X1 U23528 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n20580), .ZN(
        P1_U3182) );
  AND2_X1 U23529 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n20580), .ZN(
        P1_U3183) );
  AND2_X1 U23530 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(n20580), .ZN(
        P1_U3184) );
  AND2_X1 U23531 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n20580), .ZN(
        P1_U3185) );
  AND2_X1 U23532 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n20580), .ZN(P1_U3186) );
  AND2_X1 U23533 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n20580), .ZN(P1_U3187) );
  AND2_X1 U23534 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n20580), .ZN(P1_U3188) );
  AND2_X1 U23535 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n20580), .ZN(P1_U3189) );
  AND2_X1 U23536 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n20580), .ZN(P1_U3190) );
  AND2_X1 U23537 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n20580), .ZN(P1_U3191) );
  AND2_X1 U23538 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n20580), .ZN(P1_U3192) );
  AND2_X1 U23539 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n20580), .ZN(P1_U3193) );
  AOI21_X1 U23540 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n20590), .A(n20585), 
        .ZN(n20587) );
  NOR2_X1 U23541 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n20582) );
  NOR2_X1 U23542 ( .A1(n20582), .A2(n20581), .ZN(n20584) );
  INV_X1 U23543 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n20583) );
  AOI211_X1 U23544 ( .C1(NA), .C2(n20585), .A(n20584), .B(n20583), .ZN(n20586)
         );
  OAI22_X1 U23545 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20587), .B1(n20675), 
        .B2(n20586), .ZN(P1_U3194) );
  NAND3_X1 U23546 ( .A1(n20590), .A2(P1_STATE_REG_1__SCAN_IN), .A3(n20589), 
        .ZN(n20595) );
  INV_X1 U23547 ( .A(n20587), .ZN(n20588) );
  OAI211_X1 U23548 ( .C1(P1_STATE_REG_1__SCAN_IN), .C2(n20589), .A(
        P1_STATE_REG_2__SCAN_IN), .B(n20588), .ZN(n20594) );
  NAND2_X1 U23549 ( .A1(n20590), .A2(n20589), .ZN(n20591) );
  OAI221_X1 U23550 ( .B1(P1_REQUESTPENDING_REG_SCAN_IN), .B2(
        P1_STATE_REG_1__SCAN_IN), .C1(P1_REQUESTPENDING_REG_SCAN_IN), .C2(
        n20591), .A(n20597), .ZN(n20592) );
  NAND3_X1 U23551 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(HOLD), .A3(n20592), .ZN(
        n20593) );
  OAI211_X1 U23552 ( .C1(n20596), .C2(n20595), .A(n20594), .B(n20593), .ZN(
        P1_U3196) );
  NAND2_X1 U23553 ( .A1(n20675), .A2(n20597), .ZN(n20639) );
  INV_X1 U23554 ( .A(P1_ADDRESS_REG_0__SCAN_IN), .ZN(n20598) );
  NAND2_X1 U23555 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20675), .ZN(n20643) );
  OAI222_X1 U23556 ( .A1(n20639), .A2(n20600), .B1(n20598), .B2(n20675), .C1(
        n12917), .C2(n20643), .ZN(P1_U3197) );
  INV_X1 U23557 ( .A(n20639), .ZN(n20647) );
  AOI22_X1 U23558 ( .A1(P1_ADDRESS_REG_1__SCAN_IN), .A2(n20662), .B1(
        P1_REIP_REG_3__SCAN_IN), .B2(n20647), .ZN(n20599) );
  OAI21_X1 U23559 ( .B1(n20600), .B2(n20643), .A(n20599), .ZN(P1_U3198) );
  INV_X1 U23560 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n20602) );
  OAI222_X1 U23561 ( .A1(n20643), .A2(n20602), .B1(n20601), .B2(n20675), .C1(
        n20604), .C2(n20639), .ZN(P1_U3199) );
  INV_X1 U23562 ( .A(P1_ADDRESS_REG_3__SCAN_IN), .ZN(n20603) );
  OAI222_X1 U23563 ( .A1(n20643), .A2(n20604), .B1(n20603), .B2(n20675), .C1(
        n20606), .C2(n20639), .ZN(P1_U3200) );
  INV_X1 U23564 ( .A(P1_ADDRESS_REG_4__SCAN_IN), .ZN(n20605) );
  OAI222_X1 U23565 ( .A1(n20643), .A2(n20606), .B1(n20605), .B2(n20675), .C1(
        n20730), .C2(n20639), .ZN(P1_U3201) );
  INV_X1 U23566 ( .A(P1_ADDRESS_REG_5__SCAN_IN), .ZN(n20607) );
  OAI222_X1 U23567 ( .A1(n20643), .A2(n20730), .B1(n20607), .B2(n20675), .C1(
        n20609), .C2(n20639), .ZN(P1_U3202) );
  AOI22_X1 U23568 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(n20662), .B1(
        P1_REIP_REG_8__SCAN_IN), .B2(n20647), .ZN(n20608) );
  OAI21_X1 U23569 ( .B1(n20609), .B2(n20643), .A(n20608), .ZN(P1_U3203) );
  INV_X1 U23570 ( .A(n20643), .ZN(n20648) );
  AOI22_X1 U23571 ( .A1(P1_ADDRESS_REG_7__SCAN_IN), .A2(n20662), .B1(
        P1_REIP_REG_8__SCAN_IN), .B2(n20648), .ZN(n20610) );
  OAI21_X1 U23572 ( .B1(n20612), .B2(n20639), .A(n20610), .ZN(P1_U3204) );
  AOI22_X1 U23573 ( .A1(P1_ADDRESS_REG_8__SCAN_IN), .A2(n20662), .B1(
        P1_REIP_REG_10__SCAN_IN), .B2(n20647), .ZN(n20611) );
  OAI21_X1 U23574 ( .B1(n20612), .B2(n20643), .A(n20611), .ZN(P1_U3205) );
  AOI22_X1 U23575 ( .A1(P1_ADDRESS_REG_9__SCAN_IN), .A2(n20662), .B1(
        P1_REIP_REG_10__SCAN_IN), .B2(n20648), .ZN(n20613) );
  OAI21_X1 U23576 ( .B1(n20615), .B2(n20639), .A(n20613), .ZN(P1_U3206) );
  INV_X1 U23577 ( .A(P1_ADDRESS_REG_10__SCAN_IN), .ZN(n20614) );
  OAI222_X1 U23578 ( .A1(n20643), .A2(n20615), .B1(n20614), .B2(n20675), .C1(
        n20617), .C2(n20639), .ZN(P1_U3207) );
  INV_X1 U23579 ( .A(P1_ADDRESS_REG_11__SCAN_IN), .ZN(n20616) );
  OAI222_X1 U23580 ( .A1(n20643), .A2(n20617), .B1(n20616), .B2(n20675), .C1(
        n20619), .C2(n20639), .ZN(P1_U3208) );
  INV_X1 U23581 ( .A(P1_ADDRESS_REG_12__SCAN_IN), .ZN(n20618) );
  OAI222_X1 U23582 ( .A1(n20643), .A2(n20619), .B1(n20618), .B2(n20675), .C1(
        n20824), .C2(n20639), .ZN(P1_U3209) );
  INV_X1 U23583 ( .A(P1_ADDRESS_REG_13__SCAN_IN), .ZN(n20620) );
  OAI222_X1 U23584 ( .A1(n20639), .A2(n20622), .B1(n20620), .B2(n20675), .C1(
        n20824), .C2(n20643), .ZN(P1_U3210) );
  INV_X1 U23585 ( .A(P1_ADDRESS_REG_14__SCAN_IN), .ZN(n20621) );
  OAI222_X1 U23586 ( .A1(n20643), .A2(n20622), .B1(n20621), .B2(n20675), .C1(
        n20624), .C2(n20639), .ZN(P1_U3211) );
  INV_X1 U23587 ( .A(P1_ADDRESS_REG_15__SCAN_IN), .ZN(n20623) );
  OAI222_X1 U23588 ( .A1(n20643), .A2(n20624), .B1(n20623), .B2(n20675), .C1(
        n14333), .C2(n20639), .ZN(P1_U3212) );
  INV_X1 U23589 ( .A(P1_ADDRESS_REG_16__SCAN_IN), .ZN(n20625) );
  OAI222_X1 U23590 ( .A1(n20643), .A2(n14333), .B1(n20625), .B2(n20675), .C1(
        n20627), .C2(n20639), .ZN(P1_U3213) );
  INV_X1 U23591 ( .A(P1_ADDRESS_REG_17__SCAN_IN), .ZN(n20626) );
  OAI222_X1 U23592 ( .A1(n20643), .A2(n20627), .B1(n20626), .B2(n20675), .C1(
        n20629), .C2(n20639), .ZN(P1_U3214) );
  AOI22_X1 U23593 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(n20662), .B1(
        P1_REIP_REG_20__SCAN_IN), .B2(n20647), .ZN(n20628) );
  OAI21_X1 U23594 ( .B1(n20629), .B2(n20643), .A(n20628), .ZN(P1_U3215) );
  AOI22_X1 U23595 ( .A1(P1_ADDRESS_REG_19__SCAN_IN), .A2(n20662), .B1(
        P1_REIP_REG_20__SCAN_IN), .B2(n20648), .ZN(n20630) );
  OAI21_X1 U23596 ( .B1(n20631), .B2(n20639), .A(n20630), .ZN(P1_U3216) );
  INV_X1 U23597 ( .A(P1_ADDRESS_REG_20__SCAN_IN), .ZN(n20759) );
  OAI222_X1 U23598 ( .A1(n20643), .A2(n20631), .B1(n20759), .B2(n20675), .C1(
        n20633), .C2(n20639), .ZN(P1_U3217) );
  INV_X1 U23599 ( .A(P1_ADDRESS_REG_21__SCAN_IN), .ZN(n20911) );
  INV_X1 U23600 ( .A(P1_REIP_REG_23__SCAN_IN), .ZN(n20632) );
  OAI222_X1 U23601 ( .A1(n20643), .A2(n20633), .B1(n20911), .B2(n20675), .C1(
        n20632), .C2(n20639), .ZN(P1_U3218) );
  AOI222_X1 U23602 ( .A1(n20647), .A2(P1_REIP_REG_24__SCAN_IN), .B1(
        P1_ADDRESS_REG_22__SCAN_IN), .B2(n20662), .C1(P1_REIP_REG_23__SCAN_IN), 
        .C2(n20648), .ZN(n20634) );
  INV_X1 U23603 ( .A(n20634), .ZN(P1_U3219) );
  INV_X1 U23604 ( .A(P1_ADDRESS_REG_23__SCAN_IN), .ZN(n20635) );
  OAI222_X1 U23605 ( .A1(n20643), .A2(n20636), .B1(n20635), .B2(n20675), .C1(
        n20637), .C2(n20639), .ZN(P1_U3220) );
  INV_X1 U23606 ( .A(P1_ADDRESS_REG_24__SCAN_IN), .ZN(n20638) );
  OAI222_X1 U23607 ( .A1(n20639), .A2(n20642), .B1(n20638), .B2(n20675), .C1(
        n20637), .C2(n20643), .ZN(P1_U3221) );
  INV_X1 U23608 ( .A(P1_ADDRESS_REG_25__SCAN_IN), .ZN(n20641) );
  OAI222_X1 U23609 ( .A1(n20643), .A2(n20642), .B1(n20641), .B2(n20675), .C1(
        n20640), .C2(n20639), .ZN(P1_U3222) );
  AOI222_X1 U23610 ( .A1(n20648), .A2(P1_REIP_REG_27__SCAN_IN), .B1(
        P1_ADDRESS_REG_26__SCAN_IN), .B2(n20662), .C1(P1_REIP_REG_28__SCAN_IN), 
        .C2(n20647), .ZN(n20644) );
  INV_X1 U23611 ( .A(n20644), .ZN(P1_U3223) );
  AOI222_X1 U23612 ( .A1(n20648), .A2(P1_REIP_REG_28__SCAN_IN), .B1(
        P1_ADDRESS_REG_27__SCAN_IN), .B2(n20662), .C1(P1_REIP_REG_29__SCAN_IN), 
        .C2(n20647), .ZN(n20645) );
  INV_X1 U23613 ( .A(n20645), .ZN(P1_U3224) );
  AOI222_X1 U23614 ( .A1(n20647), .A2(P1_REIP_REG_30__SCAN_IN), .B1(
        P1_ADDRESS_REG_28__SCAN_IN), .B2(n20662), .C1(P1_REIP_REG_29__SCAN_IN), 
        .C2(n20648), .ZN(n20646) );
  INV_X1 U23615 ( .A(n20646), .ZN(P1_U3225) );
  AOI222_X1 U23616 ( .A1(n20648), .A2(P1_REIP_REG_30__SCAN_IN), .B1(
        P1_ADDRESS_REG_29__SCAN_IN), .B2(n20662), .C1(P1_REIP_REG_31__SCAN_IN), 
        .C2(n20647), .ZN(n20649) );
  INV_X1 U23617 ( .A(n20649), .ZN(P1_U3226) );
  MUX2_X1 U23618 ( .A(P1_BE_N_REG_3__SCAN_IN), .B(P1_BYTEENABLE_REG_3__SCAN_IN), .S(n20675), .Z(P1_U3458) );
  MUX2_X1 U23619 ( .A(P1_BE_N_REG_2__SCAN_IN), .B(P1_BYTEENABLE_REG_2__SCAN_IN), .S(n20675), .Z(P1_U3459) );
  MUX2_X1 U23620 ( .A(P1_BE_N_REG_1__SCAN_IN), .B(P1_BYTEENABLE_REG_1__SCAN_IN), .S(n20675), .Z(P1_U3460) );
  OAI22_X1 U23621 ( .A1(n20662), .A2(P1_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P1_BE_N_REG_0__SCAN_IN), .B2(n20675), .ZN(n20650) );
  INV_X1 U23622 ( .A(n20650), .ZN(P1_U3461) );
  OAI21_X1 U23623 ( .B1(P1_DATAWIDTH_REG_0__SCAN_IN), .B2(n20654), .A(n20652), 
        .ZN(n20651) );
  INV_X1 U23624 ( .A(n20651), .ZN(P1_U3464) );
  INV_X1 U23625 ( .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20653) );
  OAI21_X1 U23626 ( .B1(n20654), .B2(n20653), .A(n20652), .ZN(P1_U3465) );
  NOR2_X1 U23627 ( .A1(P1_DATAWIDTH_REG_1__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(n20655) );
  AOI21_X1 U23628 ( .B1(P1_DATAWIDTH_REG_0__SCAN_IN), .B2(n12475), .A(n20655), 
        .ZN(n20658) );
  OAI211_X1 U23629 ( .C1(n20659), .C2(P1_BYTEENABLE_REG_2__SCAN_IN), .A(n20656), .B(n20660), .ZN(n20657) );
  OAI21_X1 U23630 ( .B1(n20658), .B2(n20660), .A(n20657), .ZN(P1_U3481) );
  OAI22_X1 U23631 ( .A1(n20660), .A2(P1_REIP_REG_0__SCAN_IN), .B1(n20659), 
        .B2(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n20661) );
  INV_X1 U23632 ( .A(n20661), .ZN(P1_U3482) );
  AOI22_X1 U23633 ( .A1(n20675), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n20663), 
        .B2(n20662), .ZN(P1_U3483) );
  AOI211_X1 U23634 ( .C1(n20667), .C2(n20666), .A(n20665), .B(n20664), .ZN(
        n20674) );
  OAI211_X1 U23635 ( .C1(P1_STATEBS16_REG_SCAN_IN), .C2(n20669), .A(n20668), 
        .B(P1_STATE2_REG_2__SCAN_IN), .ZN(n20671) );
  AOI21_X1 U23636 ( .B1(P1_STATE2_REG_0__SCAN_IN), .B2(n20671), .A(n20670), 
        .ZN(n20673) );
  NAND2_X1 U23637 ( .A1(n20674), .A2(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n20672) );
  OAI21_X1 U23638 ( .B1(n20674), .B2(n20673), .A(n20672), .ZN(P1_U3485) );
  MUX2_X1 U23639 ( .A(P1_M_IO_N_REG_SCAN_IN), .B(P1_MEMORYFETCH_REG_SCAN_IN), 
        .S(n20675), .Z(P1_U3486) );
  AOI22_X1 U23640 ( .A1(n20677), .A2(P3_ADDRESS_REG_29__SCAN_IN), .B1(
        P2_ADDRESS_REG_29__SCAN_IN), .B2(n20676), .ZN(n20983) );
  NOR4_X1 U23641 ( .A1(P2_ADDRESS_REG_6__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(P2_M_IO_N_REG_SCAN_IN), .A4(
        P2_W_R_N_REG_SCAN_IN), .ZN(n20686) );
  NOR4_X1 U23642 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(
        P3_INSTQUEUE_REG_14__6__SCAN_IN), .A3(P3_ADDRESS_REG_9__SCAN_IN), .A4(
        P3_ADDRESS_REG_3__SCAN_IN), .ZN(n20678) );
  NAND3_X1 U23643 ( .A1(n20678), .A2(n20821), .A3(n20755), .ZN(n20684) );
  NOR4_X1 U23644 ( .A1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(
        P2_EAX_REG_11__SCAN_IN), .A3(P2_MORE_REG_SCAN_IN), .A4(
        P2_UWORD_REG_8__SCAN_IN), .ZN(n20682) );
  NOR4_X1 U23645 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_UWORD_REG_5__SCAN_IN), 
        .A3(P1_UWORD_REG_10__SCAN_IN), .A4(P1_DATAO_REG_19__SCAN_IN), .ZN(
        n20681) );
  NOR4_X1 U23646 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(
        P3_INSTQUEUE_REG_3__4__SCAN_IN), .A3(P3_INSTQUEUE_REG_1__2__SCAN_IN), 
        .A4(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n20680) );
  NOR4_X1 U23647 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(
        P3_EAX_REG_12__SCAN_IN), .A3(P3_EAX_REG_8__SCAN_IN), .A4(
        P3_DATAO_REG_22__SCAN_IN), .ZN(n20679) );
  NAND4_X1 U23648 ( .A1(n20682), .A2(n20681), .A3(n20680), .A4(n20679), .ZN(
        n20683) );
  NOR4_X1 U23649 ( .A1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_6__SCAN_IN), .A3(n20684), .A4(n20683), .ZN(n20685) );
  NAND4_X1 U23650 ( .A1(n20688), .A2(n20687), .A3(n20686), .A4(n20685), .ZN(
        n20720) );
  NOR4_X1 U23651 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(
        P1_INSTQUEUE_REG_10__4__SCAN_IN), .A3(P1_INSTQUEUE_REG_6__2__SCAN_IN), 
        .A4(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n20692) );
  NOR4_X1 U23652 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_13__5__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A4(P1_REIP_REG_6__SCAN_IN), .ZN(
        n20691) );
  NOR4_X1 U23653 ( .A1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P1_EBX_REG_29__SCAN_IN), .A3(P1_EBX_REG_21__SCAN_IN), .A4(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n20690) );
  NOR4_X1 U23654 ( .A1(P1_INSTQUEUE_REG_0__6__SCAN_IN), .A2(
        P1_REIP_REG_14__SCAN_IN), .A3(DATAI_27_), .A4(BUF1_REG_18__SCAN_IN), 
        .ZN(n20689) );
  NAND4_X1 U23655 ( .A1(n20692), .A2(n20691), .A3(n20690), .A4(n20689), .ZN(
        n20719) );
  NOR4_X1 U23656 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A3(P3_EBX_REG_10__SCAN_IN), .A4(
        P2_DATAO_REG_19__SCAN_IN), .ZN(n20696) );
  NOR4_X1 U23657 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(
        P3_INSTQUEUE_REG_13__6__SCAN_IN), .A3(P3_EBX_REG_31__SCAN_IN), .A4(
        P3_REIP_REG_2__SCAN_IN), .ZN(n20695) );
  NOR4_X1 U23658 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(
        P2_REIP_REG_26__SCAN_IN), .A3(BUF1_REG_25__SCAN_IN), .A4(
        BUF2_REG_25__SCAN_IN), .ZN(n20694) );
  NOR4_X1 U23659 ( .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A3(P2_REIP_REG_19__SCAN_IN), .A4(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n20693) );
  NAND4_X1 U23660 ( .A1(n20696), .A2(n20695), .A3(n20694), .A4(n20693), .ZN(
        n20718) );
  NAND4_X1 U23661 ( .A1(P1_INSTQUEUE_REG_12__5__SCAN_IN), .A2(
        P1_EAX_REG_23__SCAN_IN), .A3(P1_REIP_REG_17__SCAN_IN), .A4(
        P1_LWORD_REG_12__SCAN_IN), .ZN(n20700) );
  NAND4_X1 U23662 ( .A1(P2_REIP_REG_20__SCAN_IN), .A2(P1_CODEFETCH_REG_SCAN_IN), .A3(P3_DATAWIDTH_REG_15__SCAN_IN), .A4(P3_ADDRESS_REG_23__SCAN_IN), .ZN(
        n20699) );
  NAND4_X1 U23663 ( .A1(P1_EBX_REG_2__SCAN_IN), .A2(BUF1_REG_23__SCAN_IN), 
        .A3(P1_DATAO_REG_5__SCAN_IN), .A4(P3_LWORD_REG_8__SCAN_IN), .ZN(n20698) );
  NAND4_X1 U23664 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(
        P2_EAX_REG_23__SCAN_IN), .A3(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A4(
        P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n20697) );
  NOR4_X1 U23665 ( .A1(n20700), .A2(n20699), .A3(n20698), .A4(n20697), .ZN(
        n20716) );
  NAND4_X1 U23666 ( .A1(P1_INSTQUEUE_REG_4__2__SCAN_IN), .A2(
        P2_DATAO_REG_1__SCAN_IN), .A3(P1_LWORD_REG_14__SCAN_IN), .A4(
        P1_DATAO_REG_1__SCAN_IN), .ZN(n20704) );
  NAND4_X1 U23667 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(
        P2_ADDRESS_REG_10__SCAN_IN), .A3(P1_INSTADDRPOINTER_REG_2__SCAN_IN), 
        .A4(P3_DATAO_REG_30__SCAN_IN), .ZN(n20703) );
  NAND4_X1 U23668 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(
        BUF2_REG_20__SCAN_IN), .A3(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A4(
        P1_LWORD_REG_7__SCAN_IN), .ZN(n20702) );
  NAND4_X1 U23669 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(
        P1_ADDRESS_REG_20__SCAN_IN), .A3(BUF1_REG_8__SCAN_IN), .A4(
        P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n20701) );
  NOR4_X1 U23670 ( .A1(n20704), .A2(n20703), .A3(n20702), .A4(n20701), .ZN(
        n20715) );
  NAND4_X1 U23671 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(
        P1_EAX_REG_18__SCAN_IN), .A3(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A4(
        P3_REIP_REG_25__SCAN_IN), .ZN(n20708) );
  NAND4_X1 U23672 ( .A1(P1_INSTQUEUE_REG_15__2__SCAN_IN), .A2(
        P3_EAX_REG_26__SCAN_IN), .A3(P2_UWORD_REG_5__SCAN_IN), .A4(
        P3_DATAO_REG_19__SCAN_IN), .ZN(n20707) );
  NAND4_X1 U23673 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_3__2__SCAN_IN), .A3(P2_UWORD_REG_4__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20706) );
  NAND4_X1 U23674 ( .A1(P2_REIP_REG_13__SCAN_IN), .A2(DATAI_14_), .A3(
        P3_INSTQUEUE_REG_12__5__SCAN_IN), .A4(P3_ADDRESS_REG_8__SCAN_IN), .ZN(
        n20705) );
  NOR4_X1 U23675 ( .A1(n20708), .A2(n20707), .A3(n20706), .A4(n20705), .ZN(
        n20714) );
  NAND4_X1 U23676 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_24__SCAN_IN), .A3(
        P3_INSTQUEUE_REG_12__2__SCAN_IN), .A4(P2_LWORD_REG_10__SCAN_IN), .ZN(
        n20712) );
  NAND4_X1 U23677 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_1__3__SCAN_IN), .A3(P3_INSTQUEUE_REG_5__5__SCAN_IN), 
        .A4(P3_BE_N_REG_2__SCAN_IN), .ZN(n20711) );
  NAND4_X1 U23678 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_23__SCAN_IN), .A3(P1_ADDRESS_REG_21__SCAN_IN), 
        .A4(P3_EAX_REG_7__SCAN_IN), .ZN(n20710) );
  NAND4_X1 U23679 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(
        P2_REIP_REG_7__SCAN_IN), .A3(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A4(
        P3_DATAO_REG_11__SCAN_IN), .ZN(n20709) );
  NOR4_X1 U23680 ( .A1(n20712), .A2(n20711), .A3(n20710), .A4(n20709), .ZN(
        n20713) );
  NAND4_X1 U23681 ( .A1(n20716), .A2(n20715), .A3(n20714), .A4(n20713), .ZN(
        n20717) );
  NOR4_X1 U23682 ( .A1(n20720), .A2(n20719), .A3(n20718), .A4(n20717), .ZN(
        n20981) );
  AOI22_X1 U23683 ( .A1(n20723), .A2(keyinput127), .B1(n20722), .B2(
        keyinput126), .ZN(n20721) );
  OAI221_X1 U23684 ( .B1(n20723), .B2(keyinput127), .C1(n20722), .C2(
        keyinput126), .A(n20721), .ZN(n20727) );
  XNOR2_X1 U23685 ( .A(n20724), .B(keyinput105), .ZN(n20726) );
  XOR2_X1 U23686 ( .A(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B(keyinput29), .Z(
        n20725) );
  OR3_X1 U23687 ( .A1(n20727), .A2(n20726), .A3(n20725), .ZN(n20736) );
  AOI22_X1 U23688 ( .A1(n20730), .A2(keyinput94), .B1(n20729), .B2(keyinput51), 
        .ZN(n20728) );
  OAI221_X1 U23689 ( .B1(n20730), .B2(keyinput94), .C1(n20729), .C2(keyinput51), .A(n20728), .ZN(n20735) );
  AOI22_X1 U23690 ( .A1(n20733), .A2(keyinput74), .B1(n20732), .B2(keyinput33), 
        .ZN(n20731) );
  OAI221_X1 U23691 ( .B1(n20733), .B2(keyinput74), .C1(n20732), .C2(keyinput33), .A(n20731), .ZN(n20734) );
  NOR3_X1 U23692 ( .A1(n20736), .A2(n20735), .A3(n20734), .ZN(n20786) );
  AOI22_X1 U23693 ( .A1(n20739), .A2(keyinput89), .B1(keyinput2), .B2(n20738), 
        .ZN(n20737) );
  OAI221_X1 U23694 ( .B1(n20739), .B2(keyinput89), .C1(n20738), .C2(keyinput2), 
        .A(n20737), .ZN(n20752) );
  INV_X1 U23695 ( .A(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n20742) );
  AOI22_X1 U23696 ( .A1(n20742), .A2(keyinput70), .B1(keyinput86), .B2(n20741), 
        .ZN(n20740) );
  OAI221_X1 U23697 ( .B1(n20742), .B2(keyinput70), .C1(n20741), .C2(keyinput86), .A(n20740), .ZN(n20751) );
  INV_X1 U23698 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n20744) );
  AOI22_X1 U23699 ( .A1(n20745), .A2(keyinput42), .B1(keyinput92), .B2(n20744), 
        .ZN(n20743) );
  OAI221_X1 U23700 ( .B1(n20745), .B2(keyinput42), .C1(n20744), .C2(keyinput92), .A(n20743), .ZN(n20750) );
  INV_X1 U23701 ( .A(DATAI_27_), .ZN(n20748) );
  AOI22_X1 U23702 ( .A1(n20748), .A2(keyinput83), .B1(keyinput69), .B2(n20747), 
        .ZN(n20746) );
  OAI221_X1 U23703 ( .B1(n20748), .B2(keyinput83), .C1(n20747), .C2(keyinput69), .A(n20746), .ZN(n20749) );
  NOR4_X1 U23704 ( .A1(n20752), .A2(n20751), .A3(n20750), .A4(n20749), .ZN(
        n20785) );
  AOI22_X1 U23705 ( .A1(n20755), .A2(keyinput16), .B1(keyinput117), .B2(n20754), .ZN(n20753) );
  OAI221_X1 U23706 ( .B1(n20755), .B2(keyinput16), .C1(n20754), .C2(
        keyinput117), .A(n20753), .ZN(n20767) );
  AOI22_X1 U23707 ( .A1(n20757), .A2(keyinput26), .B1(keyinput72), .B2(n11896), 
        .ZN(n20756) );
  OAI221_X1 U23708 ( .B1(n20757), .B2(keyinput26), .C1(n11896), .C2(keyinput72), .A(n20756), .ZN(n20766) );
  INV_X1 U23709 ( .A(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n20760) );
  AOI22_X1 U23710 ( .A1(n20760), .A2(keyinput100), .B1(keyinput24), .B2(n20759), .ZN(n20758) );
  OAI221_X1 U23711 ( .B1(n20760), .B2(keyinput100), .C1(n20759), .C2(
        keyinput24), .A(n20758), .ZN(n20765) );
  INV_X1 U23712 ( .A(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n20763) );
  INV_X1 U23713 ( .A(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n20762) );
  AOI22_X1 U23714 ( .A1(n20763), .A2(keyinput96), .B1(n20762), .B2(keyinput67), 
        .ZN(n20761) );
  OAI221_X1 U23715 ( .B1(n20763), .B2(keyinput96), .C1(n20762), .C2(keyinput67), .A(n20761), .ZN(n20764) );
  NOR4_X1 U23716 ( .A1(n20767), .A2(n20766), .A3(n20765), .A4(n20764), .ZN(
        n20784) );
  INV_X1 U23717 ( .A(P1_LWORD_REG_7__SCAN_IN), .ZN(n20769) );
  AOI22_X1 U23718 ( .A1(n20770), .A2(keyinput22), .B1(keyinput61), .B2(n20769), 
        .ZN(n20768) );
  OAI221_X1 U23719 ( .B1(n20770), .B2(keyinput22), .C1(n20769), .C2(keyinput61), .A(n20768), .ZN(n20782) );
  AOI22_X1 U23720 ( .A1(n20772), .A2(keyinput80), .B1(n12917), .B2(keyinput13), 
        .ZN(n20771) );
  OAI221_X1 U23721 ( .B1(n20772), .B2(keyinput80), .C1(n12917), .C2(keyinput13), .A(n20771), .ZN(n20781) );
  AOI22_X1 U23722 ( .A1(n20775), .A2(keyinput64), .B1(keyinput125), .B2(n20774), .ZN(n20773) );
  OAI221_X1 U23723 ( .B1(n20775), .B2(keyinput64), .C1(n20774), .C2(
        keyinput125), .A(n20773), .ZN(n20780) );
  AOI22_X1 U23724 ( .A1(n20778), .A2(keyinput37), .B1(n20777), .B2(keyinput112), .ZN(n20776) );
  OAI221_X1 U23725 ( .B1(n20778), .B2(keyinput37), .C1(n20777), .C2(
        keyinput112), .A(n20776), .ZN(n20779) );
  NOR4_X1 U23726 ( .A1(n20782), .A2(n20781), .A3(n20780), .A4(n20779), .ZN(
        n20783) );
  NAND4_X1 U23727 ( .A1(n20786), .A2(n20785), .A3(n20784), .A4(n20783), .ZN(
        n20979) );
  INV_X1 U23728 ( .A(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n20788) );
  AOI22_X1 U23729 ( .A1(n20788), .A2(keyinput79), .B1(n11207), .B2(keyinput59), 
        .ZN(n20787) );
  OAI221_X1 U23730 ( .B1(n20788), .B2(keyinput79), .C1(n11207), .C2(keyinput59), .A(n20787), .ZN(n20792) );
  XOR2_X1 U23731 ( .A(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B(keyinput71), .Z(
        n20791) );
  XNOR2_X1 U23732 ( .A(n20789), .B(keyinput84), .ZN(n20790) );
  OR3_X1 U23733 ( .A1(n20792), .A2(n20791), .A3(n20790), .ZN(n20801) );
  INV_X1 U23734 ( .A(P3_EBX_REG_31__SCAN_IN), .ZN(n20794) );
  AOI22_X1 U23735 ( .A1(n20795), .A2(keyinput57), .B1(keyinput120), .B2(n20794), .ZN(n20793) );
  OAI221_X1 U23736 ( .B1(n20795), .B2(keyinput57), .C1(n20794), .C2(
        keyinput120), .A(n20793), .ZN(n20800) );
  AOI22_X1 U23737 ( .A1(n20798), .A2(keyinput87), .B1(keyinput102), .B2(n20797), .ZN(n20796) );
  OAI221_X1 U23738 ( .B1(n20798), .B2(keyinput87), .C1(n20797), .C2(
        keyinput102), .A(n20796), .ZN(n20799) );
  NOR3_X1 U23739 ( .A1(n20801), .A2(n20800), .A3(n20799), .ZN(n20849) );
  AOI22_X1 U23740 ( .A1(n20804), .A2(keyinput54), .B1(keyinput48), .B2(n20803), 
        .ZN(n20802) );
  OAI221_X1 U23741 ( .B1(n20804), .B2(keyinput54), .C1(n20803), .C2(keyinput48), .A(n20802), .ZN(n20816) );
  INV_X1 U23742 ( .A(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n20806) );
  AOI22_X1 U23743 ( .A1(n10050), .A2(keyinput31), .B1(keyinput90), .B2(n20806), 
        .ZN(n20805) );
  OAI221_X1 U23744 ( .B1(n10050), .B2(keyinput31), .C1(n20806), .C2(keyinput90), .A(n20805), .ZN(n20815) );
  AOI22_X1 U23745 ( .A1(n20809), .A2(keyinput81), .B1(keyinput23), .B2(n20808), 
        .ZN(n20807) );
  OAI221_X1 U23746 ( .B1(n20809), .B2(keyinput81), .C1(n20808), .C2(keyinput23), .A(n20807), .ZN(n20814) );
  INV_X1 U23747 ( .A(P1_CODEFETCH_REG_SCAN_IN), .ZN(n20811) );
  AOI22_X1 U23748 ( .A1(n20812), .A2(keyinput114), .B1(keyinput76), .B2(n20811), .ZN(n20810) );
  OAI221_X1 U23749 ( .B1(n20812), .B2(keyinput114), .C1(n20811), .C2(
        keyinput76), .A(n20810), .ZN(n20813) );
  NOR4_X1 U23750 ( .A1(n20816), .A2(n20815), .A3(n20814), .A4(n20813), .ZN(
        n20848) );
  AOI22_X1 U23751 ( .A1(n20819), .A2(keyinput113), .B1(n20818), .B2(keyinput5), 
        .ZN(n20817) );
  OAI221_X1 U23752 ( .B1(n20819), .B2(keyinput113), .C1(n20818), .C2(keyinput5), .A(n20817), .ZN(n20830) );
  INV_X1 U23753 ( .A(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n20822) );
  AOI22_X1 U23754 ( .A1(n20822), .A2(keyinput44), .B1(keyinput45), .B2(n20821), 
        .ZN(n20820) );
  OAI221_X1 U23755 ( .B1(n20822), .B2(keyinput44), .C1(n20821), .C2(keyinput45), .A(n20820), .ZN(n20829) );
  AOI22_X1 U23756 ( .A1(n20824), .A2(keyinput73), .B1(n11628), .B2(keyinput17), 
        .ZN(n20823) );
  OAI221_X1 U23757 ( .B1(n20824), .B2(keyinput73), .C1(n11628), .C2(keyinput17), .A(n20823), .ZN(n20828) );
  AOI22_X1 U23758 ( .A1(n14333), .A2(keyinput34), .B1(keyinput118), .B2(n20826), .ZN(n20825) );
  OAI221_X1 U23759 ( .B1(n14333), .B2(keyinput34), .C1(n20826), .C2(
        keyinput118), .A(n20825), .ZN(n20827) );
  NOR4_X1 U23760 ( .A1(n20830), .A2(n20829), .A3(n20828), .A4(n20827), .ZN(
        n20847) );
  AOI22_X1 U23761 ( .A1(n20833), .A2(keyinput9), .B1(n20832), .B2(keyinput108), 
        .ZN(n20831) );
  OAI221_X1 U23762 ( .B1(n20833), .B2(keyinput9), .C1(n20832), .C2(keyinput108), .A(n20831), .ZN(n20845) );
  AOI22_X1 U23763 ( .A1(n20836), .A2(keyinput98), .B1(n20835), .B2(keyinput62), 
        .ZN(n20834) );
  OAI221_X1 U23764 ( .B1(n20836), .B2(keyinput98), .C1(n20835), .C2(keyinput62), .A(n20834), .ZN(n20844) );
  INV_X1 U23765 ( .A(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n20838) );
  AOI22_X1 U23766 ( .A1(n11174), .A2(keyinput77), .B1(keyinput82), .B2(n20838), 
        .ZN(n20837) );
  OAI221_X1 U23767 ( .B1(n11174), .B2(keyinput77), .C1(n20838), .C2(keyinput82), .A(n20837), .ZN(n20843) );
  INV_X1 U23768 ( .A(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n20840) );
  AOI22_X1 U23769 ( .A1(n20841), .A2(keyinput97), .B1(keyinput58), .B2(n20840), 
        .ZN(n20839) );
  OAI221_X1 U23770 ( .B1(n20841), .B2(keyinput97), .C1(n20840), .C2(keyinput58), .A(n20839), .ZN(n20842) );
  NOR4_X1 U23771 ( .A1(n20845), .A2(n20844), .A3(n20843), .A4(n20842), .ZN(
        n20846) );
  NAND4_X1 U23772 ( .A1(n20849), .A2(n20848), .A3(n20847), .A4(n20846), .ZN(
        n20978) );
  INV_X1 U23773 ( .A(P1_UWORD_REG_5__SCAN_IN), .ZN(n20852) );
  AOI22_X1 U23774 ( .A1(n20852), .A2(keyinput21), .B1(n20851), .B2(keyinput106), .ZN(n20850) );
  OAI221_X1 U23775 ( .B1(n20852), .B2(keyinput21), .C1(n20851), .C2(
        keyinput106), .A(n20850), .ZN(n20864) );
  AOI22_X1 U23776 ( .A1(n20854), .A2(keyinput68), .B1(n14151), .B2(keyinput91), 
        .ZN(n20853) );
  OAI221_X1 U23777 ( .B1(n20854), .B2(keyinput68), .C1(n14151), .C2(keyinput91), .A(n20853), .ZN(n20863) );
  AOI22_X1 U23778 ( .A1(n20857), .A2(keyinput103), .B1(keyinput66), .B2(n20856), .ZN(n20855) );
  OAI221_X1 U23779 ( .B1(n20857), .B2(keyinput103), .C1(n20856), .C2(
        keyinput66), .A(n20855), .ZN(n20862) );
  INV_X1 U23780 ( .A(P3_LWORD_REG_8__SCAN_IN), .ZN(n20860) );
  AOI22_X1 U23781 ( .A1(n20860), .A2(keyinput8), .B1(n20859), .B2(keyinput0), 
        .ZN(n20858) );
  OAI221_X1 U23782 ( .B1(n20860), .B2(keyinput8), .C1(n20859), .C2(keyinput0), 
        .A(n20858), .ZN(n20861) );
  NOR4_X1 U23783 ( .A1(n20864), .A2(n20863), .A3(n20862), .A4(n20861), .ZN(
        n20909) );
  INV_X1 U23784 ( .A(P1_UWORD_REG_10__SCAN_IN), .ZN(n20866) );
  AOI22_X1 U23785 ( .A1(n20867), .A2(keyinput35), .B1(keyinput107), .B2(n20866), .ZN(n20865) );
  OAI221_X1 U23786 ( .B1(n20867), .B2(keyinput35), .C1(n20866), .C2(
        keyinput107), .A(n20865), .ZN(n20878) );
  AOI22_X1 U23787 ( .A1(n20870), .A2(keyinput4), .B1(n20869), .B2(keyinput7), 
        .ZN(n20868) );
  OAI221_X1 U23788 ( .B1(n20870), .B2(keyinput4), .C1(n20869), .C2(keyinput7), 
        .A(n20868), .ZN(n20877) );
  AOI22_X1 U23789 ( .A1(n20872), .A2(keyinput28), .B1(n11179), .B2(keyinput10), 
        .ZN(n20871) );
  OAI221_X1 U23790 ( .B1(n20872), .B2(keyinput28), .C1(n11179), .C2(keyinput10), .A(n20871), .ZN(n20876) );
  INV_X1 U23791 ( .A(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n20874) );
  AOI22_X1 U23792 ( .A1(n20874), .A2(keyinput95), .B1(n14174), .B2(keyinput47), 
        .ZN(n20873) );
  OAI221_X1 U23793 ( .B1(n20874), .B2(keyinput95), .C1(n14174), .C2(keyinput47), .A(n20873), .ZN(n20875) );
  NOR4_X1 U23794 ( .A1(n20878), .A2(n20877), .A3(n20876), .A4(n20875), .ZN(
        n20908) );
  AOI22_X1 U23795 ( .A1(n20881), .A2(keyinput46), .B1(keyinput39), .B2(n20880), 
        .ZN(n20879) );
  OAI221_X1 U23796 ( .B1(n20881), .B2(keyinput46), .C1(n20880), .C2(keyinput39), .A(n20879), .ZN(n20892) );
  INV_X1 U23797 ( .A(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n20883) );
  AOI22_X1 U23798 ( .A1(n20884), .A2(keyinput123), .B1(keyinput27), .B2(n20883), .ZN(n20882) );
  OAI221_X1 U23799 ( .B1(n20884), .B2(keyinput123), .C1(n20883), .C2(
        keyinput27), .A(n20882), .ZN(n20891) );
  INV_X1 U23800 ( .A(P2_LWORD_REG_10__SCAN_IN), .ZN(n20886) );
  AOI22_X1 U23801 ( .A1(n20886), .A2(keyinput1), .B1(n13758), .B2(keyinput11), 
        .ZN(n20885) );
  OAI221_X1 U23802 ( .B1(n20886), .B2(keyinput1), .C1(n13758), .C2(keyinput11), 
        .A(n20885), .ZN(n20890) );
  INV_X1 U23803 ( .A(P3_DATAO_REG_11__SCAN_IN), .ZN(n20888) );
  AOI22_X1 U23804 ( .A1(n11570), .A2(keyinput41), .B1(keyinput25), .B2(n20888), 
        .ZN(n20887) );
  OAI221_X1 U23805 ( .B1(n11570), .B2(keyinput41), .C1(n20888), .C2(keyinput25), .A(n20887), .ZN(n20889) );
  NOR4_X1 U23806 ( .A1(n20892), .A2(n20891), .A3(n20890), .A4(n20889), .ZN(
        n20907) );
  AOI22_X1 U23807 ( .A1(n20894), .A2(keyinput50), .B1(n11283), .B2(keyinput43), 
        .ZN(n20893) );
  OAI221_X1 U23808 ( .B1(n20894), .B2(keyinput50), .C1(n11283), .C2(keyinput43), .A(n20893), .ZN(n20905) );
  AOI22_X1 U23809 ( .A1(n20896), .A2(keyinput32), .B1(n11625), .B2(keyinput124), .ZN(n20895) );
  OAI221_X1 U23810 ( .B1(n20896), .B2(keyinput32), .C1(n11625), .C2(
        keyinput124), .A(n20895), .ZN(n20904) );
  AOI22_X1 U23811 ( .A1(n20898), .A2(keyinput99), .B1(keyinput122), .B2(n13046), .ZN(n20897) );
  OAI221_X1 U23812 ( .B1(n20898), .B2(keyinput99), .C1(n13046), .C2(
        keyinput122), .A(n20897), .ZN(n20903) );
  INV_X1 U23813 ( .A(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n20900) );
  AOI22_X1 U23814 ( .A1(n20901), .A2(keyinput6), .B1(keyinput119), .B2(n20900), 
        .ZN(n20899) );
  OAI221_X1 U23815 ( .B1(n20901), .B2(keyinput6), .C1(n20900), .C2(keyinput119), .A(n20899), .ZN(n20902) );
  NOR4_X1 U23816 ( .A1(n20905), .A2(n20904), .A3(n20903), .A4(n20902), .ZN(
        n20906) );
  NAND4_X1 U23817 ( .A1(n20909), .A2(n20908), .A3(n20907), .A4(n20906), .ZN(
        n20977) );
  AOI22_X1 U23818 ( .A1(n20912), .A2(keyinput15), .B1(n20911), .B2(keyinput18), 
        .ZN(n20910) );
  OAI221_X1 U23819 ( .B1(n20912), .B2(keyinput15), .C1(n20911), .C2(keyinput18), .A(n20910), .ZN(n20925) );
  INV_X1 U23820 ( .A(P2_UWORD_REG_5__SCAN_IN), .ZN(n20914) );
  AOI22_X1 U23821 ( .A1(n20915), .A2(keyinput56), .B1(n20914), .B2(keyinput60), 
        .ZN(n20913) );
  OAI221_X1 U23822 ( .B1(n20915), .B2(keyinput56), .C1(n20914), .C2(keyinput60), .A(n20913), .ZN(n20924) );
  INV_X1 U23823 ( .A(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n20917) );
  AOI22_X1 U23824 ( .A1(n20918), .A2(keyinput115), .B1(n20917), .B2(keyinput53), .ZN(n20916) );
  OAI221_X1 U23825 ( .B1(n20918), .B2(keyinput115), .C1(n20917), .C2(
        keyinput53), .A(n20916), .ZN(n20923) );
  INV_X1 U23826 ( .A(P3_DATAO_REG_19__SCAN_IN), .ZN(n20921) );
  INV_X1 U23827 ( .A(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n20920) );
  AOI22_X1 U23828 ( .A1(n20921), .A2(keyinput20), .B1(n20920), .B2(keyinput49), 
        .ZN(n20919) );
  OAI221_X1 U23829 ( .B1(n20921), .B2(keyinput20), .C1(n20920), .C2(keyinput49), .A(n20919), .ZN(n20922) );
  NOR4_X1 U23830 ( .A1(n20925), .A2(n20924), .A3(n20923), .A4(n20922), .ZN(
        n20975) );
  AOI22_X1 U23831 ( .A1(n20928), .A2(keyinput121), .B1(n20927), .B2(keyinput52), .ZN(n20926) );
  OAI221_X1 U23832 ( .B1(n20928), .B2(keyinput121), .C1(n20927), .C2(
        keyinput52), .A(n20926), .ZN(n20940) );
  AOI22_X1 U23833 ( .A1(n20931), .A2(keyinput111), .B1(keyinput88), .B2(n20930), .ZN(n20929) );
  OAI221_X1 U23834 ( .B1(n20931), .B2(keyinput111), .C1(n20930), .C2(
        keyinput88), .A(n20929), .ZN(n20939) );
  AOI22_X1 U23835 ( .A1(n20934), .A2(keyinput75), .B1(keyinput110), .B2(n20933), .ZN(n20932) );
  OAI221_X1 U23836 ( .B1(n20934), .B2(keyinput75), .C1(n20933), .C2(
        keyinput110), .A(n20932), .ZN(n20938) );
  AOI22_X1 U23837 ( .A1(n20936), .A2(keyinput19), .B1(n11215), .B2(keyinput63), 
        .ZN(n20935) );
  OAI221_X1 U23838 ( .B1(n20936), .B2(keyinput19), .C1(n11215), .C2(keyinput63), .A(n20935), .ZN(n20937) );
  NOR4_X1 U23839 ( .A1(n20940), .A2(n20939), .A3(n20938), .A4(n20937), .ZN(
        n20974) );
  AOI22_X1 U23840 ( .A1(n11602), .A2(keyinput55), .B1(keyinput78), .B2(n20942), 
        .ZN(n20941) );
  OAI221_X1 U23841 ( .B1(n11602), .B2(keyinput55), .C1(n20942), .C2(keyinput78), .A(n20941), .ZN(n20955) );
  INV_X1 U23842 ( .A(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n20945) );
  AOI22_X1 U23843 ( .A1(n20945), .A2(keyinput36), .B1(keyinput12), .B2(n20944), 
        .ZN(n20943) );
  OAI221_X1 U23844 ( .B1(n20945), .B2(keyinput36), .C1(n20944), .C2(keyinput12), .A(n20943), .ZN(n20954) );
  AOI22_X1 U23845 ( .A1(n20948), .A2(keyinput101), .B1(n20947), .B2(keyinput38), .ZN(n20946) );
  OAI221_X1 U23846 ( .B1(n20948), .B2(keyinput101), .C1(n20947), .C2(
        keyinput38), .A(n20946), .ZN(n20953) );
  INV_X1 U23847 ( .A(P3_DATAO_REG_22__SCAN_IN), .ZN(n20951) );
  AOI22_X1 U23848 ( .A1(n20951), .A2(keyinput14), .B1(keyinput30), .B2(n20950), 
        .ZN(n20949) );
  OAI221_X1 U23849 ( .B1(n20951), .B2(keyinput14), .C1(n20950), .C2(keyinput30), .A(n20949), .ZN(n20952) );
  NOR4_X1 U23850 ( .A1(n20955), .A2(n20954), .A3(n20953), .A4(n20952), .ZN(
        n20973) );
  INV_X1 U23851 ( .A(P2_UWORD_REG_8__SCAN_IN), .ZN(n20958) );
  AOI22_X1 U23852 ( .A1(n20958), .A2(keyinput109), .B1(n20957), .B2(keyinput65), .ZN(n20956) );
  OAI221_X1 U23853 ( .B1(n20958), .B2(keyinput109), .C1(n20957), .C2(
        keyinput65), .A(n20956), .ZN(n20971) );
  INV_X1 U23854 ( .A(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n20960) );
  AOI22_X1 U23855 ( .A1(n20961), .A2(keyinput93), .B1(keyinput116), .B2(n20960), .ZN(n20959) );
  OAI221_X1 U23856 ( .B1(n20961), .B2(keyinput93), .C1(n20960), .C2(
        keyinput116), .A(n20959), .ZN(n20970) );
  INV_X1 U23857 ( .A(P2_UWORD_REG_4__SCAN_IN), .ZN(n20964) );
  AOI22_X1 U23858 ( .A1(n20964), .A2(keyinput85), .B1(keyinput40), .B2(n20963), 
        .ZN(n20962) );
  OAI221_X1 U23859 ( .B1(n20964), .B2(keyinput85), .C1(n20963), .C2(keyinput40), .A(n20962), .ZN(n20969) );
  AOI22_X1 U23860 ( .A1(n20967), .A2(keyinput104), .B1(n20966), .B2(keyinput3), 
        .ZN(n20965) );
  OAI221_X1 U23861 ( .B1(n20967), .B2(keyinput104), .C1(n20966), .C2(keyinput3), .A(n20965), .ZN(n20968) );
  NOR4_X1 U23862 ( .A1(n20971), .A2(n20970), .A3(n20969), .A4(n20968), .ZN(
        n20972) );
  NAND4_X1 U23863 ( .A1(n20975), .A2(n20974), .A3(n20973), .A4(n20972), .ZN(
        n20976) );
  NOR4_X1 U23864 ( .A1(n20979), .A2(n20978), .A3(n20977), .A4(n20976), .ZN(
        n20980) );
  XOR2_X1 U23865 ( .A(n20981), .B(n20980), .Z(n20982) );
  XNOR2_X1 U23866 ( .A(n20983), .B(n20982), .ZN(U355) );
  INV_X2 U11300 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n18624) );
  INV_X2 U11166 ( .A(n19845), .ZN(n13009) );
  CLKBUF_X2 U11178 ( .A(n13718), .Z(n13769) );
  CLKBUF_X2 U11179 ( .A(n12127), .Z(n9757) );
  CLKBUF_X1 U11210 ( .A(n12119), .Z(n13437) );
  CLKBUF_X1 U11220 ( .A(n10455), .Z(n11662) );
  INV_X1 U11235 ( .A(n9785), .ZN(n15318) );
  INV_X1 U11293 ( .A(n13936), .ZN(n13971) );
  CLKBUF_X1 U11295 ( .A(n12631), .Z(n9754) );
  INV_X2 U11583 ( .A(n11164), .ZN(n10944) );
  CLKBUF_X1 U12443 ( .A(n17215), .Z(n17234) );
  CLKBUF_X1 U12468 ( .A(n16367), .Z(n16371) );
endmodule

