

module b20_C_gen_AntiSAT_k_128_4 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, keyinput_f0, 
        keyinput_f1, keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5, 
        keyinput_f6, keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10, 
        keyinput_f11, keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15, 
        keyinput_f16, keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20, 
        keyinput_f21, keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25, 
        keyinput_f26, keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30, 
        keyinput_f31, keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35, 
        keyinput_f36, keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40, 
        keyinput_f41, keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45, 
        keyinput_f46, keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50, 
        keyinput_f51, keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55, 
        keyinput_f56, keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60, 
        keyinput_f61, keyinput_f62, keyinput_f63, keyinput_g0, keyinput_g1, 
        keyinput_g2, keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, 
        keyinput_g7, keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, 
        keyinput_g12, keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, 
        keyinput_g17, keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, 
        keyinput_g22, keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, 
        keyinput_g27, keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, 
        keyinput_g32, keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, 
        keyinput_g37, keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, 
        keyinput_g42, keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, 
        keyinput_g47, keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, 
        keyinput_g52, keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, 
        keyinput_g57, keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, 
        keyinput_g62, keyinput_g63, ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, 
        ADD_1068_U57, ADD_1068_U58, ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, 
        ADD_1068_U62, ADD_1068_U63, ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, 
        ADD_1068_U50, ADD_1068_U51, ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, 
        ADD_1068_U5, ADD_1068_U46, U126, U123, P1_U3355, P1_U3354, P1_U3353, 
        P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, 
        P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, 
        P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, 
        P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, 
        P1_U3324, P1_U3439, P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, 
        P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, 
        P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, 
        P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, 
        P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, 
        P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, 
        P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, 
        P1_U3501, P1_U3504, P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, 
        P1_U3513, P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, 
        P1_U3520, P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, 
        P1_U3527, P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, 
        P1_U3534, P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, 
        P1_U3541, P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, 
        P1_U3548, P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, 
        P1_U3292, P1_U3291, P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, 
        P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, 
        P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, 
        P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, 
        P1_U3356, P1_U3264, P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, 
        P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, 
        P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, 
        P1_U3244, P1_U3243, P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, 
        P1_U3559, P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, 
        P1_U3566, P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, 
        P1_U3573, P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, 
        P1_U3580, P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, 
        P1_U3241, P1_U3240, P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, 
        P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, 
        P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, 
        P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, 
        P1_U3213, P1_U3086, P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, 
        P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, 
        P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, 
        P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, 
        P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, 
        P2_U3264, P2_U3376, P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, 
        P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, 
        P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, 
        P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, 
        P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, 
        P2_U3396, P2_U3399, P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, 
        P2_U3417, P2_U3420, P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, 
        P2_U3438, P2_U3441, P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, 
        P2_U3450, P2_U3451, P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, 
        P2_U3457, P2_U3458, P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, 
        P2_U3464, P2_U3465, P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, 
        P2_U3471, P2_U3472, P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, 
        P2_U3478, P2_U3479, P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, 
        P2_U3485, P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, 
        P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, 
        P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, 
        P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, 
        P2_U3211, P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, 
        P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, 
        P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, 
        P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, 
        P2_U3183, P2_U3182, P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, 
        P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, 
        P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, 
        P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, 
        P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, 
        P2_U3181, P2_U3180, P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, 
        P2_U3174, P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, 
        P2_U3167, P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, 
        P2_U3160, P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, 
        P2_U3153, P2_U3151, P2_U3150, P2_U3893 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, keyinput_f0, keyinput_f1, keyinput_f2,
         keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, keyinput_f7,
         keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, keyinput_f12,
         keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, keyinput_f17,
         keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, keyinput_f22,
         keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, keyinput_f27,
         keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, keyinput_f32,
         keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, keyinput_f37,
         keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, keyinput_f42,
         keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, keyinput_f47,
         keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, keyinput_f52,
         keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, keyinput_f57,
         keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, keyinput_f62,
         keyinput_f63, keyinput_g0, keyinput_g1, keyinput_g2, keyinput_g3,
         keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7, keyinput_g8,
         keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12, keyinput_g13,
         keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17, keyinput_g18,
         keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22, keyinput_g23,
         keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27, keyinput_g28,
         keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32, keyinput_g33,
         keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37, keyinput_g38,
         keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42, keyinput_g43,
         keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47, keyinput_g48,
         keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52, keyinput_g53,
         keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57, keyinput_g58,
         keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62, keyinput_g63;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4350, n4351, n4352, n4353, n4354, n4356, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4469, n4470, n4471, n4472, n4473,
         n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483,
         n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493,
         n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503,
         n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513,
         n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523,
         n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533,
         n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543,
         n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553,
         n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563,
         n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573,
         n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583,
         n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593,
         n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603,
         n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613,
         n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623,
         n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633,
         n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643,
         n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654,
         n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664,
         n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674,
         n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684,
         n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694,
         n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704,
         n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714,
         n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724,
         n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734,
         n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744,
         n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754,
         n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764,
         n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774,
         n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784,
         n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794,
         n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804,
         n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814,
         n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824,
         n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834,
         n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844,
         n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854,
         n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864,
         n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874,
         n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884,
         n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894,
         n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904,
         n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914,
         n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924,
         n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934,
         n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944,
         n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954,
         n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964,
         n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974,
         n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984,
         n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994,
         n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004,
         n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014,
         n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024,
         n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034,
         n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044,
         n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054,
         n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064,
         n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074,
         n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084,
         n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094,
         n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104,
         n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114,
         n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124,
         n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134,
         n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144,
         n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154,
         n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164,
         n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174,
         n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184,
         n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194,
         n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204,
         n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214,
         n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224,
         n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234,
         n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244,
         n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254,
         n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264,
         n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274,
         n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284,
         n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294,
         n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304,
         n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314,
         n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324,
         n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334,
         n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344,
         n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354,
         n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364,
         n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374,
         n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384,
         n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394,
         n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404,
         n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414,
         n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424,
         n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434,
         n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444,
         n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454,
         n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464,
         n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474,
         n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484,
         n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494,
         n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504,
         n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514,
         n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524,
         n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534,
         n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544,
         n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554,
         n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564,
         n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574,
         n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584,
         n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594,
         n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604,
         n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614,
         n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624,
         n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634,
         n5635, n5636, n5637, n5638, n5639, n5640, n5642, n5643, n5644, n5645,
         n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655,
         n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665,
         n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675,
         n5676, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686,
         n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5695, n5696, n5697,
         n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5707, n5708,
         n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718,
         n5719, n5720, n5721, n5723, n5724, n5725, n5726, n5729, n5730, n5731,
         n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741,
         n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751,
         n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761,
         n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771,
         n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781,
         n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791,
         n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801,
         n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811,
         n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821,
         n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831,
         n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841,
         n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851,
         n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861,
         n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871,
         n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881,
         n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891,
         n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901,
         n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911,
         n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921,
         n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931,
         n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941,
         n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951,
         n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961,
         n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971,
         n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981,
         n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991,
         n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001,
         n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011,
         n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021,
         n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031,
         n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041,
         n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051,
         n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061,
         n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071,
         n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081,
         n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091,
         n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101,
         n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111,
         n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121,
         n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131,
         n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141,
         n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151,
         n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161,
         n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171,
         n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181,
         n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191,
         n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201,
         n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211,
         n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221,
         n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231,
         n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241,
         n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251,
         n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261,
         n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271,
         n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281,
         n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291,
         n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301,
         n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311,
         n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321,
         n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331,
         n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341,
         n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351,
         n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361,
         n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371,
         n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381,
         n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391,
         n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401,
         n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411,
         n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421,
         n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431,
         n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441,
         n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451,
         n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461,
         n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471,
         n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481,
         n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491,
         n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501,
         n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511,
         n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521,
         n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531,
         n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541,
         n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551,
         n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561,
         n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571,
         n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581,
         n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591,
         n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601,
         n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611,
         n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621,
         n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631,
         n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641,
         n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651,
         n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661,
         n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671,
         n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681,
         n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691,
         n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701,
         n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711,
         n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721,
         n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731,
         n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741,
         n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751,
         n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761,
         n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771,
         n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781,
         n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791,
         n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801,
         n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811,
         n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821,
         n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831,
         n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841,
         n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851,
         n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861,
         n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871,
         n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881,
         n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891,
         n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901,
         n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911,
         n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921,
         n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931,
         n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941,
         n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951,
         n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961,
         n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971,
         n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981,
         n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991,
         n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001,
         n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011,
         n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021,
         n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031,
         n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041,
         n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051,
         n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061,
         n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071,
         n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081,
         n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091,
         n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101,
         n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111,
         n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121,
         n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131,
         n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141,
         n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151,
         n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161,
         n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171,
         n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181,
         n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191,
         n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201,
         n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211,
         n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221,
         n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231,
         n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241,
         n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251,
         n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261,
         n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271,
         n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281,
         n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291,
         n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301,
         n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311,
         n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321,
         n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331,
         n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341,
         n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351,
         n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361,
         n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371,
         n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381,
         n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391,
         n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401,
         n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411,
         n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421,
         n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431,
         n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441,
         n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451,
         n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461,
         n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471,
         n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481,
         n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491,
         n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501,
         n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511,
         n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521,
         n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531,
         n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541,
         n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551,
         n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561,
         n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571,
         n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581,
         n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591,
         n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601,
         n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611,
         n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621,
         n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631,
         n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641,
         n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651,
         n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661,
         n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671,
         n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681,
         n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691,
         n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701,
         n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711,
         n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721,
         n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731,
         n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741,
         n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751,
         n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761,
         n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771,
         n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781,
         n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791,
         n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801,
         n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811,
         n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821,
         n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831,
         n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841,
         n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851,
         n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861,
         n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871,
         n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881,
         n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891,
         n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901,
         n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911,
         n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921,
         n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931,
         n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941,
         n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951,
         n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961,
         n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971,
         n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981,
         n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991,
         n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001,
         n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011,
         n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021,
         n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031,
         n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041,
         n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051,
         n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061,
         n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071,
         n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081,
         n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091,
         n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101,
         n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111,
         n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121,
         n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131,
         n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141,
         n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151,
         n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161,
         n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171,
         n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181,
         n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191,
         n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201,
         n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211,
         n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221,
         n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231,
         n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241,
         n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251,
         n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261,
         n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271,
         n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281,
         n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291,
         n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301,
         n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311,
         n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321,
         n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331,
         n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341,
         n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351,
         n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361,
         n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371,
         n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381,
         n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391,
         n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401,
         n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411,
         n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421,
         n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431,
         n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441,
         n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451,
         n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461,
         n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471,
         n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481,
         n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491,
         n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501,
         n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511,
         n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521,
         n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531,
         n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541,
         n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551,
         n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561,
         n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571,
         n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581,
         n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591,
         n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601,
         n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611,
         n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621,
         n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631,
         n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641,
         n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651,
         n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661,
         n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671,
         n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681,
         n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691,
         n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701,
         n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711,
         n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721,
         n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731,
         n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741,
         n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751,
         n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761,
         n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771,
         n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781,
         n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791,
         n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801,
         n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811,
         n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821,
         n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831,
         n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841,
         n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851,
         n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861,
         n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871,
         n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881,
         n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891,
         n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901,
         n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911,
         n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921,
         n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931,
         n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941,
         n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951,
         n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961,
         n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971,
         n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981,
         n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991,
         n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001,
         n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011,
         n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021,
         n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031,
         n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041,
         n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051,
         n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061,
         n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071,
         n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081,
         n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091,
         n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101,
         n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111,
         n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121,
         n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131,
         n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141,
         n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151,
         n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161,
         n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171,
         n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181,
         n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191,
         n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201,
         n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211,
         n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221,
         n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231,
         n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241,
         n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251,
         n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261,
         n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271,
         n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281,
         n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291,
         n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301,
         n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311,
         n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321,
         n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331,
         n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341,
         n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351,
         n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361,
         n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371,
         n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381,
         n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391,
         n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401,
         n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411,
         n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421,
         n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431,
         n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441,
         n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451,
         n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461,
         n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471,
         n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9480, n9481, n9482,
         n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492,
         n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502,
         n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512,
         n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522,
         n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532,
         n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542,
         n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552,
         n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562,
         n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572,
         n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582,
         n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
         n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602,
         n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
         n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
         n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
         n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
         n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
         n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
         n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
         n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
         n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
         n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
         n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
         n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
         n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
         n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
         n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
         n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
         n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
         n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
         n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
         n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
         n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
         n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
         n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
         n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193,
         n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
         n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209,
         n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217,
         n10218, n10222;

  AND2_X1 U4856 ( .A1(n9307), .A2(n9309), .ZN(n9432) );
  AND2_X1 U4857 ( .A1(n9084), .A2(n8950), .ZN(n4351) );
  NAND2_X1 U4858 ( .A1(n4356), .A2(n4354), .ZN(n4859) );
  NAND2_X1 U4859 ( .A1(n4452), .A2(n5704), .ZN(n4356) );
  NOR2_X1 U4860 ( .A1(n9117), .A2(n6840), .ZN(n4354) );
  NAND2_X1 U4862 ( .A1(n7751), .A2(n6329), .ZN(n8616) );
  NAND2_X1 U4863 ( .A1(n5690), .A2(n4360), .ZN(n4359) );
  AND2_X1 U4864 ( .A1(n5689), .A2(n9113), .ZN(n4360) );
  MUX2_X1 U4865 ( .A(n5686), .B(n5685), .S(n6840), .Z(n5690) );
  OR2_X1 U4866 ( .A1(n7482), .A2(n8114), .ZN(n7484) );
  AOI21_X1 U4867 ( .B1(n5650), .B2(n5649), .A(n5648), .ZN(n5654) );
  AND2_X1 U4868 ( .A1(n4980), .A2(n6214), .ZN(n4353) );
  NAND2_X1 U4869 ( .A1(n4361), .A2(n5640), .ZN(n5646) );
  INV_X1 U4870 ( .A(n7305), .ZN(n4362) );
  INV_X1 U4871 ( .A(n6840), .ZN(n4365) );
  NAND2_X1 U4872 ( .A1(n5625), .A2(n10222), .ZN(n5623) );
  MUX2_X1 U4873 ( .A(n5621), .B(n5620), .S(n4365), .Z(n5625) );
  CLKBUF_X1 U4876 ( .A(P1_IR_REG_12__SCAN_IN), .Z(n4366) );
  NAND2_X1 U4877 ( .A1(n6181), .A2(n6182), .ZN(n6489) );
  NAND2_X1 U4878 ( .A1(n4803), .A2(n5617), .ZN(n6737) );
  INV_X1 U4879 ( .A(n5297), .ZN(n5542) );
  INV_X1 U4880 ( .A(n6182), .ZN(n6183) );
  AND4_X1 U4881 ( .A1(n6171), .A2(n6172), .A3(n6173), .A4(n6174), .ZN(n6182)
         );
  INV_X1 U4882 ( .A(n9726), .ZN(n6757) );
  AND2_X1 U4883 ( .A1(n5275), .A2(n5274), .ZN(n4895) );
  AND2_X1 U4884 ( .A1(n5272), .A2(n5273), .ZN(n4896) );
  NAND2_X2 U4885 ( .A1(n6812), .A2(n4369), .ZN(n6521) );
  INV_X1 U4886 ( .A(n5138), .ZN(n7867) );
  AND2_X1 U4888 ( .A1(n5114), .A2(n4808), .ZN(n5813) );
  AND2_X1 U4889 ( .A1(n4971), .A2(n4970), .ZN(n4969) );
  AND3_X1 U4890 ( .A1(n5116), .A2(n5115), .A3(n5576), .ZN(n5120) );
  NOR2_X1 U4891 ( .A1(P2_IR_REG_14__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .ZN(
        n6102) );
  NOR2_X1 U4892 ( .A1(n5110), .A2(n4816), .ZN(n4815) );
  NOR2_X1 U4893 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n4820) );
  NAND3_X1 U4894 ( .A1(n4352), .A2(n4350), .A3(n5801), .ZN(n5800) );
  NAND2_X1 U4895 ( .A1(n5720), .A2(n4351), .ZN(n4350) );
  NAND2_X1 U4896 ( .A1(n5726), .A2(n5725), .ZN(n4352) );
  NAND2_X1 U4897 ( .A1(n4979), .A2(n4353), .ZN(n6227) );
  OAI21_X1 U4901 ( .B1(n8473), .B2(n4648), .A(n4647), .ZN(n8452) );
  NAND2_X1 U4902 ( .A1(n4359), .A2(n5693), .ZN(n4453) );
  NAND3_X1 U4903 ( .A1(n4364), .A2(n4363), .A3(n4362), .ZN(n4361) );
  NAND2_X1 U4904 ( .A1(n5634), .A2(n6840), .ZN(n4363) );
  NAND2_X1 U4905 ( .A1(n5635), .A2(n4365), .ZN(n4364) );
  NAND2_X1 U4906 ( .A1(n6933), .A2(n5287), .ZN(n6749) );
  NAND2_X1 U4907 ( .A1(n4367), .A2(n7827), .ZN(n5683) );
  NAND4_X1 U4908 ( .A1(n5676), .A2(n5675), .A3(n5673), .A4(n5674), .ZN(n4367)
         );
  NAND2_X1 U4909 ( .A1(n5277), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n5272) );
  NOR2_X2 U4910 ( .A1(n7867), .A2(n9478), .ZN(n5277) );
  XNOR2_X2 U4911 ( .A(n9719), .B(n8823), .ZN(n6934) );
  NAND2_X4 U4912 ( .A1(n4896), .A2(n4895), .ZN(n9719) );
  INV_X1 U4913 ( .A(n5880), .ZN(n6052) );
  INV_X1 U4914 ( .A(n8289), .ZN(n8284) );
  INV_X1 U4915 ( .A(n6915), .ZN(n4488) );
  INV_X2 U4916 ( .A(n4371), .ZN(n6055) );
  NAND2_X1 U4917 ( .A1(n4639), .A2(n4638), .ZN(n4376) );
  INV_X2 U4918 ( .A(n7350), .ZN(n6475) );
  AND2_X1 U4919 ( .A1(n6015), .A2(n6014), .ZN(n8907) );
  CLKBUF_X3 U4920 ( .A(n5278), .Z(n5427) );
  NAND2_X1 U4921 ( .A1(n9207), .A2(n9211), .ZN(n9209) );
  NAND2_X1 U4922 ( .A1(n5836), .A2(n9080), .ZN(n7243) );
  AND3_X1 U4923 ( .A1(n5340), .A2(n5339), .A3(n5338), .ZN(n6857) );
  XNOR2_X1 U4924 ( .A(n5100), .B(n5099), .ZN(n5141) );
  XNOR2_X1 U4925 ( .A(n4992), .B(SI_2_), .ZN(n5294) );
  NAND2_X1 U4926 ( .A1(n5468), .A2(n5467), .ZN(n9427) );
  INV_X1 U4927 ( .A(n8582), .ZN(n8633) );
  INV_X1 U4928 ( .A(n7439), .ZN(n9746) );
  XNOR2_X1 U4929 ( .A(n5268), .B(n5267), .ZN(n8970) );
  AND2_X1 U4930 ( .A1(n4406), .A2(n4539), .ZN(n4368) );
  NAND2_X2 U4931 ( .A1(n5848), .A2(n6058), .ZN(n5862) );
  NAND2_X2 U4932 ( .A1(n7854), .A2(n7853), .ZN(n7895) );
  NAND2_X1 U4933 ( .A1(n6117), .A2(n6133), .ZN(n4369) );
  NAND2_X1 U4934 ( .A1(n6117), .A2(n6133), .ZN(n4370) );
  NAND2_X1 U4935 ( .A1(n6117), .A2(n6133), .ZN(n8415) );
  NAND3_X2 U4936 ( .A1(n9209), .A2(n9194), .A3(n9192), .ZN(n9193) );
  NAND2_X2 U4937 ( .A1(n5399), .A2(n5398), .ZN(n7437) );
  INV_X1 U4938 ( .A(n8325), .ZN(n6199) );
  NAND4_X2 U4939 ( .A1(n6191), .A2(n6190), .A3(n6189), .A4(n6188), .ZN(n8325)
         );
  OAI21_X2 U4940 ( .B1(n5396), .B2(n5395), .A(n5017), .ZN(n5360) );
  AOI21_X2 U4941 ( .B1(n8879), .B2(n8878), .A(n8877), .ZN(n8881) );
  NAND3_X2 U4942 ( .A1(n5540), .A2(n5539), .A3(n5538), .ZN(n7863) );
  OAI211_X2 U4943 ( .C1(n7231), .C2(n4757), .A(n7330), .B(n4756), .ZN(n7388)
         );
  NAND2_X2 U4944 ( .A1(n4730), .A2(n4728), .ZN(n7951) );
  AOI211_X2 U4945 ( .C1(n9320), .C2(n9143), .A(n9142), .B(n9141), .ZN(n9144)
         );
  XNOR2_X2 U4946 ( .A(n4610), .B(P2_IR_REG_2__SCAN_IN), .ZN(n8338) );
  XNOR2_X2 U4947 ( .A(n5141), .B(SI_29_), .ZN(n7866) );
  AOI22_X2 U4948 ( .A1(n7624), .A2(n7623), .B1(n9769), .B2(n9777), .ZN(n7691)
         );
  AND2_X1 U4949 ( .A1(n9322), .A2(n9321), .ZN(n4587) );
  NAND2_X1 U4950 ( .A1(n9106), .A2(n9105), .ZN(n9147) );
  NAND2_X1 U4951 ( .A1(n7917), .A2(n7916), .ZN(n8049) );
  NOR2_X1 U4952 ( .A1(n9178), .A2(n9116), .ZN(n9160) );
  OAI21_X1 U4953 ( .B1(n7906), .B2(n8537), .A(n7905), .ZN(n8028) );
  NAND2_X1 U4954 ( .A1(n6509), .A2(n8259), .ZN(n8461) );
  NOR2_X1 U4955 ( .A1(n8085), .A2(n8086), .ZN(n8083) );
  NAND2_X1 U4956 ( .A1(n5081), .A2(n5080), .ZN(n5171) );
  XNOR2_X1 U4957 ( .A(n4481), .B(n8355), .ZN(n8344) );
  NAND2_X1 U4958 ( .A1(n4865), .A2(n4866), .ZN(n5194) );
  OR2_X1 U4959 ( .A1(n7685), .A2(n7708), .ZN(n7687) );
  NAND2_X1 U4960 ( .A1(n5043), .A2(n5042), .ZN(n5494) );
  INV_X1 U4961 ( .A(n7271), .ZN(n7425) );
  INV_X4 U4962 ( .A(n7183), .ZN(n7934) );
  INV_X1 U4963 ( .A(n8107), .ZN(n8152) );
  INV_X1 U4964 ( .A(n6058), .ZN(n6011) );
  INV_X4 U4965 ( .A(n5892), .ZN(n6049) );
  NAND2_X1 U4966 ( .A1(n8960), .A2(n6867), .ZN(n5738) );
  NAND2_X1 U4967 ( .A1(n6934), .A2(n6935), .ZN(n6933) );
  NOR2_X1 U4968 ( .A1(n8961), .A2(n6954), .ZN(n5616) );
  INV_X2 U4969 ( .A(n6833), .ZN(n8960) );
  NAND2_X1 U4970 ( .A1(n5821), .A2(n5820), .ZN(n5837) );
  BUF_X1 U4971 ( .A(n5276), .Z(n4372) );
  NOR2_X2 U4972 ( .A1(n9478), .A2(n5138), .ZN(n5276) );
  AND2_X1 U4973 ( .A1(n7383), .A2(n7863), .ZN(n6080) );
  OAI21_X1 U4974 ( .B1(n8783), .B2(n8782), .A(n8936), .ZN(n8787) );
  NOR2_X1 U4975 ( .A1(n8783), .A2(n6077), .ZN(n6096) );
  AOI21_X1 U4976 ( .B1(n4841), .B2(n4553), .A(n4552), .ZN(n8782) );
  NAND2_X1 U4977 ( .A1(n4469), .A2(n4467), .ZN(n4466) );
  OAI21_X1 U4978 ( .B1(n4707), .B2(n4706), .A(n4708), .ZN(n6580) );
  AND2_X1 U4979 ( .A1(n4448), .A2(n4582), .ZN(n4581) );
  OR2_X1 U4980 ( .A1(n4587), .A2(n9796), .ZN(n4582) );
  AND2_X1 U4981 ( .A1(n4823), .A2(n4821), .ZN(n8905) );
  NAND2_X1 U4982 ( .A1(n8099), .A2(n8098), .ZN(n8679) );
  NAND2_X1 U4983 ( .A1(n4897), .A2(n9104), .ZN(n9162) );
  AND2_X1 U4984 ( .A1(n5130), .A2(n5129), .ZN(n9439) );
  NOR2_X1 U4985 ( .A1(n9160), .A2(n9161), .ZN(n9159) );
  OAI21_X1 U4986 ( .B1(n5711), .B2(n5710), .A(n5709), .ZN(n5713) );
  AOI21_X1 U4987 ( .B1(n4947), .B2(n4950), .A(n4404), .ZN(n4945) );
  OAI21_X1 U4988 ( .B1(n5564), .B2(n5563), .A(n5562), .ZN(n5568) );
  NAND2_X1 U4989 ( .A1(n8268), .A2(n8269), .ZN(n8451) );
  NAND2_X1 U4990 ( .A1(n5154), .A2(n5153), .ZN(n9318) );
  NAND2_X1 U4991 ( .A1(n5097), .A2(n5096), .ZN(n5100) );
  INV_X1 U4992 ( .A(n8692), .ZN(n8458) );
  INV_X1 U4993 ( .A(n4563), .ZN(n9237) );
  AND2_X1 U4994 ( .A1(n6450), .A2(n6449), .ZN(n8692) );
  AOI21_X1 U4995 ( .B1(n4655), .B2(n4661), .A(n4654), .ZN(n4653) );
  NAND2_X1 U4996 ( .A1(n5173), .A2(n5172), .ZN(n9164) );
  NAND2_X1 U4997 ( .A1(n4613), .A2(n4612), .ZN(n4454) );
  NAND2_X1 U4998 ( .A1(n6440), .A2(n6439), .ZN(n8698) );
  XNOR2_X1 U4999 ( .A(n5162), .B(n5161), .ZN(n7805) );
  NAND2_X1 U5000 ( .A1(n4546), .A2(n7761), .ZN(n4545) );
  NAND2_X1 U5001 ( .A1(n5087), .A2(n5086), .ZN(n5162) );
  AOI21_X1 U5002 ( .B1(n4550), .B2(n4548), .A(n4418), .ZN(n4547) );
  XNOR2_X1 U5003 ( .A(n5171), .B(n5170), .ZN(n7744) );
  AOI21_X1 U5004 ( .B1(n9098), .B2(n9097), .A(n4559), .ZN(n9286) );
  AOI21_X1 U5005 ( .B1(n4737), .B2(n4740), .A(n4736), .ZN(n4735) );
  NAND2_X1 U5006 ( .A1(n5183), .A2(n5182), .ZN(n9201) );
  OR2_X1 U5007 ( .A1(n8352), .A2(n8353), .ZN(n4775) );
  NAND2_X1 U5008 ( .A1(n5235), .A2(n5234), .ZN(n9241) );
  NAND2_X1 U5009 ( .A1(n6502), .A2(n8232), .ZN(n8548) );
  NAND2_X1 U5010 ( .A1(n6412), .A2(n6411), .ZN(n8727) );
  NAND2_X1 U5011 ( .A1(n5196), .A2(n5195), .ZN(n9363) );
  NAND2_X1 U5012 ( .A1(n6403), .A2(n6402), .ZN(n8733) );
  NAND2_X1 U5013 ( .A1(n5247), .A2(n5246), .ZN(n9388) );
  AOI21_X1 U5014 ( .B1(n4903), .B2(n4901), .A(n4415), .ZN(n4900) );
  XNOR2_X1 U5015 ( .A(n5194), .B(n5193), .ZN(n7637) );
  NOR2_X1 U5016 ( .A1(n7833), .A2(n5667), .ZN(n4784) );
  AND2_X1 U5017 ( .A1(n5587), .A2(n5586), .ZN(n7827) );
  OR2_X1 U5018 ( .A1(n9392), .A2(n9256), .ZN(n5687) );
  OR2_X1 U5019 ( .A1(n8744), .A2(n8578), .ZN(n8232) );
  NAND2_X1 U5020 ( .A1(n6392), .A2(n6391), .ZN(n8063) );
  NAND2_X1 U5021 ( .A1(n4907), .A2(n4904), .ZN(n4902) );
  NAND2_X1 U5022 ( .A1(n5521), .A2(n5520), .ZN(n9300) );
  NAND2_X1 U5023 ( .A1(n5059), .A2(n5058), .ZN(n5245) );
  NAND2_X1 U5024 ( .A1(n8861), .A2(n7824), .ZN(n5767) );
  NAND2_X1 U5025 ( .A1(n6369), .A2(n6368), .ZN(n8744) );
  NAND2_X1 U5026 ( .A1(n5507), .A2(n5506), .ZN(n9096) );
  NAND2_X1 U5027 ( .A1(n6718), .A2(n8097), .ZN(n6369) );
  NAND2_X1 U5028 ( .A1(n6378), .A2(n6377), .ZN(n8750) );
  NAND2_X1 U5029 ( .A1(n7277), .A2(n7276), .ZN(n4777) );
  XNOR2_X1 U5030 ( .A(n4642), .B(n5503), .ZN(n6718) );
  NAND2_X1 U5031 ( .A1(n5431), .A2(n7517), .ZN(n7620) );
  XNOR2_X1 U5032 ( .A(n5494), .B(n5493), .ZN(n6671) );
  OAI21_X1 U5033 ( .B1(n5494), .B2(n5044), .A(n5046), .ZN(n4642) );
  AND2_X1 U5034 ( .A1(n7280), .A2(n7279), .ZN(n7369) );
  OR2_X1 U5035 ( .A1(n7061), .A2(n7062), .ZN(n4502) );
  NAND2_X1 U5036 ( .A1(n5484), .A2(n5483), .ZN(n7819) );
  AND2_X1 U5037 ( .A1(n7619), .A2(n5656), .ZN(n5596) );
  NOR2_X1 U5038 ( .A1(n7073), .A2(n7063), .ZN(n7113) );
  NAND2_X1 U5039 ( .A1(n5438), .A2(n5437), .ZN(n9780) );
  OR2_X1 U5040 ( .A1(n7816), .A2(n9777), .ZN(n7619) );
  NOR2_X1 U5041 ( .A1(n7060), .A2(n7059), .ZN(n7095) );
  XNOR2_X1 U5042 ( .A(n4566), .B(n5447), .ZN(n6636) );
  NAND2_X1 U5043 ( .A1(n4674), .A2(n4678), .ZN(n5464) );
  OAI21_X1 U5044 ( .B1(n5433), .B2(n5034), .A(n5033), .ZN(n4566) );
  AOI21_X1 U5045 ( .B1(n5623), .B2(n5738), .A(n5622), .ZN(n5624) );
  NAND2_X1 U5046 ( .A1(n4667), .A2(n5030), .ZN(n5433) );
  XNOR2_X1 U5047 ( .A(n5419), .B(n5418), .ZN(n6628) );
  NAND2_X1 U5048 ( .A1(n7491), .A2(n8158), .ZN(n7490) );
  AND2_X1 U5049 ( .A1(n6289), .A2(n6288), .ZN(n7679) );
  NAND2_X2 U5050 ( .A1(n7163), .A2(n8624), .ZN(n8089) );
  NAND2_X1 U5051 ( .A1(n5364), .A2(n5363), .ZN(n9747) );
  AND2_X2 U5052 ( .A1(n7293), .A2(n8624), .ZN(n8582) );
  NAND2_X1 U5053 ( .A1(n5023), .A2(n4592), .ZN(n4591) );
  NAND2_X1 U5054 ( .A1(n6996), .A2(n6995), .ZN(n7000) );
  NAND2_X1 U5055 ( .A1(n7197), .A2(n8152), .ZN(n7198) );
  AND2_X1 U5056 ( .A1(n7478), .A2(n8168), .ZN(n8111) );
  NAND2_X1 U5057 ( .A1(n4558), .A2(n4860), .ZN(n5396) );
  BUF_X4 U5058 ( .A(n5848), .Z(n4371) );
  INV_X4 U5059 ( .A(n5871), .ZN(n5892) );
  AND3_X1 U5060 ( .A1(n5379), .A2(n5378), .A3(n5377), .ZN(n7311) );
  AND3_X1 U5061 ( .A1(n5371), .A2(n5370), .A3(n5369), .ZN(n7473) );
  INV_X1 U5062 ( .A(n9865), .ZN(n6181) );
  AND2_X1 U5063 ( .A1(n5318), .A2(n5317), .ZN(n6833) );
  NAND2_X1 U5064 ( .A1(n5581), .A2(n5797), .ZN(n5834) );
  XNOR2_X1 U5065 ( .A(n6532), .B(n6531), .ZN(n6542) );
  INV_X2 U5066 ( .A(n6225), .ZN(n8097) );
  NAND2_X1 U5067 ( .A1(n5816), .A2(n5815), .ZN(n7703) );
  OR2_X1 U5068 ( .A1(n6534), .A2(n6533), .ZN(n6536) );
  XNOR2_X1 U5069 ( .A(n6341), .B(P2_IR_REG_13__SCAN_IN), .ZN(n8351) );
  INV_X1 U5070 ( .A(n5830), .ZN(n5831) );
  NAND2_X2 U5071 ( .A1(n6138), .A2(n6137), .ZN(n7348) );
  AND2_X2 U5072 ( .A1(n8771), .A2(n8769), .ZN(n6170) );
  NAND2_X4 U5073 ( .A1(n8769), .A2(n6136), .ZN(n6186) );
  INV_X2 U5074 ( .A(n6521), .ZN(n6585) );
  OAI21_X1 U5075 ( .B1(n5812), .B2(n5811), .A(n5810), .ZN(n5816) );
  MUX2_X1 U5076 ( .A(n5134), .B(n5133), .S(P1_IR_REG_30__SCAN_IN), .Z(n9478)
         );
  AND2_X1 U5077 ( .A1(n4594), .A2(n5026), .ZN(n4590) );
  INV_X1 U5078 ( .A(n6137), .ZN(n6136) );
  XNOR2_X1 U5079 ( .A(n4542), .B(P2_IR_REG_29__SCAN_IN), .ZN(n6137) );
  INV_X1 U5080 ( .A(n5418), .ZN(n4594) );
  XNOR2_X1 U5081 ( .A(n5128), .B(n5127), .ZN(n9485) );
  NAND2_X1 U5082 ( .A1(n8332), .A2(n8331), .ZN(n8330) );
  XNOR2_X1 U5083 ( .A(n6222), .B(P2_IR_REG_4__SCAN_IN), .ZN(n6899) );
  NAND2_X2 U5084 ( .A1(n4810), .A2(P1_U3086), .ZN(n9487) );
  NAND2_X2 U5085 ( .A1(n4810), .A2(P2_U3151), .ZN(n8777) );
  AND2_X1 U5086 ( .A1(n4398), .A2(n4963), .ZN(n6250) );
  NOR2_X1 U5087 ( .A1(n5121), .A2(P1_IR_REG_15__SCAN_IN), .ZN(n4808) );
  NAND4_X1 U5088 ( .A1(n5120), .A2(n5119), .A3(n5118), .A4(n5117), .ZN(n5121)
         );
  NAND3_X1 U5089 ( .A1(n4636), .A2(n4635), .A3(n4634), .ZN(n4639) );
  NAND3_X1 U5090 ( .A1(n4637), .A2(P1_ADDR_REG_19__SCAN_IN), .A3(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n4638) );
  AND2_X1 U5091 ( .A1(n6194), .A2(n6099), .ZN(n4964) );
  NOR2_X2 U5092 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n6194) );
  INV_X4 U5093 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  NOR2_X1 U5094 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_13__SCAN_IN), .ZN(
        n6103) );
  INV_X1 U5095 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n4635) );
  INV_X1 U5096 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4634) );
  INV_X1 U5097 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4637) );
  INV_X1 U5098 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n5107) );
  INV_X1 U5099 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5320) );
  INV_X4 U5100 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  INV_X1 U5101 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5576) );
  XNOR2_X1 U5102 ( .A(n5136), .B(n5125), .ZN(n5822) );
  NAND2_X1 U5103 ( .A1(n9470), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5136) );
  NAND2_X2 U5104 ( .A1(n7994), .A2(n7993), .ZN(n8004) );
  NOR2_X2 U5105 ( .A1(n8083), .A2(n7899), .ZN(n7994) );
  AND2_X1 U5106 ( .A1(n9478), .A2(n5138), .ZN(n5289) );
  AOI21_X2 U5107 ( .B1(n4814), .B2(n4427), .A(n4813), .ZN(n7467) );
  NAND2_X1 U5108 ( .A1(n6622), .A2(n4810), .ZN(n4373) );
  NAND2_X1 U5109 ( .A1(n6622), .A2(n4810), .ZN(n4374) );
  NAND2_X1 U5110 ( .A1(n6622), .A2(n4810), .ZN(n5297) );
  NAND2_X1 U5111 ( .A1(n4639), .A2(n4638), .ZN(n4375) );
  NAND2_X1 U5112 ( .A1(n8258), .A2(n8257), .ZN(n4535) );
  NAND2_X1 U5113 ( .A1(n8561), .A2(n6386), .ZN(n4682) );
  OR2_X1 U5114 ( .A1(n8319), .A2(n9890), .ZN(n8187) );
  INV_X1 U5115 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n4970) );
  NAND2_X1 U5116 ( .A1(n9103), .A2(n9199), .ZN(n4577) );
  NAND2_X1 U5117 ( .A1(n7707), .A2(n9775), .ZN(n4910) );
  AND2_X1 U5118 ( .A1(n6099), .A2(n4537), .ZN(n4536) );
  INV_X1 U5119 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n4537) );
  INV_X1 U5120 ( .A(n6540), .ZN(n6115) );
  AOI21_X1 U5121 ( .B1(n7198), .B2(n8155), .A(n8154), .ZN(n8156) );
  OAI21_X1 U5122 ( .B1(n4526), .B2(n4529), .A(n8289), .ZN(n4516) );
  AOI21_X1 U5123 ( .B1(n4377), .B2(n8228), .A(n4423), .ZN(n4526) );
  OAI21_X1 U5124 ( .B1(n4534), .B2(n4533), .A(n8270), .ZN(n8279) );
  NAND2_X1 U5125 ( .A1(n8265), .A2(n8266), .ZN(n4533) );
  OR2_X1 U5126 ( .A1(n9316), .A2(n8951), .ZN(n5716) );
  AOI21_X1 U5127 ( .B1(n4679), .B2(n5034), .A(n4416), .ZN(n4678) );
  NAND2_X1 U5128 ( .A1(n5027), .A2(n10132), .ZN(n5030) );
  NAND2_X1 U5129 ( .A1(n4682), .A2(n4403), .ZN(n6387) );
  OR2_X1 U5130 ( .A1(n8324), .A2(n7507), .ZN(n8167) );
  NAND2_X1 U5131 ( .A1(n6545), .A2(n6544), .ZN(n7173) );
  OR2_X1 U5132 ( .A1(n8458), .A2(n8072), .ZN(n8268) );
  OR2_X1 U5133 ( .A1(n8704), .A2(n8486), .ZN(n8259) );
  OR2_X1 U5134 ( .A1(n8024), .A2(n8018), .ZN(n8254) );
  NAND2_X1 U5135 ( .A1(n7891), .A2(n8547), .ZN(n4973) );
  AND2_X1 U5136 ( .A1(n7975), .A2(n8547), .ZN(n8243) );
  OR2_X1 U5137 ( .A1(n8733), .A2(n8311), .ZN(n8242) );
  INV_X1 U5138 ( .A(n8421), .ZN(n6527) );
  OR2_X1 U5139 ( .A1(n8750), .A2(n8082), .ZN(n8225) );
  NAND2_X1 U5140 ( .A1(n4765), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6561) );
  AND2_X1 U5141 ( .A1(n4389), .A2(n4762), .ZN(n4761) );
  INV_X1 U5142 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n4762) );
  AND2_X1 U5143 ( .A1(n6481), .A2(n6483), .ZN(n4764) );
  NOR2_X1 U5144 ( .A1(n6106), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n4972) );
  NOR2_X1 U5145 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n6105) );
  NOR2_X1 U5146 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n6104) );
  NOR2_X1 U5147 ( .A1(n4965), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n4963) );
  NOR2_X1 U5148 ( .A1(n8829), .A2(n4828), .ZN(n4827) );
  INV_X1 U5149 ( .A(n6000), .ZN(n4828) );
  AOI21_X1 U5150 ( .B1(n4849), .B2(n4847), .A(n4408), .ZN(n4846) );
  INV_X1 U5151 ( .A(n4852), .ZN(n4847) );
  INV_X1 U5153 ( .A(n6789), .ZN(n4915) );
  NAND2_X1 U5154 ( .A1(n5093), .A2(n5092), .ZN(n5151) );
  NAND2_X1 U5155 ( .A1(n5162), .A2(n5161), .ZN(n5093) );
  NAND2_X1 U5156 ( .A1(n5071), .A2(n5070), .ZN(n5181) );
  NAND2_X1 U5157 ( .A1(n5194), .A2(n5193), .ZN(n5071) );
  INV_X1 U5158 ( .A(n5205), .ZN(n4868) );
  NAND2_X1 U5159 ( .A1(n5060), .A2(n10080), .ZN(n4876) );
  OR2_X1 U5160 ( .A1(n5480), .A2(SI_15_), .ZN(n5043) );
  AOI21_X1 U5161 ( .B1(n4862), .B2(n4864), .A(n4417), .ZN(n4860) );
  NAND2_X1 U5162 ( .A1(n5351), .A2(n4862), .ZN(n4558) );
  AND2_X1 U5163 ( .A1(n7921), .A2(n7919), .ZN(n4760) );
  OR2_X1 U5164 ( .A1(n8299), .A2(n8298), .ZN(n4539) );
  AND2_X1 U5165 ( .A1(n8296), .A2(n8298), .ZN(n4541) );
  NAND2_X1 U5166 ( .A1(n4767), .A2(n4483), .ZN(n4766) );
  OR2_X1 U5167 ( .A1(n8338), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n4483) );
  OR2_X1 U5168 ( .A1(n9836), .A2(n9835), .ZN(n4613) );
  NAND2_X1 U5169 ( .A1(n4491), .A2(n4490), .ZN(n4771) );
  INV_X1 U5170 ( .A(n9830), .ZN(n4490) );
  AND2_X1 U5171 ( .A1(n4972), .A2(n6107), .ZN(n4971) );
  INV_X1 U5172 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n6107) );
  OR2_X1 U5173 ( .A1(n6441), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n6453) );
  NAND2_X1 U5174 ( .A1(n6131), .A2(n6130), .ZN(n6441) );
  INV_X1 U5175 ( .A(n6431), .ZN(n6131) );
  AOI21_X1 U5176 ( .B1(n8118), .B2(n4722), .A(n4721), .ZN(n4720) );
  INV_X1 U5177 ( .A(n8195), .ZN(n4721) );
  XNOR2_X1 U5178 ( .A(n8323), .B(n7232), .ZN(n8158) );
  AND2_X1 U5179 ( .A1(n6512), .A2(n7294), .ZN(n7666) );
  AOI22_X1 U5180 ( .A1(n8483), .A2(n6438), .B1(n8499), .B2(n8024), .ZN(n8473)
         );
  AND2_X1 U5181 ( .A1(n6587), .A2(n6647), .ZN(n7162) );
  OAI21_X1 U5182 ( .B1(n6540), .B2(n4543), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n4542) );
  INV_X1 U5183 ( .A(n4977), .ZN(n4543) );
  AND2_X1 U5184 ( .A1(n4969), .A2(n6250), .ZN(n6156) );
  AND4_X1 U5185 ( .A1(n6111), .A2(n6110), .A3(n6109), .A4(n6108), .ZN(n6112)
         );
  AND2_X1 U5186 ( .A1(n6156), .A2(n6157), .ZN(n6482) );
  INV_X1 U5187 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n6157) );
  INV_X1 U5188 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n6481) );
  NAND2_X1 U5189 ( .A1(n4554), .A2(n5904), .ZN(n5905) );
  OAI21_X1 U5190 ( .B1(n7029), .B2(n4832), .A(n4830), .ZN(n4554) );
  NAND2_X1 U5191 ( .A1(n4834), .A2(n4833), .ZN(n4832) );
  NAND2_X1 U5192 ( .A1(n4831), .A2(n4834), .ZN(n4830) );
  AOI21_X1 U5193 ( .B1(n4837), .B2(n7031), .A(n4836), .ZN(n4835) );
  OR2_X1 U5194 ( .A1(n8922), .A2(n8923), .ZN(n4842) );
  INV_X1 U5195 ( .A(n5289), .ZN(n5559) );
  AOI21_X1 U5196 ( .B1(n4380), .B2(n4571), .A(n4421), .ZN(n4568) );
  INV_X1 U5197 ( .A(n9194), .ZN(n9190) );
  NAND2_X1 U5198 ( .A1(n4424), .A2(n4577), .ZN(n4572) );
  NAND2_X1 U5199 ( .A1(n4565), .A2(n4981), .ZN(n9251) );
  OR2_X1 U5200 ( .A1(n9392), .A2(n9396), .ZN(n9101) );
  INV_X1 U5201 ( .A(n4784), .ZN(n4783) );
  AOI21_X1 U5202 ( .B1(n4784), .B2(n4782), .A(n4781), .ZN(n4780) );
  INV_X1 U5203 ( .A(n5767), .ZN(n4781) );
  NAND2_X1 U5204 ( .A1(n4419), .A2(n4900), .ZN(n4562) );
  INV_X1 U5205 ( .A(n7719), .ZN(n4904) );
  NAND2_X1 U5206 ( .A1(n4923), .A2(n4924), .ZN(n7624) );
  AOI21_X1 U5207 ( .B1(n4925), .B2(n4931), .A(n4422), .ZN(n4924) );
  AND2_X1 U5208 ( .A1(n4927), .A2(n4926), .ZN(n4925) );
  INV_X1 U5209 ( .A(n7436), .ZN(n4930) );
  AND2_X1 U5210 ( .A1(n5746), .A2(n7264), .ZN(n6791) );
  AND2_X1 U5211 ( .A1(n9132), .A2(n9107), .ZN(n4921) );
  NAND2_X1 U5212 ( .A1(n5112), .A2(n5107), .ZN(n4816) );
  INV_X1 U5213 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5112) );
  MUX2_X1 U5214 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6116), .S(
        P2_IR_REG_27__SCAN_IN), .Z(n6117) );
  INV_X1 U5215 ( .A(n4494), .ZN(n4493) );
  OAI21_X1 U5216 ( .B1(n8400), .B2(n4495), .A(n8426), .ZN(n4494) );
  NAND2_X1 U5217 ( .A1(n8414), .A2(n4496), .ZN(n4495) );
  INV_X1 U5218 ( .A(n8398), .ZN(n4496) );
  OR2_X1 U5219 ( .A1(n6737), .A2(n5616), .ZN(n5621) );
  NAND2_X1 U5220 ( .A1(n4384), .A2(n8284), .ZN(n4514) );
  AND2_X1 U5221 ( .A1(n8191), .A2(n8179), .ZN(n4515) );
  NAND2_X1 U5222 ( .A1(n8203), .A2(n8195), .ZN(n8196) );
  NOR2_X1 U5223 ( .A1(n4524), .A2(n4523), .ZN(n4522) );
  NAND2_X1 U5224 ( .A1(n4519), .A2(n4377), .ZN(n4518) );
  INV_X1 U5225 ( .A(n4529), .ZN(n4519) );
  NAND2_X1 U5226 ( .A1(n5705), .A2(n5703), .ZN(n4452) );
  NAND2_X1 U5227 ( .A1(n4799), .A2(n4800), .ZN(n4796) );
  INV_X1 U5228 ( .A(n4799), .ZN(n4798) );
  NAND2_X1 U5229 ( .A1(n9445), .A2(n9166), .ZN(n5780) );
  NAND2_X1 U5230 ( .A1(n5243), .A2(SI_20_), .ZN(n4877) );
  AOI21_X1 U5231 ( .B1(n4894), .B2(n5039), .A(n4892), .ZN(n4891) );
  NOR2_X1 U5232 ( .A1(n4680), .A2(n5036), .ZN(n4679) );
  INV_X1 U5233 ( .A(n5033), .ZN(n4680) );
  INV_X1 U5234 ( .A(SI_10_), .ZN(n10053) );
  XNOR2_X1 U5235 ( .A(n7183), .B(n6181), .ZN(n7177) );
  NAND2_X1 U5236 ( .A1(n4608), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n6999) );
  NOR2_X1 U5237 ( .A1(n9815), .A2(n8392), .ZN(n4507) );
  NAND2_X1 U5238 ( .A1(n4511), .A2(n9815), .ZN(n4509) );
  OR2_X1 U5239 ( .A1(n8392), .A2(n4772), .ZN(n4512) );
  AND2_X1 U5240 ( .A1(n8392), .A2(n4772), .ZN(n4511) );
  INV_X1 U5241 ( .A(n4698), .ZN(n4694) );
  AND2_X1 U5242 ( .A1(n4947), .A2(n4646), .ZN(n4645) );
  NAND2_X1 U5243 ( .A1(n4647), .A2(n4648), .ZN(n4646) );
  NAND2_X1 U5244 ( .A1(n4682), .A2(n8559), .ZN(n4681) );
  NAND2_X1 U5245 ( .A1(n6388), .A2(n4955), .ZN(n4952) );
  OR2_X1 U5246 ( .A1(n9912), .A2(n8619), .ZN(n8207) );
  INV_X1 U5247 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n10067) );
  NOR2_X1 U5248 ( .A1(n6307), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n4460) );
  INV_X1 U5249 ( .A(n9869), .ZN(n6198) );
  NAND2_X1 U5250 ( .A1(n6199), .A2(n6198), .ZN(n8143) );
  NAND2_X1 U5251 ( .A1(n8143), .A2(n8144), .ZN(n8107) );
  INV_X1 U5252 ( .A(n8326), .ZN(n4689) );
  NAND2_X1 U5253 ( .A1(n9865), .A2(n6183), .ZN(n8148) );
  OR2_X1 U5254 ( .A1(n6642), .A2(n6556), .ZN(n6570) );
  NAND2_X1 U5255 ( .A1(n8263), .A2(n8264), .ZN(n4697) );
  AND2_X1 U5256 ( .A1(n6507), .A2(n8511), .ZN(n8252) );
  INV_X1 U5257 ( .A(n8508), .ZN(n4656) );
  INV_X1 U5258 ( .A(n8507), .ZN(n4654) );
  NAND2_X1 U5259 ( .A1(n8517), .A2(n4658), .ZN(n4657) );
  INV_X1 U5260 ( .A(n4662), .ZN(n4658) );
  AOI21_X1 U5261 ( .B1(n4665), .B2(n4664), .A(n4663), .ZN(n4662) );
  INV_X1 U5262 ( .A(n4973), .ZN(n4664) );
  INV_X1 U5263 ( .A(n7870), .ZN(n4974) );
  NAND2_X1 U5264 ( .A1(n4966), .A2(n6100), .ZN(n4965) );
  INV_X1 U5265 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n4966) );
  AND2_X1 U5266 ( .A1(n5147), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n5155) );
  NOR2_X1 U5267 ( .A1(n4605), .A2(n9241), .ZN(n4604) );
  INV_X1 U5268 ( .A(n4606), .ZN(n4605) );
  OR2_X1 U5269 ( .A1(n9788), .A2(n9775), .ZN(n5662) );
  AND2_X1 U5270 ( .A1(n5662), .A2(n5756), .ZN(n5599) );
  OR2_X1 U5271 ( .A1(n5440), .A2(n5439), .ZN(n5457) );
  OR2_X1 U5272 ( .A1(n9318), .A2(n9325), .ZN(n5712) );
  NAND2_X1 U5273 ( .A1(n4598), .A2(n7707), .ZN(n7712) );
  OAI21_X1 U5274 ( .B1(n5141), .B2(n10047), .A(n5101), .ZN(n5564) );
  NAND2_X1 U5275 ( .A1(n5171), .A2(n5170), .ZN(n5087) );
  AND2_X1 U5276 ( .A1(n5080), .A2(n5079), .ZN(n5218) );
  INV_X1 U5277 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5808) );
  AOI21_X1 U5278 ( .B1(n4885), .B2(n4883), .A(n4442), .ZN(n4882) );
  INV_X1 U5279 ( .A(n4885), .ZN(n4884) );
  INV_X1 U5280 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5573) );
  AOI21_X1 U5281 ( .B1(n4889), .B2(n5044), .A(n4888), .ZN(n4887) );
  INV_X1 U5282 ( .A(n5051), .ZN(n4888) );
  AND2_X1 U5283 ( .A1(n4890), .A2(n5046), .ZN(n4889) );
  INV_X1 U5284 ( .A(n5503), .ZN(n4890) );
  NAND2_X1 U5285 ( .A1(n5114), .A2(n5113), .ZN(n5504) );
  NAND2_X1 U5286 ( .A1(n4671), .A2(n4668), .ZN(n5480) );
  INV_X1 U5287 ( .A(n4669), .ZN(n4668) );
  OAI21_X1 U5288 ( .B1(n4677), .B2(n4670), .A(n4675), .ZN(n4669) );
  INV_X1 U5289 ( .A(n5432), .ZN(n5034) );
  NAND2_X1 U5290 ( .A1(n4591), .A2(n5026), .ZN(n5419) );
  XNOR2_X1 U5291 ( .A(n5025), .B(n10053), .ZN(n5403) );
  OR2_X1 U5292 ( .A1(n5382), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n5408) );
  OAI21_X1 U5293 ( .B1(n4555), .B2(n4471), .A(n4470), .ZN(n5010) );
  NAND2_X1 U5294 ( .A1(n4555), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n4470) );
  NAND2_X1 U5295 ( .A1(n5108), .A2(n5107), .ZN(n5319) );
  OR2_X1 U5296 ( .A1(n7987), .A2(n4733), .ZN(n4732) );
  INV_X1 U5297 ( .A(n7929), .ZN(n4733) );
  OR2_X1 U5298 ( .A1(n7894), .A2(n7893), .ZN(n4755) );
  NAND2_X1 U5299 ( .A1(n7236), .A2(n7230), .ZN(n4759) );
  INV_X1 U5300 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n10128) );
  AOI21_X1 U5301 ( .B1(n4739), .B2(n4738), .A(n4407), .ZN(n4737) );
  INV_X1 U5302 ( .A(n4744), .ZN(n4738) );
  NOR2_X1 U5303 ( .A1(n4378), .A2(n7957), .ZN(n4750) );
  AOI21_X1 U5304 ( .B1(n4378), .B2(n7893), .A(n4754), .ZN(n4753) );
  INV_X1 U5305 ( .A(n8037), .ZN(n4754) );
  AND3_X1 U5306 ( .A1(n6150), .A2(n6149), .A3(n6148), .ZN(n6418) );
  AND2_X1 U5307 ( .A1(n6417), .A2(n6416), .ZN(n8030) );
  NAND2_X1 U5308 ( .A1(n7126), .A2(n4489), .ZN(n6917) );
  NOR2_X1 U5309 ( .A1(n6987), .A2(n6986), .ZN(n7060) );
  NAND2_X1 U5310 ( .A1(n4779), .A2(n4778), .ZN(n7277) );
  INV_X1 U5311 ( .A(n7099), .ZN(n4778) );
  NOR2_X1 U5312 ( .A1(n8342), .A2(n8343), .ZN(n9821) );
  NOR2_X1 U5313 ( .A1(n8356), .A2(n8674), .ZN(n8393) );
  INV_X1 U5314 ( .A(n4481), .ZN(n8364) );
  XNOR2_X1 U5315 ( .A(n4454), .B(n8367), .ZN(n9854) );
  XNOR2_X1 U5316 ( .A(n8396), .B(n9847), .ZN(n9849) );
  INV_X1 U5317 ( .A(n4454), .ZN(n8368) );
  NAND2_X1 U5318 ( .A1(n4463), .A2(n10055), .ZN(n6431) );
  AND4_X1 U5319 ( .A1(n6155), .A2(n6154), .A3(n6153), .A4(n6152), .ZN(n8547)
         );
  OR2_X1 U5320 ( .A1(n6346), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n6359) );
  NAND2_X1 U5321 ( .A1(n4460), .A2(n10067), .ZN(n6334) );
  NAND2_X1 U5322 ( .A1(n4961), .A2(n4440), .ZN(n4960) );
  NAND2_X1 U5323 ( .A1(n9902), .A2(n7852), .ZN(n4962) );
  NAND2_X1 U5324 ( .A1(n4960), .A2(n4958), .ZN(n7751) );
  NOR2_X1 U5325 ( .A1(n8206), .A2(n4959), .ZN(n4958) );
  INV_X1 U5326 ( .A(n4962), .ZN(n4959) );
  OAI21_X1 U5327 ( .B1(n7454), .B2(n6495), .A(n8187), .ZN(n7559) );
  NAND2_X1 U5328 ( .A1(n4724), .A2(n8120), .ZN(n7561) );
  INV_X1 U5329 ( .A(n7559), .ZN(n4724) );
  NAND2_X1 U5330 ( .A1(n7484), .A2(n4967), .ZN(n7609) );
  NOR2_X1 U5331 ( .A1(n8179), .A2(n4968), .ZN(n4967) );
  INV_X1 U5332 ( .A(n6255), .ZN(n4968) );
  NAND2_X1 U5333 ( .A1(n4456), .A2(n4455), .ZN(n6256) );
  INV_X1 U5334 ( .A(n6241), .ZN(n4456) );
  NAND2_X1 U5335 ( .A1(n6805), .A2(n8110), .ZN(n4979) );
  NAND2_X1 U5336 ( .A1(n7206), .A2(n7205), .ZN(n7293) );
  AND2_X1 U5337 ( .A1(n7204), .A2(n7203), .ZN(n7205) );
  NAND2_X1 U5338 ( .A1(n6543), .A2(n6645), .ZN(n7202) );
  OR2_X1 U5339 ( .A1(n6642), .A2(P2_D_REG_1__SCAN_IN), .ZN(n6543) );
  OR2_X1 U5340 ( .A1(n6528), .A2(n9870), .ZN(n4985) );
  NOR2_X1 U5341 ( .A1(n8451), .A2(n8103), .ZN(n4698) );
  AND2_X1 U5342 ( .A1(n6471), .A2(n6470), .ZN(n8454) );
  OR2_X1 U5343 ( .A1(n8263), .A2(n8103), .ZN(n8462) );
  NAND2_X1 U5344 ( .A1(n8473), .A2(n8479), .ZN(n8472) );
  INV_X1 U5345 ( .A(n4703), .ZN(n4702) );
  AND2_X1 U5346 ( .A1(n4704), .A2(n8236), .ZN(n4703) );
  INV_X1 U5347 ( .A(n8252), .ZN(n4704) );
  AND2_X1 U5348 ( .A1(n6144), .A2(n6143), .ZN(n8486) );
  AND2_X1 U5349 ( .A1(n8254), .A2(n8104), .ZN(n8492) );
  AOI22_X1 U5350 ( .A1(n8497), .A2(n6426), .B1(n8485), .B2(n6507), .ZN(n8483)
         );
  OR2_X1 U5351 ( .A1(n8721), .A2(n6418), .ZN(n8236) );
  NAND2_X1 U5352 ( .A1(n8506), .A2(n8250), .ZN(n4705) );
  AND2_X1 U5353 ( .A1(n6504), .A2(n4714), .ZN(n4713) );
  NAND2_X1 U5354 ( .A1(n4974), .A2(n4973), .ZN(n4666) );
  NAND2_X1 U5355 ( .A1(n4666), .A2(n4665), .ZN(n8534) );
  OR2_X1 U5356 ( .A1(n7975), .A2(n8547), .ZN(n8531) );
  NAND2_X1 U5357 ( .A1(n4718), .A2(n4717), .ZN(n4716) );
  AOI21_X1 U5358 ( .B1(n8571), .B2(n6501), .A(n6500), .ZN(n8558) );
  AND4_X1 U5359 ( .A1(n6374), .A2(n6373), .A3(n6372), .A4(n6371), .ZN(n8578)
         );
  AND4_X1 U5360 ( .A1(n6364), .A2(n6363), .A3(n6362), .A4(n6361), .ZN(n8608)
         );
  NAND2_X1 U5361 ( .A1(n8289), .A2(n6520), .ZN(n8622) );
  INV_X1 U5362 ( .A(n8591), .ZN(n8620) );
  OR2_X1 U5363 ( .A1(n8757), .A2(n8608), .ZN(n8570) );
  AND2_X1 U5364 ( .A1(n7166), .A2(n8289), .ZN(n8591) );
  INV_X1 U5365 ( .A(n8622), .ZN(n8593) );
  AND2_X1 U5366 ( .A1(n6521), .A2(n4810), .ZN(n6247) );
  INV_X1 U5367 ( .A(n7745), .ZN(n6559) );
  NAND2_X1 U5368 ( .A1(n6545), .A2(n7745), .ZN(n6642) );
  AND2_X1 U5369 ( .A1(n6113), .A2(n4978), .ZN(n4977) );
  XNOR2_X1 U5370 ( .A(n6134), .B(P2_IR_REG_30__SCAN_IN), .ZN(n6135) );
  NAND2_X1 U5371 ( .A1(n8765), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6134) );
  AND2_X1 U5372 ( .A1(n6112), .A2(n4711), .ZN(n4710) );
  INV_X1 U5373 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n4711) );
  NAND2_X1 U5374 ( .A1(n6530), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6534) );
  INV_X1 U5375 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n6533) );
  NAND2_X1 U5376 ( .A1(n6534), .A2(n6533), .ZN(n6535) );
  XNOR2_X1 U5377 ( .A(n6485), .B(P2_IR_REG_21__SCAN_IN), .ZN(n8151) );
  NAND2_X1 U5378 ( .A1(n6482), .A2(n4764), .ZN(n6487) );
  AND2_X1 U5379 ( .A1(n6250), .A2(n4972), .ZN(n6375) );
  AND2_X1 U5380 ( .A1(n6074), .A2(n6073), .ZN(n5820) );
  INV_X1 U5381 ( .A(n7703), .ZN(n5821) );
  INV_X1 U5382 ( .A(n5155), .ZN(n5167) );
  NOR2_X1 U5383 ( .A1(n5970), .A2(n4853), .ZN(n4852) );
  INV_X1 U5384 ( .A(n5955), .ZN(n4853) );
  OR2_X1 U5385 ( .A1(n5525), .A2(n5524), .ZN(n5548) );
  INV_X1 U5386 ( .A(n4846), .ZN(n4548) );
  AND2_X1 U5387 ( .A1(n4845), .A2(n4551), .ZN(n4550) );
  NAND2_X1 U5388 ( .A1(n4846), .A2(n5952), .ZN(n4551) );
  AND2_X1 U5389 ( .A1(n4824), .A2(n4822), .ZN(n4821) );
  INV_X1 U5390 ( .A(n6014), .ZN(n4822) );
  NAND2_X1 U5391 ( .A1(n5888), .A2(n6829), .ZN(n7029) );
  INV_X1 U5392 ( .A(n5834), .ZN(n5829) );
  AND2_X1 U5393 ( .A1(n9570), .A2(n9014), .ZN(n9592) );
  AOI21_X1 U5394 ( .B1(P1_REG2_REG_4__SCAN_IN), .B2(n9013), .A(n9573), .ZN(
        n9587) );
  AOI21_X1 U5395 ( .B1(P1_REG1_REG_14__SCAN_IN), .B2(n9659), .A(n9660), .ZN(
        n9039) );
  AOI21_X1 U5396 ( .B1(P1_REG2_REG_14__SCAN_IN), .B2(n9659), .A(n9665), .ZN(
        n9050) );
  AND2_X1 U5397 ( .A1(n9696), .A2(n9053), .ZN(n9054) );
  NAND2_X1 U5398 ( .A1(n5143), .A2(n5142), .ZN(n9316) );
  NAND2_X1 U5399 ( .A1(n4607), .A2(n9445), .ZN(n9153) );
  OR2_X1 U5400 ( .A1(n9117), .A2(n9116), .ZN(n4800) );
  NAND2_X1 U5401 ( .A1(n5777), .A2(n9161), .ZN(n4799) );
  AND2_X1 U5402 ( .A1(n9185), .A2(n9334), .ZN(n9116) );
  NAND2_X1 U5403 ( .A1(n5584), .A2(n5777), .ZN(n9161) );
  OR2_X1 U5404 ( .A1(n9201), .A2(n9360), .ZN(n9176) );
  NAND2_X1 U5405 ( .A1(n4574), .A2(n4572), .ZN(n4570) );
  INV_X1 U5406 ( .A(n4572), .ZN(n4571) );
  AND2_X1 U5407 ( .A1(n9176), .A2(n5700), .ZN(n9194) );
  AND2_X1 U5408 ( .A1(n9233), .A2(n9378), .ZN(n4916) );
  AND2_X1 U5409 ( .A1(n5696), .A2(n9192), .ZN(n9211) );
  NAND2_X1 U5410 ( .A1(n9380), .A2(n9255), .ZN(n4918) );
  OAI22_X1 U5411 ( .A1(n9100), .A2(n9099), .B1(n9277), .B2(n9400), .ZN(n9267)
         );
  AND2_X1 U5412 ( .A1(n4561), .A2(n4560), .ZN(n9098) );
  NAND2_X1 U5413 ( .A1(n8861), .A2(n9406), .ZN(n4560) );
  NOR2_X1 U5414 ( .A1(n5491), .A2(n4787), .ZN(n4786) );
  INV_X1 U5415 ( .A(n4906), .ZN(n4901) );
  INV_X1 U5416 ( .A(n4902), .ZN(n4903) );
  AND2_X1 U5417 ( .A1(n5765), .A2(n5651), .ZN(n7721) );
  NAND2_X1 U5418 ( .A1(n4908), .A2(n4910), .ZN(n4907) );
  NAND2_X1 U5419 ( .A1(n4909), .A2(n7708), .ZN(n4908) );
  NAND2_X1 U5420 ( .A1(n7690), .A2(n4911), .ZN(n4909) );
  AND2_X1 U5421 ( .A1(n4910), .A2(n4911), .ZN(n4906) );
  AND2_X1 U5422 ( .A1(n5664), .A2(n5762), .ZN(n7719) );
  OR2_X1 U5423 ( .A1(n9780), .A2(n8955), .ZN(n4911) );
  INV_X1 U5424 ( .A(n5596), .ZN(n7623) );
  NAND2_X1 U5425 ( .A1(n4425), .A2(n4938), .ZN(n4927) );
  NAND2_X1 U5426 ( .A1(n4934), .A2(n4935), .ZN(n4933) );
  INV_X1 U5427 ( .A(n4936), .ZN(n4934) );
  NAND2_X1 U5428 ( .A1(n7437), .A2(n9746), .ZN(n4936) );
  NAND2_X1 U5429 ( .A1(n7303), .A2(n7302), .ZN(n7436) );
  NAND2_X1 U5430 ( .A1(n7262), .A2(n7305), .ZN(n7303) );
  OAI211_X1 U5431 ( .C1(n6773), .C2(n4915), .A(n4912), .B(n6792), .ZN(n7261)
         );
  NOR2_X1 U5432 ( .A1(n4915), .A2(n4914), .ZN(n4913) );
  INV_X1 U5433 ( .A(n6771), .ZN(n4914) );
  NAND2_X1 U5434 ( .A1(n6774), .A2(n6773), .ZN(n6790) );
  AOI21_X1 U5435 ( .B1(n9717), .B2(n6692), .A(n6691), .ZN(n6849) );
  INV_X1 U5436 ( .A(n4478), .ZN(n4477) );
  NAND2_X1 U5437 ( .A1(n9138), .A2(n4480), .ZN(n4479) );
  AOI22_X1 U5438 ( .A1(n9166), .A2(n9754), .B1(n9757), .B2(n9140), .ZN(n4478)
         );
  AND2_X1 U5439 ( .A1(n9316), .A2(n9787), .ZN(n4788) );
  OR2_X1 U5440 ( .A1(n9147), .A2(n9108), .ZN(n4922) );
  AND2_X1 U5441 ( .A1(n5429), .A2(n5428), .ZN(n9777) );
  NAND2_X1 U5442 ( .A1(n6084), .A2(n9564), .ZN(n9776) );
  INV_X1 U5443 ( .A(n9757), .ZN(n9774) );
  INV_X1 U5444 ( .A(n9776), .ZN(n9754) );
  OAI21_X1 U5445 ( .B1(n6687), .B2(P1_D_REG_0__SCAN_IN), .A(n9469), .ZN(n6854)
         );
  AOI21_X1 U5446 ( .B1(n4379), .B2(n4875), .A(n4867), .ZN(n4866) );
  INV_X1 U5447 ( .A(n5065), .ZN(n4867) );
  AND2_X1 U5448 ( .A1(n5070), .A2(n5069), .ZN(n5193) );
  NAND2_X1 U5449 ( .A1(n4869), .A2(n4873), .ZN(n5206) );
  NAND2_X1 U5450 ( .A1(n4871), .A2(n4870), .ZN(n4869) );
  NAND2_X1 U5451 ( .A1(n5108), .A2(n4940), .ZN(n4941) );
  NOR2_X1 U5452 ( .A1(n5110), .A2(P1_IR_REG_3__SCAN_IN), .ZN(n4940) );
  NAND2_X1 U5453 ( .A1(n5008), .A2(n5007), .ZN(n5351) );
  INV_X1 U5454 ( .A(n7191), .ZN(n7192) );
  NAND2_X1 U5455 ( .A1(n7178), .A2(n7180), .ZN(n7399) );
  NAND2_X1 U5456 ( .A1(n7926), .A2(n7925), .ZN(n7986) );
  INV_X1 U5457 ( .A(n8709), .ZN(n8024) );
  INV_X1 U5458 ( .A(n8317), .ZN(n7788) );
  INV_X1 U5459 ( .A(n9902), .ZN(n7801) );
  AND2_X1 U5460 ( .A1(n6460), .A2(n6459), .ZN(n8072) );
  AND2_X1 U5461 ( .A1(n7189), .A2(n7188), .ZN(n8084) );
  NAND2_X1 U5462 ( .A1(n4540), .A2(n4368), .ZN(n4538) );
  NAND2_X1 U5463 ( .A1(n8297), .A2(n4541), .ZN(n4540) );
  XNOR2_X1 U5464 ( .A(n6484), .B(P2_IR_REG_22__SCAN_IN), .ZN(n8305) );
  NAND2_X1 U5465 ( .A1(n6529), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6484) );
  NAND2_X1 U5466 ( .A1(n6482), .A2(n4389), .ZN(n6529) );
  INV_X1 U5467 ( .A(n8072), .ZN(n8465) );
  NAND2_X1 U5468 ( .A1(n6447), .A2(n6446), .ZN(n8474) );
  INV_X1 U5469 ( .A(n8486), .ZN(n8464) );
  INV_X1 U5470 ( .A(n8030), .ZN(n8538) );
  NAND4_X1 U5471 ( .A1(n6220), .A2(n6219), .A3(n6218), .A4(n6217), .ZN(n8323)
         );
  NAND4_X1 U5472 ( .A1(n6207), .A2(n6206), .A3(n6205), .A4(n6204), .ZN(n8324)
         );
  NAND2_X1 U5473 ( .A1(n6170), .A2(n10069), .ZN(n6206) );
  NOR2_X1 U5474 ( .A1(n8597), .A2(n8344), .ZN(n8365) );
  OAI21_X1 U5475 ( .B1(n4630), .B2(n4629), .A(n4628), .ZN(n4627) );
  NOR2_X1 U5476 ( .A1(n4633), .A2(n4632), .ZN(n4629) );
  NAND2_X1 U5477 ( .A1(n4630), .A2(n8417), .ZN(n4628) );
  INV_X1 U5478 ( .A(n4631), .ZN(n4630) );
  OAI21_X1 U5479 ( .B1(n8400), .B2(n8398), .A(n8416), .ZN(n4498) );
  INV_X1 U5480 ( .A(n4499), .ZN(n4497) );
  NAND2_X1 U5481 ( .A1(n6878), .A2(n6888), .ZN(n9856) );
  NAND2_X1 U5482 ( .A1(n6464), .A2(n6463), .ZN(n8687) );
  XNOR2_X1 U5483 ( .A(n6159), .B(n6481), .ZN(n8421) );
  INV_X1 U5484 ( .A(n8781), .ZN(n4553) );
  INV_X1 U5485 ( .A(n8780), .ZN(n4552) );
  INV_X1 U5486 ( .A(n7437), .ZN(n4596) );
  OAI21_X1 U5487 ( .B1(n8889), .B2(n5997), .A(n6000), .ZN(n8828) );
  AND3_X1 U5488 ( .A1(n5477), .A2(n5476), .A3(n5475), .ZN(n8939) );
  NOR2_X1 U5489 ( .A1(n5828), .A2(n4880), .ZN(n4879) );
  NOR2_X1 U5490 ( .A1(n5796), .A2(n6839), .ZN(n4880) );
  INV_X1 U5491 ( .A(n9324), .ZN(n9345) );
  NAND4_X1 U5492 ( .A1(n5293), .A2(n5292), .A3(n5291), .A4(n5290), .ZN(n8962)
         );
  NAND2_X1 U5493 ( .A1(n8983), .A2(n8984), .ZN(n9011) );
  INV_X1 U5494 ( .A(n9078), .ZN(n4474) );
  NAND2_X1 U5495 ( .A1(n4791), .A2(n4789), .ZN(n9314) );
  INV_X1 U5496 ( .A(n4790), .ZN(n4789) );
  NAND2_X1 U5497 ( .A1(n4792), .A2(n9765), .ZN(n4791) );
  OAI22_X1 U5498 ( .A1(n9325), .A2(n9776), .B1(n9122), .B2(n9121), .ZN(n4790)
         );
  AOI21_X1 U5499 ( .B1(n4921), .B2(n9108), .A(n4405), .ZN(n4920) );
  AND2_X1 U5500 ( .A1(n5215), .A2(n5214), .ZN(n9361) );
  AND2_X1 U5501 ( .A1(n5502), .A2(n5501), .ZN(n7824) );
  NAND2_X1 U5502 ( .A1(n9265), .A2(n6713), .ZN(n9273) );
  INV_X2 U5503 ( .A(n9265), .ZN(n9293) );
  OR2_X1 U5504 ( .A1(n6686), .A2(n6846), .ZN(n9242) );
  NAND2_X1 U5505 ( .A1(n4578), .A2(n4584), .ZN(n4580) );
  NAND2_X1 U5506 ( .A1(n9132), .A2(n9794), .ZN(n4584) );
  NAND2_X1 U5507 ( .A1(n4922), .A2(n4585), .ZN(n4578) );
  AND2_X1 U5508 ( .A1(n9107), .A2(n9794), .ZN(n4585) );
  NAND2_X1 U5509 ( .A1(n4922), .A2(n4921), .ZN(n9131) );
  NOR2_X1 U5510 ( .A1(n4806), .A2(n5121), .ZN(n4805) );
  NAND2_X1 U5511 ( .A1(n8194), .A2(n4513), .ZN(n8203) );
  OAI211_X1 U5512 ( .C1(n8176), .C2(n8284), .A(n4515), .B(n4514), .ZN(n4513)
         );
  NAND2_X1 U5513 ( .A1(n4530), .A2(n8209), .ZN(n8211) );
  AOI21_X1 U5514 ( .B1(n4453), .B2(n5263), .A(n5695), .ZN(n5698) );
  NAND2_X1 U5515 ( .A1(n4377), .A2(n8233), .ZN(n4520) );
  NAND2_X1 U5516 ( .A1(n4859), .A2(n4856), .ZN(n5711) );
  NAND2_X1 U5517 ( .A1(n4857), .A2(n6840), .ZN(n4856) );
  INV_X1 U5518 ( .A(n5672), .ZN(n5770) );
  INV_X1 U5519 ( .A(n5446), .ZN(n5035) );
  INV_X1 U5520 ( .A(SI_13_), .ZN(n10071) );
  INV_X1 U5521 ( .A(n8520), .ZN(n4663) );
  NOR2_X1 U5522 ( .A1(n5975), .A2(n4850), .ZN(n4849) );
  INV_X1 U5523 ( .A(n5969), .ZN(n4850) );
  NOR2_X1 U5524 ( .A1(n5391), .A2(n7645), .ZN(n5367) );
  NAND2_X1 U5525 ( .A1(n5831), .A2(n7383), .ZN(n5833) );
  AOI21_X1 U5526 ( .B1(n9178), .B2(n4797), .A(n4795), .ZN(n4794) );
  NOR2_X1 U5527 ( .A1(n4798), .A2(n9145), .ZN(n4797) );
  OAI21_X1 U5528 ( .B1(n4796), .B2(n9145), .A(n9118), .ZN(n4795) );
  NOR2_X1 U5529 ( .A1(n9388), .A2(n9392), .ZN(n4606) );
  NAND2_X1 U5530 ( .A1(n5151), .A2(n5152), .ZN(n5097) );
  AND2_X1 U5531 ( .A1(n4887), .A2(n5515), .ZN(n4885) );
  INV_X1 U5532 ( .A(n4889), .ZN(n4883) );
  INV_X1 U5533 ( .A(n5492), .ZN(n5045) );
  AOI21_X1 U5534 ( .B1(n4413), .B2(n4678), .A(n4676), .ZN(n4675) );
  INV_X1 U5535 ( .A(n5039), .ZN(n4676) );
  NAND2_X1 U5536 ( .A1(n4678), .A2(n5038), .ZN(n4677) );
  NAND2_X1 U5537 ( .A1(n5418), .A2(n5030), .ZN(n4670) );
  NOR2_X1 U5538 ( .A1(n4677), .A2(n4673), .ZN(n4672) );
  INV_X1 U5539 ( .A(n5030), .ZN(n4673) );
  NOR2_X1 U5540 ( .A1(n5024), .A2(n4593), .ZN(n4592) );
  INV_X1 U5541 ( .A(n5022), .ZN(n4593) );
  INV_X1 U5542 ( .A(n5403), .ZN(n5024) );
  OAI21_X1 U5543 ( .B1(n5009), .B2(n4864), .A(n5380), .ZN(n4863) );
  INV_X1 U5544 ( .A(n5011), .ZN(n4864) );
  OAI21_X1 U5545 ( .B1(n4376), .B2(n4641), .A(n4640), .ZN(n4989) );
  NAND2_X1 U5546 ( .A1(n4375), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n4640) );
  INV_X1 U5547 ( .A(SI_8_), .ZN(n10078) );
  INV_X1 U5548 ( .A(SI_11_), .ZN(n10132) );
  INV_X1 U5549 ( .A(SI_22_), .ZN(n10103) );
  NOR2_X1 U5550 ( .A1(n6379), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n4461) );
  OR2_X1 U5551 ( .A1(n8280), .A2(n8278), .ZN(n4532) );
  NAND2_X1 U5552 ( .A1(n6194), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6894) );
  AND2_X1 U5553 ( .A1(n6882), .A2(n4488), .ZN(n4623) );
  NAND2_X1 U5554 ( .A1(n4621), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n4620) );
  NAND2_X1 U5555 ( .A1(n7019), .A2(n6994), .ZN(n6996) );
  NOR2_X1 U5556 ( .A1(n6989), .A2(n6988), .ZN(n4464) );
  AND2_X1 U5557 ( .A1(n7581), .A2(n7580), .ZN(n8350) );
  NAND2_X1 U5558 ( .A1(n9828), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n4772) );
  NAND2_X1 U5559 ( .A1(n9843), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n4612) );
  AND2_X1 U5560 ( .A1(n4771), .A2(n4770), .ZN(n8396) );
  NAND2_X1 U5561 ( .A1(n9843), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n4770) );
  AND2_X1 U5562 ( .A1(n8445), .A2(n4948), .ZN(n4947) );
  NAND2_X1 U5563 ( .A1(n6462), .A2(n4949), .ZN(n4948) );
  INV_X1 U5564 ( .A(n6461), .ZN(n4949) );
  INV_X1 U5565 ( .A(n6462), .ZN(n4950) );
  NOR2_X1 U5566 ( .A1(n6421), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n4463) );
  NOR2_X1 U5567 ( .A1(n6404), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n4462) );
  INV_X1 U5568 ( .A(n4461), .ZN(n6381) );
  NAND2_X1 U5569 ( .A1(n6127), .A2(n10198), .ZN(n6379) );
  INV_X1 U5570 ( .A(n6359), .ZN(n6127) );
  AND2_X1 U5571 ( .A1(n8207), .A2(n8208), .ZN(n8206) );
  OR2_X1 U5572 ( .A1(n6299), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n6307) );
  INV_X1 U5573 ( .A(n8183), .ZN(n4723) );
  OR2_X1 U5574 ( .A1(n7801), .A2(n7852), .ZN(n8199) );
  NAND2_X1 U5575 ( .A1(n4381), .A2(n4651), .ZN(n4648) );
  NAND2_X1 U5576 ( .A1(n4649), .A2(n4381), .ZN(n4647) );
  AND2_X1 U5577 ( .A1(n8104), .A2(n8489), .ZN(n8253) );
  NAND2_X1 U5578 ( .A1(n4703), .A2(n4701), .ZN(n4700) );
  INV_X1 U5579 ( .A(n8250), .ZN(n4701) );
  OR2_X1 U5580 ( .A1(n8727), .A2(n8030), .ZN(n8248) );
  NAND2_X1 U5581 ( .A1(n8231), .A2(n4715), .ZN(n4714) );
  NOR2_X1 U5582 ( .A1(n6573), .A2(n6557), .ZN(n7155) );
  INV_X1 U5583 ( .A(n4837), .ZN(n4831) );
  INV_X1 U5584 ( .A(n4836), .ZN(n4834) );
  AND2_X1 U5585 ( .A1(n4838), .A2(n7032), .ZN(n4837) );
  NAND2_X1 U5586 ( .A1(n7252), .A2(n7253), .ZN(n4838) );
  NOR2_X1 U5587 ( .A1(n7252), .A2(n7253), .ZN(n4836) );
  INV_X1 U5588 ( .A(n5862), .ZN(n5880) );
  AND2_X1 U5589 ( .A1(n5843), .A2(n5842), .ZN(n5849) );
  INV_X1 U5590 ( .A(n4825), .ZN(n4824) );
  OAI21_X1 U5591 ( .B1(n8829), .B2(n4826), .A(n6007), .ZN(n4825) );
  NAND2_X1 U5592 ( .A1(n5997), .A2(n6000), .ZN(n4826) );
  INV_X1 U5593 ( .A(n4849), .ZN(n4848) );
  OR2_X1 U5594 ( .A1(n5721), .A2(n9121), .ZN(n5583) );
  AND2_X1 U5595 ( .A1(P1_REG3_REG_24__SCAN_IN), .A2(n5186), .ZN(n5188) );
  NOR2_X1 U5596 ( .A1(n5210), .A2(n8800), .ZN(n5186) );
  AND2_X1 U5597 ( .A1(n5687), .A2(n5681), .ZN(n5602) );
  INV_X1 U5598 ( .A(n4786), .ZN(n4782) );
  INV_X1 U5599 ( .A(n7514), .ZN(n4926) );
  OR2_X1 U5600 ( .A1(n9139), .A2(n5608), .ZN(n4480) );
  NAND2_X1 U5601 ( .A1(n9268), .A2(n4606), .ZN(n9257) );
  AND2_X1 U5602 ( .A1(n6767), .A2(n5738), .ZN(n6702) );
  AND2_X1 U5603 ( .A1(n5092), .A2(n5091), .ZN(n5161) );
  AND2_X1 U5604 ( .A1(n5086), .A2(n5085), .ZN(n5170) );
  AND2_X1 U5605 ( .A1(n5075), .A2(n5074), .ZN(n5180) );
  XNOR2_X1 U5606 ( .A(n5798), .B(P1_IR_REG_23__SCAN_IN), .ZN(n6621) );
  INV_X1 U5607 ( .A(n4874), .ZN(n4873) );
  OAI21_X1 U5608 ( .B1(n4877), .B2(n4875), .A(n5061), .ZN(n4874) );
  INV_X1 U5609 ( .A(n5245), .ZN(n4871) );
  NAND2_X1 U5610 ( .A1(n5320), .A2(n5109), .ZN(n5110) );
  INV_X1 U5611 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n5109) );
  INV_X1 U5612 ( .A(SI_14_), .ZN(n10058) );
  NAND2_X1 U5613 ( .A1(n5433), .A2(n4679), .ZN(n4674) );
  XNOR2_X1 U5614 ( .A(n5032), .B(n5031), .ZN(n5432) );
  OAI21_X1 U5615 ( .B1(n4555), .B2(n4996), .A(n4995), .ZN(n4998) );
  NAND2_X1 U5616 ( .A1(n4376), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n4995) );
  NAND2_X1 U5617 ( .A1(n7535), .A2(n7534), .ZN(n7591) );
  INV_X1 U5618 ( .A(n7922), .ZN(n8016) );
  NAND2_X1 U5619 ( .A1(n8049), .A2(n7919), .ZN(n8015) );
  INV_X1 U5620 ( .A(n8058), .ZN(n4741) );
  INV_X1 U5621 ( .A(n7970), .ZN(n4736) );
  NAND2_X1 U5622 ( .A1(n7771), .A2(n7770), .ZN(n7787) );
  NAND2_X1 U5623 ( .A1(n4461), .A2(n6128), .ZN(n6393) );
  NOR2_X1 U5624 ( .A1(n4746), .A2(n4745), .ZN(n4744) );
  INV_X1 U5625 ( .A(n8002), .ZN(n4745) );
  NAND2_X1 U5626 ( .A1(n8003), .A2(n4747), .ZN(n4743) );
  AND2_X1 U5627 ( .A1(n7165), .A2(n7166), .ZN(n8078) );
  INV_X1 U5628 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n4763) );
  AND2_X1 U5629 ( .A1(n7356), .A2(n7355), .ZN(n8137) );
  NAND2_X1 U5630 ( .A1(n6194), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6881) );
  NAND2_X1 U5631 ( .A1(n8334), .A2(n4766), .ZN(n8333) );
  NAND2_X1 U5632 ( .A1(n7132), .A2(n4621), .ZN(n6919) );
  NAND3_X1 U5633 ( .A1(n4484), .A2(n4486), .A3(n6915), .ZN(n7126) );
  OR2_X1 U5634 ( .A1(n6917), .A2(n6203), .ZN(n7128) );
  NAND2_X1 U5635 ( .A1(n4619), .A2(n7132), .ZN(n7134) );
  INV_X1 U5636 ( .A(n4620), .ZN(n4619) );
  OR2_X1 U5637 ( .A1(n6231), .A2(n6902), .ZN(n7009) );
  OAI21_X1 U5638 ( .B1(n6996), .B2(n6995), .A(n7000), .ZN(n7047) );
  INV_X1 U5639 ( .A(n6999), .ZN(n7046) );
  NOR2_X1 U5640 ( .A1(n7050), .A2(n4505), .ZN(n6987) );
  INV_X1 U5641 ( .A(n4504), .ZN(n4505) );
  NAND2_X1 U5642 ( .A1(n4502), .A2(n4393), .ZN(n4779) );
  INV_X1 U5643 ( .A(n4777), .ZN(n7364) );
  NAND2_X1 U5644 ( .A1(n4501), .A2(n4500), .ZN(n7581) );
  INV_X1 U5645 ( .A(n7565), .ZN(n4617) );
  OR2_X1 U5646 ( .A1(n7374), .A2(n7373), .ZN(n7566) );
  NOR2_X1 U5647 ( .A1(n8354), .A2(n6348), .ZN(n4482) );
  OAI211_X1 U5648 ( .C1(n4775), .C2(n4510), .A(n4508), .B(n4506), .ZN(n8356)
         );
  INV_X1 U5649 ( .A(n4511), .ZN(n4510) );
  AND2_X1 U5650 ( .A1(n4509), .A2(n4512), .ZN(n4508) );
  NOR2_X1 U5651 ( .A1(n9849), .A2(n9850), .ZN(n9848) );
  INV_X1 U5652 ( .A(n8371), .ZN(n4632) );
  AOI21_X1 U5653 ( .B1(n8369), .B2(n4632), .A(n8406), .ZN(n4631) );
  AOI21_X1 U5654 ( .B1(n4693), .B2(n4696), .A(n4409), .ZN(n4691) );
  AOI21_X1 U5655 ( .B1(n4694), .B2(n4695), .A(n8445), .ZN(n4693) );
  INV_X1 U5656 ( .A(n6474), .ZN(n7943) );
  OR2_X1 U5657 ( .A1(n6465), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n6474) );
  INV_X1 U5658 ( .A(n4463), .ZN(n6429) );
  OR2_X1 U5659 ( .A1(n6415), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6421) );
  NAND2_X1 U5660 ( .A1(n4462), .A2(n10126), .ZN(n6415) );
  INV_X1 U5661 ( .A(n4462), .ZN(n6413) );
  OR2_X1 U5662 ( .A1(n6393), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n6395) );
  NAND2_X1 U5663 ( .A1(n6129), .A2(n10045), .ZN(n6404) );
  INV_X1 U5664 ( .A(n6395), .ZN(n6129) );
  NAND2_X1 U5665 ( .A1(n4953), .A2(n4951), .ZN(n8545) );
  NAND2_X1 U5666 ( .A1(n4388), .A2(n4952), .ZN(n4951) );
  NAND3_X1 U5667 ( .A1(n4388), .A2(n8616), .A3(n4956), .ZN(n4953) );
  OAI21_X1 U5668 ( .B1(n8628), .B2(n6497), .A(n6498), .ZN(n8613) );
  NAND2_X1 U5669 ( .A1(n6126), .A2(n6125), .ZN(n6346) );
  INV_X1 U5670 ( .A(n6334), .ZN(n6126) );
  INV_X1 U5671 ( .A(n4460), .ZN(n6323) );
  AND4_X1 U5672 ( .A1(n6328), .A2(n6327), .A3(n6326), .A4(n6325), .ZN(n8619)
         );
  AND2_X1 U5673 ( .A1(n8199), .A2(n8197), .ZN(n8119) );
  NAND2_X1 U5674 ( .A1(n4457), .A2(n6124), .ZN(n6299) );
  INV_X1 U5675 ( .A(n6281), .ZN(n4457) );
  NAND2_X1 U5676 ( .A1(n4459), .A2(n4458), .ZN(n6281) );
  INV_X1 U5677 ( .A(n6269), .ZN(n4459) );
  AND2_X1 U5678 ( .A1(n6494), .A2(n6493), .ZN(n7454) );
  OAI21_X1 U5679 ( .B1(n7490), .B2(n4688), .A(n4685), .ZN(n7604) );
  INV_X1 U5680 ( .A(n8111), .ZN(n4688) );
  AOI21_X1 U5681 ( .B1(n8111), .B2(n4687), .A(n4686), .ZN(n4685) );
  INV_X1 U5682 ( .A(n8161), .ZN(n4687) );
  NAND2_X1 U5683 ( .A1(n7484), .A2(n6255), .ZN(n7607) );
  NAND2_X1 U5684 ( .A1(n6123), .A2(n6122), .ZN(n6269) );
  INV_X1 U5685 ( .A(n6256), .ZN(n6123) );
  AND2_X1 U5686 ( .A1(n8163), .A2(n8172), .ZN(n8114) );
  INV_X1 U5687 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n6120) );
  NAND2_X1 U5688 ( .A1(n7490), .A2(n8161), .ZN(n7323) );
  NAND2_X1 U5689 ( .A1(n7323), .A2(n8111), .ZN(n7479) );
  OAI21_X1 U5690 ( .B1(n7197), .B2(n8152), .A(n7198), .ZN(n7210) );
  AND2_X1 U5691 ( .A1(n8284), .A2(n6575), .ZN(n7201) );
  AND2_X1 U5692 ( .A1(n6573), .A2(n6572), .ZN(n7206) );
  NAND2_X1 U5693 ( .A1(n8093), .A2(n8092), .ZN(n8433) );
  NAND2_X1 U5694 ( .A1(n4652), .A2(n4653), .ZN(n8510) );
  NAND2_X1 U5695 ( .A1(n4974), .A2(n4655), .ZN(n4652) );
  NAND2_X1 U5696 ( .A1(n4659), .A2(n4657), .ZN(n8519) );
  NAND2_X1 U5697 ( .A1(n7870), .A2(n4660), .ZN(n4659) );
  AND2_X1 U5698 ( .A1(n6161), .A2(n6160), .ZN(n7891) );
  AOI21_X1 U5699 ( .B1(n8616), .B2(n4956), .A(n4954), .ZN(n8590) );
  AND3_X1 U5700 ( .A1(n6197), .A2(n6196), .A3(n6195), .ZN(n9869) );
  OR2_X1 U5701 ( .A1(n6521), .A2(n6895), .ZN(n6195) );
  NAND2_X1 U5702 ( .A1(n8149), .A2(n7207), .ZN(n9870) );
  NOR2_X1 U5703 ( .A1(n7157), .A2(n6565), .ZN(n7187) );
  INV_X1 U5704 ( .A(n7162), .ZN(n6565) );
  AND3_X1 U5705 ( .A1(n6180), .A2(n6179), .A3(n6178), .ZN(n9865) );
  OR2_X1 U5706 ( .A1(n6521), .A2(n6177), .ZN(n6178) );
  NOR2_X1 U5707 ( .A1(n7666), .A2(n9898), .ZN(n9908) );
  NAND2_X1 U5708 ( .A1(n8149), .A2(n8139), .ZN(n9901) );
  OR2_X1 U5709 ( .A1(n6330), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n6331) );
  INV_X1 U5710 ( .A(n4965), .ZN(n4684) );
  INV_X1 U5711 ( .A(n6621), .ZN(n6085) );
  NAND2_X1 U5712 ( .A1(n5834), .A2(n6080), .ZN(n5835) );
  NAND2_X1 U5713 ( .A1(n5956), .A2(n5955), .ZN(n8851) );
  AND2_X1 U5714 ( .A1(n5485), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n8870) );
  OR2_X1 U5715 ( .A1(n8791), .A2(n5952), .ZN(n5956) );
  AND2_X1 U5716 ( .A1(n5237), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n5236) );
  NAND2_X1 U5717 ( .A1(n5829), .A2(n5831), .ZN(n6699) );
  NOR2_X1 U5718 ( .A1(n5730), .A2(n7863), .ZN(n4467) );
  INV_X1 U5719 ( .A(n6080), .ZN(n6698) );
  AND3_X1 U5720 ( .A1(n5150), .A2(n5149), .A3(n5148), .ZN(n8951) );
  AOI21_X1 U5721 ( .B1(n9017), .B2(P1_REG1_REG_5__SCAN_IN), .A(n9590), .ZN(
        n9602) );
  AOI21_X1 U5722 ( .B1(P1_REG2_REG_6__SCAN_IN), .B2(n9019), .A(n9605), .ZN(
        n9506) );
  AOI21_X1 U5723 ( .B1(P1_REG2_REG_7__SCAN_IN), .B2(n9022), .A(n9505), .ZN(
        n9516) );
  AOI21_X1 U5724 ( .B1(n9022), .B2(P1_REG1_REG_7__SCAN_IN), .A(n9501), .ZN(
        n9520) );
  AOI21_X1 U5725 ( .B1(n9498), .B2(P1_REG1_REG_10__SCAN_IN), .A(n9490), .ZN(
        n9616) );
  AOI21_X1 U5726 ( .B1(P1_REG2_REG_10__SCAN_IN), .B2(n9498), .A(n9493), .ZN(
        n9620) );
  NAND2_X1 U5727 ( .A1(n9634), .A2(n9038), .ZN(n9650) );
  AOI21_X1 U5728 ( .B1(P1_REG2_REG_13__SCAN_IN), .B2(n9644), .A(n9645), .ZN(
        n9666) );
  AOI21_X1 U5729 ( .B1(n9644), .B2(P1_REG1_REG_13__SCAN_IN), .A(n9649), .ZN(
        n9662) );
  AND2_X1 U5730 ( .A1(n9066), .A2(n9065), .ZN(n9703) );
  NAND2_X1 U5731 ( .A1(n9348), .A2(n9334), .ZN(n4898) );
  NAND2_X1 U5732 ( .A1(n9200), .A2(n9348), .ZN(n9179) );
  AND2_X1 U5733 ( .A1(n5204), .A2(n5203), .ZN(n9199) );
  NOR2_X1 U5734 ( .A1(n9233), .A2(n4603), .ZN(n4602) );
  INV_X1 U5735 ( .A(n4604), .ZN(n4603) );
  AND2_X1 U5736 ( .A1(n9388), .A2(n9377), .ZN(n4564) );
  AND3_X1 U5737 ( .A1(n5529), .A2(n5528), .A3(n5527), .ZN(n9277) );
  INV_X1 U5738 ( .A(n4804), .ZN(n9280) );
  NAND2_X1 U5739 ( .A1(n9268), .A2(n9274), .ZN(n9269) );
  INV_X1 U5740 ( .A(n5602), .ZN(n9275) );
  NOR2_X1 U5741 ( .A1(n9096), .A2(n9397), .ZN(n4559) );
  NOR2_X1 U5742 ( .A1(n7712), .A2(n9427), .ZN(n7725) );
  NAND2_X1 U5743 ( .A1(n7725), .A2(n8949), .ZN(n7836) );
  INV_X1 U5744 ( .A(n5599), .ZN(n7708) );
  AND2_X1 U5745 ( .A1(n5443), .A2(n5442), .ZN(n7689) );
  NAND2_X1 U5746 ( .A1(n7269), .A2(n4382), .ZN(n7468) );
  NAND2_X1 U5747 ( .A1(n7269), .A2(n7425), .ZN(n7316) );
  NAND2_X1 U5748 ( .A1(n6772), .A2(n6771), .ZN(n6774) );
  NAND2_X1 U5749 ( .A1(n5617), .A2(n5619), .ZN(n6753) );
  INV_X1 U5750 ( .A(n6753), .ZN(n6748) );
  INV_X1 U5751 ( .A(n6934), .ZN(n6931) );
  NOR2_X1 U5752 ( .A1(n6595), .A2(n4810), .ZN(n4809) );
  NAND2_X1 U5753 ( .A1(n6581), .A2(n5837), .ZN(n6686) );
  AND2_X1 U5754 ( .A1(n5160), .A2(n5159), .ZN(n9325) );
  INV_X1 U5755 ( .A(n9300), .ZN(n9400) );
  AND3_X1 U5756 ( .A1(n5359), .A2(n5358), .A3(n5357), .ZN(n9733) );
  INV_X1 U5757 ( .A(n9768), .ZN(n9787) );
  AND2_X1 U5758 ( .A1(n5834), .A2(n7446), .ZN(n9720) );
  XNOR2_X1 U5759 ( .A(n5568), .B(n5567), .ZN(n8763) );
  XNOR2_X1 U5760 ( .A(n5564), .B(n5563), .ZN(n8768) );
  XNOR2_X1 U5761 ( .A(n5151), .B(n5152), .ZN(n7889) );
  NAND2_X1 U5762 ( .A1(n4807), .A2(n5113), .ZN(n4806) );
  AND2_X1 U5763 ( .A1(n5122), .A2(n5123), .ZN(n4807) );
  XNOR2_X1 U5764 ( .A(n5817), .B(P1_IR_REG_26__SCAN_IN), .ZN(n6074) );
  NAND2_X1 U5765 ( .A1(n5812), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5580) );
  NAND2_X1 U5766 ( .A1(n5580), .A2(n5808), .ZN(n5797) );
  XNOR2_X1 U5767 ( .A(n5582), .B(n5577), .ZN(n5830) );
  NAND2_X1 U5768 ( .A1(n5795), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5582) );
  NAND2_X1 U5769 ( .A1(n4872), .A2(n4876), .ZN(n5233) );
  NAND2_X1 U5770 ( .A1(n5505), .A2(n4854), .ZN(n4855) );
  NOR2_X1 U5771 ( .A1(n5575), .A2(P1_IR_REG_16__SCAN_IN), .ZN(n4854) );
  INV_X1 U5772 ( .A(n5504), .ZN(n5505) );
  INV_X1 U5773 ( .A(n5534), .ZN(n5533) );
  NAND2_X1 U5774 ( .A1(n4886), .A2(n4887), .ZN(n5516) );
  NAND2_X1 U5775 ( .A1(n5494), .A2(n4889), .ZN(n4886) );
  OR2_X1 U5776 ( .A1(n5408), .A2(n5407), .ZN(n5420) );
  NAND2_X1 U5777 ( .A1(n5023), .A2(n5022), .ZN(n5404) );
  AND2_X1 U5778 ( .A1(n5322), .A2(n5336), .ZN(n9013) );
  INV_X1 U5779 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n10198) );
  AOI21_X1 U5780 ( .B1(n4391), .B2(n4733), .A(n4729), .ZN(n4728) );
  INV_X1 U5781 ( .A(n8067), .ZN(n4729) );
  NAND2_X1 U5782 ( .A1(n4748), .A2(n4753), .ZN(n7958) );
  NAND2_X1 U5783 ( .A1(n7895), .A2(n4378), .ZN(n4748) );
  AND4_X1 U5784 ( .A1(n6409), .A2(n6408), .A3(n6407), .A4(n6406), .ZN(n8311)
         );
  AND2_X1 U5785 ( .A1(n6437), .A2(n6436), .ZN(n8018) );
  NAND2_X1 U5786 ( .A1(n4759), .A2(n7328), .ZN(n4756) );
  AOI21_X1 U5787 ( .B1(n8004), .B2(n8002), .A(n8003), .ZN(n8007) );
  INV_X1 U5788 ( .A(n4759), .ZN(n4758) );
  AND2_X1 U5789 ( .A1(n7231), .A2(n7230), .ZN(n7237) );
  NAND2_X1 U5790 ( .A1(n7653), .A2(n7652), .ZN(n7654) );
  AND4_X1 U5791 ( .A1(n6352), .A2(n6351), .A3(n6350), .A4(n6349), .ZN(n8621)
         );
  AOI21_X1 U5792 ( .B1(n7895), .B2(n7894), .A(n7893), .ZN(n8039) );
  NAND2_X1 U5793 ( .A1(n4725), .A2(n7180), .ZN(n7341) );
  INV_X1 U5794 ( .A(n8081), .ZN(n8009) );
  INV_X1 U5795 ( .A(n8084), .ZN(n8005) );
  NAND2_X1 U5796 ( .A1(n4742), .A2(n4743), .ZN(n8057) );
  NAND2_X1 U5797 ( .A1(n8004), .A2(n4744), .ZN(n4742) );
  NAND2_X1 U5798 ( .A1(n4731), .A2(n7929), .ZN(n8069) );
  NAND2_X1 U5799 ( .A1(n7986), .A2(n7987), .ZN(n4731) );
  NAND2_X1 U5800 ( .A1(n4753), .A2(n4752), .ZN(n4751) );
  AOI21_X1 U5801 ( .B1(n4750), .B2(n4753), .A(n4410), .ZN(n4749) );
  INV_X1 U5802 ( .A(n7957), .ZN(n4752) );
  AND4_X1 U5803 ( .A1(n6385), .A2(n6384), .A3(n6383), .A4(n6382), .ZN(n8082)
         );
  INV_X1 U5804 ( .A(n8137), .ZN(n8429) );
  OR2_X1 U5805 ( .A1(n6587), .A2(n7218), .ZN(n8383) );
  INV_X1 U5806 ( .A(n8018), .ZN(n8499) );
  INV_X1 U5807 ( .A(n6418), .ZN(n8525) );
  INV_X1 U5808 ( .A(n8608), .ZN(n8313) );
  NAND2_X1 U5809 ( .A1(n6170), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n6190) );
  NAND3_X1 U5810 ( .A1(n6164), .A2(n6166), .A3(n4401), .ZN(n8326) );
  NAND2_X1 U5811 ( .A1(n6170), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n6164) );
  OR2_X1 U5812 ( .A1(n6186), .A2(n6162), .ZN(n6166) );
  NAND2_X1 U5813 ( .A1(n4611), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4610) );
  XNOR2_X1 U5814 ( .A(n4503), .B(n7075), .ZN(n7061) );
  INV_X1 U5815 ( .A(n7095), .ZN(n4503) );
  INV_X1 U5816 ( .A(n4502), .ZN(n7096) );
  INV_X1 U5817 ( .A(n4779), .ZN(n7100) );
  XNOR2_X1 U5818 ( .A(n4777), .B(n4776), .ZN(n7278) );
  NOR2_X1 U5819 ( .A1(n7278), .A2(n6306), .ZN(n7365) );
  OAI211_X1 U5820 ( .C1(n7566), .C2(n8351), .A(n4614), .B(n4615), .ZN(n7567)
         );
  NAND2_X1 U5821 ( .A1(n4618), .A2(n4617), .ZN(n4615) );
  NAND2_X1 U5822 ( .A1(n7566), .A2(n4616), .ZN(n4614) );
  NOR2_X1 U5823 ( .A1(n4618), .A2(n4617), .ZN(n4616) );
  INV_X1 U5824 ( .A(n4775), .ZN(n9816) );
  INV_X1 U5825 ( .A(n4773), .ZN(n9814) );
  INV_X1 U5826 ( .A(n4613), .ZN(n9834) );
  INV_X1 U5827 ( .A(n4771), .ZN(n9829) );
  NAND2_X1 U5828 ( .A1(n6250), .A2(n4971), .ZN(n6365) );
  NOR2_X1 U5829 ( .A1(P2_U3150), .A2(n6817), .ZN(n9845) );
  NAND2_X1 U5830 ( .A1(n6810), .A2(n6809), .ZN(n9846) );
  AOI21_X1 U5831 ( .B1(n8400), .B2(n8399), .A(n8398), .ZN(n8410) );
  INV_X1 U5832 ( .A(n8679), .ZN(n8432) );
  NAND2_X1 U5833 ( .A1(n6453), .A2(n6442), .ZN(n8468) );
  NAND2_X1 U5834 ( .A1(n4957), .A2(n8210), .ZN(n8605) );
  OR2_X1 U5835 ( .A1(n8616), .A2(n8212), .ZN(n4957) );
  OR2_X1 U5836 ( .A1(n7207), .A2(n9901), .ZN(n8626) );
  AND2_X1 U5837 ( .A1(n6316), .A2(n6315), .ZN(n9902) );
  NAND2_X1 U5838 ( .A1(n7561), .A2(n8183), .ZN(n7665) );
  AND3_X1 U5839 ( .A1(n6278), .A2(n6277), .A3(n6276), .ZN(n9890) );
  AND3_X1 U5840 ( .A1(n6254), .A2(n6253), .A3(n6252), .ZN(n9879) );
  NAND2_X1 U5841 ( .A1(n4979), .A2(n6214), .ZN(n7493) );
  INV_X1 U5842 ( .A(n8600), .ZN(n8550) );
  AOI21_X2 U5843 ( .B1(n7456), .B2(n7455), .A(n8582), .ZN(n8630) );
  INV_X1 U5844 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n4709) );
  INV_X1 U5845 ( .A(n7942), .ZN(n4707) );
  NAND2_X1 U5846 ( .A1(n4985), .A2(n9929), .ZN(n4706) );
  INV_X1 U5847 ( .A(n8676), .ZN(n8673) );
  INV_X1 U5848 ( .A(n8433), .ZN(n8684) );
  NAND2_X1 U5849 ( .A1(n8440), .A2(n8439), .ZN(n8441) );
  NAND2_X1 U5850 ( .A1(n4692), .A2(n4695), .ZN(n8446) );
  NAND2_X1 U5851 ( .A1(n8461), .A2(n4698), .ZN(n4692) );
  OAI21_X1 U5852 ( .B1(n8461), .B2(n8263), .A(n8264), .ZN(n8450) );
  NAND2_X1 U5853 ( .A1(n8472), .A2(n4651), .ZN(n8463) );
  NAND2_X1 U5854 ( .A1(n6119), .A2(n6118), .ZN(n8704) );
  AND2_X1 U5855 ( .A1(n6428), .A2(n6427), .ZN(n8709) );
  NAND2_X1 U5856 ( .A1(n4705), .A2(n4703), .ZN(n8490) );
  NAND2_X1 U5857 ( .A1(n6420), .A2(n6419), .ZN(n8715) );
  NAND2_X1 U5858 ( .A1(n4705), .A2(n8236), .ZN(n8496) );
  NAND2_X1 U5859 ( .A1(n6146), .A2(n6145), .ZN(n8721) );
  AND2_X1 U5860 ( .A1(n4666), .A2(n4395), .ZN(n8536) );
  NAND2_X1 U5861 ( .A1(n4716), .A2(n4715), .ZN(n8532) );
  INV_X1 U5862 ( .A(n7891), .ZN(n7975) );
  NAND2_X1 U5863 ( .A1(n4716), .A2(n8233), .ZN(n7869) );
  INV_X1 U5864 ( .A(n8063), .ZN(n8741) );
  AND2_X1 U5865 ( .A1(n8581), .A2(n8580), .ZN(n8749) );
  INV_X1 U5866 ( .A(n8759), .ZN(n8753) );
  NAND2_X1 U5867 ( .A1(n6358), .A2(n6357), .ZN(n8757) );
  INV_X1 U5868 ( .A(n8740), .ZN(n8758) );
  AND3_X1 U5869 ( .A1(n6213), .A2(n6212), .A3(n6211), .ZN(n7507) );
  NAND2_X1 U5870 ( .A1(n7162), .A2(n6642), .ZN(n6651) );
  AND2_X1 U5871 ( .A1(n4977), .A2(n4976), .ZN(n4975) );
  INV_X1 U5872 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n4976) );
  BUF_X1 U5873 ( .A(n6137), .Z(n8771) );
  AND2_X1 U5874 ( .A1(n6541), .A2(n6540), .ZN(n7745) );
  NAND2_X1 U5875 ( .A1(n6156), .A2(n6112), .ZN(n6538) );
  NAND2_X1 U5876 ( .A1(n6535), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6532) );
  INV_X1 U5877 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7546) );
  INV_X1 U5878 ( .A(n8305), .ZN(n8149) );
  INV_X1 U5879 ( .A(n8151), .ZN(n8139) );
  NAND2_X1 U5880 ( .A1(n6488), .A2(n6487), .ZN(n8298) );
  INV_X1 U5881 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7223) );
  INV_X1 U5882 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n6672) );
  INV_X1 U5883 ( .A(n8395), .ZN(n9843) );
  INV_X1 U5884 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6630) );
  INV_X1 U5885 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6610) );
  INV_X1 U5886 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6606) );
  INV_X1 U5887 ( .A(n7051), .ZN(n6995) );
  INV_X1 U5888 ( .A(n6905), .ZN(n6963) );
  AND2_X1 U5889 ( .A1(n6085), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6581) );
  OR2_X1 U5890 ( .A1(n7030), .A2(n7031), .ZN(n4839) );
  AND2_X1 U5891 ( .A1(n5167), .A2(n5166), .ZN(n9148) );
  INV_X1 U5892 ( .A(n4545), .ZN(n4544) );
  AND2_X1 U5893 ( .A1(n5922), .A2(n4546), .ZN(n7760) );
  NOR2_X1 U5894 ( .A1(n8780), .A2(n8781), .ZN(n4840) );
  INV_X1 U5895 ( .A(n4844), .ZN(n4843) );
  AND3_X1 U5896 ( .A1(n5192), .A2(n5191), .A3(n5190), .ZN(n9360) );
  NOR2_X1 U5897 ( .A1(n8881), .A2(n6031), .ZN(n8844) );
  NAND2_X1 U5898 ( .A1(n6671), .A2(n5517), .ZN(n5497) );
  INV_X1 U5899 ( .A(n6857), .ZN(n6835) );
  NAND2_X1 U5900 ( .A1(n4851), .A2(n5969), .ZN(n8867) );
  NAND2_X1 U5901 ( .A1(n5956), .A2(n4852), .ZN(n4851) );
  AND3_X1 U5902 ( .A1(n5552), .A2(n5551), .A3(n5550), .ZN(n9256) );
  INV_X1 U5903 ( .A(n4550), .ZN(n4549) );
  INV_X1 U5904 ( .A(n8945), .ZN(n8899) );
  NAND2_X1 U5905 ( .A1(n6636), .A2(n5517), .ZN(n5453) );
  CLKBUF_X1 U5906 ( .A(n7029), .Z(n7030) );
  INV_X1 U5907 ( .A(n9733), .ZN(n7037) );
  AND2_X1 U5908 ( .A1(n8869), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8927) );
  INV_X1 U5909 ( .A(n9335), .ZN(n9166) );
  INV_X1 U5910 ( .A(n9256), .ZN(n9396) );
  INV_X1 U5911 ( .A(n9277), .ZN(n9405) );
  INV_X1 U5912 ( .A(n7473), .ZN(n9755) );
  OR2_X1 U5913 ( .A1(n9550), .A2(n8982), .ZN(n8983) );
  NOR2_X1 U5914 ( .A1(n9051), .A2(n9679), .ZN(n9689) );
  OR2_X1 U5915 ( .A1(n9689), .A2(n9688), .ZN(n9696) );
  INV_X1 U5916 ( .A(n9687), .ZN(n9700) );
  NAND2_X1 U5917 ( .A1(n4383), .A2(n9319), .ZN(n9307) );
  XOR2_X1 U5918 ( .A(n9084), .B(n9092), .Z(n4383) );
  OAI21_X1 U5919 ( .B1(n9178), .B2(n4800), .A(n4799), .ZN(n9146) );
  AND2_X1 U5920 ( .A1(n5179), .A2(n5178), .ZN(n9324) );
  NAND2_X1 U5921 ( .A1(n4569), .A2(n4572), .ZN(n9191) );
  OAI21_X1 U5922 ( .B1(n9223), .B2(n4571), .A(n4380), .ZN(n9189) );
  NAND2_X1 U5923 ( .A1(n9223), .A2(n4573), .ZN(n4569) );
  INV_X1 U5924 ( .A(n4916), .ZN(n4575) );
  NAND2_X1 U5925 ( .A1(n9223), .A2(n9102), .ZN(n4576) );
  INV_X1 U5926 ( .A(n9361), .ZN(n9378) );
  NAND2_X1 U5927 ( .A1(n4785), .A2(n5765), .ZN(n7831) );
  NAND2_X1 U5928 ( .A1(n7704), .A2(n4786), .ZN(n4785) );
  AND2_X1 U5929 ( .A1(n5490), .A2(n5489), .ZN(n9425) );
  OAI21_X1 U5930 ( .B1(n7691), .B2(n4902), .A(n4900), .ZN(n7820) );
  NAND2_X1 U5931 ( .A1(n7704), .A2(n5762), .ZN(n7722) );
  AND3_X1 U5932 ( .A1(n5461), .A2(n5460), .A3(n5459), .ZN(n9775) );
  NAND2_X1 U5933 ( .A1(n4905), .A2(n4907), .ZN(n7720) );
  NAND2_X1 U5934 ( .A1(n7691), .A2(n4906), .ZN(n4905) );
  NAND2_X1 U5935 ( .A1(n4928), .A2(n4927), .ZN(n7515) );
  NAND2_X1 U5936 ( .A1(n4930), .A2(n4929), .ZN(n4928) );
  NAND2_X1 U5937 ( .A1(n4932), .A2(n4935), .ZN(n7466) );
  NAND2_X1 U5938 ( .A1(n7436), .A2(n4936), .ZN(n4932) );
  NAND2_X1 U5939 ( .A1(n6790), .A2(n6789), .ZN(n6793) );
  NAND2_X1 U5940 ( .A1(n6737), .A2(n6738), .ZN(n6736) );
  INV_X1 U5941 ( .A(n9306), .ZN(n9212) );
  INV_X1 U5942 ( .A(n9284), .ZN(n9302) );
  NAND2_X1 U5943 ( .A1(n6694), .A2(n9242), .ZN(n9265) );
  INV_X1 U5944 ( .A(n9273), .ZN(n9299) );
  INV_X1 U5945 ( .A(n9314), .ZN(n4476) );
  INV_X1 U5946 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n4586) );
  INV_X1 U5947 ( .A(n7819), .ZN(n8949) );
  INV_X1 U5948 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n9471) );
  AND2_X1 U5949 ( .A1(n4943), .A2(n5122), .ZN(n4942) );
  AND2_X1 U5950 ( .A1(n5123), .A2(n5127), .ZN(n4943) );
  NOR2_X1 U5951 ( .A1(n5813), .A2(n5814), .ZN(n5815) );
  NOR2_X1 U5952 ( .A1(P1_IR_REG_24__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n5814) );
  INV_X1 U5953 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7888) );
  CLKBUF_X1 U5954 ( .A(n5830), .Z(n7446) );
  INV_X1 U5955 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7865) );
  INV_X1 U5956 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n6719) );
  INV_X1 U5957 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n6674) );
  NOR2_X1 U5958 ( .A1(n4939), .A2(n4941), .ZN(n5465) );
  INV_X1 U5959 ( .A(n5111), .ZN(n4939) );
  INV_X1 U5960 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n6612) );
  INV_X1 U5961 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6608) );
  NAND2_X1 U5962 ( .A1(n4861), .A2(n5011), .ZN(n5381) );
  NAND2_X1 U5963 ( .A1(n5351), .A2(n5009), .ZN(n4861) );
  OR2_X1 U5964 ( .A1(n5356), .A2(n5355), .ZN(n9611) );
  INV_X1 U5965 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6605) );
  INV_X1 U5966 ( .A(n5108), .ZN(n5310) );
  INV_X1 U5967 ( .A(n4727), .ZN(n7400) );
  XNOR2_X1 U5968 ( .A(n4538), .B(n8421), .ZN(n8308) );
  INV_X1 U5969 ( .A(n8425), .ZN(n4768) );
  NAND2_X1 U5970 ( .A1(n4683), .A2(n4445), .ZN(n6568) );
  AND2_X1 U5971 ( .A1(n5826), .A2(n5825), .ZN(n5827) );
  NAND2_X1 U5972 ( .A1(n9081), .A2(n7863), .ZN(n4475) );
  NAND2_X1 U5973 ( .A1(n4588), .A2(n9131), .ZN(n9323) );
  INV_X1 U5974 ( .A(n4589), .ZN(n4588) );
  OAI21_X1 U5975 ( .B1(n9432), .B2(n9811), .A(n4599), .ZN(P1_U3553) );
  AOI21_X1 U5976 ( .B1(n9084), .B2(n4601), .A(n4600), .ZN(n4599) );
  NOR2_X1 U5977 ( .A1(n9813), .A2(n9308), .ZN(n4600) );
  INV_X1 U5978 ( .A(n9423), .ZN(n4601) );
  NAND2_X1 U5979 ( .A1(n4579), .A2(n4581), .ZN(P1_U3518) );
  AND2_X1 U5980 ( .A1(n8561), .A2(n8227), .ZN(n4377) );
  INV_X1 U5981 ( .A(n4555), .ZN(n4994) );
  AND2_X1 U5982 ( .A1(n4755), .A2(n4446), .ZN(n4378) );
  AND2_X1 U5983 ( .A1(n4873), .A2(n4868), .ZN(n4379) );
  AND2_X1 U5984 ( .A1(n9190), .A2(n4570), .ZN(n4380) );
  OR2_X1 U5985 ( .A1(n8698), .A2(n8474), .ZN(n4381) );
  AND2_X1 U5986 ( .A1(n7425), .A2(n4596), .ZN(n4382) );
  INV_X1 U5987 ( .A(n4696), .ZN(n4695) );
  OAI21_X1 U5988 ( .B1(n8451), .B2(n4697), .A(n8268), .ZN(n4696) );
  NOR2_X1 U5989 ( .A1(n8612), .A2(n8124), .ZN(n4956) );
  INV_X1 U5990 ( .A(n4931), .ZN(n4929) );
  NAND2_X1 U5991 ( .A1(n4935), .A2(n4938), .ZN(n4931) );
  NAND2_X1 U5992 ( .A1(n4595), .A2(n7473), .ZN(n4938) );
  AND2_X1 U5993 ( .A1(n4657), .A2(n4656), .ZN(n4655) );
  AND2_X1 U5994 ( .A1(n8166), .A2(n8165), .ZN(n4384) );
  NAND2_X1 U5995 ( .A1(n4428), .A2(n5114), .ZN(n4385) );
  OR2_X1 U5996 ( .A1(n4499), .A2(n8416), .ZN(n4386) );
  OR2_X1 U5997 ( .A1(n9388), .A2(n9377), .ZN(n4387) );
  NAND2_X1 U5998 ( .A1(n5221), .A2(n5220), .ZN(n9185) );
  INV_X1 U5999 ( .A(n9185), .ZN(n9348) );
  INV_X1 U6000 ( .A(n7513), .ZN(n4937) );
  NAND2_X1 U6001 ( .A1(n4843), .A2(n5906), .ZN(n7547) );
  NAND2_X1 U6002 ( .A1(n6387), .A2(n4681), .ZN(n4388) );
  NAND2_X1 U6003 ( .A1(n6250), .A2(n6101), .ZN(n6264) );
  INV_X1 U6004 ( .A(n5277), .ZN(n5288) );
  INV_X1 U6005 ( .A(n4740), .ZN(n4739) );
  NAND2_X1 U6006 ( .A1(n4743), .A2(n4741), .ZN(n4740) );
  OAI21_X1 U6007 ( .B1(n8004), .B2(n4740), .A(n4737), .ZN(n7969) );
  AND2_X1 U6008 ( .A1(n4764), .A2(n4763), .ZN(n4389) );
  INV_X1 U6009 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5122) );
  OR2_X1 U6010 ( .A1(n7819), .A2(n8952), .ZN(n4390) );
  NAND2_X1 U6011 ( .A1(n4946), .A2(n6462), .ZN(n8436) );
  AND2_X1 U6012 ( .A1(n4732), .A2(n8066), .ZN(n4391) );
  AND2_X1 U6013 ( .A1(n6526), .A2(n8596), .ZN(n4392) );
  OR2_X1 U6014 ( .A1(n7112), .A2(n7095), .ZN(n4393) );
  NAND2_X1 U6015 ( .A1(n5453), .A2(n5452), .ZN(n9788) );
  INV_X1 U6016 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n6100) );
  INV_X1 U6017 ( .A(n9747), .ZN(n4595) );
  NAND2_X1 U6018 ( .A1(n5164), .A2(n5163), .ZN(n9156) );
  INV_X1 U6019 ( .A(n9156), .ZN(n9445) );
  NOR3_X1 U6020 ( .A1(n8507), .A2(n8517), .A3(n8130), .ZN(n4394) );
  NAND2_X1 U6021 ( .A1(n7975), .A2(n8537), .ZN(n4395) );
  NAND2_X1 U6022 ( .A1(n4963), .A2(n4964), .ZN(n6248) );
  OR2_X1 U6023 ( .A1(n7819), .A2(n9425), .ZN(n5765) );
  AND3_X1 U6024 ( .A1(n5394), .A2(n5393), .A3(n5392), .ZN(n7439) );
  NAND2_X1 U6025 ( .A1(n8698), .A2(n8455), .ZN(n8264) );
  NOR2_X1 U6026 ( .A1(n8256), .A2(n8479), .ZN(n4396) );
  AND2_X1 U6027 ( .A1(n5740), .A2(n5626), .ZN(n6738) );
  NAND2_X1 U6028 ( .A1(n4964), .A2(n6100), .ZN(n6221) );
  AND2_X1 U6029 ( .A1(n9363), .A2(n9369), .ZN(n4397) );
  NAND2_X1 U6030 ( .A1(n5544), .A2(n5543), .ZN(n9392) );
  AND2_X1 U6031 ( .A1(n4536), .A2(n6194), .ZN(n4398) );
  INV_X1 U6032 ( .A(n9233), .ZN(n9372) );
  NAND2_X1 U6033 ( .A1(n5208), .A2(n5207), .ZN(n9233) );
  INV_X1 U6034 ( .A(n4607), .ZN(n9163) );
  NOR2_X1 U6035 ( .A1(n9179), .A2(n9164), .ZN(n4607) );
  AND2_X1 U6036 ( .A1(n8609), .A2(n8592), .ZN(n4399) );
  AND2_X1 U6037 ( .A1(n4773), .A2(n4772), .ZN(n4400) );
  INV_X1 U6038 ( .A(n4955), .ZN(n4954) );
  AOI21_X1 U6039 ( .B1(n4956), .B2(n8212), .A(n4399), .ZN(n4955) );
  AND2_X1 U6040 ( .A1(n6165), .A2(n6167), .ZN(n4401) );
  AND2_X1 U6041 ( .A1(n7566), .A2(n7565), .ZN(n4402) );
  NAND2_X1 U6042 ( .A1(n8560), .A2(n6386), .ZN(n4403) );
  INV_X1 U6043 ( .A(n4661), .ZN(n4660) );
  NAND2_X1 U6044 ( .A1(n4665), .A2(n8517), .ZN(n4661) );
  INV_X1 U6045 ( .A(n8445), .ZN(n8437) );
  XNOR2_X1 U6046 ( .A(n8687), .B(n8454), .ZN(n8445) );
  AND2_X1 U6047 ( .A1(n8687), .A2(n8310), .ZN(n4404) );
  AND2_X1 U6048 ( .A1(n9318), .A2(n9149), .ZN(n4405) );
  OR2_X1 U6049 ( .A1(n8301), .A2(n8300), .ZN(n4406) );
  INV_X1 U6050 ( .A(n5038), .ZN(n4894) );
  INV_X1 U6051 ( .A(n4747), .ZN(n4746) );
  INV_X1 U6052 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n5113) );
  NOR2_X1 U6053 ( .A1(n7904), .A2(n8563), .ZN(n4407) );
  INV_X1 U6054 ( .A(n6667), .ZN(n7459) );
  NAND2_X1 U6055 ( .A1(n4689), .A2(n7300), .ZN(n6667) );
  NOR2_X1 U6056 ( .A1(n8865), .A2(n8864), .ZN(n4408) );
  NOR2_X1 U6057 ( .A1(n8687), .A2(n8454), .ZN(n4409) );
  NOR2_X1 U6058 ( .A1(n7897), .A2(n8592), .ZN(n4410) );
  AND2_X1 U6059 ( .A1(n8808), .A2(n5985), .ZN(n4411) );
  INV_X1 U6060 ( .A(n4651), .ZN(n4650) );
  OR2_X1 U6061 ( .A1(n8704), .A2(n8464), .ZN(n4651) );
  OR2_X1 U6062 ( .A1(n6985), .A2(n6995), .ZN(n4412) );
  NOR2_X1 U6063 ( .A1(n4679), .A2(n4894), .ZN(n4413) );
  NAND2_X1 U6064 ( .A1(n8232), .A2(n8230), .ZN(n8557) );
  NAND2_X1 U6065 ( .A1(n6482), .A2(n6481), .ZN(n4414) );
  INV_X1 U6066 ( .A(n9084), .ZN(n9435) );
  NAND2_X1 U6067 ( .A1(n5570), .A2(n5569), .ZN(n9084) );
  NOR2_X1 U6068 ( .A1(n9427), .A2(n8953), .ZN(n4415) );
  INV_X1 U6069 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n6101) );
  AND2_X1 U6070 ( .A1(n5417), .A2(n5416), .ZN(n7814) );
  AND2_X1 U6071 ( .A1(n5035), .A2(n10071), .ZN(n4416) );
  AND2_X1 U6072 ( .A1(n5013), .A2(SI_7_), .ZN(n4417) );
  NAND2_X1 U6073 ( .A1(n8806), .A2(n5987), .ZN(n4418) );
  NOR2_X1 U6074 ( .A1(n4392), .A2(n6525), .ZN(n7942) );
  INV_X1 U6075 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n5116) );
  INV_X1 U6076 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n8764) );
  INV_X1 U6077 ( .A(n8231), .ZN(n4717) );
  AND2_X1 U6078 ( .A1(n4902), .A2(n4390), .ZN(n4419) );
  AND2_X1 U6079 ( .A1(n4812), .A2(n4811), .ZN(n4420) );
  NOR2_X1 U6080 ( .A1(n9454), .A2(n9360), .ZN(n4421) );
  AND2_X1 U6081 ( .A1(n7814), .A2(n4937), .ZN(n4422) );
  NAND2_X1 U6082 ( .A1(n8233), .A2(n8230), .ZN(n4423) );
  OAI21_X1 U6083 ( .B1(n8479), .B2(n4650), .A(n6448), .ZN(n4649) );
  NAND2_X1 U6084 ( .A1(n4596), .A2(n7439), .ZN(n4935) );
  AND2_X1 U6085 ( .A1(n8535), .A2(n4395), .ZN(n4665) );
  INV_X1 U6086 ( .A(n4574), .ZN(n4573) );
  NAND2_X1 U6087 ( .A1(n9102), .A2(n4577), .ZN(n4574) );
  OR2_X1 U6088 ( .A1(n4916), .A2(n4397), .ZN(n4424) );
  AND2_X1 U6089 ( .A1(n8248), .A2(n8246), .ZN(n8521) );
  NAND2_X1 U6090 ( .A1(n4717), .A2(n8531), .ZN(n4529) );
  NAND2_X1 U6091 ( .A1(n7465), .A2(n4933), .ZN(n4425) );
  AND2_X1 U6092 ( .A1(n4576), .A2(n4575), .ZN(n4426) );
  NOR2_X1 U6093 ( .A1(n8243), .A2(n8106), .ZN(n4715) );
  NOR2_X1 U6094 ( .A1(n5592), .A2(n5638), .ZN(n4427) );
  AND2_X1 U6095 ( .A1(n4808), .A2(n5122), .ZN(n4428) );
  OR2_X1 U6096 ( .A1(n8949), .A2(n9425), .ZN(n4429) );
  AND2_X1 U6097 ( .A1(n4717), .A2(n8232), .ZN(n4430) );
  NOR2_X1 U6098 ( .A1(n8182), .A2(n4723), .ZN(n4722) );
  AND2_X1 U6099 ( .A1(n8253), .A2(n4700), .ZN(n4431) );
  AND2_X1 U6100 ( .A1(n7656), .A2(n7652), .ZN(n4432) );
  NOR2_X1 U6101 ( .A1(n9315), .A2(n4788), .ZN(n4433) );
  AND2_X1 U6102 ( .A1(n4382), .A2(n4595), .ZN(n4434) );
  XNOR2_X1 U6103 ( .A(n6210), .B(n6100), .ZN(n6915) );
  INV_X1 U6104 ( .A(n9815), .ZN(n4774) );
  AND2_X1 U6105 ( .A1(n9268), .A2(n4604), .ZN(n4435) );
  INV_X1 U6106 ( .A(n5762), .ZN(n4787) );
  OAI21_X1 U6107 ( .B1(n5504), .B2(P1_IR_REG_16__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5518) );
  INV_X1 U6108 ( .A(n6989), .ZN(n7072) );
  INV_X1 U6109 ( .A(n7112), .ZN(n7075) );
  INV_X1 U6110 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n4978) );
  AND2_X2 U6111 ( .A1(n8305), .A2(n8151), .ZN(n8289) );
  OR2_X1 U6112 ( .A1(n6579), .A2(n8740), .ZN(n4436) );
  NAND2_X1 U6113 ( .A1(n4544), .A2(n5922), .ZN(n7759) );
  AND3_X1 U6114 ( .A1(n5255), .A2(n5254), .A3(n5253), .ZN(n9278) );
  OR2_X1 U6115 ( .A1(n6579), .A2(n8667), .ZN(n4437) );
  INV_X1 U6116 ( .A(n9255), .ZN(n9368) );
  AND3_X1 U6117 ( .A1(n5242), .A2(n5241), .A3(n5240), .ZN(n9255) );
  INV_X1 U6118 ( .A(n9334), .ZN(n9196) );
  AND3_X1 U6119 ( .A1(n5229), .A2(n5228), .A3(n5227), .ZN(n9334) );
  AND3_X1 U6120 ( .A1(n5513), .A2(n5512), .A3(n5511), .ZN(n9414) );
  OR2_X1 U6121 ( .A1(n9380), .A2(n9255), .ZN(n4438) );
  INV_X1 U6122 ( .A(n4875), .ZN(n4870) );
  NAND2_X1 U6123 ( .A1(n4443), .A2(n4876), .ZN(n4875) );
  AND2_X1 U6124 ( .A1(n4785), .A2(n4784), .ZN(n4439) );
  OR2_X1 U6125 ( .A1(n7852), .A2(n9902), .ZN(n4440) );
  OR2_X1 U6126 ( .A1(n7365), .A2(n7366), .ZN(n4501) );
  INV_X1 U6127 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n10069) );
  AND2_X1 U6128 ( .A1(n4960), .A2(n4962), .ZN(n4441) );
  AND2_X1 U6129 ( .A1(n5052), .A2(SI_18_), .ZN(n4442) );
  OR2_X1 U6130 ( .A1(n5231), .A2(SI_21_), .ZN(n4443) );
  OR2_X1 U6131 ( .A1(n9445), .A2(n9465), .ZN(n4444) );
  NAND2_X1 U6132 ( .A1(n6536), .A2(n6535), .ZN(n6558) );
  INV_X1 U6133 ( .A(n7370), .ZN(n4776) );
  INV_X2 U6134 ( .A(n9811), .ZN(n9813) );
  OR2_X1 U6135 ( .A1(n9914), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n4445) );
  OAI21_X1 U6136 ( .B1(n7691), .B2(n7690), .A(n4911), .ZN(n7709) );
  NAND2_X1 U6137 ( .A1(n4839), .A2(n7032), .ZN(n7251) );
  INV_X1 U6138 ( .A(n8354), .ZN(n9828) );
  OR2_X1 U6139 ( .A1(n7896), .A2(n8314), .ZN(n4446) );
  INV_X1 U6140 ( .A(n4598), .ZN(n7692) );
  NOR2_X1 U6141 ( .A1(n7625), .A2(n9780), .ZN(n4598) );
  AND2_X1 U6142 ( .A1(n5906), .A2(n5905), .ZN(n4447) );
  OR2_X1 U6143 ( .A1(n7113), .A2(n7114), .ZN(n4609) );
  INV_X1 U6144 ( .A(SI_20_), .ZN(n10080) );
  INV_X2 U6145 ( .A(n9796), .ZN(n9798) );
  OR2_X1 U6146 ( .A1(n9798), .A2(n4586), .ZN(n4448) );
  NAND2_X1 U6147 ( .A1(n4726), .A2(n6667), .ZN(n4727) );
  AND2_X1 U6148 ( .A1(n9720), .A2(n7383), .ZN(n9319) );
  INV_X1 U6149 ( .A(n8417), .ZN(n4633) );
  AND2_X1 U6150 ( .A1(n6705), .A2(n6704), .ZN(n9783) );
  INV_X1 U6151 ( .A(n7031), .ZN(n4833) );
  INV_X1 U6152 ( .A(n7367), .ZN(n4500) );
  AND3_X1 U6153 ( .A1(n4727), .A2(n7178), .A3(n7180), .ZN(n4449) );
  AND2_X1 U6154 ( .A1(n7279), .A2(n7116), .ZN(n4450) );
  NAND2_X1 U6155 ( .A1(n4633), .A2(n4632), .ZN(n4451) );
  INV_X1 U6156 ( .A(SI_15_), .ZN(n4892) );
  INV_X1 U6157 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n4455) );
  NAND2_X1 U6158 ( .A1(n5795), .A2(n5794), .ZN(n7383) );
  NAND2_X1 U6159 ( .A1(n5813), .A2(n4942), .ZN(n9470) );
  INV_X1 U6161 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n4458) );
  INV_X1 U6162 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n4471) );
  INV_X1 U6163 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n4641) );
  INV_X1 U6164 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n4636) );
  INV_X1 U6165 ( .A(n8351), .ZN(n4618) );
  NAND2_X1 U6166 ( .A1(n4466), .A2(n4465), .ZN(n4881) );
  NAND2_X1 U6167 ( .A1(n5731), .A2(n5831), .ZN(n4469) );
  NOR2_X1 U6168 ( .A1(n6309), .A2(n7281), .ZN(n7371) );
  NOR2_X1 U6169 ( .A1(n6228), .A2(n6887), .ZN(n6990) );
  XNOR2_X1 U6170 ( .A(n7111), .B(n7112), .ZN(n7073) );
  NOR2_X1 U6171 ( .A1(n7071), .A2(n4464), .ZN(n7111) );
  NOR2_X1 U6172 ( .A1(n8372), .A2(n8371), .ZN(n8407) );
  OAI21_X1 U6173 ( .B1(n4804), .B2(n9111), .A(n9112), .ZN(n9240) );
  NOR2_X2 U6174 ( .A1(n8565), .A2(n9854), .ZN(n9853) );
  INV_X1 U6175 ( .A(n6194), .ZN(n4611) );
  OAI211_X1 U6176 ( .C1(n4498), .C2(n4497), .A(n4493), .B(n4386), .ZN(n4769)
         );
  NOR2_X1 U6177 ( .A1(n8399), .A2(n8398), .ZN(n4492) );
  INV_X1 U6178 ( .A(n9831), .ZN(n4491) );
  NAND2_X1 U6179 ( .A1(n9444), .A2(n4444), .ZN(P1_U3517) );
  NAND2_X1 U6180 ( .A1(n9237), .A2(n4918), .ZN(n4917) );
  OAI21_X1 U6181 ( .B1(n9251), .B2(n4564), .A(n4387), .ZN(n4563) );
  NAND2_X1 U6182 ( .A1(n9267), .A2(n9101), .ZN(n4565) );
  NAND2_X1 U6183 ( .A1(n9174), .A2(n4898), .ZN(n4897) );
  NAND2_X1 U6184 ( .A1(n7832), .A2(n7833), .ZN(n4561) );
  INV_X1 U6185 ( .A(n5532), .ZN(n5057) );
  AOI21_X2 U6186 ( .B1(n8274), .B2(n8284), .A(n8273), .ZN(n8280) );
  NAND2_X1 U6187 ( .A1(n5219), .A2(n5218), .ZN(n5081) );
  NOR2_X1 U6188 ( .A1(n8279), .A2(n4532), .ZN(n8290) );
  NAND2_X1 U6189 ( .A1(n7467), .A2(n7514), .ZN(n7517) );
  OR2_X1 U6190 ( .A1(n6784), .A2(n5631), .ZN(n7265) );
  INV_X1 U6191 ( .A(n5616), .ZN(n5740) );
  OAI21_X2 U6192 ( .B1(n4783), .B2(n7704), .A(n4780), .ZN(n7828) );
  NAND2_X1 U6193 ( .A1(n6886), .A2(n6963), .ZN(n7017) );
  INV_X1 U6194 ( .A(n7047), .ZN(n4608) );
  INV_X1 U6195 ( .A(n4964), .ZN(n6209) );
  NAND2_X1 U6196 ( .A1(n4545), .A2(n5922), .ZN(n7811) );
  NAND2_X1 U6197 ( .A1(n5518), .A2(n5573), .ZN(n5534) );
  NAND2_X1 U6198 ( .A1(n4844), .A2(n5906), .ZN(n7641) );
  NAND2_X1 U6199 ( .A1(n4823), .A2(n4824), .ZN(n6015) );
  INV_X1 U6200 ( .A(n5114), .ZN(n5481) );
  AND3_X4 U6201 ( .A1(n4815), .A2(n5111), .A3(n5108), .ZN(n5114) );
  INV_X2 U6202 ( .A(n7863), .ZN(n9080) );
  NAND2_X1 U6203 ( .A1(n9079), .A2(n9700), .ZN(n4473) );
  INV_X1 U6204 ( .A(n6738), .ZN(n4802) );
  NAND2_X1 U6205 ( .A1(n4475), .A2(n4472), .ZN(n9083) );
  INV_X1 U6206 ( .A(n7265), .ZN(n4814) );
  NOR2_X1 U6207 ( .A1(n9276), .A2(n9275), .ZN(n4804) );
  NAND2_X2 U6208 ( .A1(n7705), .A2(n7719), .ZN(n7704) );
  XNOR2_X1 U6209 ( .A(n4793), .B(n9109), .ZN(n4792) );
  NAND2_X1 U6210 ( .A1(n4719), .A2(n4720), .ZN(n7733) );
  NAND3_X1 U6211 ( .A1(n4969), .A2(n6250), .A3(n4710), .ZN(n6540) );
  NAND2_X1 U6212 ( .A1(n5732), .A2(n7863), .ZN(n4465) );
  NAND2_X1 U6213 ( .A1(n6749), .A2(n5619), .ZN(n4803) );
  MUX2_X1 U6214 ( .A(n5715), .B(n5714), .S(n4365), .Z(n5719) );
  INV_X1 U6215 ( .A(n4863), .ZN(n4862) );
  NAND2_X1 U6216 ( .A1(n4988), .A2(n5269), .ZN(n4557) );
  NAND2_X1 U6217 ( .A1(n4858), .A2(n5777), .ZN(n4857) );
  OAI21_X1 U6218 ( .B1(n5683), .B2(n5774), .A(n9112), .ZN(n5684) );
  OAI21_X1 U6219 ( .B1(n4881), .B2(n7383), .A(n4879), .ZN(n4878) );
  NAND2_X1 U6220 ( .A1(n5702), .A2(n5701), .ZN(n5705) );
  NAND2_X1 U6221 ( .A1(n9635), .A2(n9636), .ZN(n9634) );
  NAND3_X1 U6222 ( .A1(n4474), .A2(n9080), .A3(n4473), .ZN(n4472) );
  XNOR2_X2 U6223 ( .A(n5299), .B(P1_IR_REG_2__SCAN_IN), .ZN(n9560) );
  NAND2_X1 U6224 ( .A1(n5309), .A2(n4997), .ZN(n5000) );
  NAND2_X1 U6225 ( .A1(n4556), .A2(n4993), .ZN(n5309) );
  NAND2_X1 U6226 ( .A1(n9138), .A2(n9119), .ZN(n4793) );
  NAND3_X1 U6227 ( .A1(n9317), .A2(n4476), .A3(n4433), .ZN(n9440) );
  NAND2_X1 U6228 ( .A1(n5800), .A2(n5829), .ZN(n5731) );
  NAND3_X1 U6229 ( .A1(n5672), .A2(n5766), .A3(n6840), .ZN(n5673) );
  NAND2_X1 U6230 ( .A1(n5767), .A2(n5651), .ZN(n5672) );
  NAND2_X1 U6231 ( .A1(n4591), .A2(n4590), .ZN(n4667) );
  NAND2_X1 U6232 ( .A1(n4878), .A2(n5827), .ZN(P1_U3242) );
  AOI21_X2 U6233 ( .B1(n4479), .B2(n9765), .A(n4477), .ZN(n9322) );
  NOR2_X1 U6234 ( .A1(n5643), .A2(n5401), .ZN(n5595) );
  NAND2_X1 U6235 ( .A1(n9240), .A2(n9239), .ZN(n9238) );
  NAND2_X1 U6236 ( .A1(n4557), .A2(n4990), .ZN(n5295) );
  INV_X1 U6237 ( .A(n5750), .ZN(n4813) );
  NAND2_X1 U6238 ( .A1(n4583), .A2(n4587), .ZN(n9441) );
  NAND2_X1 U6239 ( .A1(n4376), .A2(n4986), .ZN(n5285) );
  NAND2_X4 U6240 ( .A1(n4639), .A2(n4638), .ZN(n4555) );
  OR2_X2 U6241 ( .A1(n9819), .A2(n4482), .ZN(n4481) );
  NAND2_X1 U6242 ( .A1(n4609), .A2(n4450), .ZN(n7280) );
  NAND2_X1 U6243 ( .A1(n4620), .A2(n7132), .ZN(n6883) );
  NOR2_X1 U6244 ( .A1(n8365), .A2(n8366), .ZN(n9836) );
  NAND2_X1 U6245 ( .A1(n7084), .A2(n6894), .ZN(n8334) );
  INV_X1 U6246 ( .A(n8334), .ZN(n4487) );
  NAND2_X1 U6247 ( .A1(n4485), .A2(n6896), .ZN(n4484) );
  INV_X1 U6248 ( .A(n4766), .ZN(n4485) );
  NAND2_X1 U6249 ( .A1(n4487), .A2(n6896), .ZN(n4486) );
  NAND3_X1 U6250 ( .A1(n8333), .A2(n6896), .A3(n4488), .ZN(n4489) );
  NOR2_X1 U6251 ( .A1(n4492), .A2(n8409), .ZN(n4499) );
  NAND2_X1 U6252 ( .A1(n4412), .A2(n4504), .ZN(n7048) );
  NAND2_X1 U6253 ( .A1(n6985), .A2(n6995), .ZN(n4504) );
  NAND2_X1 U6254 ( .A1(n4775), .A2(n4774), .ZN(n4773) );
  NAND2_X1 U6255 ( .A1(n4775), .A2(n4507), .ZN(n4506) );
  INV_X1 U6256 ( .A(n4516), .ZN(n4523) );
  NAND2_X1 U6257 ( .A1(n4521), .A2(n4517), .ZN(n8244) );
  AOI22_X1 U6258 ( .A1(n4524), .A2(n4520), .B1(n4523), .B2(n4518), .ZN(n4517)
         );
  OR2_X1 U6259 ( .A1(n8229), .A2(n4522), .ZN(n4521) );
  INV_X1 U6260 ( .A(n4525), .ZN(n4524) );
  OAI21_X1 U6261 ( .B1(n4527), .B2(n8106), .A(n8284), .ZN(n4525) );
  AND2_X1 U6262 ( .A1(n4430), .A2(n4528), .ZN(n4527) );
  NAND2_X1 U6263 ( .A1(n4377), .A2(n8228), .ZN(n4528) );
  INV_X1 U6264 ( .A(n8211), .ZN(n8214) );
  OAI211_X1 U6265 ( .C1(n8205), .C2(n8289), .A(n8206), .B(n4531), .ZN(n4530)
         );
  OR2_X1 U6266 ( .A1(n8204), .A2(n8284), .ZN(n4531) );
  AOI21_X1 U6267 ( .B1(n4535), .B2(n4396), .A(n8267), .ZN(n4534) );
  OR2_X2 U6268 ( .A1(n5920), .A2(n5919), .ZN(n4546) );
  OAI21_X1 U6269 ( .B1(n8791), .B2(n4549), .A(n4547), .ZN(n5992) );
  OR2_X2 U6270 ( .A1(n8924), .A2(n4842), .ZN(n4841) );
  OAI21_X2 U6271 ( .B1(n8903), .B2(n8907), .A(n8797), .ZN(n8879) );
  NOR2_X2 U6272 ( .A1(n8905), .A2(n8904), .ZN(n8903) );
  NAND2_X1 U6273 ( .A1(n4555), .A2(SI_0_), .ZN(n5284) );
  NAND2_X1 U6274 ( .A1(n4555), .A2(P1_U3086), .ZN(n9484) );
  MUX2_X1 U6275 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(P1_DATAO_REG_20__SCAN_IN), 
        .S(n4810), .Z(n5243) );
  MUX2_X1 U6276 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(P1_DATAO_REG_21__SCAN_IN), 
        .S(n4810), .Z(n5231) );
  MUX2_X1 U6277 ( .A(n7888), .B(n7546), .S(n4810), .Z(n5062) );
  MUX2_X1 U6278 ( .A(n7865), .B(n7223), .S(n4810), .Z(n5053) );
  MUX2_X1 U6279 ( .A(n7640), .B(n5066), .S(n4810), .Z(n5067) );
  MUX2_X1 U6280 ( .A(n7739), .B(n7742), .S(n4810), .Z(n5077) );
  MUX2_X1 U6281 ( .A(n7784), .B(n5082), .S(n4810), .Z(n5083) );
  MUX2_X1 U6282 ( .A(n9486), .B(n5088), .S(n4810), .Z(n5089) );
  MUX2_X1 U6283 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(P1_DATAO_REG_28__SCAN_IN), 
        .S(n4810), .Z(n5094) );
  MUX2_X1 U6284 ( .A(n7868), .B(n5098), .S(n4810), .Z(n5099) );
  MUX2_X1 U6285 ( .A(n9482), .B(n5102), .S(n4810), .Z(n5103) );
  MUX2_X1 U6286 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n4810), .Z(n5566) );
  NAND2_X1 U6287 ( .A1(n5295), .A2(n4991), .ZN(n4556) );
  NAND3_X1 U6288 ( .A1(n4562), .A2(n4899), .A3(n4429), .ZN(n7832) );
  NAND2_X1 U6289 ( .A1(n9223), .A2(n4380), .ZN(n4567) );
  NAND2_X1 U6290 ( .A1(n4567), .A2(n4568), .ZN(n9174) );
  NAND2_X1 U6291 ( .A1(n9131), .A2(n4580), .ZN(n4583) );
  NAND3_X1 U6292 ( .A1(n4580), .A2(n9131), .A3(n9798), .ZN(n4579) );
  AOI21_X1 U6293 ( .B1(n4922), .B2(n9107), .A(n9132), .ZN(n4589) );
  NOR2_X2 U6294 ( .A1(n4597), .A2(n7513), .ZN(n7523) );
  NAND2_X1 U6295 ( .A1(n4434), .A2(n7269), .ZN(n4597) );
  INV_X1 U6296 ( .A(n4597), .ZN(n7470) );
  NAND2_X1 U6297 ( .A1(n9268), .A2(n4602), .ZN(n9226) );
  NOR2_X2 U6298 ( .A1(n9218), .A2(n9201), .ZN(n9200) );
  NAND2_X2 U6299 ( .A1(n5822), .A2(n9485), .ZN(n6622) );
  MUX2_X1 U6300 ( .A(n7214), .B(P2_REG2_REG_2__SCAN_IN), .S(n8338), .Z(n8332)
         );
  NOR2_X1 U6301 ( .A1(n7567), .A2(n7569), .ZN(n8342) );
  NAND2_X1 U6302 ( .A1(n8330), .A2(n6882), .ZN(n4622) );
  NAND2_X1 U6303 ( .A1(n4623), .A2(n8330), .ZN(n4621) );
  NAND2_X2 U6304 ( .A1(n4622), .A2(n6915), .ZN(n7132) );
  OAI21_X1 U6305 ( .B1(n4625), .B2(n9853), .A(n4624), .ZN(n4626) );
  NAND2_X1 U6306 ( .A1(n9853), .A2(n4451), .ZN(n4624) );
  AND2_X1 U6307 ( .A1(n4631), .A2(n8417), .ZN(n4625) );
  NAND2_X1 U6308 ( .A1(n4626), .A2(n4627), .ZN(n8427) );
  NOR2_X1 U6309 ( .A1(n9853), .A2(n8369), .ZN(n8372) );
  NAND2_X1 U6310 ( .A1(n8473), .A2(n4647), .ZN(n4643) );
  NAND2_X1 U6311 ( .A1(n4643), .A2(n4645), .ZN(n4944) );
  NAND2_X1 U6312 ( .A1(n5419), .A2(n4672), .ZN(n4671) );
  NAND3_X1 U6313 ( .A1(n7942), .A2(n9914), .A3(n4985), .ZN(n4683) );
  AND2_X1 U6314 ( .A1(n4964), .A2(n4684), .ZN(n6236) );
  INV_X1 U6315 ( .A(n8174), .ZN(n4686) );
  NAND2_X1 U6316 ( .A1(n6489), .A2(n8148), .ZN(n8108) );
  NAND4_X1 U6317 ( .A1(n6489), .A2(n8148), .A3(n7300), .A4(n4689), .ZN(n6490)
         );
  NAND2_X1 U6318 ( .A1(n8461), .A2(n4693), .ZN(n4690) );
  NAND2_X1 U6319 ( .A1(n4690), .A2(n4691), .ZN(n8091) );
  INV_X1 U6320 ( .A(n8263), .ZN(n4699) );
  OAI21_X1 U6321 ( .B1(n8506), .B2(n4702), .A(n4431), .ZN(n6508) );
  NAND2_X1 U6322 ( .A1(n9927), .A2(n4709), .ZN(n4708) );
  INV_X1 U6323 ( .A(n8548), .ZN(n4718) );
  NAND2_X1 U6324 ( .A1(n4712), .A2(n4713), .ZN(n6505) );
  NAND2_X1 U6325 ( .A1(n8548), .A2(n4715), .ZN(n4712) );
  NAND2_X1 U6326 ( .A1(n7559), .A2(n4722), .ZN(n4719) );
  NAND4_X1 U6327 ( .A1(n6105), .A2(n6104), .A3(n6103), .A4(n6102), .ZN(n6106)
         );
  NAND2_X1 U6328 ( .A1(n7934), .A2(n7179), .ZN(n4726) );
  NAND2_X1 U6329 ( .A1(n4727), .A2(n7178), .ZN(n4725) );
  NAND2_X1 U6330 ( .A1(n7986), .A2(n4391), .ZN(n4730) );
  NAND2_X1 U6331 ( .A1(n8004), .A2(n4737), .ZN(n4734) );
  NAND2_X1 U6332 ( .A1(n4734), .A2(n4735), .ZN(n7905) );
  NAND2_X1 U6333 ( .A1(n7903), .A2(n8578), .ZN(n4747) );
  OAI21_X2 U6334 ( .B1(n7895), .B2(n4751), .A(n4749), .ZN(n8085) );
  NAND2_X1 U6335 ( .A1(n7653), .A2(n4432), .ZN(n7771) );
  NAND2_X1 U6336 ( .A1(n7231), .A2(n4758), .ZN(n7329) );
  INV_X1 U6337 ( .A(n7328), .ZN(n4757) );
  NAND2_X1 U6338 ( .A1(n8049), .A2(n4760), .ZN(n7926) );
  NAND2_X1 U6339 ( .A1(n6482), .A2(n4761), .ZN(n4765) );
  OAI21_X1 U6340 ( .B1(n8334), .B2(n4766), .A(n8333), .ZN(n8335) );
  NAND2_X1 U6341 ( .A1(n8338), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n4767) );
  OAI211_X1 U6342 ( .C1(n8427), .C2(n9856), .A(n4769), .B(n4768), .ZN(P2_U3201) );
  INV_X1 U6343 ( .A(n4794), .ZN(n9139) );
  OAI21_X1 U6344 ( .B1(n4802), .B2(n4803), .A(n4801), .ZN(n6703) );
  AOI21_X1 U6345 ( .B1(n6738), .B2(n5618), .A(n5616), .ZN(n4801) );
  NAND2_X1 U6346 ( .A1(n5114), .A2(n4805), .ZN(n5126) );
  NAND3_X1 U6347 ( .A1(n9485), .A2(n9542), .A3(n8987), .ZN(n4811) );
  NAND2_X2 U6348 ( .A1(n6622), .A2(n4555), .ZN(n5296) );
  NAND2_X1 U6349 ( .A1(n6622), .A2(n4809), .ZN(n4812) );
  AND2_X2 U6350 ( .A1(n5298), .A2(n5106), .ZN(n5108) );
  AND4_X2 U6351 ( .A1(n4820), .A2(n4819), .A3(n4818), .A4(n4817), .ZN(n5111)
         );
  NOR2_X2 U6352 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n4817) );
  NOR2_X2 U6353 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n4818) );
  NOR2_X2 U6354 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n4819) );
  NAND2_X1 U6355 ( .A1(n8889), .A2(n4827), .ZN(n4823) );
  NAND2_X1 U6356 ( .A1(n4829), .A2(n4835), .ZN(n5903) );
  NAND2_X1 U6357 ( .A1(n7029), .A2(n4837), .ZN(n4829) );
  AND2_X2 U6358 ( .A1(n4841), .A2(n4840), .ZN(n8783) );
  NOR2_X2 U6359 ( .A1(n8844), .A2(n8843), .ZN(n8924) );
  NAND2_X1 U6360 ( .A1(n5905), .A2(n7548), .ZN(n4844) );
  NAND2_X1 U6361 ( .A1(n7641), .A2(n7643), .ZN(n7642) );
  OAI21_X1 U6362 ( .B1(n5956), .B2(n4848), .A(n4846), .ZN(n8807) );
  AOI21_X1 U6363 ( .B1(n4846), .B2(n4848), .A(n4411), .ZN(n4845) );
  INV_X1 U6364 ( .A(n4855), .ZN(n5792) );
  NAND2_X1 U6365 ( .A1(n4855), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5793) );
  OAI21_X1 U6366 ( .B1(n5705), .B2(n9116), .A(n5704), .ZN(n4858) );
  NAND2_X1 U6367 ( .A1(n5245), .A2(n4379), .ZN(n4865) );
  NAND2_X1 U6368 ( .A1(n5245), .A2(n4877), .ZN(n4872) );
  OAI21_X1 U6369 ( .B1(n5494), .B2(n4884), .A(n4882), .ZN(n5532) );
  NAND2_X1 U6370 ( .A1(n4893), .A2(n4891), .ZN(n5041) );
  NAND2_X1 U6371 ( .A1(n5464), .A2(n5039), .ZN(n4893) );
  NAND2_X1 U6372 ( .A1(n6931), .A2(n6930), .ZN(n6929) );
  NAND2_X2 U6373 ( .A1(n4420), .A2(n5271), .ZN(n8823) );
  NAND3_X1 U6374 ( .A1(n7691), .A2(n4390), .A3(n4900), .ZN(n4899) );
  NAND2_X1 U6375 ( .A1(n6772), .A2(n4913), .ZN(n4912) );
  NAND2_X2 U6376 ( .A1(n4917), .A2(n4438), .ZN(n9223) );
  NAND2_X1 U6377 ( .A1(n4919), .A2(n4920), .ZN(n9110) );
  NAND2_X1 U6378 ( .A1(n9147), .A2(n4921), .ZN(n4919) );
  NAND2_X1 U6379 ( .A1(n7436), .A2(n4925), .ZN(n4923) );
  INV_X1 U6380 ( .A(n4941), .ZN(n5352) );
  NAND2_X1 U6381 ( .A1(n4944), .A2(n4945), .ZN(n6480) );
  NAND2_X1 U6382 ( .A1(n8452), .A2(n6461), .ZN(n4946) );
  INV_X1 U6383 ( .A(n7731), .ZN(n4961) );
  NAND2_X1 U6384 ( .A1(n6115), .A2(n6113), .ZN(n6133) );
  NAND2_X1 U6385 ( .A1(n6115), .A2(n4975), .ZN(n8765) );
  AND2_X2 U6386 ( .A1(n9290), .A2(n9400), .ZN(n9268) );
  NOR2_X2 U6387 ( .A1(n7834), .A2(n9096), .ZN(n9290) );
  AOI21_X1 U6388 ( .B1(n8442), .B2(n8596), .A(n8441), .ZN(n8685) );
  XNOR2_X1 U6389 ( .A(n8436), .B(n8437), .ZN(n8442) );
  NAND2_X1 U6390 ( .A1(n5887), .A2(n5886), .ZN(n6829) );
  NOR2_X2 U6391 ( .A1(n6941), .A2(n6757), .ZN(n6760) );
  NAND2_X1 U6392 ( .A1(n7173), .A2(n7172), .ZN(n7200) );
  NAND2_X1 U6393 ( .A1(n7173), .A2(n4984), .ZN(n7175) );
  INV_X1 U6394 ( .A(n5884), .ZN(n5887) );
  CLKBUF_X1 U6395 ( .A(n5822), .Z(n9542) );
  NAND2_X1 U6396 ( .A1(n7915), .A2(n7914), .ZN(n8048) );
  NAND2_X1 U6397 ( .A1(n7793), .A2(n7792), .ZN(n7854) );
  NAND2_X1 U6398 ( .A1(n7773), .A2(n7772), .ZN(n7793) );
  NOR2_X1 U6399 ( .A1(n7791), .A2(n7790), .ZN(n7792) );
  INV_X1 U6400 ( .A(n7794), .ZN(n7791) );
  XNOR2_X1 U6401 ( .A(n5840), .B(n4371), .ZN(n5850) );
  NOR2_X2 U6402 ( .A1(n6794), .A2(n7037), .ZN(n7269) );
  XNOR2_X1 U6403 ( .A(n6561), .B(n6560), .ZN(n7160) );
  NAND2_X1 U6404 ( .A1(n6561), .A2(n6560), .ZN(n6530) );
  AND2_X4 U6405 ( .A1(n6521), .A2(n4555), .ZN(n6192) );
  OAI211_X1 U6406 ( .C1(n7348), .C2(n8651), .A(n6425), .B(n6424), .ZN(n8511)
         );
  INV_X1 U6407 ( .A(n7348), .ZN(n6514) );
  OAI21_X2 U6408 ( .B1(n8518), .B2(n6506), .A(n8248), .ZN(n8506) );
  INV_X2 U6409 ( .A(n8823), .ZN(n6959) );
  NAND2_X1 U6410 ( .A1(n8028), .A2(n8029), .ZN(n7910) );
  NAND2_X1 U6411 ( .A1(n6133), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6114) );
  OR2_X1 U6412 ( .A1(n8323), .A2(n7232), .ZN(n4980) );
  OR2_X1 U6413 ( .A1(n9274), .A2(n9256), .ZN(n4981) );
  INV_X1 U6414 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n6122) );
  NAND2_X1 U6415 ( .A1(n5712), .A2(n9119), .ZN(n9132) );
  INV_X1 U6416 ( .A(n7851), .ZN(n7790) );
  AND2_X1 U6417 ( .A1(n5022), .A2(n5021), .ZN(n4982) );
  NOR3_X1 U6418 ( .A1(n9145), .A2(n9161), .A3(n5607), .ZN(n4983) );
  NAND2_X1 U6419 ( .A1(n5780), .A2(n9118), .ZN(n9145) );
  AND2_X1 U6420 ( .A1(n7172), .A2(n7171), .ZN(n4984) );
  NAND2_X1 U6421 ( .A1(n7910), .A2(n7909), .ZN(n7978) );
  INV_X1 U6422 ( .A(n8179), .ZN(n6268) );
  INV_X1 U6423 ( .A(n5780), .ZN(n5710) );
  INV_X1 U6424 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n5115) );
  INV_X1 U6425 ( .A(n9132), .ZN(n5608) );
  INV_X1 U6426 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5106) );
  INV_X1 U6427 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n6113) );
  INV_X1 U6428 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n6099) );
  NOR2_X1 U6429 ( .A1(n5473), .A2(n5472), .ZN(n5471) );
  AND2_X1 U6430 ( .A1(n5367), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n5412) );
  INV_X1 U6431 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n5018) );
  NAND2_X1 U6432 ( .A1(n7908), .A2(n8311), .ZN(n7909) );
  OAI22_X1 U6433 ( .A1(n7324), .A2(n6240), .B1(n7336), .B2(n8322), .ZN(n7482)
         );
  AND2_X1 U6434 ( .A1(n5471), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n5485) );
  NOR2_X1 U6435 ( .A1(n5548), .A2(n5146), .ZN(n5237) );
  OR2_X1 U6436 ( .A1(n5457), .A2(n5456), .ZN(n5473) );
  OR2_X1 U6437 ( .A1(n5389), .A2(n5388), .ZN(n5391) );
  INV_X1 U6438 ( .A(n9611), .ZN(n9019) );
  INV_X1 U6439 ( .A(SI_23_), .ZN(n10097) );
  INV_X1 U6440 ( .A(SI_19_), .ZN(n10120) );
  INV_X1 U6441 ( .A(SI_9_), .ZN(n10144) );
  INV_X1 U6442 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n4996) );
  INV_X1 U6443 ( .A(n8316), .ZN(n7852) );
  AND2_X1 U6444 ( .A1(n7898), .A2(n8313), .ZN(n7899) );
  OR2_X1 U6445 ( .A1(n7174), .A2(n8284), .ZN(n7294) );
  AND2_X1 U6446 ( .A1(n6292), .A2(n6291), .ZN(n6295) );
  AND2_X1 U6447 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n5315) );
  AND2_X1 U6448 ( .A1(n5188), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n5174) );
  INV_X1 U6449 ( .A(n4372), .ZN(n5199) );
  AND2_X1 U6450 ( .A1(n5158), .A2(n5157), .ZN(n9135) );
  INV_X1 U6451 ( .A(n9242), .ZN(n9291) );
  INV_X1 U6452 ( .A(n6699), .ZN(n6084) );
  INV_X1 U6453 ( .A(n7383), .ZN(n6839) );
  OR2_X1 U6454 ( .A1(n5100), .A2(n5099), .ZN(n5101) );
  INV_X1 U6455 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n5123) );
  INV_X1 U6456 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5809) );
  INV_X1 U6457 ( .A(SI_18_), .ZN(n10056) );
  INV_X1 U6458 ( .A(SI_12_), .ZN(n5031) );
  XNOR2_X1 U6459 ( .A(n7787), .B(n7788), .ZN(n7773) );
  INV_X1 U6460 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n6124) );
  AND2_X1 U6461 ( .A1(n7892), .A2(n8315), .ZN(n7893) );
  INV_X1 U6462 ( .A(n8078), .ZN(n8031) );
  OR2_X1 U6463 ( .A1(n7167), .A2(n7166), .ZN(n8081) );
  INV_X1 U6464 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n6560) );
  INV_X1 U6465 ( .A(n6186), .ZN(n6423) );
  OR2_X1 U6466 ( .A1(n6811), .A2(n8776), .ZN(n6889) );
  INV_X1 U6467 ( .A(n8206), .ZN(n7752) );
  NOR2_X1 U6468 ( .A1(n9870), .A2(n8151), .ZN(n7161) );
  INV_X1 U6469 ( .A(n7666), .ZN(n7456) );
  OR2_X1 U6470 ( .A1(n7202), .A2(n7200), .ZN(n6573) );
  INV_X1 U6471 ( .A(n8474), .ZN(n8455) );
  NAND2_X1 U6472 ( .A1(n8259), .A2(n8260), .ZN(n8479) );
  AND2_X1 U6473 ( .A1(n8217), .A2(n6499), .ZN(n8612) );
  OR2_X1 U6474 ( .A1(n8124), .A2(n8212), .ZN(n8629) );
  INV_X1 U6475 ( .A(n8596), .ZN(n8618) );
  INV_X1 U6476 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n6483) );
  AND2_X1 U6477 ( .A1(n6295), .A2(n6294), .ZN(n6318) );
  AND2_X1 U6478 ( .A1(n6044), .A2(n6043), .ZN(n8781) );
  NAND2_X1 U6479 ( .A1(n5236), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n5210) );
  OR2_X1 U6480 ( .A1(n6083), .A2(n6686), .ZN(n6082) );
  INV_X1 U6481 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n7645) );
  OR2_X1 U6482 ( .A1(n9547), .A2(n9564), .ZN(n9692) );
  NOR2_X1 U6483 ( .A1(n9300), .A2(n9405), .ZN(n9099) );
  NAND2_X1 U6484 ( .A1(n9720), .A2(n6698), .ZN(n9768) );
  OR2_X1 U6485 ( .A1(n6700), .A2(n6821), .ZN(n7259) );
  OR2_X1 U6486 ( .A1(n6840), .A2(n6839), .ZN(n9738) );
  NOR2_X1 U6487 ( .A1(n5809), .A2(n5124), .ZN(n5810) );
  INV_X1 U6488 ( .A(n8511), .ZN(n8485) );
  INV_X1 U6489 ( .A(n7978), .ZN(n7979) );
  OR2_X1 U6490 ( .A1(n7219), .A2(n7633), .ZN(n8077) );
  OR3_X1 U6491 ( .A1(n6542), .A2(n6558), .A3(n6559), .ZN(n6587) );
  INV_X1 U6492 ( .A(n9858), .ZN(n8361) );
  NOR2_X1 U6493 ( .A1(n6889), .A2(n6888), .ZN(n8426) );
  NAND2_X1 U6494 ( .A1(n7162), .A2(n7161), .ZN(n8624) );
  NAND2_X1 U6495 ( .A1(n6562), .A2(n8300), .ZN(n8596) );
  INV_X1 U6496 ( .A(n8624), .ZN(n8599) );
  NOR2_X1 U6497 ( .A1(n9927), .A2(n9908), .ZN(n8676) );
  INV_X1 U6498 ( .A(n8667), .ZN(n8675) );
  AND2_X1 U6499 ( .A1(n8234), .A2(n8531), .ZN(n8128) );
  NOR2_X1 U6500 ( .A1(n9915), .A2(n9908), .ZN(n8759) );
  INV_X1 U6501 ( .A(n9901), .ZN(n9913) );
  INV_X1 U6502 ( .A(n9870), .ZN(n9898) );
  INV_X1 U6503 ( .A(n9908), .ZN(n9906) );
  NAND2_X1 U6504 ( .A1(n7160), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7218) );
  NOR2_X1 U6505 ( .A1(n6296), .A2(n6318), .ZN(n7118) );
  AND2_X1 U6506 ( .A1(n5169), .A2(n5168), .ZN(n9335) );
  INV_X1 U6507 ( .A(n9704), .ZN(n9664) );
  INV_X1 U6508 ( .A(n9319), .ZN(n9792) );
  AND2_X1 U6509 ( .A1(n5585), .A2(n5703), .ZN(n9175) );
  AND2_X1 U6510 ( .A1(n5680), .A2(n5678), .ZN(n9287) );
  AND2_X1 U6511 ( .A1(n5749), .A2(n7516), .ZN(n7514) );
  AND2_X1 U6512 ( .A1(n9265), .A2(n7863), .ZN(n9284) );
  INV_X1 U6513 ( .A(n6854), .ZN(n6850) );
  INV_X1 U6514 ( .A(n9794), .ZN(n9760) );
  INV_X1 U6515 ( .A(n9783), .ZN(n9765) );
  NAND2_X1 U6516 ( .A1(n7259), .A2(n9738), .ZN(n9794) );
  INV_X1 U6517 ( .A(n8077), .ZN(n8061) );
  INV_X1 U6518 ( .A(n8454), .ZN(n8310) );
  INV_X1 U6519 ( .A(n8621), .ZN(n8592) );
  INV_X1 U6520 ( .A(n9845), .ZN(n8387) );
  INV_X1 U6521 ( .A(n8426), .ZN(n9860) );
  INV_X1 U6522 ( .A(n9846), .ZN(n9844) );
  INV_X1 U6523 ( .A(n8630), .ZN(n8603) );
  NAND2_X1 U6524 ( .A1(n9929), .A2(n9913), .ZN(n8667) );
  INV_X1 U6525 ( .A(n9929), .ZN(n9927) );
  AND2_X2 U6526 ( .A1(n7206), .A2(n6578), .ZN(n9929) );
  NAND2_X1 U6527 ( .A1(n9914), .A2(n9913), .ZN(n8740) );
  AND3_X1 U6528 ( .A1(n9893), .A2(n9892), .A3(n9891), .ZN(n9923) );
  AND2_X1 U6529 ( .A1(n6567), .A2(n6566), .ZN(n9915) );
  INV_X2 U6530 ( .A(n9915), .ZN(n9914) );
  INV_X1 U6531 ( .A(n7218), .ZN(n6647) );
  INV_X1 U6532 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n6720) );
  INV_X1 U6533 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6617) );
  INV_X1 U6534 ( .A(n8936), .ZN(n8920) );
  INV_X1 U6535 ( .A(n9199), .ZN(n9369) );
  OR2_X1 U6536 ( .A1(n9547), .A2(n9561), .ZN(n9704) );
  NAND2_X1 U6537 ( .A1(n9265), .A2(n6701), .ZN(n9306) );
  NAND2_X1 U6538 ( .A1(n9813), .A2(n9787), .ZN(n9423) );
  NAND2_X1 U6539 ( .A1(n6855), .A2(n6850), .ZN(n9811) );
  NAND2_X1 U6540 ( .A1(n9798), .A2(n9787), .ZN(n9465) );
  NAND2_X1 U6541 ( .A1(n6855), .A2(n6854), .ZN(n9796) );
  NAND2_X2 U6542 ( .A1(n6687), .A2(n6689), .ZN(n9717) );
  INV_X1 U6543 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7701) );
  INV_X1 U6544 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6629) );
  INV_X2 U6545 ( .A(n8383), .ZN(P2_U3893) );
  AND2_X2 U6546 ( .A1(n6582), .A2(n6581), .ZN(P1_U3973) );
  XNOR2_X1 U6547 ( .A(n4989), .B(SI_1_), .ZN(n5270) );
  INV_X1 U6548 ( .A(n5270), .ZN(n4988) );
  AND2_X1 U6549 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n4986) );
  NAND3_X1 U6550 ( .A1(n4994), .A2(SI_0_), .A3(P1_DATAO_REG_0__SCAN_IN), .ZN(
        n4987) );
  NAND2_X1 U6551 ( .A1(n5285), .A2(n4987), .ZN(n5269) );
  NAND2_X1 U6552 ( .A1(n4989), .A2(SI_1_), .ZN(n4990) );
  MUX2_X1 U6553 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .S(n4376), .Z(n4992) );
  INV_X1 U6554 ( .A(n5294), .ZN(n4991) );
  NAND2_X1 U6555 ( .A1(n4992), .A2(SI_2_), .ZN(n4993) );
  XNOR2_X1 U6556 ( .A(n4998), .B(SI_3_), .ZN(n5308) );
  INV_X1 U6557 ( .A(n5308), .ZN(n4997) );
  NAND2_X1 U6558 ( .A1(n4998), .A2(SI_3_), .ZN(n4999) );
  NAND2_X1 U6559 ( .A1(n5000), .A2(n4999), .ZN(n5324) );
  INV_X1 U6560 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6598) );
  MUX2_X1 U6561 ( .A(n6598), .B(n6605), .S(n4555), .Z(n5001) );
  XNOR2_X1 U6562 ( .A(n5001), .B(SI_4_), .ZN(n5323) );
  NAND2_X1 U6563 ( .A1(n5324), .A2(n5323), .ZN(n5004) );
  INV_X1 U6564 ( .A(n5001), .ZN(n5002) );
  NAND2_X1 U6565 ( .A1(n5002), .A2(SI_4_), .ZN(n5003) );
  NAND2_X1 U6566 ( .A1(n5004), .A2(n5003), .ZN(n5335) );
  MUX2_X1 U6567 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n4555), .Z(n5006) );
  INV_X1 U6568 ( .A(SI_5_), .ZN(n5005) );
  XNOR2_X1 U6569 ( .A(n5006), .B(n5005), .ZN(n5334) );
  NAND2_X1 U6570 ( .A1(n5335), .A2(n5334), .ZN(n5008) );
  NAND2_X1 U6571 ( .A1(n5006), .A2(SI_5_), .ZN(n5007) );
  XNOR2_X1 U6572 ( .A(n5010), .B(SI_6_), .ZN(n5350) );
  INV_X1 U6573 ( .A(n5350), .ZN(n5009) );
  NAND2_X1 U6574 ( .A1(n5010), .A2(SI_6_), .ZN(n5011) );
  MUX2_X1 U6575 ( .A(n6606), .B(n6608), .S(n4555), .Z(n5012) );
  XNOR2_X1 U6576 ( .A(n5012), .B(SI_7_), .ZN(n5380) );
  INV_X1 U6577 ( .A(n5012), .ZN(n5013) );
  MUX2_X1 U6578 ( .A(n6610), .B(n6612), .S(n4555), .Z(n5014) );
  NAND2_X1 U6579 ( .A1(n5014), .A2(n10078), .ZN(n5017) );
  INV_X1 U6580 ( .A(n5014), .ZN(n5015) );
  NAND2_X1 U6581 ( .A1(n5015), .A2(SI_8_), .ZN(n5016) );
  NAND2_X1 U6582 ( .A1(n5017), .A2(n5016), .ZN(n5395) );
  MUX2_X1 U6583 ( .A(n6617), .B(n5018), .S(n4555), .Z(n5019) );
  NAND2_X1 U6584 ( .A1(n5019), .A2(n10144), .ZN(n5022) );
  INV_X1 U6585 ( .A(n5019), .ZN(n5020) );
  NAND2_X1 U6586 ( .A1(n5020), .A2(SI_9_), .ZN(n5021) );
  NAND2_X1 U6587 ( .A1(n5360), .A2(n4982), .ZN(n5023) );
  MUX2_X1 U6588 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .S(n4555), .Z(n5025) );
  NAND2_X1 U6589 ( .A1(n5025), .A2(SI_10_), .ZN(n5026) );
  MUX2_X1 U6590 ( .A(n6630), .B(n6629), .S(n4555), .Z(n5027) );
  INV_X1 U6591 ( .A(n5027), .ZN(n5028) );
  NAND2_X1 U6592 ( .A1(n5028), .A2(SI_11_), .ZN(n5029) );
  NAND2_X1 U6593 ( .A1(n5030), .A2(n5029), .ZN(n5418) );
  MUX2_X1 U6594 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .S(n4555), .Z(n5032) );
  NAND2_X1 U6595 ( .A1(n5032), .A2(SI_12_), .ZN(n5033) );
  MUX2_X1 U6596 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n4555), .Z(n5446) );
  NOR2_X1 U6597 ( .A1(n5035), .A2(n10071), .ZN(n5036) );
  MUX2_X1 U6598 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n4555), .Z(n5462) );
  INV_X1 U6599 ( .A(n5462), .ZN(n5037) );
  NAND2_X1 U6600 ( .A1(n5037), .A2(n10058), .ZN(n5038) );
  NAND2_X1 U6601 ( .A1(n5462), .A2(SI_14_), .ZN(n5039) );
  MUX2_X1 U6602 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .S(n4555), .Z(n5478) );
  INV_X1 U6603 ( .A(n5478), .ZN(n5040) );
  NAND2_X1 U6604 ( .A1(n5041), .A2(n5040), .ZN(n5042) );
  MUX2_X1 U6605 ( .A(n6672), .B(n6674), .S(n4555), .Z(n5492) );
  NOR2_X1 U6606 ( .A1(n5045), .A2(SI_16_), .ZN(n5044) );
  NAND2_X1 U6607 ( .A1(n5045), .A2(SI_16_), .ZN(n5046) );
  MUX2_X1 U6608 ( .A(n6720), .B(n6719), .S(n4555), .Z(n5048) );
  INV_X1 U6609 ( .A(SI_17_), .ZN(n5047) );
  NAND2_X1 U6610 ( .A1(n5048), .A2(n5047), .ZN(n5051) );
  INV_X1 U6611 ( .A(n5048), .ZN(n5049) );
  NAND2_X1 U6612 ( .A1(n5049), .A2(SI_17_), .ZN(n5050) );
  NAND2_X1 U6613 ( .A1(n5051), .A2(n5050), .ZN(n5503) );
  MUX2_X1 U6614 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n4555), .Z(n5052) );
  XNOR2_X1 U6615 ( .A(n5052), .B(n10056), .ZN(n5515) );
  NAND2_X1 U6616 ( .A1(n5053), .A2(n10120), .ZN(n5058) );
  INV_X1 U6617 ( .A(n5053), .ZN(n5054) );
  NAND2_X1 U6618 ( .A1(n5054), .A2(SI_19_), .ZN(n5055) );
  NAND2_X1 U6619 ( .A1(n5058), .A2(n5055), .ZN(n5531) );
  INV_X1 U6620 ( .A(n5531), .ZN(n5056) );
  NAND2_X1 U6621 ( .A1(n5057), .A2(n5056), .ZN(n5059) );
  INV_X1 U6622 ( .A(n5243), .ZN(n5060) );
  NAND2_X1 U6623 ( .A1(n5231), .A2(SI_21_), .ZN(n5061) );
  NAND2_X1 U6624 ( .A1(n5062), .A2(n10103), .ZN(n5065) );
  INV_X1 U6625 ( .A(n5062), .ZN(n5063) );
  NAND2_X1 U6626 ( .A1(n5063), .A2(SI_22_), .ZN(n5064) );
  NAND2_X1 U6627 ( .A1(n5065), .A2(n5064), .ZN(n5205) );
  INV_X1 U6628 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n5066) );
  INV_X1 U6629 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n7640) );
  NAND2_X1 U6630 ( .A1(n5067), .A2(n10097), .ZN(n5070) );
  INV_X1 U6631 ( .A(n5067), .ZN(n5068) );
  NAND2_X1 U6632 ( .A1(n5068), .A2(SI_23_), .ZN(n5069) );
  INV_X1 U6633 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7700) );
  MUX2_X1 U6634 ( .A(n7700), .B(n7701), .S(n4555), .Z(n5072) );
  INV_X1 U6635 ( .A(SI_24_), .ZN(n10141) );
  NAND2_X1 U6636 ( .A1(n5072), .A2(n10141), .ZN(n5075) );
  INV_X1 U6637 ( .A(n5072), .ZN(n5073) );
  NAND2_X1 U6638 ( .A1(n5073), .A2(SI_24_), .ZN(n5074) );
  NAND2_X1 U6639 ( .A1(n5181), .A2(n5180), .ZN(n5076) );
  NAND2_X1 U6640 ( .A1(n5076), .A2(n5075), .ZN(n5219) );
  INV_X1 U6641 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7742) );
  INV_X1 U6642 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7739) );
  INV_X1 U6643 ( .A(SI_25_), .ZN(n10146) );
  NAND2_X1 U6644 ( .A1(n5077), .A2(n10146), .ZN(n5080) );
  INV_X1 U6645 ( .A(n5077), .ZN(n5078) );
  NAND2_X1 U6646 ( .A1(n5078), .A2(SI_25_), .ZN(n5079) );
  INV_X1 U6647 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n5082) );
  INV_X1 U6648 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n7784) );
  INV_X1 U6649 ( .A(SI_26_), .ZN(n10131) );
  NAND2_X1 U6650 ( .A1(n5083), .A2(n10131), .ZN(n5086) );
  INV_X1 U6651 ( .A(n5083), .ZN(n5084) );
  NAND2_X1 U6652 ( .A1(n5084), .A2(SI_26_), .ZN(n5085) );
  INV_X1 U6653 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n5088) );
  INV_X1 U6654 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n9486) );
  INV_X1 U6655 ( .A(SI_27_), .ZN(n10115) );
  NAND2_X1 U6656 ( .A1(n5089), .A2(n10115), .ZN(n5092) );
  INV_X1 U6657 ( .A(n5089), .ZN(n5090) );
  NAND2_X1 U6658 ( .A1(n5090), .A2(SI_27_), .ZN(n5091) );
  INV_X1 U6659 ( .A(SI_28_), .ZN(n10112) );
  XNOR2_X1 U6660 ( .A(n5094), .B(n10112), .ZN(n5152) );
  INV_X1 U6661 ( .A(n5094), .ZN(n5095) );
  NAND2_X1 U6662 ( .A1(n5095), .A2(n10112), .ZN(n5096) );
  INV_X1 U6663 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n5098) );
  INV_X1 U6664 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n7868) );
  INV_X1 U6665 ( .A(SI_29_), .ZN(n10047) );
  INV_X1 U6666 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n5102) );
  INV_X1 U6667 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n9482) );
  INV_X1 U6668 ( .A(SI_30_), .ZN(n10117) );
  NAND2_X1 U6669 ( .A1(n5103), .A2(n10117), .ZN(n5562) );
  INV_X1 U6670 ( .A(n5103), .ZN(n5104) );
  NAND2_X1 U6671 ( .A1(n5104), .A2(SI_30_), .ZN(n5105) );
  NAND2_X1 U6672 ( .A1(n5562), .A2(n5105), .ZN(n5563) );
  NOR2_X2 U6673 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5298) );
  NOR2_X1 U6674 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), .ZN(
        n5119) );
  NOR2_X1 U6675 ( .A1(P1_IR_REG_24__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), .ZN(
        n5118) );
  NOR2_X1 U6676 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .ZN(
        n5117) );
  INV_X1 U6677 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n5124) );
  INV_X1 U6678 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5125) );
  NAND2_X1 U6679 ( .A1(n5126), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5128) );
  INV_X1 U6680 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5127) );
  INV_X2 U6681 ( .A(n5296), .ZN(n5517) );
  NAND2_X1 U6682 ( .A1(n8768), .A2(n5517), .ZN(n5130) );
  OR2_X1 U6683 ( .A1(n5297), .A2(n9482), .ZN(n5129) );
  INV_X1 U6684 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n9308) );
  INV_X1 U6685 ( .A(n9470), .ZN(n5132) );
  NOR2_X1 U6686 ( .A1(P1_IR_REG_29__SCAN_IN), .A2(P1_IR_REG_28__SCAN_IN), .ZN(
        n5131) );
  AOI21_X1 U6687 ( .B1(n5132), .B2(n5131), .A(n5124), .ZN(n5133) );
  INV_X1 U6688 ( .A(n5133), .ZN(n5134) );
  NAND2_X1 U6689 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_28__SCAN_IN), 
        .ZN(n5135) );
  NAND2_X1 U6690 ( .A1(n5136), .A2(n5135), .ZN(n5137) );
  XNOR2_X2 U6691 ( .A(n5137), .B(n9471), .ZN(n5138) );
  INV_X4 U6692 ( .A(n5199), .ZN(n5556) );
  NAND2_X1 U6693 ( .A1(n5556), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n5140) );
  AND2_X2 U6694 ( .A1(n9478), .A2(n7867), .ZN(n5278) );
  NAND2_X1 U6695 ( .A1(n5427), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n5139) );
  OAI211_X1 U6696 ( .C1(n9308), .C2(n5559), .A(n5140), .B(n5139), .ZN(n9088)
         );
  NAND2_X1 U6697 ( .A1(n7866), .A2(n5517), .ZN(n5143) );
  OR2_X1 U6698 ( .A1(n5297), .A2(n7868), .ZN(n5142) );
  INV_X4 U6699 ( .A(n5559), .ZN(n5545) );
  NAND2_X1 U6700 ( .A1(n5545), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n5145) );
  NAND2_X1 U6701 ( .A1(n5427), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n5144) );
  AND2_X1 U6702 ( .A1(n5145), .A2(n5144), .ZN(n5150) );
  INV_X2 U6703 ( .A(n5288), .ZN(n5549) );
  NAND2_X1 U6704 ( .A1(n5315), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n5344) );
  INV_X1 U6705 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n5343) );
  NOR2_X1 U6706 ( .A1(n5344), .A2(n5343), .ZN(n5342) );
  NAND2_X1 U6707 ( .A1(n5342), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5389) );
  INV_X1 U6708 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n5388) );
  NAND2_X1 U6709 ( .A1(n5412), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5440) );
  INV_X1 U6710 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n5439) );
  INV_X1 U6711 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n5456) );
  INV_X1 U6712 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n5472) );
  NAND2_X1 U6713 ( .A1(n8870), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n5525) );
  INV_X1 U6714 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n5524) );
  NAND2_X1 U6715 ( .A1(P1_REG3_REG_20__SCAN_IN), .A2(P1_REG3_REG_19__SCAN_IN), 
        .ZN(n5146) );
  INV_X1 U6716 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n8800) );
  NAND2_X1 U6717 ( .A1(n5174), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n5177) );
  INV_X1 U6718 ( .A(n5177), .ZN(n5147) );
  NAND2_X1 U6719 ( .A1(n5155), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n5158) );
  INV_X1 U6720 ( .A(n5158), .ZN(n9124) );
  NAND2_X1 U6721 ( .A1(n5549), .A2(n9124), .ZN(n5149) );
  NAND2_X1 U6722 ( .A1(n5556), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n5148) );
  NAND2_X1 U6723 ( .A1(n7889), .A2(n5517), .ZN(n5154) );
  INV_X1 U6724 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n7890) );
  OR2_X1 U6725 ( .A1(n5297), .A2(n7890), .ZN(n5153) );
  AOI22_X1 U6726 ( .A1(n5556), .A2(P1_REG2_REG_28__SCAN_IN), .B1(n5545), .B2(
        P1_REG1_REG_28__SCAN_IN), .ZN(n5160) );
  INV_X1 U6727 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n5156) );
  NAND2_X1 U6728 ( .A1(n5167), .A2(n5156), .ZN(n5157) );
  AOI22_X1 U6729 ( .A1(n5549), .A2(n9135), .B1(n5427), .B2(
        P1_REG0_REG_28__SCAN_IN), .ZN(n5159) );
  NAND2_X1 U6730 ( .A1(n5716), .A2(n5712), .ZN(n5785) );
  NAND2_X1 U6731 ( .A1(n9318), .A2(n9325), .ZN(n9119) );
  NAND2_X1 U6732 ( .A1(n7805), .A2(n5517), .ZN(n5164) );
  OR2_X1 U6733 ( .A1(n5297), .A2(n9486), .ZN(n5163) );
  AOI22_X1 U6734 ( .A1(n5556), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n5545), .B2(
        P1_REG1_REG_27__SCAN_IN), .ZN(n5169) );
  INV_X1 U6735 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n5165) );
  NAND2_X1 U6736 ( .A1(n5177), .A2(n5165), .ZN(n5166) );
  AOI22_X1 U6737 ( .A1(n5549), .A2(n9148), .B1(n5427), .B2(
        P1_REG0_REG_27__SCAN_IN), .ZN(n5168) );
  NAND2_X1 U6738 ( .A1(n9156), .A2(n9335), .ZN(n9118) );
  AND2_X1 U6739 ( .A1(n9119), .A2(n9118), .ZN(n5709) );
  INV_X1 U6740 ( .A(n5709), .ZN(n5262) );
  NAND2_X1 U6741 ( .A1(n7744), .A2(n5517), .ZN(n5173) );
  OR2_X1 U6742 ( .A1(n5297), .A2(n7784), .ZN(n5172) );
  AOI22_X1 U6743 ( .A1(n5556), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n5545), .B2(
        P1_REG1_REG_26__SCAN_IN), .ZN(n5179) );
  INV_X1 U6744 ( .A(n5174), .ZN(n5226) );
  INV_X1 U6745 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n5175) );
  NAND2_X1 U6746 ( .A1(n5226), .A2(n5175), .ZN(n5176) );
  AND2_X1 U6747 ( .A1(n5177), .A2(n5176), .ZN(n9165) );
  AOI22_X1 U6748 ( .A1(n5549), .A2(n9165), .B1(n5427), .B2(
        P1_REG0_REG_26__SCAN_IN), .ZN(n5178) );
  OR2_X1 U6749 ( .A1(n9164), .A2(n9324), .ZN(n5584) );
  XNOR2_X1 U6750 ( .A(n5181), .B(n5180), .ZN(n7699) );
  NAND2_X1 U6751 ( .A1(n7699), .A2(n5517), .ZN(n5183) );
  OR2_X1 U6752 ( .A1(n5297), .A2(n7701), .ZN(n5182) );
  NAND2_X1 U6753 ( .A1(n5545), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n5185) );
  NAND2_X1 U6754 ( .A1(n5427), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n5184) );
  AND2_X1 U6755 ( .A1(n5185), .A2(n5184), .ZN(n5192) );
  INV_X1 U6756 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n5187) );
  INV_X1 U6757 ( .A(n5186), .ZN(n5197) );
  NAND2_X1 U6758 ( .A1(n5187), .A2(n5197), .ZN(n5189) );
  INV_X1 U6759 ( .A(n5188), .ZN(n5224) );
  AND2_X1 U6760 ( .A1(n5189), .A2(n5224), .ZN(n9202) );
  NAND2_X1 U6761 ( .A1(n5549), .A2(n9202), .ZN(n5191) );
  NAND2_X1 U6762 ( .A1(n5556), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n5190) );
  NAND2_X1 U6763 ( .A1(n9201), .A2(n9360), .ZN(n5700) );
  NAND2_X1 U6764 ( .A1(n7637), .A2(n5517), .ZN(n5196) );
  OR2_X1 U6765 ( .A1(n5297), .A2(n7640), .ZN(n5195) );
  NAND2_X1 U6766 ( .A1(n5210), .A2(n8800), .ZN(n5198) );
  NAND2_X1 U6767 ( .A1(n5198), .A2(n5197), .ZN(n9213) );
  OR2_X1 U6768 ( .A1(n9213), .A2(n5288), .ZN(n5204) );
  INV_X1 U6769 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n9214) );
  NAND2_X1 U6770 ( .A1(n5545), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n5201) );
  NAND2_X1 U6771 ( .A1(n5278), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n5200) );
  OAI211_X1 U6772 ( .C1(n5199), .C2(n9214), .A(n5201), .B(n5200), .ZN(n5202)
         );
  INV_X1 U6773 ( .A(n5202), .ZN(n5203) );
  NAND2_X1 U6774 ( .A1(n9363), .A2(n9199), .ZN(n9192) );
  OR2_X1 U6775 ( .A1(n9363), .A2(n9199), .ZN(n5696) );
  XNOR2_X1 U6776 ( .A(n5206), .B(n5205), .ZN(n7545) );
  NAND2_X1 U6777 ( .A1(n7545), .A2(n5517), .ZN(n5208) );
  OR2_X1 U6778 ( .A1(n5297), .A2(n7888), .ZN(n5207) );
  OR2_X1 U6779 ( .A1(n5236), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n5209) );
  AND2_X1 U6780 ( .A1(n5210), .A2(n5209), .ZN(n9227) );
  NAND2_X1 U6781 ( .A1(n9227), .A2(n5549), .ZN(n5215) );
  INV_X1 U6782 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n9229) );
  NAND2_X1 U6783 ( .A1(n5427), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n5212) );
  NAND2_X1 U6784 ( .A1(n5545), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n5211) );
  OAI211_X1 U6785 ( .C1(n5199), .C2(n9229), .A(n5212), .B(n5211), .ZN(n5213)
         );
  INV_X1 U6786 ( .A(n5213), .ZN(n5214) );
  OR2_X1 U6787 ( .A1(n9233), .A2(n9361), .ZN(n5216) );
  NAND2_X1 U6788 ( .A1(n5696), .A2(n5216), .ZN(n5613) );
  NAND3_X1 U6789 ( .A1(n5700), .A2(n9192), .A3(n5613), .ZN(n5217) );
  AND2_X1 U6790 ( .A1(n5217), .A2(n9176), .ZN(n5264) );
  XNOR2_X1 U6791 ( .A(n5219), .B(n5218), .ZN(n7738) );
  NAND2_X1 U6792 ( .A1(n7738), .A2(n5517), .ZN(n5221) );
  OR2_X1 U6793 ( .A1(n5297), .A2(n7739), .ZN(n5220) );
  NAND2_X1 U6794 ( .A1(n5545), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n5223) );
  NAND2_X1 U6795 ( .A1(n5427), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n5222) );
  AND2_X1 U6796 ( .A1(n5223), .A2(n5222), .ZN(n5229) );
  INV_X1 U6797 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n8845) );
  NAND2_X1 U6798 ( .A1(n5224), .A2(n8845), .ZN(n5225) );
  AND2_X1 U6799 ( .A1(n5226), .A2(n5225), .ZN(n8846) );
  NAND2_X1 U6800 ( .A1(n5549), .A2(n8846), .ZN(n5228) );
  NAND2_X1 U6801 ( .A1(n5556), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n5227) );
  OR2_X1 U6802 ( .A1(n9185), .A2(n9334), .ZN(n5585) );
  INV_X1 U6803 ( .A(SI_21_), .ZN(n5230) );
  XNOR2_X1 U6804 ( .A(n5231), .B(n5230), .ZN(n5232) );
  XNOR2_X1 U6805 ( .A(n5233), .B(n5232), .ZN(n7407) );
  NAND2_X1 U6806 ( .A1(n7407), .A2(n5517), .ZN(n5235) );
  INV_X1 U6807 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7447) );
  OR2_X1 U6808 ( .A1(n5297), .A2(n7447), .ZN(n5234) );
  INV_X1 U6809 ( .A(n5236), .ZN(n5239) );
  INV_X1 U6810 ( .A(n5237), .ZN(n5249) );
  INV_X1 U6811 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n8830) );
  NAND2_X1 U6812 ( .A1(n5249), .A2(n8830), .ZN(n5238) );
  AND2_X1 U6813 ( .A1(n5239), .A2(n5238), .ZN(n8831) );
  NAND2_X1 U6814 ( .A1(n8831), .A2(n5549), .ZN(n5242) );
  AOI22_X1 U6815 ( .A1(n5556), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n5545), .B2(
        P1_REG1_REG_21__SCAN_IN), .ZN(n5241) );
  NAND2_X1 U6816 ( .A1(n5427), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n5240) );
  OR2_X1 U6817 ( .A1(n9241), .A2(n9255), .ZN(n5263) );
  INV_X1 U6818 ( .A(n5263), .ZN(n5692) );
  NAND2_X1 U6819 ( .A1(n9241), .A2(n9255), .ZN(n9113) );
  XNOR2_X1 U6820 ( .A(n5243), .B(n10080), .ZN(n5244) );
  XNOR2_X1 U6821 ( .A(n5245), .B(n5244), .ZN(n7381) );
  NAND2_X1 U6822 ( .A1(n7381), .A2(n5517), .ZN(n5247) );
  INV_X1 U6823 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7382) );
  OR2_X1 U6824 ( .A1(n5297), .A2(n7382), .ZN(n5246) );
  INV_X1 U6825 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n5248) );
  INV_X1 U6826 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n8890) );
  OAI21_X1 U6827 ( .B1(n5548), .B2(n5248), .A(n8890), .ZN(n5250) );
  NAND2_X1 U6828 ( .A1(n5250), .A2(n5249), .ZN(n9259) );
  OR2_X1 U6829 ( .A1(n5288), .A2(n9259), .ZN(n5255) );
  NAND2_X1 U6830 ( .A1(n5545), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n5252) );
  NAND2_X1 U6831 ( .A1(n5427), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n5251) );
  AND2_X1 U6832 ( .A1(n5252), .A2(n5251), .ZN(n5254) );
  NAND2_X1 U6833 ( .A1(n5556), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n5253) );
  NAND2_X1 U6834 ( .A1(n9388), .A2(n9278), .ZN(n9112) );
  NAND2_X1 U6835 ( .A1(n9113), .A2(n9112), .ZN(n5691) );
  INV_X1 U6836 ( .A(n5691), .ZN(n5257) );
  NAND2_X1 U6837 ( .A1(n9233), .A2(n9361), .ZN(n9114) );
  NAND2_X1 U6838 ( .A1(n9192), .A2(n9114), .ZN(n5612) );
  INV_X1 U6839 ( .A(n5612), .ZN(n5256) );
  OAI211_X1 U6840 ( .C1(n5692), .C2(n5257), .A(n5700), .B(n5256), .ZN(n5258)
         );
  NAND3_X1 U6841 ( .A1(n5264), .A2(n5585), .A3(n5258), .ZN(n5259) );
  INV_X1 U6842 ( .A(n9116), .ZN(n5703) );
  NAND2_X1 U6843 ( .A1(n5259), .A2(n5703), .ZN(n5260) );
  AND3_X1 U6844 ( .A1(n5780), .A2(n5584), .A3(n5260), .ZN(n5261) );
  OR2_X1 U6845 ( .A1(n5262), .A2(n5261), .ZN(n5783) );
  AND2_X1 U6846 ( .A1(n5584), .A2(n5585), .ZN(n5704) );
  INV_X1 U6847 ( .A(n5704), .ZN(n5266) );
  OR2_X1 U6848 ( .A1(n9388), .A2(n9278), .ZN(n5688) );
  NAND2_X1 U6849 ( .A1(n5263), .A2(n5688), .ZN(n5614) );
  INV_X1 U6850 ( .A(n5264), .ZN(n5265) );
  OR3_X1 U6851 ( .A1(n5266), .A2(n5614), .A3(n5265), .ZN(n5779) );
  INV_X1 U6852 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n5268) );
  NAND2_X1 U6853 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5267) );
  XNOR2_X1 U6854 ( .A(n5270), .B(n5269), .ZN(n6175) );
  INV_X1 U6855 ( .A(n6175), .ZN(n6595) );
  INV_X1 U6856 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6588) );
  OR2_X1 U6857 ( .A1(n4373), .A2(n6588), .ZN(n5271) );
  NAND2_X1 U6858 ( .A1(n5289), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5275) );
  NAND2_X1 U6859 ( .A1(n5278), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n5274) );
  NAND2_X1 U6860 ( .A1(n5276), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5273) );
  NAND2_X1 U6861 ( .A1(n4372), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n5282) );
  NAND2_X1 U6862 ( .A1(n5277), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n5281) );
  NAND2_X1 U6863 ( .A1(n5289), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5280) );
  NAND2_X1 U6864 ( .A1(n5278), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5279) );
  NAND4_X2 U6865 ( .A1(n5282), .A2(n5281), .A3(n5280), .A4(n5279), .ZN(n8822)
         );
  INV_X1 U6866 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n9544) );
  INV_X1 U6867 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5283) );
  NAND2_X1 U6868 ( .A1(n5284), .A2(n5283), .ZN(n5286) );
  NAND2_X1 U6869 ( .A1(n5286), .A2(n5285), .ZN(n9488) );
  MUX2_X1 U6870 ( .A(n9544), .B(n9488), .S(n6622), .Z(n6942) );
  NOR2_X1 U6871 ( .A1(n8822), .A2(n6942), .ZN(n6935) );
  INV_X1 U6872 ( .A(n9719), .ZN(n6680) );
  NAND2_X1 U6873 ( .A1(n6680), .A2(n8823), .ZN(n5287) );
  NAND2_X1 U6874 ( .A1(n5277), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n5293) );
  NAND2_X1 U6875 ( .A1(n4372), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5292) );
  NAND2_X1 U6876 ( .A1(n5289), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5291) );
  NAND2_X1 U6877 ( .A1(n5278), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5290) );
  XNOR2_X1 U6878 ( .A(n5295), .B(n5294), .ZN(n6193) );
  INV_X1 U6879 ( .A(n6193), .ZN(n6602) );
  OR2_X1 U6880 ( .A1(n5296), .A2(n6602), .ZN(n5302) );
  INV_X1 U6881 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6603) );
  OR2_X1 U6882 ( .A1(n4374), .A2(n6603), .ZN(n5301) );
  INV_X4 U6883 ( .A(n6622), .ZN(n5541) );
  OR2_X1 U6884 ( .A1(n5298), .A2(n5124), .ZN(n5299) );
  NAND2_X1 U6885 ( .A1(n5541), .A2(n9560), .ZN(n5300) );
  AND3_X2 U6886 ( .A1(n5302), .A2(n5301), .A3(n5300), .ZN(n9726) );
  NAND2_X1 U6887 ( .A1(n8962), .A2(n9726), .ZN(n5619) );
  INV_X1 U6888 ( .A(n8962), .ZN(n6936) );
  NAND2_X1 U6889 ( .A1(n6936), .A2(n6757), .ZN(n5617) );
  INV_X1 U6890 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n5303) );
  NAND2_X1 U6891 ( .A1(n5277), .A2(n5303), .ZN(n5307) );
  NAND2_X1 U6892 ( .A1(n4372), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5306) );
  NAND2_X1 U6893 ( .A1(n5289), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n5305) );
  NAND2_X1 U6894 ( .A1(n5278), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5304) );
  NAND4_X2 U6895 ( .A1(n5307), .A2(n5306), .A3(n5305), .A4(n5304), .ZN(n8961)
         );
  XNOR2_X1 U6896 ( .A(n5309), .B(n5308), .ZN(n6208) );
  INV_X1 U6897 ( .A(n6208), .ZN(n6597) );
  OR2_X1 U6898 ( .A1(n5296), .A2(n6597), .ZN(n5314) );
  INV_X1 U6899 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6590) );
  OR2_X1 U6900 ( .A1(n4374), .A2(n6590), .ZN(n5313) );
  NAND2_X1 U6901 ( .A1(n5310), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5311) );
  XNOR2_X1 U6902 ( .A(n5311), .B(P1_IR_REG_3__SCAN_IN), .ZN(n9009) );
  NAND2_X1 U6903 ( .A1(n5541), .A2(n9009), .ZN(n5312) );
  AND3_X2 U6904 ( .A1(n5314), .A2(n5313), .A3(n5312), .ZN(n6954) );
  NAND2_X1 U6905 ( .A1(n8961), .A2(n6954), .ZN(n5626) );
  AOI22_X1 U6906 ( .A1(n4372), .A2(P1_REG2_REG_4__SCAN_IN), .B1(n5545), .B2(
        P1_REG1_REG_4__SCAN_IN), .ZN(n5318) );
  INV_X1 U6907 ( .A(n5315), .ZN(n5328) );
  OAI21_X1 U6908 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(n5328), .ZN(n6726) );
  INV_X1 U6909 ( .A(n6726), .ZN(n5316) );
  AOI22_X1 U6910 ( .A1(n5549), .A2(n5316), .B1(n5278), .B2(
        P1_REG0_REG_4__SCAN_IN), .ZN(n5317) );
  NAND2_X1 U6911 ( .A1(n5319), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5321) );
  OR2_X1 U6912 ( .A1(n5321), .A2(n5320), .ZN(n5322) );
  NAND2_X1 U6913 ( .A1(n5321), .A2(n5320), .ZN(n5336) );
  INV_X1 U6914 ( .A(n9013), .ZN(n9579) );
  XNOR2_X1 U6915 ( .A(n5324), .B(n5323), .ZN(n6604) );
  OR2_X1 U6916 ( .A1(n5296), .A2(n6604), .ZN(n5326) );
  OR2_X1 U6917 ( .A1(n5297), .A2(n6605), .ZN(n5325) );
  OAI211_X1 U6918 ( .C1(n6622), .C2(n9579), .A(n5326), .B(n5325), .ZN(n6727)
         );
  INV_X1 U6919 ( .A(n6727), .ZN(n6867) );
  NAND2_X1 U6920 ( .A1(n6703), .A2(n5738), .ZN(n6768) );
  NAND2_X1 U6921 ( .A1(n6833), .A2(n6727), .ZN(n6767) );
  NAND2_X1 U6922 ( .A1(n6768), .A2(n6767), .ZN(n5341) );
  NAND2_X1 U6923 ( .A1(n4372), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n5333) );
  INV_X1 U6924 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n5327) );
  NAND2_X1 U6925 ( .A1(n5328), .A2(n5327), .ZN(n5329) );
  AND2_X1 U6926 ( .A1(n5344), .A2(n5329), .ZN(n6832) );
  NAND2_X1 U6927 ( .A1(n5549), .A2(n6832), .ZN(n5332) );
  NAND2_X1 U6928 ( .A1(n5545), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5331) );
  NAND2_X1 U6929 ( .A1(n5278), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n5330) );
  NAND4_X1 U6930 ( .A1(n5333), .A2(n5332), .A3(n5331), .A4(n5330), .ZN(n8959)
         );
  XNOR2_X1 U6931 ( .A(n5335), .B(n5334), .ZN(n6594) );
  OR2_X1 U6932 ( .A1(n5296), .A2(n6594), .ZN(n5340) );
  INV_X1 U6933 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6592) );
  OR2_X1 U6934 ( .A1(n5297), .A2(n6592), .ZN(n5339) );
  NAND2_X1 U6935 ( .A1(n5336), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5337) );
  XNOR2_X1 U6936 ( .A(n5337), .B(P1_IR_REG_5__SCAN_IN), .ZN(n9017) );
  NAND2_X1 U6937 ( .A1(n5541), .A2(n9017), .ZN(n5338) );
  NOR2_X1 U6938 ( .A1(n8959), .A2(n6857), .ZN(n5622) );
  INV_X1 U6939 ( .A(n5622), .ZN(n5627) );
  NAND2_X1 U6940 ( .A1(n8959), .A2(n6857), .ZN(n5743) );
  AND2_X1 U6941 ( .A1(n5627), .A2(n5743), .ZN(n6766) );
  NAND2_X1 U6942 ( .A1(n5341), .A2(n6766), .ZN(n6770) );
  NAND2_X1 U6943 ( .A1(n6770), .A2(n5627), .ZN(n6784) );
  NAND2_X1 U6944 ( .A1(n4372), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n5349) );
  INV_X1 U6945 ( .A(n5342), .ZN(n5375) );
  NAND2_X1 U6946 ( .A1(n5344), .A2(n5343), .ZN(n5345) );
  AND2_X1 U6947 ( .A1(n5375), .A2(n5345), .ZN(n7034) );
  NAND2_X1 U6948 ( .A1(n5549), .A2(n7034), .ZN(n5348) );
  NAND2_X1 U6949 ( .A1(n5545), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n5347) );
  NAND2_X1 U6950 ( .A1(n5278), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5346) );
  NAND4_X1 U6951 ( .A1(n5349), .A2(n5348), .A3(n5347), .A4(n5346), .ZN(n8958)
         );
  INV_X1 U6952 ( .A(n8958), .ZN(n7263) );
  XNOR2_X1 U6953 ( .A(n5351), .B(n5350), .ZN(n6596) );
  NAND2_X1 U6954 ( .A1(n5517), .A2(n6596), .ZN(n5359) );
  NOR2_X1 U6955 ( .A1(n5352), .A2(n5124), .ZN(n5353) );
  MUX2_X1 U6956 ( .A(n5124), .B(n5353), .S(P1_IR_REG_6__SCAN_IN), .Z(n5356) );
  INV_X1 U6957 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5354) );
  NAND2_X1 U6958 ( .A1(n5352), .A2(n5354), .ZN(n5382) );
  INV_X1 U6959 ( .A(n5382), .ZN(n5355) );
  NAND2_X1 U6960 ( .A1(n5541), .A2(n9019), .ZN(n5358) );
  INV_X1 U6961 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6600) );
  OR2_X1 U6962 ( .A1(n5297), .A2(n6600), .ZN(n5357) );
  NAND2_X1 U6963 ( .A1(n7263), .A2(n7037), .ZN(n5746) );
  INV_X1 U6964 ( .A(n5746), .ZN(n5631) );
  XNOR2_X1 U6965 ( .A(n5360), .B(n4982), .ZN(n6613) );
  NAND2_X1 U6966 ( .A1(n6613), .A2(n5517), .ZN(n5364) );
  NAND2_X1 U6967 ( .A1(n5408), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5397) );
  INV_X1 U6968 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n5406) );
  NAND2_X1 U6969 ( .A1(n5397), .A2(n5406), .ZN(n5361) );
  NAND2_X1 U6970 ( .A1(n5361), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5362) );
  XNOR2_X1 U6971 ( .A(n5362), .B(P1_IR_REG_9__SCAN_IN), .ZN(n9045) );
  AOI22_X1 U6972 ( .A1(n5542), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n5541), .B2(
        n9045), .ZN(n5363) );
  NAND2_X1 U6973 ( .A1(n5545), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n5366) );
  NAND2_X1 U6974 ( .A1(n5427), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5365) );
  AND2_X1 U6975 ( .A1(n5366), .A2(n5365), .ZN(n5371) );
  INV_X1 U6976 ( .A(n5367), .ZN(n5414) );
  NAND2_X1 U6977 ( .A1(n5391), .A2(n7645), .ZN(n5368) );
  AND2_X1 U6978 ( .A1(n5414), .A2(n5368), .ZN(n7646) );
  NAND2_X1 U6979 ( .A1(n5549), .A2(n7646), .ZN(n5370) );
  NAND2_X1 U6980 ( .A1(n5556), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5369) );
  NAND2_X1 U6981 ( .A1(n9747), .A2(n7473), .ZN(n7429) );
  INV_X1 U6982 ( .A(n7429), .ZN(n5592) );
  NAND2_X1 U6983 ( .A1(n5545), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5373) );
  NAND2_X1 U6984 ( .A1(n5427), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5372) );
  AND2_X1 U6985 ( .A1(n5373), .A2(n5372), .ZN(n5379) );
  INV_X1 U6986 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n5374) );
  NAND2_X1 U6987 ( .A1(n5375), .A2(n5374), .ZN(n5376) );
  AND2_X1 U6988 ( .A1(n5389), .A2(n5376), .ZN(n7270) );
  NAND2_X1 U6989 ( .A1(n5549), .A2(n7270), .ZN(n5378) );
  NAND2_X1 U6990 ( .A1(n5556), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n5377) );
  XNOR2_X1 U6991 ( .A(n5381), .B(n5380), .ZN(n6607) );
  OR2_X1 U6992 ( .A1(n6607), .A2(n5296), .ZN(n5385) );
  NAND2_X1 U6993 ( .A1(n5382), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5383) );
  XNOR2_X1 U6994 ( .A(n5383), .B(P1_IR_REG_7__SCAN_IN), .ZN(n9022) );
  AOI22_X1 U6995 ( .A1(n5542), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n5541), .B2(
        n9022), .ZN(n5384) );
  NAND2_X1 U6996 ( .A1(n5385), .A2(n5384), .ZN(n7271) );
  NAND2_X1 U6997 ( .A1(n7311), .A2(n7271), .ZN(n7307) );
  NAND2_X1 U6998 ( .A1(n5545), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5387) );
  NAND2_X1 U6999 ( .A1(n5427), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n5386) );
  AND2_X1 U7000 ( .A1(n5387), .A2(n5386), .ZN(n5394) );
  NAND2_X1 U7001 ( .A1(n5389), .A2(n5388), .ZN(n5390) );
  AND2_X1 U7002 ( .A1(n5391), .A2(n5390), .ZN(n7549) );
  NAND2_X1 U7003 ( .A1(n5549), .A2(n7549), .ZN(n5393) );
  NAND2_X1 U7004 ( .A1(n5556), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n5392) );
  XNOR2_X1 U7005 ( .A(n5396), .B(n5395), .ZN(n6609) );
  NAND2_X1 U7006 ( .A1(n6609), .A2(n5517), .ZN(n5399) );
  XNOR2_X1 U7007 ( .A(n5397), .B(P1_IR_REG_8__SCAN_IN), .ZN(n9025) );
  AOI22_X1 U7008 ( .A1(n5542), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n5541), .B2(
        n9025), .ZN(n5398) );
  NAND2_X1 U7009 ( .A1(n7439), .A2(n7437), .ZN(n7431) );
  NAND2_X1 U7010 ( .A1(n7307), .A2(n7431), .ZN(n5638) );
  OR2_X1 U7011 ( .A1(n7473), .A2(n9747), .ZN(n7430) );
  NAND2_X1 U7012 ( .A1(n4596), .A2(n9746), .ZN(n7432) );
  NAND2_X1 U7013 ( .A1(n7430), .A2(n7432), .ZN(n5643) );
  INV_X1 U7014 ( .A(n5643), .ZN(n5400) );
  AOI21_X1 U7015 ( .B1(n5400), .B2(n5638), .A(n5592), .ZN(n5747) );
  INV_X1 U7016 ( .A(n7311), .ZN(n8957) );
  NAND2_X1 U7017 ( .A1(n8957), .A2(n7425), .ZN(n5636) );
  INV_X1 U7018 ( .A(n5636), .ZN(n5401) );
  NAND2_X1 U7019 ( .A1(n8958), .A2(n9733), .ZN(n7264) );
  NAND2_X1 U7020 ( .A1(n5595), .A2(n7264), .ZN(n5402) );
  NAND2_X1 U7021 ( .A1(n5747), .A2(n5402), .ZN(n5750) );
  XNOR2_X1 U7022 ( .A(n5404), .B(n5403), .ZN(n6615) );
  NAND2_X1 U7023 ( .A1(n6615), .A2(n5517), .ZN(n5411) );
  INV_X1 U7024 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n5405) );
  NAND2_X1 U7025 ( .A1(n5406), .A2(n5405), .ZN(n5407) );
  NAND2_X1 U7026 ( .A1(n5420), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5409) );
  XNOR2_X1 U7027 ( .A(n5409), .B(P1_IR_REG_10__SCAN_IN), .ZN(n9498) );
  AOI22_X1 U7028 ( .A1(n5542), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n5541), .B2(
        n9498), .ZN(n5410) );
  NAND2_X1 U7029 ( .A1(n5411), .A2(n5410), .ZN(n7513) );
  AOI22_X1 U7030 ( .A1(n5556), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n5545), .B2(
        P1_REG1_REG_10__SCAN_IN), .ZN(n5417) );
  INV_X1 U7031 ( .A(n5412), .ZN(n5425) );
  INV_X1 U7032 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n5413) );
  NAND2_X1 U7033 ( .A1(n5414), .A2(n5413), .ZN(n5415) );
  AND2_X1 U7034 ( .A1(n5425), .A2(n5415), .ZN(n7762) );
  AOI22_X1 U7035 ( .A1(n5549), .A2(n7762), .B1(n5427), .B2(
        P1_REG0_REG_10__SCAN_IN), .ZN(n5416) );
  OR2_X1 U7036 ( .A1(n7513), .A2(n7814), .ZN(n5749) );
  NAND2_X1 U7037 ( .A1(n7513), .A2(n7814), .ZN(n7516) );
  NAND2_X1 U7038 ( .A1(n6628), .A2(n5517), .ZN(n5423) );
  NOR2_X1 U7039 ( .A1(n5420), .A2(P1_IR_REG_10__SCAN_IN), .ZN(n5435) );
  OR2_X1 U7040 ( .A1(n5435), .A2(n5124), .ZN(n5421) );
  XNOR2_X1 U7041 ( .A(n5421), .B(P1_IR_REG_11__SCAN_IN), .ZN(n9047) );
  AOI22_X1 U7042 ( .A1(n5542), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n5541), .B2(
        n9047), .ZN(n5422) );
  NAND2_X1 U7043 ( .A1(n5423), .A2(n5422), .ZN(n7816) );
  AOI22_X1 U7044 ( .A1(n5556), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n5545), .B2(
        P1_REG1_REG_11__SCAN_IN), .ZN(n5429) );
  INV_X1 U7045 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n5424) );
  NAND2_X1 U7046 ( .A1(n5425), .A2(n5424), .ZN(n5426) );
  AND2_X1 U7047 ( .A1(n5440), .A2(n5426), .ZN(n7812) );
  AOI22_X1 U7048 ( .A1(n5549), .A2(n7812), .B1(n5427), .B2(
        P1_REG0_REG_11__SCAN_IN), .ZN(n5428) );
  NAND2_X1 U7049 ( .A1(n7816), .A2(n9777), .ZN(n5656) );
  INV_X1 U7050 ( .A(n7516), .ZN(n5430) );
  NOR2_X1 U7051 ( .A1(n7623), .A2(n5430), .ZN(n5431) );
  XNOR2_X1 U7052 ( .A(n5433), .B(n5432), .ZN(n6632) );
  NAND2_X1 U7053 ( .A1(n6632), .A2(n5517), .ZN(n5438) );
  INV_X1 U7054 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n5434) );
  NAND2_X1 U7055 ( .A1(n5435), .A2(n5434), .ZN(n5436) );
  NAND2_X1 U7056 ( .A1(n5436), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5449) );
  XNOR2_X1 U7057 ( .A(n5449), .B(n4366), .ZN(n9629) );
  AOI22_X1 U7058 ( .A1(n5542), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n5541), .B2(
        n9629), .ZN(n5437) );
  AOI22_X1 U7059 ( .A1(n5556), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n5545), .B2(
        P1_REG1_REG_12__SCAN_IN), .ZN(n5443) );
  NAND2_X1 U7060 ( .A1(n5440), .A2(n5439), .ZN(n5441) );
  AND2_X1 U7061 ( .A1(n5457), .A2(n5441), .ZN(n8838) );
  AOI22_X1 U7062 ( .A1(n5549), .A2(n8838), .B1(n5278), .B2(
        P1_REG0_REG_12__SCAN_IN), .ZN(n5442) );
  NOR2_X1 U7063 ( .A1(n9780), .A2(n7689), .ZN(n5653) );
  INV_X1 U7064 ( .A(n5653), .ZN(n5658) );
  NAND2_X1 U7065 ( .A1(n9780), .A2(n7689), .ZN(n5757) );
  NAND2_X1 U7066 ( .A1(n5658), .A2(n5757), .ZN(n7618) );
  INV_X1 U7067 ( .A(n7619), .ZN(n5444) );
  NOR2_X1 U7068 ( .A1(n7618), .A2(n5444), .ZN(n5445) );
  NAND2_X1 U7069 ( .A1(n7620), .A2(n5445), .ZN(n7617) );
  NAND2_X1 U7070 ( .A1(n7617), .A2(n5757), .ZN(n7685) );
  XNOR2_X1 U7071 ( .A(n5446), .B(SI_13_), .ZN(n5447) );
  INV_X1 U7072 ( .A(n4366), .ZN(n5448) );
  NAND2_X1 U7073 ( .A1(n5449), .A2(n5448), .ZN(n5450) );
  NAND2_X1 U7074 ( .A1(n5450), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5451) );
  XNOR2_X1 U7075 ( .A(n5451), .B(P1_IR_REG_13__SCAN_IN), .ZN(n9644) );
  AOI22_X1 U7076 ( .A1(n5542), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n5541), .B2(
        n9644), .ZN(n5452) );
  NAND2_X1 U7077 ( .A1(n5545), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n5455) );
  NAND2_X1 U7078 ( .A1(n5427), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n5454) );
  AND2_X1 U7079 ( .A1(n5455), .A2(n5454), .ZN(n5461) );
  NAND2_X1 U7080 ( .A1(n5457), .A2(n5456), .ZN(n5458) );
  AND2_X1 U7081 ( .A1(n5473), .A2(n5458), .ZN(n8897) );
  NAND2_X1 U7082 ( .A1(n5549), .A2(n8897), .ZN(n5460) );
  NAND2_X1 U7083 ( .A1(n5556), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n5459) );
  NAND2_X1 U7084 ( .A1(n9788), .A2(n9775), .ZN(n5756) );
  AND2_X2 U7085 ( .A1(n7687), .A2(n5662), .ZN(n7705) );
  XNOR2_X1 U7086 ( .A(n5462), .B(n10058), .ZN(n5463) );
  XNOR2_X1 U7087 ( .A(n5464), .B(n5463), .ZN(n6640) );
  NAND2_X1 U7088 ( .A1(n6640), .A2(n5517), .ZN(n5468) );
  OR2_X1 U7089 ( .A1(n5465), .A2(n5124), .ZN(n5466) );
  XNOR2_X1 U7090 ( .A(n5466), .B(P1_IR_REG_14__SCAN_IN), .ZN(n9659) );
  AOI22_X1 U7091 ( .A1(n5542), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n5541), .B2(
        n9659), .ZN(n5467) );
  NAND2_X1 U7092 ( .A1(n5545), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n5470) );
  NAND2_X1 U7093 ( .A1(n5427), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5469) );
  AND2_X1 U7094 ( .A1(n5470), .A2(n5469), .ZN(n5477) );
  INV_X1 U7095 ( .A(n5471), .ZN(n5487) );
  NAND2_X1 U7096 ( .A1(n5473), .A2(n5472), .ZN(n5474) );
  AND2_X1 U7097 ( .A1(n5487), .A2(n5474), .ZN(n8792) );
  NAND2_X1 U7098 ( .A1(n5549), .A2(n8792), .ZN(n5476) );
  NAND2_X1 U7099 ( .A1(n5556), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n5475) );
  OR2_X1 U7100 ( .A1(n9427), .A2(n8939), .ZN(n5664) );
  NAND2_X1 U7101 ( .A1(n9427), .A2(n8939), .ZN(n5762) );
  XNOR2_X1 U7102 ( .A(n5478), .B(SI_15_), .ZN(n5479) );
  XNOR2_X1 U7103 ( .A(n5480), .B(n5479), .ZN(n6652) );
  NAND2_X1 U7104 ( .A1(n6652), .A2(n5517), .ZN(n5484) );
  NAND2_X1 U7105 ( .A1(n5481), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5482) );
  XNOR2_X1 U7106 ( .A(n5482), .B(P1_IR_REG_15__SCAN_IN), .ZN(n9684) );
  AOI22_X1 U7107 ( .A1(n5542), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n5541), .B2(
        n9684), .ZN(n5483) );
  AOI22_X1 U7108 ( .A1(n5556), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n5545), .B2(
        P1_REG1_REG_15__SCAN_IN), .ZN(n5490) );
  INV_X1 U7109 ( .A(n5485), .ZN(n5499) );
  INV_X1 U7110 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n5486) );
  NAND2_X1 U7111 ( .A1(n5487), .A2(n5486), .ZN(n5488) );
  AND2_X1 U7112 ( .A1(n5499), .A2(n5488), .ZN(n8938) );
  AOI22_X1 U7113 ( .A1(n5549), .A2(n8938), .B1(n5427), .B2(
        P1_REG0_REG_15__SCAN_IN), .ZN(n5489) );
  NAND2_X1 U7114 ( .A1(n7819), .A2(n9425), .ZN(n5651) );
  INV_X1 U7115 ( .A(n7721), .ZN(n5491) );
  XNOR2_X1 U7116 ( .A(n5492), .B(SI_16_), .ZN(n5493) );
  NAND2_X1 U7117 ( .A1(n5504), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5495) );
  XNOR2_X1 U7118 ( .A(n5495), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9052) );
  AOI22_X1 U7119 ( .A1(n5542), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n5541), .B2(
        n9052), .ZN(n5496) );
  NAND2_X2 U7120 ( .A1(n5497), .A2(n5496), .ZN(n8861) );
  AOI22_X1 U7121 ( .A1(n5556), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n5545), .B2(
        P1_REG1_REG_16__SCAN_IN), .ZN(n5502) );
  INV_X1 U7122 ( .A(n8870), .ZN(n8868) );
  INV_X1 U7123 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n5498) );
  NAND2_X1 U7124 ( .A1(n5499), .A2(n5498), .ZN(n5500) );
  AND2_X1 U7125 ( .A1(n8868), .A2(n5500), .ZN(n8858) );
  AOI22_X1 U7126 ( .A1(n5549), .A2(n8858), .B1(n5427), .B2(
        P1_REG0_REG_16__SCAN_IN), .ZN(n5501) );
  NAND2_X1 U7127 ( .A1(n5766), .A2(n5767), .ZN(n7833) );
  NAND2_X1 U7128 ( .A1(n6718), .A2(n5517), .ZN(n5507) );
  XNOR2_X1 U7129 ( .A(n5518), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9071) );
  AOI22_X1 U7130 ( .A1(n5542), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n5541), .B2(
        n9071), .ZN(n5506) );
  NAND2_X1 U7131 ( .A1(n5545), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n5509) );
  NAND2_X1 U7132 ( .A1(n5427), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n5508) );
  AND2_X1 U7133 ( .A1(n5509), .A2(n5508), .ZN(n5513) );
  INV_X1 U7134 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n9057) );
  NAND2_X1 U7135 ( .A1(n8868), .A2(n9057), .ZN(n5510) );
  AND2_X1 U7136 ( .A1(n5525), .A2(n5510), .ZN(n7821) );
  NAND2_X1 U7137 ( .A1(n5549), .A2(n7821), .ZN(n5512) );
  NAND2_X1 U7138 ( .A1(n5556), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n5511) );
  OR2_X1 U7139 ( .A1(n9096), .A2(n9414), .ZN(n5587) );
  NAND2_X1 U7140 ( .A1(n9096), .A2(n9414), .ZN(n5586) );
  NAND2_X1 U7141 ( .A1(n7828), .A2(n7827), .ZN(n5514) );
  NAND2_X1 U7142 ( .A1(n5514), .A2(n5586), .ZN(n9288) );
  XNOR2_X1 U7143 ( .A(n5516), .B(n5515), .ZN(n6733) );
  NAND2_X1 U7144 ( .A1(n6733), .A2(n5517), .ZN(n5521) );
  NAND2_X1 U7145 ( .A1(n5534), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5519) );
  XNOR2_X1 U7146 ( .A(n5519), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9708) );
  AOI22_X1 U7147 ( .A1(n5542), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n5541), .B2(
        n9708), .ZN(n5520) );
  NAND2_X1 U7148 ( .A1(n5545), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n5523) );
  NAND2_X1 U7149 ( .A1(n5427), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n5522) );
  AND2_X1 U7150 ( .A1(n5523), .A2(n5522), .ZN(n5529) );
  NAND2_X1 U7151 ( .A1(n5525), .A2(n5524), .ZN(n5526) );
  AND2_X1 U7152 ( .A1(n5548), .A2(n5526), .ZN(n9292) );
  NAND2_X1 U7153 ( .A1(n5549), .A2(n9292), .ZN(n5528) );
  NAND2_X1 U7154 ( .A1(n5556), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n5527) );
  OR2_X1 U7155 ( .A1(n9300), .A2(n9277), .ZN(n5680) );
  NAND2_X1 U7156 ( .A1(n9300), .A2(n9277), .ZN(n5678) );
  NAND2_X1 U7157 ( .A1(n9288), .A2(n9287), .ZN(n5530) );
  NAND2_X1 U7158 ( .A1(n5530), .A2(n5678), .ZN(n9276) );
  XNOR2_X1 U7159 ( .A(n5532), .B(n5531), .ZN(n7222) );
  NAND2_X1 U7160 ( .A1(n7222), .A2(n5517), .ZN(n5544) );
  NOR2_X1 U7161 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n5574) );
  NAND2_X1 U7162 ( .A1(n5533), .A2(n5574), .ZN(n5540) );
  NAND3_X1 U7163 ( .A1(n5534), .A2(P1_IR_REG_31__SCAN_IN), .A3(
        P1_IR_REG_19__SCAN_IN), .ZN(n5539) );
  INV_X1 U7164 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5537) );
  NAND2_X1 U7165 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), 
        .ZN(n5535) );
  NAND2_X1 U7166 ( .A1(n5535), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5536) );
  OAI21_X1 U7167 ( .B1(n5537), .B2(P1_IR_REG_31__SCAN_IN), .A(n5536), .ZN(
        n5538) );
  AOI22_X1 U7168 ( .A1(n5542), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n9080), .B2(
        n5541), .ZN(n5543) );
  NAND2_X1 U7169 ( .A1(n5545), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n5547) );
  NAND2_X1 U7170 ( .A1(n5427), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n5546) );
  AND2_X1 U7171 ( .A1(n5547), .A2(n5546), .ZN(n5552) );
  XNOR2_X1 U7172 ( .A(n5548), .B(P1_REG3_REG_19__SCAN_IN), .ZN(n9271) );
  NAND2_X1 U7173 ( .A1(n9271), .A2(n5549), .ZN(n5551) );
  NAND2_X1 U7174 ( .A1(n5556), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n5550) );
  NAND2_X1 U7175 ( .A1(n9392), .A2(n9256), .ZN(n5681) );
  NAND2_X1 U7176 ( .A1(n9280), .A2(n5687), .ZN(n9252) );
  NAND2_X1 U7177 ( .A1(n9164), .A2(n9324), .ZN(n5777) );
  OAI21_X1 U7178 ( .B1(n5779), .B2(n9252), .A(n5777), .ZN(n5553) );
  AND2_X1 U7179 ( .A1(n5553), .A2(n5780), .ZN(n5554) );
  NOR2_X1 U7180 ( .A1(n5783), .A2(n5554), .ZN(n5555) );
  NOR2_X1 U7181 ( .A1(n5785), .A2(n5555), .ZN(n5560) );
  INV_X1 U7182 ( .A(n9439), .ZN(n5721) );
  INV_X1 U7183 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n9311) );
  NAND2_X1 U7184 ( .A1(n5556), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n5558) );
  NAND2_X1 U7185 ( .A1(n5427), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n5557) );
  OAI211_X1 U7186 ( .C1(n9311), .C2(n5559), .A(n5558), .B(n5557), .ZN(n8950)
         );
  INV_X1 U7187 ( .A(n8950), .ZN(n9121) );
  NAND2_X1 U7188 ( .A1(n5721), .A2(n9121), .ZN(n5609) );
  NAND2_X1 U7189 ( .A1(n9316), .A2(n8951), .ZN(n5717) );
  NAND2_X1 U7190 ( .A1(n5609), .A2(n5717), .ZN(n5786) );
  INV_X1 U7191 ( .A(n9088), .ZN(n5571) );
  OAI22_X1 U7192 ( .A1(n5560), .A2(n5786), .B1(n5571), .B2(n5583), .ZN(n5561)
         );
  OAI21_X1 U7193 ( .B1(n9439), .B2(n9088), .A(n5561), .ZN(n5572) );
  INV_X1 U7194 ( .A(SI_31_), .ZN(n5565) );
  XNOR2_X1 U7195 ( .A(n5566), .B(n5565), .ZN(n5567) );
  NAND2_X1 U7196 ( .A1(n8763), .A2(n5517), .ZN(n5570) );
  INV_X1 U7197 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n9473) );
  OR2_X1 U7198 ( .A1(n5297), .A2(n9473), .ZN(n5569) );
  NAND2_X1 U7199 ( .A1(n9084), .A2(n5571), .ZN(n5801) );
  AND2_X1 U7200 ( .A1(n9435), .A2(n9088), .ZN(n5790) );
  AOI21_X1 U7201 ( .B1(n5572), .B2(n5801), .A(n5790), .ZN(n5611) );
  NAND2_X1 U7202 ( .A1(n5574), .A2(n5573), .ZN(n5575) );
  NAND2_X1 U7203 ( .A1(n5792), .A2(n5576), .ZN(n5795) );
  INV_X1 U7204 ( .A(n5795), .ZN(n5578) );
  INV_X1 U7205 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5577) );
  NAND2_X1 U7206 ( .A1(n5578), .A2(n5577), .ZN(n5812) );
  INV_X1 U7207 ( .A(n5580), .ZN(n5579) );
  NAND2_X1 U7208 ( .A1(n5579), .A2(P1_IR_REG_22__SCAN_IN), .ZN(n5581) );
  NAND2_X1 U7209 ( .A1(n5801), .A2(n5583), .ZN(n5789) );
  XNOR2_X1 U7210 ( .A(n9388), .B(n9278), .ZN(n9253) );
  AND2_X1 U7211 ( .A1(n5678), .A2(n5586), .ZN(n5682) );
  AND2_X1 U7212 ( .A1(n5680), .A2(n5587), .ZN(n5772) );
  INV_X1 U7213 ( .A(n6942), .ZN(n9721) );
  XNOR2_X1 U7214 ( .A(n8822), .B(n9721), .ZN(n9718) );
  NAND4_X1 U7215 ( .A1(n6738), .A2(n6748), .A3(n9718), .A4(n7446), .ZN(n5589)
         );
  NAND2_X1 U7216 ( .A1(n6702), .A2(n6934), .ZN(n5588) );
  NOR2_X1 U7217 ( .A1(n5589), .A2(n5588), .ZN(n5591) );
  INV_X1 U7218 ( .A(n5638), .ZN(n5590) );
  NAND4_X1 U7219 ( .A1(n5591), .A2(n5590), .A3(n6791), .A4(n6766), .ZN(n5593)
         );
  NOR2_X1 U7220 ( .A1(n5593), .A2(n5592), .ZN(n5594) );
  NAND4_X1 U7221 ( .A1(n5596), .A2(n5595), .A3(n7514), .A4(n5594), .ZN(n5597)
         );
  NOR2_X1 U7222 ( .A1(n7618), .A2(n5597), .ZN(n5598) );
  NAND4_X1 U7223 ( .A1(n7721), .A2(n7719), .A3(n5599), .A4(n5598), .ZN(n5600)
         );
  NOR2_X1 U7224 ( .A1(n7833), .A2(n5600), .ZN(n5601) );
  NAND4_X1 U7225 ( .A1(n5602), .A2(n5682), .A3(n5772), .A4(n5601), .ZN(n5603)
         );
  NOR2_X1 U7226 ( .A1(n9253), .A2(n5603), .ZN(n5604) );
  XNOR2_X1 U7227 ( .A(n9233), .B(n9378), .ZN(n9224) );
  XNOR2_X1 U7228 ( .A(n9241), .B(n9368), .ZN(n9239) );
  NAND4_X1 U7229 ( .A1(n9211), .A2(n5604), .A3(n9224), .A4(n9239), .ZN(n5605)
         );
  NOR2_X1 U7230 ( .A1(n9190), .A2(n5605), .ZN(n5606) );
  NAND2_X1 U7231 ( .A1(n9175), .A2(n5606), .ZN(n5607) );
  NAND2_X1 U7232 ( .A1(n5716), .A2(n5717), .ZN(n9120) );
  INV_X1 U7233 ( .A(n9120), .ZN(n9109) );
  NAND4_X1 U7234 ( .A1(n4983), .A2(n5609), .A3(n9109), .A4(n5608), .ZN(n5610)
         );
  OR3_X1 U7235 ( .A1(n5790), .A2(n5789), .A3(n5610), .ZN(n5729) );
  OAI21_X1 U7236 ( .B1(n5611), .B2(n6699), .A(n5729), .ZN(n5732) );
  NAND2_X1 U7237 ( .A1(n5834), .A2(n9080), .ZN(n6840) );
  MUX2_X1 U7238 ( .A(n5613), .B(n5612), .S(n6840), .Z(n5699) );
  NAND3_X1 U7239 ( .A1(n5614), .A2(n9113), .A3(n6840), .ZN(n5615) );
  NAND2_X1 U7240 ( .A1(n9224), .A2(n5615), .ZN(n5695) );
  INV_X1 U7241 ( .A(n5617), .ZN(n5618) );
  OR2_X1 U7242 ( .A1(n6749), .A2(n5618), .ZN(n5737) );
  AND2_X1 U7243 ( .A1(n5626), .A2(n5619), .ZN(n5735) );
  NAND2_X1 U7244 ( .A1(n5737), .A2(n5735), .ZN(n5620) );
  NAND2_X1 U7245 ( .A1(n7264), .A2(n5743), .ZN(n5630) );
  OAI21_X1 U7246 ( .B1(n5624), .B2(n5630), .A(n5746), .ZN(n5635) );
  INV_X1 U7247 ( .A(n5625), .ZN(n5629) );
  NAND2_X1 U7248 ( .A1(n5738), .A2(n5626), .ZN(n5628) );
  AND2_X1 U7249 ( .A1(n5627), .A2(n6767), .ZN(n5742) );
  OAI21_X1 U7250 ( .B1(n5629), .B2(n5628), .A(n5742), .ZN(n5633) );
  INV_X1 U7251 ( .A(n5630), .ZN(n5632) );
  AOI21_X1 U7252 ( .B1(n5633), .B2(n5632), .A(n5631), .ZN(n5634) );
  NAND2_X1 U7253 ( .A1(n7307), .A2(n5636), .ZN(n7305) );
  NAND2_X1 U7254 ( .A1(n7432), .A2(n5636), .ZN(n5637) );
  MUX2_X1 U7255 ( .A(n5638), .B(n5637), .S(n4365), .Z(n5639) );
  INV_X1 U7256 ( .A(n5639), .ZN(n5640) );
  NAND2_X1 U7257 ( .A1(n7429), .A2(n7431), .ZN(n5642) );
  MUX2_X1 U7258 ( .A(n5643), .B(n5642), .S(n4365), .Z(n5644) );
  INV_X1 U7259 ( .A(n5644), .ZN(n5645) );
  NAND2_X1 U7260 ( .A1(n5646), .A2(n5645), .ZN(n5655) );
  NAND2_X1 U7261 ( .A1(n5655), .A2(n7430), .ZN(n5647) );
  NAND2_X1 U7262 ( .A1(n5647), .A2(n7516), .ZN(n5650) );
  AND2_X1 U7263 ( .A1(n7619), .A2(n5749), .ZN(n5649) );
  NAND2_X1 U7264 ( .A1(n5757), .A2(n5656), .ZN(n5648) );
  AND3_X1 U7265 ( .A1(n5762), .A2(n4365), .A3(n5756), .ZN(n5652) );
  OAI211_X1 U7266 ( .C1(n5654), .C2(n5653), .A(n5770), .B(n5652), .ZN(n5676)
         );
  NAND2_X1 U7267 ( .A1(n5655), .A2(n7429), .ZN(n5657) );
  NAND2_X1 U7268 ( .A1(n5656), .A2(n7516), .ZN(n5752) );
  AOI21_X1 U7269 ( .B1(n5657), .B2(n5749), .A(n5752), .ZN(n5659) );
  NAND2_X1 U7270 ( .A1(n5658), .A2(n7619), .ZN(n5753) );
  OAI21_X1 U7271 ( .B1(n5659), .B2(n5753), .A(n5757), .ZN(n5661) );
  AND4_X1 U7272 ( .A1(n5765), .A2(n5664), .A3(n5662), .A4(n6840), .ZN(n5660)
         );
  NAND3_X1 U7273 ( .A1(n5661), .A2(n5660), .A3(n5766), .ZN(n5675) );
  NAND2_X1 U7274 ( .A1(n5664), .A2(n5662), .ZN(n5761) );
  NAND3_X1 U7275 ( .A1(n5761), .A2(n4365), .A3(n5762), .ZN(n5670) );
  NAND2_X1 U7276 ( .A1(n5762), .A2(n5756), .ZN(n5663) );
  NAND4_X1 U7277 ( .A1(n5765), .A2(n5664), .A3(n6840), .A4(n5663), .ZN(n5665)
         );
  NAND2_X1 U7278 ( .A1(n5766), .A2(n5665), .ZN(n5666) );
  OAI21_X1 U7279 ( .B1(n5766), .B2(n4365), .A(n5666), .ZN(n5669) );
  INV_X1 U7280 ( .A(n5765), .ZN(n5667) );
  NAND3_X1 U7281 ( .A1(n5767), .A2(n5667), .A3(n4365), .ZN(n5668) );
  OAI211_X1 U7282 ( .C1(n5672), .C2(n5670), .A(n5669), .B(n5668), .ZN(n5671)
         );
  INV_X1 U7283 ( .A(n5671), .ZN(n5674) );
  NAND2_X1 U7284 ( .A1(n5683), .A2(n5772), .ZN(n5679) );
  NAND3_X1 U7285 ( .A1(n5679), .A2(n5681), .A3(n5678), .ZN(n5686) );
  NAND2_X1 U7286 ( .A1(n5687), .A2(n5680), .ZN(n5774) );
  OAI21_X1 U7287 ( .B1(n5774), .B2(n5682), .A(n5681), .ZN(n5776) );
  NOR2_X1 U7288 ( .A1(n5776), .A2(n5684), .ZN(n5685) );
  NAND2_X1 U7289 ( .A1(n5688), .A2(n5687), .ZN(n9111) );
  NAND2_X1 U7290 ( .A1(n9111), .A2(n4365), .ZN(n5689) );
  NAND2_X1 U7291 ( .A1(n5691), .A2(n4365), .ZN(n5693) );
  MUX2_X1 U7292 ( .A(n5696), .B(n9192), .S(n4365), .Z(n5697) );
  OAI211_X1 U7293 ( .C1(n5699), .C2(n5698), .A(n9194), .B(n5697), .ZN(n5702)
         );
  MUX2_X1 U7294 ( .A(n9176), .B(n5700), .S(n6840), .Z(n5701) );
  INV_X1 U7295 ( .A(n5777), .ZN(n9117) );
  NAND2_X1 U7296 ( .A1(n5711), .A2(n5780), .ZN(n5708) );
  INV_X1 U7297 ( .A(n5712), .ZN(n5707) );
  AOI21_X1 U7298 ( .B1(n5708), .B2(n5709), .A(n5707), .ZN(n5715) );
  NAND2_X1 U7299 ( .A1(n5713), .A2(n5712), .ZN(n5714) );
  MUX2_X1 U7300 ( .A(n5717), .B(n5716), .S(n6840), .Z(n5718) );
  OAI21_X1 U7301 ( .B1(n5719), .B2(n9120), .A(n5718), .ZN(n5723) );
  MUX2_X1 U7302 ( .A(n5723), .B(n6840), .S(n9439), .Z(n5720) );
  MUX2_X1 U7303 ( .A(n5723), .B(n4365), .S(n5721), .Z(n5726) );
  NAND2_X1 U7304 ( .A1(n9084), .A2(n9121), .ZN(n5724) );
  NAND2_X1 U7305 ( .A1(n5724), .A2(n9088), .ZN(n5725) );
  INV_X1 U7306 ( .A(n5729), .ZN(n5730) );
  NAND2_X1 U7307 ( .A1(n9719), .A2(n6959), .ZN(n5734) );
  NAND2_X1 U7308 ( .A1(n8822), .A2(n6942), .ZN(n5733) );
  AND3_X1 U7309 ( .A1(n5734), .A2(n5733), .A3(n5831), .ZN(n5736) );
  OAI21_X1 U7310 ( .B1(n5737), .B2(n5736), .A(n5735), .ZN(n5741) );
  INV_X1 U7311 ( .A(n5738), .ZN(n5739) );
  AOI21_X1 U7312 ( .B1(n5741), .B2(n5740), .A(n5739), .ZN(n5745) );
  INV_X1 U7313 ( .A(n5742), .ZN(n5744) );
  OAI21_X1 U7314 ( .B1(n5745), .B2(n5744), .A(n5743), .ZN(n5748) );
  NAND3_X1 U7315 ( .A1(n5748), .A2(n5747), .A3(n5746), .ZN(n5751) );
  NAND3_X1 U7316 ( .A1(n5751), .A2(n5750), .A3(n5749), .ZN(n5755) );
  INV_X1 U7317 ( .A(n5752), .ZN(n5754) );
  AOI21_X1 U7318 ( .B1(n5755), .B2(n5754), .A(n5753), .ZN(n5760) );
  INV_X1 U7319 ( .A(n5756), .ZN(n5759) );
  INV_X1 U7320 ( .A(n5757), .ZN(n5758) );
  OR3_X1 U7321 ( .A1(n5760), .A2(n5759), .A3(n5758), .ZN(n5764) );
  INV_X1 U7322 ( .A(n5761), .ZN(n5763) );
  AOI21_X1 U7323 ( .B1(n5764), .B2(n5763), .A(n4787), .ZN(n5769) );
  NAND2_X1 U7324 ( .A1(n5766), .A2(n5765), .ZN(n5768) );
  AOI22_X1 U7325 ( .A1(n5770), .A2(n5769), .B1(n5768), .B2(n5767), .ZN(n5771)
         );
  NAND2_X1 U7326 ( .A1(n5772), .A2(n5771), .ZN(n5773) );
  NOR2_X1 U7327 ( .A1(n5774), .A2(n5773), .ZN(n5775) );
  NOR2_X1 U7328 ( .A1(n5776), .A2(n5775), .ZN(n5778) );
  OAI21_X1 U7329 ( .B1(n5779), .B2(n5778), .A(n5777), .ZN(n5781) );
  AND2_X1 U7330 ( .A1(n5781), .A2(n5780), .ZN(n5782) );
  NOR2_X1 U7331 ( .A1(n5783), .A2(n5782), .ZN(n5784) );
  NOR2_X1 U7332 ( .A1(n5785), .A2(n5784), .ZN(n5787) );
  NOR2_X1 U7333 ( .A1(n5787), .A2(n5786), .ZN(n5788) );
  OR2_X1 U7334 ( .A1(n5789), .A2(n5788), .ZN(n5791) );
  INV_X1 U7335 ( .A(n5790), .ZN(n5806) );
  NAND2_X1 U7336 ( .A1(n5791), .A2(n5806), .ZN(n5799) );
  NAND2_X1 U7337 ( .A1(n5799), .A2(n9080), .ZN(n5796) );
  MUX2_X1 U7338 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5793), .S(
        P1_IR_REG_20__SCAN_IN), .Z(n5794) );
  NAND2_X1 U7339 ( .A1(n5797), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5798) );
  AND2_X1 U7340 ( .A1(n6621), .A2(P1_STATE_REG_SCAN_IN), .ZN(n5802) );
  OAI21_X1 U7341 ( .B1(n5799), .B2(n6698), .A(n5802), .ZN(n5828) );
  OAI21_X1 U7342 ( .B1(n5801), .B2(n7863), .A(n5800), .ZN(n5805) );
  INV_X1 U7343 ( .A(n5802), .ZN(n7638) );
  NAND3_X1 U7344 ( .A1(n5834), .A2(n5831), .A3(n6839), .ZN(n5803) );
  NOR2_X1 U7345 ( .A1(n7638), .A2(n5803), .ZN(n5804) );
  OAI211_X1 U7346 ( .C1(n5806), .C2(n7863), .A(n5805), .B(n5804), .ZN(n5826)
         );
  INV_X1 U7347 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n5807) );
  NAND2_X1 U7348 ( .A1(n5808), .A2(n5807), .ZN(n5811) );
  INV_X1 U7349 ( .A(n5813), .ZN(n5818) );
  NAND2_X1 U7350 ( .A1(n4385), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5817) );
  NAND2_X1 U7351 ( .A1(n5818), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5819) );
  XNOR2_X1 U7352 ( .A(n5819), .B(P1_IR_REG_25__SCAN_IN), .ZN(n6073) );
  INV_X1 U7353 ( .A(n9542), .ZN(n9564) );
  NOR4_X1 U7354 ( .A1(n6686), .A2(n9776), .A3(n9485), .A4(n6698), .ZN(n5824)
         );
  OAI21_X1 U7355 ( .B1(n7638), .B2(n5829), .A(P1_B_REG_SCAN_IN), .ZN(n5823) );
  OR2_X1 U7356 ( .A1(n5824), .A2(n5823), .ZN(n5825) );
  NAND2_X1 U7357 ( .A1(n5829), .A2(n7863), .ZN(n6695) );
  AND2_X1 U7358 ( .A1(n6695), .A2(n5833), .ZN(n5832) );
  NAND2_X1 U7359 ( .A1(n5832), .A2(n5837), .ZN(n5848) );
  INV_X1 U7360 ( .A(n5833), .ZN(n5836) );
  NAND3_X4 U7361 ( .A1(n5837), .A2(n7243), .A3(n5835), .ZN(n6058) );
  NAND2_X1 U7362 ( .A1(n5862), .A2(n8823), .ZN(n5839) );
  AND2_X2 U7363 ( .A1(n5837), .A2(n5836), .ZN(n5871) );
  NAND2_X1 U7364 ( .A1(n9719), .A2(n5871), .ZN(n5838) );
  NAND2_X1 U7365 ( .A1(n5839), .A2(n5838), .ZN(n5840) );
  AND2_X1 U7366 ( .A1(n8823), .A2(n5871), .ZN(n5841) );
  AOI21_X1 U7367 ( .B1(n9719), .B2(n6011), .A(n5841), .ZN(n5851) );
  XNOR2_X1 U7368 ( .A(n5850), .B(n5851), .ZN(n8820) );
  NAND2_X1 U7369 ( .A1(n9721), .A2(n5862), .ZN(n5843) );
  NAND2_X1 U7370 ( .A1(n8822), .A2(n5871), .ZN(n5842) );
  INV_X1 U7371 ( .A(n5837), .ZN(n6582) );
  NAND2_X1 U7372 ( .A1(n6582), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5844) );
  NAND2_X1 U7373 ( .A1(n5849), .A2(n5844), .ZN(n6657) );
  NAND2_X1 U7374 ( .A1(n8822), .A2(n6011), .ZN(n5847) );
  OAI22_X1 U7375 ( .A1(n6942), .A2(n5892), .B1(n9544), .B2(n5837), .ZN(n5845)
         );
  INV_X1 U7376 ( .A(n5845), .ZN(n5846) );
  NAND2_X1 U7377 ( .A1(n5847), .A2(n5846), .ZN(n6656) );
  AOI22_X1 U7378 ( .A1(n6657), .A2(n6656), .B1(n5849), .B2(n6055), .ZN(n8819)
         );
  NAND2_X1 U7379 ( .A1(n8820), .A2(n8819), .ZN(n8818) );
  INV_X1 U7380 ( .A(n5850), .ZN(n5852) );
  NAND2_X1 U7381 ( .A1(n5852), .A2(n5851), .ZN(n5853) );
  NAND2_X1 U7382 ( .A1(n8818), .A2(n5853), .ZN(n6675) );
  NAND2_X1 U7383 ( .A1(n8962), .A2(n5871), .ZN(n5855) );
  NAND2_X1 U7384 ( .A1(n6757), .A2(n5862), .ZN(n5854) );
  NAND2_X1 U7385 ( .A1(n5855), .A2(n5854), .ZN(n5856) );
  XNOR2_X1 U7386 ( .A(n5856), .B(n4371), .ZN(n5857) );
  AOI22_X1 U7387 ( .A1(n8962), .A2(n6011), .B1(n6757), .B2(n6049), .ZN(n5858)
         );
  XNOR2_X1 U7388 ( .A(n5857), .B(n5858), .ZN(n6676) );
  NAND2_X1 U7389 ( .A1(n6675), .A2(n6676), .ZN(n5861) );
  INV_X1 U7390 ( .A(n5857), .ZN(n5859) );
  NAND2_X1 U7391 ( .A1(n5859), .A2(n5858), .ZN(n5860) );
  NAND2_X1 U7392 ( .A1(n5861), .A2(n5860), .ZN(n6661) );
  NAND2_X1 U7393 ( .A1(n8961), .A2(n6049), .ZN(n5864) );
  INV_X1 U7394 ( .A(n6954), .ZN(n6744) );
  NAND2_X1 U7395 ( .A1(n6744), .A2(n5862), .ZN(n5863) );
  NAND2_X1 U7396 ( .A1(n5864), .A2(n5863), .ZN(n5865) );
  XNOR2_X1 U7397 ( .A(n5865), .B(n4371), .ZN(n5866) );
  AOI22_X1 U7398 ( .A1(n8961), .A2(n6011), .B1(n6744), .B2(n6049), .ZN(n5867)
         );
  XNOR2_X1 U7399 ( .A(n5866), .B(n5867), .ZN(n6662) );
  NAND2_X1 U7400 ( .A1(n6661), .A2(n6662), .ZN(n5870) );
  INV_X1 U7401 ( .A(n5866), .ZN(n5868) );
  NAND2_X1 U7402 ( .A1(n5868), .A2(n5867), .ZN(n5869) );
  NAND2_X1 U7403 ( .A1(n5870), .A2(n5869), .ZN(n6722) );
  INV_X1 U7404 ( .A(n6722), .ZN(n5876) );
  OAI22_X1 U7405 ( .A1(n6833), .A2(n5892), .B1(n6867), .B2(n5880), .ZN(n5872)
         );
  XNOR2_X1 U7406 ( .A(n5872), .B(n4371), .ZN(n5878) );
  OR2_X1 U7407 ( .A1(n6833), .A2(n6058), .ZN(n5874) );
  NAND2_X1 U7408 ( .A1(n6727), .A2(n6049), .ZN(n5873) );
  NAND2_X1 U7409 ( .A1(n5874), .A2(n5873), .ZN(n5877) );
  XNOR2_X1 U7410 ( .A(n5878), .B(n5877), .ZN(n6725) );
  INV_X1 U7411 ( .A(n6725), .ZN(n5875) );
  NAND2_X1 U7412 ( .A1(n5876), .A2(n5875), .ZN(n6723) );
  NAND2_X1 U7413 ( .A1(n5878), .A2(n5877), .ZN(n5879) );
  NAND2_X1 U7414 ( .A1(n6723), .A2(n5879), .ZN(n5884) );
  NAND2_X1 U7415 ( .A1(n8959), .A2(n5871), .ZN(n5882) );
  NAND2_X1 U7416 ( .A1(n6835), .A2(n6052), .ZN(n5881) );
  NAND2_X1 U7417 ( .A1(n5882), .A2(n5881), .ZN(n5883) );
  XNOR2_X1 U7418 ( .A(n5883), .B(n4371), .ZN(n5885) );
  NAND2_X1 U7419 ( .A1(n5884), .A2(n5885), .ZN(n6828) );
  AOI22_X1 U7420 ( .A1(n8959), .A2(n6011), .B1(n6835), .B2(n6049), .ZN(n6830)
         );
  NAND2_X1 U7421 ( .A1(n6828), .A2(n6830), .ZN(n5888) );
  INV_X1 U7422 ( .A(n5885), .ZN(n5886) );
  NAND2_X1 U7423 ( .A1(n8958), .A2(n6049), .ZN(n5890) );
  NAND2_X1 U7424 ( .A1(n7037), .A2(n6052), .ZN(n5889) );
  NAND2_X1 U7425 ( .A1(n5890), .A2(n5889), .ZN(n5891) );
  XNOR2_X1 U7426 ( .A(n5891), .B(n6055), .ZN(n5895) );
  NAND2_X1 U7427 ( .A1(n8958), .A2(n6011), .ZN(n5894) );
  NAND2_X1 U7428 ( .A1(n7037), .A2(n6049), .ZN(n5893) );
  AND2_X1 U7429 ( .A1(n5894), .A2(n5893), .ZN(n5896) );
  AND2_X1 U7430 ( .A1(n5895), .A2(n5896), .ZN(n7031) );
  INV_X1 U7431 ( .A(n5895), .ZN(n5898) );
  INV_X1 U7432 ( .A(n5896), .ZN(n5897) );
  NAND2_X1 U7433 ( .A1(n5898), .A2(n5897), .ZN(n7032) );
  OAI22_X1 U7434 ( .A1(n7311), .A2(n6058), .B1(n7425), .B2(n5892), .ZN(n7253)
         );
  OAI22_X1 U7435 ( .A1(n7311), .A2(n5892), .B1(n7425), .B2(n5880), .ZN(n5899)
         );
  XNOR2_X1 U7436 ( .A(n5899), .B(n4371), .ZN(n7252) );
  NAND2_X1 U7437 ( .A1(n7437), .A2(n6052), .ZN(n5900) );
  OAI21_X1 U7438 ( .B1(n7439), .B2(n5892), .A(n5900), .ZN(n5901) );
  XNOR2_X1 U7439 ( .A(n5901), .B(n4371), .ZN(n5904) );
  INV_X1 U7440 ( .A(n5904), .ZN(n5902) );
  NAND2_X1 U7441 ( .A1(n5903), .A2(n5902), .ZN(n5906) );
  AOI22_X1 U7442 ( .A1(n9746), .A2(n6011), .B1(n6049), .B2(n7437), .ZN(n7548)
         );
  NAND2_X1 U7443 ( .A1(n9747), .A2(n6052), .ZN(n5908) );
  NAND2_X1 U7444 ( .A1(n9755), .A2(n6049), .ZN(n5907) );
  NAND2_X1 U7445 ( .A1(n5908), .A2(n5907), .ZN(n5909) );
  XNOR2_X1 U7446 ( .A(n5909), .B(n6055), .ZN(n5914) );
  NAND2_X1 U7447 ( .A1(n9747), .A2(n6049), .ZN(n5911) );
  NAND2_X1 U7448 ( .A1(n9755), .A2(n6011), .ZN(n5910) );
  NAND2_X1 U7449 ( .A1(n5911), .A2(n5910), .ZN(n5912) );
  XNOR2_X1 U7450 ( .A(n5914), .B(n5912), .ZN(n7643) );
  INV_X1 U7451 ( .A(n5912), .ZN(n5913) );
  NAND2_X1 U7452 ( .A1(n5914), .A2(n5913), .ZN(n5915) );
  NAND2_X1 U7453 ( .A1(n7642), .A2(n5915), .ZN(n5920) );
  NAND2_X1 U7454 ( .A1(n7513), .A2(n6052), .ZN(n5917) );
  OR2_X1 U7455 ( .A1(n7814), .A2(n5892), .ZN(n5916) );
  NAND2_X1 U7456 ( .A1(n5917), .A2(n5916), .ZN(n5918) );
  XNOR2_X1 U7457 ( .A(n5918), .B(n6055), .ZN(n5919) );
  NAND2_X1 U7458 ( .A1(n5920), .A2(n5919), .ZN(n5922) );
  NOR2_X1 U7459 ( .A1(n7814), .A2(n6058), .ZN(n5921) );
  AOI21_X1 U7460 ( .B1(n7513), .B2(n6049), .A(n5921), .ZN(n7761) );
  NAND2_X1 U7461 ( .A1(n7816), .A2(n6052), .ZN(n5924) );
  OR2_X1 U7462 ( .A1(n9777), .A2(n5892), .ZN(n5923) );
  NAND2_X1 U7463 ( .A1(n5924), .A2(n5923), .ZN(n5925) );
  XNOR2_X1 U7464 ( .A(n5925), .B(n6055), .ZN(n5928) );
  NOR2_X1 U7465 ( .A1(n9777), .A2(n6058), .ZN(n5926) );
  AOI21_X1 U7466 ( .B1(n7816), .B2(n6049), .A(n5926), .ZN(n5927) );
  OR2_X1 U7467 ( .A1(n5928), .A2(n5927), .ZN(n7809) );
  NAND2_X1 U7468 ( .A1(n7811), .A2(n7809), .ZN(n5929) );
  NAND2_X1 U7469 ( .A1(n5928), .A2(n5927), .ZN(n7808) );
  NAND2_X1 U7470 ( .A1(n5929), .A2(n7808), .ZN(n8837) );
  NAND2_X1 U7471 ( .A1(n9780), .A2(n6052), .ZN(n5931) );
  OR2_X1 U7472 ( .A1(n7689), .A2(n5892), .ZN(n5930) );
  NAND2_X1 U7473 ( .A1(n5931), .A2(n5930), .ZN(n5932) );
  XNOR2_X1 U7474 ( .A(n5932), .B(n4371), .ZN(n5934) );
  NOR2_X1 U7475 ( .A1(n7689), .A2(n6058), .ZN(n5933) );
  AOI21_X1 U7476 ( .B1(n9780), .B2(n6049), .A(n5933), .ZN(n5935) );
  XNOR2_X1 U7477 ( .A(n5934), .B(n5935), .ZN(n8836) );
  NAND2_X1 U7478 ( .A1(n8837), .A2(n8836), .ZN(n5938) );
  INV_X1 U7479 ( .A(n5934), .ZN(n5936) );
  NAND2_X1 U7480 ( .A1(n5936), .A2(n5935), .ZN(n5937) );
  NAND2_X1 U7481 ( .A1(n5938), .A2(n5937), .ZN(n8896) );
  NAND2_X1 U7482 ( .A1(n9788), .A2(n6052), .ZN(n5940) );
  INV_X1 U7483 ( .A(n9775), .ZN(n8954) );
  NAND2_X1 U7484 ( .A1(n8954), .A2(n5871), .ZN(n5939) );
  NAND2_X1 U7485 ( .A1(n5940), .A2(n5939), .ZN(n5941) );
  XNOR2_X1 U7486 ( .A(n5941), .B(n4371), .ZN(n5943) );
  NOR2_X1 U7487 ( .A1(n9775), .A2(n6058), .ZN(n5942) );
  AOI21_X1 U7488 ( .B1(n9788), .B2(n6049), .A(n5942), .ZN(n5944) );
  XNOR2_X1 U7489 ( .A(n5943), .B(n5944), .ZN(n8895) );
  NAND2_X1 U7490 ( .A1(n8896), .A2(n8895), .ZN(n5947) );
  INV_X1 U7491 ( .A(n5943), .ZN(n5945) );
  NAND2_X1 U7492 ( .A1(n5945), .A2(n5944), .ZN(n5946) );
  NAND2_X1 U7493 ( .A1(n5947), .A2(n5946), .ZN(n8791) );
  NAND2_X1 U7494 ( .A1(n9427), .A2(n6052), .ZN(n5949) );
  INV_X1 U7495 ( .A(n8939), .ZN(n8953) );
  NAND2_X1 U7496 ( .A1(n8953), .A2(n5871), .ZN(n5948) );
  NAND2_X1 U7497 ( .A1(n5949), .A2(n5948), .ZN(n5950) );
  XNOR2_X1 U7498 ( .A(n5950), .B(n6055), .ZN(n8789) );
  NOR2_X1 U7499 ( .A1(n8939), .A2(n6058), .ZN(n5951) );
  AOI21_X1 U7500 ( .B1(n9427), .B2(n6049), .A(n5951), .ZN(n8788) );
  AND2_X1 U7501 ( .A1(n8789), .A2(n8788), .ZN(n5952) );
  INV_X1 U7502 ( .A(n8789), .ZN(n5954) );
  INV_X1 U7503 ( .A(n8788), .ZN(n5953) );
  NAND2_X1 U7504 ( .A1(n5954), .A2(n5953), .ZN(n5955) );
  NAND2_X1 U7505 ( .A1(n8861), .A2(n6052), .ZN(n5958) );
  OR2_X1 U7506 ( .A1(n7824), .A2(n5892), .ZN(n5957) );
  NAND2_X1 U7507 ( .A1(n5958), .A2(n5957), .ZN(n5959) );
  XNOR2_X1 U7508 ( .A(n5959), .B(n6055), .ZN(n8855) );
  NOR2_X1 U7509 ( .A1(n7824), .A2(n6058), .ZN(n5960) );
  AOI21_X1 U7510 ( .B1(n8861), .B2(n6049), .A(n5960), .ZN(n8854) );
  NAND2_X1 U7511 ( .A1(n7819), .A2(n6052), .ZN(n5962) );
  OR2_X1 U7512 ( .A1(n9425), .A2(n5892), .ZN(n5961) );
  NAND2_X1 U7513 ( .A1(n5962), .A2(n5961), .ZN(n5963) );
  XNOR2_X1 U7514 ( .A(n5963), .B(n6055), .ZN(n8852) );
  NOR2_X1 U7515 ( .A1(n9425), .A2(n6058), .ZN(n5964) );
  AOI21_X1 U7516 ( .B1(n7819), .B2(n6049), .A(n5964), .ZN(n8935) );
  OAI22_X1 U7517 ( .A1(n8855), .A2(n8854), .B1(n8852), .B2(n8935), .ZN(n5970)
         );
  NAND2_X1 U7518 ( .A1(n8852), .A2(n8935), .ZN(n5966) );
  INV_X1 U7519 ( .A(n8854), .ZN(n5965) );
  NAND2_X1 U7520 ( .A1(n5966), .A2(n5965), .ZN(n5968) );
  INV_X1 U7521 ( .A(n5966), .ZN(n5967) );
  AOI22_X1 U7522 ( .A1(n8855), .A2(n5968), .B1(n8854), .B2(n5967), .ZN(n5969)
         );
  NAND2_X1 U7523 ( .A1(n9096), .A2(n6052), .ZN(n5972) );
  INV_X1 U7524 ( .A(n9414), .ZN(n9397) );
  NAND2_X1 U7525 ( .A1(n9397), .A2(n5871), .ZN(n5971) );
  NAND2_X1 U7526 ( .A1(n5972), .A2(n5971), .ZN(n5973) );
  XNOR2_X1 U7527 ( .A(n5973), .B(n6055), .ZN(n8865) );
  NOR2_X1 U7528 ( .A1(n9414), .A2(n6058), .ZN(n5974) );
  AOI21_X1 U7529 ( .B1(n9096), .B2(n6049), .A(n5974), .ZN(n8864) );
  AND2_X1 U7530 ( .A1(n8865), .A2(n8864), .ZN(n5975) );
  NAND2_X1 U7531 ( .A1(n9300), .A2(n6052), .ZN(n5977) );
  NAND2_X1 U7532 ( .A1(n9405), .A2(n5871), .ZN(n5976) );
  NAND2_X1 U7533 ( .A1(n5977), .A2(n5976), .ZN(n5978) );
  XNOR2_X1 U7534 ( .A(n5978), .B(n6055), .ZN(n8808) );
  NOR2_X1 U7535 ( .A1(n9277), .A2(n6058), .ZN(n5979) );
  AOI21_X1 U7536 ( .B1(n9300), .B2(n6049), .A(n5979), .ZN(n5985) );
  NAND2_X1 U7537 ( .A1(n9392), .A2(n6052), .ZN(n5981) );
  NAND2_X1 U7538 ( .A1(n9396), .A2(n5871), .ZN(n5980) );
  NAND2_X1 U7539 ( .A1(n5981), .A2(n5980), .ZN(n5982) );
  XNOR2_X1 U7540 ( .A(n5982), .B(n4371), .ZN(n5988) );
  NAND2_X1 U7541 ( .A1(n9392), .A2(n5871), .ZN(n5984) );
  NAND2_X1 U7542 ( .A1(n9396), .A2(n6011), .ZN(n5983) );
  NAND2_X1 U7543 ( .A1(n5984), .A2(n5983), .ZN(n5989) );
  NAND2_X1 U7544 ( .A1(n5988), .A2(n5989), .ZN(n8806) );
  INV_X1 U7545 ( .A(n8808), .ZN(n5986) );
  INV_X1 U7546 ( .A(n5985), .ZN(n8916) );
  NAND2_X1 U7547 ( .A1(n5986), .A2(n8916), .ZN(n5987) );
  INV_X1 U7548 ( .A(n5988), .ZN(n5991) );
  INV_X1 U7549 ( .A(n5989), .ZN(n5990) );
  NAND2_X1 U7550 ( .A1(n5991), .A2(n5990), .ZN(n8805) );
  NAND2_X1 U7551 ( .A1(n5992), .A2(n8805), .ZN(n8889) );
  NAND2_X1 U7552 ( .A1(n9388), .A2(n6052), .ZN(n5994) );
  INV_X1 U7553 ( .A(n9278), .ZN(n9377) );
  NAND2_X1 U7554 ( .A1(n9377), .A2(n6049), .ZN(n5993) );
  NAND2_X1 U7555 ( .A1(n5994), .A2(n5993), .ZN(n5995) );
  XNOR2_X1 U7556 ( .A(n5995), .B(n6055), .ZN(n8887) );
  NOR2_X1 U7557 ( .A1(n9278), .A2(n6058), .ZN(n5996) );
  AOI21_X1 U7558 ( .B1(n9388), .B2(n6049), .A(n5996), .ZN(n8886) );
  AND2_X1 U7559 ( .A1(n8887), .A2(n8886), .ZN(n5997) );
  INV_X1 U7560 ( .A(n8887), .ZN(n5999) );
  INV_X1 U7561 ( .A(n8886), .ZN(n5998) );
  NAND2_X1 U7562 ( .A1(n5999), .A2(n5998), .ZN(n6000) );
  NAND2_X1 U7563 ( .A1(n9241), .A2(n6052), .ZN(n6002) );
  OR2_X1 U7564 ( .A1(n9255), .A2(n5892), .ZN(n6001) );
  NAND2_X1 U7565 ( .A1(n6002), .A2(n6001), .ZN(n6003) );
  XNOR2_X1 U7566 ( .A(n6003), .B(n6055), .ZN(n6006) );
  NOR2_X1 U7567 ( .A1(n9255), .A2(n6058), .ZN(n6004) );
  AOI21_X1 U7568 ( .B1(n9241), .B2(n6049), .A(n6004), .ZN(n6005) );
  XNOR2_X1 U7569 ( .A(n6006), .B(n6005), .ZN(n8829) );
  NAND2_X1 U7570 ( .A1(n6006), .A2(n6005), .ZN(n6007) );
  NAND2_X1 U7571 ( .A1(n9233), .A2(n6052), .ZN(n6009) );
  NAND2_X1 U7572 ( .A1(n9378), .A2(n5871), .ZN(n6008) );
  NAND2_X1 U7573 ( .A1(n6009), .A2(n6008), .ZN(n6010) );
  XNOR2_X1 U7574 ( .A(n6010), .B(n6055), .ZN(n6014) );
  NAND2_X1 U7575 ( .A1(n9233), .A2(n5871), .ZN(n6013) );
  NAND2_X1 U7576 ( .A1(n9378), .A2(n6011), .ZN(n6012) );
  NAND2_X1 U7577 ( .A1(n6013), .A2(n6012), .ZN(n8904) );
  NAND2_X1 U7578 ( .A1(n9363), .A2(n6052), .ZN(n6017) );
  OR2_X1 U7579 ( .A1(n9199), .A2(n5892), .ZN(n6016) );
  NAND2_X1 U7580 ( .A1(n6017), .A2(n6016), .ZN(n6018) );
  XNOR2_X1 U7581 ( .A(n6018), .B(n6055), .ZN(n6021) );
  NOR2_X1 U7582 ( .A1(n9199), .A2(n6058), .ZN(n6019) );
  AOI21_X1 U7583 ( .B1(n9363), .B2(n6049), .A(n6019), .ZN(n6020) );
  NAND2_X1 U7584 ( .A1(n6021), .A2(n6020), .ZN(n8878) );
  OR2_X1 U7585 ( .A1(n6021), .A2(n6020), .ZN(n6022) );
  AND2_X1 U7586 ( .A1(n8878), .A2(n6022), .ZN(n8797) );
  NAND2_X1 U7587 ( .A1(n9201), .A2(n6052), .ZN(n6024) );
  INV_X1 U7588 ( .A(n9360), .ZN(n9344) );
  NAND2_X1 U7589 ( .A1(n9344), .A2(n5871), .ZN(n6023) );
  NAND2_X1 U7590 ( .A1(n6024), .A2(n6023), .ZN(n6025) );
  XNOR2_X1 U7591 ( .A(n6025), .B(n6055), .ZN(n6028) );
  NOR2_X1 U7592 ( .A1(n9360), .A2(n6058), .ZN(n6026) );
  AOI21_X1 U7593 ( .B1(n9201), .B2(n6049), .A(n6026), .ZN(n6027) );
  NAND2_X1 U7594 ( .A1(n6028), .A2(n6027), .ZN(n6030) );
  OR2_X1 U7595 ( .A1(n6028), .A2(n6027), .ZN(n6029) );
  NAND2_X1 U7596 ( .A1(n6030), .A2(n6029), .ZN(n8877) );
  INV_X1 U7597 ( .A(n6030), .ZN(n6031) );
  NAND2_X1 U7598 ( .A1(n9185), .A2(n6052), .ZN(n6033) );
  NAND2_X1 U7599 ( .A1(n9196), .A2(n5871), .ZN(n6032) );
  NAND2_X1 U7600 ( .A1(n6033), .A2(n6032), .ZN(n6034) );
  XNOR2_X1 U7601 ( .A(n6034), .B(n4371), .ZN(n6036) );
  OAI22_X1 U7602 ( .A1(n9348), .A2(n5892), .B1(n9334), .B2(n6058), .ZN(n6035)
         );
  XNOR2_X1 U7603 ( .A(n6036), .B(n6035), .ZN(n8843) );
  NOR2_X1 U7604 ( .A1(n6036), .A2(n6035), .ZN(n8923) );
  NAND2_X1 U7605 ( .A1(n9164), .A2(n6052), .ZN(n6038) );
  OR2_X1 U7606 ( .A1(n9324), .A2(n5892), .ZN(n6037) );
  NAND2_X1 U7607 ( .A1(n6038), .A2(n6037), .ZN(n6039) );
  XNOR2_X1 U7608 ( .A(n6039), .B(n6055), .ZN(n6041) );
  NOR2_X1 U7609 ( .A1(n9324), .A2(n6058), .ZN(n6040) );
  AOI21_X1 U7610 ( .B1(n9164), .B2(n6049), .A(n6040), .ZN(n6042) );
  XNOR2_X1 U7611 ( .A(n6041), .B(n6042), .ZN(n8922) );
  INV_X1 U7612 ( .A(n6041), .ZN(n6044) );
  INV_X1 U7613 ( .A(n6042), .ZN(n6043) );
  NAND2_X1 U7614 ( .A1(n9156), .A2(n6052), .ZN(n6046) );
  OR2_X1 U7615 ( .A1(n9335), .A2(n5892), .ZN(n6045) );
  NAND2_X1 U7616 ( .A1(n6046), .A2(n6045), .ZN(n6047) );
  XNOR2_X1 U7617 ( .A(n6047), .B(n6055), .ZN(n6051) );
  NOR2_X1 U7618 ( .A1(n9335), .A2(n6058), .ZN(n6048) );
  AOI21_X1 U7619 ( .B1(n9156), .B2(n6049), .A(n6048), .ZN(n6050) );
  NAND2_X1 U7620 ( .A1(n6051), .A2(n6050), .ZN(n6090) );
  OAI21_X1 U7621 ( .B1(n6051), .B2(n6050), .A(n6090), .ZN(n8780) );
  NAND2_X1 U7622 ( .A1(n9318), .A2(n6052), .ZN(n6054) );
  OR2_X1 U7623 ( .A1(n9325), .A2(n5892), .ZN(n6053) );
  NAND2_X1 U7624 ( .A1(n6054), .A2(n6053), .ZN(n6056) );
  XNOR2_X1 U7625 ( .A(n6056), .B(n6055), .ZN(n6060) );
  NAND2_X1 U7626 ( .A1(n9318), .A2(n5871), .ZN(n6057) );
  OAI21_X1 U7627 ( .B1(n9325), .B2(n6058), .A(n6057), .ZN(n6059) );
  XNOR2_X1 U7628 ( .A(n6060), .B(n6059), .ZN(n6076) );
  NOR2_X1 U7629 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .ZN(
        n6064) );
  NOR4_X1 U7630 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n6063) );
  NOR4_X1 U7631 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n6062) );
  NOR4_X1 U7632 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n6061) );
  NAND4_X1 U7633 ( .A1(n6064), .A2(n6063), .A3(n6062), .A4(n6061), .ZN(n6070)
         );
  NOR4_X1 U7634 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n6068) );
  NOR4_X1 U7635 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n6067) );
  NOR4_X1 U7636 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n6066) );
  NOR4_X1 U7637 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n6065) );
  NAND4_X1 U7638 ( .A1(n6068), .A2(n6067), .A3(n6066), .A4(n6065), .ZN(n6069)
         );
  NOR2_X1 U7639 ( .A1(n6070), .A2(n6069), .ZN(n6688) );
  INV_X1 U7640 ( .A(n6073), .ZN(n7740) );
  NAND2_X1 U7641 ( .A1(n7740), .A2(P1_B_REG_SCAN_IN), .ZN(n6071) );
  MUX2_X1 U7642 ( .A(P1_B_REG_SCAN_IN), .B(n6071), .S(n7703), .Z(n6072) );
  NAND2_X1 U7643 ( .A1(n6072), .A2(n6074), .ZN(n6687) );
  INV_X1 U7644 ( .A(n6074), .ZN(n7786) );
  NAND2_X1 U7645 ( .A1(n7703), .A2(n7786), .ZN(n9469) );
  OR2_X1 U7646 ( .A1(n6074), .A2(n6073), .ZN(n9468) );
  OAI21_X1 U7647 ( .B1(n6687), .B2(P1_D_REG_1__SCAN_IN), .A(n9468), .ZN(n6847)
         );
  INV_X1 U7648 ( .A(n6847), .ZN(n6693) );
  OAI211_X1 U7649 ( .C1(n6688), .C2(n6687), .A(n6850), .B(n6693), .ZN(n6083)
         );
  NAND2_X1 U7650 ( .A1(n9768), .A2(n6699), .ZN(n6075) );
  NOR2_X2 U7651 ( .A1(n6082), .A2(n6075), .ZN(n8936) );
  NAND3_X1 U7652 ( .A1(n8783), .A2(n6076), .A3(n8936), .ZN(n6098) );
  INV_X1 U7653 ( .A(n6076), .ZN(n6091) );
  NAND3_X1 U7654 ( .A1(n6091), .A2(n8936), .A3(n6090), .ZN(n6077) );
  NAND2_X1 U7655 ( .A1(n9720), .A2(n6839), .ZN(n6712) );
  OR2_X1 U7656 ( .A1(n6082), .A2(n6712), .ZN(n6078) );
  NAND2_X1 U7657 ( .A1(n9319), .A2(n9080), .ZN(n6846) );
  NAND2_X2 U7658 ( .A1(n6078), .A2(n9242), .ZN(n8928) );
  NOR2_X2 U7659 ( .A1(n6699), .A2(n9564), .ZN(n9757) );
  NAND2_X1 U7660 ( .A1(n9757), .A2(n6080), .ZN(n6079) );
  NOR2_X2 U7661 ( .A1(n6082), .A2(n6079), .ZN(n8945) );
  NAND2_X1 U7662 ( .A1(n9754), .A2(n6080), .ZN(n6081) );
  NOR2_X2 U7663 ( .A1(n6082), .A2(n6081), .ZN(n8926) );
  AOI22_X1 U7664 ( .A1(n8926), .A2(n9166), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3086), .ZN(n6089) );
  NAND2_X1 U7665 ( .A1(n6083), .A2(n6846), .ZN(n6087) );
  NAND2_X1 U7666 ( .A1(n6084), .A2(n6698), .ZN(n6690) );
  AND3_X1 U7667 ( .A1(n6690), .A2(n6085), .A3(n5837), .ZN(n6086) );
  NAND2_X1 U7668 ( .A1(n6087), .A2(n6086), .ZN(n8869) );
  NAND2_X1 U7669 ( .A1(n8927), .A2(n9135), .ZN(n6088) );
  OAI211_X1 U7670 ( .C1(n8899), .C2(n8951), .A(n6089), .B(n6088), .ZN(n6093)
         );
  NOR3_X1 U7671 ( .A1(n6091), .A2(n6090), .A3(n8920), .ZN(n6092) );
  AOI211_X1 U7672 ( .C1(n9318), .C2(n8928), .A(n6093), .B(n6092), .ZN(n6094)
         );
  INV_X1 U7673 ( .A(n6094), .ZN(n6095) );
  NOR2_X1 U7674 ( .A1(n6096), .A2(n6095), .ZN(n6097) );
  NAND2_X1 U7675 ( .A1(n6098), .A2(n6097), .ZN(P1_U3220) );
  NOR2_X1 U7676 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_25__SCAN_IN), .ZN(
        n6111) );
  NOR2_X1 U7677 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), .ZN(
        n6110) );
  NOR2_X1 U7678 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_23__SCAN_IN), .ZN(
        n6109) );
  NOR2_X1 U7679 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), .ZN(
        n6108) );
  XNOR2_X2 U7680 ( .A(n6114), .B(n4978), .ZN(n6812) );
  NAND2_X1 U7681 ( .A1(n6540), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6116) );
  NAND2_X1 U7682 ( .A1(n7738), .A2(n8097), .ZN(n6119) );
  NAND2_X1 U7683 ( .A1(n6192), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n6118) );
  NAND2_X1 U7684 ( .A1(n10069), .A2(n10128), .ZN(n6229) );
  INV_X1 U7685 ( .A(n6229), .ZN(n6121) );
  NAND2_X1 U7686 ( .A1(n6121), .A2(n6120), .ZN(n6241) );
  INV_X1 U7687 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n6125) );
  INV_X1 U7688 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n6128) );
  INV_X1 U7689 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n10045) );
  INV_X1 U7690 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n10055) );
  INV_X1 U7691 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n6130) );
  NAND2_X1 U7692 ( .A1(n6431), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n6132) );
  NAND2_X1 U7693 ( .A1(n6441), .A2(n6132), .ZN(n8478) );
  NAND2_X1 U7694 ( .A1(n8478), .A2(n6170), .ZN(n6144) );
  INV_X1 U7695 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n6141) );
  INV_X1 U7696 ( .A(n6135), .ZN(n6138) );
  NAND2_X2 U7697 ( .A1(n6138), .A2(n6136), .ZN(n7350) );
  NAND2_X1 U7698 ( .A1(n6475), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n6140) );
  NAND2_X1 U7699 ( .A1(n6514), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n6139) );
  OAI211_X1 U7700 ( .C1(n6141), .C2(n6186), .A(n6140), .B(n6139), .ZN(n6142)
         );
  INV_X1 U7701 ( .A(n6142), .ZN(n6143) );
  NAND2_X1 U7702 ( .A1(n7545), .A2(n8097), .ZN(n6146) );
  NAND2_X1 U7703 ( .A1(n6192), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n6145) );
  NAND2_X1 U7704 ( .A1(n6415), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6147) );
  NAND2_X1 U7705 ( .A1(n6421), .A2(n6147), .ZN(n8514) );
  NAND2_X1 U7706 ( .A1(n8514), .A2(n6170), .ZN(n6150) );
  AOI22_X1 U7707 ( .A1(n6514), .A2(P2_REG1_REG_22__SCAN_IN), .B1(n6475), .B2(
        P2_REG0_REG_22__SCAN_IN), .ZN(n6149) );
  NAND2_X1 U7708 ( .A1(n6423), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n6148) );
  NAND2_X1 U7709 ( .A1(n6475), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n6155) );
  INV_X1 U7710 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n7878) );
  OR2_X1 U7711 ( .A1(n7348), .A2(n7878), .ZN(n6154) );
  INV_X1 U7712 ( .A(n6170), .ZN(n6396) );
  NAND2_X1 U7713 ( .A1(n6395), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n6151) );
  AND2_X1 U7714 ( .A1(n6404), .A2(n6151), .ZN(n7973) );
  OR2_X1 U7715 ( .A1(n6396), .A2(n7973), .ZN(n6153) );
  INV_X1 U7716 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n7882) );
  OR2_X1 U7717 ( .A1(n6186), .A2(n7882), .ZN(n6152) );
  INV_X1 U7718 ( .A(n8547), .ZN(n8537) );
  NAND2_X1 U7719 ( .A1(n7222), .A2(n8097), .ZN(n6161) );
  INV_X1 U7720 ( .A(n6482), .ZN(n6158) );
  NAND2_X1 U7721 ( .A1(n6158), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6159) );
  AOI22_X1 U7722 ( .A1(n6192), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n6527), .B2(
        n6585), .ZN(n6160) );
  INV_X1 U7723 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n7226) );
  OR2_X1 U7724 ( .A1(n7350), .A2(n7226), .ZN(n6167) );
  INV_X1 U7725 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n6162) );
  INV_X1 U7726 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n6163) );
  OR2_X1 U7727 ( .A1(n7348), .A2(n6163), .ZN(n6165) );
  INV_X1 U7728 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n7297) );
  NAND2_X1 U7729 ( .A1(n4810), .A2(SI_0_), .ZN(n6168) );
  XNOR2_X1 U7730 ( .A(n6168), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n8779) );
  MUX2_X1 U7731 ( .A(P2_IR_REG_0__SCAN_IN), .B(n8779), .S(n6521), .Z(n7300) );
  NAND2_X1 U7732 ( .A1(n8326), .A2(n7300), .ZN(n7460) );
  INV_X1 U7733 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n6871) );
  OR2_X1 U7734 ( .A1(n7348), .A2(n6871), .ZN(n6174) );
  INV_X1 U7735 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n6169) );
  OR2_X1 U7736 ( .A1(n7350), .A2(n6169), .ZN(n6173) );
  NAND2_X1 U7737 ( .A1(n6170), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n6172) );
  INV_X1 U7738 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n7462) );
  OR2_X1 U7739 ( .A1(n6186), .A2(n7462), .ZN(n6171) );
  NAND2_X1 U7740 ( .A1(n6192), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n6180) );
  NAND2_X1 U7741 ( .A1(n6247), .A2(n6175), .ZN(n6179) );
  NAND2_X1 U7742 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n6176) );
  XNOR2_X1 U7743 ( .A(n6176), .B(P2_IR_REG_1__SCAN_IN), .ZN(n6892) );
  INV_X1 U7744 ( .A(n6892), .ZN(n6177) );
  NAND2_X1 U7745 ( .A1(n7460), .A2(n8108), .ZN(n6185) );
  OR2_X1 U7746 ( .A1(n6183), .A2(n6181), .ZN(n6184) );
  NAND2_X1 U7747 ( .A1(n6185), .A2(n6184), .ZN(n7208) );
  NAND2_X1 U7748 ( .A1(n6475), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n6191) );
  INV_X1 U7749 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n7346) );
  INV_X1 U7750 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n7214) );
  OR2_X1 U7751 ( .A1(n6186), .A2(n7214), .ZN(n6189) );
  INV_X1 U7752 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n6187) );
  OR2_X1 U7753 ( .A1(n7348), .A2(n6187), .ZN(n6188) );
  NAND2_X1 U7754 ( .A1(n6192), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n6197) );
  NAND2_X1 U7755 ( .A1(n6247), .A2(n6193), .ZN(n6196) );
  NAND2_X1 U7756 ( .A1(n8325), .A2(n9869), .ZN(n8144) );
  NAND2_X1 U7757 ( .A1(n7208), .A2(n8107), .ZN(n6201) );
  OR2_X1 U7758 ( .A1(n8325), .A2(n6198), .ZN(n6200) );
  NAND2_X1 U7759 ( .A1(n6201), .A2(n6200), .ZN(n6805) );
  NAND2_X1 U7760 ( .A1(n6475), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n6207) );
  INV_X1 U7761 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n6202) );
  OR2_X1 U7762 ( .A1(n6186), .A2(n6202), .ZN(n6205) );
  INV_X1 U7763 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n6203) );
  OR2_X1 U7764 ( .A1(n7348), .A2(n6203), .ZN(n6204) );
  NAND2_X1 U7765 ( .A1(n6192), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n6213) );
  NAND2_X1 U7766 ( .A1(n6247), .A2(n6208), .ZN(n6212) );
  NAND2_X1 U7767 ( .A1(n6209), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6210) );
  NAND2_X1 U7768 ( .A1(n6585), .A2(n4488), .ZN(n6211) );
  NAND2_X1 U7769 ( .A1(n8324), .A2(n7507), .ZN(n8160) );
  NAND2_X1 U7770 ( .A1(n8167), .A2(n8160), .ZN(n8110) );
  INV_X1 U7771 ( .A(n7507), .ZN(n7170) );
  OR2_X1 U7772 ( .A1(n8324), .A2(n7170), .ZN(n6214) );
  NAND2_X1 U7773 ( .A1(n6514), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6220) );
  INV_X1 U7774 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n6215) );
  OR2_X1 U7775 ( .A1(n7350), .A2(n6215), .ZN(n6219) );
  NAND2_X1 U7776 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n6216) );
  AND2_X1 U7777 ( .A1(n6229), .A2(n6216), .ZN(n7492) );
  OR2_X1 U7778 ( .A1(n6396), .A2(n7492), .ZN(n6218) );
  INV_X1 U7779 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n6884) );
  OR2_X1 U7780 ( .A1(n6186), .A2(n6884), .ZN(n6217) );
  INV_X1 U7781 ( .A(n6247), .ZN(n6225) );
  NAND2_X1 U7782 ( .A1(n6192), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n6224) );
  NAND2_X1 U7783 ( .A1(n6221), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6222) );
  NAND2_X1 U7784 ( .A1(n6585), .A2(n6899), .ZN(n6223) );
  OAI211_X1 U7785 ( .C1(n6225), .C2(n6604), .A(n6224), .B(n6223), .ZN(n7232)
         );
  NAND2_X1 U7786 ( .A1(n8323), .A2(n7232), .ZN(n6226) );
  NAND2_X1 U7787 ( .A1(n6227), .A2(n6226), .ZN(n7324) );
  NAND2_X1 U7788 ( .A1(n6475), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n6235) );
  INV_X1 U7789 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n6228) );
  OR2_X1 U7790 ( .A1(n6186), .A2(n6228), .ZN(n6234) );
  NAND2_X1 U7791 ( .A1(n6229), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n6230) );
  AND2_X1 U7792 ( .A1(n6241), .A2(n6230), .ZN(n7500) );
  OR2_X1 U7793 ( .A1(n6396), .A2(n7500), .ZN(n6233) );
  INV_X1 U7794 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n6231) );
  OR2_X1 U7795 ( .A1(n7348), .A2(n6231), .ZN(n6232) );
  NAND4_X1 U7796 ( .A1(n6235), .A2(n6234), .A3(n6233), .A4(n6232), .ZN(n8322)
         );
  NAND2_X1 U7797 ( .A1(n6192), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n6239) );
  OR2_X1 U7798 ( .A1(n6236), .A2(n8764), .ZN(n6237) );
  XNOR2_X1 U7799 ( .A(n6237), .B(P2_IR_REG_5__SCAN_IN), .ZN(n6905) );
  NAND2_X1 U7800 ( .A1(n6585), .A2(n6905), .ZN(n6238) );
  OAI211_X1 U7801 ( .C1(n6225), .C2(n6594), .A(n6239), .B(n6238), .ZN(n7336)
         );
  AND2_X1 U7802 ( .A1(n8322), .A2(n7336), .ZN(n6240) );
  NAND2_X1 U7803 ( .A1(n6475), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n6246) );
  OR2_X1 U7804 ( .A1(n7348), .A2(n9919), .ZN(n6245) );
  NAND2_X1 U7805 ( .A1(n6241), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n6242) );
  AND2_X1 U7806 ( .A1(n6256), .A2(n6242), .ZN(n7481) );
  OR2_X1 U7807 ( .A1(n6396), .A2(n7481), .ZN(n6244) );
  INV_X1 U7808 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n6992) );
  OR2_X1 U7809 ( .A1(n6186), .A2(n6992), .ZN(n6243) );
  NAND4_X1 U7810 ( .A1(n6246), .A2(n6245), .A3(n6244), .A4(n6243), .ZN(n8321)
         );
  NAND2_X1 U7811 ( .A1(n6247), .A2(n6596), .ZN(n6254) );
  NAND2_X1 U7812 ( .A1(n6192), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n6253) );
  NAND2_X1 U7813 ( .A1(n6248), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6249) );
  MUX2_X1 U7814 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6249), .S(
        P2_IR_REG_6__SCAN_IN), .Z(n6251) );
  INV_X1 U7815 ( .A(n6250), .ZN(n6262) );
  AND2_X1 U7816 ( .A1(n6251), .A2(n6262), .ZN(n6993) );
  NAND2_X1 U7817 ( .A1(n6585), .A2(n6993), .ZN(n6252) );
  OR2_X1 U7818 ( .A1(n8321), .A2(n9879), .ZN(n8163) );
  NAND2_X1 U7819 ( .A1(n8321), .A2(n9879), .ZN(n8172) );
  INV_X1 U7820 ( .A(n9879), .ZN(n7396) );
  NAND2_X1 U7821 ( .A1(n8321), .A2(n7396), .ZN(n6255) );
  NAND2_X1 U7822 ( .A1(n6475), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n6261) );
  INV_X1 U7823 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n6969) );
  OR2_X1 U7824 ( .A1(n7348), .A2(n6969), .ZN(n6260) );
  NAND2_X1 U7825 ( .A1(n6256), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n6257) );
  AND2_X1 U7826 ( .A1(n6269), .A2(n6257), .ZN(n7606) );
  OR2_X1 U7827 ( .A1(n6396), .A2(n7606), .ZN(n6259) );
  INV_X1 U7828 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n6970) );
  OR2_X1 U7829 ( .A1(n6186), .A2(n6970), .ZN(n6258) );
  NAND4_X1 U7830 ( .A1(n6261), .A2(n6260), .A3(n6259), .A4(n6258), .ZN(n8320)
         );
  NAND2_X1 U7831 ( .A1(n6192), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n6267) );
  NAND2_X1 U7832 ( .A1(n6262), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6263) );
  MUX2_X1 U7833 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6263), .S(
        P2_IR_REG_7__SCAN_IN), .Z(n6265) );
  AND2_X1 U7834 ( .A1(n6265), .A2(n6264), .ZN(n7051) );
  NAND2_X1 U7835 ( .A1(n6585), .A2(n7051), .ZN(n6266) );
  OAI211_X1 U7836 ( .C1(n6225), .C2(n6607), .A(n6267), .B(n6266), .ZN(n7542)
         );
  XNOR2_X1 U7837 ( .A(n8320), .B(n7542), .ZN(n8179) );
  NAND2_X1 U7838 ( .A1(n6475), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n6274) );
  INV_X1 U7839 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n9922) );
  OR2_X1 U7840 ( .A1(n7348), .A2(n9922), .ZN(n6273) );
  NAND2_X1 U7841 ( .A1(n6269), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n6270) );
  AND2_X1 U7842 ( .A1(n6281), .A2(n6270), .ZN(n7603) );
  OR2_X1 U7843 ( .A1(n6396), .A2(n7603), .ZN(n6272) );
  INV_X1 U7844 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n6988) );
  OR2_X1 U7845 ( .A1(n6186), .A2(n6988), .ZN(n6271) );
  NAND4_X1 U7846 ( .A1(n6274), .A2(n6273), .A3(n6272), .A4(n6271), .ZN(n8319)
         );
  NAND2_X1 U7847 ( .A1(n8097), .A2(n6609), .ZN(n6278) );
  NAND2_X1 U7848 ( .A1(n6192), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n6277) );
  NAND2_X1 U7849 ( .A1(n6264), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6275) );
  XNOR2_X1 U7850 ( .A(n6275), .B(P2_IR_REG_8__SCAN_IN), .ZN(n6989) );
  NAND2_X1 U7851 ( .A1(n6585), .A2(n6989), .ZN(n6276) );
  NAND2_X1 U7852 ( .A1(n8319), .A2(n9890), .ZN(n8181) );
  NAND2_X1 U7853 ( .A1(n8187), .A2(n8181), .ZN(n8116) );
  OR2_X1 U7854 ( .A1(n8320), .A2(n7542), .ZN(n7448) );
  AND2_X1 U7855 ( .A1(n8116), .A2(n7448), .ZN(n6279) );
  NAND2_X1 U7856 ( .A1(n7609), .A2(n6279), .ZN(n7449) );
  INV_X1 U7857 ( .A(n9890), .ZN(n7600) );
  NAND2_X1 U7858 ( .A1(n8319), .A2(n7600), .ZN(n6280) );
  NAND2_X1 U7859 ( .A1(n6475), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n6286) );
  INV_X1 U7860 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7063) );
  OR2_X1 U7861 ( .A1(n6186), .A2(n7063), .ZN(n6285) );
  NAND2_X1 U7862 ( .A1(n6281), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n6282) );
  AND2_X1 U7863 ( .A1(n6299), .A2(n6282), .ZN(n7663) );
  OR2_X1 U7864 ( .A1(n6396), .A2(n7663), .ZN(n6284) );
  INV_X1 U7865 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n7062) );
  OR2_X1 U7866 ( .A1(n7348), .A2(n7062), .ZN(n6283) );
  NAND4_X1 U7867 ( .A1(n6286), .A2(n6285), .A3(n6284), .A4(n6283), .ZN(n8318)
         );
  NAND2_X1 U7868 ( .A1(n6613), .A2(n8097), .ZN(n6289) );
  NOR2_X1 U7869 ( .A1(n6264), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n6292) );
  OR2_X1 U7870 ( .A1(n6292), .A2(n8764), .ZN(n6287) );
  XNOR2_X1 U7871 ( .A(n6287), .B(P2_IR_REG_9__SCAN_IN), .ZN(n7112) );
  AOI22_X1 U7872 ( .A1(n6192), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6585), .B2(
        n7112), .ZN(n6288) );
  OR2_X1 U7873 ( .A1(n8318), .A2(n7679), .ZN(n8188) );
  NAND2_X1 U7874 ( .A1(n8318), .A2(n7679), .ZN(n8183) );
  NAND2_X1 U7875 ( .A1(n8188), .A2(n8183), .ZN(n8118) );
  NAND2_X1 U7876 ( .A1(n7557), .A2(n8118), .ZN(n7556) );
  INV_X1 U7877 ( .A(n7679), .ZN(n7682) );
  OR2_X1 U7878 ( .A1(n8318), .A2(n7682), .ZN(n6290) );
  NAND2_X1 U7879 ( .A1(n7556), .A2(n6290), .ZN(n7664) );
  NAND2_X1 U7880 ( .A1(n6615), .A2(n8097), .ZN(n6298) );
  INV_X1 U7881 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n6291) );
  NOR2_X1 U7882 ( .A1(n6295), .A2(n8764), .ZN(n6293) );
  MUX2_X1 U7883 ( .A(n8764), .B(n6293), .S(P2_IR_REG_10__SCAN_IN), .Z(n6296)
         );
  INV_X1 U7884 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n6294) );
  AOI22_X1 U7885 ( .A1(n6192), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6585), .B2(
        n7118), .ZN(n6297) );
  NAND2_X1 U7886 ( .A1(n6298), .A2(n6297), .ZN(n7776) );
  NAND2_X1 U7887 ( .A1(n6475), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n6304) );
  INV_X1 U7888 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7115) );
  OR2_X1 U7889 ( .A1(n6186), .A2(n7115), .ZN(n6303) );
  NAND2_X1 U7890 ( .A1(n6299), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n6300) );
  AND2_X1 U7891 ( .A1(n6307), .A2(n6300), .ZN(n7670) );
  OR2_X1 U7892 ( .A1(n6396), .A2(n7670), .ZN(n6302) );
  INV_X1 U7893 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n9924) );
  OR2_X1 U7894 ( .A1(n7348), .A2(n9924), .ZN(n6301) );
  NAND4_X1 U7895 ( .A1(n6304), .A2(n6303), .A3(n6302), .A4(n6301), .ZN(n8317)
         );
  NOR2_X1 U7896 ( .A1(n7776), .A2(n8317), .ZN(n6305) );
  INV_X1 U7897 ( .A(n7776), .ZN(n9895) );
  OAI22_X1 U7898 ( .A1(n7664), .A2(n6305), .B1(n9895), .B2(n7788), .ZN(n7731)
         );
  NAND2_X1 U7899 ( .A1(n6475), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n6313) );
  INV_X1 U7900 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n6306) );
  OR2_X1 U7901 ( .A1(n7348), .A2(n6306), .ZN(n6312) );
  NAND2_X1 U7902 ( .A1(n6307), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6308) );
  AND2_X1 U7903 ( .A1(n6323), .A2(n6308), .ZN(n7795) );
  OR2_X1 U7904 ( .A1(n6396), .A2(n7795), .ZN(n6311) );
  INV_X1 U7905 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n6309) );
  OR2_X1 U7906 ( .A1(n6186), .A2(n6309), .ZN(n6310) );
  NAND4_X1 U7907 ( .A1(n6313), .A2(n6312), .A3(n6311), .A4(n6310), .ZN(n8316)
         );
  NAND2_X1 U7908 ( .A1(n6628), .A2(n8097), .ZN(n6316) );
  OR2_X1 U7909 ( .A1(n6318), .A2(n8764), .ZN(n6314) );
  XNOR2_X1 U7910 ( .A(n6314), .B(P2_IR_REG_11__SCAN_IN), .ZN(n7370) );
  AOI22_X1 U7911 ( .A1(n6192), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n6585), .B2(
        n7370), .ZN(n6315) );
  NAND2_X1 U7912 ( .A1(n6632), .A2(n8097), .ZN(n6321) );
  INV_X1 U7913 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n6317) );
  NAND2_X1 U7914 ( .A1(n6318), .A2(n6317), .ZN(n6330) );
  NAND2_X1 U7915 ( .A1(n6330), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6319) );
  XNOR2_X1 U7916 ( .A(n6319), .B(P2_IR_REG_12__SCAN_IN), .ZN(n7579) );
  AOI22_X1 U7917 ( .A1(n6192), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6585), .B2(
        n7579), .ZN(n6320) );
  NAND2_X1 U7918 ( .A1(n6321), .A2(n6320), .ZN(n9912) );
  NAND2_X1 U7919 ( .A1(n6514), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n6328) );
  INV_X1 U7920 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n6322) );
  OR2_X1 U7921 ( .A1(n7350), .A2(n6322), .ZN(n6327) );
  NAND2_X1 U7922 ( .A1(n6323), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n6324) );
  AND2_X1 U7923 ( .A1(n6334), .A2(n6324), .ZN(n7855) );
  OR2_X1 U7924 ( .A1(n6396), .A2(n7855), .ZN(n6326) );
  INV_X1 U7925 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n7755) );
  OR2_X1 U7926 ( .A1(n6186), .A2(n7755), .ZN(n6325) );
  NAND2_X1 U7927 ( .A1(n9912), .A2(n8619), .ZN(n8208) );
  INV_X1 U7928 ( .A(n8619), .ZN(n8315) );
  NAND2_X1 U7929 ( .A1(n9912), .A2(n8315), .ZN(n6329) );
  NAND2_X1 U7930 ( .A1(n6636), .A2(n8097), .ZN(n6333) );
  NAND2_X1 U7931 ( .A1(n6331), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6341) );
  AOI22_X1 U7932 ( .A1(n6192), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6585), .B2(
        n8351), .ZN(n6332) );
  NAND2_X1 U7933 ( .A1(n6333), .A2(n6332), .ZN(n8623) );
  NAND2_X1 U7934 ( .A1(n6475), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n6339) );
  INV_X1 U7935 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n7568) );
  OR2_X1 U7936 ( .A1(n7348), .A2(n7568), .ZN(n6338) );
  NAND2_X1 U7937 ( .A1(n6334), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n6335) );
  AND2_X1 U7938 ( .A1(n6346), .A2(n6335), .ZN(n8625) );
  OR2_X1 U7939 ( .A1(n6396), .A2(n8625), .ZN(n6337) );
  INV_X1 U7940 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n7569) );
  OR2_X1 U7941 ( .A1(n6186), .A2(n7569), .ZN(n6336) );
  NAND4_X1 U7942 ( .A1(n6339), .A2(n6338), .A3(n6337), .A4(n6336), .ZN(n8314)
         );
  AND2_X1 U7943 ( .A1(n8623), .A2(n8314), .ZN(n8212) );
  OR2_X1 U7944 ( .A1(n8623), .A2(n8314), .ZN(n8210) );
  NAND2_X1 U7945 ( .A1(n6640), .A2(n8097), .ZN(n6344) );
  INV_X1 U7946 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n6340) );
  NAND2_X1 U7947 ( .A1(n6341), .A2(n6340), .ZN(n6342) );
  NAND2_X1 U7948 ( .A1(n6342), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6354) );
  XNOR2_X1 U7949 ( .A(n6354), .B(P2_IR_REG_14__SCAN_IN), .ZN(n8354) );
  AOI22_X1 U7950 ( .A1(n6192), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n6585), .B2(
        n8354), .ZN(n6343) );
  NAND2_X1 U7951 ( .A1(n6344), .A2(n6343), .ZN(n8609) );
  NAND2_X1 U7952 ( .A1(n6475), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n6352) );
  INV_X1 U7953 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n6345) );
  OR2_X1 U7954 ( .A1(n7348), .A2(n6345), .ZN(n6351) );
  NAND2_X1 U7955 ( .A1(n6346), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n6347) );
  AND2_X1 U7956 ( .A1(n6359), .A2(n6347), .ZN(n8610) );
  OR2_X1 U7957 ( .A1(n6396), .A2(n8610), .ZN(n6350) );
  INV_X1 U7958 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n6348) );
  OR2_X1 U7959 ( .A1(n6186), .A2(n6348), .ZN(n6349) );
  OR2_X1 U7960 ( .A1(n8609), .A2(n8621), .ZN(n8217) );
  NAND2_X1 U7961 ( .A1(n8609), .A2(n8621), .ZN(n6499) );
  NAND2_X1 U7962 ( .A1(n6652), .A2(n8097), .ZN(n6358) );
  INV_X1 U7963 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n6353) );
  NAND2_X1 U7964 ( .A1(n6354), .A2(n6353), .ZN(n6355) );
  NAND2_X1 U7965 ( .A1(n6355), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6356) );
  XNOR2_X1 U7966 ( .A(n6356), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8392) );
  AOI22_X1 U7967 ( .A1(n6192), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n8392), .B2(
        n6585), .ZN(n6357) );
  NAND2_X1 U7968 ( .A1(n6475), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n6364) );
  INV_X1 U7969 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n8674) );
  OR2_X1 U7970 ( .A1(n7348), .A2(n8674), .ZN(n6363) );
  NAND2_X1 U7971 ( .A1(n6359), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n6360) );
  AND2_X1 U7972 ( .A1(n6379), .A2(n6360), .ZN(n8076) );
  OR2_X1 U7973 ( .A1(n6396), .A2(n8076), .ZN(n6362) );
  INV_X1 U7974 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n8597) );
  OR2_X1 U7975 ( .A1(n6186), .A2(n8597), .ZN(n6361) );
  NAND2_X1 U7976 ( .A1(n8757), .A2(n8608), .ZN(n8223) );
  NAND2_X1 U7977 ( .A1(n8570), .A2(n8223), .ZN(n8589) );
  NAND2_X1 U7978 ( .A1(n6365), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6366) );
  MUX2_X1 U7979 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6366), .S(
        P2_IR_REG_17__SCAN_IN), .Z(n6367) );
  INV_X1 U7980 ( .A(n6156), .ZN(n6389) );
  AND2_X1 U7981 ( .A1(n6367), .A2(n6389), .ZN(n9847) );
  AOI22_X1 U7982 ( .A1(n6192), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n6585), .B2(
        n9847), .ZN(n6368) );
  NAND2_X1 U7983 ( .A1(n6475), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n6374) );
  INV_X1 U7984 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n9850) );
  OR2_X1 U7985 ( .A1(n7348), .A2(n9850), .ZN(n6373) );
  NAND2_X1 U7986 ( .A1(n6381), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n6370) );
  AND2_X1 U7987 ( .A1(n6393), .A2(n6370), .ZN(n8008) );
  OR2_X1 U7988 ( .A1(n6396), .A2(n8008), .ZN(n6372) );
  INV_X1 U7989 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8565) );
  OR2_X1 U7990 ( .A1(n6186), .A2(n8565), .ZN(n6371) );
  INV_X1 U7991 ( .A(n8578), .ZN(n8312) );
  NAND2_X1 U7992 ( .A1(n8744), .A2(n8312), .ZN(n6386) );
  NAND2_X1 U7993 ( .A1(n8744), .A2(n8578), .ZN(n8230) );
  NAND2_X1 U7994 ( .A1(n6671), .A2(n8097), .ZN(n6378) );
  OR2_X1 U7995 ( .A1(n6375), .A2(n8764), .ZN(n6376) );
  XNOR2_X1 U7996 ( .A(n6376), .B(P2_IR_REG_16__SCAN_IN), .ZN(n8395) );
  AOI22_X1 U7997 ( .A1(n6192), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n6585), .B2(
        n8395), .ZN(n6377) );
  NAND2_X1 U7998 ( .A1(n6475), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n6385) );
  INV_X1 U7999 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8670) );
  OR2_X1 U8000 ( .A1(n7348), .A2(n8670), .ZN(n6384) );
  NAND2_X1 U8001 ( .A1(n6379), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n6380) );
  AND2_X1 U8002 ( .A1(n6381), .A2(n6380), .ZN(n7996) );
  OR2_X1 U8003 ( .A1(n6396), .A2(n7996), .ZN(n6383) );
  INV_X1 U8004 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8583) );
  OR2_X1 U8005 ( .A1(n6186), .A2(n8583), .ZN(n6382) );
  INV_X1 U8006 ( .A(n8082), .ZN(n8594) );
  NAND2_X1 U8007 ( .A1(n8750), .A2(n8594), .ZN(n8560) );
  AND2_X1 U8008 ( .A1(n8589), .A2(n6387), .ZN(n6388) );
  NAND2_X1 U8009 ( .A1(n8750), .A2(n8082), .ZN(n8226) );
  NAND2_X1 U8010 ( .A1(n8225), .A2(n8226), .ZN(n8222) );
  OR2_X1 U8011 ( .A1(n8757), .A2(n8313), .ZN(n8573) );
  AND2_X1 U8012 ( .A1(n8222), .A2(n8573), .ZN(n8559) );
  NAND2_X1 U8013 ( .A1(n6733), .A2(n8097), .ZN(n6392) );
  NAND2_X1 U8014 ( .A1(n6389), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6390) );
  XNOR2_X1 U8015 ( .A(n6390), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8412) );
  AOI22_X1 U8016 ( .A1(n6192), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6585), .B2(
        n8412), .ZN(n6391) );
  NAND2_X1 U8017 ( .A1(n6475), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n6400) );
  INV_X1 U8018 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8665) );
  OR2_X1 U8019 ( .A1(n7348), .A2(n8665), .ZN(n6399) );
  NAND2_X1 U8020 ( .A1(n6393), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n6394) );
  AND2_X1 U8021 ( .A1(n6395), .A2(n6394), .ZN(n8551) );
  OR2_X1 U8022 ( .A1(n6396), .A2(n8551), .ZN(n6398) );
  INV_X1 U8023 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8552) );
  OR2_X1 U8024 ( .A1(n6186), .A2(n8552), .ZN(n6397) );
  NAND4_X1 U8025 ( .A1(n6400), .A2(n6399), .A3(n6398), .A4(n6397), .ZN(n8563)
         );
  AND2_X1 U8026 ( .A1(n8063), .A2(n8563), .ZN(n6401) );
  OAI22_X1 U8027 ( .A1(n8545), .A2(n6401), .B1(n8063), .B2(n8563), .ZN(n7870)
         );
  NAND2_X1 U8028 ( .A1(n7381), .A2(n8097), .ZN(n6403) );
  NAND2_X1 U8029 ( .A1(n6192), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n6402) );
  NAND2_X1 U8030 ( .A1(n6404), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n6405) );
  NAND2_X1 U8031 ( .A1(n6413), .A2(n6405), .ZN(n8541) );
  NAND2_X1 U8032 ( .A1(n6170), .A2(n8541), .ZN(n6409) );
  INV_X1 U8033 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n8660) );
  OR2_X1 U8034 ( .A1(n7348), .A2(n8660), .ZN(n6408) );
  INV_X1 U8035 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n8732) );
  OR2_X1 U8036 ( .A1(n7350), .A2(n8732), .ZN(n6407) );
  INV_X1 U8037 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n8540) );
  OR2_X1 U8038 ( .A1(n6186), .A2(n8540), .ZN(n6406) );
  NAND2_X1 U8039 ( .A1(n8733), .A2(n8311), .ZN(n8245) );
  NAND2_X1 U8040 ( .A1(n8242), .A2(n8245), .ZN(n8535) );
  INV_X1 U8041 ( .A(n8733), .ZN(n6410) );
  NAND2_X1 U8042 ( .A1(n6410), .A2(n8311), .ZN(n8520) );
  NAND2_X1 U8043 ( .A1(n7407), .A2(n8097), .ZN(n6412) );
  NAND2_X1 U8044 ( .A1(n6192), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n6411) );
  NAND2_X1 U8045 ( .A1(n6413), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n6414) );
  NAND2_X1 U8046 ( .A1(n6415), .A2(n6414), .ZN(n8528) );
  AOI22_X1 U8047 ( .A1(n8528), .A2(n6170), .B1(n6423), .B2(
        P2_REG2_REG_21__SCAN_IN), .ZN(n6417) );
  AOI22_X1 U8048 ( .A1(n6514), .A2(P2_REG1_REG_21__SCAN_IN), .B1(n6475), .B2(
        P2_REG0_REG_21__SCAN_IN), .ZN(n6416) );
  NAND2_X1 U8049 ( .A1(n8727), .A2(n8030), .ZN(n8246) );
  NOR2_X1 U8050 ( .A1(n8727), .A2(n8538), .ZN(n8508) );
  NAND2_X1 U8051 ( .A1(n8721), .A2(n6418), .ZN(n8250) );
  NAND2_X1 U8052 ( .A1(n8236), .A2(n8250), .ZN(n8507) );
  OAI21_X1 U8053 ( .B1(n8721), .B2(n8525), .A(n8510), .ZN(n8497) );
  NAND2_X1 U8054 ( .A1(n7637), .A2(n8097), .ZN(n6420) );
  NAND2_X1 U8055 ( .A1(n6192), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n6419) );
  INV_X1 U8056 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n8651) );
  NAND2_X1 U8057 ( .A1(n6421), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6422) );
  NAND2_X1 U8058 ( .A1(n6429), .A2(n6422), .ZN(n8502) );
  NAND2_X1 U8059 ( .A1(n8502), .A2(n6170), .ZN(n6425) );
  AOI22_X1 U8060 ( .A1(n6423), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n6475), .B2(
        P2_REG0_REG_23__SCAN_IN), .ZN(n6424) );
  NAND2_X1 U8061 ( .A1(n8715), .A2(n8511), .ZN(n6426) );
  INV_X1 U8062 ( .A(n8715), .ZN(n6507) );
  NAND2_X1 U8063 ( .A1(n7699), .A2(n8097), .ZN(n6428) );
  NAND2_X1 U8064 ( .A1(n6192), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n6427) );
  NAND2_X1 U8065 ( .A1(n6429), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n6430) );
  NAND2_X1 U8066 ( .A1(n6431), .A2(n6430), .ZN(n8488) );
  NAND2_X1 U8067 ( .A1(n8488), .A2(n6170), .ZN(n6437) );
  INV_X1 U8068 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n6434) );
  NAND2_X1 U8069 ( .A1(n6514), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n6433) );
  NAND2_X1 U8070 ( .A1(n6475), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n6432) );
  OAI211_X1 U8071 ( .C1(n6434), .C2(n6186), .A(n6433), .B(n6432), .ZN(n6435)
         );
  INV_X1 U8072 ( .A(n6435), .ZN(n6436) );
  NAND2_X1 U8073 ( .A1(n8709), .A2(n8018), .ZN(n6438) );
  NAND2_X1 U8074 ( .A1(n8704), .A2(n8486), .ZN(n8260) );
  NAND2_X1 U8075 ( .A1(n7744), .A2(n8097), .ZN(n6440) );
  NAND2_X1 U8076 ( .A1(n6192), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n6439) );
  NAND2_X1 U8077 ( .A1(n6441), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n6442) );
  NAND2_X1 U8078 ( .A1(n8468), .A2(n6170), .ZN(n6447) );
  INV_X1 U8079 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n8467) );
  NAND2_X1 U8080 ( .A1(n6514), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n6444) );
  NAND2_X1 U8081 ( .A1(n6475), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n6443) );
  OAI211_X1 U8082 ( .C1(n8467), .C2(n6186), .A(n6444), .B(n6443), .ZN(n6445)
         );
  INV_X1 U8083 ( .A(n6445), .ZN(n6446) );
  NAND2_X1 U8084 ( .A1(n8698), .A2(n8474), .ZN(n6448) );
  NAND2_X1 U8085 ( .A1(n7805), .A2(n8097), .ZN(n6450) );
  NAND2_X1 U8086 ( .A1(n6192), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n6449) );
  INV_X1 U8087 ( .A(n6453), .ZN(n6452) );
  INV_X1 U8088 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n6451) );
  NAND2_X1 U8089 ( .A1(n6452), .A2(n6451), .ZN(n6465) );
  NAND2_X1 U8090 ( .A1(n6453), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n6454) );
  NAND2_X1 U8091 ( .A1(n6465), .A2(n6454), .ZN(n8457) );
  NAND2_X1 U8092 ( .A1(n8457), .A2(n6170), .ZN(n6460) );
  INV_X1 U8093 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n6457) );
  NAND2_X1 U8094 ( .A1(n6514), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n6456) );
  NAND2_X1 U8095 ( .A1(n6475), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n6455) );
  OAI211_X1 U8096 ( .C1(n6457), .C2(n6186), .A(n6456), .B(n6455), .ZN(n6458)
         );
  INV_X1 U8097 ( .A(n6458), .ZN(n6459) );
  NAND2_X1 U8098 ( .A1(n8692), .A2(n8072), .ZN(n6461) );
  NAND2_X1 U8099 ( .A1(n8458), .A2(n8465), .ZN(n6462) );
  NAND2_X1 U8100 ( .A1(n7889), .A2(n8097), .ZN(n6464) );
  NAND2_X1 U8101 ( .A1(n6192), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n6463) );
  NAND2_X1 U8102 ( .A1(n6465), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n6466) );
  NAND2_X1 U8103 ( .A1(n6474), .A2(n6466), .ZN(n8444) );
  NAND2_X1 U8104 ( .A1(n8444), .A2(n6170), .ZN(n6471) );
  INV_X1 U8105 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n8443) );
  NAND2_X1 U8106 ( .A1(n6514), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n6468) );
  NAND2_X1 U8107 ( .A1(n6475), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n6467) );
  OAI211_X1 U8108 ( .C1(n8443), .C2(n6186), .A(n6468), .B(n6467), .ZN(n6469)
         );
  INV_X1 U8109 ( .A(n6469), .ZN(n6470) );
  NAND2_X1 U8110 ( .A1(n7866), .A2(n8097), .ZN(n6473) );
  NAND2_X1 U8111 ( .A1(n6192), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n6472) );
  NAND2_X2 U8112 ( .A1(n6473), .A2(n6472), .ZN(n8272) );
  NAND2_X1 U8113 ( .A1(n7943), .A2(n6170), .ZN(n7356) );
  INV_X1 U8114 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n7945) );
  NAND2_X1 U8115 ( .A1(n6475), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n6477) );
  NAND2_X1 U8116 ( .A1(n6514), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n6476) );
  OAI211_X1 U8117 ( .C1(n6186), .C2(n7945), .A(n6477), .B(n6476), .ZN(n6478)
         );
  INV_X1 U8118 ( .A(n6478), .ZN(n6479) );
  NAND2_X1 U8119 ( .A1(n7356), .A2(n6479), .ZN(n8438) );
  XNOR2_X1 U8120 ( .A(n8272), .B(n8438), .ZN(n8134) );
  XNOR2_X1 U8121 ( .A(n6480), .B(n8134), .ZN(n6526) );
  NAND2_X1 U8122 ( .A1(n8305), .A2(n6527), .ZN(n6562) );
  NAND2_X1 U8123 ( .A1(n6487), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6485) );
  NAND2_X1 U8124 ( .A1(n4414), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6486) );
  MUX2_X1 U8125 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6486), .S(
        P2_IR_REG_20__SCAN_IN), .Z(n6488) );
  INV_X1 U8126 ( .A(n8298), .ZN(n6574) );
  NAND2_X1 U8127 ( .A1(n8151), .A2(n6574), .ZN(n8300) );
  INV_X1 U8128 ( .A(n7300), .ZN(n7179) );
  NAND2_X1 U8129 ( .A1(n6490), .A2(n6489), .ZN(n7197) );
  NAND2_X1 U8130 ( .A1(n7198), .A2(n8143), .ZN(n6803) );
  INV_X1 U8131 ( .A(n8110), .ZN(n6804) );
  NAND2_X1 U8132 ( .A1(n6803), .A2(n6804), .ZN(n6802) );
  NAND2_X1 U8133 ( .A1(n6802), .A2(n8167), .ZN(n7491) );
  INV_X1 U8134 ( .A(n7232), .ZN(n9875) );
  OR2_X1 U8135 ( .A1(n8323), .A2(n9875), .ZN(n8161) );
  INV_X1 U8136 ( .A(n7336), .ZN(n7501) );
  OR2_X1 U8137 ( .A1(n8322), .A2(n7501), .ZN(n7478) );
  NAND2_X1 U8138 ( .A1(n8322), .A2(n7501), .ZN(n8168) );
  AND2_X1 U8139 ( .A1(n7478), .A2(n8163), .ZN(n8174) );
  INV_X1 U8140 ( .A(n7542), .ZN(n9884) );
  NAND2_X1 U8141 ( .A1(n8320), .A2(n9884), .ZN(n8180) );
  AND2_X1 U8142 ( .A1(n8172), .A2(n8180), .ZN(n6491) );
  NAND2_X1 U8143 ( .A1(n7604), .A2(n6491), .ZN(n6494) );
  INV_X1 U8144 ( .A(n8180), .ZN(n6492) );
  OR2_X1 U8145 ( .A1(n6492), .A2(n8179), .ZN(n6493) );
  INV_X1 U8146 ( .A(n8181), .ZN(n6495) );
  AND2_X1 U8147 ( .A1(n9895), .A2(n8317), .ZN(n8182) );
  NAND2_X1 U8148 ( .A1(n7788), .A2(n7776), .ZN(n8195) );
  NAND2_X1 U8149 ( .A1(n7801), .A2(n7852), .ZN(n8197) );
  NAND2_X1 U8150 ( .A1(n7733), .A2(n8119), .ZN(n7747) );
  INV_X1 U8151 ( .A(n8197), .ZN(n8201) );
  NOR2_X1 U8152 ( .A1(n7752), .A2(n8201), .ZN(n6496) );
  NAND2_X1 U8153 ( .A1(n7747), .A2(n6496), .ZN(n7749) );
  NAND2_X1 U8154 ( .A1(n7749), .A2(n8207), .ZN(n8628) );
  INV_X1 U8155 ( .A(n8314), .ZN(n8607) );
  NOR2_X1 U8156 ( .A1(n8623), .A2(n8607), .ZN(n6497) );
  NAND2_X1 U8157 ( .A1(n8623), .A2(n8607), .ZN(n6498) );
  INV_X1 U8158 ( .A(n6499), .ZN(n8219) );
  AOI21_X1 U8159 ( .B1(n8613), .B2(n8217), .A(n8219), .ZN(n8587) );
  NAND2_X1 U8160 ( .A1(n8587), .A2(n8223), .ZN(n8571) );
  AND2_X1 U8161 ( .A1(n8570), .A2(n8225), .ZN(n6501) );
  INV_X1 U8162 ( .A(n8226), .ZN(n6500) );
  NAND2_X1 U8163 ( .A1(n8558), .A2(n8230), .ZN(n6502) );
  AND2_X1 U8164 ( .A1(n8741), .A2(n8563), .ZN(n8231) );
  INV_X1 U8165 ( .A(n8563), .ZN(n6503) );
  NAND2_X1 U8166 ( .A1(n8063), .A2(n6503), .ZN(n8233) );
  AND2_X1 U8167 ( .A1(n8242), .A2(n8531), .ZN(n6504) );
  NAND2_X1 U8168 ( .A1(n6505), .A2(n8245), .ZN(n8518) );
  INV_X1 U8169 ( .A(n8246), .ZN(n6506) );
  NAND2_X1 U8170 ( .A1(n8024), .A2(n8018), .ZN(n8104) );
  NAND2_X1 U8171 ( .A1(n8715), .A2(n8485), .ZN(n8489) );
  NAND2_X1 U8172 ( .A1(n6508), .A2(n8254), .ZN(n8480) );
  NAND2_X1 U8173 ( .A1(n8480), .A2(n8260), .ZN(n6509) );
  NOR2_X1 U8174 ( .A1(n8698), .A2(n8455), .ZN(n8263) );
  NAND2_X1 U8175 ( .A1(n8458), .A2(n8072), .ZN(n8269) );
  INV_X1 U8176 ( .A(n8134), .ZN(n6510) );
  XNOR2_X1 U8177 ( .A(n8091), .B(n6510), .ZN(n7948) );
  OAI211_X1 U8178 ( .C1(n8305), .C2(n8298), .A(n9901), .B(n8421), .ZN(n6511)
         );
  INV_X1 U8179 ( .A(n6511), .ZN(n6512) );
  NAND2_X1 U8180 ( .A1(n8298), .A2(n8421), .ZN(n7174) );
  NAND2_X1 U8181 ( .A1(n7948), .A2(n7666), .ZN(n6524) );
  INV_X1 U8182 ( .A(n6812), .ZN(n8302) );
  INV_X1 U8183 ( .A(n8415), .ZN(n6888) );
  NAND2_X1 U8184 ( .A1(n8302), .A2(n6888), .ZN(n6513) );
  NAND2_X1 U8185 ( .A1(n6521), .A2(n6513), .ZN(n6520) );
  INV_X1 U8186 ( .A(n6520), .ZN(n7166) );
  INV_X1 U8187 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n6517) );
  NAND2_X1 U8188 ( .A1(n6514), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n6516) );
  NAND2_X1 U8189 ( .A1(n6475), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n6515) );
  OAI211_X1 U8190 ( .C1(n6517), .C2(n6186), .A(n6516), .B(n6515), .ZN(n6518)
         );
  INV_X1 U8191 ( .A(n6518), .ZN(n6519) );
  NAND2_X1 U8192 ( .A1(n7356), .A2(n6519), .ZN(n8309) );
  AND2_X1 U8193 ( .A1(n6521), .A2(P2_B_REG_SCAN_IN), .ZN(n6522) );
  NOR2_X1 U8194 ( .A1(n8622), .A2(n6522), .ZN(n8428) );
  AOI22_X1 U8195 ( .A1(n8591), .A2(n8310), .B1(n8309), .B2(n8428), .ZN(n6523)
         );
  NAND2_X1 U8196 ( .A1(n6524), .A2(n6523), .ZN(n6525) );
  INV_X1 U8197 ( .A(n7948), .ZN(n6528) );
  AND2_X1 U8198 ( .A1(n8298), .A2(n6527), .ZN(n7207) );
  INV_X1 U8199 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n6531) );
  XNOR2_X1 U8200 ( .A(n6558), .B(P2_B_REG_SCAN_IN), .ZN(n6537) );
  NAND2_X1 U8201 ( .A1(n6542), .A2(n6537), .ZN(n6545) );
  NAND2_X1 U8202 ( .A1(n6538), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6539) );
  MUX2_X1 U8203 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6539), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n6541) );
  NAND2_X1 U8204 ( .A1(n6542), .A2(n6559), .ZN(n6645) );
  INV_X1 U8205 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n6644) );
  AND2_X1 U8206 ( .A1(n7745), .A2(n6644), .ZN(n6544) );
  NAND2_X1 U8207 ( .A1(n6558), .A2(n6559), .ZN(n7172) );
  NOR2_X1 U8208 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .ZN(
        n6549) );
  NOR4_X1 U8209 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_22__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n6548) );
  NOR4_X1 U8210 ( .A1(P2_D_REG_12__SCAN_IN), .A2(P2_D_REG_25__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_23__SCAN_IN), .ZN(n6547) );
  NOR4_X1 U8211 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_28__SCAN_IN), .A3(
        P2_D_REG_27__SCAN_IN), .A4(P2_D_REG_26__SCAN_IN), .ZN(n6546) );
  NAND4_X1 U8212 ( .A1(n6549), .A2(n6548), .A3(n6547), .A4(n6546), .ZN(n6555)
         );
  NOR4_X1 U8213 ( .A1(P2_D_REG_14__SCAN_IN), .A2(P2_D_REG_13__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n6553) );
  NOR4_X1 U8214 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_9__SCAN_IN), .A3(
        P2_D_REG_17__SCAN_IN), .A4(P2_D_REG_15__SCAN_IN), .ZN(n6552) );
  NOR4_X1 U8215 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n6551) );
  NOR4_X1 U8216 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_19__SCAN_IN), .ZN(n6550) );
  NAND4_X1 U8217 ( .A1(n6553), .A2(n6552), .A3(n6551), .A4(n6550), .ZN(n6554)
         );
  NOR2_X1 U8218 ( .A1(n6555), .A2(n6554), .ZN(n6556) );
  INV_X1 U8219 ( .A(n6570), .ZN(n6557) );
  NAND2_X1 U8220 ( .A1(n7155), .A2(n7162), .ZN(n7185) );
  NAND2_X1 U8221 ( .A1(n8139), .A2(n6574), .ZN(n6563) );
  OR2_X1 U8222 ( .A1(n6563), .A2(n6562), .ZN(n7151) );
  AND2_X1 U8223 ( .A1(n7151), .A2(n7294), .ZN(n6564) );
  OR2_X1 U8224 ( .A1(n7185), .A2(n6564), .ZN(n6567) );
  NAND3_X1 U8225 ( .A1(n7202), .A2(n7200), .A3(n6570), .ZN(n7157) );
  NAND3_X1 U8226 ( .A1(n8284), .A2(n7151), .A3(n9901), .ZN(n7184) );
  NAND2_X1 U8227 ( .A1(n7184), .A2(n8626), .ZN(n7150) );
  NAND2_X1 U8228 ( .A1(n7187), .A2(n7150), .ZN(n6566) );
  INV_X1 U8229 ( .A(n8272), .ZN(n6579) );
  NAND2_X1 U8230 ( .A1(n6568), .A2(n4436), .ZN(P2_U3456) );
  NAND2_X1 U8231 ( .A1(n8289), .A2(n7174), .ZN(n6569) );
  NAND2_X1 U8232 ( .A1(n6587), .A2(n6569), .ZN(n7152) );
  NOR2_X1 U8233 ( .A1(n7152), .A2(n7218), .ZN(n6571) );
  AND2_X1 U8234 ( .A1(n6571), .A2(n6570), .ZN(n6572) );
  NAND3_X1 U8235 ( .A1(n8305), .A2(n6574), .A3(n8421), .ZN(n6575) );
  OAI21_X1 U8236 ( .B1(n7200), .B2(n7161), .A(n7201), .ZN(n6577) );
  INV_X1 U8237 ( .A(n7201), .ZN(n7199) );
  NAND2_X1 U8238 ( .A1(n7202), .A2(n7199), .ZN(n6576) );
  AND2_X1 U8239 ( .A1(n6577), .A2(n6576), .ZN(n6578) );
  NAND2_X1 U8240 ( .A1(n6580), .A2(n4437), .ZN(P2_U3488) );
  INV_X1 U8241 ( .A(n6587), .ZN(n6583) );
  NAND2_X1 U8242 ( .A1(n6583), .A2(n7160), .ZN(n6816) );
  NAND2_X1 U8243 ( .A1(n7160), .A2(n8289), .ZN(n6584) );
  NAND2_X1 U8244 ( .A1(n6816), .A2(n6584), .ZN(n6811) );
  OR2_X1 U8245 ( .A1(n6811), .A2(n6585), .ZN(n6586) );
  NAND2_X1 U8246 ( .A1(n6586), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3150) );
  OAI222_X1 U8247 ( .A1(n9487), .A2(n6588), .B1(n9484), .B2(n6595), .C1(
        P1_U3086), .C2(n8970), .ZN(P1_U3354) );
  INV_X1 U8248 ( .A(n9009), .ZN(n6589) );
  OAI222_X1 U8249 ( .A1(n9487), .A2(n6590), .B1(n9484), .B2(n6597), .C1(
        P1_U3086), .C2(n6589), .ZN(P1_U3352) );
  NOR2_X1 U8250 ( .A1(n4810), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8774) );
  INV_X1 U8251 ( .A(n8774), .ZN(n7741) );
  INV_X1 U8252 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6591) );
  INV_X1 U8253 ( .A(n8338), .ZN(n6895) );
  OAI222_X1 U8254 ( .A1(n7741), .A2(n6591), .B1(n8777), .B2(n6602), .C1(n6895), 
        .C2(P2_U3151), .ZN(P2_U3293) );
  INV_X1 U8255 ( .A(n9017), .ZN(n9596) );
  OAI222_X1 U8256 ( .A1(n9487), .A2(n6592), .B1(n9484), .B2(n6594), .C1(
        P1_U3086), .C2(n9596), .ZN(P1_U3350) );
  INV_X1 U8257 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6593) );
  OAI222_X1 U8258 ( .A1(n6963), .A2(P2_U3151), .B1(n8777), .B2(n6594), .C1(
        n6593), .C2(n7741), .ZN(P2_U3290) );
  OAI222_X1 U8259 ( .A1(n7741), .A2(n4641), .B1(n8777), .B2(n6595), .C1(n6177), 
        .C2(P2_U3151), .ZN(P2_U3294) );
  INV_X1 U8260 ( .A(n6993), .ZN(n7020) );
  INV_X1 U8261 ( .A(n6596), .ZN(n6599) );
  OAI222_X1 U8262 ( .A1(n7020), .A2(P2_U3151), .B1(n8777), .B2(n6599), .C1(
        n4471), .C2(n7741), .ZN(P2_U3289) );
  OAI222_X1 U8263 ( .A1(n7741), .A2(n4996), .B1(n8777), .B2(n6597), .C1(n6915), 
        .C2(P2_U3151), .ZN(P2_U3292) );
  INV_X1 U8264 ( .A(n6899), .ZN(n7138) );
  OAI222_X1 U8265 ( .A1(n7138), .A2(P2_U3151), .B1(n8777), .B2(n6604), .C1(
        n6598), .C2(n7741), .ZN(P2_U3291) );
  INV_X1 U8266 ( .A(n9484), .ZN(n7636) );
  INV_X1 U8267 ( .A(n7636), .ZN(n9481) );
  OAI222_X1 U8268 ( .A1(n9487), .A2(n6600), .B1(n9481), .B2(n6599), .C1(
        P1_U3086), .C2(n9611), .ZN(P1_U3349) );
  INV_X1 U8269 ( .A(n9560), .ZN(n6601) );
  OAI222_X1 U8270 ( .A1(n9487), .A2(n6603), .B1(n9481), .B2(n6602), .C1(
        P1_U3086), .C2(n6601), .ZN(P1_U3353) );
  OAI222_X1 U8271 ( .A1(n9487), .A2(n6605), .B1(n9481), .B2(n6604), .C1(
        P1_U3086), .C2(n9579), .ZN(P1_U3351) );
  OAI222_X1 U8272 ( .A1(n6995), .A2(P2_U3151), .B1(n8777), .B2(n6607), .C1(
        n6606), .C2(n7741), .ZN(P2_U3288) );
  INV_X1 U8273 ( .A(n9022), .ZN(n9511) );
  OAI222_X1 U8274 ( .A1(n9487), .A2(n6608), .B1(n9484), .B2(n6607), .C1(
        P1_U3086), .C2(n9511), .ZN(P1_U3348) );
  INV_X1 U8275 ( .A(n6609), .ZN(n6611) );
  OAI222_X1 U8276 ( .A1(n7072), .A2(P2_U3151), .B1(n8777), .B2(n6611), .C1(
        n6610), .C2(n7741), .ZN(P2_U3287) );
  INV_X1 U8277 ( .A(n9025), .ZN(n9525) );
  OAI222_X1 U8278 ( .A1(n9487), .A2(n6612), .B1(n9481), .B2(n6611), .C1(
        P1_U3086), .C2(n9525), .ZN(P1_U3347) );
  INV_X1 U8279 ( .A(n6613), .ZN(n6618) );
  INV_X1 U8280 ( .A(n9487), .ZN(n6734) );
  AOI22_X1 U8281 ( .A1(n9045), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n6734), .ZN(n6614) );
  OAI21_X1 U8282 ( .B1(n6618), .B2(n9481), .A(n6614), .ZN(P1_U3346) );
  INV_X1 U8283 ( .A(n6615), .ZN(n6620) );
  AOI22_X1 U8284 ( .A1(n9498), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n6734), .ZN(n6616) );
  OAI21_X1 U8285 ( .B1(n6620), .B2(n9481), .A(n6616), .ZN(P1_U3345) );
  OAI222_X1 U8286 ( .A1(P2_U3151), .A2(n7075), .B1(n8777), .B2(n6618), .C1(
        n6617), .C2(n7741), .ZN(P2_U3286) );
  INV_X1 U8287 ( .A(n7118), .ZN(n7103) );
  INV_X1 U8288 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6619) );
  OAI222_X1 U8289 ( .A1(P2_U3151), .A2(n7103), .B1(n8777), .B2(n6620), .C1(
        n6619), .C2(n7741), .ZN(P2_U3285) );
  NAND2_X1 U8290 ( .A1(n6686), .A2(n7638), .ZN(n8965) );
  OR2_X1 U8291 ( .A1(n6699), .A2(n6621), .ZN(n6623) );
  NAND2_X1 U8292 ( .A1(n6623), .A2(n6622), .ZN(n8963) );
  AND2_X1 U8293 ( .A1(n8965), .A2(n8963), .ZN(n9581) );
  NOR2_X1 U8294 ( .A1(n9581), .A2(P1_U3973), .ZN(P1_U3085) );
  INV_X1 U8295 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n6625) );
  NAND2_X1 U8296 ( .A1(n8822), .A2(P1_U3973), .ZN(n6624) );
  OAI21_X1 U8297 ( .B1(P1_U3973), .B2(n6625), .A(n6624), .ZN(P1_U3554) );
  INV_X1 U8298 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n6627) );
  NAND2_X1 U8299 ( .A1(n9088), .A2(P1_U3973), .ZN(n6626) );
  OAI21_X1 U8300 ( .B1(P1_U3973), .B2(n6627), .A(n6626), .ZN(P1_U3585) );
  INV_X1 U8301 ( .A(n6628), .ZN(n6631) );
  INV_X1 U8302 ( .A(n9047), .ZN(n9625) );
  OAI222_X1 U8303 ( .A1(n9487), .A2(n6629), .B1(n9484), .B2(n6631), .C1(
        P1_U3086), .C2(n9625), .ZN(P1_U3344) );
  OAI222_X1 U8304 ( .A1(n4776), .A2(P2_U3151), .B1(n8777), .B2(n6631), .C1(
        n6630), .C2(n7741), .ZN(P2_U3284) );
  INV_X1 U8305 ( .A(n6632), .ZN(n6635) );
  AOI22_X1 U8306 ( .A1(n9629), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n6734), .ZN(n6633) );
  OAI21_X1 U8307 ( .B1(n6635), .B2(n9481), .A(n6633), .ZN(P1_U3343) );
  INV_X1 U8308 ( .A(n7579), .ZN(n7360) );
  INV_X1 U8309 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6634) );
  OAI222_X1 U8310 ( .A1(P2_U3151), .A2(n7360), .B1(n8777), .B2(n6635), .C1(
        n6634), .C2(n7741), .ZN(P2_U3283) );
  INV_X1 U8311 ( .A(n6636), .ZN(n6639) );
  AOI22_X1 U8312 ( .A1(n9644), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n6734), .ZN(n6637) );
  OAI21_X1 U8313 ( .B1(n6639), .B2(n9481), .A(n6637), .ZN(P1_U3342) );
  AOI22_X1 U8314 ( .A1(n8351), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_13__SCAN_IN), .B2(n8774), .ZN(n6638) );
  OAI21_X1 U8315 ( .B1(n6639), .B2(n8777), .A(n6638), .ZN(P2_U3282) );
  INV_X1 U8316 ( .A(n6640), .ZN(n6650) );
  AOI22_X1 U8317 ( .A1(n9659), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n6734), .ZN(n6641) );
  OAI21_X1 U8318 ( .B1(n6650), .B2(n9481), .A(n6641), .ZN(P1_U3341) );
  INV_X1 U8319 ( .A(n7172), .ZN(n6643) );
  AOI22_X1 U8320 ( .A1(n6651), .A2(n6644), .B1(n6647), .B2(n6643), .ZN(
        P2_U3376) );
  INV_X1 U8321 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n6648) );
  INV_X1 U8322 ( .A(n6645), .ZN(n6646) );
  AOI22_X1 U8323 ( .A1(n6651), .A2(n6648), .B1(n6647), .B2(n6646), .ZN(
        P2_U3377) );
  INV_X1 U8324 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6649) );
  OAI222_X1 U8325 ( .A1(P2_U3151), .A2(n9828), .B1(n8777), .B2(n6650), .C1(
        n6649), .C2(n7741), .ZN(P2_U3281) );
  AND2_X1 U8326 ( .A1(n6651), .A2(P2_D_REG_5__SCAN_IN), .ZN(P2_U3260) );
  AND2_X1 U8327 ( .A1(n6651), .A2(P2_D_REG_2__SCAN_IN), .ZN(P2_U3263) );
  AND2_X1 U8328 ( .A1(n6651), .A2(P2_D_REG_20__SCAN_IN), .ZN(P2_U3245) );
  AND2_X1 U8329 ( .A1(n6651), .A2(P2_D_REG_31__SCAN_IN), .ZN(P2_U3234) );
  AND2_X1 U8330 ( .A1(n6651), .A2(P2_D_REG_10__SCAN_IN), .ZN(P2_U3255) );
  AND2_X1 U8331 ( .A1(n6651), .A2(P2_D_REG_6__SCAN_IN), .ZN(P2_U3259) );
  AND2_X1 U8332 ( .A1(n6651), .A2(P2_D_REG_7__SCAN_IN), .ZN(P2_U3258) );
  AND2_X1 U8333 ( .A1(n6651), .A2(P2_D_REG_13__SCAN_IN), .ZN(P2_U3252) );
  AND2_X1 U8334 ( .A1(n6651), .A2(P2_D_REG_26__SCAN_IN), .ZN(P2_U3239) );
  AND2_X1 U8335 ( .A1(n6651), .A2(P2_D_REG_27__SCAN_IN), .ZN(P2_U3238) );
  AND2_X1 U8336 ( .A1(n6651), .A2(P2_D_REG_28__SCAN_IN), .ZN(P2_U3237) );
  AND2_X1 U8337 ( .A1(n6651), .A2(P2_D_REG_29__SCAN_IN), .ZN(P2_U3236) );
  AND2_X1 U8338 ( .A1(n6651), .A2(P2_D_REG_3__SCAN_IN), .ZN(P2_U3262) );
  AND2_X1 U8339 ( .A1(n6651), .A2(P2_D_REG_4__SCAN_IN), .ZN(P2_U3261) );
  AND2_X1 U8340 ( .A1(n6651), .A2(P2_D_REG_17__SCAN_IN), .ZN(P2_U3248) );
  AND2_X1 U8341 ( .A1(n6651), .A2(P2_D_REG_18__SCAN_IN), .ZN(P2_U3247) );
  AND2_X1 U8342 ( .A1(n6651), .A2(P2_D_REG_19__SCAN_IN), .ZN(P2_U3246) );
  AND2_X1 U8343 ( .A1(n6651), .A2(P2_D_REG_8__SCAN_IN), .ZN(P2_U3257) );
  AND2_X1 U8344 ( .A1(n6651), .A2(P2_D_REG_9__SCAN_IN), .ZN(P2_U3256) );
  AND2_X1 U8345 ( .A1(n6651), .A2(P2_D_REG_22__SCAN_IN), .ZN(P2_U3243) );
  AND2_X1 U8346 ( .A1(n6651), .A2(P2_D_REG_11__SCAN_IN), .ZN(P2_U3254) );
  AND2_X1 U8347 ( .A1(n6651), .A2(P2_D_REG_12__SCAN_IN), .ZN(P2_U3253) );
  AND2_X1 U8348 ( .A1(n6651), .A2(P2_D_REG_25__SCAN_IN), .ZN(P2_U3240) );
  AND2_X1 U8349 ( .A1(n6651), .A2(P2_D_REG_14__SCAN_IN), .ZN(P2_U3251) );
  AND2_X1 U8350 ( .A1(n6651), .A2(P2_D_REG_15__SCAN_IN), .ZN(P2_U3250) );
  AND2_X1 U8351 ( .A1(n6651), .A2(P2_D_REG_16__SCAN_IN), .ZN(P2_U3249) );
  AND2_X1 U8352 ( .A1(n6651), .A2(P2_D_REG_24__SCAN_IN), .ZN(P2_U3241) );
  AND2_X1 U8353 ( .A1(n6651), .A2(P2_D_REG_30__SCAN_IN), .ZN(P2_U3235) );
  AND2_X1 U8354 ( .A1(n6651), .A2(P2_D_REG_21__SCAN_IN), .ZN(P2_U3244) );
  AND2_X1 U8355 ( .A1(n6651), .A2(P2_D_REG_23__SCAN_IN), .ZN(P2_U3242) );
  INV_X1 U8356 ( .A(n8392), .ZN(n8355) );
  INV_X1 U8357 ( .A(n6652), .ZN(n6654) );
  INV_X1 U8358 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n6653) );
  OAI222_X1 U8359 ( .A1(n8355), .A2(P2_U3151), .B1(n8777), .B2(n6654), .C1(
        n6653), .C2(n7741), .ZN(P2_U3280) );
  INV_X1 U8360 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n6655) );
  INV_X1 U8361 ( .A(n9684), .ZN(n9049) );
  OAI222_X1 U8362 ( .A1(n9487), .A2(n6655), .B1(n9484), .B2(n6654), .C1(
        P1_U3086), .C2(n9049), .ZN(P1_U3340) );
  XNOR2_X1 U8363 ( .A(n6657), .B(n6656), .ZN(n9563) );
  INV_X1 U8364 ( .A(n8869), .ZN(n6658) );
  NAND2_X1 U8365 ( .A1(n6658), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8824) );
  AOI22_X1 U8366 ( .A1(n8824), .A2(P1_REG3_REG_0__SCAN_IN), .B1(n8945), .B2(
        n9719), .ZN(n6660) );
  NAND2_X1 U8367 ( .A1(n8928), .A2(n9721), .ZN(n6659) );
  OAI211_X1 U8368 ( .C1(n9563), .C2(n8920), .A(n6660), .B(n6659), .ZN(P1_U3232) );
  XOR2_X1 U8369 ( .A(n6661), .B(n6662), .Z(n6666) );
  INV_X1 U8370 ( .A(n8926), .ZN(n8940) );
  NAND2_X1 U8371 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_U3086), .ZN(n8975) );
  OAI21_X1 U8372 ( .B1(n8940), .B2(n6936), .A(n8975), .ZN(n6664) );
  INV_X1 U8373 ( .A(n8927), .ZN(n8941) );
  OAI22_X1 U8374 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(n8941), .B1(n8899), .B2(
        n6833), .ZN(n6663) );
  AOI211_X1 U8375 ( .C1(n6744), .C2(n8928), .A(n6664), .B(n6663), .ZN(n6665)
         );
  OAI21_X1 U8376 ( .B1(n6666), .B2(n8920), .A(n6665), .ZN(P1_U3218) );
  NAND2_X1 U8377 ( .A1(n8326), .A2(n7179), .ZN(n8147) );
  NAND2_X1 U8378 ( .A1(n6667), .A2(n8147), .ZN(n8109) );
  NAND2_X1 U8379 ( .A1(n9908), .A2(n8618), .ZN(n6668) );
  NAND2_X1 U8380 ( .A1(n8109), .A2(n6668), .ZN(n6669) );
  NAND2_X1 U8381 ( .A1(n6183), .A2(n8593), .ZN(n7296) );
  OAI211_X1 U8382 ( .C1(n9901), .C2(n7179), .A(n6669), .B(n7296), .ZN(n7224)
         );
  NAND2_X1 U8383 ( .A1(n9929), .A2(n7224), .ZN(n6670) );
  OAI21_X1 U8384 ( .B1(n9929), .B2(n6163), .A(n6670), .ZN(P2_U3459) );
  INV_X1 U8385 ( .A(n6671), .ZN(n6673) );
  OAI222_X1 U8386 ( .A1(P2_U3151), .A2(n9843), .B1(n8777), .B2(n6673), .C1(
        n6672), .C2(n7741), .ZN(P2_U3279) );
  INV_X1 U8387 ( .A(n9052), .ZN(n9693) );
  OAI222_X1 U8388 ( .A1(n9487), .A2(n6674), .B1(n9484), .B2(n6673), .C1(n9693), 
        .C2(P1_U3086), .ZN(P1_U3339) );
  XOR2_X1 U8389 ( .A(n6675), .B(n6676), .Z(n6679) );
  AOI22_X1 U8390 ( .A1(n8926), .A2(n9719), .B1(n8945), .B2(n8961), .ZN(n6678)
         );
  AOI22_X1 U8391 ( .A1(P1_REG3_REG_2__SCAN_IN), .A2(n8824), .B1(n8928), .B2(
        n6757), .ZN(n6677) );
  OAI211_X1 U8392 ( .C1(n6679), .C2(n8920), .A(n6678), .B(n6677), .ZN(P1_U3237) );
  NAND2_X1 U8393 ( .A1(n8822), .A2(n9721), .ZN(n6930) );
  NAND2_X1 U8394 ( .A1(n6680), .A2(n6959), .ZN(n6681) );
  NAND2_X1 U8395 ( .A1(n6929), .A2(n6681), .ZN(n6754) );
  NAND2_X1 U8396 ( .A1(n6754), .A2(n6753), .ZN(n6756) );
  NAND2_X1 U8397 ( .A1(n6936), .A2(n9726), .ZN(n6682) );
  NAND2_X1 U8398 ( .A1(n6756), .A2(n6682), .ZN(n6741) );
  NAND2_X1 U8399 ( .A1(n6741), .A2(n4802), .ZN(n6740) );
  INV_X1 U8400 ( .A(n8961), .ZN(n6729) );
  NAND2_X1 U8401 ( .A1(n6729), .A2(n6954), .ZN(n6683) );
  NAND2_X1 U8402 ( .A1(n6740), .A2(n6683), .ZN(n6685) );
  INV_X1 U8403 ( .A(n6702), .ZN(n6684) );
  NAND2_X1 U8404 ( .A1(n6685), .A2(n6684), .ZN(n6772) );
  OAI21_X1 U8405 ( .B1(n6685), .B2(n6684), .A(n6772), .ZN(n6863) );
  INV_X1 U8406 ( .A(n6863), .ZN(n6717) );
  INV_X1 U8407 ( .A(n6686), .ZN(n6689) );
  NAND2_X1 U8408 ( .A1(n6689), .A2(n6688), .ZN(n6692) );
  INV_X1 U8409 ( .A(n6690), .ZN(n6691) );
  NAND3_X1 U8410 ( .A1(n6849), .A2(n6693), .A3(n6854), .ZN(n6694) );
  NAND2_X1 U8411 ( .A1(n6695), .A2(n6698), .ZN(n6697) );
  INV_X1 U8412 ( .A(n9720), .ZN(n6696) );
  NAND2_X1 U8413 ( .A1(n6697), .A2(n6696), .ZN(n6700) );
  NOR2_X1 U8414 ( .A1(n6699), .A2(n6698), .ZN(n6821) );
  NAND2_X1 U8415 ( .A1(n7259), .A2(n7243), .ZN(n6701) );
  INV_X1 U8416 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6710) );
  XNOR2_X1 U8417 ( .A(n6703), .B(n6702), .ZN(n6706) );
  NAND2_X1 U8418 ( .A1(n5829), .A2(n9080), .ZN(n6705) );
  OR2_X1 U8419 ( .A1(n7446), .A2(n7383), .ZN(n6704) );
  NAND2_X1 U8420 ( .A1(n6706), .A2(n9765), .ZN(n6708) );
  AOI22_X1 U8421 ( .A1(n9754), .A2(n8961), .B1(n8959), .B2(n9757), .ZN(n6707)
         );
  NAND2_X1 U8422 ( .A1(n6708), .A2(n6707), .ZN(n6861) );
  INV_X1 U8423 ( .A(n6861), .ZN(n6709) );
  MUX2_X1 U8424 ( .A(n6710), .B(n6709), .S(n9265), .Z(n6716) );
  NAND2_X1 U8425 ( .A1(n6959), .A2(n6942), .ZN(n6941) );
  NAND2_X1 U8426 ( .A1(n6760), .A2(n6954), .ZN(n6742) );
  AOI21_X1 U8427 ( .B1(n6742), .B2(n6727), .A(n9792), .ZN(n6711) );
  OR2_X1 U8428 ( .A1(n6742), .A2(n6727), .ZN(n6775) );
  AND2_X1 U8429 ( .A1(n6711), .A2(n6775), .ZN(n6862) );
  INV_X1 U8430 ( .A(n6712), .ZN(n6713) );
  OAI22_X1 U8431 ( .A1(n9273), .A2(n6867), .B1(n6726), .B2(n9242), .ZN(n6714)
         );
  AOI21_X1 U8432 ( .B1(n9284), .B2(n6862), .A(n6714), .ZN(n6715) );
  OAI211_X1 U8433 ( .C1(n6717), .C2(n9306), .A(n6716), .B(n6715), .ZN(P1_U3289) );
  INV_X1 U8434 ( .A(n6718), .ZN(n6721) );
  INV_X1 U8435 ( .A(n9071), .ZN(n9064) );
  OAI222_X1 U8436 ( .A1(n9487), .A2(n6719), .B1(n9484), .B2(n6721), .C1(
        P1_U3086), .C2(n9064), .ZN(P1_U3338) );
  INV_X1 U8437 ( .A(n9847), .ZN(n8367) );
  OAI222_X1 U8438 ( .A1(n8367), .A2(P2_U3151), .B1(n8777), .B2(n6721), .C1(
        n6720), .C2(n7741), .ZN(P2_U3278) );
  INV_X1 U8439 ( .A(n6723), .ZN(n6724) );
  AOI211_X1 U8440 ( .C1(n6725), .C2(n6722), .A(n8920), .B(n6724), .ZN(n6732)
         );
  INV_X1 U8441 ( .A(n8959), .ZN(n6788) );
  OAI22_X1 U8442 ( .A1(n8941), .A2(n6726), .B1(n8899), .B2(n6788), .ZN(n6731)
         );
  NAND2_X1 U8443 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_U3086), .ZN(n9584) );
  NAND2_X1 U8444 ( .A1(n8928), .A2(n6727), .ZN(n6728) );
  OAI211_X1 U8445 ( .C1(n8940), .C2(n6729), .A(n9584), .B(n6728), .ZN(n6730)
         );
  OR3_X1 U8446 ( .A1(n6732), .A2(n6731), .A3(n6730), .ZN(P1_U3230) );
  INV_X1 U8447 ( .A(n6733), .ZN(n6826) );
  AOI22_X1 U8448 ( .A1(n9708), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n6734), .ZN(n6735) );
  OAI21_X1 U8449 ( .B1(n6826), .B2(n9481), .A(n6735), .ZN(P1_U3337) );
  OAI21_X1 U8450 ( .B1(n6738), .B2(n6737), .A(n6736), .ZN(n6739) );
  AOI222_X1 U8451 ( .A1(n9765), .A2(n6739), .B1(n8960), .B2(n9757), .C1(n8962), 
        .C2(n9754), .ZN(n6948) );
  OAI21_X1 U8452 ( .B1(n6741), .B2(n4802), .A(n6740), .ZN(n6946) );
  OAI211_X1 U8453 ( .C1(n6760), .C2(n6954), .A(n6742), .B(n9319), .ZN(n6947)
         );
  INV_X1 U8454 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n8985) );
  OAI22_X1 U8455 ( .A1(n9265), .A2(n8985), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        n9242), .ZN(n6743) );
  AOI21_X1 U8456 ( .B1(n9299), .B2(n6744), .A(n6743), .ZN(n6745) );
  OAI21_X1 U8457 ( .B1(n9302), .B2(n6947), .A(n6745), .ZN(n6746) );
  AOI21_X1 U8458 ( .B1(n6946), .B2(n9212), .A(n6746), .ZN(n6747) );
  OAI21_X1 U8459 ( .B1(n6948), .B2(n9293), .A(n6747), .ZN(P1_U3290) );
  XNOR2_X1 U8460 ( .A(n6749), .B(n6748), .ZN(n6750) );
  NAND2_X1 U8461 ( .A1(n6750), .A2(n9765), .ZN(n6752) );
  AOI22_X1 U8462 ( .A1(n9754), .A2(n9719), .B1(n8961), .B2(n9757), .ZN(n6751)
         );
  AND2_X1 U8463 ( .A1(n6752), .A2(n6751), .ZN(n9729) );
  OR2_X1 U8464 ( .A1(n6754), .A2(n6753), .ZN(n6755) );
  NAND2_X1 U8465 ( .A1(n6756), .A2(n6755), .ZN(n9728) );
  AOI22_X1 U8466 ( .A1(n9293), .A2(P1_REG2_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(n9291), .ZN(n6763) );
  NAND2_X1 U8467 ( .A1(n6941), .A2(n6757), .ZN(n6758) );
  NAND2_X1 U8468 ( .A1(n6758), .A2(n9319), .ZN(n6759) );
  OR2_X1 U8469 ( .A1(n6760), .A2(n6759), .ZN(n9725) );
  INV_X1 U8470 ( .A(n9725), .ZN(n6761) );
  NAND2_X1 U8471 ( .A1(n9284), .A2(n6761), .ZN(n6762) );
  OAI211_X1 U8472 ( .C1(n9726), .C2(n9273), .A(n6763), .B(n6762), .ZN(n6764)
         );
  AOI21_X1 U8473 ( .B1(n9212), .B2(n9728), .A(n6764), .ZN(n6765) );
  OAI21_X1 U8474 ( .B1(n9293), .B2(n9729), .A(n6765), .ZN(P1_U3291) );
  INV_X1 U8475 ( .A(n6766), .ZN(n6773) );
  NAND3_X1 U8476 ( .A1(n6768), .A2(n6767), .A3(n6773), .ZN(n6769) );
  AND2_X1 U8477 ( .A1(n6770), .A2(n6769), .ZN(n6843) );
  NAND2_X1 U8478 ( .A1(n9265), .A2(n9765), .ZN(n9173) );
  NAND2_X1 U8479 ( .A1(n6833), .A2(n6867), .ZN(n6771) );
  OAI21_X1 U8480 ( .B1(n6774), .B2(n6773), .A(n6790), .ZN(n6845) );
  NAND2_X1 U8481 ( .A1(n6845), .A2(n9212), .ZN(n6783) );
  INV_X1 U8482 ( .A(n6775), .ZN(n6776) );
  OR2_X2 U8483 ( .A1(n6775), .A2(n6835), .ZN(n6794) );
  OAI211_X1 U8484 ( .C1(n6776), .C2(n6857), .A(n9319), .B(n6794), .ZN(n6841)
         );
  INV_X1 U8485 ( .A(n6841), .ZN(n6781) );
  AOI22_X1 U8486 ( .A1(n9293), .A2(P1_REG2_REG_5__SCAN_IN), .B1(n6832), .B2(
        n9291), .ZN(n6777) );
  OAI21_X1 U8487 ( .B1(n6857), .B2(n9273), .A(n6777), .ZN(n6780) );
  AND2_X1 U8488 ( .A1(n9265), .A2(n9757), .ZN(n9294) );
  INV_X1 U8489 ( .A(n9294), .ZN(n6778) );
  NAND2_X1 U8490 ( .A1(n9265), .A2(n9754), .ZN(n9297) );
  OAI22_X1 U8491 ( .A1(n6778), .A2(n7263), .B1(n6833), .B2(n9297), .ZN(n6779)
         );
  AOI211_X1 U8492 ( .C1(n9284), .C2(n6781), .A(n6780), .B(n6779), .ZN(n6782)
         );
  OAI211_X1 U8493 ( .C1(n6843), .C2(n9173), .A(n6783), .B(n6782), .ZN(P1_U3288) );
  XNOR2_X1 U8494 ( .A(n6784), .B(n6791), .ZN(n6785) );
  NAND2_X1 U8495 ( .A1(n6785), .A2(n9765), .ZN(n6787) );
  AOI22_X1 U8496 ( .A1(n8957), .A2(n9757), .B1(n9754), .B2(n8959), .ZN(n6786)
         );
  NAND2_X1 U8497 ( .A1(n6787), .A2(n6786), .ZN(n9734) );
  INV_X1 U8498 ( .A(n9734), .ZN(n6801) );
  NAND2_X1 U8499 ( .A1(n6788), .A2(n6857), .ZN(n6789) );
  INV_X1 U8500 ( .A(n6791), .ZN(n6792) );
  OAI21_X1 U8501 ( .B1(n6793), .B2(n6792), .A(n7261), .ZN(n9736) );
  INV_X1 U8502 ( .A(n6794), .ZN(n6796) );
  INV_X1 U8503 ( .A(n7269), .ZN(n6795) );
  OAI211_X1 U8504 ( .C1(n9733), .C2(n6796), .A(n6795), .B(n9319), .ZN(n9732)
         );
  AOI22_X1 U8505 ( .A1(n9293), .A2(P1_REG2_REG_6__SCAN_IN), .B1(n7034), .B2(
        n9291), .ZN(n6798) );
  NAND2_X1 U8506 ( .A1(n9299), .A2(n7037), .ZN(n6797) );
  OAI211_X1 U8507 ( .C1(n9732), .C2(n9302), .A(n6798), .B(n6797), .ZN(n6799)
         );
  AOI21_X1 U8508 ( .B1(n9736), .B2(n9212), .A(n6799), .ZN(n6800) );
  OAI21_X1 U8509 ( .B1(n9293), .B2(n6801), .A(n6800), .ZN(P1_U3287) );
  OAI21_X1 U8510 ( .B1(n6803), .B2(n6804), .A(n6802), .ZN(n7511) );
  INV_X1 U8511 ( .A(n8323), .ZN(n7333) );
  XNOR2_X1 U8512 ( .A(n6805), .B(n6804), .ZN(n6806) );
  OAI222_X1 U8513 ( .A1(n8622), .A2(n7333), .B1(n8620), .B2(n6199), .C1(n8618), 
        .C2(n6806), .ZN(n7508) );
  AOI21_X1 U8514 ( .B1(n9906), .B2(n7511), .A(n7508), .ZN(n7416) );
  AOI22_X1 U8515 ( .A1(n8675), .A2(n7170), .B1(n9927), .B2(
        P2_REG1_REG_3__SCAN_IN), .ZN(n6807) );
  OAI21_X1 U8516 ( .B1(n7416), .B2(n9927), .A(n6807), .ZN(P2_U3462) );
  NOR2_X1 U8517 ( .A1(n4370), .A2(P2_U3151), .ZN(n7806) );
  NAND2_X1 U8518 ( .A1(n7806), .A2(n6812), .ZN(n6808) );
  OR2_X1 U8519 ( .A1(n6811), .A2(n6808), .ZN(n6810) );
  OR2_X1 U8520 ( .A1(n6812), .A2(P2_U3151), .ZN(n8776) );
  OR2_X1 U8521 ( .A1(n6816), .A2(n8776), .ZN(n6809) );
  INV_X1 U8522 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n6890) );
  NAND2_X1 U8523 ( .A1(P2_U3893), .A2(n6812), .ZN(n9858) );
  MUX2_X1 U8524 ( .A(P2_REG2_REG_0__SCAN_IN), .B(P2_REG1_REG_0__SCAN_IN), .S(
        n4370), .Z(n6813) );
  NOR2_X1 U8525 ( .A1(n6813), .A2(n6890), .ZN(n7090) );
  AOI21_X1 U8526 ( .B1(n6890), .B2(n6813), .A(n7090), .ZN(n6814) );
  AOI21_X1 U8527 ( .B1(n6889), .B2(n9858), .A(n6814), .ZN(n6815) );
  AOI21_X1 U8528 ( .B1(P2_REG3_REG_0__SCAN_IN), .B2(P2_U3151), .A(n6815), .ZN(
        n6819) );
  INV_X1 U8529 ( .A(n6816), .ZN(n6817) );
  NAND2_X1 U8530 ( .A1(n9845), .A2(P2_ADDR_REG_0__SCAN_IN), .ZN(n6818) );
  OAI211_X1 U8531 ( .C1(n9844), .C2(n6890), .A(n6819), .B(n6818), .ZN(P2_U3182) );
  INV_X1 U8532 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n9543) );
  INV_X1 U8533 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n6820) );
  OAI22_X1 U8534 ( .A1(n9265), .A2(n9543), .B1(n6820), .B2(n9242), .ZN(n6823)
         );
  NOR4_X1 U8535 ( .A1(n9293), .A2(n9718), .A3(n6821), .A4(n9720), .ZN(n6822)
         );
  AOI211_X1 U8536 ( .C1(n9294), .C2(n9719), .A(n6823), .B(n6822), .ZN(n6825)
         );
  NOR2_X1 U8537 ( .A1(n9302), .A2(n9792), .ZN(n9143) );
  OAI21_X1 U8538 ( .B1(n9143), .B2(n9299), .A(n9721), .ZN(n6824) );
  NAND2_X1 U8539 ( .A1(n6825), .A2(n6824), .ZN(P1_U3293) );
  INV_X1 U8540 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n6827) );
  INV_X1 U8541 ( .A(n8412), .ZN(n8370) );
  OAI222_X1 U8542 ( .A1(n7741), .A2(n6827), .B1(n8777), .B2(n6826), .C1(
        P2_U3151), .C2(n8370), .ZN(P2_U3277) );
  NAND2_X1 U8543 ( .A1(n6829), .A2(n6828), .ZN(n6831) );
  XNOR2_X1 U8544 ( .A(n6831), .B(n6830), .ZN(n6838) );
  AOI22_X1 U8545 ( .A1(n8927), .A2(n6832), .B1(n8945), .B2(n8958), .ZN(n6837)
         );
  NAND2_X1 U8546 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n9598) );
  OAI21_X1 U8547 ( .B1(n8940), .B2(n6833), .A(n9598), .ZN(n6834) );
  AOI21_X1 U8548 ( .B1(n6835), .B2(n8928), .A(n6834), .ZN(n6836) );
  OAI211_X1 U8549 ( .C1(n6838), .C2(n8920), .A(n6837), .B(n6836), .ZN(P1_U3227) );
  AOI22_X1 U8550 ( .A1(n8960), .A2(n9754), .B1(n9757), .B2(n8958), .ZN(n6842)
         );
  OAI211_X1 U8551 ( .C1(n6843), .C2(n9783), .A(n6842), .B(n6841), .ZN(n6844)
         );
  AOI21_X1 U8552 ( .B1(n9794), .B2(n6845), .A(n6844), .ZN(n6860) );
  AND2_X1 U8553 ( .A1(n6847), .A2(n6846), .ZN(n6848) );
  AND2_X1 U8554 ( .A1(n6849), .A2(n6848), .ZN(n6855) );
  INV_X1 U8555 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n6851) );
  OAI22_X1 U8556 ( .A1(n9423), .A2(n6857), .B1(n9813), .B2(n6851), .ZN(n6852)
         );
  INV_X1 U8557 ( .A(n6852), .ZN(n6853) );
  OAI21_X1 U8558 ( .B1(n6860), .B2(n9811), .A(n6853), .ZN(P1_U3527) );
  INV_X1 U8559 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n6856) );
  OAI22_X1 U8560 ( .A1(n9465), .A2(n6857), .B1(n9798), .B2(n6856), .ZN(n6858)
         );
  INV_X1 U8561 ( .A(n6858), .ZN(n6859) );
  OAI21_X1 U8562 ( .B1(n6860), .B2(n9796), .A(n6859), .ZN(P1_U3468) );
  AOI211_X1 U8563 ( .C1(n9794), .C2(n6863), .A(n6862), .B(n6861), .ZN(n6870)
         );
  INV_X1 U8564 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n9012) );
  OAI22_X1 U8565 ( .A1(n9423), .A2(n6867), .B1(n9813), .B2(n9012), .ZN(n6864)
         );
  INV_X1 U8566 ( .A(n6864), .ZN(n6865) );
  OAI21_X1 U8567 ( .B1(n6870), .B2(n9811), .A(n6865), .ZN(P1_U3526) );
  INV_X1 U8568 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n6866) );
  OAI22_X1 U8569 ( .A1(n9465), .A2(n6867), .B1(n9798), .B2(n6866), .ZN(n6868)
         );
  INV_X1 U8570 ( .A(n6868), .ZN(n6869) );
  OAI21_X1 U8571 ( .B1(n6870), .B2(n9796), .A(n6869), .ZN(P1_U3465) );
  MUX2_X1 U8572 ( .A(P2_REG2_REG_5__SCAN_IN), .B(P2_REG1_REG_5__SCAN_IN), .S(
        n8415), .Z(n6964) );
  XNOR2_X1 U8573 ( .A(n6964), .B(n6905), .ZN(n6965) );
  MUX2_X1 U8574 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n4370), .Z(n6876) );
  INV_X1 U8575 ( .A(n6876), .ZN(n6877) );
  MUX2_X1 U8576 ( .A(n7462), .B(n6871), .S(n8415), .Z(n6872) );
  XNOR2_X1 U8577 ( .A(n6872), .B(n6892), .ZN(n7089) );
  OAI22_X1 U8578 ( .A1(n7089), .A2(n7090), .B1(n6892), .B2(n6872), .ZN(n8327)
         );
  MUX2_X1 U8579 ( .A(P2_REG2_REG_2__SCAN_IN), .B(P2_REG1_REG_2__SCAN_IN), .S(
        n8415), .Z(n6873) );
  XNOR2_X1 U8580 ( .A(n6873), .B(n8338), .ZN(n8328) );
  AOI22_X1 U8581 ( .A1(n8327), .A2(n8328), .B1(n6873), .B2(n6895), .ZN(n6925)
         );
  MUX2_X1 U8582 ( .A(P2_REG2_REG_3__SCAN_IN), .B(P2_REG1_REG_3__SCAN_IN), .S(
        n8415), .Z(n6874) );
  XNOR2_X1 U8583 ( .A(n6874), .B(n4488), .ZN(n6924) );
  NAND2_X1 U8584 ( .A1(n6925), .A2(n6924), .ZN(n7143) );
  INV_X1 U8585 ( .A(n6874), .ZN(n6875) );
  NAND2_X1 U8586 ( .A1(n6875), .A2(n4488), .ZN(n7142) );
  XNOR2_X1 U8587 ( .A(n6876), .B(n6899), .ZN(n7145) );
  NAND3_X1 U8588 ( .A1(n7143), .A2(n7142), .A3(n7145), .ZN(n7144) );
  OAI21_X1 U8589 ( .B1(n6899), .B2(n6877), .A(n7144), .ZN(n6966) );
  XOR2_X1 U8590 ( .A(n6965), .B(n6966), .Z(n6912) );
  INV_X1 U8591 ( .A(n6889), .ZN(n6878) );
  NAND2_X1 U8592 ( .A1(n6890), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6879) );
  NAND2_X1 U8593 ( .A1(n6892), .A2(n6879), .ZN(n6880) );
  NAND2_X1 U8594 ( .A1(n6880), .A2(n6881), .ZN(n7083) );
  OR2_X1 U8595 ( .A1(n7083), .A2(n7462), .ZN(n7081) );
  NAND2_X1 U8596 ( .A1(n7081), .A2(n6881), .ZN(n8331) );
  NAND2_X1 U8597 ( .A1(n6895), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6882) );
  MUX2_X1 U8598 ( .A(n6884), .B(P2_REG2_REG_4__SCAN_IN), .S(n6899), .Z(n7131)
         );
  NAND2_X1 U8599 ( .A1(n6883), .A2(n7131), .ZN(n7136) );
  OR2_X1 U8600 ( .A1(n6899), .A2(n6884), .ZN(n6885) );
  NAND2_X1 U8601 ( .A1(n7136), .A2(n6885), .ZN(n6886) );
  OAI21_X1 U8602 ( .B1(n6886), .B2(n6963), .A(n7017), .ZN(n6887) );
  AOI21_X1 U8603 ( .B1(n6887), .B2(n6228), .A(n6990), .ZN(n6908) );
  NAND2_X1 U8604 ( .A1(n6890), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6891) );
  NAND2_X1 U8605 ( .A1(n6892), .A2(n6891), .ZN(n6893) );
  NAND2_X1 U8606 ( .A1(n6893), .A2(n6894), .ZN(n7086) );
  OR2_X1 U8607 ( .A1(n7086), .A2(n6871), .ZN(n7084) );
  NAND2_X1 U8608 ( .A1(n6895), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6896) );
  NAND2_X1 U8609 ( .A1(n7128), .A2(n7126), .ZN(n6897) );
  MUX2_X1 U8610 ( .A(n6898), .B(P2_REG1_REG_4__SCAN_IN), .S(n6899), .Z(n7125)
         );
  NAND2_X1 U8611 ( .A1(n6897), .A2(n7125), .ZN(n7130) );
  INV_X1 U8612 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6898) );
  OR2_X1 U8613 ( .A1(n6899), .A2(n6898), .ZN(n6900) );
  NAND2_X1 U8614 ( .A1(n7130), .A2(n6900), .ZN(n6901) );
  NAND2_X1 U8615 ( .A1(n6901), .A2(n6963), .ZN(n7011) );
  OAI21_X1 U8616 ( .B1(n6901), .B2(n6963), .A(n7011), .ZN(n6902) );
  NAND2_X1 U8617 ( .A1(n6902), .A2(n6231), .ZN(n6903) );
  NAND2_X1 U8618 ( .A1(n6903), .A2(n7009), .ZN(n6904) );
  NAND2_X1 U8619 ( .A1(n8426), .A2(n6904), .ZN(n6907) );
  AND2_X1 U8620 ( .A1(P2_U3151), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n7335) );
  AOI21_X1 U8621 ( .B1(n9846), .B2(n6905), .A(n7335), .ZN(n6906) );
  OAI211_X1 U8622 ( .C1(n9856), .C2(n6908), .A(n6907), .B(n6906), .ZN(n6911)
         );
  INV_X1 U8623 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n6909) );
  NOR2_X1 U8624 ( .A1(n8387), .A2(n6909), .ZN(n6910) );
  AOI211_X1 U8625 ( .C1(n6912), .C2(n8361), .A(n6911), .B(n6910), .ZN(n6913)
         );
  INV_X1 U8626 ( .A(n6913), .ZN(P2_U3187) );
  NOR2_X1 U8627 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10069), .ZN(n7169) );
  INV_X1 U8628 ( .A(n7169), .ZN(n6914) );
  OAI21_X1 U8629 ( .B1(n9844), .B2(n6915), .A(n6914), .ZN(n6923) );
  INV_X1 U8630 ( .A(n7128), .ZN(n6916) );
  AOI21_X1 U8631 ( .B1(n6203), .B2(n6917), .A(n6916), .ZN(n6921) );
  INV_X1 U8632 ( .A(n7134), .ZN(n6918) );
  AOI21_X1 U8633 ( .B1(n6202), .B2(n6919), .A(n6918), .ZN(n6920) );
  OAI22_X1 U8634 ( .A1(n9860), .A2(n6921), .B1(n6920), .B2(n9856), .ZN(n6922)
         );
  AOI211_X1 U8635 ( .C1(n9845), .C2(P2_ADDR_REG_3__SCAN_IN), .A(n6923), .B(
        n6922), .ZN(n6928) );
  OAI21_X1 U8636 ( .B1(n6925), .B2(n6924), .A(n7143), .ZN(n6926) );
  NAND2_X1 U8637 ( .A1(n6926), .A2(n8361), .ZN(n6927) );
  NAND2_X1 U8638 ( .A1(n6928), .A2(n6927), .ZN(P2_U3185) );
  OAI21_X1 U8639 ( .B1(n6931), .B2(n6930), .A(n6929), .ZN(n6932) );
  INV_X1 U8640 ( .A(n6932), .ZN(n7245) );
  OAI21_X1 U8641 ( .B1(n6935), .B2(n6934), .A(n6933), .ZN(n6940) );
  INV_X1 U8642 ( .A(n8822), .ZN(n6937) );
  OAI22_X1 U8643 ( .A1(n6937), .A2(n9776), .B1(n6936), .B2(n9774), .ZN(n6939)
         );
  NOR2_X1 U8644 ( .A1(n7245), .A2(n7259), .ZN(n6938) );
  AOI211_X1 U8645 ( .C1(n9765), .C2(n6940), .A(n6939), .B(n6938), .ZN(n7250)
         );
  OAI211_X1 U8646 ( .C1(n6959), .C2(n6942), .A(n9319), .B(n6941), .ZN(n7244)
         );
  OAI211_X1 U8647 ( .C1(n7245), .C2(n9738), .A(n7250), .B(n7244), .ZN(n6961)
         );
  INV_X1 U8648 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n6943) );
  OAI22_X1 U8649 ( .A1(n9423), .A2(n6959), .B1(n9813), .B2(n6943), .ZN(n6944)
         );
  AOI21_X1 U8650 ( .B1(n6961), .B2(n9813), .A(n6944), .ZN(n6945) );
  INV_X1 U8651 ( .A(n6945), .ZN(P1_U3523) );
  INV_X1 U8652 ( .A(n6946), .ZN(n6949) );
  OAI211_X1 U8653 ( .C1(n9760), .C2(n6949), .A(n6948), .B(n6947), .ZN(n6956)
         );
  INV_X1 U8654 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6950) );
  OAI22_X1 U8655 ( .A1(n9423), .A2(n6954), .B1(n9813), .B2(n6950), .ZN(n6951)
         );
  AOI21_X1 U8656 ( .B1(n6956), .B2(n9813), .A(n6951), .ZN(n6952) );
  INV_X1 U8657 ( .A(n6952), .ZN(P1_U3525) );
  INV_X1 U8658 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n6953) );
  OAI22_X1 U8659 ( .A1(n9465), .A2(n6954), .B1(n9798), .B2(n6953), .ZN(n6955)
         );
  AOI21_X1 U8660 ( .B1(n6956), .B2(n9798), .A(n6955), .ZN(n6957) );
  INV_X1 U8661 ( .A(n6957), .ZN(P1_U3462) );
  INV_X1 U8662 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n6958) );
  OAI22_X1 U8663 ( .A1(n9465), .A2(n6959), .B1(n9798), .B2(n6958), .ZN(n6960)
         );
  AOI21_X1 U8664 ( .B1(n6961), .B2(n9798), .A(n6960), .ZN(n6962) );
  INV_X1 U8665 ( .A(n6962), .ZN(P1_U3456) );
  AOI22_X1 U8666 ( .A1(n6966), .A2(n6965), .B1(n6964), .B2(n6963), .ZN(n7025)
         );
  MUX2_X1 U8667 ( .A(P2_REG2_REG_6__SCAN_IN), .B(P2_REG1_REG_6__SCAN_IN), .S(
        n4370), .Z(n6967) );
  NOR2_X1 U8668 ( .A1(n6967), .A2(n7020), .ZN(n6968) );
  AOI21_X1 U8669 ( .B1(n6967), .B2(n7020), .A(n6968), .ZN(n7024) );
  NAND2_X1 U8670 ( .A1(n7025), .A2(n7024), .ZN(n7043) );
  INV_X1 U8671 ( .A(n6968), .ZN(n7042) );
  MUX2_X1 U8672 ( .A(n6970), .B(n6969), .S(n8415), .Z(n6971) );
  NAND2_X1 U8673 ( .A1(n6971), .A2(n7051), .ZN(n6974) );
  INV_X1 U8674 ( .A(n6971), .ZN(n6972) );
  NAND2_X1 U8675 ( .A1(n6972), .A2(n6995), .ZN(n6973) );
  NAND2_X1 U8676 ( .A1(n6974), .A2(n6973), .ZN(n7041) );
  AOI21_X1 U8677 ( .B1(n7043), .B2(n7042), .A(n7041), .ZN(n7045) );
  INV_X1 U8678 ( .A(n6974), .ZN(n6979) );
  MUX2_X1 U8679 ( .A(n6988), .B(n9922), .S(n8415), .Z(n6975) );
  NAND2_X1 U8680 ( .A1(n6975), .A2(n6989), .ZN(n7068) );
  INV_X1 U8681 ( .A(n6975), .ZN(n6976) );
  NAND2_X1 U8682 ( .A1(n6976), .A2(n7072), .ZN(n6977) );
  AND2_X1 U8683 ( .A1(n7068), .A2(n6977), .ZN(n6978) );
  OAI21_X1 U8684 ( .B1(n7045), .B2(n6979), .A(n6978), .ZN(n7069) );
  INV_X1 U8685 ( .A(n7069), .ZN(n6981) );
  NOR3_X1 U8686 ( .A1(n7045), .A2(n6979), .A3(n6978), .ZN(n6980) );
  OAI21_X1 U8687 ( .B1(n6981), .B2(n6980), .A(n8361), .ZN(n7007) );
  NOR2_X1 U8688 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n4458), .ZN(n7599) );
  INV_X1 U8689 ( .A(n7599), .ZN(n6982) );
  OAI21_X1 U8690 ( .B1(n9844), .B2(n7072), .A(n6982), .ZN(n7005) );
  NAND2_X1 U8691 ( .A1(n7011), .A2(n7009), .ZN(n6983) );
  XNOR2_X1 U8692 ( .A(n6993), .B(P2_REG1_REG_6__SCAN_IN), .ZN(n7008) );
  NAND2_X1 U8693 ( .A1(n6983), .A2(n7008), .ZN(n7013) );
  OR2_X1 U8694 ( .A1(n6993), .A2(n9919), .ZN(n6984) );
  NAND2_X1 U8695 ( .A1(n7013), .A2(n6984), .ZN(n6985) );
  NOR2_X1 U8696 ( .A1(n6969), .A2(n7048), .ZN(n7050) );
  NAND2_X1 U8697 ( .A1(n7072), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n7058) );
  OAI21_X1 U8698 ( .B1(n7072), .B2(P2_REG1_REG_8__SCAN_IN), .A(n7058), .ZN(
        n6986) );
  AOI21_X1 U8699 ( .B1(n6987), .B2(n6986), .A(n7060), .ZN(n7003) );
  XNOR2_X1 U8700 ( .A(n6989), .B(n6988), .ZN(n6998) );
  INV_X1 U8701 ( .A(n6998), .ZN(n6997) );
  INV_X1 U8702 ( .A(n6990), .ZN(n7015) );
  NAND2_X1 U8703 ( .A1(n7017), .A2(n7015), .ZN(n6991) );
  XNOR2_X1 U8704 ( .A(n6993), .B(P2_REG2_REG_6__SCAN_IN), .ZN(n7014) );
  NAND2_X1 U8705 ( .A1(n6991), .A2(n7014), .ZN(n7019) );
  OR2_X1 U8706 ( .A1(n6993), .A2(n6992), .ZN(n6994) );
  NOR2_X1 U8707 ( .A1(n6997), .A2(n7046), .ZN(n7001) );
  AOI21_X1 U8708 ( .B1(n7000), .B2(n6999), .A(n6998), .ZN(n7071) );
  AOI21_X1 U8709 ( .B1(n7001), .B2(n7000), .A(n7071), .ZN(n7002) );
  OAI22_X1 U8710 ( .A1(n9860), .A2(n7003), .B1(n7002), .B2(n9856), .ZN(n7004)
         );
  AOI211_X1 U8711 ( .C1(n9845), .C2(P2_ADDR_REG_8__SCAN_IN), .A(n7005), .B(
        n7004), .ZN(n7006) );
  NAND2_X1 U8712 ( .A1(n7007), .A2(n7006), .ZN(P2_U3190) );
  INV_X1 U8713 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n9944) );
  INV_X1 U8714 ( .A(n7008), .ZN(n7010) );
  NAND3_X1 U8715 ( .A1(n7011), .A2(n7010), .A3(n7009), .ZN(n7012) );
  AOI21_X1 U8716 ( .B1(n7013), .B2(n7012), .A(n9860), .ZN(n7023) );
  INV_X1 U8717 ( .A(n7014), .ZN(n7016) );
  NAND3_X1 U8718 ( .A1(n7017), .A2(n7016), .A3(n7015), .ZN(n7018) );
  AOI21_X1 U8719 ( .B1(n7019), .B2(n7018), .A(n9856), .ZN(n7022) );
  NOR2_X1 U8720 ( .A1(n9844), .A2(n7020), .ZN(n7021) );
  NOR2_X1 U8721 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n4455), .ZN(n7395) );
  NOR4_X1 U8722 ( .A1(n7023), .A2(n7022), .A3(n7021), .A4(n7395), .ZN(n7028)
         );
  OAI21_X1 U8723 ( .B1(n7025), .B2(n7024), .A(n7043), .ZN(n7026) );
  NAND2_X1 U8724 ( .A1(n7026), .A2(n8361), .ZN(n7027) );
  OAI211_X1 U8725 ( .C1(n9944), .C2(n8387), .A(n7028), .B(n7027), .ZN(P2_U3188) );
  NAND2_X1 U8726 ( .A1(n4833), .A2(n7032), .ZN(n7033) );
  XNOR2_X1 U8727 ( .A(n7030), .B(n7033), .ZN(n7040) );
  AOI22_X1 U8728 ( .A1(n7034), .A2(n8927), .B1(n8926), .B2(n8959), .ZN(n7039)
         );
  NAND2_X1 U8729 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n9613) );
  INV_X1 U8730 ( .A(n9613), .ZN(n7036) );
  NOR2_X1 U8731 ( .A1(n8899), .A2(n7311), .ZN(n7035) );
  AOI211_X1 U8732 ( .C1(n7037), .C2(n8928), .A(n7036), .B(n7035), .ZN(n7038)
         );
  OAI211_X1 U8733 ( .C1(n7040), .C2(n8920), .A(n7039), .B(n7038), .ZN(P1_U3239) );
  INV_X1 U8734 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n9948) );
  AND3_X1 U8735 ( .A1(n7043), .A2(n7042), .A3(n7041), .ZN(n7044) );
  OAI21_X1 U8736 ( .B1(n7045), .B2(n7044), .A(n8361), .ZN(n7057) );
  AOI21_X1 U8737 ( .B1(n7047), .B2(n6970), .A(n7046), .ZN(n7054) );
  AND2_X1 U8738 ( .A1(n7048), .A2(n6969), .ZN(n7049) );
  OAI21_X1 U8739 ( .B1(n7050), .B2(n7049), .A(n8426), .ZN(n7053) );
  NOR2_X1 U8740 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6122), .ZN(n7541) );
  AOI21_X1 U8741 ( .B1(n9846), .B2(n7051), .A(n7541), .ZN(n7052) );
  OAI211_X1 U8742 ( .C1(n7054), .C2(n9856), .A(n7053), .B(n7052), .ZN(n7055)
         );
  INV_X1 U8743 ( .A(n7055), .ZN(n7056) );
  OAI211_X1 U8744 ( .C1(n9948), .C2(n8387), .A(n7057), .B(n7056), .ZN(P2_U3189) );
  INV_X1 U8745 ( .A(n7058), .ZN(n7059) );
  AOI21_X1 U8746 ( .B1(n7062), .B2(n7061), .A(n7096), .ZN(n7080) );
  MUX2_X1 U8747 ( .A(n7063), .B(n7062), .S(n4370), .Z(n7064) );
  NAND2_X1 U8748 ( .A1(n7064), .A2(n7112), .ZN(n7101) );
  INV_X1 U8749 ( .A(n7064), .ZN(n7065) );
  NAND2_X1 U8750 ( .A1(n7065), .A2(n7075), .ZN(n7066) );
  NAND2_X1 U8751 ( .A1(n7101), .A2(n7066), .ZN(n7067) );
  AOI21_X1 U8752 ( .B1(n7069), .B2(n7068), .A(n7067), .ZN(n7108) );
  AND3_X1 U8753 ( .A1(n7069), .A2(n7068), .A3(n7067), .ZN(n7070) );
  OAI21_X1 U8754 ( .B1(n7108), .B2(n7070), .A(n8361), .ZN(n7079) );
  AOI21_X1 U8755 ( .B1(n7063), .B2(n7073), .A(n7113), .ZN(n7074) );
  NOR2_X1 U8756 ( .A1(n7074), .A2(n9856), .ZN(n7077) );
  NOR2_X1 U8757 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6124), .ZN(n7660) );
  INV_X1 U8758 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n9954) );
  OAI22_X1 U8759 ( .A1(n9844), .A2(n7075), .B1(n8387), .B2(n9954), .ZN(n7076)
         );
  NOR3_X1 U8760 ( .A1(n7077), .A2(n7660), .A3(n7076), .ZN(n7078) );
  OAI211_X1 U8761 ( .C1(n7080), .C2(n9860), .A(n7079), .B(n7078), .ZN(P2_U3191) );
  INV_X1 U8762 ( .A(n7081), .ZN(n7082) );
  AOI21_X1 U8763 ( .B1(n7462), .B2(n7083), .A(n7082), .ZN(n7094) );
  INV_X1 U8764 ( .A(n7084), .ZN(n7085) );
  AOI21_X1 U8765 ( .B1(n6871), .B2(n7086), .A(n7085), .ZN(n7087) );
  OAI22_X1 U8766 ( .A1(n9860), .A2(n7087), .B1(n9844), .B2(n6177), .ZN(n7088)
         );
  AOI21_X1 U8767 ( .B1(n9845), .B2(P2_ADDR_REG_1__SCAN_IN), .A(n7088), .ZN(
        n7093) );
  XOR2_X1 U8768 ( .A(n7090), .B(n7089), .Z(n7091) );
  INV_X1 U8769 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n10105) );
  AOI22_X1 U8770 ( .A1(n8361), .A2(n7091), .B1(P2_U3151), .B2(
        P2_REG3_REG_1__SCAN_IN), .ZN(n7092) );
  OAI211_X1 U8771 ( .C1(n7094), .C2(n9856), .A(n7093), .B(n7092), .ZN(P2_U3183) );
  OR2_X1 U8772 ( .A1(n7118), .A2(n9924), .ZN(n7276) );
  NAND2_X1 U8773 ( .A1(n7118), .A2(n9924), .ZN(n7097) );
  NAND2_X1 U8774 ( .A1(n7276), .A2(n7097), .ZN(n7099) );
  INV_X1 U8775 ( .A(n7277), .ZN(n7098) );
  AOI21_X1 U8776 ( .B1(n7100), .B2(n7099), .A(n7098), .ZN(n7124) );
  INV_X1 U8777 ( .A(n7101), .ZN(n7107) );
  MUX2_X1 U8778 ( .A(n7115), .B(n9924), .S(n8415), .Z(n7102) );
  NAND2_X1 U8779 ( .A1(n7102), .A2(n7118), .ZN(n7285) );
  INV_X1 U8780 ( .A(n7102), .ZN(n7104) );
  NAND2_X1 U8781 ( .A1(n7104), .A2(n7103), .ZN(n7105) );
  AND2_X1 U8782 ( .A1(n7285), .A2(n7105), .ZN(n7106) );
  OAI21_X1 U8783 ( .B1(n7108), .B2(n7107), .A(n7106), .ZN(n7286) );
  INV_X1 U8784 ( .A(n7286), .ZN(n7110) );
  NOR3_X1 U8785 ( .A1(n7108), .A2(n7107), .A3(n7106), .ZN(n7109) );
  OAI21_X1 U8786 ( .B1(n7110), .B2(n7109), .A(n8361), .ZN(n7123) );
  NOR2_X1 U8787 ( .A1(n7112), .A2(n7111), .ZN(n7114) );
  OR2_X1 U8788 ( .A1(n7118), .A2(n7115), .ZN(n7279) );
  NAND2_X1 U8789 ( .A1(n7118), .A2(n7115), .ZN(n7116) );
  OAI21_X1 U8790 ( .B1(n4609), .B2(n4450), .A(n7280), .ZN(n7121) );
  INV_X1 U8791 ( .A(n9856), .ZN(n8337) );
  INV_X1 U8792 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n9958) );
  INV_X1 U8793 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n7117) );
  NOR2_X1 U8794 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7117), .ZN(n7775) );
  AOI21_X1 U8795 ( .B1(n9846), .B2(n7118), .A(n7775), .ZN(n7119) );
  OAI21_X1 U8796 ( .B1(n8387), .B2(n9958), .A(n7119), .ZN(n7120) );
  AOI21_X1 U8797 ( .B1(n7121), .B2(n8337), .A(n7120), .ZN(n7122) );
  OAI211_X1 U8798 ( .C1(n7124), .C2(n9860), .A(n7123), .B(n7122), .ZN(P2_U3192) );
  INV_X1 U8799 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n7149) );
  INV_X1 U8800 ( .A(n7125), .ZN(n7127) );
  NAND3_X1 U8801 ( .A1(n7128), .A2(n7127), .A3(n7126), .ZN(n7129) );
  AOI21_X1 U8802 ( .B1(n7130), .B2(n7129), .A(n9860), .ZN(n7141) );
  INV_X1 U8803 ( .A(n7131), .ZN(n7133) );
  NAND3_X1 U8804 ( .A1(n7134), .A2(n7133), .A3(n7132), .ZN(n7135) );
  AOI21_X1 U8805 ( .B1(n7136), .B2(n7135), .A(n9856), .ZN(n7140) );
  NOR2_X1 U8806 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10128), .ZN(n7228) );
  INV_X1 U8807 ( .A(n7228), .ZN(n7137) );
  OAI21_X1 U8808 ( .B1(n9844), .B2(n7138), .A(n7137), .ZN(n7139) );
  NOR3_X1 U8809 ( .A1(n7141), .A2(n7140), .A3(n7139), .ZN(n7148) );
  AND2_X1 U8810 ( .A1(n7143), .A2(n7142), .ZN(n7146) );
  OAI211_X1 U8811 ( .C1(n7146), .C2(n7145), .A(n8361), .B(n7144), .ZN(n7147)
         );
  OAI211_X1 U8812 ( .C1(n8387), .C2(n7149), .A(n7148), .B(n7147), .ZN(P2_U3186) );
  INV_X1 U8813 ( .A(n7150), .ZN(n7154) );
  INV_X1 U8814 ( .A(n7151), .ZN(n7186) );
  AOI21_X1 U8815 ( .B1(n7157), .B2(n7186), .A(n7152), .ZN(n7153) );
  OAI21_X1 U8816 ( .B1(n7155), .B2(n7154), .A(n7153), .ZN(n7156) );
  NAND2_X1 U8817 ( .A1(n7156), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7159) );
  INV_X1 U8818 ( .A(n7294), .ZN(n7164) );
  AND2_X1 U8819 ( .A1(n7162), .A2(n7164), .ZN(n8303) );
  NAND2_X1 U8820 ( .A1(n7157), .A2(n8303), .ZN(n7158) );
  NAND2_X1 U8821 ( .A1(n7159), .A2(n7158), .ZN(n7219) );
  OR2_X1 U8822 ( .A1(n7160), .A2(P2_U3151), .ZN(n8307) );
  INV_X1 U8823 ( .A(n8307), .ZN(n7633) );
  OR2_X1 U8824 ( .A1(n7185), .A2(n9901), .ZN(n7163) );
  AND2_X1 U8825 ( .A1(n7187), .A2(n7164), .ZN(n7165) );
  INV_X1 U8826 ( .A(n7165), .ZN(n7167) );
  OAI22_X1 U8827 ( .A1(n8031), .A2(n6199), .B1(n7333), .B2(n8081), .ZN(n7168)
         );
  AOI211_X1 U8828 ( .C1(n7170), .C2(n8089), .A(n7169), .B(n7168), .ZN(n7196)
         );
  XNOR2_X1 U8829 ( .A(n8151), .B(n8298), .ZN(n7171) );
  NAND2_X4 U8830 ( .A1(n7175), .A2(n7174), .ZN(n7183) );
  INV_X1 U8831 ( .A(n7177), .ZN(n7176) );
  NAND2_X1 U8832 ( .A1(n7176), .A2(n6183), .ZN(n7178) );
  NAND2_X1 U8833 ( .A1(n7177), .A2(n6182), .ZN(n7180) );
  XNOR2_X1 U8834 ( .A(n7183), .B(n6198), .ZN(n7181) );
  XNOR2_X1 U8835 ( .A(n7181), .B(n8325), .ZN(n7342) );
  NAND2_X1 U8836 ( .A1(n7341), .A2(n7342), .ZN(n7340) );
  NAND2_X1 U8837 ( .A1(n7181), .A2(n6199), .ZN(n7182) );
  NAND2_X1 U8838 ( .A1(n7340), .A2(n7182), .ZN(n7190) );
  XNOR2_X1 U8839 ( .A(n7183), .B(n7507), .ZN(n7229) );
  XNOR2_X1 U8840 ( .A(n7229), .B(n8324), .ZN(n7191) );
  OR2_X1 U8841 ( .A1(n7185), .A2(n7184), .ZN(n7189) );
  NAND2_X1 U8842 ( .A1(n7187), .A2(n7186), .ZN(n7188) );
  AOI21_X1 U8843 ( .B1(n7190), .B2(n7191), .A(n8084), .ZN(n7194) );
  INV_X1 U8844 ( .A(n7190), .ZN(n7193) );
  NAND2_X1 U8845 ( .A1(n7193), .A2(n7192), .ZN(n7231) );
  NAND2_X1 U8846 ( .A1(n7194), .A2(n7231), .ZN(n7195) );
  OAI211_X1 U8847 ( .C1(P2_REG3_REG_3__SCAN_IN), .C2(n8061), .A(n7196), .B(
        n7195), .ZN(P2_U3158) );
  INV_X1 U8848 ( .A(n7210), .ZN(n9871) );
  NAND2_X1 U8849 ( .A1(n7200), .A2(n7199), .ZN(n7204) );
  NAND2_X1 U8850 ( .A1(n7202), .A2(n7201), .ZN(n7203) );
  NAND2_X1 U8851 ( .A1(n7207), .A2(n8151), .ZN(n7455) );
  NOR2_X1 U8852 ( .A1(n8582), .A2(n7455), .ZN(n7947) );
  INV_X1 U8853 ( .A(n7947), .ZN(n7217) );
  XNOR2_X1 U8854 ( .A(n7208), .B(n8152), .ZN(n7212) );
  INV_X1 U8855 ( .A(n8324), .ZN(n7496) );
  OAI22_X1 U8856 ( .A1(n6182), .A2(n8620), .B1(n7496), .B2(n8622), .ZN(n7209)
         );
  AOI21_X1 U8857 ( .B1(n7210), .B2(n7666), .A(n7209), .ZN(n7211) );
  OAI21_X1 U8858 ( .B1(n8618), .B2(n7212), .A(n7211), .ZN(n9873) );
  OAI22_X1 U8859 ( .A1(n8624), .A2(n7346), .B1(n9869), .B2(n8626), .ZN(n7213)
         );
  NOR2_X1 U8860 ( .A1(n9873), .A2(n7213), .ZN(n7215) );
  MUX2_X1 U8861 ( .A(n7215), .B(n7214), .S(n8582), .Z(n7216) );
  OAI21_X1 U8862 ( .B1(n9871), .B2(n7217), .A(n7216), .ZN(P2_U3231) );
  NOR2_X1 U8863 ( .A1(n7219), .A2(n7218), .ZN(n7401) );
  AOI22_X1 U8864 ( .A1(n8005), .A2(n8109), .B1(n7300), .B2(n8089), .ZN(n7221)
         );
  NAND2_X1 U8865 ( .A1(n8009), .A2(n6183), .ZN(n7220) );
  OAI211_X1 U8866 ( .C1(n7401), .C2(n7297), .A(n7221), .B(n7220), .ZN(P2_U3172) );
  INV_X1 U8867 ( .A(n7222), .ZN(n7864) );
  OAI222_X1 U8868 ( .A1(P2_U3151), .A2(n8421), .B1(n8777), .B2(n7864), .C1(
        n7223), .C2(n7741), .ZN(P2_U3276) );
  NAND2_X1 U8869 ( .A1(n9914), .A2(n7224), .ZN(n7225) );
  OAI21_X1 U8870 ( .B1(n9914), .B2(n7226), .A(n7225), .ZN(P2_U3390) );
  INV_X1 U8871 ( .A(n8322), .ZN(n7495) );
  OAI22_X1 U8872 ( .A1(n8031), .A2(n7496), .B1(n7495), .B2(n8081), .ZN(n7227)
         );
  AOI211_X1 U8873 ( .C1(n7232), .C2(n8089), .A(n7228), .B(n7227), .ZN(n7240)
         );
  NAND2_X1 U8874 ( .A1(n7229), .A2(n8324), .ZN(n7230) );
  XNOR2_X1 U8875 ( .A(n7183), .B(n7232), .ZN(n7233) );
  NAND2_X1 U8876 ( .A1(n7233), .A2(n7333), .ZN(n7328) );
  INV_X1 U8877 ( .A(n7233), .ZN(n7234) );
  NAND2_X1 U8878 ( .A1(n7234), .A2(n8323), .ZN(n7235) );
  AND2_X1 U8879 ( .A1(n7328), .A2(n7235), .ZN(n7236) );
  OAI21_X1 U8880 ( .B1(n7237), .B2(n7236), .A(n7329), .ZN(n7238) );
  NAND2_X1 U8881 ( .A1(n7238), .A2(n8005), .ZN(n7239) );
  OAI211_X1 U8882 ( .C1(n7492), .C2(n8061), .A(n7240), .B(n7239), .ZN(P2_U3170) );
  INV_X1 U8883 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n7242) );
  INV_X1 U8884 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n7241) );
  OAI22_X1 U8885 ( .A1(n9265), .A2(n7242), .B1(n7241), .B2(n9242), .ZN(n7248)
         );
  NOR2_X1 U8886 ( .A1(n9293), .A2(n7243), .ZN(n7321) );
  INV_X1 U8887 ( .A(n7321), .ZN(n7246) );
  OAI22_X1 U8888 ( .A1(n7246), .A2(n7245), .B1(n9302), .B2(n7244), .ZN(n7247)
         );
  AOI211_X1 U8889 ( .C1(n9299), .C2(n8823), .A(n7248), .B(n7247), .ZN(n7249)
         );
  OAI21_X1 U8890 ( .B1(n7250), .B2(n9293), .A(n7249), .ZN(P1_U3292) );
  XOR2_X1 U8891 ( .A(n7253), .B(n7252), .Z(n7254) );
  XNOR2_X1 U8892 ( .A(n7251), .B(n7254), .ZN(n7258) );
  AOI22_X1 U8893 ( .A1(n7270), .A2(n8927), .B1(n8945), .B2(n9746), .ZN(n7255)
         );
  NAND2_X1 U8894 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3086), .ZN(n9513) );
  OAI211_X1 U8895 ( .C1(n7263), .C2(n8940), .A(n7255), .B(n9513), .ZN(n7256)
         );
  AOI21_X1 U8896 ( .B1(n7271), .B2(n8928), .A(n7256), .ZN(n7257) );
  OAI21_X1 U8897 ( .B1(n7258), .B2(n8920), .A(n7257), .ZN(P1_U3213) );
  INV_X1 U8898 ( .A(n7259), .ZN(n7304) );
  NAND2_X1 U8899 ( .A1(n7263), .A2(n9733), .ZN(n7260) );
  NAND2_X1 U8900 ( .A1(n7261), .A2(n7260), .ZN(n7262) );
  OAI21_X1 U8901 ( .B1(n7262), .B2(n7305), .A(n7303), .ZN(n7417) );
  OAI22_X1 U8902 ( .A1(n7263), .A2(n9776), .B1(n7439), .B2(n9774), .ZN(n7268)
         );
  NAND2_X1 U8903 ( .A1(n7265), .A2(n7264), .ZN(n7306) );
  XOR2_X1 U8904 ( .A(n7305), .B(n7306), .Z(n7266) );
  NOR2_X1 U8905 ( .A1(n7266), .A2(n9783), .ZN(n7267) );
  AOI211_X1 U8906 ( .C1(n7304), .C2(n7417), .A(n7268), .B(n7267), .ZN(n7419)
         );
  OAI211_X1 U8907 ( .C1(n7269), .C2(n7425), .A(n7316), .B(n9319), .ZN(n7418)
         );
  AOI22_X1 U8908 ( .A1(n9293), .A2(P1_REG2_REG_7__SCAN_IN), .B1(n7270), .B2(
        n9291), .ZN(n7273) );
  NAND2_X1 U8909 ( .A1(n9299), .A2(n7271), .ZN(n7272) );
  OAI211_X1 U8910 ( .C1(n7418), .C2(n9302), .A(n7273), .B(n7272), .ZN(n7274)
         );
  AOI21_X1 U8911 ( .B1(n7417), .B2(n7321), .A(n7274), .ZN(n7275) );
  OAI21_X1 U8912 ( .B1(n7419), .B2(n9293), .A(n7275), .ZN(P1_U3286) );
  AOI21_X1 U8913 ( .B1(n6306), .B2(n7278), .A(n7365), .ZN(n7292) );
  XNOR2_X1 U8914 ( .A(n7370), .B(n7369), .ZN(n7281) );
  AOI21_X1 U8915 ( .B1(n6309), .B2(n7281), .A(n7371), .ZN(n7282) );
  NOR2_X1 U8916 ( .A1(n7282), .A2(n9856), .ZN(n7284) );
  INV_X1 U8917 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n10072) );
  NOR2_X1 U8918 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10072), .ZN(n7797) );
  INV_X1 U8919 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n9962) );
  OAI22_X1 U8920 ( .A1(n9844), .A2(n4776), .B1(n8387), .B2(n9962), .ZN(n7283)
         );
  NOR3_X1 U8921 ( .A1(n7284), .A2(n7797), .A3(n7283), .ZN(n7291) );
  NAND2_X1 U8922 ( .A1(n7286), .A2(n7285), .ZN(n7288) );
  MUX2_X1 U8923 ( .A(P2_REG2_REG_11__SCAN_IN), .B(P2_REG1_REG_11__SCAN_IN), 
        .S(n4370), .Z(n7359) );
  XNOR2_X1 U8924 ( .A(n7359), .B(n7370), .ZN(n7287) );
  NAND2_X1 U8925 ( .A1(n7288), .A2(n7287), .ZN(n7358) );
  OAI21_X1 U8926 ( .B1(n7288), .B2(n7287), .A(n7358), .ZN(n7289) );
  NAND2_X1 U8927 ( .A1(n7289), .A2(n8361), .ZN(n7290) );
  OAI211_X1 U8928 ( .C1(n7292), .C2(n9860), .A(n7291), .B(n7290), .ZN(P2_U3193) );
  NOR2_X2 U8929 ( .A1(n7293), .A2(n8626), .ZN(n8600) );
  NAND3_X1 U8930 ( .A1(n8109), .A2(n7294), .A3(n9901), .ZN(n7295) );
  OAI211_X1 U8931 ( .C1(n8624), .C2(n7297), .A(n7296), .B(n7295), .ZN(n7298)
         );
  MUX2_X1 U8932 ( .A(n7298), .B(P2_REG2_REG_0__SCAN_IN), .S(n8582), .Z(n7299)
         );
  AOI21_X1 U8933 ( .B1(n8600), .B2(n7300), .A(n7299), .ZN(n7301) );
  INV_X1 U8934 ( .A(n7301), .ZN(P2_U3233) );
  NAND2_X1 U8935 ( .A1(n7311), .A2(n7425), .ZN(n7302) );
  XNOR2_X1 U8936 ( .A(n7439), .B(n7437), .ZN(n7309) );
  XNOR2_X1 U8937 ( .A(n7436), .B(n7309), .ZN(n9742) );
  NAND2_X1 U8938 ( .A1(n9742), .A2(n7304), .ZN(n7315) );
  OR2_X1 U8939 ( .A1(n7306), .A2(n7305), .ZN(n7308) );
  NAND2_X1 U8940 ( .A1(n7308), .A2(n7307), .ZN(n7434) );
  INV_X1 U8941 ( .A(n7309), .ZN(n7310) );
  XNOR2_X1 U8942 ( .A(n7434), .B(n7310), .ZN(n7313) );
  OAI22_X1 U8943 ( .A1(n7473), .A2(n9774), .B1(n7311), .B2(n9776), .ZN(n7312)
         );
  AOI21_X1 U8944 ( .B1(n7313), .B2(n9765), .A(n7312), .ZN(n7314) );
  AND2_X1 U8945 ( .A1(n7315), .A2(n7314), .ZN(n9744) );
  AOI21_X1 U8946 ( .B1(n7316), .B2(n7437), .A(n9792), .ZN(n7317) );
  NAND2_X1 U8947 ( .A1(n7317), .A2(n7468), .ZN(n9739) );
  AOI22_X1 U8948 ( .A1(n9293), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n7549), .B2(
        n9291), .ZN(n7319) );
  NAND2_X1 U8949 ( .A1(n9299), .A2(n7437), .ZN(n7318) );
  OAI211_X1 U8950 ( .C1(n9739), .C2(n9302), .A(n7319), .B(n7318), .ZN(n7320)
         );
  AOI21_X1 U8951 ( .B1(n9742), .B2(n7321), .A(n7320), .ZN(n7322) );
  OAI21_X1 U8952 ( .B1(n9744), .B2(n9293), .A(n7322), .ZN(P1_U3285) );
  OAI21_X1 U8953 ( .B1(n7323), .B2(n8111), .A(n7479), .ZN(n7505) );
  INV_X1 U8954 ( .A(n8321), .ZN(n7539) );
  XOR2_X1 U8955 ( .A(n7324), .B(n8111), .Z(n7325) );
  OAI222_X1 U8956 ( .A1(n8622), .A2(n7539), .B1(n8620), .B2(n7333), .C1(n7325), 
        .C2(n8618), .ZN(n7502) );
  AOI21_X1 U8957 ( .B1(n9906), .B2(n7505), .A(n7502), .ZN(n7412) );
  AOI22_X1 U8958 ( .A1(n8675), .A2(n7336), .B1(n9927), .B2(
        P2_REG1_REG_5__SCAN_IN), .ZN(n7326) );
  OAI21_X1 U8959 ( .B1(n7412), .B2(n9927), .A(n7326), .ZN(P2_U3464) );
  INV_X1 U8960 ( .A(n7329), .ZN(n7327) );
  XNOR2_X1 U8961 ( .A(n7183), .B(n7336), .ZN(n7386) );
  XNOR2_X1 U8962 ( .A(n7386), .B(n8322), .ZN(n7330) );
  NOR3_X1 U8963 ( .A1(n7327), .A2(n4757), .A3(n7330), .ZN(n7332) );
  INV_X1 U8964 ( .A(n7388), .ZN(n7331) );
  OAI21_X1 U8965 ( .B1(n7332), .B2(n7331), .A(n8005), .ZN(n7338) );
  OAI22_X1 U8966 ( .A1(n8031), .A2(n7333), .B1(n7539), .B2(n8081), .ZN(n7334)
         );
  AOI211_X1 U8967 ( .C1(n7336), .C2(n8089), .A(n7335), .B(n7334), .ZN(n7337)
         );
  OAI211_X1 U8968 ( .C1(n7500), .C2(n8061), .A(n7338), .B(n7337), .ZN(P2_U3167) );
  INV_X1 U8969 ( .A(n8089), .ZN(n8055) );
  OAI22_X1 U8970 ( .A1(n8031), .A2(n6182), .B1(n8055), .B2(n9869), .ZN(n7339)
         );
  AOI21_X1 U8971 ( .B1(n8009), .B2(n8324), .A(n7339), .ZN(n7345) );
  OAI21_X1 U8972 ( .B1(n7342), .B2(n7341), .A(n7340), .ZN(n7343) );
  NAND2_X1 U8973 ( .A1(n7343), .A2(n8005), .ZN(n7344) );
  OAI211_X1 U8974 ( .C1(n7401), .C2(n7346), .A(n7345), .B(n7344), .ZN(P2_U3177) );
  INV_X1 U8975 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n7353) );
  INV_X1 U8976 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n7347) );
  OR2_X1 U8977 ( .A1(n7348), .A2(n7347), .ZN(n7352) );
  INV_X1 U8978 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n7349) );
  OR2_X1 U8979 ( .A1(n7350), .A2(n7349), .ZN(n7351) );
  OAI211_X1 U8980 ( .C1(n6186), .C2(n7353), .A(n7352), .B(n7351), .ZN(n7354)
         );
  INV_X1 U8981 ( .A(n7354), .ZN(n7355) );
  NAND2_X1 U8982 ( .A1(n8429), .A2(P2_U3893), .ZN(n7357) );
  OAI21_X1 U8983 ( .B1(P2_U3893), .B2(n9473), .A(n7357), .ZN(P2_U3522) );
  OAI21_X1 U8984 ( .B1(n7359), .B2(n4776), .A(n7358), .ZN(n7572) );
  MUX2_X1 U8985 ( .A(P2_REG2_REG_12__SCAN_IN), .B(P2_REG1_REG_12__SCAN_IN), 
        .S(n8415), .Z(n7361) );
  NOR2_X1 U8986 ( .A1(n7361), .A2(n7360), .ZN(n7571) );
  INV_X1 U8987 ( .A(n7571), .ZN(n7362) );
  NAND2_X1 U8988 ( .A1(n7361), .A2(n7360), .ZN(n7570) );
  NAND2_X1 U8989 ( .A1(n7362), .A2(n7570), .ZN(n7363) );
  XNOR2_X1 U8990 ( .A(n7572), .B(n7363), .ZN(n7380) );
  NOR2_X1 U8991 ( .A1(n7370), .A2(n7364), .ZN(n7366) );
  INV_X1 U8992 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n7578) );
  MUX2_X1 U8993 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n7578), .S(n7579), .Z(n7367)
         );
  OAI21_X1 U8994 ( .B1(n4501), .B2(n4500), .A(n7581), .ZN(n7378) );
  INV_X1 U8995 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n9966) );
  NOR2_X1 U8996 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10067), .ZN(n7857) );
  AOI21_X1 U8997 ( .B1(n9846), .B2(n7579), .A(n7857), .ZN(n7368) );
  OAI21_X1 U8998 ( .B1(n8387), .B2(n9966), .A(n7368), .ZN(n7377) );
  NOR2_X1 U8999 ( .A1(n7370), .A2(n7369), .ZN(n7372) );
  NOR2_X1 U9000 ( .A1(n7372), .A2(n7371), .ZN(n7374) );
  MUX2_X1 U9001 ( .A(P2_REG2_REG_12__SCAN_IN), .B(n7755), .S(n7579), .Z(n7373)
         );
  NAND2_X1 U9002 ( .A1(n7374), .A2(n7373), .ZN(n7375) );
  AOI21_X1 U9003 ( .B1(n7566), .B2(n7375), .A(n9856), .ZN(n7376) );
  AOI211_X1 U9004 ( .C1(n8426), .C2(n7378), .A(n7377), .B(n7376), .ZN(n7379)
         );
  OAI21_X1 U9005 ( .B1(n9858), .B2(n7380), .A(n7379), .ZN(P2_U3194) );
  INV_X1 U9006 ( .A(n7381), .ZN(n7385) );
  OAI222_X1 U9007 ( .A1(P1_U3086), .A2(n7383), .B1(n9484), .B2(n7385), .C1(
        n7382), .C2(n9487), .ZN(P1_U3335) );
  INV_X1 U9008 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7384) );
  OAI222_X1 U9009 ( .A1(n8298), .A2(P2_U3151), .B1(n8777), .B2(n7385), .C1(
        n7384), .C2(n7741), .ZN(P2_U3275) );
  NAND2_X1 U9010 ( .A1(n7386), .A2(n7495), .ZN(n7387) );
  NAND2_X1 U9011 ( .A1(n7388), .A2(n7387), .ZN(n7389) );
  XNOR2_X1 U9012 ( .A(n7183), .B(n9879), .ZN(n7529) );
  XNOR2_X1 U9013 ( .A(n7529), .B(n8321), .ZN(n7390) );
  AOI21_X1 U9014 ( .B1(n7389), .B2(n7390), .A(n8084), .ZN(n7393) );
  INV_X1 U9015 ( .A(n7389), .ZN(n7392) );
  INV_X1 U9016 ( .A(n7390), .ZN(n7391) );
  NAND2_X1 U9017 ( .A1(n7392), .A2(n7391), .ZN(n7535) );
  NAND2_X1 U9018 ( .A1(n7393), .A2(n7535), .ZN(n7398) );
  INV_X1 U9019 ( .A(n8320), .ZN(n7597) );
  OAI22_X1 U9020 ( .A1(n8031), .A2(n7495), .B1(n7597), .B2(n8081), .ZN(n7394)
         );
  AOI211_X1 U9021 ( .C1(n7396), .C2(n8089), .A(n7395), .B(n7394), .ZN(n7397)
         );
  OAI211_X1 U9022 ( .C1(n7481), .C2(n8061), .A(n7398), .B(n7397), .ZN(P2_U3179) );
  AOI21_X1 U9023 ( .B1(n7400), .B2(n7399), .A(n4449), .ZN(n7406) );
  INV_X1 U9024 ( .A(n7401), .ZN(n7404) );
  AOI22_X1 U9025 ( .A1(n8078), .A2(n8326), .B1(n8089), .B2(n6181), .ZN(n7402)
         );
  OAI21_X1 U9026 ( .B1(n6199), .B2(n8081), .A(n7402), .ZN(n7403) );
  AOI21_X1 U9027 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(n7404), .A(n7403), .ZN(
        n7405) );
  OAI21_X1 U9028 ( .B1(n8084), .B2(n7406), .A(n7405), .ZN(P2_U3162) );
  INV_X1 U9029 ( .A(n7407), .ZN(n7445) );
  INV_X1 U9030 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7408) );
  OAI222_X1 U9031 ( .A1(n8139), .A2(P2_U3151), .B1(n8777), .B2(n7445), .C1(
        n7408), .C2(n7741), .ZN(P2_U3274) );
  INV_X1 U9032 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n7409) );
  OAI22_X1 U9033 ( .A1(n8740), .A2(n7501), .B1(n7409), .B2(n9914), .ZN(n7410)
         );
  INV_X1 U9034 ( .A(n7410), .ZN(n7411) );
  OAI21_X1 U9035 ( .B1(n7412), .B2(n9915), .A(n7411), .ZN(P2_U3405) );
  INV_X1 U9036 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n7413) );
  OAI22_X1 U9037 ( .A1(n8740), .A2(n7507), .B1(n7413), .B2(n9914), .ZN(n7414)
         );
  INV_X1 U9038 ( .A(n7414), .ZN(n7415) );
  OAI21_X1 U9039 ( .B1(n7416), .B2(n9915), .A(n7415), .ZN(P2_U3399) );
  INV_X1 U9040 ( .A(n7417), .ZN(n7420) );
  OAI211_X1 U9041 ( .C1(n7420), .C2(n9738), .A(n7419), .B(n7418), .ZN(n7427)
         );
  INV_X1 U9042 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n7421) );
  OAI22_X1 U9043 ( .A1(n9465), .A2(n7425), .B1(n9798), .B2(n7421), .ZN(n7422)
         );
  AOI21_X1 U9044 ( .B1(n7427), .B2(n9798), .A(n7422), .ZN(n7423) );
  INV_X1 U9045 ( .A(n7423), .ZN(P1_U3474) );
  INV_X1 U9046 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n7424) );
  OAI22_X1 U9047 ( .A1(n9423), .A2(n7425), .B1(n9813), .B2(n7424), .ZN(n7426)
         );
  AOI21_X1 U9048 ( .B1(n7427), .B2(n9813), .A(n7426), .ZN(n7428) );
  INV_X1 U9049 ( .A(n7428), .ZN(P1_U3529) );
  NAND2_X1 U9050 ( .A1(n7430), .A2(n7429), .ZN(n7465) );
  INV_X1 U9051 ( .A(n7431), .ZN(n7433) );
  OAI21_X1 U9052 ( .B1(n7434), .B2(n7433), .A(n7432), .ZN(n7435) );
  XOR2_X1 U9053 ( .A(n7465), .B(n7435), .Z(n9750) );
  XNOR2_X1 U9054 ( .A(n7466), .B(n7465), .ZN(n9752) );
  NAND2_X1 U9055 ( .A1(n9752), .A2(n9212), .ZN(n7444) );
  AOI22_X1 U9056 ( .A1(n9293), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n7646), .B2(
        n9291), .ZN(n7438) );
  OAI21_X1 U9057 ( .B1(n7439), .B2(n9297), .A(n7438), .ZN(n7442) );
  XNOR2_X1 U9058 ( .A(n7468), .B(n4595), .ZN(n7440) );
  INV_X1 U9059 ( .A(n7814), .ZN(n8956) );
  AOI22_X1 U9060 ( .A1(n7440), .A2(n9319), .B1(n9757), .B2(n8956), .ZN(n9749)
         );
  NOR2_X1 U9061 ( .A1(n9749), .A2(n9302), .ZN(n7441) );
  AOI211_X1 U9062 ( .C1(n9299), .C2(n9747), .A(n7442), .B(n7441), .ZN(n7443)
         );
  OAI211_X1 U9063 ( .C1(n9750), .C2(n9173), .A(n7444), .B(n7443), .ZN(P1_U3284) );
  OAI222_X1 U9064 ( .A1(n9487), .A2(n7447), .B1(P1_U3086), .B2(n7446), .C1(
        n9481), .C2(n7445), .ZN(P1_U3334) );
  AND2_X1 U9065 ( .A1(n7609), .A2(n7448), .ZN(n7450) );
  OAI211_X1 U9066 ( .C1(n7450), .C2(n8116), .A(n7449), .B(n8596), .ZN(n7452)
         );
  AOI22_X1 U9067 ( .A1(n8591), .A2(n8320), .B1(n8318), .B2(n8593), .ZN(n7451)
         );
  AND2_X1 U9068 ( .A1(n7452), .A2(n7451), .ZN(n9893) );
  OAI22_X1 U9069 ( .A1(n8550), .A2(n9890), .B1(n7603), .B2(n8624), .ZN(n7453)
         );
  AOI21_X1 U9070 ( .B1(P2_REG2_REG_8__SCAN_IN), .B2(n8582), .A(n7453), .ZN(
        n7458) );
  XNOR2_X1 U9071 ( .A(n7454), .B(n8116), .ZN(n9889) );
  NAND2_X1 U9072 ( .A1(n9889), .A2(n8630), .ZN(n7457) );
  OAI211_X1 U9073 ( .C1(n9893), .C2(n8582), .A(n7458), .B(n7457), .ZN(P2_U3225) );
  XNOR2_X1 U9074 ( .A(n8108), .B(n7459), .ZN(n9866) );
  AOI22_X1 U9075 ( .A1(n8600), .A2(n6181), .B1(n8599), .B2(
        P2_REG3_REG_1__SCAN_IN), .ZN(n7464) );
  XNOR2_X1 U9076 ( .A(n8108), .B(n7460), .ZN(n7461) );
  AOI222_X1 U9077 ( .A1(n8596), .A2(n7461), .B1(n8325), .B2(n8593), .C1(n8326), 
        .C2(n8591), .ZN(n9864) );
  MUX2_X1 U9078 ( .A(n9864), .B(n7462), .S(n8582), .Z(n7463) );
  OAI211_X1 U9079 ( .C1(n8603), .C2(n9866), .A(n7464), .B(n7463), .ZN(P2_U3232) );
  XOR2_X1 U9080 ( .A(n7514), .B(n7515), .Z(n9761) );
  OAI21_X1 U9081 ( .B1(n7467), .B2(n7514), .A(n7517), .ZN(n9764) );
  INV_X1 U9082 ( .A(n9173), .ZN(n9304) );
  INV_X1 U9083 ( .A(n7523), .ZN(n7469) );
  OAI211_X1 U9084 ( .C1(n4937), .C2(n7470), .A(n7469), .B(n9319), .ZN(n9759)
         );
  AOI22_X1 U9085 ( .A1(n9293), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n7762), .B2(
        n9291), .ZN(n7472) );
  INV_X1 U9086 ( .A(n9777), .ZN(n9756) );
  NAND2_X1 U9087 ( .A1(n9294), .A2(n9756), .ZN(n7471) );
  OAI211_X1 U9088 ( .C1(n7473), .C2(n9297), .A(n7472), .B(n7471), .ZN(n7474)
         );
  AOI21_X1 U9089 ( .B1(n9299), .B2(n7513), .A(n7474), .ZN(n7475) );
  OAI21_X1 U9090 ( .B1(n9759), .B2(n9302), .A(n7475), .ZN(n7476) );
  AOI21_X1 U9091 ( .B1(n9764), .B2(n9304), .A(n7476), .ZN(n7477) );
  OAI21_X1 U9092 ( .B1(n9761), .B2(n9306), .A(n7477), .ZN(P1_U3283) );
  NAND2_X1 U9093 ( .A1(n7479), .A2(n7478), .ZN(n7480) );
  XNOR2_X1 U9094 ( .A(n7480), .B(n8114), .ZN(n9882) );
  OAI22_X1 U9095 ( .A1(n8550), .A2(n9879), .B1(n7481), .B2(n8624), .ZN(n7488)
         );
  NAND2_X1 U9096 ( .A1(n7482), .A2(n8114), .ZN(n7483) );
  NAND3_X1 U9097 ( .A1(n7484), .A2(n8596), .A3(n7483), .ZN(n7486) );
  AOI22_X1 U9098 ( .A1(n8593), .A2(n8320), .B1(n8322), .B2(n8591), .ZN(n7485)
         );
  NAND2_X1 U9099 ( .A1(n7486), .A2(n7485), .ZN(n9880) );
  MUX2_X1 U9100 ( .A(n9880), .B(P2_REG2_REG_6__SCAN_IN), .S(n8582), .Z(n7487)
         );
  AOI211_X1 U9101 ( .C1(n8630), .C2(n9882), .A(n7488), .B(n7487), .ZN(n7489)
         );
  INV_X1 U9102 ( .A(n7489), .ZN(P2_U3227) );
  OAI21_X1 U9103 ( .B1(n7491), .B2(n8158), .A(n7490), .ZN(n9878) );
  OAI22_X1 U9104 ( .A1(n8550), .A2(n9875), .B1(n7492), .B2(n8624), .ZN(n7498)
         );
  XNOR2_X1 U9105 ( .A(n7493), .B(n8158), .ZN(n7494) );
  OAI222_X1 U9106 ( .A1(n8620), .A2(n7496), .B1(n8622), .B2(n7495), .C1(n7494), 
        .C2(n8618), .ZN(n9876) );
  MUX2_X1 U9107 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n9876), .S(n8633), .Z(n7497)
         );
  AOI211_X1 U9108 ( .C1(n8630), .C2(n9878), .A(n7498), .B(n7497), .ZN(n7499)
         );
  INV_X1 U9109 ( .A(n7499), .ZN(P2_U3229) );
  OAI22_X1 U9110 ( .A1(n8550), .A2(n7501), .B1(n7500), .B2(n8624), .ZN(n7504)
         );
  MUX2_X1 U9111 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n7502), .S(n8633), .Z(n7503)
         );
  AOI211_X1 U9112 ( .C1(n8630), .C2(n7505), .A(n7504), .B(n7503), .ZN(n7506)
         );
  INV_X1 U9113 ( .A(n7506), .ZN(P2_U3228) );
  OAI22_X1 U9114 ( .A1(n8550), .A2(n7507), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        n8624), .ZN(n7510) );
  MUX2_X1 U9115 ( .A(n7508), .B(P2_REG2_REG_3__SCAN_IN), .S(n8582), .Z(n7509)
         );
  AOI211_X1 U9116 ( .C1(n8630), .C2(n7511), .A(n7510), .B(n7509), .ZN(n7512)
         );
  INV_X1 U9117 ( .A(n7512), .ZN(P2_U3230) );
  XNOR2_X1 U9118 ( .A(n7624), .B(n7623), .ZN(n9772) );
  INV_X1 U9119 ( .A(n9772), .ZN(n7528) );
  NAND2_X1 U9120 ( .A1(n7517), .A2(n7516), .ZN(n7518) );
  NAND2_X1 U9121 ( .A1(n7518), .A2(n7623), .ZN(n7519) );
  NAND3_X1 U9122 ( .A1(n7519), .A2(n7620), .A3(n9765), .ZN(n7522) );
  OAI22_X1 U9123 ( .A1(n7814), .A2(n9776), .B1(n7689), .B2(n9774), .ZN(n7520)
         );
  INV_X1 U9124 ( .A(n7520), .ZN(n7521) );
  NAND2_X1 U9125 ( .A1(n7522), .A2(n7521), .ZN(n9771) );
  INV_X1 U9126 ( .A(n7816), .ZN(n9769) );
  NAND2_X1 U9127 ( .A1(n7523), .A2(n9769), .ZN(n7625) );
  OAI211_X1 U9128 ( .C1(n7523), .C2(n9769), .A(n9319), .B(n7625), .ZN(n9767)
         );
  AOI22_X1 U9129 ( .A1(n9293), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n7812), .B2(
        n9291), .ZN(n7525) );
  NAND2_X1 U9130 ( .A1(n7816), .A2(n9299), .ZN(n7524) );
  OAI211_X1 U9131 ( .C1(n9767), .C2(n9302), .A(n7525), .B(n7524), .ZN(n7526)
         );
  AOI21_X1 U9132 ( .B1(n9771), .B2(n9265), .A(n7526), .ZN(n7527) );
  OAI21_X1 U9133 ( .B1(n7528), .B2(n9306), .A(n7527), .ZN(P1_U3282) );
  NAND2_X1 U9134 ( .A1(n7529), .A2(n8321), .ZN(n7533) );
  AND2_X1 U9135 ( .A1(n7535), .A2(n7533), .ZN(n7537) );
  XNOR2_X1 U9136 ( .A(n7183), .B(n7542), .ZN(n7530) );
  NAND2_X1 U9137 ( .A1(n7530), .A2(n7597), .ZN(n7590) );
  INV_X1 U9138 ( .A(n7530), .ZN(n7531) );
  NAND2_X1 U9139 ( .A1(n7531), .A2(n8320), .ZN(n7532) );
  AND2_X1 U9140 ( .A1(n7590), .A2(n7532), .ZN(n7536) );
  AND2_X1 U9141 ( .A1(n7533), .A2(n7536), .ZN(n7534) );
  OAI21_X1 U9142 ( .B1(n7537), .B2(n7536), .A(n7591), .ZN(n7538) );
  NAND2_X1 U9143 ( .A1(n7538), .A2(n8005), .ZN(n7544) );
  INV_X1 U9144 ( .A(n8319), .ZN(n7658) );
  OAI22_X1 U9145 ( .A1(n8031), .A2(n7539), .B1(n7658), .B2(n8081), .ZN(n7540)
         );
  AOI211_X1 U9146 ( .C1(n7542), .C2(n8089), .A(n7541), .B(n7540), .ZN(n7543)
         );
  OAI211_X1 U9147 ( .C1(n7606), .C2(n8061), .A(n7544), .B(n7543), .ZN(P2_U3153) );
  INV_X1 U9148 ( .A(n7545), .ZN(n7887) );
  OAI222_X1 U9149 ( .A1(P2_U3151), .A2(n8149), .B1(n8777), .B2(n7887), .C1(
        n7546), .C2(n7741), .ZN(P2_U3273) );
  OAI21_X1 U9150 ( .B1(n7548), .B2(n4447), .A(n7547), .ZN(n7554) );
  INV_X1 U9151 ( .A(n8928), .ZN(n8948) );
  AOI22_X1 U9152 ( .A1(n8927), .A2(n7549), .B1(n8926), .B2(n8957), .ZN(n7552)
         );
  NAND2_X1 U9153 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n9527) );
  INV_X1 U9154 ( .A(n9527), .ZN(n7550) );
  AOI21_X1 U9155 ( .B1(n8945), .B2(n9755), .A(n7550), .ZN(n7551) );
  OAI211_X1 U9156 ( .C1(n4596), .C2(n8948), .A(n7552), .B(n7551), .ZN(n7553)
         );
  AOI21_X1 U9157 ( .B1(n7554), .B2(n8936), .A(n7553), .ZN(n7555) );
  INV_X1 U9158 ( .A(n7555), .ZN(P1_U3221) );
  OAI21_X1 U9159 ( .B1(n7557), .B2(n8118), .A(n7556), .ZN(n7558) );
  AOI222_X1 U9160 ( .A1(n8596), .A2(n7558), .B1(n8317), .B2(n8593), .C1(n8319), 
        .C2(n8591), .ZN(n7675) );
  NAND2_X1 U9161 ( .A1(n7559), .A2(n8118), .ZN(n7560) );
  AND2_X1 U9162 ( .A1(n7561), .A2(n7560), .ZN(n7677) );
  NOR2_X1 U9163 ( .A1(n8550), .A2(n7679), .ZN(n7563) );
  OAI22_X1 U9164 ( .A1(n8633), .A2(n7063), .B1(n7663), .B2(n8624), .ZN(n7562)
         );
  AOI211_X1 U9165 ( .C1(n7677), .C2(n8630), .A(n7563), .B(n7562), .ZN(n7564)
         );
  OAI21_X1 U9166 ( .B1(n7675), .B2(n8582), .A(n7564), .ZN(P2_U3224) );
  OR2_X1 U9167 ( .A1(n7579), .A2(n7755), .ZN(n7565) );
  AOI21_X1 U9168 ( .B1(n7567), .B2(n7569), .A(n8342), .ZN(n7587) );
  MUX2_X1 U9169 ( .A(n7569), .B(n7568), .S(n8415), .Z(n8346) );
  XNOR2_X1 U9170 ( .A(n8346), .B(n8351), .ZN(n7574) );
  OAI21_X1 U9171 ( .B1(n7572), .B2(n7571), .A(n7570), .ZN(n7573) );
  NOR2_X1 U9172 ( .A1(n7573), .A2(n7574), .ZN(n8345) );
  AOI21_X1 U9173 ( .B1(n7574), .B2(n7573), .A(n8345), .ZN(n7577) );
  AND2_X1 U9174 ( .A1(P2_U3151), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n8041) );
  INV_X1 U9175 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n9970) );
  NOR2_X1 U9176 ( .A1(n8387), .A2(n9970), .ZN(n7575) );
  AOI211_X1 U9177 ( .C1(n8351), .C2(n9846), .A(n8041), .B(n7575), .ZN(n7576)
         );
  OAI21_X1 U9178 ( .B1(n7577), .B2(n9858), .A(n7576), .ZN(n7585) );
  OR2_X1 U9179 ( .A1(n7579), .A2(n7578), .ZN(n7580) );
  XNOR2_X1 U9180 ( .A(n8351), .B(n8350), .ZN(n7582) );
  NOR2_X1 U9181 ( .A1(n7568), .A2(n7582), .ZN(n8352) );
  AOI21_X1 U9182 ( .B1(n7568), .B2(n7582), .A(n8352), .ZN(n7583) );
  NOR2_X1 U9183 ( .A1(n7583), .A2(n9860), .ZN(n7584) );
  NOR2_X1 U9184 ( .A1(n7585), .A2(n7584), .ZN(n7586) );
  OAI21_X1 U9185 ( .B1(n7587), .B2(n9856), .A(n7586), .ZN(P2_U3195) );
  INV_X1 U9186 ( .A(n7591), .ZN(n7589) );
  INV_X1 U9187 ( .A(n7590), .ZN(n7588) );
  XNOR2_X1 U9188 ( .A(n7183), .B(n7600), .ZN(n7651) );
  XNOR2_X1 U9189 ( .A(n7651), .B(n8319), .ZN(n7592) );
  NOR3_X1 U9190 ( .A1(n7589), .A2(n7588), .A3(n7592), .ZN(n7595) );
  NAND2_X1 U9191 ( .A1(n7591), .A2(n7590), .ZN(n7593) );
  NAND2_X1 U9192 ( .A1(n7593), .A2(n7592), .ZN(n7653) );
  INV_X1 U9193 ( .A(n7653), .ZN(n7594) );
  OAI21_X1 U9194 ( .B1(n7595), .B2(n7594), .A(n8005), .ZN(n7602) );
  INV_X1 U9195 ( .A(n8318), .ZN(n7596) );
  OAI22_X1 U9196 ( .A1(n8031), .A2(n7597), .B1(n7596), .B2(n8081), .ZN(n7598)
         );
  AOI211_X1 U9197 ( .C1(n7600), .C2(n8089), .A(n7599), .B(n7598), .ZN(n7601)
         );
  OAI211_X1 U9198 ( .C1(n7603), .C2(n8061), .A(n7602), .B(n7601), .ZN(P2_U3161) );
  NAND2_X1 U9199 ( .A1(n7604), .A2(n8172), .ZN(n7605) );
  XNOR2_X1 U9200 ( .A(n7605), .B(n6268), .ZN(n9887) );
  OAI22_X1 U9201 ( .A1(n8550), .A2(n9884), .B1(n7606), .B2(n8624), .ZN(n7615)
         );
  NAND2_X1 U9202 ( .A1(n9887), .A2(n7666), .ZN(n7613) );
  NAND2_X1 U9203 ( .A1(n7607), .A2(n8179), .ZN(n7608) );
  NAND2_X1 U9204 ( .A1(n7609), .A2(n7608), .ZN(n7610) );
  NAND2_X1 U9205 ( .A1(n7610), .A2(n8596), .ZN(n7612) );
  AOI22_X1 U9206 ( .A1(n8591), .A2(n8321), .B1(n8319), .B2(n8593), .ZN(n7611)
         );
  NAND3_X1 U9207 ( .A1(n7613), .A2(n7612), .A3(n7611), .ZN(n9885) );
  MUX2_X1 U9208 ( .A(n9885), .B(P2_REG2_REG_7__SCAN_IN), .S(n8582), .Z(n7614)
         );
  AOI211_X1 U9209 ( .C1(n9887), .C2(n7947), .A(n7615), .B(n7614), .ZN(n7616)
         );
  INV_X1 U9210 ( .A(n7616), .ZN(P2_U3226) );
  INV_X1 U9211 ( .A(n7617), .ZN(n7622) );
  INV_X1 U9212 ( .A(n7618), .ZN(n7690) );
  AOI21_X1 U9213 ( .B1(n7620), .B2(n7619), .A(n7690), .ZN(n7621) );
  NOR2_X1 U9214 ( .A1(n7622), .A2(n7621), .ZN(n9782) );
  XNOR2_X1 U9215 ( .A(n7691), .B(n7690), .ZN(n9785) );
  NAND2_X1 U9216 ( .A1(n9785), .A2(n9212), .ZN(n7632) );
  AOI211_X1 U9217 ( .C1(n9780), .C2(n7625), .A(n9792), .B(n4598), .ZN(n9778)
         );
  INV_X1 U9218 ( .A(n9780), .ZN(n7626) );
  NOR2_X1 U9219 ( .A1(n7626), .A2(n9273), .ZN(n7630) );
  AOI22_X1 U9220 ( .A1(n9293), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n8838), .B2(
        n9291), .ZN(n7628) );
  NAND2_X1 U9221 ( .A1(n9294), .A2(n8954), .ZN(n7627) );
  OAI211_X1 U9222 ( .C1(n9777), .C2(n9297), .A(n7628), .B(n7627), .ZN(n7629)
         );
  AOI211_X1 U9223 ( .C1(n9778), .C2(n9284), .A(n7630), .B(n7629), .ZN(n7631)
         );
  OAI211_X1 U9224 ( .C1(n9782), .C2(n9173), .A(n7632), .B(n7631), .ZN(P1_U3281) );
  INV_X1 U9225 ( .A(n7637), .ZN(n7635) );
  AOI21_X1 U9226 ( .B1(P1_DATAO_REG_23__SCAN_IN), .B2(n8774), .A(n7633), .ZN(
        n7634) );
  OAI21_X1 U9227 ( .B1(n7635), .B2(n8777), .A(n7634), .ZN(P2_U3272) );
  NAND2_X1 U9228 ( .A1(n7637), .A2(n7636), .ZN(n7639) );
  OAI211_X1 U9229 ( .C1(n7640), .C2(n9487), .A(n7639), .B(n7638), .ZN(P1_U3332) );
  OAI21_X1 U9230 ( .B1(n7643), .B2(n7641), .A(n7642), .ZN(n7644) );
  NAND2_X1 U9231 ( .A1(n7644), .A2(n8936), .ZN(n7650) );
  NOR2_X1 U9232 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7645), .ZN(n9007) );
  INV_X1 U9233 ( .A(n7646), .ZN(n7647) );
  OAI22_X1 U9234 ( .A1(n8941), .A2(n7647), .B1(n8899), .B2(n7814), .ZN(n7648)
         );
  AOI211_X1 U9235 ( .C1(n8926), .C2(n9746), .A(n9007), .B(n7648), .ZN(n7649)
         );
  OAI211_X1 U9236 ( .C1(n4595), .C2(n8948), .A(n7650), .B(n7649), .ZN(P1_U3231) );
  NAND2_X1 U9237 ( .A1(n7651), .A2(n7658), .ZN(n7652) );
  XNOR2_X1 U9238 ( .A(n7183), .B(n7679), .ZN(n7769) );
  XNOR2_X1 U9239 ( .A(n7769), .B(n8318), .ZN(n7655) );
  AOI21_X1 U9240 ( .B1(n7654), .B2(n7655), .A(n8084), .ZN(n7657) );
  INV_X1 U9241 ( .A(n7655), .ZN(n7656) );
  NAND2_X1 U9242 ( .A1(n7657), .A2(n7771), .ZN(n7662) );
  OAI22_X1 U9243 ( .A1(n8031), .A2(n7658), .B1(n7788), .B2(n8081), .ZN(n7659)
         );
  AOI211_X1 U9244 ( .C1(n7682), .C2(n8089), .A(n7660), .B(n7659), .ZN(n7661)
         );
  OAI211_X1 U9245 ( .C1(n7663), .C2(n8061), .A(n7662), .B(n7661), .ZN(P2_U3171) );
  XNOR2_X1 U9246 ( .A(n7788), .B(n7776), .ZN(n8122) );
  XOR2_X1 U9247 ( .A(n8122), .B(n7664), .Z(n7669) );
  AOI22_X1 U9248 ( .A1(n8593), .A2(n8316), .B1(n8318), .B2(n8591), .ZN(n7668)
         );
  XNOR2_X1 U9249 ( .A(n7665), .B(n8122), .ZN(n9899) );
  NAND2_X1 U9250 ( .A1(n9899), .A2(n7666), .ZN(n7667) );
  OAI211_X1 U9251 ( .C1(n7669), .C2(n8618), .A(n7668), .B(n7667), .ZN(n9896)
         );
  INV_X1 U9252 ( .A(n9896), .ZN(n7674) );
  INV_X1 U9253 ( .A(n7670), .ZN(n7774) );
  AOI22_X1 U9254 ( .A1(n8582), .A2(P2_REG2_REG_10__SCAN_IN), .B1(n8599), .B2(
        n7774), .ZN(n7671) );
  OAI21_X1 U9255 ( .B1(n8550), .B2(n9895), .A(n7671), .ZN(n7672) );
  AOI21_X1 U9256 ( .B1(n9899), .B2(n7947), .A(n7672), .ZN(n7673) );
  OAI21_X1 U9257 ( .B1(n7674), .B2(n8582), .A(n7673), .ZN(P2_U3223) );
  INV_X1 U9258 ( .A(n7675), .ZN(n7676) );
  AOI21_X1 U9259 ( .B1(n7677), .B2(n9906), .A(n7676), .ZN(n7684) );
  INV_X1 U9260 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n7678) );
  OAI22_X1 U9261 ( .A1(n8740), .A2(n7679), .B1(n7678), .B2(n9914), .ZN(n7680)
         );
  INV_X1 U9262 ( .A(n7680), .ZN(n7681) );
  OAI21_X1 U9263 ( .B1(n7684), .B2(n9915), .A(n7681), .ZN(P2_U3417) );
  AOI22_X1 U9264 ( .A1(n8675), .A2(n7682), .B1(n9927), .B2(
        P2_REG1_REG_9__SCAN_IN), .ZN(n7683) );
  OAI21_X1 U9265 ( .B1(n7684), .B2(n9927), .A(n7683), .ZN(P2_U3468) );
  AOI21_X1 U9266 ( .B1(n7685), .B2(n7708), .A(n9783), .ZN(n7688) );
  OAI22_X1 U9267 ( .A1(n7689), .A2(n9776), .B1(n8939), .B2(n9774), .ZN(n7686)
         );
  AOI21_X1 U9268 ( .B1(n7688), .B2(n7687), .A(n7686), .ZN(n9790) );
  INV_X1 U9269 ( .A(n7689), .ZN(n8955) );
  XNOR2_X1 U9270 ( .A(n7709), .B(n7708), .ZN(n9795) );
  NAND2_X1 U9271 ( .A1(n9795), .A2(n9212), .ZN(n7698) );
  NAND2_X1 U9272 ( .A1(n7692), .A2(n9788), .ZN(n7693) );
  NAND2_X1 U9273 ( .A1(n7712), .A2(n7693), .ZN(n9791) );
  INV_X1 U9274 ( .A(n9791), .ZN(n7696) );
  INV_X1 U9275 ( .A(n9788), .ZN(n7707) );
  AOI22_X1 U9276 ( .A1(n9293), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n8897), .B2(
        n9291), .ZN(n7694) );
  OAI21_X1 U9277 ( .B1(n7707), .B2(n9273), .A(n7694), .ZN(n7695) );
  AOI21_X1 U9278 ( .B1(n7696), .B2(n9143), .A(n7695), .ZN(n7697) );
  OAI211_X1 U9279 ( .C1(n9293), .C2(n9790), .A(n7698), .B(n7697), .ZN(P1_U3280) );
  INV_X1 U9280 ( .A(n7699), .ZN(n7702) );
  OAI222_X1 U9281 ( .A1(n6558), .A2(P2_U3151), .B1(n8777), .B2(n7702), .C1(
        n7700), .C2(n7741), .ZN(P2_U3271) );
  OAI222_X1 U9282 ( .A1(n7703), .A2(P1_U3086), .B1(n9484), .B2(n7702), .C1(
        n7701), .C2(n9487), .ZN(P1_U3331) );
  OAI21_X1 U9283 ( .B1(n7719), .B2(n7705), .A(n7704), .ZN(n7706) );
  NAND2_X1 U9284 ( .A1(n7706), .A2(n9765), .ZN(n9429) );
  XNOR2_X1 U9285 ( .A(n7720), .B(n7719), .ZN(n9424) );
  NAND2_X1 U9286 ( .A1(n9424), .A2(n9212), .ZN(n7718) );
  AOI22_X1 U9287 ( .A1(n9293), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n8792), .B2(
        n9291), .ZN(n7711) );
  INV_X1 U9288 ( .A(n9425), .ZN(n8952) );
  NAND2_X1 U9289 ( .A1(n9294), .A2(n8952), .ZN(n7710) );
  OAI211_X1 U9290 ( .C1(n9775), .C2(n9297), .A(n7711), .B(n7710), .ZN(n7716)
         );
  INV_X1 U9291 ( .A(n7725), .ZN(n7714) );
  AOI21_X1 U9292 ( .B1(n7712), .B2(n9427), .A(n9792), .ZN(n7713) );
  NAND2_X1 U9293 ( .A1(n7714), .A2(n7713), .ZN(n9428) );
  NOR2_X1 U9294 ( .A1(n9428), .A2(n9302), .ZN(n7715) );
  AOI211_X1 U9295 ( .C1(n9299), .C2(n9427), .A(n7716), .B(n7715), .ZN(n7717)
         );
  OAI211_X1 U9296 ( .C1(n9293), .C2(n9429), .A(n7718), .B(n7717), .ZN(P1_U3279) );
  XNOR2_X1 U9297 ( .A(n7820), .B(n7721), .ZN(n7845) );
  XNOR2_X1 U9298 ( .A(n7722), .B(n7721), .ZN(n7724) );
  OAI22_X1 U9299 ( .A1(n7824), .A2(n9774), .B1(n8939), .B2(n9776), .ZN(n7723)
         );
  AOI21_X1 U9300 ( .B1(n7724), .B2(n9765), .A(n7723), .ZN(n7844) );
  INV_X1 U9301 ( .A(n7844), .ZN(n7729) );
  OAI211_X1 U9302 ( .C1(n7725), .C2(n8949), .A(n7836), .B(n9319), .ZN(n7843)
         );
  AOI22_X1 U9303 ( .A1(n9293), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n8938), .B2(
        n9291), .ZN(n7727) );
  NAND2_X1 U9304 ( .A1(n7819), .A2(n9299), .ZN(n7726) );
  OAI211_X1 U9305 ( .C1(n7843), .C2(n9302), .A(n7727), .B(n7726), .ZN(n7728)
         );
  AOI21_X1 U9306 ( .B1(n7729), .B2(n9265), .A(n7728), .ZN(n7730) );
  OAI21_X1 U9307 ( .B1(n7845), .B2(n9306), .A(n7730), .ZN(P1_U3278) );
  XOR2_X1 U9308 ( .A(n7731), .B(n8119), .Z(n7732) );
  OAI222_X1 U9309 ( .A1(n8622), .A2(n8619), .B1(n8620), .B2(n7788), .C1(n7732), 
        .C2(n8618), .ZN(n9903) );
  INV_X1 U9310 ( .A(n9903), .ZN(n7737) );
  OAI21_X1 U9311 ( .B1(n7733), .B2(n8119), .A(n7747), .ZN(n9905) );
  NOR2_X1 U9312 ( .A1(n8550), .A2(n9902), .ZN(n7735) );
  OAI22_X1 U9313 ( .A1(n8633), .A2(n6309), .B1(n7795), .B2(n8624), .ZN(n7734)
         );
  AOI211_X1 U9314 ( .C1(n9905), .C2(n8630), .A(n7735), .B(n7734), .ZN(n7736)
         );
  OAI21_X1 U9315 ( .B1(n7737), .B2(n8582), .A(n7736), .ZN(P2_U3222) );
  INV_X1 U9316 ( .A(n7738), .ZN(n7743) );
  OAI222_X1 U9317 ( .A1(n7740), .A2(P1_U3086), .B1(n9484), .B2(n7743), .C1(
        n7739), .C2(n9487), .ZN(P1_U3330) );
  OAI222_X1 U9318 ( .A1(n6542), .A2(P2_U3151), .B1(n8777), .B2(n7743), .C1(
        n7742), .C2(n7741), .ZN(P2_U3270) );
  INV_X1 U9319 ( .A(n7744), .ZN(n7785) );
  AOI22_X1 U9320 ( .A1(n7745), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_26__SCAN_IN), .B2(n8774), .ZN(n7746) );
  OAI21_X1 U9321 ( .B1(n7785), .B2(n8777), .A(n7746), .ZN(P2_U3269) );
  INV_X1 U9322 ( .A(n7747), .ZN(n7748) );
  OAI21_X1 U9323 ( .B1(n7748), .B2(n8201), .A(n7752), .ZN(n7750) );
  NAND2_X1 U9324 ( .A1(n7750), .A2(n7749), .ZN(n9909) );
  OAI211_X1 U9325 ( .C1(n4441), .C2(n7752), .A(n8596), .B(n7751), .ZN(n7754)
         );
  AOI22_X1 U9326 ( .A1(n8591), .A2(n8316), .B1(n8314), .B2(n8593), .ZN(n7753)
         );
  NAND2_X1 U9327 ( .A1(n7754), .A2(n7753), .ZN(n9910) );
  NAND2_X1 U9328 ( .A1(n9910), .A2(n8633), .ZN(n7758) );
  OAI22_X1 U9329 ( .A1(n8633), .A2(n7755), .B1(n7855), .B2(n8624), .ZN(n7756)
         );
  AOI21_X1 U9330 ( .B1(n8600), .B2(n9912), .A(n7756), .ZN(n7757) );
  OAI211_X1 U9331 ( .C1(n8603), .C2(n9909), .A(n7758), .B(n7757), .ZN(P2_U3221) );
  OAI21_X1 U9332 ( .B1(n7761), .B2(n7760), .A(n7759), .ZN(n7767) );
  AOI22_X1 U9333 ( .A1(n7762), .A2(n8927), .B1(n8926), .B2(n9755), .ZN(n7765)
         );
  NAND2_X1 U9334 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n9499) );
  INV_X1 U9335 ( .A(n9499), .ZN(n7763) );
  AOI21_X1 U9336 ( .B1(n8945), .B2(n9756), .A(n7763), .ZN(n7764) );
  OAI211_X1 U9337 ( .C1(n4937), .C2(n8948), .A(n7765), .B(n7764), .ZN(n7766)
         );
  AOI21_X1 U9338 ( .B1(n7767), .B2(n8936), .A(n7766), .ZN(n7768) );
  INV_X1 U9339 ( .A(n7768), .ZN(P1_U3217) );
  NAND2_X1 U9340 ( .A1(n7769), .A2(n8318), .ZN(n7770) );
  XNOR2_X1 U9341 ( .A(n7183), .B(n7776), .ZN(n7772) );
  OAI21_X1 U9342 ( .B1(n7773), .B2(n7772), .A(n7793), .ZN(n7782) );
  NAND2_X1 U9343 ( .A1(n8077), .A2(n7774), .ZN(n7780) );
  AOI21_X1 U9344 ( .B1(n8078), .B2(n8318), .A(n7775), .ZN(n7779) );
  NAND2_X1 U9345 ( .A1(n8089), .A2(n7776), .ZN(n7778) );
  OR2_X1 U9346 ( .A1(n8081), .A2(n7852), .ZN(n7777) );
  NAND4_X1 U9347 ( .A1(n7780), .A2(n7779), .A3(n7778), .A4(n7777), .ZN(n7781)
         );
  AOI21_X1 U9348 ( .B1(n7782), .B2(n8005), .A(n7781), .ZN(n7783) );
  INV_X1 U9349 ( .A(n7783), .ZN(P2_U3157) );
  OAI222_X1 U9350 ( .A1(n7786), .A2(P1_U3086), .B1(n9484), .B2(n7785), .C1(
        n7784), .C2(n9487), .ZN(P1_U3329) );
  INV_X1 U9351 ( .A(n7787), .ZN(n7789) );
  NAND2_X1 U9352 ( .A1(n7789), .A2(n7788), .ZN(n7794) );
  XNOR2_X1 U9353 ( .A(n8119), .B(n7183), .ZN(n7851) );
  NAND2_X1 U9354 ( .A1(n7854), .A2(n8005), .ZN(n7804) );
  AOI21_X1 U9355 ( .B1(n7793), .B2(n7794), .A(n7851), .ZN(n7803) );
  INV_X1 U9356 ( .A(n7795), .ZN(n7796) );
  NAND2_X1 U9357 ( .A1(n8077), .A2(n7796), .ZN(n7799) );
  AOI21_X1 U9358 ( .B1(n8078), .B2(n8317), .A(n7797), .ZN(n7798) );
  OAI211_X1 U9359 ( .C1(n8619), .C2(n8081), .A(n7799), .B(n7798), .ZN(n7800)
         );
  AOI21_X1 U9360 ( .B1(n7801), .B2(n8089), .A(n7800), .ZN(n7802) );
  OAI21_X1 U9361 ( .B1(n7804), .B2(n7803), .A(n7802), .ZN(P2_U3176) );
  INV_X1 U9362 ( .A(n7805), .ZN(n9483) );
  AOI21_X1 U9363 ( .B1(n8774), .B2(P1_DATAO_REG_27__SCAN_IN), .A(n7806), .ZN(
        n7807) );
  OAI21_X1 U9364 ( .B1(n9483), .B2(n8777), .A(n7807), .ZN(P2_U3268) );
  NAND2_X1 U9365 ( .A1(n7809), .A2(n7808), .ZN(n7810) );
  XNOR2_X1 U9366 ( .A(n7811), .B(n7810), .ZN(n7818) );
  AOI22_X1 U9367 ( .A1(n8927), .A2(n7812), .B1(n8945), .B2(n8955), .ZN(n7813)
         );
  NAND2_X1 U9368 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n9627) );
  OAI211_X1 U9369 ( .C1(n7814), .C2(n8940), .A(n7813), .B(n9627), .ZN(n7815)
         );
  AOI21_X1 U9370 ( .B1(n7816), .B2(n8928), .A(n7815), .ZN(n7817) );
  OAI21_X1 U9371 ( .B1(n7818), .B2(n8920), .A(n7817), .ZN(P1_U3236) );
  INV_X1 U9372 ( .A(n7824), .ZN(n9406) );
  XNOR2_X1 U9373 ( .A(n9098), .B(n7827), .ZN(n9413) );
  OR2_X2 U9374 ( .A1(n7836), .A2(n8861), .ZN(n7834) );
  AOI211_X1 U9375 ( .C1(n9096), .C2(n7834), .A(n9792), .B(n9290), .ZN(n9410)
         );
  INV_X1 U9376 ( .A(n9096), .ZN(n9408) );
  NOR2_X1 U9377 ( .A1(n9408), .A2(n9273), .ZN(n7826) );
  AOI22_X1 U9378 ( .A1(n9293), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n7821), .B2(
        n9291), .ZN(n7823) );
  NAND2_X1 U9379 ( .A1(n9294), .A2(n9405), .ZN(n7822) );
  OAI211_X1 U9380 ( .C1(n7824), .C2(n9297), .A(n7823), .B(n7822), .ZN(n7825)
         );
  AOI211_X1 U9381 ( .C1(n9410), .C2(n9284), .A(n7826), .B(n7825), .ZN(n7830)
         );
  XNOR2_X1 U9382 ( .A(n7828), .B(n7827), .ZN(n9411) );
  NAND2_X1 U9383 ( .A1(n9411), .A2(n9304), .ZN(n7829) );
  OAI211_X1 U9384 ( .C1(n9413), .C2(n9306), .A(n7830), .B(n7829), .ZN(P1_U3276) );
  AOI21_X1 U9385 ( .B1(n7833), .B2(n7831), .A(n4439), .ZN(n9418) );
  XOR2_X1 U9386 ( .A(n7833), .B(n7832), .Z(n9420) );
  NAND2_X1 U9387 ( .A1(n9420), .A2(n9212), .ZN(n7842) );
  INV_X1 U9388 ( .A(n7834), .ZN(n7835) );
  AOI211_X1 U9389 ( .C1(n8861), .C2(n7836), .A(n9792), .B(n7835), .ZN(n9416)
         );
  INV_X1 U9390 ( .A(n8861), .ZN(n9466) );
  NOR2_X1 U9391 ( .A1(n9466), .A2(n9273), .ZN(n7840) );
  AOI22_X1 U9392 ( .A1(n9293), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n8858), .B2(
        n9291), .ZN(n7838) );
  NAND2_X1 U9393 ( .A1(n9294), .A2(n9397), .ZN(n7837) );
  OAI211_X1 U9394 ( .C1(n9425), .C2(n9297), .A(n7838), .B(n7837), .ZN(n7839)
         );
  AOI211_X1 U9395 ( .C1(n9416), .C2(n9284), .A(n7840), .B(n7839), .ZN(n7841)
         );
  OAI211_X1 U9396 ( .C1(n9418), .C2(n9173), .A(n7842), .B(n7841), .ZN(P1_U3277) );
  INV_X1 U9397 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n7847) );
  OAI211_X1 U9398 ( .C1(n7845), .C2(n9760), .A(n7844), .B(n7843), .ZN(n7846)
         );
  INV_X1 U9399 ( .A(n7846), .ZN(n7849) );
  MUX2_X1 U9400 ( .A(n7847), .B(n7849), .S(n9798), .Z(n7848) );
  OAI21_X1 U9401 ( .B1(n8949), .B2(n9465), .A(n7848), .ZN(P1_U3498) );
  INV_X1 U9402 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n9677) );
  MUX2_X1 U9403 ( .A(n9677), .B(n7849), .S(n9813), .Z(n7850) );
  OAI21_X1 U9404 ( .B1(n8949), .B2(n9423), .A(n7850), .ZN(P1_U3537) );
  NAND2_X1 U9405 ( .A1(n7790), .A2(n8316), .ZN(n7853) );
  XNOR2_X1 U9406 ( .A(n9912), .B(n7934), .ZN(n7892) );
  XNOR2_X1 U9407 ( .A(n7892), .B(n8619), .ZN(n7894) );
  XNOR2_X1 U9408 ( .A(n7895), .B(n7894), .ZN(n7862) );
  INV_X1 U9409 ( .A(n7855), .ZN(n7856) );
  NAND2_X1 U9410 ( .A1(n8077), .A2(n7856), .ZN(n7859) );
  AOI21_X1 U9411 ( .B1(n8078), .B2(n8316), .A(n7857), .ZN(n7858) );
  OAI211_X1 U9412 ( .C1(n8607), .C2(n8081), .A(n7859), .B(n7858), .ZN(n7860)
         );
  AOI21_X1 U9413 ( .B1(n9912), .B2(n8089), .A(n7860), .ZN(n7861) );
  OAI21_X1 U9414 ( .B1(n7862), .B2(n8084), .A(n7861), .ZN(P2_U3164) );
  OAI222_X1 U9415 ( .A1(n9487), .A2(n7865), .B1(n9481), .B2(n7864), .C1(n7863), 
        .C2(P1_U3086), .ZN(P1_U3336) );
  INV_X1 U9416 ( .A(n7866), .ZN(n8773) );
  OAI222_X1 U9417 ( .A1(n9487), .A2(n7868), .B1(P1_U3086), .B2(n7867), .C1(
        n9484), .C2(n8773), .ZN(P1_U3326) );
  INV_X1 U9418 ( .A(n8243), .ZN(n8234) );
  XOR2_X1 U9419 ( .A(n8128), .B(n7869), .Z(n7886) );
  INV_X1 U9420 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n7875) );
  INV_X1 U9421 ( .A(n8128), .ZN(n7871) );
  XNOR2_X1 U9422 ( .A(n7870), .B(n7871), .ZN(n7874) );
  NAND2_X1 U9423 ( .A1(n8563), .A2(n8591), .ZN(n7872) );
  OAI21_X1 U9424 ( .B1(n8311), .B2(n8622), .A(n7872), .ZN(n7873) );
  AOI21_X1 U9425 ( .B1(n7874), .B2(n8596), .A(n7873), .ZN(n7881) );
  MUX2_X1 U9426 ( .A(n7875), .B(n7881), .S(n9914), .Z(n7877) );
  NAND2_X1 U9427 ( .A1(n7975), .A2(n8758), .ZN(n7876) );
  OAI211_X1 U9428 ( .C1(n7886), .C2(n8753), .A(n7877), .B(n7876), .ZN(P2_U3446) );
  MUX2_X1 U9429 ( .A(n7878), .B(n7881), .S(n9929), .Z(n7880) );
  NAND2_X1 U9430 ( .A1(n7975), .A2(n8675), .ZN(n7879) );
  OAI211_X1 U9431 ( .C1(n8673), .C2(n7886), .A(n7880), .B(n7879), .ZN(P2_U3478) );
  MUX2_X1 U9432 ( .A(n7882), .B(n7881), .S(n8633), .Z(n7885) );
  INV_X1 U9433 ( .A(n7973), .ZN(n7883) );
  AOI22_X1 U9434 ( .A1(n7975), .A2(n8600), .B1(n8599), .B2(n7883), .ZN(n7884)
         );
  OAI211_X1 U9435 ( .C1(n7886), .C2(n8603), .A(n7885), .B(n7884), .ZN(P2_U3214) );
  OAI222_X1 U9436 ( .A1(n9487), .A2(n7888), .B1(n9481), .B2(n7887), .C1(
        P1_U3086), .C2(n5834), .ZN(P1_U3333) );
  INV_X1 U9437 ( .A(n7889), .ZN(n8778) );
  OAI222_X1 U9438 ( .A1(n9487), .A2(n7890), .B1(P1_U3086), .B2(n9542), .C1(
        n9484), .C2(n8778), .ZN(P1_U3327) );
  XNOR2_X1 U9439 ( .A(n7891), .B(n7183), .ZN(n7906) );
  XNOR2_X1 U9440 ( .A(n8744), .B(n7934), .ZN(n7902) );
  INV_X1 U9441 ( .A(n7902), .ZN(n7903) );
  XNOR2_X1 U9442 ( .A(n8623), .B(n7934), .ZN(n7896) );
  NAND2_X1 U9443 ( .A1(n7896), .A2(n8314), .ZN(n8037) );
  XNOR2_X1 U9444 ( .A(n8609), .B(n7934), .ZN(n7897) );
  XNOR2_X1 U9445 ( .A(n7897), .B(n8592), .ZN(n7957) );
  XNOR2_X1 U9446 ( .A(n8757), .B(n7934), .ZN(n7898) );
  XNOR2_X1 U9447 ( .A(n7898), .B(n8313), .ZN(n8086) );
  XNOR2_X1 U9448 ( .A(n8750), .B(n7934), .ZN(n7900) );
  XNOR2_X1 U9449 ( .A(n7900), .B(n8082), .ZN(n7993) );
  INV_X1 U9450 ( .A(n7900), .ZN(n7901) );
  NAND2_X1 U9451 ( .A1(n7901), .A2(n8082), .ZN(n8002) );
  XNOR2_X1 U9452 ( .A(n7902), .B(n8312), .ZN(n8003) );
  XNOR2_X1 U9453 ( .A(n8063), .B(n7934), .ZN(n7904) );
  XNOR2_X1 U9454 ( .A(n7904), .B(n8563), .ZN(n8058) );
  XNOR2_X1 U9455 ( .A(n7906), .B(n8547), .ZN(n7970) );
  XNOR2_X1 U9456 ( .A(n8733), .B(n7934), .ZN(n7907) );
  XNOR2_X1 U9457 ( .A(n7907), .B(n8311), .ZN(n8029) );
  INV_X1 U9458 ( .A(n7907), .ZN(n7908) );
  XNOR2_X1 U9459 ( .A(n8727), .B(n7934), .ZN(n7912) );
  XNOR2_X1 U9460 ( .A(n7912), .B(n8538), .ZN(n7980) );
  INV_X1 U9461 ( .A(n7980), .ZN(n7911) );
  NAND2_X1 U9462 ( .A1(n7978), .A2(n7911), .ZN(n7915) );
  INV_X1 U9463 ( .A(n7912), .ZN(n7913) );
  NAND2_X1 U9464 ( .A1(n7913), .A2(n8030), .ZN(n7914) );
  INV_X1 U9465 ( .A(n8048), .ZN(n7917) );
  XNOR2_X1 U9466 ( .A(n8721), .B(n7934), .ZN(n7918) );
  XNOR2_X1 U9467 ( .A(n7918), .B(n8525), .ZN(n8047) );
  INV_X1 U9468 ( .A(n8047), .ZN(n7916) );
  NAND2_X1 U9469 ( .A1(n7918), .A2(n8525), .ZN(n7919) );
  XNOR2_X1 U9470 ( .A(n8709), .B(n7934), .ZN(n8019) );
  XNOR2_X1 U9471 ( .A(n8715), .B(n7183), .ZN(n7922) );
  OAI22_X1 U9472 ( .A1(n8019), .A2(n8018), .B1(n8485), .B2(n7922), .ZN(n7920)
         );
  INV_X1 U9473 ( .A(n7920), .ZN(n7921) );
  OAI21_X1 U9474 ( .B1(n8016), .B2(n8511), .A(n8499), .ZN(n7924) );
  NOR3_X1 U9475 ( .A1(n8016), .A2(n8511), .A3(n8499), .ZN(n7923) );
  AOI21_X1 U9476 ( .B1(n8019), .B2(n7924), .A(n7923), .ZN(n7925) );
  XNOR2_X1 U9477 ( .A(n8704), .B(n7934), .ZN(n7927) );
  XNOR2_X1 U9478 ( .A(n7927), .B(n8486), .ZN(n7987) );
  INV_X1 U9479 ( .A(n7927), .ZN(n7928) );
  NAND2_X1 U9480 ( .A1(n7928), .A2(n8486), .ZN(n7929) );
  XNOR2_X1 U9481 ( .A(n8698), .B(n7934), .ZN(n7930) );
  NAND2_X1 U9482 ( .A1(n7930), .A2(n8474), .ZN(n8066) );
  INV_X1 U9483 ( .A(n7930), .ZN(n7931) );
  NAND2_X1 U9484 ( .A1(n7931), .A2(n8455), .ZN(n8067) );
  XNOR2_X1 U9485 ( .A(n8692), .B(n7183), .ZN(n7932) );
  XNOR2_X1 U9486 ( .A(n7932), .B(n8465), .ZN(n7950) );
  INV_X1 U9487 ( .A(n7932), .ZN(n7933) );
  OAI22_X1 U9488 ( .A1(n7951), .A2(n7950), .B1(n8072), .B2(n7933), .ZN(n7936)
         );
  XNOR2_X1 U9489 ( .A(n8445), .B(n7934), .ZN(n7935) );
  XNOR2_X1 U9490 ( .A(n7936), .B(n7935), .ZN(n7941) );
  INV_X1 U9491 ( .A(n8438), .ZN(n8274) );
  AOI22_X1 U9492 ( .A1(n8465), .A2(n8078), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3151), .ZN(n7938) );
  NAND2_X1 U9493 ( .A1(n8077), .A2(n8444), .ZN(n7937) );
  OAI211_X1 U9494 ( .C1(n8274), .C2(n8081), .A(n7938), .B(n7937), .ZN(n7939)
         );
  AOI21_X1 U9495 ( .B1(n8687), .B2(n8089), .A(n7939), .ZN(n7940) );
  OAI21_X1 U9496 ( .B1(n7941), .B2(n8084), .A(n7940), .ZN(P2_U3160) );
  NAND2_X1 U9497 ( .A1(n8272), .A2(n8600), .ZN(n7944) );
  NAND2_X1 U9498 ( .A1(n7943), .A2(n8599), .ZN(n8430) );
  OAI211_X1 U9499 ( .C1(n8633), .C2(n7945), .A(n7944), .B(n8430), .ZN(n7946)
         );
  AOI21_X1 U9500 ( .B1(n7948), .B2(n7947), .A(n7946), .ZN(n7949) );
  OAI21_X1 U9501 ( .B1(n7942), .B2(n8582), .A(n7949), .ZN(P2_U3204) );
  XNOR2_X1 U9502 ( .A(n7951), .B(n7950), .ZN(n7956) );
  AOI22_X1 U9503 ( .A1(n8310), .A2(n8009), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3151), .ZN(n7953) );
  NAND2_X1 U9504 ( .A1(n8077), .A2(n8457), .ZN(n7952) );
  OAI211_X1 U9505 ( .C1(n8455), .C2(n8031), .A(n7953), .B(n7952), .ZN(n7954)
         );
  AOI21_X1 U9506 ( .B1(n8458), .B2(n8089), .A(n7954), .ZN(n7955) );
  OAI21_X1 U9507 ( .B1(n7956), .B2(n8084), .A(n7955), .ZN(P2_U3154) );
  XOR2_X1 U9508 ( .A(n7958), .B(n7957), .Z(n7963) );
  AOI22_X1 U9509 ( .A1(n8009), .A2(n8313), .B1(P2_REG3_REG_14__SCAN_IN), .B2(
        P2_U3151), .ZN(n7960) );
  NAND2_X1 U9510 ( .A1(n8078), .A2(n8314), .ZN(n7959) );
  OAI211_X1 U9511 ( .C1(n8061), .C2(n8610), .A(n7960), .B(n7959), .ZN(n7961)
         );
  AOI21_X1 U9512 ( .B1(n8609), .B2(n8089), .A(n7961), .ZN(n7962) );
  OAI21_X1 U9513 ( .B1(n7963), .B2(n8084), .A(n7962), .ZN(P2_U3155) );
  XNOR2_X1 U9514 ( .A(n8015), .B(n8016), .ZN(n8017) );
  XNOR2_X1 U9515 ( .A(n8017), .B(n8485), .ZN(n7968) );
  AOI22_X1 U9516 ( .A1(n8078), .A2(n8525), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3151), .ZN(n7965) );
  NAND2_X1 U9517 ( .A1(n8077), .A2(n8502), .ZN(n7964) );
  OAI211_X1 U9518 ( .C1(n8018), .C2(n8081), .A(n7965), .B(n7964), .ZN(n7966)
         );
  AOI21_X1 U9519 ( .B1(n8715), .B2(n8089), .A(n7966), .ZN(n7967) );
  OAI21_X1 U9520 ( .B1(n7968), .B2(n8084), .A(n7967), .ZN(P2_U3156) );
  XOR2_X1 U9521 ( .A(n7970), .B(n7969), .Z(n7977) );
  OAI22_X1 U9522 ( .A1(n8081), .A2(n8311), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10045), .ZN(n7971) );
  AOI21_X1 U9523 ( .B1(n8078), .B2(n8563), .A(n7971), .ZN(n7972) );
  OAI21_X1 U9524 ( .B1(n7973), .B2(n8061), .A(n7972), .ZN(n7974) );
  AOI21_X1 U9525 ( .B1(n7975), .B2(n8089), .A(n7974), .ZN(n7976) );
  OAI21_X1 U9526 ( .B1(n7977), .B2(n8084), .A(n7976), .ZN(P2_U3159) );
  XOR2_X1 U9527 ( .A(n7980), .B(n7979), .Z(n7985) );
  AOI22_X1 U9528 ( .A1(n8009), .A2(n8525), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3151), .ZN(n7982) );
  NAND2_X1 U9529 ( .A1(n8077), .A2(n8528), .ZN(n7981) );
  OAI211_X1 U9530 ( .C1(n8311), .C2(n8031), .A(n7982), .B(n7981), .ZN(n7983)
         );
  AOI21_X1 U9531 ( .B1(n8727), .B2(n8089), .A(n7983), .ZN(n7984) );
  OAI21_X1 U9532 ( .B1(n7985), .B2(n8084), .A(n7984), .ZN(P2_U3163) );
  XOR2_X1 U9533 ( .A(n7987), .B(n7986), .Z(n7992) );
  AOI22_X1 U9534 ( .A1(n8009), .A2(n8474), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3151), .ZN(n7989) );
  NAND2_X1 U9535 ( .A1(n8077), .A2(n8478), .ZN(n7988) );
  OAI211_X1 U9536 ( .C1(n8018), .C2(n8031), .A(n7989), .B(n7988), .ZN(n7990)
         );
  AOI21_X1 U9537 ( .B1(n8704), .B2(n8089), .A(n7990), .ZN(n7991) );
  OAI21_X1 U9538 ( .B1(n7992), .B2(n8084), .A(n7991), .ZN(P2_U3165) );
  INV_X1 U9539 ( .A(n8750), .ZN(n8001) );
  OAI21_X1 U9540 ( .B1(n7994), .B2(n7993), .A(n8004), .ZN(n7995) );
  NAND2_X1 U9541 ( .A1(n7995), .A2(n8005), .ZN(n8000) );
  INV_X1 U9542 ( .A(n7996), .ZN(n8584) );
  AOI22_X1 U9543 ( .A1(n8009), .A2(n8312), .B1(P2_REG3_REG_16__SCAN_IN), .B2(
        P2_U3151), .ZN(n7997) );
  OAI21_X1 U9544 ( .B1(n8608), .B2(n8031), .A(n7997), .ZN(n7998) );
  AOI21_X1 U9545 ( .B1(n8584), .B2(n8077), .A(n7998), .ZN(n7999) );
  OAI211_X1 U9546 ( .C1(n8001), .C2(n8055), .A(n8000), .B(n7999), .ZN(P2_U3166) );
  INV_X1 U9547 ( .A(n8744), .ZN(n8014) );
  AND3_X1 U9548 ( .A1(n8004), .A2(n8003), .A3(n8002), .ZN(n8006) );
  OAI21_X1 U9549 ( .B1(n8007), .B2(n8006), .A(n8005), .ZN(n8013) );
  INV_X1 U9550 ( .A(n8008), .ZN(n8566) );
  AOI22_X1 U9551 ( .A1(n8009), .A2(n8563), .B1(P2_REG3_REG_17__SCAN_IN), .B2(
        P2_U3151), .ZN(n8010) );
  OAI21_X1 U9552 ( .B1(n8082), .B2(n8031), .A(n8010), .ZN(n8011) );
  AOI21_X1 U9553 ( .B1(n8566), .B2(n8077), .A(n8011), .ZN(n8012) );
  OAI211_X1 U9554 ( .C1(n8014), .C2(n8055), .A(n8013), .B(n8012), .ZN(P2_U3168) );
  OAI22_X1 U9555 ( .A1(n8017), .A2(n8511), .B1(n8016), .B2(n8015), .ZN(n8021)
         );
  XNOR2_X1 U9556 ( .A(n8019), .B(n8018), .ZN(n8020) );
  XNOR2_X1 U9557 ( .A(n8021), .B(n8020), .ZN(n8027) );
  OAI22_X1 U9558 ( .A1(n8081), .A2(n8486), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10055), .ZN(n8023) );
  NOR2_X1 U9559 ( .A1(n8031), .A2(n8485), .ZN(n8022) );
  AOI211_X1 U9560 ( .C1(n8488), .C2(n8077), .A(n8023), .B(n8022), .ZN(n8026)
         );
  NAND2_X1 U9561 ( .A1(n8024), .A2(n8089), .ZN(n8025) );
  OAI211_X1 U9562 ( .C1(n8027), .C2(n8084), .A(n8026), .B(n8025), .ZN(P2_U3169) );
  XOR2_X1 U9563 ( .A(n8029), .B(n8028), .Z(n8036) );
  INV_X1 U9564 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n10113) );
  OAI22_X1 U9565 ( .A1(n8081), .A2(n8030), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10113), .ZN(n8033) );
  NOR2_X1 U9566 ( .A1(n8031), .A2(n8547), .ZN(n8032) );
  AOI211_X1 U9567 ( .C1(n8541), .C2(n8077), .A(n8033), .B(n8032), .ZN(n8035)
         );
  NAND2_X1 U9568 ( .A1(n8733), .A2(n8089), .ZN(n8034) );
  OAI211_X1 U9569 ( .C1(n8036), .C2(n8084), .A(n8035), .B(n8034), .ZN(P2_U3173) );
  NAND2_X1 U9570 ( .A1(n4446), .A2(n8037), .ZN(n8038) );
  XNOR2_X1 U9571 ( .A(n8039), .B(n8038), .ZN(n8046) );
  INV_X1 U9572 ( .A(n8625), .ZN(n8040) );
  NAND2_X1 U9573 ( .A1(n8077), .A2(n8040), .ZN(n8043) );
  AOI21_X1 U9574 ( .B1(n8078), .B2(n8315), .A(n8041), .ZN(n8042) );
  OAI211_X1 U9575 ( .C1(n8621), .C2(n8081), .A(n8043), .B(n8042), .ZN(n8044)
         );
  AOI21_X1 U9576 ( .B1(n8623), .B2(n8089), .A(n8044), .ZN(n8045) );
  OAI21_X1 U9577 ( .B1(n8046), .B2(n8084), .A(n8045), .ZN(P2_U3174) );
  INV_X1 U9578 ( .A(n8721), .ZN(n8056) );
  AOI21_X1 U9579 ( .B1(n8048), .B2(n8047), .A(n8084), .ZN(n8050) );
  NAND2_X1 U9580 ( .A1(n8050), .A2(n8049), .ZN(n8054) );
  AOI22_X1 U9581 ( .A1(n8078), .A2(n8538), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3151), .ZN(n8051) );
  OAI21_X1 U9582 ( .B1(n8485), .B2(n8081), .A(n8051), .ZN(n8052) );
  AOI21_X1 U9583 ( .B1(n8514), .B2(n8077), .A(n8052), .ZN(n8053) );
  OAI211_X1 U9584 ( .C1(n8056), .C2(n8055), .A(n8054), .B(n8053), .ZN(P2_U3175) );
  XOR2_X1 U9585 ( .A(n8058), .B(n8057), .Z(n8065) );
  NAND2_X1 U9586 ( .A1(P2_U3151), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8385) );
  OAI21_X1 U9587 ( .B1(n8081), .B2(n8547), .A(n8385), .ZN(n8059) );
  AOI21_X1 U9588 ( .B1(n8078), .B2(n8312), .A(n8059), .ZN(n8060) );
  OAI21_X1 U9589 ( .B1(n8551), .B2(n8061), .A(n8060), .ZN(n8062) );
  AOI21_X1 U9590 ( .B1(n8063), .B2(n8089), .A(n8062), .ZN(n8064) );
  OAI21_X1 U9591 ( .B1(n8065), .B2(n8084), .A(n8064), .ZN(P2_U3178) );
  NAND2_X1 U9592 ( .A1(n8067), .A2(n8066), .ZN(n8068) );
  XNOR2_X1 U9593 ( .A(n8069), .B(n8068), .ZN(n8075) );
  AOI22_X1 U9594 ( .A1(n8078), .A2(n8464), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3151), .ZN(n8071) );
  NAND2_X1 U9595 ( .A1(n8077), .A2(n8468), .ZN(n8070) );
  OAI211_X1 U9596 ( .C1(n8072), .C2(n8081), .A(n8071), .B(n8070), .ZN(n8073)
         );
  AOI21_X1 U9597 ( .B1(n8698), .B2(n8089), .A(n8073), .ZN(n8074) );
  OAI21_X1 U9598 ( .B1(n8075), .B2(n8084), .A(n8074), .ZN(P2_U3180) );
  INV_X1 U9599 ( .A(n8076), .ZN(n8598) );
  NAND2_X1 U9600 ( .A1(n8077), .A2(n8598), .ZN(n8080) );
  AND2_X1 U9601 ( .A1(P2_U3151), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8348) );
  AOI21_X1 U9602 ( .B1(n8078), .B2(n8592), .A(n8348), .ZN(n8079) );
  OAI211_X1 U9603 ( .C1(n8082), .C2(n8081), .A(n8080), .B(n8079), .ZN(n8088)
         );
  AOI211_X1 U9604 ( .C1(n8086), .C2(n8085), .A(n8084), .B(n8083), .ZN(n8087)
         );
  AOI211_X1 U9605 ( .C1(n8757), .C2(n8089), .A(n8088), .B(n8087), .ZN(n8090)
         );
  INV_X1 U9606 ( .A(n8090), .ZN(P2_U3181) );
  INV_X1 U9607 ( .A(n8091), .ZN(n8096) );
  NOR2_X1 U9608 ( .A1(n8272), .A2(n8274), .ZN(n8282) );
  INV_X1 U9609 ( .A(n8282), .ZN(n8095) );
  NAND2_X1 U9610 ( .A1(n8768), .A2(n8097), .ZN(n8093) );
  NAND2_X1 U9611 ( .A1(n6192), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n8092) );
  INV_X1 U9612 ( .A(n8309), .ZN(n8285) );
  NAND2_X1 U9613 ( .A1(n8433), .A2(n8285), .ZN(n8102) );
  NAND2_X1 U9614 ( .A1(n8272), .A2(n8274), .ZN(n8094) );
  NAND2_X1 U9615 ( .A1(n8102), .A2(n8094), .ZN(n8288) );
  AOI21_X1 U9616 ( .B1(n8096), .B2(n8095), .A(n8288), .ZN(n8101) );
  NAND2_X1 U9617 ( .A1(n8763), .A2(n8097), .ZN(n8099) );
  NAND2_X1 U9618 ( .A1(n6192), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n8098) );
  OAI21_X1 U9619 ( .B1(n8429), .B2(n8433), .A(n8432), .ZN(n8100) );
  NOR2_X1 U9620 ( .A1(n8433), .A2(n8285), .ZN(n8281) );
  AOI22_X1 U9621 ( .A1(n8101), .A2(n8100), .B1(n8281), .B2(n8679), .ZN(n8301)
         );
  INV_X1 U9622 ( .A(n8102), .ZN(n8133) );
  INV_X1 U9623 ( .A(n8264), .ZN(n8103) );
  INV_X1 U9624 ( .A(n8489), .ZN(n8105) );
  NOR2_X1 U9625 ( .A1(n8252), .A2(n8105), .ZN(n8498) );
  INV_X1 U9626 ( .A(n8521), .ZN(n8517) );
  INV_X1 U9627 ( .A(n8535), .ZN(n8129) );
  INV_X1 U9628 ( .A(n8233), .ZN(n8106) );
  NOR2_X1 U9629 ( .A1(n8231), .A2(n8106), .ZN(n8549) );
  NOR2_X1 U9630 ( .A1(n8108), .A2(n8107), .ZN(n8113) );
  NOR2_X1 U9631 ( .A1(n8110), .A2(n8109), .ZN(n8112) );
  NAND4_X1 U9632 ( .A1(n8113), .A2(n8112), .A3(n8111), .A4(n8158), .ZN(n8117)
         );
  INV_X1 U9633 ( .A(n8114), .ZN(n8115) );
  NOR3_X1 U9634 ( .A1(n8117), .A2(n8116), .A3(n8115), .ZN(n8121) );
  INV_X1 U9635 ( .A(n8118), .ZN(n8120) );
  NAND4_X1 U9636 ( .A1(n8121), .A2(n8120), .A3(n8119), .A4(n8179), .ZN(n8123)
         );
  NOR2_X1 U9637 ( .A1(n8123), .A2(n8122), .ZN(n8125) );
  INV_X1 U9638 ( .A(n8210), .ZN(n8124) );
  NAND4_X1 U9639 ( .A1(n8612), .A2(n8206), .A3(n8125), .A4(n8629), .ZN(n8126)
         );
  NOR4_X1 U9640 ( .A1(n8557), .A2(n8222), .A3(n8589), .A4(n8126), .ZN(n8127)
         );
  NAND4_X1 U9641 ( .A1(n8129), .A2(n8128), .A3(n8549), .A4(n8127), .ZN(n8130)
         );
  NAND3_X1 U9642 ( .A1(n8492), .A2(n8498), .A3(n4394), .ZN(n8131) );
  OR3_X1 U9643 ( .A1(n8462), .A2(n8479), .A3(n8131), .ZN(n8132) );
  NOR4_X1 U9644 ( .A1(n8133), .A2(n8445), .A3(n8451), .A4(n8132), .ZN(n8136)
         );
  INV_X1 U9645 ( .A(n8281), .ZN(n8135) );
  NAND2_X1 U9646 ( .A1(n8432), .A2(n8429), .ZN(n8296) );
  NAND4_X1 U9647 ( .A1(n8136), .A2(n8135), .A3(n8296), .A4(n8134), .ZN(n8140)
         );
  NAND2_X1 U9648 ( .A1(n8679), .A2(n8137), .ZN(n8293) );
  INV_X1 U9649 ( .A(n8293), .ZN(n8138) );
  AOI21_X1 U9650 ( .B1(n8140), .B2(n8139), .A(n8138), .ZN(n8299) );
  INV_X1 U9651 ( .A(n8253), .ZN(n8241) );
  NOR2_X1 U9652 ( .A1(n8236), .A2(n8289), .ZN(n8141) );
  OAI21_X1 U9653 ( .B1(n8252), .B2(n8141), .A(n8253), .ZN(n8142) );
  OAI211_X1 U9654 ( .C1(n8284), .C2(n8250), .A(n8142), .B(n8254), .ZN(n8240)
         );
  NAND2_X1 U9655 ( .A1(n8167), .A2(n8143), .ZN(n8146) );
  NAND2_X1 U9656 ( .A1(n8160), .A2(n8144), .ZN(n8145) );
  MUX2_X1 U9657 ( .A(n8146), .B(n8145), .S(n8289), .Z(n8157) );
  NAND2_X1 U9658 ( .A1(n8148), .A2(n8147), .ZN(n8153) );
  NAND2_X1 U9659 ( .A1(n8153), .A2(n8149), .ZN(n8150) );
  NAND3_X1 U9660 ( .A1(n8152), .A2(n8151), .A3(n8150), .ZN(n8155) );
  AOI21_X1 U9661 ( .B1(n8153), .B2(n6489), .A(n8284), .ZN(n8154) );
  OR2_X1 U9662 ( .A1(n8157), .A2(n8156), .ZN(n8159) );
  NAND2_X1 U9663 ( .A1(n8159), .A2(n8158), .ZN(n8171) );
  INV_X1 U9664 ( .A(n8160), .ZN(n8162) );
  OAI211_X1 U9665 ( .C1(n8171), .C2(n8162), .A(n8174), .B(n8161), .ZN(n8166)
         );
  NAND2_X1 U9666 ( .A1(n8172), .A2(n8168), .ZN(n8164) );
  NAND2_X1 U9667 ( .A1(n8164), .A2(n8163), .ZN(n8165) );
  INV_X1 U9668 ( .A(n8167), .ZN(n8170) );
  NAND2_X1 U9669 ( .A1(n8323), .A2(n9875), .ZN(n8169) );
  OAI211_X1 U9670 ( .C1(n8171), .C2(n8170), .A(n8169), .B(n8168), .ZN(n8175)
         );
  INV_X1 U9671 ( .A(n8172), .ZN(n8173) );
  AOI21_X1 U9672 ( .B1(n8175), .B2(n8174), .A(n8173), .ZN(n8176) );
  NAND2_X1 U9673 ( .A1(n8187), .A2(n8188), .ZN(n8178) );
  NAND2_X1 U9674 ( .A1(n8183), .A2(n8181), .ZN(n8177) );
  MUX2_X1 U9675 ( .A(n8178), .B(n8177), .S(n8289), .Z(n8185) );
  INV_X1 U9676 ( .A(n8185), .ZN(n8191) );
  AND2_X1 U9677 ( .A1(n8181), .A2(n8180), .ZN(n8184) );
  INV_X1 U9678 ( .A(n8182), .ZN(n8200) );
  OAI211_X1 U9679 ( .C1(n8185), .C2(n8184), .A(n8200), .B(n8183), .ZN(n8186)
         );
  INV_X1 U9680 ( .A(n8186), .ZN(n8193) );
  OAI21_X1 U9681 ( .B1(n9884), .B2(n8320), .A(n8187), .ZN(n8190) );
  NAND2_X1 U9682 ( .A1(n8195), .A2(n8188), .ZN(n8189) );
  AOI21_X1 U9683 ( .B1(n8191), .B2(n8190), .A(n8189), .ZN(n8192) );
  MUX2_X1 U9684 ( .A(n8193), .B(n8192), .S(n8289), .Z(n8194) );
  NAND2_X1 U9685 ( .A1(n8196), .A2(n8199), .ZN(n8198) );
  NAND2_X1 U9686 ( .A1(n8198), .A2(n8197), .ZN(n8205) );
  AND2_X1 U9687 ( .A1(n8200), .A2(n8199), .ZN(n8202) );
  AOI21_X1 U9688 ( .B1(n8203), .B2(n8202), .A(n8201), .ZN(n8204) );
  MUX2_X1 U9689 ( .A(n8208), .B(n8207), .S(n8289), .Z(n8209) );
  NOR2_X1 U9690 ( .A1(n8211), .A2(n8210), .ZN(n8216) );
  MUX2_X1 U9691 ( .A(n8314), .B(n8623), .S(n8289), .Z(n8215) );
  INV_X1 U9692 ( .A(n8212), .ZN(n8213) );
  OAI22_X1 U9693 ( .A1(n8216), .A2(n8215), .B1(n8214), .B2(n8213), .ZN(n8221)
         );
  INV_X1 U9694 ( .A(n8217), .ZN(n8218) );
  MUX2_X1 U9695 ( .A(n8219), .B(n8218), .S(n8289), .Z(n8220) );
  AOI211_X1 U9696 ( .C1(n8221), .C2(n8612), .A(n8220), .B(n8589), .ZN(n8229)
         );
  INV_X1 U9697 ( .A(n8222), .ZN(n8574) );
  MUX2_X1 U9698 ( .A(n8223), .B(n8570), .S(n8284), .Z(n8224) );
  NAND2_X1 U9699 ( .A1(n8574), .A2(n8224), .ZN(n8228) );
  INV_X1 U9700 ( .A(n8557), .ZN(n8561) );
  MUX2_X1 U9701 ( .A(n8226), .B(n8225), .S(n8289), .Z(n8227) );
  NAND3_X1 U9702 ( .A1(n8244), .A2(n8245), .A3(n8234), .ZN(n8235) );
  NAND3_X1 U9703 ( .A1(n8235), .A2(n8248), .A3(n8242), .ZN(n8238) );
  INV_X1 U9704 ( .A(n8236), .ZN(n8237) );
  AOI211_X1 U9705 ( .C1(n8238), .C2(n8246), .A(n8237), .B(n8284), .ZN(n8239)
         );
  AOI211_X1 U9706 ( .C1(n8289), .C2(n8241), .A(n8240), .B(n8239), .ZN(n8258)
         );
  OAI211_X1 U9707 ( .C1(n8244), .C2(n8243), .A(n8242), .B(n8531), .ZN(n8247)
         );
  NAND3_X1 U9708 ( .A1(n8247), .A2(n8246), .A3(n8245), .ZN(n8249) );
  NAND2_X1 U9709 ( .A1(n8249), .A2(n8248), .ZN(n8251) );
  NAND4_X1 U9710 ( .A1(n8251), .A2(n8253), .A3(n8284), .A4(n8250), .ZN(n8257)
         );
  NAND2_X1 U9711 ( .A1(n8253), .A2(n8252), .ZN(n8255) );
  AOI21_X1 U9712 ( .B1(n8255), .B2(n8254), .A(n8284), .ZN(n8256) );
  INV_X1 U9713 ( .A(n8462), .ZN(n8262) );
  MUX2_X1 U9714 ( .A(n8260), .B(n8259), .S(n8284), .Z(n8261) );
  NAND2_X1 U9715 ( .A1(n8262), .A2(n8261), .ZN(n8267) );
  INV_X1 U9716 ( .A(n8451), .ZN(n8266) );
  MUX2_X1 U9717 ( .A(n8264), .B(n4699), .S(n8289), .Z(n8265) );
  MUX2_X1 U9718 ( .A(n8269), .B(n8268), .S(n8284), .Z(n8270) );
  INV_X1 U9719 ( .A(n8279), .ZN(n8277) );
  INV_X1 U9720 ( .A(n8687), .ZN(n8271) );
  MUX2_X1 U9721 ( .A(n8454), .B(n8271), .S(n8284), .Z(n8278) );
  INV_X1 U9722 ( .A(n8278), .ZN(n8276) );
  MUX2_X1 U9723 ( .A(n8289), .B(n8438), .S(n8272), .Z(n8273) );
  INV_X1 U9724 ( .A(n8280), .ZN(n8275) );
  OAI21_X1 U9725 ( .B1(n8277), .B2(n8276), .A(n8275), .ZN(n8292) );
  NOR3_X1 U9726 ( .A1(n8290), .A2(n8282), .A3(n8281), .ZN(n8283) );
  OAI21_X1 U9727 ( .B1(n8687), .B2(n8292), .A(n8283), .ZN(n8287) );
  OAI21_X1 U9728 ( .B1(n8285), .B2(n8284), .A(n8433), .ZN(n8286) );
  OAI211_X1 U9729 ( .C1(n8289), .C2(n8309), .A(n8287), .B(n8286), .ZN(n8295)
         );
  NOR3_X1 U9730 ( .A1(n8290), .A2(n8289), .A3(n8288), .ZN(n8291) );
  OAI21_X1 U9731 ( .B1(n8310), .B2(n8292), .A(n8291), .ZN(n8294) );
  NAND3_X1 U9732 ( .A1(n8295), .A2(n8294), .A3(n8293), .ZN(n8297) );
  NAND3_X1 U9733 ( .A1(n8303), .A2(n8302), .A3(n4370), .ZN(n8304) );
  OAI211_X1 U9734 ( .C1(n8305), .C2(n8307), .A(n8304), .B(P2_B_REG_SCAN_IN), 
        .ZN(n8306) );
  OAI21_X1 U9735 ( .B1(n8308), .B2(n8307), .A(n8306), .ZN(P2_U3296) );
  MUX2_X1 U9736 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n8309), .S(P2_U3893), .Z(
        P2_U3521) );
  MUX2_X1 U9737 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n8438), .S(P2_U3893), .Z(
        P2_U3520) );
  MUX2_X1 U9738 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n8310), .S(P2_U3893), .Z(
        P2_U3519) );
  MUX2_X1 U9739 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8465), .S(P2_U3893), .Z(
        P2_U3518) );
  MUX2_X1 U9740 ( .A(n8474), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8383), .Z(
        P2_U3517) );
  MUX2_X1 U9741 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8464), .S(P2_U3893), .Z(
        P2_U3516) );
  MUX2_X1 U9742 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n8499), .S(P2_U3893), .Z(
        P2_U3515) );
  MUX2_X1 U9743 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(n8511), .S(P2_U3893), .Z(
        P2_U3514) );
  MUX2_X1 U9744 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8525), .S(P2_U3893), .Z(
        P2_U3513) );
  MUX2_X1 U9745 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8538), .S(P2_U3893), .Z(
        P2_U3512) );
  INV_X1 U9746 ( .A(n8311), .ZN(n8524) );
  MUX2_X1 U9747 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8524), .S(P2_U3893), .Z(
        P2_U3511) );
  MUX2_X1 U9748 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8537), .S(P2_U3893), .Z(
        P2_U3510) );
  MUX2_X1 U9749 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n8563), .S(P2_U3893), .Z(
        P2_U3509) );
  MUX2_X1 U9750 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8312), .S(P2_U3893), .Z(
        P2_U3508) );
  MUX2_X1 U9751 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8594), .S(P2_U3893), .Z(
        P2_U3507) );
  MUX2_X1 U9752 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n8313), .S(P2_U3893), .Z(
        P2_U3506) );
  MUX2_X1 U9753 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n8592), .S(P2_U3893), .Z(
        P2_U3505) );
  MUX2_X1 U9754 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n8314), .S(P2_U3893), .Z(
        P2_U3504) );
  MUX2_X1 U9755 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n8315), .S(P2_U3893), .Z(
        P2_U3503) );
  MUX2_X1 U9756 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n8316), .S(P2_U3893), .Z(
        P2_U3502) );
  MUX2_X1 U9757 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n8317), .S(P2_U3893), .Z(
        P2_U3501) );
  MUX2_X1 U9758 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n8318), .S(P2_U3893), .Z(
        P2_U3500) );
  MUX2_X1 U9759 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n8319), .S(P2_U3893), .Z(
        P2_U3499) );
  MUX2_X1 U9760 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n8320), .S(P2_U3893), .Z(
        P2_U3498) );
  MUX2_X1 U9761 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n8321), .S(P2_U3893), .Z(
        P2_U3497) );
  MUX2_X1 U9762 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(n8322), .S(P2_U3893), .Z(
        P2_U3496) );
  MUX2_X1 U9763 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n8323), .S(P2_U3893), .Z(
        P2_U3495) );
  MUX2_X1 U9764 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(n8324), .S(P2_U3893), .Z(
        P2_U3494) );
  MUX2_X1 U9765 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(n8325), .S(P2_U3893), .Z(
        P2_U3493) );
  MUX2_X1 U9766 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n6183), .S(P2_U3893), .Z(
        P2_U3492) );
  MUX2_X1 U9767 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n8326), .S(P2_U3893), .Z(
        P2_U3491) );
  XOR2_X1 U9768 ( .A(n8328), .B(n8327), .Z(n8329) );
  AOI22_X1 U9769 ( .A1(n9845), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(n8361), .B2(
        n8329), .ZN(n8341) );
  OAI21_X1 U9770 ( .B1(n8332), .B2(n8331), .A(n8330), .ZN(n8336) );
  AOI22_X1 U9771 ( .A1(n8337), .A2(n8336), .B1(n8426), .B2(n8335), .ZN(n8340)
         );
  AOI22_X1 U9772 ( .A1(n9846), .A2(n8338), .B1(P2_U3151), .B2(
        P2_REG3_REG_2__SCAN_IN), .ZN(n8339) );
  NAND3_X1 U9773 ( .A1(n8341), .A2(n8340), .A3(n8339), .ZN(P2_U3184) );
  NOR2_X1 U9774 ( .A1(n8351), .A2(n4402), .ZN(n8343) );
  AOI22_X1 U9775 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n8354), .B1(n9828), .B2(
        n6348), .ZN(n9820) );
  NOR2_X1 U9776 ( .A1(n9821), .A2(n9820), .ZN(n9819) );
  AOI21_X1 U9777 ( .B1(n8344), .B2(n8597), .A(n8365), .ZN(n8363) );
  AOI21_X1 U9778 ( .B1(n8351), .B2(n8346), .A(n8345), .ZN(n9817) );
  MUX2_X1 U9779 ( .A(P2_REG2_REG_14__SCAN_IN), .B(P2_REG1_REG_14__SCAN_IN), 
        .S(n4370), .Z(n8347) );
  XNOR2_X1 U9780 ( .A(n8347), .B(n9828), .ZN(n9818) );
  OAI22_X1 U9781 ( .A1(n9817), .A2(n9818), .B1(n8347), .B2(n9828), .ZN(n8376)
         );
  MUX2_X1 U9782 ( .A(P2_REG2_REG_15__SCAN_IN), .B(P2_REG1_REG_15__SCAN_IN), 
        .S(n8415), .Z(n8373) );
  XNOR2_X1 U9783 ( .A(n8373), .B(n8392), .ZN(n8375) );
  XNOR2_X1 U9784 ( .A(n8376), .B(n8375), .ZN(n8360) );
  INV_X1 U9785 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n9976) );
  AOI21_X1 U9786 ( .B1(n9846), .B2(n8392), .A(n8348), .ZN(n8349) );
  OAI21_X1 U9787 ( .B1(n8387), .B2(n9976), .A(n8349), .ZN(n8359) );
  NOR2_X1 U9788 ( .A1(n8351), .A2(n8350), .ZN(n8353) );
  AOI22_X1 U9789 ( .A1(P2_REG1_REG_14__SCAN_IN), .A2(n8354), .B1(n9828), .B2(
        n6345), .ZN(n9815) );
  AOI21_X1 U9790 ( .B1(n8674), .B2(n8356), .A(n8393), .ZN(n8357) );
  NOR2_X1 U9791 ( .A1(n8357), .A2(n9860), .ZN(n8358) );
  AOI211_X1 U9792 ( .C1(n8361), .C2(n8360), .A(n8359), .B(n8358), .ZN(n8362)
         );
  OAI21_X1 U9793 ( .B1(n8363), .B2(n9856), .A(n8362), .ZN(P2_U3197) );
  NOR2_X1 U9794 ( .A1(n8392), .A2(n8364), .ZN(n8366) );
  AOI22_X1 U9795 ( .A1(P2_REG2_REG_16__SCAN_IN), .A2(n8395), .B1(n9843), .B2(
        n8583), .ZN(n9835) );
  NOR2_X1 U9796 ( .A1(n9847), .A2(n8368), .ZN(n8369) );
  NAND2_X1 U9797 ( .A1(n8370), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n8405) );
  OAI21_X1 U9798 ( .B1(n8370), .B2(P2_REG2_REG_18__SCAN_IN), .A(n8405), .ZN(
        n8371) );
  AOI21_X1 U9799 ( .B1(n8372), .B2(n8371), .A(n8407), .ZN(n8404) );
  INV_X1 U9800 ( .A(n8373), .ZN(n8374) );
  AOI22_X1 U9801 ( .A1(n8376), .A2(n8375), .B1(n8392), .B2(n8374), .ZN(n9832)
         );
  MUX2_X1 U9802 ( .A(P2_REG2_REG_16__SCAN_IN), .B(P2_REG1_REG_16__SCAN_IN), 
        .S(n4370), .Z(n8377) );
  XNOR2_X1 U9803 ( .A(n8377), .B(n9843), .ZN(n9833) );
  OAI22_X1 U9804 ( .A1(n9832), .A2(n9833), .B1(n8377), .B2(n9843), .ZN(n9851)
         );
  MUX2_X1 U9805 ( .A(P2_REG2_REG_17__SCAN_IN), .B(P2_REG1_REG_17__SCAN_IN), 
        .S(n8415), .Z(n8378) );
  XNOR2_X1 U9806 ( .A(n8378), .B(n9847), .ZN(n9852) );
  INV_X1 U9807 ( .A(n8378), .ZN(n8379) );
  AOI22_X1 U9808 ( .A1(n9851), .A2(n9852), .B1(n9847), .B2(n8379), .ZN(n8381)
         );
  MUX2_X1 U9809 ( .A(P2_REG2_REG_18__SCAN_IN), .B(P2_REG1_REG_18__SCAN_IN), 
        .S(n8415), .Z(n8380) );
  NOR2_X1 U9810 ( .A1(n8381), .A2(n8380), .ZN(n8413) );
  NAND2_X1 U9811 ( .A1(n8381), .A2(n8380), .ZN(n8411) );
  INV_X1 U9812 ( .A(n8411), .ZN(n8382) );
  NOR2_X1 U9813 ( .A1(n8413), .A2(n8382), .ZN(n8388) );
  INV_X1 U9814 ( .A(n8388), .ZN(n8384) );
  OAI21_X1 U9815 ( .B1(n8384), .B2(n8383), .A(n9844), .ZN(n8391) );
  INV_X1 U9816 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n8386) );
  OAI21_X1 U9817 ( .B1(n8387), .B2(n8386), .A(n8385), .ZN(n8390) );
  NOR3_X1 U9818 ( .A1(n8388), .A2(n8412), .A3(n9858), .ZN(n8389) );
  AOI211_X1 U9819 ( .C1(n8412), .C2(n8391), .A(n8390), .B(n8389), .ZN(n8403)
         );
  NOR2_X1 U9820 ( .A1(n8392), .A2(n4400), .ZN(n8394) );
  NOR2_X1 U9821 ( .A1(n8394), .A2(n8393), .ZN(n9831) );
  AOI22_X1 U9822 ( .A1(P2_REG1_REG_16__SCAN_IN), .A2(n8395), .B1(n9843), .B2(
        n8670), .ZN(n9830) );
  INV_X1 U9823 ( .A(n9848), .ZN(n8400) );
  OR2_X1 U9824 ( .A1(n8396), .A2(n9847), .ZN(n8399) );
  OR2_X1 U9825 ( .A1(n8412), .A2(n8665), .ZN(n8408) );
  NAND2_X1 U9826 ( .A1(n8412), .A2(n8665), .ZN(n8397) );
  NAND2_X1 U9827 ( .A1(n8408), .A2(n8397), .ZN(n8398) );
  AND3_X1 U9828 ( .A1(n8400), .A2(n8399), .A3(n8398), .ZN(n8401) );
  OAI21_X1 U9829 ( .B1(n8410), .B2(n8401), .A(n8426), .ZN(n8402) );
  OAI211_X1 U9830 ( .C1(n8404), .C2(n9856), .A(n8403), .B(n8402), .ZN(P2_U3200) );
  INV_X1 U9831 ( .A(n8405), .ZN(n8406) );
  MUX2_X1 U9832 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n7882), .S(n8421), .Z(n8417)
         );
  INV_X1 U9833 ( .A(n8408), .ZN(n8409) );
  XNOR2_X1 U9834 ( .A(n8421), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n8414) );
  OAI21_X1 U9835 ( .B1(n8413), .B2(n8412), .A(n8411), .ZN(n8419) );
  INV_X1 U9836 ( .A(n8414), .ZN(n8416) );
  MUX2_X1 U9837 ( .A(n8417), .B(n8416), .S(n4370), .Z(n8418) );
  XNOR2_X1 U9838 ( .A(n8419), .B(n8418), .ZN(n8424) );
  NAND2_X1 U9839 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(P2_U3151), .ZN(n8420) );
  OAI21_X1 U9840 ( .B1(n9844), .B2(n8421), .A(n8420), .ZN(n8422) );
  AOI21_X1 U9841 ( .B1(P2_ADDR_REG_19__SCAN_IN), .B2(n9845), .A(n8422), .ZN(
        n8423) );
  OAI21_X1 U9842 ( .B1(n8424), .B2(n9858), .A(n8423), .ZN(n8425) );
  NAND2_X1 U9843 ( .A1(n8429), .A2(n8428), .ZN(n8634) );
  AOI21_X1 U9844 ( .B1(n8430), .B2(n8634), .A(n8582), .ZN(n8434) );
  AOI21_X1 U9845 ( .B1(n8582), .B2(P2_REG2_REG_31__SCAN_IN), .A(n8434), .ZN(
        n8431) );
  OAI21_X1 U9846 ( .B1(n8432), .B2(n8550), .A(n8431), .ZN(P2_U3202) );
  AOI21_X1 U9847 ( .B1(n8582), .B2(P2_REG2_REG_30__SCAN_IN), .A(n8434), .ZN(
        n8435) );
  OAI21_X1 U9848 ( .B1(n8684), .B2(n8550), .A(n8435), .ZN(P2_U3203) );
  NAND2_X1 U9849 ( .A1(n8438), .A2(n8593), .ZN(n8440) );
  NAND2_X1 U9850 ( .A1(n8465), .A2(n8591), .ZN(n8439) );
  MUX2_X1 U9851 ( .A(n8443), .B(n8685), .S(n8633), .Z(n8449) );
  AOI22_X1 U9852 ( .A1(n8687), .A2(n8600), .B1(n8599), .B2(n8444), .ZN(n8448)
         );
  XNOR2_X1 U9853 ( .A(n8446), .B(n8445), .ZN(n8688) );
  NAND2_X1 U9854 ( .A1(n8688), .A2(n8630), .ZN(n8447) );
  NAND3_X1 U9855 ( .A1(n8449), .A2(n8448), .A3(n8447), .ZN(P2_U3205) );
  XNOR2_X1 U9856 ( .A(n8450), .B(n8451), .ZN(n8693) );
  XNOR2_X1 U9857 ( .A(n8452), .B(n8451), .ZN(n8453) );
  OAI222_X1 U9858 ( .A1(n8620), .A2(n8455), .B1(n8622), .B2(n8454), .C1(n8618), 
        .C2(n8453), .ZN(n8691) );
  MUX2_X1 U9859 ( .A(P2_REG2_REG_27__SCAN_IN), .B(n8691), .S(n8633), .Z(n8456)
         );
  INV_X1 U9860 ( .A(n8456), .ZN(n8460) );
  AOI22_X1 U9861 ( .A1(n8458), .A2(n8600), .B1(n8599), .B2(n8457), .ZN(n8459)
         );
  OAI211_X1 U9862 ( .C1(n8693), .C2(n8603), .A(n8460), .B(n8459), .ZN(P2_U3206) );
  XOR2_X1 U9863 ( .A(n8462), .B(n8461), .Z(n8701) );
  XNOR2_X1 U9864 ( .A(n8463), .B(n8462), .ZN(n8466) );
  AOI222_X1 U9865 ( .A1(n8596), .A2(n8466), .B1(n8465), .B2(n8593), .C1(n8464), 
        .C2(n8591), .ZN(n8696) );
  MUX2_X1 U9866 ( .A(n8467), .B(n8696), .S(n8633), .Z(n8470) );
  AOI22_X1 U9867 ( .A1(n8698), .A2(n8600), .B1(n8599), .B2(n8468), .ZN(n8469)
         );
  OAI211_X1 U9868 ( .C1(n8701), .C2(n8603), .A(n8470), .B(n8469), .ZN(P2_U3207) );
  INV_X1 U9869 ( .A(n8704), .ZN(n8471) );
  NOR2_X1 U9870 ( .A1(n8471), .A2(n8626), .ZN(n8477) );
  OAI21_X1 U9871 ( .B1(n8473), .B2(n8479), .A(n8472), .ZN(n8475) );
  AOI222_X1 U9872 ( .A1(n8596), .A2(n8475), .B1(n8474), .B2(n8593), .C1(n8499), 
        .C2(n8591), .ZN(n8702) );
  INV_X1 U9873 ( .A(n8702), .ZN(n8476) );
  AOI211_X1 U9874 ( .C1(n8599), .C2(n8478), .A(n8477), .B(n8476), .ZN(n8482)
         );
  XNOR2_X1 U9875 ( .A(n8480), .B(n8479), .ZN(n8705) );
  AOI22_X1 U9876 ( .A1(n8705), .A2(n8630), .B1(P2_REG2_REG_25__SCAN_IN), .B2(
        n8582), .ZN(n8481) );
  OAI21_X1 U9877 ( .B1(n8482), .B2(n8582), .A(n8481), .ZN(P2_U3208) );
  NOR2_X1 U9878 ( .A1(n8709), .A2(n8626), .ZN(n8487) );
  XOR2_X1 U9879 ( .A(n8492), .B(n8483), .Z(n8484) );
  OAI222_X1 U9880 ( .A1(n8622), .A2(n8486), .B1(n8620), .B2(n8485), .C1(n8618), 
        .C2(n8484), .ZN(n8708) );
  AOI211_X1 U9881 ( .C1(n8599), .C2(n8488), .A(n8487), .B(n8708), .ZN(n8495)
         );
  NAND2_X1 U9882 ( .A1(n8490), .A2(n8489), .ZN(n8491) );
  XOR2_X1 U9883 ( .A(n8492), .B(n8491), .Z(n8710) );
  INV_X1 U9884 ( .A(n8710), .ZN(n8493) );
  AOI22_X1 U9885 ( .A1(n8493), .A2(n8630), .B1(P2_REG2_REG_24__SCAN_IN), .B2(
        n8582), .ZN(n8494) );
  OAI21_X1 U9886 ( .B1(n8495), .B2(n8582), .A(n8494), .ZN(P2_U3209) );
  XOR2_X1 U9887 ( .A(n8496), .B(n8498), .Z(n8716) );
  INV_X1 U9888 ( .A(n8716), .ZN(n8505) );
  INV_X1 U9889 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n8501) );
  XOR2_X1 U9890 ( .A(n8497), .B(n8498), .Z(n8500) );
  AOI222_X1 U9891 ( .A1(n8596), .A2(n8500), .B1(n8499), .B2(n8593), .C1(n8525), 
        .C2(n8591), .ZN(n8713) );
  MUX2_X1 U9892 ( .A(n8501), .B(n8713), .S(n8633), .Z(n8504) );
  AOI22_X1 U9893 ( .A1(n8715), .A2(n8600), .B1(n8599), .B2(n8502), .ZN(n8503)
         );
  OAI211_X1 U9894 ( .C1(n8505), .C2(n8603), .A(n8504), .B(n8503), .ZN(P2_U3210) );
  XOR2_X1 U9895 ( .A(n8506), .B(n8507), .Z(n8724) );
  INV_X1 U9896 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n8513) );
  OR3_X1 U9897 ( .A1(n8519), .A2(n8508), .A3(n8507), .ZN(n8509) );
  NAND2_X1 U9898 ( .A1(n8510), .A2(n8509), .ZN(n8512) );
  AOI222_X1 U9899 ( .A1(n8596), .A2(n8512), .B1(n8511), .B2(n8593), .C1(n8538), 
        .C2(n8591), .ZN(n8719) );
  MUX2_X1 U9900 ( .A(n8513), .B(n8719), .S(n8633), .Z(n8516) );
  AOI22_X1 U9901 ( .A1(n8721), .A2(n8600), .B1(n8599), .B2(n8514), .ZN(n8515)
         );
  OAI211_X1 U9902 ( .C1(n8724), .C2(n8603), .A(n8516), .B(n8515), .ZN(P2_U3211) );
  XNOR2_X1 U9903 ( .A(n8518), .B(n8517), .ZN(n8730) );
  INV_X1 U9904 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n8527) );
  INV_X1 U9905 ( .A(n8519), .ZN(n8523) );
  NAND3_X1 U9906 ( .A1(n8534), .A2(n8521), .A3(n8520), .ZN(n8522) );
  NAND2_X1 U9907 ( .A1(n8523), .A2(n8522), .ZN(n8526) );
  AOI222_X1 U9908 ( .A1(n8596), .A2(n8526), .B1(n8525), .B2(n8593), .C1(n8524), 
        .C2(n8591), .ZN(n8725) );
  MUX2_X1 U9909 ( .A(n8527), .B(n8725), .S(n8633), .Z(n8530) );
  AOI22_X1 U9910 ( .A1(n8727), .A2(n8600), .B1(n8599), .B2(n8528), .ZN(n8529)
         );
  OAI211_X1 U9911 ( .C1(n8730), .C2(n8603), .A(n8530), .B(n8529), .ZN(P2_U3212) );
  NAND2_X1 U9912 ( .A1(n8532), .A2(n8531), .ZN(n8533) );
  XNOR2_X1 U9913 ( .A(n8533), .B(n8535), .ZN(n8734) );
  INV_X1 U9914 ( .A(n8734), .ZN(n8544) );
  OAI21_X1 U9915 ( .B1(n8536), .B2(n8535), .A(n8534), .ZN(n8539) );
  AOI222_X1 U9916 ( .A1(n8596), .A2(n8539), .B1(n8538), .B2(n8593), .C1(n8537), 
        .C2(n8591), .ZN(n8731) );
  MUX2_X1 U9917 ( .A(n8540), .B(n8731), .S(n8633), .Z(n8543) );
  AOI22_X1 U9918 ( .A1(n8733), .A2(n8600), .B1(n8599), .B2(n8541), .ZN(n8542)
         );
  OAI211_X1 U9919 ( .C1(n8544), .C2(n8603), .A(n8543), .B(n8542), .ZN(P2_U3213) );
  XOR2_X1 U9920 ( .A(n8545), .B(n8549), .Z(n8546) );
  OAI222_X1 U9921 ( .A1(n8622), .A2(n8547), .B1(n8620), .B2(n8578), .C1(n8546), 
        .C2(n8618), .ZN(n8663) );
  INV_X1 U9922 ( .A(n8663), .ZN(n8556) );
  XOR2_X1 U9923 ( .A(n8549), .B(n8548), .Z(n8664) );
  NOR2_X1 U9924 ( .A1(n8741), .A2(n8550), .ZN(n8554) );
  OAI22_X1 U9925 ( .A1(n8633), .A2(n8552), .B1(n8551), .B2(n8624), .ZN(n8553)
         );
  AOI211_X1 U9926 ( .C1(n8664), .C2(n8630), .A(n8554), .B(n8553), .ZN(n8555)
         );
  OAI21_X1 U9927 ( .B1(n8556), .B2(n8582), .A(n8555), .ZN(P2_U3215) );
  XNOR2_X1 U9928 ( .A(n8558), .B(n8557), .ZN(n8745) );
  INV_X1 U9929 ( .A(n8745), .ZN(n8569) );
  NAND2_X1 U9930 ( .A1(n8590), .A2(n8589), .ZN(n8588) );
  NAND2_X1 U9931 ( .A1(n8588), .A2(n8559), .ZN(n8576) );
  NAND2_X1 U9932 ( .A1(n8576), .A2(n8560), .ZN(n8562) );
  XNOR2_X1 U9933 ( .A(n8562), .B(n8561), .ZN(n8564) );
  AOI222_X1 U9934 ( .A1(n8596), .A2(n8564), .B1(n8563), .B2(n8593), .C1(n8594), 
        .C2(n8591), .ZN(n8742) );
  MUX2_X1 U9935 ( .A(n8565), .B(n8742), .S(n8633), .Z(n8568) );
  AOI22_X1 U9936 ( .A1(n8744), .A2(n8600), .B1(n8599), .B2(n8566), .ZN(n8567)
         );
  OAI211_X1 U9937 ( .C1(n8569), .C2(n8603), .A(n8568), .B(n8567), .ZN(P2_U3216) );
  NAND2_X1 U9938 ( .A1(n8571), .A2(n8570), .ZN(n8572) );
  XNOR2_X1 U9939 ( .A(n8572), .B(n8574), .ZN(n8754) );
  NAND2_X1 U9940 ( .A1(n8588), .A2(n8573), .ZN(n8575) );
  NAND2_X1 U9941 ( .A1(n8575), .A2(n8574), .ZN(n8577) );
  NAND3_X1 U9942 ( .A1(n8577), .A2(n8596), .A3(n8576), .ZN(n8581) );
  OAI22_X1 U9943 ( .A1(n8608), .A2(n8620), .B1(n8578), .B2(n8622), .ZN(n8579)
         );
  INV_X1 U9944 ( .A(n8579), .ZN(n8580) );
  MUX2_X1 U9945 ( .A(n8749), .B(n8583), .S(n8582), .Z(n8586) );
  AOI22_X1 U9946 ( .A1(n8750), .A2(n8600), .B1(n8599), .B2(n8584), .ZN(n8585)
         );
  OAI211_X1 U9947 ( .C1(n8754), .C2(n8603), .A(n8586), .B(n8585), .ZN(P2_U3217) );
  XNOR2_X1 U9948 ( .A(n8587), .B(n8589), .ZN(n8760) );
  INV_X1 U9949 ( .A(n8760), .ZN(n8604) );
  OAI21_X1 U9950 ( .B1(n8590), .B2(n8589), .A(n8588), .ZN(n8595) );
  AOI222_X1 U9951 ( .A1(n8596), .A2(n8595), .B1(n8594), .B2(n8593), .C1(n8592), 
        .C2(n8591), .ZN(n8755) );
  MUX2_X1 U9952 ( .A(n8597), .B(n8755), .S(n8633), .Z(n8602) );
  AOI22_X1 U9953 ( .A1(n8757), .A2(n8600), .B1(n8599), .B2(n8598), .ZN(n8601)
         );
  OAI211_X1 U9954 ( .C1(n8604), .C2(n8603), .A(n8602), .B(n8601), .ZN(P2_U3218) );
  XNOR2_X1 U9955 ( .A(n8605), .B(n8612), .ZN(n8606) );
  OAI222_X1 U9956 ( .A1(n8622), .A2(n8608), .B1(n8620), .B2(n8607), .C1(n8618), 
        .C2(n8606), .ZN(n9531) );
  INV_X1 U9957 ( .A(n8609), .ZN(n9530) );
  OAI22_X1 U9958 ( .A1(n9530), .A2(n8626), .B1(n8610), .B2(n8624), .ZN(n8611)
         );
  OAI21_X1 U9959 ( .B1(n9531), .B2(n8611), .A(n8633), .ZN(n8615) );
  XNOR2_X1 U9960 ( .A(n8613), .B(n8612), .ZN(n9533) );
  NAND2_X1 U9961 ( .A1(n9533), .A2(n8630), .ZN(n8614) );
  OAI211_X1 U9962 ( .C1(n6348), .C2(n8633), .A(n8615), .B(n8614), .ZN(P2_U3219) );
  XOR2_X1 U9963 ( .A(n8629), .B(n8616), .Z(n8617) );
  OAI222_X1 U9964 ( .A1(n8622), .A2(n8621), .B1(n8620), .B2(n8619), .C1(n8618), 
        .C2(n8617), .ZN(n9535) );
  INV_X1 U9965 ( .A(n8623), .ZN(n9534) );
  OAI22_X1 U9966 ( .A1(n9534), .A2(n8626), .B1(n8625), .B2(n8624), .ZN(n8627)
         );
  OAI21_X1 U9967 ( .B1(n9535), .B2(n8627), .A(n8633), .ZN(n8632) );
  XOR2_X1 U9968 ( .A(n8629), .B(n8628), .Z(n9537) );
  NAND2_X1 U9969 ( .A1(n9537), .A2(n8630), .ZN(n8631) );
  OAI211_X1 U9970 ( .C1(n7569), .C2(n8633), .A(n8632), .B(n8631), .ZN(P2_U3220) );
  NAND2_X1 U9971 ( .A1(n8679), .A2(n8675), .ZN(n8635) );
  INV_X1 U9972 ( .A(n8634), .ZN(n8680) );
  NAND2_X1 U9973 ( .A1(n8680), .A2(n9929), .ZN(n8636) );
  OAI211_X1 U9974 ( .C1(n9929), .C2(n7347), .A(n8635), .B(n8636), .ZN(P2_U3490) );
  NAND2_X1 U9975 ( .A1(n9927), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n8637) );
  OAI211_X1 U9976 ( .C1(n8684), .C2(n8667), .A(n8637), .B(n8636), .ZN(P2_U3489) );
  INV_X1 U9977 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n8638) );
  MUX2_X1 U9978 ( .A(n8638), .B(n8685), .S(n9929), .Z(n8640) );
  AOI22_X1 U9979 ( .A1(n8688), .A2(n8676), .B1(n8675), .B2(n8687), .ZN(n8639)
         );
  NAND2_X1 U9980 ( .A1(n8640), .A2(n8639), .ZN(P2_U3487) );
  MUX2_X1 U9981 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n8691), .S(n9929), .Z(n8642)
         );
  OAI22_X1 U9982 ( .A1(n8693), .A2(n8673), .B1(n8692), .B2(n8667), .ZN(n8641)
         );
  OR2_X1 U9983 ( .A1(n8642), .A2(n8641), .ZN(P2_U3486) );
  INV_X1 U9984 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n8643) );
  MUX2_X1 U9985 ( .A(n8643), .B(n8696), .S(n9929), .Z(n8645) );
  NAND2_X1 U9986 ( .A1(n8698), .A2(n8675), .ZN(n8644) );
  OAI211_X1 U9987 ( .C1(n8701), .C2(n8673), .A(n8645), .B(n8644), .ZN(P2_U3485) );
  INV_X1 U9988 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n8646) );
  MUX2_X1 U9989 ( .A(n8646), .B(n8702), .S(n9929), .Z(n8648) );
  AOI22_X1 U9990 ( .A1(n8705), .A2(n8676), .B1(n8675), .B2(n8704), .ZN(n8647)
         );
  NAND2_X1 U9991 ( .A1(n8648), .A2(n8647), .ZN(P2_U3484) );
  MUX2_X1 U9992 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n8708), .S(n9929), .Z(n8650)
         );
  OAI22_X1 U9993 ( .A1(n8710), .A2(n8673), .B1(n8709), .B2(n8667), .ZN(n8649)
         );
  OR2_X1 U9994 ( .A1(n8650), .A2(n8649), .ZN(P2_U3483) );
  MUX2_X1 U9995 ( .A(n8651), .B(n8713), .S(n9929), .Z(n8653) );
  AOI22_X1 U9996 ( .A1(n8716), .A2(n8676), .B1(n8675), .B2(n8715), .ZN(n8652)
         );
  NAND2_X1 U9997 ( .A1(n8653), .A2(n8652), .ZN(P2_U3482) );
  INV_X1 U9998 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n8654) );
  MUX2_X1 U9999 ( .A(n8654), .B(n8719), .S(n9929), .Z(n8656) );
  NAND2_X1 U10000 ( .A1(n8721), .A2(n8675), .ZN(n8655) );
  OAI211_X1 U10001 ( .C1(n8724), .C2(n8673), .A(n8656), .B(n8655), .ZN(
        P2_U3481) );
  INV_X1 U10002 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n8657) );
  MUX2_X1 U10003 ( .A(n8657), .B(n8725), .S(n9929), .Z(n8659) );
  NAND2_X1 U10004 ( .A1(n8727), .A2(n8675), .ZN(n8658) );
  OAI211_X1 U10005 ( .C1(n8673), .C2(n8730), .A(n8659), .B(n8658), .ZN(
        P2_U3480) );
  MUX2_X1 U10006 ( .A(n8660), .B(n8731), .S(n9929), .Z(n8662) );
  AOI22_X1 U10007 ( .A1(n8734), .A2(n8676), .B1(n8675), .B2(n8733), .ZN(n8661)
         );
  NAND2_X1 U10008 ( .A1(n8662), .A2(n8661), .ZN(P2_U3479) );
  AOI21_X1 U10009 ( .B1(n9906), .B2(n8664), .A(n8663), .ZN(n8737) );
  MUX2_X1 U10010 ( .A(n8665), .B(n8737), .S(n9929), .Z(n8666) );
  OAI21_X1 U10011 ( .B1(n8741), .B2(n8667), .A(n8666), .ZN(P2_U3477) );
  MUX2_X1 U10012 ( .A(n9850), .B(n8742), .S(n9929), .Z(n8669) );
  AOI22_X1 U10013 ( .A1(n8745), .A2(n8676), .B1(n8675), .B2(n8744), .ZN(n8668)
         );
  NAND2_X1 U10014 ( .A1(n8669), .A2(n8668), .ZN(P2_U3476) );
  MUX2_X1 U10015 ( .A(n8749), .B(n8670), .S(n9927), .Z(n8672) );
  NAND2_X1 U10016 ( .A1(n8750), .A2(n8675), .ZN(n8671) );
  OAI211_X1 U10017 ( .C1(n8754), .C2(n8673), .A(n8672), .B(n8671), .ZN(
        P2_U3475) );
  MUX2_X1 U10018 ( .A(n8674), .B(n8755), .S(n9929), .Z(n8678) );
  AOI22_X1 U10019 ( .A1(n8760), .A2(n8676), .B1(n8675), .B2(n8757), .ZN(n8677)
         );
  NAND2_X1 U10020 ( .A1(n8678), .A2(n8677), .ZN(P2_U3474) );
  NAND2_X1 U10021 ( .A1(n8679), .A2(n8758), .ZN(n8681) );
  NAND2_X1 U10022 ( .A1(n8680), .A2(n9914), .ZN(n8682) );
  OAI211_X1 U10023 ( .C1(n7349), .C2(n9914), .A(n8681), .B(n8682), .ZN(
        P2_U3458) );
  NAND2_X1 U10024 ( .A1(n9915), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n8683) );
  OAI211_X1 U10025 ( .C1(n8684), .C2(n8740), .A(n8683), .B(n8682), .ZN(
        P2_U3457) );
  INV_X1 U10026 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n8686) );
  MUX2_X1 U10027 ( .A(n8686), .B(n8685), .S(n9914), .Z(n8690) );
  AOI22_X1 U10028 ( .A1(n8688), .A2(n8759), .B1(n8758), .B2(n8687), .ZN(n8689)
         );
  NAND2_X1 U10029 ( .A1(n8690), .A2(n8689), .ZN(P2_U3455) );
  MUX2_X1 U10030 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n8691), .S(n9914), .Z(n8695) );
  OAI22_X1 U10031 ( .A1(n8693), .A2(n8753), .B1(n8692), .B2(n8740), .ZN(n8694)
         );
  OR2_X1 U10032 ( .A1(n8695), .A2(n8694), .ZN(P2_U3454) );
  INV_X1 U10033 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n8697) );
  MUX2_X1 U10034 ( .A(n8697), .B(n8696), .S(n9914), .Z(n8700) );
  NAND2_X1 U10035 ( .A1(n8698), .A2(n8758), .ZN(n8699) );
  OAI211_X1 U10036 ( .C1(n8701), .C2(n8753), .A(n8700), .B(n8699), .ZN(
        P2_U3453) );
  INV_X1 U10037 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n8703) );
  MUX2_X1 U10038 ( .A(n8703), .B(n8702), .S(n9914), .Z(n8707) );
  AOI22_X1 U10039 ( .A1(n8705), .A2(n8759), .B1(n8758), .B2(n8704), .ZN(n8706)
         );
  NAND2_X1 U10040 ( .A1(n8707), .A2(n8706), .ZN(P2_U3452) );
  MUX2_X1 U10041 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n8708), .S(n9914), .Z(n8712) );
  OAI22_X1 U10042 ( .A1(n8710), .A2(n8753), .B1(n8709), .B2(n8740), .ZN(n8711)
         );
  OR2_X1 U10043 ( .A1(n8712), .A2(n8711), .ZN(P2_U3451) );
  INV_X1 U10044 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n8714) );
  MUX2_X1 U10045 ( .A(n8714), .B(n8713), .S(n9914), .Z(n8718) );
  AOI22_X1 U10046 ( .A1(n8716), .A2(n8759), .B1(n8758), .B2(n8715), .ZN(n8717)
         );
  NAND2_X1 U10047 ( .A1(n8718), .A2(n8717), .ZN(P2_U3450) );
  INV_X1 U10048 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n8720) );
  MUX2_X1 U10049 ( .A(n8720), .B(n8719), .S(n9914), .Z(n8723) );
  NAND2_X1 U10050 ( .A1(n8721), .A2(n8758), .ZN(n8722) );
  OAI211_X1 U10051 ( .C1(n8724), .C2(n8753), .A(n8723), .B(n8722), .ZN(
        P2_U3449) );
  INV_X1 U10052 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n8726) );
  MUX2_X1 U10053 ( .A(n8726), .B(n8725), .S(n9914), .Z(n8729) );
  NAND2_X1 U10054 ( .A1(n8727), .A2(n8758), .ZN(n8728) );
  OAI211_X1 U10055 ( .C1(n8730), .C2(n8753), .A(n8729), .B(n8728), .ZN(
        P2_U3448) );
  MUX2_X1 U10056 ( .A(n8732), .B(n8731), .S(n9914), .Z(n8736) );
  AOI22_X1 U10057 ( .A1(n8734), .A2(n8759), .B1(n8758), .B2(n8733), .ZN(n8735)
         );
  NAND2_X1 U10058 ( .A1(n8736), .A2(n8735), .ZN(P2_U3447) );
  INV_X1 U10059 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n8738) );
  MUX2_X1 U10060 ( .A(n8738), .B(n8737), .S(n9914), .Z(n8739) );
  OAI21_X1 U10061 ( .B1(n8741), .B2(n8740), .A(n8739), .ZN(P2_U3444) );
  INV_X1 U10062 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n8743) );
  MUX2_X1 U10063 ( .A(n8743), .B(n8742), .S(n9914), .Z(n8747) );
  AOI22_X1 U10064 ( .A1(n8745), .A2(n8759), .B1(n8758), .B2(n8744), .ZN(n8746)
         );
  NAND2_X1 U10065 ( .A1(n8747), .A2(n8746), .ZN(P2_U3441) );
  INV_X1 U10066 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n8748) );
  MUX2_X1 U10067 ( .A(n8749), .B(n8748), .S(n9915), .Z(n8752) );
  NAND2_X1 U10068 ( .A1(n8750), .A2(n8758), .ZN(n8751) );
  OAI211_X1 U10069 ( .C1(n8754), .C2(n8753), .A(n8752), .B(n8751), .ZN(
        P2_U3438) );
  INV_X1 U10070 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n8756) );
  MUX2_X1 U10071 ( .A(n8756), .B(n8755), .S(n9914), .Z(n8762) );
  AOI22_X1 U10072 ( .A1(n8760), .A2(n8759), .B1(n8758), .B2(n8757), .ZN(n8761)
         );
  NAND2_X1 U10073 ( .A1(n8762), .A2(n8761), .ZN(P2_U3435) );
  INV_X1 U10074 ( .A(n8763), .ZN(n9477) );
  NOR4_X1 U10075 ( .A1(n8765), .A2(P2_IR_REG_30__SCAN_IN), .A3(P2_U3151), .A4(
        n8764), .ZN(n8766) );
  AOI21_X1 U10076 ( .B1(n8774), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n8766), .ZN(
        n8767) );
  OAI21_X1 U10077 ( .B1(n9477), .B2(n8777), .A(n8767), .ZN(P2_U3264) );
  INV_X1 U10078 ( .A(n8768), .ZN(n9480) );
  AOI22_X1 U10079 ( .A1(n8769), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n8774), .ZN(n8770) );
  OAI21_X1 U10080 ( .B1(n9480), .B2(n8777), .A(n8770), .ZN(P2_U3265) );
  AOI22_X1 U10081 ( .A1(n8771), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_29__SCAN_IN), .B2(n8774), .ZN(n8772) );
  OAI21_X1 U10082 ( .B1(n8773), .B2(n8777), .A(n8772), .ZN(P2_U3266) );
  NAND2_X1 U10083 ( .A1(n8774), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n8775) );
  OAI211_X1 U10084 ( .C1(n8778), .C2(n8777), .A(n8776), .B(n8775), .ZN(
        P2_U3267) );
  MUX2_X1 U10085 ( .A(n8779), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  AOI22_X1 U10086 ( .A1(n8926), .A2(n9345), .B1(P1_REG3_REG_27__SCAN_IN), .B2(
        P1_U3086), .ZN(n8786) );
  INV_X1 U10087 ( .A(n9325), .ZN(n9149) );
  AOI22_X1 U10088 ( .A1(n9148), .A2(n8927), .B1(n8945), .B2(n9149), .ZN(n8785)
         );
  NAND2_X1 U10089 ( .A1(n9156), .A2(n8928), .ZN(n8784) );
  NAND4_X1 U10090 ( .A1(n8787), .A2(n8786), .A3(n8785), .A4(n8784), .ZN(
        P1_U3214) );
  XNOR2_X1 U10091 ( .A(n8789), .B(n8788), .ZN(n8790) );
  XNOR2_X1 U10092 ( .A(n8791), .B(n8790), .ZN(n8796) );
  AOI22_X1 U10093 ( .A1(n8927), .A2(n8792), .B1(n8945), .B2(n8952), .ZN(n8793)
         );
  NAND2_X1 U10094 ( .A1(P1_U3086), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n9673) );
  OAI211_X1 U10095 ( .C1(n9775), .C2(n8940), .A(n8793), .B(n9673), .ZN(n8794)
         );
  AOI21_X1 U10096 ( .B1(n9427), .B2(n8928), .A(n8794), .ZN(n8795) );
  OAI21_X1 U10097 ( .B1(n8796), .B2(n8920), .A(n8795), .ZN(P1_U3215) );
  INV_X1 U10098 ( .A(n8879), .ZN(n8799) );
  NOR3_X1 U10099 ( .A1(n8903), .A2(n8907), .A3(n8797), .ZN(n8798) );
  OAI21_X1 U10100 ( .B1(n8799), .B2(n8798), .A(n8936), .ZN(n8804) );
  OAI22_X1 U10101 ( .A1(n8899), .A2(n9360), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8800), .ZN(n8802) );
  OAI22_X1 U10102 ( .A1(n9213), .A2(n8941), .B1(n8940), .B2(n9361), .ZN(n8801)
         );
  AOI211_X1 U10103 ( .C1(n9363), .C2(n8928), .A(n8802), .B(n8801), .ZN(n8803)
         );
  NAND2_X1 U10104 ( .A1(n8804), .A2(n8803), .ZN(P1_U3216) );
  NAND2_X1 U10105 ( .A1(n8806), .A2(n8805), .ZN(n8813) );
  INV_X1 U10106 ( .A(n8807), .ZN(n8809) );
  NAND2_X1 U10107 ( .A1(n8809), .A2(n8808), .ZN(n8810) );
  OAI21_X1 U10108 ( .B1(n8809), .B2(n8808), .A(n8810), .ZN(n8915) );
  NOR2_X1 U10109 ( .A1(n8915), .A2(n8916), .ZN(n8914) );
  INV_X1 U10110 ( .A(n8810), .ZN(n8811) );
  NOR2_X1 U10111 ( .A1(n8914), .A2(n8811), .ZN(n8812) );
  XOR2_X1 U10112 ( .A(n8813), .B(n8812), .Z(n8817) );
  AOI22_X1 U10113 ( .A1(n9271), .A2(n8927), .B1(n8926), .B2(n9405), .ZN(n8814)
         );
  NAND2_X1 U10114 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9082) );
  OAI211_X1 U10115 ( .C1(n9278), .C2(n8899), .A(n8814), .B(n9082), .ZN(n8815)
         );
  AOI21_X1 U10116 ( .B1(n9392), .B2(n8928), .A(n8815), .ZN(n8816) );
  OAI21_X1 U10117 ( .B1(n8817), .B2(n8920), .A(n8816), .ZN(P1_U3219) );
  OAI21_X1 U10118 ( .B1(n8820), .B2(n8819), .A(n8818), .ZN(n8821) );
  NAND2_X1 U10119 ( .A1(n8821), .A2(n8936), .ZN(n8827) );
  AOI22_X1 U10120 ( .A1(n8926), .A2(n8822), .B1(n8945), .B2(n8962), .ZN(n8826)
         );
  AOI22_X1 U10121 ( .A1(P1_REG3_REG_1__SCAN_IN), .A2(n8824), .B1(n8928), .B2(
        n8823), .ZN(n8825) );
  NAND3_X1 U10122 ( .A1(n8827), .A2(n8826), .A3(n8825), .ZN(P1_U3222) );
  XOR2_X1 U10123 ( .A(n8829), .B(n8828), .Z(n8835) );
  OAI22_X1 U10124 ( .A1(n8899), .A2(n9361), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8830), .ZN(n8833) );
  INV_X1 U10125 ( .A(n8831), .ZN(n9243) );
  OAI22_X1 U10126 ( .A1(n8941), .A2(n9243), .B1(n8940), .B2(n9278), .ZN(n8832)
         );
  AOI211_X1 U10127 ( .C1(n9241), .C2(n8928), .A(n8833), .B(n8832), .ZN(n8834)
         );
  OAI21_X1 U10128 ( .B1(n8835), .B2(n8920), .A(n8834), .ZN(P1_U3223) );
  XOR2_X1 U10129 ( .A(n8837), .B(n8836), .Z(n8842) );
  AOI22_X1 U10130 ( .A1(n8838), .A2(n8927), .B1(n8926), .B2(n9756), .ZN(n8839)
         );
  NAND2_X1 U10131 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n9642) );
  OAI211_X1 U10132 ( .C1(n9775), .C2(n8899), .A(n8839), .B(n9642), .ZN(n8840)
         );
  AOI21_X1 U10133 ( .B1(n9780), .B2(n8928), .A(n8840), .ZN(n8841) );
  OAI21_X1 U10134 ( .B1(n8842), .B2(n8920), .A(n8841), .ZN(P1_U3224) );
  AOI21_X1 U10135 ( .B1(n8844), .B2(n8843), .A(n8924), .ZN(n8850) );
  OAI22_X1 U10136 ( .A1(n8899), .A2(n9324), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8845), .ZN(n8848) );
  INV_X1 U10137 ( .A(n8846), .ZN(n9180) );
  OAI22_X1 U10138 ( .A1(n9180), .A2(n8941), .B1(n8940), .B2(n9360), .ZN(n8847)
         );
  AOI211_X1 U10139 ( .C1(n9185), .C2(n8928), .A(n8848), .B(n8847), .ZN(n8849)
         );
  OAI21_X1 U10140 ( .B1(n8850), .B2(n8920), .A(n8849), .ZN(P1_U3225) );
  INV_X1 U10141 ( .A(n8852), .ZN(n8853) );
  XNOR2_X1 U10142 ( .A(n8851), .B(n8852), .ZN(n8934) );
  NAND2_X1 U10143 ( .A1(n8934), .A2(n8935), .ZN(n8933) );
  OAI21_X1 U10144 ( .B1(n8853), .B2(n8851), .A(n8933), .ZN(n8857) );
  XNOR2_X1 U10145 ( .A(n8855), .B(n8854), .ZN(n8856) );
  XNOR2_X1 U10146 ( .A(n8857), .B(n8856), .ZN(n8863) );
  AOI22_X1 U10147 ( .A1(n8858), .A2(n8927), .B1(n8926), .B2(n8952), .ZN(n8859)
         );
  NAND2_X1 U10148 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9698) );
  OAI211_X1 U10149 ( .C1(n9414), .C2(n8899), .A(n8859), .B(n9698), .ZN(n8860)
         );
  AOI21_X1 U10150 ( .B1(n8861), .B2(n8928), .A(n8860), .ZN(n8862) );
  OAI21_X1 U10151 ( .B1(n8863), .B2(n8920), .A(n8862), .ZN(P1_U3226) );
  XNOR2_X1 U10152 ( .A(n8865), .B(n8864), .ZN(n8866) );
  XNOR2_X1 U10153 ( .A(n8867), .B(n8866), .ZN(n8876) );
  AOI21_X1 U10154 ( .B1(n8869), .B2(n8868), .A(P1_U3086), .ZN(n8873) );
  AOI22_X1 U10155 ( .A1(n8926), .A2(n9406), .B1(n8945), .B2(n9405), .ZN(n8872)
         );
  NAND3_X1 U10156 ( .A1(n8927), .A2(n8870), .A3(n9057), .ZN(n8871) );
  OAI211_X1 U10157 ( .C1(n8873), .C2(n9057), .A(n8872), .B(n8871), .ZN(n8874)
         );
  AOI21_X1 U10158 ( .B1(n9096), .B2(n8928), .A(n8874), .ZN(n8875) );
  OAI21_X1 U10159 ( .B1(n8876), .B2(n8920), .A(n8875), .ZN(P1_U3228) );
  AND3_X1 U10160 ( .A1(n8879), .A2(n8878), .A3(n8877), .ZN(n8880) );
  OAI21_X1 U10161 ( .B1(n8881), .B2(n8880), .A(n8936), .ZN(n8885) );
  AOI22_X1 U10162 ( .A1(n8945), .A2(n9196), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3086), .ZN(n8884) );
  AOI22_X1 U10163 ( .A1(n9202), .A2(n8927), .B1(n8926), .B2(n9369), .ZN(n8883)
         );
  NAND2_X1 U10164 ( .A1(n9201), .A2(n8928), .ZN(n8882) );
  NAND4_X1 U10165 ( .A1(n8885), .A2(n8884), .A3(n8883), .A4(n8882), .ZN(
        P1_U3229) );
  XNOR2_X1 U10166 ( .A(n8887), .B(n8886), .ZN(n8888) );
  XNOR2_X1 U10167 ( .A(n8889), .B(n8888), .ZN(n8894) );
  OAI22_X1 U10168 ( .A1(n8899), .A2(n9255), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8890), .ZN(n8892) );
  OAI22_X1 U10169 ( .A1(n8941), .A2(n9259), .B1(n8940), .B2(n9256), .ZN(n8891)
         );
  AOI211_X1 U10170 ( .C1(n9388), .C2(n8928), .A(n8892), .B(n8891), .ZN(n8893)
         );
  OAI21_X1 U10171 ( .B1(n8894), .B2(n8920), .A(n8893), .ZN(P1_U3233) );
  XOR2_X1 U10172 ( .A(n8896), .B(n8895), .Z(n8902) );
  AOI22_X1 U10173 ( .A1(n8897), .A2(n8927), .B1(n8926), .B2(n8955), .ZN(n8898)
         );
  NAND2_X1 U10174 ( .A1(P1_U3086), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n9657) );
  OAI211_X1 U10175 ( .C1(n8939), .C2(n8899), .A(n8898), .B(n9657), .ZN(n8900)
         );
  AOI21_X1 U10176 ( .B1(n9788), .B2(n8928), .A(n8900), .ZN(n8901) );
  OAI21_X1 U10177 ( .B1(n8902), .B2(n8920), .A(n8901), .ZN(P1_U3234) );
  INV_X1 U10178 ( .A(n8903), .ZN(n8908) );
  OAI21_X1 U10179 ( .B1(n8905), .B2(n8907), .A(n8904), .ZN(n8906) );
  OAI21_X1 U10180 ( .B1(n8908), .B2(n8907), .A(n8906), .ZN(n8909) );
  NAND2_X1 U10181 ( .A1(n8909), .A2(n8936), .ZN(n8913) );
  AOI22_X1 U10182 ( .A1(n8945), .A2(n9369), .B1(P1_REG3_REG_22__SCAN_IN), .B2(
        P1_U3086), .ZN(n8912) );
  AOI22_X1 U10183 ( .A1(n8927), .A2(n9227), .B1(n8926), .B2(n9368), .ZN(n8911)
         );
  NAND2_X1 U10184 ( .A1(n9233), .A2(n8928), .ZN(n8910) );
  NAND4_X1 U10185 ( .A1(n8913), .A2(n8912), .A3(n8911), .A4(n8910), .ZN(
        P1_U3235) );
  AOI21_X1 U10186 ( .B1(n8916), .B2(n8915), .A(n8914), .ZN(n8921) );
  AOI22_X1 U10187 ( .A1(n8927), .A2(n9292), .B1(n8945), .B2(n9396), .ZN(n8917)
         );
  NAND2_X1 U10188 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9713) );
  OAI211_X1 U10189 ( .C1(n9414), .C2(n8940), .A(n8917), .B(n9713), .ZN(n8918)
         );
  AOI21_X1 U10190 ( .B1(n9300), .B2(n8928), .A(n8918), .ZN(n8919) );
  OAI21_X1 U10191 ( .B1(n8921), .B2(n8920), .A(n8919), .ZN(P1_U3238) );
  OAI21_X1 U10192 ( .B1(n8924), .B2(n8923), .A(n8922), .ZN(n8925) );
  NAND3_X1 U10193 ( .A1(n4841), .A2(n8936), .A3(n8925), .ZN(n8932) );
  AOI22_X1 U10194 ( .A1(n8926), .A2(n9196), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3086), .ZN(n8931) );
  AOI22_X1 U10195 ( .A1(n8927), .A2(n9165), .B1(n8945), .B2(n9166), .ZN(n8930)
         );
  NAND2_X1 U10196 ( .A1(n9164), .A2(n8928), .ZN(n8929) );
  NAND4_X1 U10197 ( .A1(n8932), .A2(n8931), .A3(n8930), .A4(n8929), .ZN(
        P1_U3240) );
  OAI21_X1 U10198 ( .B1(n8935), .B2(n8934), .A(n8933), .ZN(n8937) );
  NAND2_X1 U10199 ( .A1(n8937), .A2(n8936), .ZN(n8947) );
  NAND2_X1 U10200 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9685) );
  INV_X1 U10201 ( .A(n9685), .ZN(n8944) );
  INV_X1 U10202 ( .A(n8938), .ZN(n8942) );
  OAI22_X1 U10203 ( .A1(n8942), .A2(n8941), .B1(n8940), .B2(n8939), .ZN(n8943)
         );
  AOI211_X1 U10204 ( .C1(n8945), .C2(n9406), .A(n8944), .B(n8943), .ZN(n8946)
         );
  OAI211_X1 U10205 ( .C1(n8949), .C2(n8948), .A(n8947), .B(n8946), .ZN(
        P1_U3241) );
  MUX2_X1 U10206 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n8950), .S(P1_U3973), .Z(
        P1_U3584) );
  INV_X1 U10207 ( .A(n8951), .ZN(n9140) );
  MUX2_X1 U10208 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n9140), .S(P1_U3973), .Z(
        P1_U3583) );
  MUX2_X1 U10209 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9149), .S(P1_U3973), .Z(
        P1_U3582) );
  MUX2_X1 U10210 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9166), .S(P1_U3973), .Z(
        P1_U3581) );
  MUX2_X1 U10211 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9345), .S(P1_U3973), .Z(
        P1_U3580) );
  MUX2_X1 U10212 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9196), .S(P1_U3973), .Z(
        P1_U3579) );
  MUX2_X1 U10213 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9344), .S(P1_U3973), .Z(
        P1_U3578) );
  MUX2_X1 U10214 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9369), .S(P1_U3973), .Z(
        P1_U3577) );
  MUX2_X1 U10215 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9378), .S(P1_U3973), .Z(
        P1_U3576) );
  MUX2_X1 U10216 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9368), .S(P1_U3973), .Z(
        P1_U3575) );
  MUX2_X1 U10217 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9377), .S(P1_U3973), .Z(
        P1_U3574) );
  MUX2_X1 U10218 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9396), .S(P1_U3973), .Z(
        P1_U3573) );
  MUX2_X1 U10219 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9405), .S(P1_U3973), .Z(
        P1_U3572) );
  MUX2_X1 U10220 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9397), .S(P1_U3973), .Z(
        P1_U3571) );
  MUX2_X1 U10221 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9406), .S(P1_U3973), .Z(
        P1_U3570) );
  MUX2_X1 U10222 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n8952), .S(P1_U3973), .Z(
        P1_U3569) );
  MUX2_X1 U10223 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n8953), .S(P1_U3973), .Z(
        P1_U3568) );
  MUX2_X1 U10224 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n8954), .S(P1_U3973), .Z(
        P1_U3567) );
  MUX2_X1 U10225 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n8955), .S(P1_U3973), .Z(
        P1_U3566) );
  MUX2_X1 U10226 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n9756), .S(P1_U3973), .Z(
        P1_U3565) );
  MUX2_X1 U10227 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n8956), .S(P1_U3973), .Z(
        P1_U3564) );
  MUX2_X1 U10228 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n9755), .S(P1_U3973), .Z(
        P1_U3563) );
  MUX2_X1 U10229 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9746), .S(P1_U3973), .Z(
        P1_U3562) );
  MUX2_X1 U10230 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n8957), .S(P1_U3973), .Z(
        P1_U3561) );
  MUX2_X1 U10231 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n8958), .S(P1_U3973), .Z(
        P1_U3560) );
  MUX2_X1 U10232 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n8959), .S(P1_U3973), .Z(
        P1_U3559) );
  MUX2_X1 U10233 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n8960), .S(P1_U3973), .Z(
        P1_U3558) );
  MUX2_X1 U10234 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n8961), .S(P1_U3973), .Z(
        P1_U3557) );
  MUX2_X1 U10235 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n8962), .S(P1_U3973), .Z(
        P1_U3556) );
  MUX2_X1 U10236 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n9719), .S(P1_U3973), .Z(
        P1_U3555) );
  XNOR2_X1 U10237 ( .A(n8970), .B(P1_REG2_REG_1__SCAN_IN), .ZN(n8967) );
  AND2_X1 U10238 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n9562) );
  INV_X1 U10239 ( .A(n8963), .ZN(n8964) );
  NAND2_X1 U10240 ( .A1(n8965), .A2(n8964), .ZN(n9547) );
  INV_X1 U10241 ( .A(n9485), .ZN(n9561) );
  NAND2_X1 U10242 ( .A1(n9564), .A2(n9561), .ZN(n8966) );
  OR2_X1 U10243 ( .A1(n9547), .A2(n8966), .ZN(n9687) );
  NAND2_X1 U10244 ( .A1(n8967), .A2(n9562), .ZN(n8989) );
  OAI211_X1 U10245 ( .C1(n8967), .C2(n9562), .A(n9700), .B(n8989), .ZN(n8974)
         );
  XNOR2_X1 U10246 ( .A(n8970), .B(P1_REG1_REG_1__SCAN_IN), .ZN(n8969) );
  AND2_X1 U10247 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n8968) );
  NAND2_X1 U10248 ( .A1(n8969), .A2(n8968), .ZN(n8980) );
  OAI211_X1 U10249 ( .C1(n8969), .C2(n8968), .A(n9664), .B(n8980), .ZN(n8973)
         );
  AOI22_X1 U10250 ( .A1(n9581), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n8972) );
  INV_X1 U10251 ( .A(n9692), .ZN(n9707) );
  INV_X1 U10252 ( .A(n8970), .ZN(n8987) );
  NAND2_X1 U10253 ( .A1(n9707), .A2(n8987), .ZN(n8971) );
  NAND4_X1 U10254 ( .A1(n8974), .A2(n8973), .A3(n8972), .A4(n8971), .ZN(
        P1_U3244) );
  INV_X1 U10255 ( .A(n9581), .ZN(n9716) );
  INV_X1 U10256 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n8976) );
  OAI21_X1 U10257 ( .B1(n9716), .B2(n8976), .A(n8975), .ZN(n8977) );
  AOI21_X1 U10258 ( .B1(n9009), .B2(n9707), .A(n8977), .ZN(n8996) );
  XNOR2_X1 U10259 ( .A(n9009), .B(n6950), .ZN(n8984) );
  NAND2_X1 U10260 ( .A1(n9560), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n8978) );
  OAI21_X1 U10261 ( .B1(n9560), .B2(P1_REG1_REG_2__SCAN_IN), .A(n8978), .ZN(
        n9551) );
  INV_X1 U10262 ( .A(n9551), .ZN(n8981) );
  NAND2_X1 U10263 ( .A1(n8987), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n8979) );
  NAND2_X1 U10264 ( .A1(n8980), .A2(n8979), .ZN(n9549) );
  AND2_X1 U10265 ( .A1(n8981), .A2(n9549), .ZN(n9550) );
  AND2_X1 U10266 ( .A1(n9560), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n8982) );
  OAI211_X1 U10267 ( .C1(n8984), .C2(n8983), .A(n9664), .B(n9011), .ZN(n8995)
         );
  XNOR2_X1 U10268 ( .A(n9009), .B(n8985), .ZN(n8993) );
  INV_X1 U10269 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n8986) );
  XNOR2_X1 U10270 ( .A(n9560), .B(n8986), .ZN(n9554) );
  NAND2_X1 U10271 ( .A1(n8987), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n8988) );
  NAND2_X1 U10272 ( .A1(n8989), .A2(n8988), .ZN(n9553) );
  AND2_X1 U10273 ( .A1(n9554), .A2(n9553), .ZN(n9555) );
  INV_X1 U10274 ( .A(n9555), .ZN(n8991) );
  NAND2_X1 U10275 ( .A1(n9560), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n8990) );
  NAND2_X1 U10276 ( .A1(n8991), .A2(n8990), .ZN(n8992) );
  NAND2_X1 U10277 ( .A1(n8992), .A2(n8993), .ZN(n8999) );
  OAI211_X1 U10278 ( .C1(n8993), .C2(n8992), .A(n9700), .B(n8999), .ZN(n8994)
         );
  NAND3_X1 U10279 ( .A1(n8996), .A2(n8995), .A3(n8994), .ZN(P1_U3246) );
  NOR2_X1 U10280 ( .A1(n9045), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n8997) );
  AOI21_X1 U10281 ( .B1(P1_REG2_REG_9__SCAN_IN), .B2(n9045), .A(n8997), .ZN(
        n9005) );
  NAND2_X1 U10282 ( .A1(n9009), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n8998) );
  NAND2_X1 U10283 ( .A1(n8999), .A2(n8998), .ZN(n9575) );
  MUX2_X1 U10284 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n6710), .S(n9013), .Z(n9576)
         );
  AND2_X1 U10285 ( .A1(n9575), .A2(n9576), .ZN(n9573) );
  NAND2_X1 U10286 ( .A1(n9017), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n9000) );
  OAI21_X1 U10287 ( .B1(n9017), .B2(P1_REG2_REG_5__SCAN_IN), .A(n9000), .ZN(
        n9588) );
  NOR2_X1 U10288 ( .A1(n9587), .A2(n9588), .ZN(n9586) );
  AOI21_X1 U10289 ( .B1(P1_REG2_REG_5__SCAN_IN), .B2(n9017), .A(n9586), .ZN(
        n9606) );
  INV_X1 U10290 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n9001) );
  AOI22_X1 U10291 ( .A1(n9019), .A2(n9001), .B1(P1_REG2_REG_6__SCAN_IN), .B2(
        n9611), .ZN(n9607) );
  NOR2_X1 U10292 ( .A1(n9606), .A2(n9607), .ZN(n9605) );
  NAND2_X1 U10293 ( .A1(n9022), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n9002) );
  OAI21_X1 U10294 ( .B1(n9022), .B2(P1_REG2_REG_7__SCAN_IN), .A(n9002), .ZN(
        n9507) );
  NOR2_X1 U10295 ( .A1(n9506), .A2(n9507), .ZN(n9505) );
  NAND2_X1 U10296 ( .A1(n9025), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n9003) );
  OAI21_X1 U10297 ( .B1(n9025), .B2(P1_REG2_REG_8__SCAN_IN), .A(n9003), .ZN(
        n9517) );
  NOR2_X1 U10298 ( .A1(n9516), .A2(n9517), .ZN(n9515) );
  AOI21_X1 U10299 ( .B1(P1_REG2_REG_8__SCAN_IN), .B2(n9025), .A(n9515), .ZN(
        n9004) );
  NAND2_X1 U10300 ( .A1(n9005), .A2(n9004), .ZN(n9044) );
  OAI21_X1 U10301 ( .B1(n9005), .B2(n9004), .A(n9044), .ZN(n9006) );
  NAND2_X1 U10302 ( .A1(n9006), .A2(n9700), .ZN(n9032) );
  AOI21_X1 U10303 ( .B1(n9581), .B2(P1_ADDR_REG_9__SCAN_IN), .A(n9007), .ZN(
        n9031) );
  NOR2_X1 U10304 ( .A1(n9045), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n9008) );
  AOI21_X1 U10305 ( .B1(P1_REG1_REG_9__SCAN_IN), .B2(n9045), .A(n9008), .ZN(
        n9027) );
  NAND2_X1 U10306 ( .A1(n9009), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n9010) );
  NAND2_X1 U10307 ( .A1(n9011), .A2(n9010), .ZN(n9571) );
  MUX2_X1 U10308 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n9012), .S(n9013), .Z(n9572)
         );
  NAND2_X1 U10309 ( .A1(n9571), .A2(n9572), .ZN(n9570) );
  NAND2_X1 U10310 ( .A1(n9013), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n9014) );
  OR2_X1 U10311 ( .A1(n9017), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n9016) );
  NAND2_X1 U10312 ( .A1(n9017), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n9015) );
  NAND2_X1 U10313 ( .A1(n9016), .A2(n9015), .ZN(n9591) );
  NOR2_X1 U10314 ( .A1(n9592), .A2(n9591), .ZN(n9590) );
  INV_X1 U10315 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n9018) );
  MUX2_X1 U10316 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n9018), .S(n9611), .Z(n9603)
         );
  NOR2_X1 U10317 ( .A1(n9602), .A2(n9603), .ZN(n9601) );
  AOI21_X1 U10318 ( .B1(n9019), .B2(P1_REG1_REG_6__SCAN_IN), .A(n9601), .ZN(
        n9503) );
  OR2_X1 U10319 ( .A1(n9022), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n9021) );
  NAND2_X1 U10320 ( .A1(n9022), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n9020) );
  NAND2_X1 U10321 ( .A1(n9021), .A2(n9020), .ZN(n9502) );
  NOR2_X1 U10322 ( .A1(n9503), .A2(n9502), .ZN(n9501) );
  OR2_X1 U10323 ( .A1(n9025), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n9024) );
  NAND2_X1 U10324 ( .A1(n9025), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n9023) );
  NAND2_X1 U10325 ( .A1(n9024), .A2(n9023), .ZN(n9521) );
  NOR2_X1 U10326 ( .A1(n9520), .A2(n9521), .ZN(n9519) );
  AOI21_X1 U10327 ( .B1(P1_REG1_REG_8__SCAN_IN), .B2(n9025), .A(n9519), .ZN(
        n9026) );
  NAND2_X1 U10328 ( .A1(n9027), .A2(n9026), .ZN(n9035) );
  OAI21_X1 U10329 ( .B1(n9027), .B2(n9026), .A(n9035), .ZN(n9028) );
  NAND2_X1 U10330 ( .A1(n9028), .A2(n9664), .ZN(n9030) );
  NAND2_X1 U10331 ( .A1(n9707), .A2(n9045), .ZN(n9029) );
  NAND4_X1 U10332 ( .A1(n9032), .A2(n9031), .A3(n9030), .A4(n9029), .ZN(
        P1_U3252) );
  XNOR2_X1 U10333 ( .A(n9071), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n9072) );
  INV_X1 U10334 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n9033) );
  MUX2_X1 U10335 ( .A(n9033), .B(P1_REG1_REG_13__SCAN_IN), .S(n9644), .Z(n9651) );
  OR2_X1 U10336 ( .A1(n9629), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n9038) );
  INV_X1 U10337 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n9034) );
  MUX2_X1 U10338 ( .A(n9034), .B(P1_REG1_REG_10__SCAN_IN), .S(n9498), .Z(n9491) );
  OAI21_X1 U10339 ( .B1(n9045), .B2(P1_REG1_REG_9__SCAN_IN), .A(n9035), .ZN(
        n9492) );
  NOR2_X1 U10340 ( .A1(n9491), .A2(n9492), .ZN(n9490) );
  INV_X1 U10341 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n9036) );
  MUX2_X1 U10342 ( .A(n9036), .B(P1_REG1_REG_11__SCAN_IN), .S(n9047), .Z(n9617) );
  NOR2_X1 U10343 ( .A1(n9616), .A2(n9617), .ZN(n9615) );
  AOI21_X1 U10344 ( .B1(n9047), .B2(P1_REG1_REG_11__SCAN_IN), .A(n9615), .ZN(
        n9635) );
  INV_X1 U10345 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n9037) );
  MUX2_X1 U10346 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n9037), .S(n9629), .Z(n9636) );
  NOR2_X1 U10347 ( .A1(n9651), .A2(n9650), .ZN(n9649) );
  XNOR2_X1 U10348 ( .A(n9659), .B(P1_REG1_REG_14__SCAN_IN), .ZN(n9661) );
  NOR2_X1 U10349 ( .A1(n9662), .A2(n9661), .ZN(n9660) );
  NOR2_X1 U10350 ( .A1(n9039), .A2(n9049), .ZN(n9040) );
  XNOR2_X1 U10351 ( .A(n9049), .B(n9039), .ZN(n9678) );
  NOR2_X1 U10352 ( .A1(n9677), .A2(n9678), .ZN(n9676) );
  NOR2_X1 U10353 ( .A1(n9040), .A2(n9676), .ZN(n9690) );
  INV_X1 U10354 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9421) );
  XNOR2_X1 U10355 ( .A(n9052), .B(n9421), .ZN(n9691) );
  AOI22_X1 U10356 ( .A1(n9690), .A2(n9691), .B1(n9421), .B2(n9693), .ZN(n9073)
         );
  XOR2_X1 U10357 ( .A(n9072), .B(n9073), .Z(n9062) );
  INV_X1 U10358 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n9063) );
  XNOR2_X1 U10359 ( .A(n9071), .B(n9063), .ZN(n9055) );
  NAND2_X1 U10360 ( .A1(n9644), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n9041) );
  OAI21_X1 U10361 ( .B1(n9644), .B2(P1_REG2_REG_13__SCAN_IN), .A(n9041), .ZN(
        n9647) );
  NOR2_X1 U10362 ( .A1(n9629), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n9042) );
  AOI21_X1 U10363 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(n9629), .A(n9042), .ZN(
        n9632) );
  NAND2_X1 U10364 ( .A1(n9498), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n9043) );
  OAI21_X1 U10365 ( .B1(n9498), .B2(P1_REG2_REG_10__SCAN_IN), .A(n9043), .ZN(
        n9494) );
  OAI21_X1 U10366 ( .B1(n9045), .B2(P1_REG2_REG_9__SCAN_IN), .A(n9044), .ZN(
        n9495) );
  NOR2_X1 U10367 ( .A1(n9494), .A2(n9495), .ZN(n9493) );
  NAND2_X1 U10368 ( .A1(n9047), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n9046) );
  OAI21_X1 U10369 ( .B1(n9047), .B2(P1_REG2_REG_11__SCAN_IN), .A(n9046), .ZN(
        n9621) );
  NOR2_X1 U10370 ( .A1(n9620), .A2(n9621), .ZN(n9619) );
  AOI21_X1 U10371 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n9047), .A(n9619), .ZN(
        n9631) );
  NAND2_X1 U10372 ( .A1(n9632), .A2(n9631), .ZN(n9630) );
  OAI21_X1 U10373 ( .B1(n9629), .B2(P1_REG2_REG_12__SCAN_IN), .A(n9630), .ZN(
        n9646) );
  NOR2_X1 U10374 ( .A1(n9647), .A2(n9646), .ZN(n9645) );
  NAND2_X1 U10375 ( .A1(n9659), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n9048) );
  OAI21_X1 U10376 ( .B1(n9659), .B2(P1_REG2_REG_14__SCAN_IN), .A(n9048), .ZN(
        n9667) );
  NOR2_X1 U10377 ( .A1(n9666), .A2(n9667), .ZN(n9665) );
  NOR2_X1 U10378 ( .A1(n9050), .A2(n9049), .ZN(n9051) );
  INV_X1 U10379 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n9680) );
  XOR2_X1 U10380 ( .A(n9684), .B(n9050), .Z(n9681) );
  NOR2_X1 U10381 ( .A1(n9680), .A2(n9681), .ZN(n9679) );
  XNOR2_X1 U10382 ( .A(n9052), .B(P1_REG2_REG_16__SCAN_IN), .ZN(n9688) );
  NAND2_X1 U10383 ( .A1(n9052), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n9053) );
  NAND2_X1 U10384 ( .A1(n9054), .A2(n9055), .ZN(n9066) );
  OAI21_X1 U10385 ( .B1(n9055), .B2(n9054), .A(n9066), .ZN(n9056) );
  NAND2_X1 U10386 ( .A1(n9056), .A2(n9700), .ZN(n9061) );
  INV_X1 U10387 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n9058) );
  OAI22_X1 U10388 ( .A1(n9716), .A2(n9058), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9057), .ZN(n9059) );
  AOI21_X1 U10389 ( .B1(n9071), .B2(n9707), .A(n9059), .ZN(n9060) );
  OAI211_X1 U10390 ( .C1(n9704), .C2(n9062), .A(n9061), .B(n9060), .ZN(
        P1_U3260) );
  NAND2_X1 U10391 ( .A1(n9064), .A2(n9063), .ZN(n9065) );
  NAND2_X1 U10392 ( .A1(n9708), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9068) );
  OAI21_X1 U10393 ( .B1(n9708), .B2(P1_REG2_REG_18__SCAN_IN), .A(n9068), .ZN(
        n9067) );
  INV_X1 U10394 ( .A(n9067), .ZN(n9702) );
  NAND2_X1 U10395 ( .A1(n9703), .A2(n9702), .ZN(n9701) );
  NAND2_X1 U10396 ( .A1(n9701), .A2(n9068), .ZN(n9070) );
  INV_X1 U10397 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n9069) );
  XNOR2_X1 U10398 ( .A(n9070), .B(n9069), .ZN(n9076) );
  OAI22_X1 U10399 ( .A1(n9073), .A2(n9072), .B1(P1_REG1_REG_17__SCAN_IN), .B2(
        n9071), .ZN(n9706) );
  NAND2_X1 U10400 ( .A1(n9708), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n9074) );
  OAI21_X1 U10401 ( .B1(n9708), .B2(P1_REG1_REG_18__SCAN_IN), .A(n9074), .ZN(
        n9705) );
  OR2_X1 U10402 ( .A1(n9706), .A2(n9705), .ZN(n9709) );
  NAND2_X1 U10403 ( .A1(n9709), .A2(n9074), .ZN(n9075) );
  XOR2_X1 U10404 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9075), .Z(n9077) );
  AOI22_X1 U10405 ( .A1(n9076), .A2(n9700), .B1(n9664), .B2(n9077), .ZN(n9081)
         );
  INV_X1 U10406 ( .A(n9076), .ZN(n9079) );
  OAI21_X1 U10407 ( .B1(n9077), .B2(n9704), .A(n9692), .ZN(n9078) );
  OAI211_X1 U10408 ( .C1(n4636), .C2(n9716), .A(n9083), .B(n9082), .ZN(
        P1_U3262) );
  INV_X1 U10409 ( .A(n9392), .ZN(n9274) );
  OR2_X2 U10410 ( .A1(n9226), .A2(n9363), .ZN(n9218) );
  OR2_X2 U10411 ( .A1(n9153), .A2(n9318), .ZN(n9133) );
  NOR2_X2 U10412 ( .A1(n9316), .A2(n9133), .ZN(n9123) );
  NAND2_X1 U10413 ( .A1(n9123), .A2(n9439), .ZN(n9092) );
  INV_X1 U10414 ( .A(P1_B_REG_SCAN_IN), .ZN(n9085) );
  OR2_X1 U10415 ( .A1(n9485), .A2(n9085), .ZN(n9086) );
  NAND2_X1 U10416 ( .A1(n9757), .A2(n9086), .ZN(n9122) );
  INV_X1 U10417 ( .A(n9122), .ZN(n9087) );
  NAND2_X1 U10418 ( .A1(n9088), .A2(n9087), .ZN(n9309) );
  NOR2_X1 U10419 ( .A1(n9293), .A2(n9309), .ZN(n9094) );
  NOR2_X1 U10420 ( .A1(n9435), .A2(n9273), .ZN(n9089) );
  AOI211_X1 U10421 ( .C1(n9293), .C2(P1_REG2_REG_31__SCAN_IN), .A(n9094), .B(
        n9089), .ZN(n9090) );
  OAI21_X1 U10422 ( .B1(n9307), .B2(n9302), .A(n9090), .ZN(P1_U3263) );
  OR2_X1 U10423 ( .A1(n9439), .A2(n9123), .ZN(n9091) );
  NAND3_X1 U10424 ( .A1(n9092), .A2(n9319), .A3(n9091), .ZN(n9310) );
  NOR2_X1 U10425 ( .A1(n9439), .A2(n9273), .ZN(n9093) );
  AOI211_X1 U10426 ( .C1(n9293), .C2(P1_REG2_REG_30__SCAN_IN), .A(n9094), .B(
        n9093), .ZN(n9095) );
  OAI21_X1 U10427 ( .B1(n9302), .B2(n9310), .A(n9095), .ZN(P1_U3264) );
  INV_X1 U10428 ( .A(n9201), .ZN(n9454) );
  INV_X1 U10429 ( .A(n9241), .ZN(n9380) );
  INV_X1 U10430 ( .A(n9388), .ZN(n9263) );
  NAND2_X1 U10431 ( .A1(n9096), .A2(n9397), .ZN(n9097) );
  INV_X1 U10432 ( .A(n9286), .ZN(n9100) );
  NAND2_X1 U10433 ( .A1(n9372), .A2(n9361), .ZN(n9102) );
  INV_X1 U10434 ( .A(n9363), .ZN(n9103) );
  NAND2_X1 U10435 ( .A1(n9185), .A2(n9196), .ZN(n9104) );
  NAND2_X1 U10436 ( .A1(n9162), .A2(n9161), .ZN(n9106) );
  NAND2_X1 U10437 ( .A1(n9164), .A2(n9345), .ZN(n9105) );
  INV_X1 U10438 ( .A(n9145), .ZN(n9108) );
  NAND2_X1 U10439 ( .A1(n9445), .A2(n9335), .ZN(n9107) );
  XNOR2_X1 U10440 ( .A(n9110), .B(n9109), .ZN(n9313) );
  INV_X1 U10441 ( .A(n9313), .ZN(n9130) );
  NAND2_X1 U10442 ( .A1(n9238), .A2(n9113), .ZN(n9225) );
  NAND2_X1 U10443 ( .A1(n9225), .A2(n9224), .ZN(n9115) );
  NAND2_X1 U10444 ( .A1(n9115), .A2(n9114), .ZN(n9207) );
  AND3_X2 U10445 ( .A1(n9193), .A2(n9175), .A3(n9176), .ZN(n9178) );
  NAND2_X1 U10446 ( .A1(n9139), .A2(n5608), .ZN(n9138) );
  INV_X1 U10447 ( .A(n9316), .ZN(n9127) );
  AOI211_X1 U10448 ( .C1(n9316), .C2(n9133), .A(n9792), .B(n9123), .ZN(n9315)
         );
  NAND2_X1 U10449 ( .A1(n9315), .A2(n9284), .ZN(n9126) );
  AOI22_X1 U10450 ( .A1(n9293), .A2(P1_REG2_REG_29__SCAN_IN), .B1(n9124), .B2(
        n9291), .ZN(n9125) );
  OAI211_X1 U10451 ( .C1(n9127), .C2(n9273), .A(n9126), .B(n9125), .ZN(n9128)
         );
  AOI21_X1 U10452 ( .B1(n9314), .B2(n9265), .A(n9128), .ZN(n9129) );
  OAI21_X1 U10453 ( .B1(n9130), .B2(n9306), .A(n9129), .ZN(P1_U3356) );
  INV_X1 U10454 ( .A(n9133), .ZN(n9134) );
  AOI21_X1 U10455 ( .B1(n9318), .B2(n9153), .A(n9134), .ZN(n9320) );
  INV_X1 U10456 ( .A(n9318), .ZN(n9137) );
  AOI22_X1 U10457 ( .A1(n9293), .A2(P1_REG2_REG_28__SCAN_IN), .B1(n9135), .B2(
        n9291), .ZN(n9136) );
  OAI21_X1 U10458 ( .B1(n9137), .B2(n9273), .A(n9136), .ZN(n9142) );
  NOR2_X1 U10459 ( .A1(n9322), .A2(n9293), .ZN(n9141) );
  OAI21_X1 U10460 ( .B1(n9323), .B2(n9306), .A(n9144), .ZN(P1_U3265) );
  XNOR2_X1 U10461 ( .A(n9146), .B(n9108), .ZN(n9329) );
  XNOR2_X1 U10462 ( .A(n9147), .B(n9108), .ZN(n9331) );
  NAND2_X1 U10463 ( .A1(n9331), .A2(n9212), .ZN(n9158) );
  AOI22_X1 U10464 ( .A1(n9293), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n9148), .B2(
        n9291), .ZN(n9151) );
  NAND2_X1 U10465 ( .A1(n9294), .A2(n9149), .ZN(n9150) );
  OAI211_X1 U10466 ( .C1(n9324), .C2(n9297), .A(n9151), .B(n9150), .ZN(n9155)
         );
  NAND2_X1 U10467 ( .A1(n9156), .A2(n9163), .ZN(n9152) );
  NAND3_X1 U10468 ( .A1(n9153), .A2(n9319), .A3(n9152), .ZN(n9327) );
  NOR2_X1 U10469 ( .A1(n9327), .A2(n9302), .ZN(n9154) );
  AOI211_X1 U10470 ( .C1(n9299), .C2(n9156), .A(n9155), .B(n9154), .ZN(n9157)
         );
  OAI211_X1 U10471 ( .C1(n9329), .C2(n9173), .A(n9158), .B(n9157), .ZN(
        P1_U3266) );
  AOI21_X1 U10472 ( .B1(n9160), .B2(n9161), .A(n9159), .ZN(n9339) );
  XOR2_X1 U10473 ( .A(n9162), .B(n9161), .Z(n9341) );
  NAND2_X1 U10474 ( .A1(n9341), .A2(n9212), .ZN(n9172) );
  AOI211_X1 U10475 ( .C1(n9164), .C2(n9179), .A(n9792), .B(n4607), .ZN(n9337)
         );
  INV_X1 U10476 ( .A(n9164), .ZN(n9449) );
  NOR2_X1 U10477 ( .A1(n9449), .A2(n9273), .ZN(n9170) );
  AOI22_X1 U10478 ( .A1(n9293), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n9165), .B2(
        n9291), .ZN(n9168) );
  NAND2_X1 U10479 ( .A1(n9294), .A2(n9166), .ZN(n9167) );
  OAI211_X1 U10480 ( .C1(n9334), .C2(n9297), .A(n9168), .B(n9167), .ZN(n9169)
         );
  AOI211_X1 U10481 ( .C1(n9337), .C2(n9284), .A(n9170), .B(n9169), .ZN(n9171)
         );
  OAI211_X1 U10482 ( .C1(n9339), .C2(n9173), .A(n9172), .B(n9171), .ZN(
        P1_U3267) );
  XOR2_X1 U10483 ( .A(n9174), .B(n9175), .Z(n9352) );
  AOI21_X1 U10484 ( .B1(n9193), .B2(n9176), .A(n9175), .ZN(n9177) );
  OR2_X1 U10485 ( .A1(n9178), .A2(n9177), .ZN(n9350) );
  OAI211_X1 U10486 ( .C1(n9348), .C2(n9200), .A(n9319), .B(n9179), .ZN(n9347)
         );
  INV_X1 U10487 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n9181) );
  OAI22_X1 U10488 ( .A1(n9265), .A2(n9181), .B1(n9180), .B2(n9242), .ZN(n9182)
         );
  AOI21_X1 U10489 ( .B1(n9294), .B2(n9345), .A(n9182), .ZN(n9183) );
  OAI21_X1 U10490 ( .B1(n9360), .B2(n9297), .A(n9183), .ZN(n9184) );
  AOI21_X1 U10491 ( .B1(n9185), .B2(n9299), .A(n9184), .ZN(n9186) );
  OAI21_X1 U10492 ( .B1(n9347), .B2(n9302), .A(n9186), .ZN(n9187) );
  AOI21_X1 U10493 ( .B1(n9350), .B2(n9304), .A(n9187), .ZN(n9188) );
  OAI21_X1 U10494 ( .B1(n9352), .B2(n9306), .A(n9188), .ZN(P1_U3268) );
  OAI21_X1 U10495 ( .B1(n9191), .B2(n9190), .A(n9189), .ZN(n9353) );
  AND2_X1 U10496 ( .A1(n9209), .A2(n9192), .ZN(n9195) );
  OAI211_X1 U10497 ( .C1(n9195), .C2(n9194), .A(n9193), .B(n9765), .ZN(n9198)
         );
  NAND2_X1 U10498 ( .A1(n9196), .A2(n9757), .ZN(n9197) );
  OAI211_X1 U10499 ( .C1(n9199), .C2(n9776), .A(n9198), .B(n9197), .ZN(n9354)
         );
  AOI211_X1 U10500 ( .C1(n9201), .C2(n9218), .A(n9792), .B(n9200), .ZN(n9355)
         );
  NAND2_X1 U10501 ( .A1(n9355), .A2(n9284), .ZN(n9204) );
  AOI22_X1 U10502 ( .A1(n9293), .A2(P1_REG2_REG_24__SCAN_IN), .B1(n9202), .B2(
        n9291), .ZN(n9203) );
  OAI211_X1 U10503 ( .C1(n9454), .C2(n9273), .A(n9204), .B(n9203), .ZN(n9205)
         );
  AOI21_X1 U10504 ( .B1(n9354), .B2(n9265), .A(n9205), .ZN(n9206) );
  OAI21_X1 U10505 ( .B1(n9353), .B2(n9306), .A(n9206), .ZN(P1_U3269) );
  OR2_X1 U10506 ( .A1(n9207), .A2(n9211), .ZN(n9208) );
  NAND2_X1 U10507 ( .A1(n9209), .A2(n9208), .ZN(n9210) );
  NAND2_X1 U10508 ( .A1(n9210), .A2(n9765), .ZN(n9365) );
  XOR2_X1 U10509 ( .A(n9211), .B(n4426), .Z(n9359) );
  NAND2_X1 U10510 ( .A1(n9359), .A2(n9212), .ZN(n9222) );
  OAI22_X1 U10511 ( .A1(n9265), .A2(n9214), .B1(n9213), .B2(n9242), .ZN(n9215)
         );
  AOI21_X1 U10512 ( .B1(n9294), .B2(n9344), .A(n9215), .ZN(n9216) );
  OAI21_X1 U10513 ( .B1(n9361), .B2(n9297), .A(n9216), .ZN(n9220) );
  NAND2_X1 U10514 ( .A1(n9226), .A2(n9363), .ZN(n9217) );
  NAND3_X1 U10515 ( .A1(n9218), .A2(n9319), .A3(n9217), .ZN(n9364) );
  NOR2_X1 U10516 ( .A1(n9364), .A2(n9302), .ZN(n9219) );
  AOI211_X1 U10517 ( .C1(n9299), .C2(n9363), .A(n9220), .B(n9219), .ZN(n9221)
         );
  OAI211_X1 U10518 ( .C1(n9293), .C2(n9365), .A(n9222), .B(n9221), .ZN(
        P1_U3270) );
  XOR2_X1 U10519 ( .A(n9224), .B(n9223), .Z(n9376) );
  XNOR2_X1 U10520 ( .A(n9225), .B(n9224), .ZN(n9374) );
  OAI211_X1 U10521 ( .C1(n9372), .C2(n4435), .A(n9319), .B(n9226), .ZN(n9371)
         );
  INV_X1 U10522 ( .A(n9227), .ZN(n9228) );
  OAI22_X1 U10523 ( .A1(n9265), .A2(n9229), .B1(n9228), .B2(n9242), .ZN(n9230)
         );
  AOI21_X1 U10524 ( .B1(n9294), .B2(n9369), .A(n9230), .ZN(n9231) );
  OAI21_X1 U10525 ( .B1(n9255), .B2(n9297), .A(n9231), .ZN(n9232) );
  AOI21_X1 U10526 ( .B1(n9233), .B2(n9299), .A(n9232), .ZN(n9234) );
  OAI21_X1 U10527 ( .B1(n9371), .B2(n9302), .A(n9234), .ZN(n9235) );
  AOI21_X1 U10528 ( .B1(n9374), .B2(n9304), .A(n9235), .ZN(n9236) );
  OAI21_X1 U10529 ( .B1(n9376), .B2(n9306), .A(n9236), .ZN(P1_U3271) );
  XOR2_X1 U10530 ( .A(n9239), .B(n9237), .Z(n9385) );
  OAI21_X1 U10531 ( .B1(n9240), .B2(n9239), .A(n9238), .ZN(n9383) );
  AOI211_X1 U10532 ( .C1(n9241), .C2(n9257), .A(n9792), .B(n4435), .ZN(n9381)
         );
  NAND2_X1 U10533 ( .A1(n9381), .A2(n9284), .ZN(n9248) );
  INV_X1 U10534 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n9244) );
  OAI22_X1 U10535 ( .A1(n9265), .A2(n9244), .B1(n9243), .B2(n9242), .ZN(n9246)
         );
  NOR2_X1 U10536 ( .A1(n9297), .A2(n9278), .ZN(n9245) );
  AOI211_X1 U10537 ( .C1(n9294), .C2(n9378), .A(n9246), .B(n9245), .ZN(n9247)
         );
  OAI211_X1 U10538 ( .C1(n9380), .C2(n9273), .A(n9248), .B(n9247), .ZN(n9249)
         );
  AOI21_X1 U10539 ( .B1(n9304), .B2(n9383), .A(n9249), .ZN(n9250) );
  OAI21_X1 U10540 ( .B1(n9385), .B2(n9306), .A(n9250), .ZN(P1_U3272) );
  XNOR2_X1 U10541 ( .A(n9251), .B(n9253), .ZN(n9390) );
  XOR2_X1 U10542 ( .A(n9253), .B(n9252), .Z(n9254) );
  OAI222_X1 U10543 ( .A1(n9776), .A2(n9256), .B1(n9774), .B2(n9255), .C1(n9254), .C2(n9783), .ZN(n9386) );
  INV_X1 U10544 ( .A(n9257), .ZN(n9258) );
  AOI211_X1 U10545 ( .C1(n9388), .C2(n9269), .A(n9792), .B(n9258), .ZN(n9387)
         );
  NAND2_X1 U10546 ( .A1(n9387), .A2(n9284), .ZN(n9262) );
  INV_X1 U10547 ( .A(n9259), .ZN(n9260) );
  AOI22_X1 U10548 ( .A1(n9293), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9260), .B2(
        n9291), .ZN(n9261) );
  OAI211_X1 U10549 ( .C1(n9263), .C2(n9273), .A(n9262), .B(n9261), .ZN(n9264)
         );
  AOI21_X1 U10550 ( .B1(n9386), .B2(n9265), .A(n9264), .ZN(n9266) );
  OAI21_X1 U10551 ( .B1(n9390), .B2(n9306), .A(n9266), .ZN(P1_U3273) );
  XNOR2_X1 U10552 ( .A(n9267), .B(n9275), .ZN(n9395) );
  INV_X1 U10553 ( .A(n9268), .ZN(n9289) );
  INV_X1 U10554 ( .A(n9269), .ZN(n9270) );
  AOI211_X1 U10555 ( .C1(n9392), .C2(n9289), .A(n9792), .B(n9270), .ZN(n9391)
         );
  AOI22_X1 U10556 ( .A1(n9293), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9271), .B2(
        n9291), .ZN(n9272) );
  OAI21_X1 U10557 ( .B1(n9274), .B2(n9273), .A(n9272), .ZN(n9283) );
  AOI21_X1 U10558 ( .B1(n9276), .B2(n9275), .A(n9783), .ZN(n9281) );
  OAI22_X1 U10559 ( .A1(n9278), .A2(n9774), .B1(n9277), .B2(n9776), .ZN(n9279)
         );
  AOI21_X1 U10560 ( .B1(n9281), .B2(n9280), .A(n9279), .ZN(n9394) );
  NOR2_X1 U10561 ( .A1(n9394), .A2(n9293), .ZN(n9282) );
  AOI211_X1 U10562 ( .C1(n9391), .C2(n9284), .A(n9283), .B(n9282), .ZN(n9285)
         );
  OAI21_X1 U10563 ( .B1(n9395), .B2(n9306), .A(n9285), .ZN(P1_U3274) );
  XOR2_X1 U10564 ( .A(n9286), .B(n9287), .Z(n9404) );
  XNOR2_X1 U10565 ( .A(n9288), .B(n9287), .ZN(n9402) );
  OAI211_X1 U10566 ( .C1(n9400), .C2(n9290), .A(n9289), .B(n9319), .ZN(n9399)
         );
  AOI22_X1 U10567 ( .A1(n9293), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9292), .B2(
        n9291), .ZN(n9296) );
  NAND2_X1 U10568 ( .A1(n9294), .A2(n9396), .ZN(n9295) );
  OAI211_X1 U10569 ( .C1(n9414), .C2(n9297), .A(n9296), .B(n9295), .ZN(n9298)
         );
  AOI21_X1 U10570 ( .B1(n9300), .B2(n9299), .A(n9298), .ZN(n9301) );
  OAI21_X1 U10571 ( .B1(n9399), .B2(n9302), .A(n9301), .ZN(n9303) );
  AOI21_X1 U10572 ( .B1(n9402), .B2(n9304), .A(n9303), .ZN(n9305) );
  OAI21_X1 U10573 ( .B1(n9404), .B2(n9306), .A(n9305), .ZN(P1_U3275) );
  AND2_X1 U10574 ( .A1(n9310), .A2(n9309), .ZN(n9436) );
  MUX2_X1 U10575 ( .A(n9311), .B(n9436), .S(n9813), .Z(n9312) );
  OAI21_X1 U10576 ( .B1(n9439), .B2(n9423), .A(n9312), .ZN(P1_U3552) );
  NAND2_X1 U10577 ( .A1(n9313), .A2(n9794), .ZN(n9317) );
  MUX2_X1 U10578 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n9440), .S(n9813), .Z(
        P1_U3551) );
  AOI22_X1 U10579 ( .A1(n9320), .A2(n9319), .B1(n9787), .B2(n9318), .ZN(n9321)
         );
  MUX2_X1 U10580 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9441), .S(n9813), .Z(
        P1_U3550) );
  INV_X1 U10581 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n9332) );
  OAI22_X1 U10582 ( .A1(n9325), .A2(n9774), .B1(n9324), .B2(n9776), .ZN(n9326)
         );
  INV_X1 U10583 ( .A(n9326), .ZN(n9328) );
  OAI211_X1 U10584 ( .C1(n9329), .C2(n9783), .A(n9328), .B(n9327), .ZN(n9330)
         );
  AOI21_X1 U10585 ( .B1(n9331), .B2(n9794), .A(n9330), .ZN(n9442) );
  MUX2_X1 U10586 ( .A(n9332), .B(n9442), .S(n9813), .Z(n9333) );
  OAI21_X1 U10587 ( .B1(n9445), .B2(n9423), .A(n9333), .ZN(P1_U3549) );
  INV_X1 U10588 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n9342) );
  OAI22_X1 U10589 ( .A1(n9335), .A2(n9774), .B1(n9334), .B2(n9776), .ZN(n9336)
         );
  NOR2_X1 U10590 ( .A1(n9337), .A2(n9336), .ZN(n9338) );
  OAI21_X1 U10591 ( .B1(n9339), .B2(n9783), .A(n9338), .ZN(n9340) );
  AOI21_X1 U10592 ( .B1(n9341), .B2(n9794), .A(n9340), .ZN(n9446) );
  MUX2_X1 U10593 ( .A(n9342), .B(n9446), .S(n9813), .Z(n9343) );
  OAI21_X1 U10594 ( .B1(n9449), .B2(n9423), .A(n9343), .ZN(P1_U3548) );
  AOI22_X1 U10595 ( .A1(n9757), .A2(n9345), .B1(n9344), .B2(n9754), .ZN(n9346)
         );
  OAI211_X1 U10596 ( .C1(n9348), .C2(n9768), .A(n9347), .B(n9346), .ZN(n9349)
         );
  AOI21_X1 U10597 ( .B1(n9350), .B2(n9765), .A(n9349), .ZN(n9351) );
  OAI21_X1 U10598 ( .B1(n9352), .B2(n9760), .A(n9351), .ZN(n9450) );
  MUX2_X1 U10599 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9450), .S(n9813), .Z(
        P1_U3547) );
  INV_X1 U10600 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n9357) );
  INV_X1 U10601 ( .A(n9353), .ZN(n9356) );
  AOI211_X1 U10602 ( .C1(n9356), .C2(n9794), .A(n9355), .B(n9354), .ZN(n9451)
         );
  MUX2_X1 U10603 ( .A(n9357), .B(n9451), .S(n9813), .Z(n9358) );
  OAI21_X1 U10604 ( .B1(n9454), .B2(n9423), .A(n9358), .ZN(P1_U3546) );
  NAND2_X1 U10605 ( .A1(n9359), .A2(n9794), .ZN(n9367) );
  OAI22_X1 U10606 ( .A1(n9361), .A2(n9776), .B1(n9360), .B2(n9774), .ZN(n9362)
         );
  AOI21_X1 U10607 ( .B1(n9363), .B2(n9787), .A(n9362), .ZN(n9366) );
  NAND4_X1 U10608 ( .A1(n9367), .A2(n9366), .A3(n9365), .A4(n9364), .ZN(n9455)
         );
  MUX2_X1 U10609 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9455), .S(n9813), .Z(
        P1_U3545) );
  AOI22_X1 U10610 ( .A1(n9369), .A2(n9757), .B1(n9754), .B2(n9368), .ZN(n9370)
         );
  OAI211_X1 U10611 ( .C1(n9372), .C2(n9768), .A(n9371), .B(n9370), .ZN(n9373)
         );
  AOI21_X1 U10612 ( .B1(n9374), .B2(n9765), .A(n9373), .ZN(n9375) );
  OAI21_X1 U10613 ( .B1(n9376), .B2(n9760), .A(n9375), .ZN(n9456) );
  MUX2_X1 U10614 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9456), .S(n9813), .Z(
        P1_U3544) );
  AOI22_X1 U10615 ( .A1(n9378), .A2(n9757), .B1(n9754), .B2(n9377), .ZN(n9379)
         );
  OAI21_X1 U10616 ( .B1(n9380), .B2(n9768), .A(n9379), .ZN(n9382) );
  AOI211_X1 U10617 ( .C1(n9383), .C2(n9765), .A(n9382), .B(n9381), .ZN(n9384)
         );
  OAI21_X1 U10618 ( .B1(n9385), .B2(n9760), .A(n9384), .ZN(n9457) );
  MUX2_X1 U10619 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9457), .S(n9813), .Z(
        P1_U3543) );
  AOI211_X1 U10620 ( .C1(n9787), .C2(n9388), .A(n9387), .B(n9386), .ZN(n9389)
         );
  OAI21_X1 U10621 ( .B1(n9390), .B2(n9760), .A(n9389), .ZN(n9458) );
  MUX2_X1 U10622 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9458), .S(n9813), .Z(
        P1_U3542) );
  AOI21_X1 U10623 ( .B1(n9787), .B2(n9392), .A(n9391), .ZN(n9393) );
  OAI211_X1 U10624 ( .C1(n9395), .C2(n9760), .A(n9394), .B(n9393), .ZN(n9459)
         );
  MUX2_X1 U10625 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9459), .S(n9813), .Z(
        P1_U3541) );
  AOI22_X1 U10626 ( .A1(n9754), .A2(n9397), .B1(n9396), .B2(n9757), .ZN(n9398)
         );
  OAI211_X1 U10627 ( .C1(n9400), .C2(n9768), .A(n9399), .B(n9398), .ZN(n9401)
         );
  AOI21_X1 U10628 ( .B1(n9402), .B2(n9765), .A(n9401), .ZN(n9403) );
  OAI21_X1 U10629 ( .B1(n9404), .B2(n9760), .A(n9403), .ZN(n9460) );
  MUX2_X1 U10630 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9460), .S(n9813), .Z(
        P1_U3540) );
  AOI22_X1 U10631 ( .A1(n9754), .A2(n9406), .B1(n9405), .B2(n9757), .ZN(n9407)
         );
  OAI21_X1 U10632 ( .B1(n9408), .B2(n9768), .A(n9407), .ZN(n9409) );
  AOI211_X1 U10633 ( .C1(n9411), .C2(n9765), .A(n9410), .B(n9409), .ZN(n9412)
         );
  OAI21_X1 U10634 ( .B1(n9413), .B2(n9760), .A(n9412), .ZN(n9461) );
  MUX2_X1 U10635 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9461), .S(n9813), .Z(
        P1_U3539) );
  OAI22_X1 U10636 ( .A1(n9425), .A2(n9776), .B1(n9414), .B2(n9774), .ZN(n9415)
         );
  NOR2_X1 U10637 ( .A1(n9416), .A2(n9415), .ZN(n9417) );
  OAI21_X1 U10638 ( .B1(n9418), .B2(n9783), .A(n9417), .ZN(n9419) );
  AOI21_X1 U10639 ( .B1(n9420), .B2(n9794), .A(n9419), .ZN(n9462) );
  MUX2_X1 U10640 ( .A(n9421), .B(n9462), .S(n9813), .Z(n9422) );
  OAI21_X1 U10641 ( .B1(n9466), .B2(n9423), .A(n9422), .ZN(P1_U3538) );
  NAND2_X1 U10642 ( .A1(n9424), .A2(n9794), .ZN(n9431) );
  OAI22_X1 U10643 ( .A1(n9425), .A2(n9774), .B1(n9775), .B2(n9776), .ZN(n9426)
         );
  AOI21_X1 U10644 ( .B1(n9427), .B2(n9787), .A(n9426), .ZN(n9430) );
  NAND4_X1 U10645 ( .A1(n9431), .A2(n9430), .A3(n9429), .A4(n9428), .ZN(n9467)
         );
  MUX2_X1 U10646 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n9467), .S(n9813), .Z(
        P1_U3536) );
  INV_X1 U10647 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n9433) );
  MUX2_X1 U10648 ( .A(n9433), .B(n9432), .S(n9798), .Z(n9434) );
  OAI21_X1 U10649 ( .B1(n9435), .B2(n9465), .A(n9434), .ZN(P1_U3521) );
  INV_X1 U10650 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n9437) );
  MUX2_X1 U10651 ( .A(n9437), .B(n9436), .S(n9798), .Z(n9438) );
  OAI21_X1 U10652 ( .B1(n9439), .B2(n9465), .A(n9438), .ZN(P1_U3520) );
  MUX2_X1 U10653 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n9440), .S(n9798), .Z(
        P1_U3519) );
  INV_X1 U10654 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n9443) );
  MUX2_X1 U10655 ( .A(n9443), .B(n9442), .S(n9798), .Z(n9444) );
  INV_X1 U10656 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n9447) );
  MUX2_X1 U10657 ( .A(n9447), .B(n9446), .S(n9798), .Z(n9448) );
  OAI21_X1 U10658 ( .B1(n9449), .B2(n9465), .A(n9448), .ZN(P1_U3516) );
  MUX2_X1 U10659 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9450), .S(n9798), .Z(
        P1_U3515) );
  INV_X1 U10660 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n9452) );
  MUX2_X1 U10661 ( .A(n9452), .B(n9451), .S(n9798), .Z(n9453) );
  OAI21_X1 U10662 ( .B1(n9454), .B2(n9465), .A(n9453), .ZN(P1_U3514) );
  MUX2_X1 U10663 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9455), .S(n9798), .Z(
        P1_U3513) );
  MUX2_X1 U10664 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9456), .S(n9798), .Z(
        P1_U3512) );
  MUX2_X1 U10665 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9457), .S(n9798), .Z(
        P1_U3511) );
  MUX2_X1 U10666 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9458), .S(n9798), .Z(
        P1_U3510) );
  MUX2_X1 U10667 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9459), .S(n9798), .Z(
        P1_U3509) );
  MUX2_X1 U10668 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9460), .S(n9798), .Z(
        P1_U3507) );
  MUX2_X1 U10669 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9461), .S(n9798), .Z(
        P1_U3504) );
  INV_X1 U10670 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n9463) );
  MUX2_X1 U10671 ( .A(n9463), .B(n9462), .S(n9798), .Z(n9464) );
  OAI21_X1 U10672 ( .B1(n9466), .B2(n9465), .A(n9464), .ZN(P1_U3501) );
  MUX2_X1 U10673 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n9467), .S(n9798), .Z(
        P1_U3495) );
  MUX2_X1 U10674 ( .A(n9468), .B(P1_D_REG_1__SCAN_IN), .S(n9717), .Z(P1_U3440)
         );
  MUX2_X1 U10675 ( .A(n9469), .B(P1_D_REG_0__SCAN_IN), .S(n9717), .Z(P1_U3439)
         );
  NOR2_X1 U10676 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(P1_IR_REG_30__SCAN_IN), 
        .ZN(n9472) );
  NAND4_X1 U10677 ( .A1(n9472), .A2(P1_IR_REG_31__SCAN_IN), .A3(
        P1_STATE_REG_SCAN_IN), .A4(n9471), .ZN(n9474) );
  OAI22_X1 U10678 ( .A1(n9470), .A2(n9474), .B1(n9473), .B2(n9487), .ZN(n9475)
         );
  INV_X1 U10679 ( .A(n9475), .ZN(n9476) );
  OAI21_X1 U10680 ( .B1(n9477), .B2(n9481), .A(n9476), .ZN(P1_U3324) );
  OAI222_X1 U10681 ( .A1(n9482), .A2(n9487), .B1(n9481), .B2(n9480), .C1(
        P1_U3086), .C2(n9478), .ZN(P1_U3325) );
  OAI222_X1 U10682 ( .A1(n9487), .A2(n9486), .B1(P1_U3086), .B2(n9485), .C1(
        n9484), .C2(n9483), .ZN(P1_U3328) );
  INV_X1 U10683 ( .A(n9488), .ZN(n9489) );
  MUX2_X1 U10684 ( .A(n9489), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  INV_X1 U10685 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n9959) );
  AOI211_X1 U10686 ( .C1(n9492), .C2(n9491), .A(n9490), .B(n9704), .ZN(n9497)
         );
  AOI211_X1 U10687 ( .C1(n9495), .C2(n9494), .A(n9493), .B(n9687), .ZN(n9496)
         );
  AOI211_X1 U10688 ( .C1(n9707), .C2(n9498), .A(n9497), .B(n9496), .ZN(n9500)
         );
  OAI211_X1 U10689 ( .C1(n9716), .C2(n9959), .A(n9500), .B(n9499), .ZN(
        P1_U3253) );
  INV_X1 U10690 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n9949) );
  AOI21_X1 U10691 ( .B1(n9503), .B2(n9502), .A(n9501), .ZN(n9504) );
  NAND2_X1 U10692 ( .A1(n9664), .A2(n9504), .ZN(n9510) );
  AOI21_X1 U10693 ( .B1(n9507), .B2(n9506), .A(n9505), .ZN(n9508) );
  NAND2_X1 U10694 ( .A1(n9700), .A2(n9508), .ZN(n9509) );
  OAI211_X1 U10695 ( .C1(n9692), .C2(n9511), .A(n9510), .B(n9509), .ZN(n9512)
         );
  INV_X1 U10696 ( .A(n9512), .ZN(n9514) );
  OAI211_X1 U10697 ( .C1(n9716), .C2(n9949), .A(n9514), .B(n9513), .ZN(
        P1_U3250) );
  INV_X1 U10698 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n9529) );
  AOI21_X1 U10699 ( .B1(n9517), .B2(n9516), .A(n9515), .ZN(n9518) );
  NAND2_X1 U10700 ( .A1(n9700), .A2(n9518), .ZN(n9524) );
  AOI21_X1 U10701 ( .B1(n9521), .B2(n9520), .A(n9519), .ZN(n9522) );
  NAND2_X1 U10702 ( .A1(n9664), .A2(n9522), .ZN(n9523) );
  OAI211_X1 U10703 ( .C1(n9692), .C2(n9525), .A(n9524), .B(n9523), .ZN(n9526)
         );
  INV_X1 U10704 ( .A(n9526), .ZN(n9528) );
  OAI211_X1 U10705 ( .C1(n9716), .C2(n9529), .A(n9528), .B(n9527), .ZN(
        P1_U3251) );
  NOR2_X1 U10706 ( .A1(n9530), .A2(n9901), .ZN(n9532) );
  AOI211_X1 U10707 ( .C1(n9533), .C2(n9906), .A(n9532), .B(n9531), .ZN(n9538)
         );
  AOI22_X1 U10708 ( .A1(n9929), .A2(n9538), .B1(n6345), .B2(n9927), .ZN(
        P2_U3473) );
  NOR2_X1 U10709 ( .A1(n9534), .A2(n9901), .ZN(n9536) );
  AOI211_X1 U10710 ( .C1(n9537), .C2(n9906), .A(n9536), .B(n9535), .ZN(n9540)
         );
  AOI22_X1 U10711 ( .A1(n9929), .A2(n9540), .B1(n7568), .B2(n9927), .ZN(
        P2_U3472) );
  INV_X1 U10712 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n9539) );
  AOI22_X1 U10713 ( .A1(n9915), .A2(n9539), .B1(n9538), .B2(n9914), .ZN(
        P2_U3432) );
  INV_X1 U10714 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n9541) );
  AOI22_X1 U10715 ( .A1(n9915), .A2(n9541), .B1(n9540), .B2(n9914), .ZN(
        P2_U3429) );
  XNOR2_X1 U10716 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U10717 ( .A(P2_RD_REG_SCAN_IN), .B(P1_RD_REG_SCAN_IN), .ZN(U126) );
  AOI21_X1 U10718 ( .B1(n9561), .B2(n9543), .A(n9542), .ZN(n9567) );
  OAI21_X1 U10719 ( .B1(n9561), .B2(P1_REG1_REG_0__SCAN_IN), .A(n9567), .ZN(
        n9545) );
  XNOR2_X1 U10720 ( .A(n9545), .B(n9544), .ZN(n9548) );
  AOI22_X1 U10721 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(n9581), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n9546) );
  OAI21_X1 U10722 ( .B1(n9548), .B2(n9547), .A(n9546), .ZN(P1_U3243) );
  AOI22_X1 U10723 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(n9581), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n9569) );
  INV_X1 U10724 ( .A(n9549), .ZN(n9552) );
  AOI211_X1 U10725 ( .C1(n9552), .C2(n9551), .A(n9550), .B(n9704), .ZN(n9559)
         );
  INV_X1 U10726 ( .A(n9553), .ZN(n9557) );
  INV_X1 U10727 ( .A(n9554), .ZN(n9556) );
  AOI211_X1 U10728 ( .C1(n9557), .C2(n9556), .A(n9555), .B(n9687), .ZN(n9558)
         );
  AOI211_X1 U10729 ( .C1(n9707), .C2(n9560), .A(n9559), .B(n9558), .ZN(n9568)
         );
  MUX2_X1 U10730 ( .A(n9563), .B(n9562), .S(n9561), .Z(n9565) );
  NAND2_X1 U10731 ( .A1(n9565), .A2(n9564), .ZN(n9566) );
  OAI211_X1 U10732 ( .C1(P1_IR_REG_0__SCAN_IN), .C2(n9567), .A(n9566), .B(
        P1_U3973), .ZN(n9583) );
  NAND3_X1 U10733 ( .A1(n9569), .A2(n9568), .A3(n9583), .ZN(P1_U3245) );
  OAI211_X1 U10734 ( .C1(n9572), .C2(n9571), .A(n9664), .B(n9570), .ZN(n9578)
         );
  INV_X1 U10735 ( .A(n9573), .ZN(n9574) );
  OAI211_X1 U10736 ( .C1(n9576), .C2(n9575), .A(n9700), .B(n9574), .ZN(n9577)
         );
  OAI211_X1 U10737 ( .C1(n9692), .C2(n9579), .A(n9578), .B(n9577), .ZN(n9580)
         );
  INV_X1 U10738 ( .A(n9580), .ZN(n9585) );
  NAND2_X1 U10739 ( .A1(n9581), .A2(P1_ADDR_REG_4__SCAN_IN), .ZN(n9582) );
  NAND4_X1 U10740 ( .A1(n9585), .A2(n9584), .A3(n9583), .A4(n9582), .ZN(
        P1_U3247) );
  INV_X1 U10741 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n9600) );
  AOI21_X1 U10742 ( .B1(n9588), .B2(n9587), .A(n9586), .ZN(n9589) );
  NAND2_X1 U10743 ( .A1(n9700), .A2(n9589), .ZN(n9595) );
  AOI21_X1 U10744 ( .B1(n9592), .B2(n9591), .A(n9590), .ZN(n9593) );
  NAND2_X1 U10745 ( .A1(n9664), .A2(n9593), .ZN(n9594) );
  OAI211_X1 U10746 ( .C1(n9692), .C2(n9596), .A(n9595), .B(n9594), .ZN(n9597)
         );
  INV_X1 U10747 ( .A(n9597), .ZN(n9599) );
  OAI211_X1 U10748 ( .C1(n9716), .C2(n9600), .A(n9599), .B(n9598), .ZN(
        P1_U3248) );
  INV_X1 U10749 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n9945) );
  AOI21_X1 U10750 ( .B1(n9603), .B2(n9602), .A(n9601), .ZN(n9604) );
  NAND2_X1 U10751 ( .A1(n9664), .A2(n9604), .ZN(n9610) );
  AOI21_X1 U10752 ( .B1(n9607), .B2(n9606), .A(n9605), .ZN(n9608) );
  NAND2_X1 U10753 ( .A1(n9700), .A2(n9608), .ZN(n9609) );
  OAI211_X1 U10754 ( .C1(n9692), .C2(n9611), .A(n9610), .B(n9609), .ZN(n9612)
         );
  INV_X1 U10755 ( .A(n9612), .ZN(n9614) );
  OAI211_X1 U10756 ( .C1(n9716), .C2(n9945), .A(n9614), .B(n9613), .ZN(
        P1_U3249) );
  INV_X1 U10757 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n9963) );
  AOI21_X1 U10758 ( .B1(n9617), .B2(n9616), .A(n9615), .ZN(n9618) );
  NAND2_X1 U10759 ( .A1(n9664), .A2(n9618), .ZN(n9624) );
  AOI21_X1 U10760 ( .B1(n9621), .B2(n9620), .A(n9619), .ZN(n9622) );
  NAND2_X1 U10761 ( .A1(n9700), .A2(n9622), .ZN(n9623) );
  OAI211_X1 U10762 ( .C1(n9692), .C2(n9625), .A(n9624), .B(n9623), .ZN(n9626)
         );
  INV_X1 U10763 ( .A(n9626), .ZN(n9628) );
  OAI211_X1 U10764 ( .C1(n9716), .C2(n9963), .A(n9628), .B(n9627), .ZN(
        P1_U3254) );
  INV_X1 U10765 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n9967) );
  INV_X1 U10766 ( .A(n9629), .ZN(n9640) );
  OAI21_X1 U10767 ( .B1(n9632), .B2(n9631), .A(n9630), .ZN(n9633) );
  NAND2_X1 U10768 ( .A1(n9700), .A2(n9633), .ZN(n9639) );
  OAI21_X1 U10769 ( .B1(n9636), .B2(n9635), .A(n9634), .ZN(n9637) );
  NAND2_X1 U10770 ( .A1(n9664), .A2(n9637), .ZN(n9638) );
  OAI211_X1 U10771 ( .C1(n9692), .C2(n9640), .A(n9639), .B(n9638), .ZN(n9641)
         );
  INV_X1 U10772 ( .A(n9641), .ZN(n9643) );
  OAI211_X1 U10773 ( .C1(n9716), .C2(n9967), .A(n9643), .B(n9642), .ZN(
        P1_U3255) );
  INV_X1 U10774 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n9971) );
  INV_X1 U10775 ( .A(n9644), .ZN(n9655) );
  AOI21_X1 U10776 ( .B1(n9647), .B2(n9646), .A(n9645), .ZN(n9648) );
  NAND2_X1 U10777 ( .A1(n9700), .A2(n9648), .ZN(n9654) );
  AOI21_X1 U10778 ( .B1(n9651), .B2(n9650), .A(n9649), .ZN(n9652) );
  NAND2_X1 U10779 ( .A1(n9664), .A2(n9652), .ZN(n9653) );
  OAI211_X1 U10780 ( .C1(n9692), .C2(n9655), .A(n9654), .B(n9653), .ZN(n9656)
         );
  INV_X1 U10781 ( .A(n9656), .ZN(n9658) );
  OAI211_X1 U10782 ( .C1(n9716), .C2(n9971), .A(n9658), .B(n9657), .ZN(
        P1_U3256) );
  INV_X1 U10783 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n9675) );
  INV_X1 U10784 ( .A(n9659), .ZN(n9671) );
  AOI21_X1 U10785 ( .B1(n9662), .B2(n9661), .A(n9660), .ZN(n9663) );
  NAND2_X1 U10786 ( .A1(n9664), .A2(n9663), .ZN(n9670) );
  AOI21_X1 U10787 ( .B1(n9667), .B2(n9666), .A(n9665), .ZN(n9668) );
  NAND2_X1 U10788 ( .A1(n9700), .A2(n9668), .ZN(n9669) );
  OAI211_X1 U10789 ( .C1(n9692), .C2(n9671), .A(n9670), .B(n9669), .ZN(n9672)
         );
  INV_X1 U10790 ( .A(n9672), .ZN(n9674) );
  OAI211_X1 U10791 ( .C1(n9716), .C2(n9675), .A(n9674), .B(n9673), .ZN(
        P1_U3257) );
  INV_X1 U10792 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n9977) );
  AOI211_X1 U10793 ( .C1(n9678), .C2(n9677), .A(n9676), .B(n9704), .ZN(n9683)
         );
  AOI211_X1 U10794 ( .C1(n9681), .C2(n9680), .A(n9679), .B(n9687), .ZN(n9682)
         );
  AOI211_X1 U10795 ( .C1(n9707), .C2(n9684), .A(n9683), .B(n9682), .ZN(n9686)
         );
  OAI211_X1 U10796 ( .C1(n9716), .C2(n9977), .A(n9686), .B(n9685), .ZN(
        P1_U3258) );
  INV_X1 U10797 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n9981) );
  AOI21_X1 U10798 ( .B1(n9689), .B2(n9688), .A(n9687), .ZN(n9697) );
  XOR2_X1 U10799 ( .A(n9691), .B(n9690), .Z(n9694) );
  OAI22_X1 U10800 ( .A1(n9694), .A2(n9704), .B1(n9693), .B2(n9692), .ZN(n9695)
         );
  AOI21_X1 U10801 ( .B1(n9697), .B2(n9696), .A(n9695), .ZN(n9699) );
  OAI211_X1 U10802 ( .C1(n9716), .C2(n9981), .A(n9699), .B(n9698), .ZN(
        P1_U3259) );
  INV_X1 U10803 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n9715) );
  OAI211_X1 U10804 ( .C1(n9703), .C2(n9702), .A(n9701), .B(n9700), .ZN(n9712)
         );
  AOI21_X1 U10805 ( .B1(n9706), .B2(n9705), .A(n9704), .ZN(n9710) );
  AOI22_X1 U10806 ( .A1(n9710), .A2(n9709), .B1(n9708), .B2(n9707), .ZN(n9711)
         );
  AND2_X1 U10807 ( .A1(n9712), .A2(n9711), .ZN(n9714) );
  OAI211_X1 U10808 ( .C1(n9716), .C2(n9715), .A(n9714), .B(n9713), .ZN(
        P1_U3261) );
  AND2_X1 U10809 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n9717), .ZN(P1_U3294) );
  AND2_X1 U10810 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n9717), .ZN(P1_U3295) );
  AND2_X1 U10811 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n9717), .ZN(P1_U3296) );
  AND2_X1 U10812 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n9717), .ZN(P1_U3297) );
  AND2_X1 U10813 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n9717), .ZN(P1_U3298) );
  AND2_X1 U10814 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n9717), .ZN(P1_U3299) );
  AND2_X1 U10815 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n9717), .ZN(P1_U3300) );
  AND2_X1 U10816 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9717), .ZN(P1_U3301) );
  AND2_X1 U10817 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n9717), .ZN(P1_U3302) );
  AND2_X1 U10818 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n9717), .ZN(P1_U3303) );
  AND2_X1 U10819 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n9717), .ZN(P1_U3304) );
  AND2_X1 U10820 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n9717), .ZN(P1_U3305) );
  AND2_X1 U10821 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n9717), .ZN(P1_U3306) );
  AND2_X1 U10822 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n9717), .ZN(P1_U3307) );
  AND2_X1 U10823 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n9717), .ZN(P1_U3308) );
  AND2_X1 U10824 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n9717), .ZN(P1_U3309) );
  AND2_X1 U10825 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n9717), .ZN(P1_U3310) );
  AND2_X1 U10826 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n9717), .ZN(P1_U3311) );
  AND2_X1 U10827 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n9717), .ZN(P1_U3312) );
  AND2_X1 U10828 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n9717), .ZN(P1_U3313) );
  AND2_X1 U10829 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n9717), .ZN(P1_U3314) );
  AND2_X1 U10830 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n9717), .ZN(P1_U3315) );
  AND2_X1 U10831 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n9717), .ZN(P1_U3316) );
  AND2_X1 U10832 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n9717), .ZN(P1_U3317) );
  AND2_X1 U10833 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n9717), .ZN(P1_U3318) );
  AND2_X1 U10834 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n9717), .ZN(P1_U3319) );
  AND2_X1 U10835 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n9717), .ZN(P1_U3320) );
  AND2_X1 U10836 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n9717), .ZN(P1_U3321) );
  AND2_X1 U10837 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n9717), .ZN(P1_U3322) );
  AND2_X1 U10838 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n9717), .ZN(P1_U3323) );
  NAND2_X1 U10839 ( .A1(n9760), .A2(n9783), .ZN(n9723) );
  INV_X1 U10840 ( .A(n9718), .ZN(n9722) );
  AOI222_X1 U10841 ( .A1(n9723), .A2(n9722), .B1(n9721), .B2(n9720), .C1(n9719), .C2(n9757), .ZN(n9800) );
  INV_X1 U10842 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n9724) );
  AOI22_X1 U10843 ( .A1(n9798), .A2(n9800), .B1(n9724), .B2(n9796), .ZN(
        P1_U3453) );
  OAI21_X1 U10844 ( .B1(n9726), .B2(n9768), .A(n9725), .ZN(n9727) );
  AOI21_X1 U10845 ( .B1(n9728), .B2(n9794), .A(n9727), .ZN(n9730) );
  AND2_X1 U10846 ( .A1(n9730), .A2(n9729), .ZN(n9802) );
  INV_X1 U10847 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n9731) );
  AOI22_X1 U10848 ( .A1(n9798), .A2(n9802), .B1(n9731), .B2(n9796), .ZN(
        P1_U3459) );
  OAI21_X1 U10849 ( .B1(n9733), .B2(n9768), .A(n9732), .ZN(n9735) );
  AOI211_X1 U10850 ( .C1(n9794), .C2(n9736), .A(n9735), .B(n9734), .ZN(n9803)
         );
  INV_X1 U10851 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n9737) );
  AOI22_X1 U10852 ( .A1(n9798), .A2(n9803), .B1(n9737), .B2(n9796), .ZN(
        P1_U3471) );
  INV_X1 U10853 ( .A(n9738), .ZN(n9741) );
  OAI21_X1 U10854 ( .B1(n4596), .B2(n9768), .A(n9739), .ZN(n9740) );
  AOI21_X1 U10855 ( .B1(n9742), .B2(n9741), .A(n9740), .ZN(n9743) );
  AND2_X1 U10856 ( .A1(n9744), .A2(n9743), .ZN(n9805) );
  INV_X1 U10857 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n9745) );
  AOI22_X1 U10858 ( .A1(n9798), .A2(n9805), .B1(n9745), .B2(n9796), .ZN(
        P1_U3477) );
  AOI22_X1 U10859 ( .A1(n9747), .A2(n9787), .B1(n9746), .B2(n9754), .ZN(n9748)
         );
  OAI211_X1 U10860 ( .C1(n9750), .C2(n9783), .A(n9749), .B(n9748), .ZN(n9751)
         );
  AOI21_X1 U10861 ( .B1(n9794), .B2(n9752), .A(n9751), .ZN(n9807) );
  INV_X1 U10862 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n9753) );
  AOI22_X1 U10863 ( .A1(n9798), .A2(n9807), .B1(n9753), .B2(n9796), .ZN(
        P1_U3480) );
  AOI22_X1 U10864 ( .A1(n9757), .A2(n9756), .B1(n9755), .B2(n9754), .ZN(n9758)
         );
  OAI211_X1 U10865 ( .C1(n4937), .C2(n9768), .A(n9759), .B(n9758), .ZN(n9763)
         );
  NOR2_X1 U10866 ( .A1(n9761), .A2(n9760), .ZN(n9762) );
  AOI211_X1 U10867 ( .C1(n9765), .C2(n9764), .A(n9763), .B(n9762), .ZN(n9808)
         );
  INV_X1 U10868 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n9766) );
  AOI22_X1 U10869 ( .A1(n9798), .A2(n9808), .B1(n9766), .B2(n9796), .ZN(
        P1_U3483) );
  OAI21_X1 U10870 ( .B1(n9769), .B2(n9768), .A(n9767), .ZN(n9770) );
  AOI211_X1 U10871 ( .C1(n9772), .C2(n9794), .A(n9771), .B(n9770), .ZN(n9809)
         );
  INV_X1 U10872 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n9773) );
  AOI22_X1 U10873 ( .A1(n9798), .A2(n9809), .B1(n9773), .B2(n9796), .ZN(
        P1_U3486) );
  OAI22_X1 U10874 ( .A1(n9777), .A2(n9776), .B1(n9775), .B2(n9774), .ZN(n9779)
         );
  AOI211_X1 U10875 ( .C1(n9787), .C2(n9780), .A(n9779), .B(n9778), .ZN(n9781)
         );
  OAI21_X1 U10876 ( .B1(n9783), .B2(n9782), .A(n9781), .ZN(n9784) );
  AOI21_X1 U10877 ( .B1(n9785), .B2(n9794), .A(n9784), .ZN(n9810) );
  INV_X1 U10878 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n9786) );
  AOI22_X1 U10879 ( .A1(n9798), .A2(n9810), .B1(n9786), .B2(n9796), .ZN(
        P1_U3489) );
  NAND2_X1 U10880 ( .A1(n9788), .A2(n9787), .ZN(n9789) );
  OAI211_X1 U10881 ( .C1(n9792), .C2(n9791), .A(n9790), .B(n9789), .ZN(n9793)
         );
  AOI21_X1 U10882 ( .B1(n9795), .B2(n9794), .A(n9793), .ZN(n9812) );
  INV_X1 U10883 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n9797) );
  AOI22_X1 U10884 ( .A1(n9798), .A2(n9812), .B1(n9797), .B2(n9796), .ZN(
        P1_U3492) );
  INV_X1 U10885 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n9799) );
  AOI22_X1 U10886 ( .A1(n9813), .A2(n9800), .B1(n9799), .B2(n9811), .ZN(
        P1_U3522) );
  INV_X1 U10887 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n9801) );
  AOI22_X1 U10888 ( .A1(n9813), .A2(n9802), .B1(n9801), .B2(n9811), .ZN(
        P1_U3524) );
  AOI22_X1 U10889 ( .A1(n9813), .A2(n9803), .B1(n9018), .B2(n9811), .ZN(
        P1_U3528) );
  INV_X1 U10890 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n9804) );
  AOI22_X1 U10891 ( .A1(n9813), .A2(n9805), .B1(n9804), .B2(n9811), .ZN(
        P1_U3530) );
  INV_X1 U10892 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n9806) );
  AOI22_X1 U10893 ( .A1(n9813), .A2(n9807), .B1(n9806), .B2(n9811), .ZN(
        P1_U3531) );
  AOI22_X1 U10894 ( .A1(n9813), .A2(n9808), .B1(n9034), .B2(n9811), .ZN(
        P1_U3532) );
  AOI22_X1 U10895 ( .A1(n9813), .A2(n9809), .B1(n9036), .B2(n9811), .ZN(
        P1_U3533) );
  AOI22_X1 U10896 ( .A1(n9813), .A2(n9810), .B1(n9037), .B2(n9811), .ZN(
        P1_U3534) );
  AOI22_X1 U10897 ( .A1(n9813), .A2(n9812), .B1(n9033), .B2(n9811), .ZN(
        P1_U3535) );
  AOI22_X1 U10898 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(n9845), .B1(
        P2_REG3_REG_14__SCAN_IN), .B2(P2_U3151), .ZN(n9827) );
  AOI21_X1 U10899 ( .B1(n9816), .B2(n9815), .A(n9814), .ZN(n9824) );
  XOR2_X1 U10900 ( .A(n9818), .B(n9817), .Z(n9823) );
  AOI21_X1 U10901 ( .B1(n9821), .B2(n9820), .A(n9819), .ZN(n9822) );
  OAI222_X1 U10902 ( .A1(n9860), .A2(n9824), .B1(n9858), .B2(n9823), .C1(n9856), .C2(n9822), .ZN(n9825) );
  INV_X1 U10903 ( .A(n9825), .ZN(n9826) );
  OAI211_X1 U10904 ( .C1(n9844), .C2(n9828), .A(n9827), .B(n9826), .ZN(
        P2_U3196) );
  AOI22_X1 U10905 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(n9845), .B1(
        P2_REG3_REG_16__SCAN_IN), .B2(P2_U3151), .ZN(n9842) );
  AOI21_X1 U10906 ( .B1(n9831), .B2(n9830), .A(n9829), .ZN(n9839) );
  XOR2_X1 U10907 ( .A(n9833), .B(n9832), .Z(n9838) );
  AOI21_X1 U10908 ( .B1(n9836), .B2(n9835), .A(n9834), .ZN(n9837) );
  OAI222_X1 U10909 ( .A1(n9860), .A2(n9839), .B1(n9858), .B2(n9838), .C1(n9856), .C2(n9837), .ZN(n9840) );
  INV_X1 U10910 ( .A(n9840), .ZN(n9841) );
  OAI211_X1 U10911 ( .C1(n9844), .C2(n9843), .A(n9842), .B(n9841), .ZN(
        P2_U3198) );
  AOI22_X1 U10912 ( .A1(n9847), .A2(n9846), .B1(n9845), .B2(
        P2_ADDR_REG_17__SCAN_IN), .ZN(n9863) );
  AOI21_X1 U10913 ( .B1(n9850), .B2(n9849), .A(n9848), .ZN(n9859) );
  XOR2_X1 U10914 ( .A(n9852), .B(n9851), .Z(n9857) );
  AOI21_X1 U10915 ( .B1(n8565), .B2(n9854), .A(n9853), .ZN(n9855) );
  OAI222_X1 U10916 ( .A1(n9860), .A2(n9859), .B1(n9858), .B2(n9857), .C1(n9856), .C2(n9855), .ZN(n9861) );
  INV_X1 U10917 ( .A(n9861), .ZN(n9862) );
  OAI211_X1 U10918 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n6128), .A(n9863), .B(
        n9862), .ZN(P2_U3199) );
  INV_X1 U10919 ( .A(n9864), .ZN(n9868) );
  OAI22_X1 U10920 ( .A1(n9866), .A2(n9908), .B1(n9865), .B2(n9901), .ZN(n9867)
         );
  NOR2_X1 U10921 ( .A1(n9868), .A2(n9867), .ZN(n9916) );
  AOI22_X1 U10922 ( .A1(n9915), .A2(n6169), .B1(n9916), .B2(n9914), .ZN(
        P2_U3393) );
  INV_X1 U10923 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n9874) );
  OAI22_X1 U10924 ( .A1(n9871), .A2(n9870), .B1(n9869), .B2(n9901), .ZN(n9872)
         );
  NOR2_X1 U10925 ( .A1(n9873), .A2(n9872), .ZN(n9917) );
  AOI22_X1 U10926 ( .A1(n9915), .A2(n9874), .B1(n9917), .B2(n9914), .ZN(
        P2_U3396) );
  NOR2_X1 U10927 ( .A1(n9875), .A2(n9901), .ZN(n9877) );
  AOI211_X1 U10928 ( .C1(n9906), .C2(n9878), .A(n9877), .B(n9876), .ZN(n9918)
         );
  AOI22_X1 U10929 ( .A1(n9915), .A2(n6215), .B1(n9918), .B2(n9914), .ZN(
        P2_U3402) );
  INV_X1 U10930 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n9883) );
  NOR2_X1 U10931 ( .A1(n9879), .A2(n9901), .ZN(n9881) );
  AOI211_X1 U10932 ( .C1(n9882), .C2(n9906), .A(n9881), .B(n9880), .ZN(n9920)
         );
  AOI22_X1 U10933 ( .A1(n9915), .A2(n9883), .B1(n9920), .B2(n9914), .ZN(
        P2_U3408) );
  INV_X1 U10934 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n9888) );
  NOR2_X1 U10935 ( .A1(n9884), .A2(n9901), .ZN(n9886) );
  AOI211_X1 U10936 ( .C1(n9887), .C2(n9898), .A(n9886), .B(n9885), .ZN(n9921)
         );
  AOI22_X1 U10937 ( .A1(n9915), .A2(n9888), .B1(n9921), .B2(n9914), .ZN(
        P2_U3411) );
  INV_X1 U10938 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n9894) );
  NAND2_X1 U10939 ( .A1(n9889), .A2(n9906), .ZN(n9892) );
  OR2_X1 U10940 ( .A1(n9890), .A2(n9901), .ZN(n9891) );
  AOI22_X1 U10941 ( .A1(n9915), .A2(n9894), .B1(n9923), .B2(n9914), .ZN(
        P2_U3414) );
  INV_X1 U10942 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n9900) );
  NOR2_X1 U10943 ( .A1(n9895), .A2(n9901), .ZN(n9897) );
  AOI211_X1 U10944 ( .C1(n9899), .C2(n9898), .A(n9897), .B(n9896), .ZN(n9925)
         );
  AOI22_X1 U10945 ( .A1(n9915), .A2(n9900), .B1(n9925), .B2(n9914), .ZN(
        P2_U3420) );
  INV_X1 U10946 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n9907) );
  NOR2_X1 U10947 ( .A1(n9902), .A2(n9901), .ZN(n9904) );
  AOI211_X1 U10948 ( .C1(n9906), .C2(n9905), .A(n9904), .B(n9903), .ZN(n9926)
         );
  AOI22_X1 U10949 ( .A1(n9915), .A2(n9907), .B1(n9926), .B2(n9914), .ZN(
        P2_U3423) );
  NOR2_X1 U10950 ( .A1(n9909), .A2(n9908), .ZN(n9911) );
  AOI211_X1 U10951 ( .C1(n9913), .C2(n9912), .A(n9911), .B(n9910), .ZN(n9928)
         );
  AOI22_X1 U10952 ( .A1(n9915), .A2(n6322), .B1(n9928), .B2(n9914), .ZN(
        P2_U3426) );
  AOI22_X1 U10953 ( .A1(n9929), .A2(n9916), .B1(n6871), .B2(n9927), .ZN(
        P2_U3460) );
  AOI22_X1 U10954 ( .A1(n9929), .A2(n9917), .B1(n6187), .B2(n9927), .ZN(
        P2_U3461) );
  AOI22_X1 U10955 ( .A1(n9929), .A2(n9918), .B1(n6898), .B2(n9927), .ZN(
        P2_U3463) );
  INV_X1 U10956 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n9919) );
  AOI22_X1 U10957 ( .A1(n9929), .A2(n9920), .B1(n9919), .B2(n9927), .ZN(
        P2_U3465) );
  AOI22_X1 U10958 ( .A1(n9929), .A2(n9921), .B1(n6969), .B2(n9927), .ZN(
        P2_U3466) );
  AOI22_X1 U10959 ( .A1(n9929), .A2(n9923), .B1(n9922), .B2(n9927), .ZN(
        P2_U3467) );
  AOI22_X1 U10960 ( .A1(n9929), .A2(n9925), .B1(n9924), .B2(n9927), .ZN(
        P2_U3469) );
  AOI22_X1 U10961 ( .A1(n9929), .A2(n9926), .B1(n6306), .B2(n9927), .ZN(
        P2_U3470) );
  AOI22_X1 U10962 ( .A1(n9929), .A2(n9928), .B1(n7578), .B2(n9927), .ZN(
        P2_U3471) );
  AOI21_X1 U10963 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(P2_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n9935) );
  INV_X1 U10964 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n9931) );
  NAND2_X1 U10965 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .ZN(n9930) );
  NOR2_X1 U10966 ( .A1(n9931), .A2(n9930), .ZN(n9933) );
  NOR2_X1 U10967 ( .A1(n9935), .A2(n9933), .ZN(n9932) );
  XOR2_X1 U10968 ( .A(P2_ADDR_REG_1__SCAN_IN), .B(n9932), .Z(ADD_1068_U5) );
  XOR2_X1 U10969 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1068_U46) );
  NOR2_X1 U10970 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n9985) );
  NOR2_X1 U10971 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n9983) );
  NOR2_X1 U10972 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n9979) );
  NOR2_X1 U10973 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n9975) );
  NOR2_X1 U10974 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n9973) );
  NOR2_X1 U10975 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n9969) );
  NOR2_X1 U10976 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n9965) );
  NOR2_X1 U10977 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n9961) );
  NOR2_X1 U10978 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n9957) );
  NOR2_X1 U10979 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n9953) );
  NOR2_X1 U10980 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n9951) );
  NOR2_X1 U10981 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n9947) );
  NOR2_X1 U10982 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(P2_ADDR_REG_5__SCAN_IN), 
        .ZN(n9943) );
  NOR2_X1 U10983 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n9941) );
  NAND2_X1 U10984 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n9939) );
  XOR2_X1 U10985 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(P2_ADDR_REG_3__SCAN_IN), .Z(
        n10216) );
  NAND2_X1 U10986 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n9937) );
  NOR2_X1 U10987 ( .A1(P2_ADDR_REG_1__SCAN_IN), .A2(n9933), .ZN(n9934) );
  NOR2_X1 U10988 ( .A1(n9935), .A2(n9934), .ZN(n10204) );
  XOR2_X1 U10989 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(P2_ADDR_REG_2__SCAN_IN), .Z(
        n10203) );
  NAND2_X1 U10990 ( .A1(n10204), .A2(n10203), .ZN(n9936) );
  NAND2_X1 U10991 ( .A1(n9937), .A2(n9936), .ZN(n10215) );
  NAND2_X1 U10992 ( .A1(n10216), .A2(n10215), .ZN(n9938) );
  NAND2_X1 U10993 ( .A1(n9939), .A2(n9938), .ZN(n10218) );
  XNOR2_X1 U10994 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10217) );
  NOR2_X1 U10995 ( .A1(n10218), .A2(n10217), .ZN(n9940) );
  NOR2_X1 U10996 ( .A1(n9941), .A2(n9940), .ZN(n10214) );
  XNOR2_X1 U10997 ( .A(P1_ADDR_REG_5__SCAN_IN), .B(P2_ADDR_REG_5__SCAN_IN), 
        .ZN(n10213) );
  NOR2_X1 U10998 ( .A1(n10214), .A2(n10213), .ZN(n9942) );
  NOR2_X1 U10999 ( .A1(n9943), .A2(n9942), .ZN(n10212) );
  AOI22_X1 U11000 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(n9945), .B1(
        P1_ADDR_REG_6__SCAN_IN), .B2(n9944), .ZN(n10211) );
  NOR2_X1 U11001 ( .A1(n10212), .A2(n10211), .ZN(n9946) );
  NOR2_X1 U11002 ( .A1(n9947), .A2(n9946), .ZN(n10210) );
  AOI22_X1 U11003 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n9949), .B1(
        P1_ADDR_REG_7__SCAN_IN), .B2(n9948), .ZN(n10209) );
  NOR2_X1 U11004 ( .A1(n10210), .A2(n10209), .ZN(n9950) );
  NOR2_X1 U11005 ( .A1(n9951), .A2(n9950), .ZN(n10208) );
  XNOR2_X1 U11006 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n10207) );
  NOR2_X1 U11007 ( .A1(n10208), .A2(n10207), .ZN(n9952) );
  NOR2_X1 U11008 ( .A1(n9953), .A2(n9952), .ZN(n10206) );
  INV_X1 U11009 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n9955) );
  AOI22_X1 U11010 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n9955), .B1(
        P1_ADDR_REG_9__SCAN_IN), .B2(n9954), .ZN(n10205) );
  NOR2_X1 U11011 ( .A1(n10206), .A2(n10205), .ZN(n9956) );
  NOR2_X1 U11012 ( .A1(n9957), .A2(n9956), .ZN(n10003) );
  AOI22_X1 U11013 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(n9959), .B1(
        P1_ADDR_REG_10__SCAN_IN), .B2(n9958), .ZN(n10002) );
  NOR2_X1 U11014 ( .A1(n10003), .A2(n10002), .ZN(n9960) );
  NOR2_X1 U11015 ( .A1(n9961), .A2(n9960), .ZN(n10001) );
  AOI22_X1 U11016 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(n9963), .B1(
        P1_ADDR_REG_11__SCAN_IN), .B2(n9962), .ZN(n10000) );
  NOR2_X1 U11017 ( .A1(n10001), .A2(n10000), .ZN(n9964) );
  NOR2_X1 U11018 ( .A1(n9965), .A2(n9964), .ZN(n9999) );
  AOI22_X1 U11019 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(n9967), .B1(
        P1_ADDR_REG_12__SCAN_IN), .B2(n9966), .ZN(n9998) );
  NOR2_X1 U11020 ( .A1(n9999), .A2(n9998), .ZN(n9968) );
  NOR2_X1 U11021 ( .A1(n9969), .A2(n9968), .ZN(n9997) );
  AOI22_X1 U11022 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(n9971), .B1(
        P1_ADDR_REG_13__SCAN_IN), .B2(n9970), .ZN(n9996) );
  NOR2_X1 U11023 ( .A1(n9997), .A2(n9996), .ZN(n9972) );
  NOR2_X1 U11024 ( .A1(n9973), .A2(n9972), .ZN(n9995) );
  XNOR2_X1 U11025 ( .A(P2_ADDR_REG_14__SCAN_IN), .B(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n9994) );
  NOR2_X1 U11026 ( .A1(n9995), .A2(n9994), .ZN(n9974) );
  NOR2_X1 U11027 ( .A1(n9975), .A2(n9974), .ZN(n9993) );
  AOI22_X1 U11028 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(n9977), .B1(
        P1_ADDR_REG_15__SCAN_IN), .B2(n9976), .ZN(n9992) );
  NOR2_X1 U11029 ( .A1(n9993), .A2(n9992), .ZN(n9978) );
  NOR2_X1 U11030 ( .A1(n9979), .A2(n9978), .ZN(n9991) );
  INV_X1 U11031 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n9980) );
  AOI22_X1 U11032 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(n9981), .B1(
        P1_ADDR_REG_16__SCAN_IN), .B2(n9980), .ZN(n9990) );
  NOR2_X1 U11033 ( .A1(n9991), .A2(n9990), .ZN(n9982) );
  NOR2_X1 U11034 ( .A1(n9983), .A2(n9982), .ZN(n9989) );
  XNOR2_X1 U11035 ( .A(P2_ADDR_REG_17__SCAN_IN), .B(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n9988) );
  NOR2_X1 U11036 ( .A1(n9989), .A2(n9988), .ZN(n9984) );
  NOR2_X1 U11037 ( .A1(n9985), .A2(n9984), .ZN(n9986) );
  NOR2_X1 U11038 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n9986), .ZN(n10006) );
  AND2_X1 U11039 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n9986), .ZN(n10004) );
  NOR2_X1 U11040 ( .A1(n10006), .A2(n10004), .ZN(n9987) );
  XOR2_X1 U11041 ( .A(P2_ADDR_REG_18__SCAN_IN), .B(n9987), .Z(ADD_1068_U55) );
  XNOR2_X1 U11042 ( .A(n9989), .B(n9988), .ZN(ADD_1068_U56) );
  XNOR2_X1 U11043 ( .A(n9991), .B(n9990), .ZN(ADD_1068_U57) );
  XNOR2_X1 U11044 ( .A(n9993), .B(n9992), .ZN(ADD_1068_U58) );
  XNOR2_X1 U11045 ( .A(n9995), .B(n9994), .ZN(ADD_1068_U59) );
  XNOR2_X1 U11046 ( .A(n9997), .B(n9996), .ZN(ADD_1068_U60) );
  XNOR2_X1 U11047 ( .A(n9999), .B(n9998), .ZN(ADD_1068_U61) );
  XNOR2_X1 U11048 ( .A(n10001), .B(n10000), .ZN(ADD_1068_U62) );
  XNOR2_X1 U11049 ( .A(n10003), .B(n10002), .ZN(ADD_1068_U63) );
  NOR2_X1 U11050 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(n10004), .ZN(n10005) );
  NOR2_X1 U11051 ( .A1(n10006), .A2(n10005), .ZN(n10202) );
  XNOR2_X1 U11052 ( .A(P1_ADDR_REG_19__SCAN_IN), .B(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n10200) );
  AOI22_X1 U11053 ( .A1(SI_31_), .A2(keyinput_f1), .B1(SI_27_), .B2(
        keyinput_f5), .ZN(n10007) );
  OAI221_X1 U11054 ( .B1(SI_31_), .B2(keyinput_f1), .C1(SI_27_), .C2(
        keyinput_f5), .A(n10007), .ZN(n10014) );
  AOI22_X1 U11055 ( .A1(SI_28_), .A2(keyinput_f4), .B1(SI_23_), .B2(
        keyinput_f9), .ZN(n10008) );
  OAI221_X1 U11056 ( .B1(SI_28_), .B2(keyinput_f4), .C1(SI_23_), .C2(
        keyinput_f9), .A(n10008), .ZN(n10013) );
  AOI22_X1 U11057 ( .A1(P2_REG3_REG_20__SCAN_IN), .A2(keyinput_f55), .B1(
        P2_REG3_REG_28__SCAN_IN), .B2(keyinput_f42), .ZN(n10009) );
  OAI221_X1 U11058 ( .B1(P2_REG3_REG_20__SCAN_IN), .B2(keyinput_f55), .C1(
        P2_REG3_REG_28__SCAN_IN), .C2(keyinput_f42), .A(n10009), .ZN(n10012)
         );
  AOI22_X1 U11059 ( .A1(P2_REG3_REG_2__SCAN_IN), .A2(keyinput_f59), .B1(SI_12_), .B2(keyinput_f20), .ZN(n10010) );
  OAI221_X1 U11060 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(keyinput_f59), .C1(
        SI_12_), .C2(keyinput_f20), .A(n10010), .ZN(n10011) );
  NOR4_X1 U11061 ( .A1(n10014), .A2(n10013), .A3(n10012), .A4(n10011), .ZN(
        n10041) );
  XOR2_X1 U11062 ( .A(SI_24_), .B(keyinput_f8), .Z(n10021) );
  AOI22_X1 U11063 ( .A1(SI_6_), .A2(keyinput_f26), .B1(SI_26_), .B2(
        keyinput_f6), .ZN(n10015) );
  OAI221_X1 U11064 ( .B1(SI_6_), .B2(keyinput_f26), .C1(SI_26_), .C2(
        keyinput_f6), .A(n10015), .ZN(n10020) );
  AOI22_X1 U11065 ( .A1(SI_30_), .A2(keyinput_f2), .B1(P2_STATE_REG_SCAN_IN), 
        .B2(keyinput_f34), .ZN(n10016) );
  OAI221_X1 U11066 ( .B1(SI_30_), .B2(keyinput_f2), .C1(P2_STATE_REG_SCAN_IN), 
        .C2(keyinput_f34), .A(n10016), .ZN(n10019) );
  AOI22_X1 U11067 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(keyinput_f39), .B1(SI_5_), .B2(keyinput_f27), .ZN(n10017) );
  OAI221_X1 U11068 ( .B1(P2_REG3_REG_10__SCAN_IN), .B2(keyinput_f39), .C1(
        SI_5_), .C2(keyinput_f27), .A(n10017), .ZN(n10018) );
  NOR4_X1 U11069 ( .A1(n10021), .A2(n10020), .A3(n10019), .A4(n10018), .ZN(
        n10040) );
  AOI22_X1 U11070 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(keyinput_f37), .B1(
        SI_19_), .B2(keyinput_f13), .ZN(n10022) );
  OAI221_X1 U11071 ( .B1(P2_REG3_REG_14__SCAN_IN), .B2(keyinput_f37), .C1(
        SI_19_), .C2(keyinput_f13), .A(n10022), .ZN(n10029) );
  AOI22_X1 U11072 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(keyinput_f56), .B1(SI_2_), .B2(keyinput_f30), .ZN(n10023) );
  OAI221_X1 U11073 ( .B1(P2_REG3_REG_13__SCAN_IN), .B2(keyinput_f56), .C1(
        SI_2_), .C2(keyinput_f30), .A(n10023), .ZN(n10028) );
  INV_X1 U11074 ( .A(SI_16_), .ZN(n10100) );
  AOI22_X1 U11075 ( .A1(n10100), .A2(keyinput_f16), .B1(keyinput_f53), .B2(
        n6124), .ZN(n10024) );
  OAI221_X1 U11076 ( .B1(n10100), .B2(keyinput_f16), .C1(n6124), .C2(
        keyinput_f53), .A(n10024), .ZN(n10027) );
  AOI22_X1 U11077 ( .A1(P2_REG3_REG_23__SCAN_IN), .A2(keyinput_f38), .B1(
        SI_17_), .B2(keyinput_f15), .ZN(n10025) );
  OAI221_X1 U11078 ( .B1(P2_REG3_REG_23__SCAN_IN), .B2(keyinput_f38), .C1(
        SI_17_), .C2(keyinput_f15), .A(n10025), .ZN(n10026) );
  NOR4_X1 U11079 ( .A1(n10029), .A2(n10028), .A3(n10027), .A4(n10026), .ZN(
        n10039) );
  AOI22_X1 U11080 ( .A1(P2_REG3_REG_26__SCAN_IN), .A2(keyinput_f62), .B1(
        P2_REG3_REG_27__SCAN_IN), .B2(keyinput_f36), .ZN(n10030) );
  OAI221_X1 U11081 ( .B1(P2_REG3_REG_26__SCAN_IN), .B2(keyinput_f62), .C1(
        P2_REG3_REG_27__SCAN_IN), .C2(keyinput_f36), .A(n10030), .ZN(n10037)
         );
  AOI22_X1 U11082 ( .A1(P2_REG3_REG_1__SCAN_IN), .A2(keyinput_f44), .B1(SI_9_), 
        .B2(keyinput_f23), .ZN(n10031) );
  OAI221_X1 U11083 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(keyinput_f44), .C1(SI_9_), .C2(keyinput_f23), .A(n10031), .ZN(n10036) );
  AOI22_X1 U11084 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(keyinput_f43), .B1(
        P2_REG3_REG_22__SCAN_IN), .B2(keyinput_f57), .ZN(n10032) );
  OAI221_X1 U11085 ( .B1(P2_REG3_REG_8__SCAN_IN), .B2(keyinput_f43), .C1(
        P2_REG3_REG_22__SCAN_IN), .C2(keyinput_f57), .A(n10032), .ZN(n10035)
         );
  AOI22_X1 U11086 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(keyinput_f49), .B1(
        P2_RD_REG_SCAN_IN), .B2(keyinput_f33), .ZN(n10033) );
  OAI221_X1 U11087 ( .B1(P2_REG3_REG_5__SCAN_IN), .B2(keyinput_f49), .C1(
        P2_RD_REG_SCAN_IN), .C2(keyinput_f33), .A(n10033), .ZN(n10034) );
  NOR4_X1 U11088 ( .A1(n10037), .A2(n10036), .A3(n10035), .A4(n10034), .ZN(
        n10038) );
  NAND4_X1 U11089 ( .A1(n10041), .A2(n10040), .A3(n10039), .A4(n10038), .ZN(
        n10093) );
  INV_X1 U11090 ( .A(SI_3_), .ZN(n10106) );
  INV_X1 U11091 ( .A(SI_7_), .ZN(n10096) );
  AOI22_X1 U11092 ( .A1(n10106), .A2(keyinput_f29), .B1(n10096), .B2(
        keyinput_f25), .ZN(n10042) );
  OAI221_X1 U11093 ( .B1(n10106), .B2(keyinput_f29), .C1(n10096), .C2(
        keyinput_f25), .A(n10042), .ZN(n10051) );
  INV_X1 U11094 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n10133) );
  INV_X1 U11095 ( .A(P2_WR_REG_SCAN_IN), .ZN(n10102) );
  AOI22_X1 U11096 ( .A1(n10133), .A2(keyinput_f48), .B1(keyinput_f0), .B2(
        n10102), .ZN(n10043) );
  OAI221_X1 U11097 ( .B1(n10133), .B2(keyinput_f48), .C1(n10102), .C2(
        keyinput_f0), .A(n10043), .ZN(n10050) );
  AOI22_X1 U11098 ( .A1(n10045), .A2(keyinput_f41), .B1(n10132), .B2(
        keyinput_f21), .ZN(n10044) );
  OAI221_X1 U11099 ( .B1(n10045), .B2(keyinput_f41), .C1(n10132), .C2(
        keyinput_f21), .A(n10044), .ZN(n10049) );
  INV_X1 U11100 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n10099) );
  AOI22_X1 U11101 ( .A1(n10099), .A2(keyinput_f60), .B1(keyinput_f3), .B2(
        n10047), .ZN(n10046) );
  OAI221_X1 U11102 ( .B1(n10099), .B2(keyinput_f60), .C1(n10047), .C2(
        keyinput_f3), .A(n10046), .ZN(n10048) );
  NOR4_X1 U11103 ( .A1(n10051), .A2(n10050), .A3(n10049), .A4(n10048), .ZN(
        n10091) );
  AOI22_X1 U11104 ( .A1(n10053), .A2(keyinput_f22), .B1(keyinput_f52), .B2(
        n10128), .ZN(n10052) );
  OAI221_X1 U11105 ( .B1(n10053), .B2(keyinput_f22), .C1(n10128), .C2(
        keyinput_f52), .A(n10052), .ZN(n10064) );
  AOI22_X1 U11106 ( .A1(n10056), .A2(keyinput_f14), .B1(keyinput_f51), .B2(
        n10055), .ZN(n10054) );
  OAI221_X1 U11107 ( .B1(n10056), .B2(keyinput_f14), .C1(n10055), .C2(
        keyinput_f51), .A(n10054), .ZN(n10063) );
  INV_X1 U11108 ( .A(SI_4_), .ZN(n10129) );
  AOI22_X1 U11109 ( .A1(n10058), .A2(keyinput_f18), .B1(keyinput_f28), .B2(
        n10129), .ZN(n10057) );
  OAI221_X1 U11110 ( .B1(n10058), .B2(keyinput_f18), .C1(n10129), .C2(
        keyinput_f28), .A(n10057), .ZN(n10062) );
  XNOR2_X1 U11111 ( .A(P2_REG3_REG_0__SCAN_IN), .B(keyinput_f54), .ZN(n10060)
         );
  XNOR2_X1 U11112 ( .A(SI_25_), .B(keyinput_f7), .ZN(n10059) );
  NAND2_X1 U11113 ( .A1(n10060), .A2(n10059), .ZN(n10061) );
  NOR4_X1 U11114 ( .A1(n10064), .A2(n10063), .A3(n10062), .A4(n10061), .ZN(
        n10090) );
  AOI22_X1 U11115 ( .A1(n6130), .A2(keyinput_f47), .B1(keyinput_f35), .B2(
        n6122), .ZN(n10065) );
  OAI221_X1 U11116 ( .B1(n6130), .B2(keyinput_f47), .C1(n6122), .C2(
        keyinput_f35), .A(n10065), .ZN(n10076) );
  AOI22_X1 U11117 ( .A1(n10103), .A2(keyinput_f10), .B1(keyinput_f46), .B2(
        n10067), .ZN(n10066) );
  OAI221_X1 U11118 ( .B1(n10103), .B2(keyinput_f10), .C1(n10067), .C2(
        keyinput_f46), .A(n10066), .ZN(n10075) );
  AOI22_X1 U11119 ( .A1(n10069), .A2(keyinput_f40), .B1(n4455), .B2(
        keyinput_f61), .ZN(n10068) );
  OAI221_X1 U11120 ( .B1(n10069), .B2(keyinput_f40), .C1(n4455), .C2(
        keyinput_f61), .A(n10068), .ZN(n10074) );
  AOI22_X1 U11121 ( .A1(n10072), .A2(keyinput_f58), .B1(n10071), .B2(
        keyinput_f19), .ZN(n10070) );
  OAI221_X1 U11122 ( .B1(n10072), .B2(keyinput_f58), .C1(n10071), .C2(
        keyinput_f19), .A(n10070), .ZN(n10073) );
  NOR4_X1 U11123 ( .A1(n10076), .A2(n10075), .A3(n10074), .A4(n10073), .ZN(
        n10089) );
  AOI22_X1 U11124 ( .A1(n6128), .A2(keyinput_f50), .B1(n10078), .B2(
        keyinput_f24), .ZN(n10077) );
  OAI221_X1 U11125 ( .B1(n6128), .B2(keyinput_f50), .C1(n10078), .C2(
        keyinput_f24), .A(n10077), .ZN(n10087) );
  AOI22_X1 U11126 ( .A1(n10080), .A2(keyinput_f12), .B1(keyinput_f17), .B2(
        n4892), .ZN(n10079) );
  OAI221_X1 U11127 ( .B1(n10080), .B2(keyinput_f12), .C1(n4892), .C2(
        keyinput_f17), .A(n10079), .ZN(n10086) );
  INV_X1 U11128 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n10126) );
  XOR2_X1 U11129 ( .A(n10126), .B(keyinput_f45), .Z(n10084) );
  XNOR2_X1 U11130 ( .A(SI_0_), .B(keyinput_f32), .ZN(n10083) );
  XNOR2_X1 U11131 ( .A(SI_21_), .B(keyinput_f11), .ZN(n10082) );
  XNOR2_X1 U11132 ( .A(SI_1_), .B(keyinput_f31), .ZN(n10081) );
  NAND4_X1 U11133 ( .A1(n10084), .A2(n10083), .A3(n10082), .A4(n10081), .ZN(
        n10085) );
  NOR3_X1 U11134 ( .A1(n10087), .A2(n10086), .A3(n10085), .ZN(n10088) );
  NAND4_X1 U11135 ( .A1(n10091), .A2(n10090), .A3(n10089), .A4(n10088), .ZN(
        n10092) );
  OAI22_X1 U11136 ( .A1(n10093), .A2(n10092), .B1(keyinput_f63), .B2(
        P2_REG3_REG_15__SCAN_IN), .ZN(n10094) );
  AOI21_X1 U11137 ( .B1(keyinput_f63), .B2(P2_REG3_REG_15__SCAN_IN), .A(n10094), .ZN(n10197) );
  AOI22_X1 U11138 ( .A1(n10097), .A2(keyinput_g9), .B1(keyinput_g25), .B2(
        n10096), .ZN(n10095) );
  OAI221_X1 U11139 ( .B1(n10097), .B2(keyinput_g9), .C1(n10096), .C2(
        keyinput_g25), .A(n10095), .ZN(n10110) );
  AOI22_X1 U11140 ( .A1(n10100), .A2(keyinput_g16), .B1(keyinput_g60), .B2(
        n10099), .ZN(n10098) );
  OAI221_X1 U11141 ( .B1(n10100), .B2(keyinput_g16), .C1(n10099), .C2(
        keyinput_g60), .A(n10098), .ZN(n10109) );
  AOI22_X1 U11142 ( .A1(n10103), .A2(keyinput_g10), .B1(keyinput_g0), .B2(
        n10102), .ZN(n10101) );
  OAI221_X1 U11143 ( .B1(n10103), .B2(keyinput_g10), .C1(n10102), .C2(
        keyinput_g0), .A(n10101), .ZN(n10108) );
  AOI22_X1 U11144 ( .A1(n10106), .A2(keyinput_g29), .B1(keyinput_g44), .B2(
        n10105), .ZN(n10104) );
  OAI221_X1 U11145 ( .B1(n10106), .B2(keyinput_g29), .C1(n10105), .C2(
        keyinput_g44), .A(n10104), .ZN(n10107) );
  NOR4_X1 U11146 ( .A1(n10110), .A2(n10109), .A3(n10108), .A4(n10107), .ZN(
        n10156) );
  AOI22_X1 U11147 ( .A1(n10113), .A2(keyinput_g55), .B1(n10112), .B2(
        keyinput_g4), .ZN(n10111) );
  OAI221_X1 U11148 ( .B1(n10113), .B2(keyinput_g55), .C1(n10112), .C2(
        keyinput_g4), .A(n10111), .ZN(n10124) );
  AOI22_X1 U11149 ( .A1(n10115), .A2(keyinput_g5), .B1(keyinput_g34), .B2(
        P2_U3151), .ZN(n10114) );
  OAI221_X1 U11150 ( .B1(n10115), .B2(keyinput_g5), .C1(P2_U3151), .C2(
        keyinput_g34), .A(n10114), .ZN(n10123) );
  AOI22_X1 U11151 ( .A1(n6128), .A2(keyinput_g50), .B1(keyinput_g2), .B2(
        n10117), .ZN(n10116) );
  OAI221_X1 U11152 ( .B1(n6128), .B2(keyinput_g50), .C1(n10117), .C2(
        keyinput_g2), .A(n10116), .ZN(n10122) );
  INV_X1 U11153 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n10119) );
  AOI22_X1 U11154 ( .A1(n10120), .A2(keyinput_g13), .B1(keyinput_g62), .B2(
        n10119), .ZN(n10118) );
  OAI221_X1 U11155 ( .B1(n10120), .B2(keyinput_g13), .C1(n10119), .C2(
        keyinput_g62), .A(n10118), .ZN(n10121) );
  NOR4_X1 U11156 ( .A1(n10124), .A2(n10123), .A3(n10122), .A4(n10121), .ZN(
        n10155) );
  AOI22_X1 U11157 ( .A1(n10126), .A2(keyinput_g45), .B1(keyinput_g59), .B2(
        n7346), .ZN(n10125) );
  OAI221_X1 U11158 ( .B1(n10126), .B2(keyinput_g45), .C1(n7346), .C2(
        keyinput_g59), .A(n10125), .ZN(n10139) );
  AOI22_X1 U11159 ( .A1(n10129), .A2(keyinput_g28), .B1(keyinput_g52), .B2(
        n10128), .ZN(n10127) );
  OAI221_X1 U11160 ( .B1(n10129), .B2(keyinput_g28), .C1(n10128), .C2(
        keyinput_g52), .A(n10127), .ZN(n10138) );
  AOI22_X1 U11161 ( .A1(n10132), .A2(keyinput_g21), .B1(n10131), .B2(
        keyinput_g6), .ZN(n10130) );
  OAI221_X1 U11162 ( .B1(n10132), .B2(keyinput_g21), .C1(n10131), .C2(
        keyinput_g6), .A(n10130), .ZN(n10137) );
  XOR2_X1 U11163 ( .A(n10133), .B(keyinput_g48), .Z(n10135) );
  XNOR2_X1 U11164 ( .A(SI_2_), .B(keyinput_g30), .ZN(n10134) );
  NAND2_X1 U11165 ( .A1(n10135), .A2(n10134), .ZN(n10136) );
  NOR4_X1 U11166 ( .A1(n10139), .A2(n10138), .A3(n10137), .A4(n10136), .ZN(
        n10154) );
  AOI22_X1 U11167 ( .A1(n10141), .A2(keyinput_g8), .B1(keyinput_g35), .B2(
        n6122), .ZN(n10140) );
  OAI221_X1 U11168 ( .B1(n10141), .B2(keyinput_g8), .C1(n6122), .C2(
        keyinput_g35), .A(n10140), .ZN(n10152) );
  INV_X1 U11169 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n10143) );
  AOI22_X1 U11170 ( .A1(n10144), .A2(keyinput_g23), .B1(keyinput_g42), .B2(
        n10143), .ZN(n10142) );
  OAI221_X1 U11171 ( .B1(n10144), .B2(keyinput_g23), .C1(n10143), .C2(
        keyinput_g42), .A(n10142), .ZN(n10151) );
  AOI22_X1 U11172 ( .A1(n4892), .A2(keyinput_g17), .B1(n10146), .B2(
        keyinput_g7), .ZN(n10145) );
  OAI221_X1 U11173 ( .B1(n4892), .B2(keyinput_g17), .C1(n10146), .C2(
        keyinput_g7), .A(n10145), .ZN(n10150) );
  XNOR2_X1 U11174 ( .A(P2_REG3_REG_6__SCAN_IN), .B(keyinput_g61), .ZN(n10148)
         );
  XNOR2_X1 U11175 ( .A(SI_0_), .B(keyinput_g32), .ZN(n10147) );
  NAND2_X1 U11176 ( .A1(n10148), .A2(n10147), .ZN(n10149) );
  NOR4_X1 U11177 ( .A1(n10152), .A2(n10151), .A3(n10150), .A4(n10149), .ZN(
        n10153) );
  NAND4_X1 U11178 ( .A1(n10156), .A2(n10155), .A3(n10154), .A4(n10153), .ZN(
        n10195) );
  AOI22_X1 U11179 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(keyinput_g56), .B1(
        P2_REG3_REG_25__SCAN_IN), .B2(keyinput_g47), .ZN(n10157) );
  OAI221_X1 U11180 ( .B1(P2_REG3_REG_13__SCAN_IN), .B2(keyinput_g56), .C1(
        P2_REG3_REG_25__SCAN_IN), .C2(keyinput_g47), .A(n10157), .ZN(n10164)
         );
  AOI22_X1 U11181 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(keyinput_g37), .B1(
        SI_21_), .B2(keyinput_g11), .ZN(n10158) );
  OAI221_X1 U11182 ( .B1(P2_REG3_REG_14__SCAN_IN), .B2(keyinput_g37), .C1(
        SI_21_), .C2(keyinput_g11), .A(n10158), .ZN(n10163) );
  AOI22_X1 U11183 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(keyinput_g39), .B1(
        SI_10_), .B2(keyinput_g22), .ZN(n10159) );
  OAI221_X1 U11184 ( .B1(P2_REG3_REG_10__SCAN_IN), .B2(keyinput_g39), .C1(
        SI_10_), .C2(keyinput_g22), .A(n10159), .ZN(n10162) );
  AOI22_X1 U11185 ( .A1(SI_29_), .A2(keyinput_g3), .B1(P2_REG3_REG_11__SCAN_IN), .B2(keyinput_g58), .ZN(n10160) );
  OAI221_X1 U11186 ( .B1(SI_29_), .B2(keyinput_g3), .C1(
        P2_REG3_REG_11__SCAN_IN), .C2(keyinput_g58), .A(n10160), .ZN(n10161)
         );
  NOR4_X1 U11187 ( .A1(n10164), .A2(n10163), .A3(n10162), .A4(n10161), .ZN(
        n10193) );
  XOR2_X1 U11188 ( .A(SI_17_), .B(keyinput_g15), .Z(n10171) );
  AOI22_X1 U11189 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(keyinput_g46), .B1(SI_5_), .B2(keyinput_g27), .ZN(n10165) );
  OAI221_X1 U11190 ( .B1(P2_REG3_REG_12__SCAN_IN), .B2(keyinput_g46), .C1(
        SI_5_), .C2(keyinput_g27), .A(n10165), .ZN(n10170) );
  AOI22_X1 U11191 ( .A1(SI_12_), .A2(keyinput_g20), .B1(SI_18_), .B2(
        keyinput_g14), .ZN(n10166) );
  OAI221_X1 U11192 ( .B1(SI_12_), .B2(keyinput_g20), .C1(SI_18_), .C2(
        keyinput_g14), .A(n10166), .ZN(n10169) );
  AOI22_X1 U11193 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(keyinput_g41), .B1(SI_8_), .B2(keyinput_g24), .ZN(n10167) );
  OAI221_X1 U11194 ( .B1(P2_REG3_REG_19__SCAN_IN), .B2(keyinput_g41), .C1(
        SI_8_), .C2(keyinput_g24), .A(n10167), .ZN(n10168) );
  NOR4_X1 U11195 ( .A1(n10171), .A2(n10170), .A3(n10169), .A4(n10168), .ZN(
        n10192) );
  INV_X1 U11196 ( .A(SI_6_), .ZN(n10173) );
  AOI22_X1 U11197 ( .A1(n5565), .A2(keyinput_g1), .B1(n10173), .B2(
        keyinput_g26), .ZN(n10172) );
  OAI221_X1 U11198 ( .B1(n5565), .B2(keyinput_g1), .C1(n10173), .C2(
        keyinput_g26), .A(n10172), .ZN(n10181) );
  AOI22_X1 U11199 ( .A1(SI_14_), .A2(keyinput_g18), .B1(SI_20_), .B2(
        keyinput_g12), .ZN(n10174) );
  OAI221_X1 U11200 ( .B1(SI_14_), .B2(keyinput_g18), .C1(SI_20_), .C2(
        keyinput_g12), .A(n10174), .ZN(n10180) );
  XNOR2_X1 U11201 ( .A(SI_1_), .B(keyinput_g31), .ZN(n10178) );
  XNOR2_X1 U11202 ( .A(P2_REG3_REG_22__SCAN_IN), .B(keyinput_g57), .ZN(n10177)
         );
  XNOR2_X1 U11203 ( .A(P2_REG3_REG_0__SCAN_IN), .B(keyinput_g54), .ZN(n10176)
         );
  XNOR2_X1 U11204 ( .A(P2_REG3_REG_27__SCAN_IN), .B(keyinput_g36), .ZN(n10175)
         );
  NAND4_X1 U11205 ( .A1(n10178), .A2(n10177), .A3(n10176), .A4(n10175), .ZN(
        n10179) );
  NOR3_X1 U11206 ( .A1(n10181), .A2(n10180), .A3(n10179), .ZN(n10191) );
  AOI22_X1 U11207 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(keyinput_g43), .B1(
        P2_REG3_REG_24__SCAN_IN), .B2(keyinput_g51), .ZN(n10182) );
  OAI221_X1 U11208 ( .B1(P2_REG3_REG_8__SCAN_IN), .B2(keyinput_g43), .C1(
        P2_REG3_REG_24__SCAN_IN), .C2(keyinput_g51), .A(n10182), .ZN(n10189)
         );
  AOI22_X1 U11209 ( .A1(P2_REG3_REG_23__SCAN_IN), .A2(keyinput_g38), .B1(
        SI_13_), .B2(keyinput_g19), .ZN(n10183) );
  OAI221_X1 U11210 ( .B1(P2_REG3_REG_23__SCAN_IN), .B2(keyinput_g38), .C1(
        SI_13_), .C2(keyinput_g19), .A(n10183), .ZN(n10188) );
  AOI22_X1 U11211 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(keyinput_g40), .B1(
        P2_REG3_REG_9__SCAN_IN), .B2(keyinput_g53), .ZN(n10184) );
  OAI221_X1 U11212 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(keyinput_g40), .C1(
        P2_REG3_REG_9__SCAN_IN), .C2(keyinput_g53), .A(n10184), .ZN(n10187) );
  AOI22_X1 U11213 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(keyinput_g49), .B1(
        P2_RD_REG_SCAN_IN), .B2(keyinput_g33), .ZN(n10185) );
  OAI221_X1 U11214 ( .B1(P2_REG3_REG_5__SCAN_IN), .B2(keyinput_g49), .C1(
        P2_RD_REG_SCAN_IN), .C2(keyinput_g33), .A(n10185), .ZN(n10186) );
  NOR4_X1 U11215 ( .A1(n10189), .A2(n10188), .A3(n10187), .A4(n10186), .ZN(
        n10190) );
  NAND4_X1 U11216 ( .A1(n10193), .A2(n10192), .A3(n10191), .A4(n10190), .ZN(
        n10194) );
  OAI22_X1 U11217 ( .A1(keyinput_g63), .A2(n10198), .B1(n10195), .B2(n10194), 
        .ZN(n10196) );
  AOI211_X1 U11218 ( .C1(keyinput_g63), .C2(n10198), .A(n10197), .B(n10196), 
        .ZN(n10199) );
  XOR2_X1 U11219 ( .A(n10200), .B(n10199), .Z(n10201) );
  XNOR2_X1 U11220 ( .A(n10202), .B(n10201), .ZN(ADD_1068_U4) );
  XOR2_X1 U11221 ( .A(n10204), .B(n10203), .Z(ADD_1068_U54) );
  XNOR2_X1 U11222 ( .A(n10206), .B(n10205), .ZN(ADD_1068_U47) );
  XNOR2_X1 U11223 ( .A(n10208), .B(n10207), .ZN(ADD_1068_U48) );
  XNOR2_X1 U11224 ( .A(n10210), .B(n10209), .ZN(ADD_1068_U49) );
  XNOR2_X1 U11225 ( .A(n10212), .B(n10211), .ZN(ADD_1068_U50) );
  XNOR2_X1 U11226 ( .A(n10214), .B(n10213), .ZN(ADD_1068_U51) );
  XOR2_X1 U11227 ( .A(n10216), .B(n10215), .Z(ADD_1068_U53) );
  XNOR2_X1 U11228 ( .A(n10218), .B(n10217), .ZN(ADD_1068_U52) );
  INV_X1 U4887 ( .A(n4555), .ZN(n4810) );
  AND2_X1 U4898 ( .A1(n7449), .A2(n6280), .ZN(n7557) );
  OR2_X1 U4861 ( .A1(n8861), .A2(n7824), .ZN(n5766) );
  CLKBUF_X2 U4874 ( .A(n6135), .Z(n8769) );
  AND2_X1 U4875 ( .A1(n6767), .A2(n5740), .ZN(n10222) );
endmodule

