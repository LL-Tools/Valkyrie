

module b14_C_2inp_gates_syn ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, U3352, U3351, U3350, U3349, 
        U3348, U3347, U3346, U3345, U3344, U3343, U3342, U3341, U3340, U3339, 
        U3338, U3337, U3336, U3335, U3334, U3333, U3332, U3331, U3330, U3329, 
        U3328, U3327, U3326, U3325, U3324, U3323, U3322, U3321, U3458, U3459, 
        U3320, U3319, U3318, U3317, U3316, U3315, U3314, U3313, U3312, U3311, 
        U3310, U3309, U3308, U3307, U3306, U3305, U3304, U3303, U3302, U3301, 
        U3300, U3299, U3298, U3297, U3296, U3295, U3294, U3293, U3292, U3291, 
        U3467, U3469, U3471, U3473, U3475, U3477, U3479, U3481, U3483, U3485, 
        U3487, U3489, U3491, U3493, U3495, U3497, U3499, U3501, U3503, U3505, 
        U3506, U3507, U3508, U3509, U3510, U3511, U3512, U3513, U3514, U3515, 
        U3516, U3517, U3518, U3519, U3520, U3521, U3522, U3523, U3524, U3525, 
        U3526, U3527, U3528, U3529, U3530, U3531, U3532, U3533, U3534, U3535, 
        U3536, U3537, U3538, U3539, U3540, U3541, U3542, U3543, U3544, U3545, 
        U3546, U3547, U3548, U3549, U3290, U3289, U3288, U3287, U3286, U3285, 
        U3284, U3283, U3282, U3281, U3280, U3279, U3278, U3277, U3276, U3275, 
        U3274, U3273, U3272, U3271, U3270, U3269, U3268, U3267, U3266, U3265, 
        U3264, U3263, U3262, U3354, U3261, U3260, U3259, U3258, U3257, U3256, 
        U3255, U3254, U3253, U3252, U3251, U3250, U3249, U3248, U3247, U3246, 
        U3245, U3244, U3243, U3242, U3241, U3240, U3550, U3551, U3552, U3553, 
        U3554, U3555, U3556, U3557, U3558, U3559, U3560, U3561, U3562, U3563, 
        U3564, U3565, U3566, U3567, U3568, U3569, U3570, U3571, U3572, U3573, 
        U3574, U3575, U3576, U3577, U3578, U3579, U3580, U3581, U3239, U3238, 
        U3237, U3236, U3235, U3234, U3233, U3232, U3231, U3230, U3229, U3228, 
        U3227, U3226, U3225, U3224, U3223, U3222, U3221, U3220, U3219, U3218, 
        U3217, U3216, U3215, U3214, U3213, U3212, U3211, U3210, U3149, U3148, 
        U4043, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, 
        keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, 
        keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, 
        keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, 
        keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, 
        keyinput29, keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, 
        keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, 
        keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, 
        keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, 
        keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, 
        keyinput59, keyinput60, keyinput61, keyinput62, keyinput63 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016,
         n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026,
         n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036,
         n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046,
         n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056,
         n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066,
         n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076,
         n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086,
         n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096,
         n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106,
         n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116,
         n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126,
         n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136,
         n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146,
         n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156,
         n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166,
         n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176,
         n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186,
         n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196,
         n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206,
         n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216,
         n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226,
         n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236,
         n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246,
         n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256,
         n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266,
         n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276,
         n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286,
         n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296,
         n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306,
         n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316,
         n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326,
         n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336,
         n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346,
         n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356,
         n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366,
         n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376,
         n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386,
         n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396,
         n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406,
         n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416,
         n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426,
         n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436,
         n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446,
         n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456,
         n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466,
         n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476,
         n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486,
         n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496,
         n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506,
         n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516,
         n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526,
         n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536,
         n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546,
         n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556,
         n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566,
         n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576,
         n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586,
         n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596,
         n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606,
         n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616,
         n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626,
         n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636,
         n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646,
         n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656,
         n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666,
         n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676,
         n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686,
         n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696,
         n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706,
         n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716,
         n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726,
         n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736,
         n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746,
         n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756,
         n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766,
         n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776,
         n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786,
         n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796,
         n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806,
         n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816,
         n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826,
         n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836,
         n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846,
         n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856,
         n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866,
         n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876,
         n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886,
         n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896,
         n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906,
         n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916,
         n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926,
         n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936,
         n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946,
         n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956,
         n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966,
         n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976,
         n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986,
         n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996,
         n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006,
         n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016,
         n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026,
         n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036,
         n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046,
         n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056,
         n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066,
         n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076,
         n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086,
         n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096,
         n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106,
         n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116,
         n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126,
         n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136,
         n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146,
         n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156,
         n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166,
         n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176,
         n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186,
         n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196,
         n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206,
         n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216,
         n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226,
         n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236,
         n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246,
         n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256,
         n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266,
         n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276,
         n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286,
         n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296,
         n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306,
         n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316,
         n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326,
         n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336,
         n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346,
         n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356,
         n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366,
         n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376,
         n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386,
         n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396,
         n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406,
         n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416,
         n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426,
         n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436,
         n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446,
         n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456,
         n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466,
         n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476,
         n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486,
         n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496,
         n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506,
         n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516,
         n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526,
         n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536,
         n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546,
         n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556,
         n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566,
         n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576,
         n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586,
         n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596,
         n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606,
         n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616,
         n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626,
         n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636,
         n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646,
         n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656,
         n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666,
         n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676,
         n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686,
         n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696,
         n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706,
         n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716,
         n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726,
         n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736,
         n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746,
         n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756,
         n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766,
         n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776,
         n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786,
         n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796,
         n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806,
         n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816,
         n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826,
         n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836,
         n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846,
         n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856,
         n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866,
         n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876,
         n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886,
         n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896,
         n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906,
         n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916,
         n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926,
         n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936,
         n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946,
         n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956,
         n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966,
         n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976,
         n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986,
         n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996,
         n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006,
         n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016,
         n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026,
         n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036,
         n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046,
         n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056,
         n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066,
         n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076,
         n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086,
         n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096,
         n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106,
         n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116,
         n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126,
         n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136,
         n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146,
         n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156,
         n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166,
         n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176,
         n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186,
         n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196,
         n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206,
         n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216,
         n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226,
         n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236,
         n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246,
         n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256,
         n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266,
         n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276,
         n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286,
         n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296,
         n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306,
         n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316,
         n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326,
         n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336,
         n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346,
         n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356,
         n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366,
         n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376,
         n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386,
         n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396,
         n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406,
         n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416,
         n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426,
         n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436,
         n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446,
         n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456,
         n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466,
         n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476,
         n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486,
         n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496,
         n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506,
         n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516,
         n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526,
         n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536,
         n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546,
         n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556,
         n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566,
         n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576,
         n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586,
         n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596,
         n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606,
         n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616,
         n4617, n4618, n4619, n4620, n4621, n4623, n4624, n4625, n4626, n4627,
         n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637,
         n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647,
         n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657,
         n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667,
         n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677,
         n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687,
         n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697,
         n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707,
         n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717,
         n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727,
         n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737,
         n4738, n4739, n4740, n4741;

  NAND2_X1 U2249 ( .A1(n2153), .A2(n2157), .ZN(n3672) );
  INV_X2 U2250 ( .A(n2741), .ZN(n3556) );
  NAND2_X1 U2251 ( .A1(n3027), .A2(n3223), .ZN(n3787) );
  NAND2_X1 U2252 ( .A1(n2620), .A2(n3803), .ZN(n3385) );
  INV_X1 U2253 ( .A(n2754), .ZN(n3557) );
  NAND2_X1 U2254 ( .A1(n3270), .A2(n3269), .ZN(n3341) );
  OAI21_X1 U2255 ( .B1(n3385), .B2(n3383), .A(n3806), .ZN(n3395) );
  INV_X1 U2256 ( .A(n2344), .ZN(n3722) );
  INV_X1 U2257 ( .A(n2720), .ZN(n3027) );
  NAND2_X1 U2258 ( .A1(n2012), .A2(n2608), .ZN(n3766) );
  INV_X1 U2259 ( .A(n2315), .ZN(n2745) );
  XNOR2_X1 U2260 ( .A(n2093), .B(n2092), .ZN(n2940) );
  BUF_X1 U2261 ( .A(n2940), .Z(n2007) );
  AOI21_X2 U2262 ( .B1(n3037), .B2(REG2_REG_6__SCAN_IN), .A(n3036), .ZN(n3039)
         );
  AND3_X1 U2263 ( .A1(n2317), .A2(n2235), .A3(n2236), .ZN(n2376) );
  AOI21_X2 U2264 ( .B1(n3296), .B2(n2395), .A(n2394), .ZN(n3384) );
  OAI21_X2 U2265 ( .B1(n4167), .B2(n4442), .A(n4166), .ZN(n4475) );
  NOR2_X2 U2266 ( .A1(n2495), .A2(IR_REG_18__SCAN_IN), .ZN(n2606) );
  OAI22_X2 U2267 ( .A1(n3114), .A2(n2356), .B1(n2355), .B2(n2354), .ZN(n3283)
         );
  NAND2_X2 U2268 ( .A1(n4059), .A2(n4058), .ZN(n4636) );
  NAND2_X1 U2269 ( .A1(n4647), .A2(n4648), .ZN(n4646) );
  OAI21_X1 U2270 ( .B1(n4075), .B2(REG1_REG_16__SCAN_IN), .A(n2101), .ZN(n4647) );
  CLKBUF_X1 U2271 ( .A(n2720), .Z(n3082) );
  INV_X2 U2272 ( .A(n3561), .ZN(n3533) );
  INV_X1 U2273 ( .A(n4016), .ZN(n3168) );
  AND4_X2 U2274 ( .A1(n2313), .A2(n2312), .A3(n2311), .A4(n2310), .ZN(n2315)
         );
  NAND4_X1 U2275 ( .A1(n2325), .A2(n2324), .A3(n2323), .A4(n2322), .ZN(n4016)
         );
  NAND2_X2 U2276 ( .A1(n2611), .A2(n2644), .ZN(n3131) );
  XNOR2_X1 U2277 ( .A(n2928), .B(n2319), .ZN(n2991) );
  INV_X2 U2278 ( .A(n2447), .ZN(n2329) );
  AOI21_X1 U2279 ( .B1(n2023), .B2(n4665), .A(n4664), .ZN(n4672) );
  MUX2_X1 U2280 ( .A(n4481), .B(n4556), .S(n4741), .Z(n4482) );
  MUX2_X1 U2281 ( .A(n4557), .B(n4556), .S(n4731), .Z(n4558) );
  AOI21_X1 U2282 ( .B1(n4659), .B2(n4658), .A(n4657), .ZN(n4665) );
  AOI21_X1 U2283 ( .B1(n4124), .B2(n4393), .A(n4123), .ZN(n4469) );
  OAI21_X1 U2284 ( .B1(n2228), .B2(n3482), .A(n3485), .ZN(n4495) );
  AND3_X1 U2285 ( .A1(n4468), .A2(n4467), .A3(n4466), .ZN(n4470) );
  AND2_X1 U2286 ( .A1(n3484), .A2(n3481), .ZN(n2228) );
  OAI21_X1 U2287 ( .B1(n4079), .B2(n2136), .A(n2134), .ZN(n4667) );
  AND2_X1 U2288 ( .A1(n4181), .A2(n4180), .ZN(n4206) );
  NOR2_X1 U2289 ( .A1(n4051), .A2(n2044), .ZN(n4056) );
  AND2_X1 U2290 ( .A1(n3466), .A2(n3467), .ZN(n4051) );
  AOI21_X1 U2291 ( .B1(n4465), .B2(n4721), .A(n4464), .ZN(n4466) );
  NAND2_X1 U2292 ( .A1(n2187), .A2(n2032), .ZN(n4375) );
  AND2_X1 U2293 ( .A1(n3051), .A2(n2740), .ZN(n3094) );
  XNOR2_X1 U2294 ( .A(n3030), .B(n4619), .ZN(n3032) );
  NAND2_X2 U2295 ( .A1(n3129), .A2(n4360), .ZN(n4682) );
  AOI21_X1 U2296 ( .B1(n2999), .B2(REG1_REG_4__SCAN_IN), .A(n2998), .ZN(n3017)
         );
  AND2_X1 U2297 ( .A1(n3796), .A2(n3794), .ZN(n3755) );
  XNOR2_X1 U2298 ( .A(n2997), .B(n2947), .ZN(n2999) );
  BUF_X4 U2299 ( .A(n2741), .Z(n3560) );
  INV_X1 U2300 ( .A(n3502), .ZN(n2985) );
  NAND4_X2 U2301 ( .A1(n2375), .A2(n2374), .A3(n2373), .A4(n2372), .ZN(n4015)
         );
  OAI21_X2 U2302 ( .B1(n2378), .B2(n2933), .A(n2294), .ZN(n3223) );
  NAND2_X2 U2303 ( .A1(n2892), .A2(n3131), .ZN(n3561) );
  AND4_X1 U2304 ( .A1(n2335), .A2(n2334), .A3(n2333), .A4(n2332), .ZN(n3502)
         );
  BUF_X4 U2305 ( .A(n2330), .Z(n2009) );
  NAND2_X2 U2306 ( .A1(n2257), .A2(n2256), .ZN(n2378) );
  AND2_X2 U2307 ( .A1(n4608), .A2(n2965), .ZN(n2331) );
  NAND2_X1 U2308 ( .A1(n2679), .A2(IR_REG_31__SCAN_IN), .ZN(n2670) );
  INV_X1 U2309 ( .A(n2274), .ZN(n2965) );
  INV_X4 U2310 ( .A(n2301), .ZN(n2008) );
  NAND2_X1 U2311 ( .A1(n2510), .A2(n2509), .ZN(n2602) );
  NAND2_X1 U2312 ( .A1(n2272), .A2(n3580), .ZN(n2274) );
  MUX2_X1 U2313 ( .A(IR_REG_31__SCAN_IN), .B(n2270), .S(IR_REG_29__SCAN_IN), 
        .Z(n2272) );
  OR2_X1 U2314 ( .A1(n2271), .A2(n2267), .ZN(n2268) );
  NOR2_X1 U2315 ( .A1(n2269), .A2(IR_REG_29__SCAN_IN), .ZN(n2271) );
  INV_X1 U2316 ( .A(IR_REG_8__SCAN_IN), .ZN(n2385) );
  INV_X1 U2317 ( .A(IR_REG_7__SCAN_IN), .ZN(n2358) );
  NOR2_X1 U2318 ( .A1(IR_REG_11__SCAN_IN), .A2(IR_REG_16__SCAN_IN), .ZN(n2242)
         );
  NOR2_X1 U2319 ( .A1(IR_REG_13__SCAN_IN), .A2(IR_REG_10__SCAN_IN), .ZN(n2243)
         );
  NOR2_X1 U2320 ( .A1(IR_REG_15__SCAN_IN), .A2(IR_REG_14__SCAN_IN), .ZN(n2244)
         );
  NOR2_X2 U2321 ( .A1(IR_REG_0__SCAN_IN), .A2(IR_REG_1__SCAN_IN), .ZN(n2317)
         );
  INV_X1 U2322 ( .A(IR_REG_19__SCAN_IN), .ZN(n2509) );
  AOI21_X1 U2323 ( .B1(n3337), .B2(REG2_REG_10__SCAN_IN), .A(n3336), .ZN(n3340) );
  NAND2_X1 U2324 ( .A1(n2273), .A2(n2274), .ZN(n2301) );
  INV_X1 U2325 ( .A(n2024), .ZN(n2082) );
  NAND2_X1 U2326 ( .A1(n2163), .A2(n2837), .ZN(n2162) );
  INV_X1 U2327 ( .A(n2840), .ZN(n2163) );
  INV_X1 U2328 ( .A(n2582), .ZN(n2201) );
  NAND2_X1 U2329 ( .A1(n2266), .A2(n2265), .ZN(n2659) );
  OR2_X1 U2330 ( .A1(n2028), .A2(n2082), .ZN(n2079) );
  NOR2_X1 U2331 ( .A1(n3831), .A2(n2090), .ZN(n2089) );
  OR2_X1 U2332 ( .A1(n2191), .A2(n2190), .ZN(n2189) );
  NAND2_X1 U2333 ( .A1(n4387), .A2(n4424), .ZN(n2197) );
  NAND2_X1 U2334 ( .A1(n2985), .A2(n3120), .ZN(n3796) );
  NAND2_X1 U2335 ( .A1(n4329), .A2(n2485), .ZN(n2205) );
  NAND2_X1 U2336 ( .A1(n2484), .A2(n2483), .ZN(n2485) );
  OR2_X1 U2337 ( .A1(n2975), .A2(n2692), .ZN(n2877) );
  INV_X1 U2338 ( .A(IR_REG_27__SCAN_IN), .ZN(n2264) );
  INV_X1 U2339 ( .A(IR_REG_22__SCAN_IN), .ZN(n2666) );
  OAI21_X1 U2340 ( .B1(n3653), .B2(n2181), .A(n2180), .ZN(n3660) );
  NAND2_X1 U2341 ( .A1(n2185), .A2(n2182), .ZN(n2181) );
  NAND2_X1 U2342 ( .A1(n2185), .A2(n2183), .ZN(n2180) );
  INV_X1 U2343 ( .A(n3508), .ZN(n2185) );
  INV_X1 U2344 ( .A(n2158), .ZN(n2157) );
  OAI21_X1 U2345 ( .B1(n2160), .B2(n3632), .A(n3633), .ZN(n2158) );
  INV_X1 U2346 ( .A(n4172), .ZN(n3686) );
  INV_X1 U2347 ( .A(n2894), .ZN(n2900) );
  AND2_X1 U2348 ( .A1(n3560), .A2(n2893), .ZN(n2896) );
  INV_X1 U2349 ( .A(n2331), .ZN(n2646) );
  NOR2_X1 U2350 ( .A1(n2676), .A2(n2976), .ZN(n2678) );
  NOR2_X1 U2351 ( .A1(n3015), .A2(n3000), .ZN(n3030) );
  NOR2_X1 U2352 ( .A1(n3019), .A2(n4737), .ZN(n3000) );
  NAND2_X1 U2353 ( .A1(n4057), .A2(n4614), .ZN(n4058) );
  INV_X1 U2354 ( .A(n4056), .ZN(n4057) );
  INV_X1 U2355 ( .A(n4093), .ZN(n4119) );
  AND2_X1 U2356 ( .A1(n4156), .A2(n2580), .ZN(n2581) );
  OR2_X1 U2357 ( .A1(n2553), .A2(n3645), .ZN(n2555) );
  AND2_X1 U2358 ( .A1(n2645), .A2(n3863), .ZN(n4442) );
  AND2_X1 U2359 ( .A1(n4609), .A2(n2917), .ZN(n4386) );
  OR2_X1 U2360 ( .A1(n3026), .A2(n2611), .ZN(n4391) );
  NAND2_X1 U2361 ( .A1(n2591), .A2(n2590), .ZN(n4165) );
  NAND2_X1 U2362 ( .A1(n3087), .A2(n2745), .ZN(n3791) );
  NOR2_X1 U2363 ( .A1(n4116), .A2(n2080), .ZN(n2076) );
  INV_X1 U2364 ( .A(n2149), .ZN(n2148) );
  AND2_X1 U2365 ( .A1(n2162), .A2(n2161), .ZN(n2159) );
  NOR2_X1 U2366 ( .A1(n2440), .A2(n2439), .ZN(n2260) );
  OR2_X1 U2367 ( .A1(n2723), .A2(n4611), .ZN(n2892) );
  OR2_X1 U2368 ( .A1(n3268), .A2(n3952), .ZN(n3269) );
  NOR2_X1 U2369 ( .A1(n2082), .A2(n2081), .ZN(n2080) );
  INV_X1 U2370 ( .A(n3851), .ZN(n2081) );
  NOR2_X1 U2371 ( .A1(n3738), .A2(n2084), .ZN(n2083) );
  NAND2_X1 U2372 ( .A1(n4346), .A2(n3748), .ZN(n2091) );
  NOR2_X1 U2373 ( .A1(n2190), .A2(n2194), .ZN(n2188) );
  AOI21_X1 U2374 ( .B1(n2210), .B2(n2222), .A(n2030), .ZN(n2209) );
  NOR2_X1 U2375 ( .A1(n2227), .A2(n2410), .ZN(n2210) );
  INV_X1 U2376 ( .A(n2227), .ZN(n2211) );
  NOR2_X1 U2377 ( .A1(n4323), .A2(n2204), .ZN(n2203) );
  INV_X1 U2378 ( .A(n2486), .ZN(n2204) );
  INV_X1 U2379 ( .A(IR_REG_25__SCAN_IN), .ZN(n2265) );
  INV_X1 U2380 ( .A(IR_REG_17__SCAN_IN), .ZN(n2246) );
  INV_X1 U2381 ( .A(IR_REG_24__SCAN_IN), .ZN(n2249) );
  OR3_X1 U2382 ( .A1(n2411), .A2(IR_REG_12__SCAN_IN), .A3(IR_REG_11__SCAN_IN), 
        .ZN(n2435) );
  NAND2_X1 U2383 ( .A1(n3135), .A2(n3136), .ZN(n2149) );
  NAND2_X1 U2384 ( .A1(n2152), .A2(n2151), .ZN(n2150) );
  INV_X1 U2385 ( .A(n3136), .ZN(n2151) );
  INV_X1 U2386 ( .A(n3135), .ZN(n2152) );
  NOR2_X1 U2387 ( .A1(n2171), .A2(n2167), .ZN(n2166) );
  XNOR2_X1 U2388 ( .A(n2753), .B(n3533), .ZN(n2759) );
  OR2_X1 U2389 ( .A1(n2148), .A2(n2150), .ZN(n2146) );
  AND2_X1 U2390 ( .A1(n2148), .A2(n3212), .ZN(n2144) );
  AND2_X1 U2391 ( .A1(n2731), .A2(n2730), .ZN(n2735) );
  NAND2_X1 U2392 ( .A1(n2162), .A2(n2841), .ZN(n2160) );
  OR2_X1 U2393 ( .A1(n2397), .A2(n2396), .ZN(n2399) );
  NAND2_X1 U2394 ( .A1(n2908), .A2(n2263), .ZN(n2257) );
  NAND2_X1 U2395 ( .A1(n3598), .A2(n3515), .ZN(n3597) );
  AND2_X1 U2396 ( .A1(n3543), .A2(n3542), .ZN(n3544) );
  NAND2_X1 U2397 ( .A1(n2926), .A2(n2925), .ZN(n4037) );
  NOR2_X1 U2398 ( .A1(n3002), .A2(n3005), .ZN(n2129) );
  NOR2_X1 U2399 ( .A1(n3060), .A2(n3059), .ZN(n3145) );
  AND2_X1 U2400 ( .A1(n4618), .A2(REG2_REG_7__SCAN_IN), .ZN(n3059) );
  NAND2_X1 U2401 ( .A1(n2104), .A2(n2103), .ZN(n3154) );
  NAND2_X1 U2402 ( .A1(n2105), .A2(n2022), .ZN(n2104) );
  NAND2_X1 U2403 ( .A1(n2107), .A2(n3065), .ZN(n2105) );
  INV_X1 U2404 ( .A(n3152), .ZN(n3149) );
  NAND2_X1 U2405 ( .A1(n3266), .A2(n3265), .ZN(n3335) );
  OR2_X1 U2406 ( .A1(n3268), .A2(n3264), .ZN(n3265) );
  XNOR2_X1 U2407 ( .A(n3335), .B(n3334), .ZN(n3337) );
  NOR2_X1 U2408 ( .A1(n3344), .A2(n2115), .ZN(n2114) );
  XNOR2_X1 U2409 ( .A(n3341), .B(n3334), .ZN(n3271) );
  NOR2_X1 U2410 ( .A1(n3434), .A2(n3433), .ZN(n3464) );
  AND2_X1 U2411 ( .A1(n4616), .A2(REG1_REG_11__SCAN_IN), .ZN(n3433) );
  NOR2_X1 U2412 ( .A1(n2121), .A2(n3456), .ZN(n2120) );
  INV_X1 U2413 ( .A(n2123), .ZN(n2121) );
  NAND2_X1 U2414 ( .A1(n2118), .A2(n2045), .ZN(n2122) );
  OAI22_X1 U2415 ( .A1(n4046), .A2(n4045), .B1(REG2_REG_13__SCAN_IN), .B2(
        n4615), .ZN(n4063) );
  AND2_X1 U2416 ( .A1(n4635), .A2(n4612), .ZN(n2096) );
  INV_X1 U2417 ( .A(n4635), .ZN(n2098) );
  NOR2_X1 U2418 ( .A1(n4060), .A2(n4612), .ZN(n2100) );
  AND2_X1 U2419 ( .A1(n4612), .A2(REG2_REG_16__SCAN_IN), .ZN(n2141) );
  AND2_X1 U2420 ( .A1(n2918), .A2(n3722), .ZN(n2919) );
  OR2_X1 U2421 ( .A1(n4612), .A2(REG2_REG_16__SCAN_IN), .ZN(n2142) );
  NAND2_X1 U2422 ( .A1(n4631), .A2(n2052), .ZN(n4079) );
  NOR2_X1 U2423 ( .A1(n2141), .A2(n2139), .ZN(n2138) );
  INV_X1 U2424 ( .A(n4651), .ZN(n2139) );
  NAND2_X1 U2425 ( .A1(n2920), .A2(n2919), .ZN(n4626) );
  NAND2_X1 U2426 ( .A1(n4634), .A2(n2095), .ZN(n2101) );
  NOR2_X1 U2427 ( .A1(n4060), .A2(n4612), .ZN(n2095) );
  INV_X1 U2428 ( .A(n2216), .ZN(n2213) );
  OR2_X1 U2429 ( .A1(n2584), .A2(n2583), .ZN(n2595) );
  NOR2_X1 U2430 ( .A1(n2581), .A2(n2021), .ZN(n2199) );
  OR2_X1 U2431 ( .A1(n2555), .A2(n3967), .ZN(n2573) );
  AOI21_X1 U2432 ( .B1(n2060), .B2(n2562), .A(n2031), .ZN(n4156) );
  NAND2_X1 U2433 ( .A1(n4182), .A2(n4180), .ZN(n2060) );
  INV_X1 U2434 ( .A(REG3_REG_24__SCAN_IN), .ZN(n3645) );
  NAND2_X1 U2435 ( .A1(n2513), .A2(n2016), .ZN(n2539) );
  NAND2_X1 U2436 ( .A1(n3482), .A2(n3481), .ZN(n2059) );
  INV_X1 U2437 ( .A(n2089), .ZN(n2088) );
  AND2_X1 U2438 ( .A1(n3714), .A2(n2087), .ZN(n2086) );
  INV_X1 U2439 ( .A(n3663), .ZN(n4273) );
  AND3_X1 U2440 ( .A1(n2277), .A2(n2276), .A3(n2275), .ZN(n4414) );
  NAND2_X1 U2441 ( .A1(n2034), .A2(n2197), .ZN(n2191) );
  NAND2_X1 U2442 ( .A1(n2409), .A2(n3389), .ZN(n2410) );
  AND2_X1 U2443 ( .A1(n3298), .A2(n3319), .ZN(n2394) );
  AOI21_X1 U2444 ( .B1(n2064), .B2(n2067), .A(n2063), .ZN(n2062) );
  INV_X1 U2445 ( .A(n3804), .ZN(n2063) );
  INV_X1 U2446 ( .A(n4611), .ZN(n4088) );
  AND4_X1 U2447 ( .A1(n2352), .A2(n2351), .A3(n2350), .A4(n2349), .ZN(n3277)
         );
  NAND2_X1 U2448 ( .A1(n2216), .A2(n2215), .ZN(n2214) );
  NOR2_X1 U2449 ( .A1(n3686), .A2(n4119), .ZN(n2215) );
  OR2_X1 U2450 ( .A1(n4196), .A2(n3527), .ZN(n4197) );
  INV_X1 U2451 ( .A(n3268), .ZN(n2408) );
  NAND2_X1 U2452 ( .A1(n3722), .A2(n2406), .ZN(n2407) );
  INV_X1 U2453 ( .A(n2742), .ZN(n3087) );
  NOR2_X1 U2454 ( .A1(n3223), .A2(n3221), .ZN(n3220) );
  NAND2_X1 U2455 ( .A1(n2675), .A2(n2979), .ZN(n2975) );
  INV_X1 U2456 ( .A(n4690), .ZN(n2681) );
  INV_X1 U2457 ( .A(n2674), .ZN(n2254) );
  AOI21_X1 U2458 ( .B1(n2669), .B2(n2668), .A(n2667), .ZN(n2679) );
  NOR2_X1 U2459 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_23__SCAN_IN), .ZN(n2667)
         );
  AND3_X1 U2460 ( .A1(n2666), .A2(n2665), .A3(n2664), .ZN(n2668) );
  INV_X1 U2461 ( .A(IR_REG_20__SCAN_IN), .ZN(n2603) );
  NAND2_X1 U2462 ( .A1(n2602), .A2(IR_REG_31__SCAN_IN), .ZN(n2604) );
  NAND2_X1 U2463 ( .A1(n2507), .A2(IR_REG_31__SCAN_IN), .ZN(n2510) );
  OR2_X1 U2464 ( .A1(n2357), .A2(n2237), .ZN(n2481) );
  NAND2_X1 U2465 ( .A1(n2289), .A2(IR_REG_31__SCAN_IN), .ZN(n2290) );
  AND2_X1 U2466 ( .A1(n2579), .A2(n2578), .ZN(n4142) );
  OR2_X1 U2467 ( .A1(n4169), .A2(n2646), .ZN(n2579) );
  NOR2_X1 U2468 ( .A1(n3654), .A2(n2884), .ZN(n3510) );
  AND2_X1 U2469 ( .A1(n2560), .A2(n2559), .ZN(n4191) );
  AND2_X1 U2470 ( .A1(n2494), .A2(n2493), .ZN(n4295) );
  AND2_X1 U2471 ( .A1(n2900), .A2(n2898), .ZN(n3691) );
  NOR2_X1 U2472 ( .A1(n3017), .A2(n3016), .ZN(n3015) );
  NOR2_X1 U2473 ( .A1(n3340), .A2(n3339), .ZN(n3428) );
  NAND2_X1 U2474 ( .A1(n4633), .A2(n4632), .ZN(n4631) );
  OAI21_X1 U2475 ( .B1(n2054), .B2(n2011), .A(n2111), .ZN(n2110) );
  NAND2_X1 U2476 ( .A1(n2018), .A2(n2053), .ZN(n2111) );
  OR2_X1 U2477 ( .A1(n4626), .A2(n4624), .ZN(n4657) );
  INV_X1 U2478 ( .A(n3470), .ZN(n4670) );
  OAI21_X1 U2479 ( .B1(n2658), .B2(n4442), .A(n2229), .ZN(n4136) );
  XNOR2_X1 U2480 ( .A(n4109), .B(n3783), .ZN(n4130) );
  AND2_X1 U2481 ( .A1(n2611), .A2(n4611), .ZN(n4674) );
  AOI21_X1 U2482 ( .B1(n4130), .B2(n4724), .A(n4136), .ZN(n2718) );
  INV_X1 U2483 ( .A(n3589), .ZN(n2161) );
  NAND2_X1 U2484 ( .A1(n2642), .A2(n3716), .ZN(n2085) );
  INV_X1 U2485 ( .A(IR_REG_6__SCAN_IN), .ZN(n2247) );
  NOR2_X1 U2486 ( .A1(n3358), .A2(n2172), .ZN(n2171) );
  INV_X1 U2487 ( .A(n2177), .ZN(n2167) );
  NOR2_X1 U2488 ( .A1(n2173), .A2(n2171), .ZN(n2165) );
  NOR2_X1 U2489 ( .A1(n3359), .A2(n2174), .ZN(n2173) );
  NAND2_X1 U2490 ( .A1(n2175), .A2(n3440), .ZN(n2174) );
  NAND2_X1 U2491 ( .A1(n2179), .A2(n2178), .ZN(n2177) );
  INV_X1 U2492 ( .A(n3306), .ZN(n2179) );
  INV_X1 U2493 ( .A(n3307), .ZN(n2178) );
  NAND2_X1 U2494 ( .A1(n3509), .A2(n2184), .ZN(n2183) );
  NOR2_X1 U2495 ( .A1(n2417), .A2(n2416), .ZN(n2415) );
  AND2_X1 U2496 ( .A1(n2159), .A2(n2155), .ZN(n2154) );
  NAND2_X1 U2497 ( .A1(n3003), .A2(REG2_REG_4__SCAN_IN), .ZN(n2133) );
  NAND2_X1 U2498 ( .A1(n2059), .A2(n2564), .ZN(n2565) );
  NOR2_X1 U2499 ( .A1(n3978), .A2(n2058), .ZN(n2057) );
  NAND2_X1 U2500 ( .A1(n2089), .A2(n4353), .ZN(n2087) );
  NOR2_X1 U2501 ( .A1(n2487), .A2(n3675), .ZN(n2499) );
  AND2_X1 U2502 ( .A1(n2260), .A2(n2048), .ZN(n2471) );
  AND2_X1 U2503 ( .A1(n3800), .A2(n2379), .ZN(n2380) );
  OR2_X1 U2504 ( .A1(n4015), .A2(n3282), .ZN(n2379) );
  NAND2_X1 U2505 ( .A1(n2699), .A2(n2367), .ZN(n3804) );
  AOI21_X1 U2506 ( .B1(n2071), .B2(n2069), .A(n2068), .ZN(n2067) );
  CLKBUF_X1 U2507 ( .A(n3071), .Z(n3072) );
  NOR2_X1 U2508 ( .A1(n3845), .A2(n4110), .ZN(n2216) );
  AOI21_X1 U2509 ( .B1(n2079), .B2(n2076), .A(n2075), .ZN(n2074) );
  NAND2_X1 U2510 ( .A1(n2079), .A2(n4114), .ZN(n2077) );
  INV_X1 U2511 ( .A(n4115), .ZN(n2075) );
  AND2_X1 U2512 ( .A1(n3722), .A2(DATAI_20_), .ZN(n4270) );
  NAND2_X1 U2513 ( .A1(n4347), .A2(n4336), .ZN(n2486) );
  OR2_X1 U2514 ( .A1(n2218), .A2(n4336), .ZN(n2217) );
  NAND2_X1 U2515 ( .A1(n4376), .A2(n4399), .ZN(n2220) );
  NOR2_X1 U2516 ( .A1(n3398), .A2(n3389), .ZN(n2212) );
  NOR2_X1 U2517 ( .A1(n3246), .A2(n2701), .ZN(n3195) );
  INV_X1 U2518 ( .A(n3196), .ZN(n2700) );
  INV_X1 U2519 ( .A(IR_REG_28__SCAN_IN), .ZN(n2263) );
  AND2_X1 U2520 ( .A1(n2652), .A2(n2253), .ZN(n2908) );
  AND2_X1 U2521 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_27__SCAN_IN), .ZN(n2255)
         );
  INV_X1 U2522 ( .A(IR_REG_23__SCAN_IN), .ZN(n2664) );
  INV_X1 U2523 ( .A(IR_REG_21__SCAN_IN), .ZN(n2665) );
  INV_X1 U2524 ( .A(IR_REG_14__SCAN_IN), .ZN(n3884) );
  INV_X1 U2525 ( .A(IR_REG_1__SCAN_IN), .ZN(n2289) );
  NAND2_X1 U2526 ( .A1(n2260), .A2(REG3_REG_14__SCAN_IN), .ZN(n2448) );
  NAND2_X1 U2527 ( .A1(n2795), .A2(n2794), .ZN(n3374) );
  INV_X1 U2528 ( .A(REG3_REG_8__SCAN_IN), .ZN(n2387) );
  AND2_X1 U2529 ( .A1(n3722), .A2(DATAI_25_), .ZN(n3527) );
  NAND2_X1 U2530 ( .A1(n2260), .A2(n2015), .ZN(n2458) );
  INV_X1 U2531 ( .A(n2726), .ZN(n3554) );
  OR2_X1 U2532 ( .A1(n2388), .A2(n2387), .ZN(n2397) );
  INV_X1 U2533 ( .A(REG3_REG_9__SCAN_IN), .ZN(n2396) );
  NAND2_X1 U2534 ( .A1(n3306), .A2(n3307), .ZN(n2175) );
  INV_X1 U2535 ( .A(REG3_REG_11__SCAN_IN), .ZN(n2416) );
  NAND2_X1 U2536 ( .A1(n2258), .A2(n2013), .ZN(n2371) );
  AND2_X1 U2537 ( .A1(n2601), .A2(n2600), .ZN(n4145) );
  OR2_X1 U2538 ( .A1(n4132), .A2(n2646), .ZN(n2601) );
  AND2_X1 U2539 ( .A1(n2545), .A2(n2544), .ZN(n4215) );
  OR2_X1 U2540 ( .A1(n2447), .A2(n2309), .ZN(n2312) );
  NAND4_X2 U2541 ( .A1(n2298), .A2(n2297), .A3(n2296), .A4(n2020), .ZN(n2720)
         );
  NAND2_X1 U2542 ( .A1(n2331), .A2(REG3_REG_1__SCAN_IN), .ZN(n2297) );
  OR2_X1 U2543 ( .A1(n2447), .A2(n2923), .ZN(n2296) );
  INV_X1 U2544 ( .A(n3013), .ZN(n2130) );
  NAND2_X1 U2545 ( .A1(n2133), .A2(n2132), .ZN(n2131) );
  INV_X1 U2546 ( .A(n3002), .ZN(n2132) );
  NAND2_X1 U2547 ( .A1(n2946), .A2(n2945), .ZN(n2997) );
  NAND2_X1 U2548 ( .A1(n3157), .A2(n3156), .ZN(n3159) );
  NAND2_X1 U2549 ( .A1(n3154), .A2(n3061), .ZN(n3156) );
  OR2_X1 U2550 ( .A1(n2481), .A2(IR_REG_9__SCAN_IN), .ZN(n2278) );
  INV_X1 U2551 ( .A(IR_REG_10__SCAN_IN), .ZN(n2279) );
  NAND2_X1 U2552 ( .A1(n3427), .A2(n3435), .ZN(n2123) );
  NAND2_X1 U2553 ( .A1(n4636), .A2(n4635), .ZN(n4634) );
  NAND2_X1 U2554 ( .A1(n4079), .A2(n2142), .ZN(n2140) );
  INV_X1 U2555 ( .A(n4076), .ZN(n2112) );
  NAND2_X1 U2556 ( .A1(n2073), .A2(n2079), .ZN(n4117) );
  AND2_X1 U2557 ( .A1(n2595), .A2(n2585), .ZN(n4150) );
  AND2_X1 U2558 ( .A1(n2565), .A2(n3745), .ZN(n4225) );
  AND2_X1 U2559 ( .A1(n3722), .A2(DATAI_22_), .ZN(n3491) );
  NAND2_X1 U2560 ( .A1(n2091), .A2(n2089), .ZN(n4267) );
  INV_X1 U2561 ( .A(REG3_REG_18__SCAN_IN), .ZN(n3675) );
  INV_X1 U2562 ( .A(n2499), .ZN(n2501) );
  INV_X1 U2563 ( .A(n2471), .ZN(n2473) );
  NAND2_X1 U2564 ( .A1(n4356), .A2(n2469), .ZN(n2470) );
  NAND2_X1 U2565 ( .A1(n2091), .A2(n3828), .ZN(n4330) );
  NAND2_X1 U2566 ( .A1(n2219), .A2(n4349), .ZN(n2218) );
  INV_X1 U2567 ( .A(n2220), .ZN(n2219) );
  OR2_X1 U2568 ( .A1(n4011), .A2(n3592), .ZN(n2196) );
  AND2_X1 U2569 ( .A1(n2195), .A2(n2198), .ZN(n4415) );
  NAND2_X1 U2570 ( .A1(n4445), .A2(n2434), .ZN(n2195) );
  INV_X1 U2571 ( .A(n2209), .ZN(n2207) );
  AND2_X1 U2572 ( .A1(n3819), .A2(n3806), .ZN(n3751) );
  NAND2_X1 U2573 ( .A1(n2618), .A2(n3804), .ZN(n3800) );
  NAND2_X1 U2574 ( .A1(n2070), .A2(n3809), .ZN(n3278) );
  OR2_X1 U2575 ( .A1(n3242), .A2(n3797), .ZN(n2070) );
  AND4_X1 U2576 ( .A1(n2366), .A2(n2365), .A3(n2364), .A4(n2363), .ZN(n3292)
         );
  OR2_X1 U2577 ( .A1(n3755), .A2(n2354), .ZN(n2356) );
  NAND2_X1 U2578 ( .A1(n2258), .A2(REG3_REG_5__SCAN_IN), .ZN(n2369) );
  INV_X1 U2579 ( .A(n2615), .ZN(n3247) );
  NAND2_X1 U2580 ( .A1(REG3_REG_4__SCAN_IN), .A2(REG3_REG_3__SCAN_IN), .ZN(
        n2347) );
  INV_X1 U2581 ( .A(n3165), .ZN(n3120) );
  AND2_X1 U2582 ( .A1(n3793), .A2(n3790), .ZN(n3754) );
  NAND2_X1 U2583 ( .A1(n2610), .A2(n4088), .ZN(n4417) );
  OAI21_X1 U2584 ( .B1(n2378), .B2(n2319), .A(n2318), .ZN(n3187) );
  NAND2_X1 U2585 ( .A1(n2378), .A2(DATAI_3_), .ZN(n2318) );
  INV_X1 U2586 ( .A(n3078), .ZN(n3750) );
  OAI21_X1 U2587 ( .B1(n2378), .B2(n2300), .A(n2299), .ZN(n3221) );
  NAND2_X1 U2588 ( .A1(n2378), .A2(DATAI_0_), .ZN(n2299) );
  AND2_X1 U2589 ( .A1(n2877), .A2(n2876), .ZN(n3127) );
  INV_X1 U2590 ( .A(n4388), .ZN(n4436) );
  INV_X1 U2591 ( .A(n4442), .ZN(n4393) );
  AND2_X1 U2592 ( .A1(n2697), .A2(n2696), .ZN(n2878) );
  NOR2_X1 U2593 ( .A1(n2019), .A2(n4102), .ZN(n4101) );
  NAND2_X1 U2594 ( .A1(n4109), .A2(n4108), .ZN(n4461) );
  INV_X1 U2595 ( .A(n3026), .ZN(n2706) );
  INV_X1 U2596 ( .A(n3527), .ZN(n4198) );
  NAND2_X1 U2597 ( .A1(n3722), .A2(DATAI_24_), .ZN(n4214) );
  NAND2_X1 U2598 ( .A1(n4278), .A2(n4280), .ZN(n4279) );
  INV_X1 U2599 ( .A(n3614), .ZN(n4301) );
  INV_X1 U2600 ( .A(n4314), .ZN(n4338) );
  INV_X1 U2601 ( .A(n4373), .ZN(n4376) );
  NOR2_X1 U2602 ( .A1(n4426), .A2(n3592), .ZN(n4397) );
  OR2_X1 U2603 ( .A1(n4423), .A2(n4424), .ZN(n4426) );
  INV_X1 U2604 ( .A(n4440), .ZN(n4446) );
  NAND2_X1 U2605 ( .A1(n3220), .A2(n3087), .ZN(n3186) );
  INV_X1 U2606 ( .A(n2878), .ZN(n3128) );
  AND3_X1 U2607 ( .A1(n2694), .A2(n2693), .A3(n2877), .ZN(n2713) );
  INV_X1 U2608 ( .A(n2266), .ZN(n2660) );
  NAND2_X1 U2609 ( .A1(n2680), .A2(n2679), .ZN(n2916) );
  XNOR2_X1 U2610 ( .A(n2609), .B(n2666), .ZN(n2723) );
  MUX2_X1 U2611 ( .A(IR_REG_31__SCAN_IN), .B(n2607), .S(IR_REG_21__SCAN_IN), 
        .Z(n2608) );
  AND2_X1 U2612 ( .A1(n2497), .A2(n2507), .ZN(n4083) );
  INV_X1 U2613 ( .A(IR_REG_13__SCAN_IN), .ZN(n2239) );
  NOR2_X1 U2614 ( .A1(n2317), .A2(n2267), .ZN(n2093) );
  NAND2_X1 U2615 ( .A1(n3138), .A2(n2150), .ZN(n2147) );
  XOR2_X1 U2616 ( .A(n3563), .B(n3564), .Z(n3581) );
  NAND2_X1 U2617 ( .A1(n2820), .A2(n2819), .ZN(n3591) );
  NAND2_X1 U2618 ( .A1(n3722), .A2(DATAI_23_), .ZN(n4241) );
  AND4_X1 U2619 ( .A1(n2403), .A2(n2402), .A3(n2401), .A4(n2400), .ZN(n3396)
         );
  AOI21_X1 U2620 ( .B1(n2146), .B2(n2144), .A(n2029), .ZN(n2143) );
  NAND2_X1 U2621 ( .A1(n2378), .A2(DATAI_1_), .ZN(n2294) );
  AND2_X1 U2622 ( .A1(n2536), .A2(n2535), .ZN(n4236) );
  NAND2_X1 U2623 ( .A1(n2176), .A2(n2175), .ZN(n3362) );
  AOI21_X1 U2624 ( .B1(n3640), .B2(n3643), .A(n3641), .ZN(n3526) );
  AND2_X1 U2625 ( .A1(n3173), .A2(n2769), .ZN(n2770) );
  NOR2_X1 U2626 ( .A1(n2025), .A2(n2156), .ZN(n3635) );
  INV_X1 U2627 ( .A(n2160), .ZN(n2156) );
  NAND2_X1 U2628 ( .A1(n2232), .A2(n2857), .ZN(n2858) );
  INV_X1 U2629 ( .A(n3610), .ZN(n2857) );
  NOR2_X1 U2630 ( .A1(n3653), .A2(n3651), .ZN(n3654) );
  NAND2_X1 U2631 ( .A1(n2168), .A2(n3358), .ZN(n3443) );
  NAND2_X1 U2632 ( .A1(n2176), .A2(n2169), .ZN(n2168) );
  NOR2_X1 U2633 ( .A1(n3359), .A2(n2170), .ZN(n2169) );
  INV_X1 U2634 ( .A(n2175), .ZN(n2170) );
  AND4_X1 U2635 ( .A1(n2287), .A2(n2286), .A3(n2285), .A4(n2284), .ZN(n3386)
         );
  NAND2_X1 U2636 ( .A1(n2900), .A2(n2897), .ZN(n3655) );
  NAND2_X1 U2637 ( .A1(n2378), .A2(DATAI_2_), .ZN(n2307) );
  NAND2_X1 U2638 ( .A1(n2902), .A2(n4360), .ZN(n3700) );
  INV_X1 U2639 ( .A(n3700), .ZN(n3677) );
  INV_X1 U2640 ( .A(n3655), .ZN(n3701) );
  NAND2_X1 U2641 ( .A1(n3553), .A2(n2230), .ZN(n3685) );
  NAND2_X1 U2642 ( .A1(n2900), .A2(n2883), .ZN(n3707) );
  INV_X1 U2643 ( .A(n3691), .ZN(n3703) );
  INV_X1 U2644 ( .A(n2896), .ZN(n3867) );
  INV_X1 U2645 ( .A(n4145), .ZN(n4111) );
  INV_X1 U2646 ( .A(n4142), .ZN(n4193) );
  NAND2_X1 U2647 ( .A1(n2552), .A2(n2551), .ZN(n4217) );
  INV_X1 U2648 ( .A(n4215), .ZN(n3874) );
  INV_X1 U2649 ( .A(n4236), .ZN(n4254) );
  NAND2_X1 U2650 ( .A1(n2528), .A2(n2527), .ZN(n3663) );
  NAND2_X1 U2651 ( .A1(n2521), .A2(n2520), .ZN(n4297) );
  INV_X1 U2652 ( .A(n4414), .ZN(n4011) );
  INV_X1 U2653 ( .A(n4437), .ZN(n4387) );
  INV_X1 U2654 ( .A(n3387), .ZN(n3319) );
  OR2_X1 U2655 ( .A1(n2447), .A2(n2321), .ZN(n2324) );
  NAND2_X1 U2656 ( .A1(n2331), .A2(REG3_REG_0__SCAN_IN), .ZN(n2304) );
  OR2_X1 U2657 ( .A1(n2447), .A2(n2302), .ZN(n2305) );
  OR2_X1 U2658 ( .A1(n2890), .A2(n4690), .ZN(n4017) );
  OAI21_X1 U2659 ( .B1(n2933), .B2(REG2_REG_1__SCAN_IN), .A(n2924), .ZN(n4019)
         );
  AND2_X1 U2660 ( .A1(n2131), .A2(n2130), .ZN(n3012) );
  INV_X1 U2661 ( .A(n2131), .ZN(n3014) );
  AND2_X1 U2662 ( .A1(n2106), .A2(n2107), .ZN(n3066) );
  NAND2_X1 U2663 ( .A1(n3032), .A2(REG1_REG_6__SCAN_IN), .ZN(n2106) );
  XNOR2_X1 U2664 ( .A(n3154), .B(n3155), .ZN(n3067) );
  AND2_X1 U2665 ( .A1(n3271), .A2(REG1_REG_10__SCAN_IN), .ZN(n3343) );
  AND2_X1 U2666 ( .A1(n3335), .A2(n4617), .ZN(n3336) );
  NAND2_X1 U2667 ( .A1(n3342), .A2(n2117), .ZN(n2116) );
  INV_X1 U2668 ( .A(n3344), .ZN(n2117) );
  NOR2_X1 U2669 ( .A1(n3343), .A2(n3342), .ZN(n3345) );
  NAND2_X1 U2670 ( .A1(n2125), .A2(n2124), .ZN(n4046) );
  NAND2_X1 U2671 ( .A1(n2118), .A2(n2127), .ZN(n2126) );
  INV_X1 U2672 ( .A(n2100), .ZN(n2099) );
  AOI21_X1 U2673 ( .B1(n2100), .B2(n2098), .A(n2046), .ZN(n2097) );
  XNOR2_X1 U2674 ( .A(n4079), .B(n4612), .ZN(n4080) );
  NAND2_X1 U2675 ( .A1(n2140), .A2(n2138), .ZN(n4649) );
  AND2_X1 U2676 ( .A1(n2140), .A2(n2137), .ZN(n4650) );
  INV_X1 U2677 ( .A(n2141), .ZN(n2137) );
  INV_X1 U2678 ( .A(n2138), .ZN(n2136) );
  AOI21_X1 U2679 ( .B1(n2135), .B2(n2138), .A(n4081), .ZN(n2134) );
  INV_X1 U2680 ( .A(n2142), .ZN(n2135) );
  AND2_X1 U2681 ( .A1(n2019), .A2(n4113), .ZN(n4465) );
  NAND2_X1 U2682 ( .A1(n2202), .A2(n2582), .ZN(n4139) );
  AND2_X1 U2683 ( .A1(n2555), .A2(n2554), .ZN(n4220) );
  INV_X1 U2684 ( .A(n2059), .ZN(n3483) );
  NAND2_X1 U2685 ( .A1(n4384), .A2(n4383), .ZN(n4382) );
  NAND2_X1 U2686 ( .A1(n2192), .A2(n2191), .ZN(n4384) );
  NAND2_X1 U2687 ( .A1(n4445), .A2(n2193), .ZN(n2192) );
  NAND2_X1 U2688 ( .A1(n2208), .A2(n2222), .ZN(n3401) );
  NAND2_X1 U2689 ( .A1(n3384), .A2(n2410), .ZN(n2208) );
  INV_X1 U2690 ( .A(n4344), .ZN(n4452) );
  INV_X1 U2691 ( .A(n4358), .ZN(n4450) );
  OR2_X1 U2692 ( .A1(n3123), .A2(n2901), .ZN(n4360) );
  AND2_X1 U2693 ( .A1(n4326), .A2(n4721), .ZN(n4358) );
  AND2_X1 U2694 ( .A1(n4682), .A2(n3132), .ZN(n4680) );
  INV_X1 U2695 ( .A(n4360), .ZN(n4678) );
  INV_X1 U2696 ( .A(IR_REG_30__SCAN_IN), .ZN(n3577) );
  AND2_X1 U2697 ( .A1(n2654), .A2(n2269), .ZN(n4609) );
  INV_X1 U2698 ( .A(n4095), .ZN(n4624) );
  INV_X1 U2699 ( .A(n2676), .ZN(n2979) );
  AND2_X1 U2700 ( .A1(n2511), .A2(n2602), .ZN(n4611) );
  INV_X1 U2701 ( .A(IR_REG_9__SCAN_IN), .ZN(n2404) );
  AND2_X1 U2702 ( .A1(n2384), .A2(n2360), .ZN(n4618) );
  OR3_X1 U2703 ( .A1(n2340), .A2(IR_REG_3__SCAN_IN), .A3(IR_REG_4__SCAN_IN), 
        .ZN(n2341) );
  INV_X1 U2704 ( .A(n2110), .ZN(n2109) );
  AND2_X1 U2705 ( .A1(n2710), .A2(n2709), .ZN(n2711) );
  NAND2_X1 U2706 ( .A1(n2708), .A2(n2707), .ZN(n2710) );
  AOI21_X1 U2707 ( .B1(n2708), .B2(n2716), .A(n2715), .ZN(n2717) );
  NOR2_X1 U2708 ( .A1(n4731), .A2(n2714), .ZN(n2715) );
  AND3_X1 U2709 ( .A1(n2061), .A2(n2376), .A3(n2014), .ZN(n2266) );
  AND2_X1 U2710 ( .A1(n2212), .A2(n3420), .ZN(n2010) );
  NOR2_X1 U2711 ( .A1(n4658), .A2(n2112), .ZN(n2011) );
  NAND2_X1 U2712 ( .A1(n2061), .A2(n2376), .ZN(n2495) );
  OR2_X1 U2713 ( .A1(n2663), .A2(IR_REG_21__SCAN_IN), .ZN(n2012) );
  AND2_X1 U2714 ( .A1(n4278), .A2(n2047), .ZN(n3490) );
  INV_X1 U2715 ( .A(n4383), .ZN(n2190) );
  OAI21_X1 U2716 ( .B1(n2378), .B2(n2308), .A(n2307), .ZN(n2742) );
  AND2_X1 U2717 ( .A1(REG3_REG_5__SCAN_IN), .A2(REG3_REG_6__SCAN_IN), .ZN(
        n2013) );
  AND4_X1 U2718 ( .A1(n2252), .A2(n2251), .A3(n2250), .A4(n2249), .ZN(n2014)
         );
  AND2_X1 U2719 ( .A1(n4170), .A2(n4148), .ZN(n2703) );
  AND2_X1 U2720 ( .A1(n4446), .A2(n4413), .ZN(n2433) );
  AND2_X1 U2721 ( .A1(n2051), .A2(n2212), .ZN(n3402) );
  NAND2_X1 U2722 ( .A1(n2051), .A2(n3382), .ZN(n3381) );
  AND2_X1 U2723 ( .A1(n3722), .A2(DATAI_27_), .ZN(n3845) );
  INV_X1 U2724 ( .A(REG3_REG_14__SCAN_IN), .ZN(n2261) );
  AND2_X1 U2725 ( .A1(n2051), .A2(n2010), .ZN(n3419) );
  INV_X1 U2726 ( .A(n3809), .ZN(n2069) );
  AND2_X1 U2727 ( .A1(REG3_REG_14__SCAN_IN), .A2(REG3_REG_15__SCAN_IN), .ZN(
        n2015) );
  NOR2_X1 U2728 ( .A1(n4426), .A2(n2217), .ZN(n4314) );
  AND2_X1 U2729 ( .A1(n2057), .A2(REG3_REG_22__SCAN_IN), .ZN(n2016) );
  INV_X1 U2730 ( .A(n3741), .ZN(n2084) );
  AND2_X1 U2731 ( .A1(n4280), .A2(n4251), .ZN(n2017) );
  XOR2_X1 U2732 ( .A(n4611), .B(REG1_REG_19__SCAN_IN), .Z(n2018) );
  XNOR2_X1 U2733 ( .A(n2604), .B(n2603), .ZN(n2611) );
  OR2_X1 U2734 ( .A1(n4197), .A2(n2214), .ZN(n2019) );
  OR2_X1 U2735 ( .A1(n2301), .A2(n2295), .ZN(n2020) );
  INV_X1 U2736 ( .A(n2378), .ZN(n2344) );
  NAND2_X1 U2737 ( .A1(n3660), .A2(n3661), .ZN(n3598) );
  OAI21_X1 U2738 ( .B1(n3722), .B2(n2408), .A(n2407), .ZN(n3382) );
  OR2_X1 U2739 ( .A1(n2592), .A2(n2201), .ZN(n2021) );
  NAND2_X1 U2740 ( .A1(n3064), .A2(n4739), .ZN(n2022) );
  NAND2_X1 U2741 ( .A1(n4646), .A2(n2011), .ZN(n2023) );
  NAND2_X1 U2742 ( .A1(n2890), .A2(n3131), .ZN(n2729) );
  NAND2_X1 U2743 ( .A1(n2085), .A2(n3741), .ZN(n4210) );
  OR2_X1 U2744 ( .A1(n4165), .A2(n4148), .ZN(n2024) );
  AND3_X1 U2745 ( .A1(n2820), .A2(n2819), .A3(n2159), .ZN(n2025) );
  AND2_X1 U2746 ( .A1(n3746), .A2(n4437), .ZN(n2026) );
  AND3_X1 U2747 ( .A1(n2820), .A2(n2819), .A3(n2161), .ZN(n2027) );
  AND2_X1 U2748 ( .A1(n4140), .A2(n3844), .ZN(n2028) );
  NAND2_X1 U2749 ( .A1(n2205), .A2(n2486), .ZN(n4320) );
  OAI21_X1 U2750 ( .B1(n4157), .B2(n2021), .A(n2200), .ZN(n4109) );
  AND2_X1 U2751 ( .A1(n2785), .A2(n2784), .ZN(n2029) );
  INV_X1 U2752 ( .A(n3213), .ZN(n2699) );
  INV_X1 U2753 ( .A(IR_REG_2__SCAN_IN), .ZN(n2092) );
  AND2_X1 U2754 ( .A1(n3398), .A2(n4014), .ZN(n2030) );
  AND2_X1 U2755 ( .A1(n4217), .A2(n3527), .ZN(n2031) );
  AND2_X1 U2756 ( .A1(n2189), .A2(n2196), .ZN(n2032) );
  INV_X1 U2757 ( .A(n2194), .ZN(n2193) );
  NAND2_X1 U2758 ( .A1(n2197), .A2(n2434), .ZN(n2194) );
  OR3_X1 U2759 ( .A1(n4197), .A2(n2213), .A3(n3686), .ZN(n2033) );
  OR2_X1 U2760 ( .A1(n2433), .A2(n2026), .ZN(n2034) );
  AND2_X1 U2761 ( .A1(n4165), .A2(n3845), .ZN(n2035) );
  AND2_X1 U2762 ( .A1(n2146), .A2(n3212), .ZN(n2036) );
  OR2_X1 U2763 ( .A1(n3005), .A2(n2130), .ZN(n2037) );
  AND2_X1 U2764 ( .A1(n2222), .A2(n2211), .ZN(n2038) );
  AND2_X1 U2765 ( .A1(n2022), .A2(REG1_REG_6__SCAN_IN), .ZN(n2039) );
  AND2_X1 U2766 ( .A1(n2265), .A2(n2186), .ZN(n2040) );
  INV_X1 U2767 ( .A(IR_REG_26__SCAN_IN), .ZN(n2186) );
  INV_X1 U2768 ( .A(IR_REG_31__SCAN_IN), .ZN(n2267) );
  XNOR2_X1 U2769 ( .A(n2468), .B(IR_REG_16__SCAN_IN), .ZN(n4612) );
  INV_X1 U2770 ( .A(n3440), .ZN(n2172) );
  INV_X1 U2771 ( .A(n3651), .ZN(n2182) );
  XNOR2_X1 U2772 ( .A(n2670), .B(IR_REG_24__SCAN_IN), .ZN(n2677) );
  NOR2_X1 U2773 ( .A1(n4316), .A2(n3614), .ZN(n4278) );
  NAND2_X1 U2774 ( .A1(n2145), .A2(n2143), .ZN(n3256) );
  NAND2_X1 U2775 ( .A1(n4278), .A2(n2017), .ZN(n2041) );
  NOR2_X1 U2776 ( .A1(n4426), .A2(n2220), .ZN(n4355) );
  INV_X1 U2777 ( .A(n3632), .ZN(n2155) );
  INV_X1 U2778 ( .A(n3427), .ZN(n2127) );
  AND2_X1 U2779 ( .A1(n4616), .A2(REG2_REG_11__SCAN_IN), .ZN(n3427) );
  NAND4_X1 U2780 ( .A1(n2306), .A2(n2305), .A3(n2304), .A4(n2303), .ZN(n3024)
         );
  AND2_X1 U2781 ( .A1(n3490), .A2(n4241), .ZN(n4208) );
  NAND2_X1 U2782 ( .A1(n2147), .A2(n2149), .ZN(n3211) );
  INV_X1 U2783 ( .A(n3828), .ZN(n2090) );
  INV_X1 U2784 ( .A(n3766), .ZN(n2644) );
  INV_X1 U2785 ( .A(n3810), .ZN(n2072) );
  INV_X1 U2786 ( .A(n3799), .ZN(n2068) );
  AND2_X1 U2787 ( .A1(n3722), .A2(DATAI_28_), .ZN(n4110) );
  INV_X1 U2788 ( .A(n2884), .ZN(n2184) );
  AND2_X1 U2789 ( .A1(n3722), .A2(DATAI_21_), .ZN(n4257) );
  NAND2_X1 U2790 ( .A1(n3173), .A2(n3172), .ZN(n2042) );
  NAND2_X1 U2791 ( .A1(n3375), .A2(n3374), .ZN(n2043) );
  AND2_X1 U2792 ( .A1(n4615), .A2(REG1_REG_13__SCAN_IN), .ZN(n2044) );
  AND2_X1 U2793 ( .A1(n3429), .A2(n2127), .ZN(n2045) );
  NOR2_X1 U2794 ( .A1(n4061), .A2(n2102), .ZN(n2046) );
  INV_X1 U2795 ( .A(REG3_REG_16__SCAN_IN), .ZN(n2457) );
  AOI21_X1 U2796 ( .B1(n3797), .B2(n3809), .A(n2072), .ZN(n2071) );
  AND2_X1 U2797 ( .A1(n2017), .A2(n2702), .ZN(n2047) );
  AND2_X1 U2798 ( .A1(n2015), .A2(REG3_REG_16__SCAN_IN), .ZN(n2048) );
  INV_X1 U2799 ( .A(n2433), .ZN(n2198) );
  OR2_X1 U2800 ( .A1(n4426), .A2(n2218), .ZN(n2049) );
  NAND2_X1 U2801 ( .A1(n2706), .A2(n2611), .ZN(n2725) );
  NOR2_X1 U2802 ( .A1(n3186), .A2(n3187), .ZN(n3119) );
  NOR2_X1 U2803 ( .A1(n3246), .A2(n3247), .ZN(n2050) );
  AND2_X1 U2804 ( .A1(n3195), .A2(n2787), .ZN(n2051) );
  INV_X1 U2805 ( .A(REG3_REG_20__SCAN_IN), .ZN(n2058) );
  OR2_X1 U2806 ( .A1(n4639), .A2(n4066), .ZN(n2052) );
  NAND2_X1 U2807 ( .A1(n4417), .A2(n4703), .ZN(n4724) );
  NAND2_X1 U2808 ( .A1(n2674), .A2(n2255), .ZN(n2907) );
  INV_X1 U2809 ( .A(REG3_REG_15__SCAN_IN), .ZN(n2056) );
  INV_X1 U2810 ( .A(n3845), .ZN(n4148) );
  NAND2_X1 U2811 ( .A1(n2937), .A2(n2936), .ZN(n4021) );
  AND2_X1 U2812 ( .A1(n4083), .A2(REG1_REG_18__SCAN_IN), .ZN(n2053) );
  OR2_X1 U2813 ( .A1(n2018), .A2(n2053), .ZN(n2054) );
  AND2_X1 U2814 ( .A1(n2011), .A2(n2018), .ZN(n2055) );
  INV_X1 U2815 ( .A(REG1_REG_10__SCAN_IN), .ZN(n2115) );
  NAND2_X1 U2816 ( .A1(n2916), .A2(STATE_REG_SCAN_IN), .ZN(n4690) );
  NAND2_X1 U2817 ( .A1(n2678), .A2(n2677), .ZN(n2890) );
  NAND2_X1 U2818 ( .A1(n2513), .A2(n2057), .ZN(n2530) );
  NAND2_X1 U2819 ( .A1(n2513), .A2(REG3_REG_20__SCAN_IN), .ZN(n2522) );
  NAND3_X1 U2820 ( .A1(n2258), .A2(n2013), .A3(REG3_REG_7__SCAN_IN), .ZN(n2388) );
  NAND4_X1 U2821 ( .A1(n2061), .A2(n2376), .A3(n2221), .A4(n2014), .ZN(n2269)
         );
  NOR2_X2 U2822 ( .A1(n2480), .A2(n2248), .ZN(n2061) );
  NAND2_X1 U2823 ( .A1(n2065), .A2(n2062), .ZN(n3291) );
  NOR2_X1 U2824 ( .A1(n2071), .A2(n2619), .ZN(n2064) );
  NAND3_X1 U2825 ( .A1(n3242), .A2(n2067), .A3(n2618), .ZN(n2065) );
  OAI21_X1 U2826 ( .B1(n3242), .B2(n2066), .A(n2067), .ZN(n3191) );
  INV_X1 U2827 ( .A(n2071), .ZN(n2066) );
  NAND2_X1 U2828 ( .A1(n4160), .A2(n2080), .ZN(n2073) );
  OAI21_X1 U2829 ( .B1(n4160), .B2(n2077), .A(n2074), .ZN(n2078) );
  AOI21_X1 U2830 ( .B1(n4160), .B2(n3851), .A(n3731), .ZN(n4141) );
  XNOR2_X1 U2831 ( .A(n2078), .B(n4118), .ZN(n4124) );
  NAND2_X1 U2832 ( .A1(n2085), .A2(n2083), .ZN(n4186) );
  OAI21_X1 U2833 ( .B1(n4346), .B2(n2088), .A(n2086), .ZN(n2639) );
  NAND2_X1 U2834 ( .A1(n4636), .A2(n2096), .ZN(n2094) );
  OAI211_X1 U2835 ( .C1(n4636), .C2(n2099), .A(n2097), .B(n2094), .ZN(n4075)
         );
  INV_X1 U2836 ( .A(n4612), .ZN(n2102) );
  NAND2_X1 U2837 ( .A1(n3032), .A2(n2039), .ZN(n2103) );
  NAND2_X1 U2838 ( .A1(n3031), .A2(n4619), .ZN(n2107) );
  NAND2_X1 U2839 ( .A1(n4646), .A2(n2055), .ZN(n2108) );
  OAI211_X1 U2840 ( .C1(n4646), .C2(n2054), .A(n2109), .B(n2108), .ZN(n4092)
         );
  NAND2_X1 U2841 ( .A1(n4646), .A2(n4076), .ZN(n4659) );
  NAND2_X1 U2842 ( .A1(n3271), .A2(n2114), .ZN(n2113) );
  NAND2_X1 U2843 ( .A1(n2116), .A2(n2113), .ZN(n3434) );
  NAND3_X1 U2844 ( .A1(n2122), .A2(n2120), .A3(n2119), .ZN(n2125) );
  NAND2_X1 U2845 ( .A1(n3428), .A2(n3435), .ZN(n2119) );
  INV_X1 U2846 ( .A(n3428), .ZN(n2118) );
  NAND3_X1 U2847 ( .A1(n2122), .A2(n2123), .A3(n2119), .ZN(n3457) );
  NAND2_X1 U2848 ( .A1(n2126), .A2(n3435), .ZN(n2124) );
  NAND2_X1 U2849 ( .A1(n2129), .A2(n2133), .ZN(n2128) );
  NAND2_X1 U2850 ( .A1(n2128), .A2(n2037), .ZN(n3035) );
  NAND2_X1 U2851 ( .A1(n3138), .A2(n2036), .ZN(n2145) );
  NAND3_X1 U2852 ( .A1(n2820), .A2(n2819), .A3(n2154), .ZN(n2153) );
  NAND2_X1 U2853 ( .A1(n3309), .A2(n2177), .ZN(n2176) );
  INV_X1 U2854 ( .A(n2164), .ZN(n2817) );
  AOI21_X1 U2855 ( .B1(n3309), .B2(n2166), .A(n2165), .ZN(n2164) );
  NAND2_X1 U2856 ( .A1(n2266), .A2(n2040), .ZN(n2674) );
  NAND2_X1 U2857 ( .A1(n4445), .A2(n2188), .ZN(n2187) );
  NOR2_X1 U2858 ( .A1(n2199), .A2(n2035), .ZN(n2200) );
  NAND2_X1 U2859 ( .A1(n4157), .A2(n2581), .ZN(n2202) );
  NAND2_X1 U2860 ( .A1(n2205), .A2(n2203), .ZN(n4321) );
  INV_X1 U2861 ( .A(n3384), .ZN(n2206) );
  AOI21_X1 U2862 ( .B1(n2206), .B2(n2038), .A(n2207), .ZN(n3413) );
  INV_X1 U2863 ( .A(n3223), .ZN(n2698) );
  INV_X1 U2864 ( .A(n3221), .ZN(n3023) );
  NAND3_X1 U2865 ( .A1(n2051), .A2(n2010), .A3(n4446), .ZN(n4423) );
  NOR2_X1 U2866 ( .A1(n4197), .A2(n3686), .ZN(n4170) );
  NAND2_X1 U2867 ( .A1(n4226), .A2(n3745), .ZN(n4249) );
  NAND2_X1 U2868 ( .A1(n2890), .A2(n2681), .ZN(n3123) );
  NAND2_X1 U2869 ( .A1(n2606), .A2(n2605), .ZN(n2663) );
  XNOR2_X1 U2870 ( .A(n2724), .B(n3561), .ZN(n2739) );
  NAND2_X1 U2871 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n2288)
         );
  NAND2_X1 U2872 ( .A1(n3500), .A2(n2775), .ZN(n3138) );
  NAND2_X1 U2873 ( .A1(n3067), .A2(REG1_REG_8__SCAN_IN), .ZN(n3157) );
  NAND2_X1 U2874 ( .A1(n4037), .A2(n2927), .ZN(n2928) );
  OR2_X1 U2875 ( .A1(n4461), .A2(n4460), .ZN(n4468) );
  XNOR2_X1 U2876 ( .A(n4117), .B(n3783), .ZN(n2658) );
  AOI21_X1 U2877 ( .B1(n3597), .B2(n3539), .A(n3549), .ZN(n3641) );
  NAND2_X1 U2878 ( .A1(n3766), .A2(n2723), .ZN(n3026) );
  AND2_X1 U2879 ( .A1(n4674), .A2(n2723), .ZN(n4712) );
  INV_X1 U2880 ( .A(n2723), .ZN(n3868) );
  AND2_X1 U2881 ( .A1(n3001), .A2(n4621), .ZN(n3002) );
  XNOR2_X1 U2882 ( .A(n3001), .B(n2947), .ZN(n3003) );
  XNOR2_X1 U2883 ( .A(n3145), .B(n3061), .ZN(n3144) );
  NAND2_X1 U2884 ( .A1(n4314), .A2(n3676), .ZN(n4316) );
  OAI21_X2 U2885 ( .B1(n3112), .B2(n2614), .A(n3796), .ZN(n3242) );
  INV_X1 U2886 ( .A(n4682), .ZN(n4431) );
  INV_X1 U2887 ( .A(n4682), .ZN(n4684) );
  AND2_X2 U2888 ( .A1(n2713), .A2(n3128), .ZN(n4731) );
  INV_X1 U2889 ( .A(n4606), .ZN(n2716) );
  AND2_X2 U2890 ( .A1(n2713), .A2(n2878), .ZN(n4741) );
  INV_X1 U2891 ( .A(n4741), .ZN(n2712) );
  INV_X1 U2892 ( .A(n4540), .ZN(n2707) );
  AND4_X1 U2893 ( .A1(n2186), .A2(n2265), .A3(n2264), .A4(n2263), .ZN(n2221)
         );
  INV_X1 U2894 ( .A(n3396), .ZN(n2409) );
  INV_X1 U2895 ( .A(n3382), .ZN(n3389) );
  INV_X1 U2896 ( .A(n4435), .ZN(n4013) );
  AND4_X1 U2897 ( .A1(n2422), .A2(n2421), .A3(n2420), .A4(n2419), .ZN(n4435)
         );
  INV_X1 U2898 ( .A(REG1_REG_5__SCAN_IN), .ZN(n4737) );
  AND2_X1 U2899 ( .A1(n2464), .A2(n2463), .ZN(n4367) );
  INV_X1 U2900 ( .A(n4367), .ZN(n2469) );
  INV_X1 U2901 ( .A(REG1_REG_7__SCAN_IN), .ZN(n4739) );
  OR2_X1 U2902 ( .A1(n2409), .A2(n3389), .ZN(n2222) );
  NAND2_X1 U2903 ( .A1(n2479), .A2(n2478), .ZN(n4347) );
  INV_X1 U2904 ( .A(n4347), .ZN(n2484) );
  OR2_X1 U2905 ( .A1(n4191), .A2(n4214), .ZN(n2223) );
  AND2_X1 U2906 ( .A1(n2382), .A2(n2381), .ZN(n2224) );
  NOR2_X1 U2907 ( .A1(n2802), .A2(n3372), .ZN(n2225) );
  NOR2_X1 U2908 ( .A1(n3316), .A2(n2802), .ZN(n2226) );
  AND2_X1 U2909 ( .A1(n3404), .A2(n3386), .ZN(n2227) );
  INV_X2 U2910 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  INV_X1 U2911 ( .A(n4336), .ZN(n2483) );
  AND2_X1 U2912 ( .A1(n2657), .A2(n2656), .ZN(n2229) );
  AND2_X1 U2913 ( .A1(n3552), .A2(n3551), .ZN(n2230) );
  OR2_X1 U2914 ( .A1(n4217), .A2(n3527), .ZN(n2231) );
  INV_X1 U2915 ( .A(n3310), .ZN(n3420) );
  AND2_X1 U2916 ( .A1(n4115), .A2(n4114), .ZN(n3783) );
  OR3_X1 U2917 ( .A1(n3611), .A2(n3607), .A3(n3670), .ZN(n2232) );
  AND2_X1 U2918 ( .A1(n3221), .A2(n3024), .ZN(n2233) );
  NAND2_X1 U2919 ( .A1(n3480), .A2(n2564), .ZN(n2234) );
  INV_X1 U2920 ( .A(n2762), .ZN(n2763) );
  INV_X1 U2921 ( .A(n3491), .ZN(n2702) );
  INV_X1 U2922 ( .A(IR_REG_0__SCAN_IN), .ZN(n2300) );
  INV_X1 U2923 ( .A(n3377), .ZN(n2794) );
  NOR2_X1 U2924 ( .A1(IR_REG_20__SCAN_IN), .A2(IR_REG_19__SCAN_IN), .ZN(n2605)
         );
  NAND2_X1 U2925 ( .A1(n2940), .A2(n2938), .ZN(n2939) );
  NAND2_X1 U2926 ( .A1(n3374), .A2(n2798), .ZN(n2802) );
  OR2_X1 U2927 ( .A1(n3547), .A2(n3546), .ZN(n3552) );
  INV_X1 U2928 ( .A(REG3_REG_27__SCAN_IN), .ZN(n2583) );
  INV_X1 U2929 ( .A(REG3_REG_25__SCAN_IN), .ZN(n3967) );
  NOR2_X1 U2930 ( .A1(n3019), .A2(n3004), .ZN(n3005) );
  INV_X1 U2931 ( .A(REG3_REG_19__SCAN_IN), .ZN(n2500) );
  INV_X1 U2932 ( .A(n3292), .ZN(n2367) );
  INV_X1 U2933 ( .A(n4110), .ZN(n3535) );
  AND2_X1 U2934 ( .A1(n3599), .A2(n3600), .ZN(n3515) );
  INV_X1 U2935 ( .A(REG3_REG_13__SCAN_IN), .ZN(n2439) );
  INV_X1 U2936 ( .A(REG3_REG_22__SCAN_IN), .ZN(n2529) );
  AND2_X1 U2937 ( .A1(n3868), .A2(n2644), .ZN(n2917) );
  INV_X1 U2938 ( .A(n4060), .ZN(n4061) );
  AND2_X1 U2939 ( .A1(n2573), .A2(n2546), .ZN(n4200) );
  NAND2_X1 U2940 ( .A1(n2565), .A2(n2234), .ZN(n4227) );
  NAND2_X1 U2941 ( .A1(n2640), .A2(n4230), .ZN(n3482) );
  NAND2_X1 U2942 ( .A1(n2499), .A2(REG3_REG_19__SCAN_IN), .ZN(n2514) );
  NAND2_X1 U2943 ( .A1(n3420), .A2(n4435), .ZN(n2423) );
  INV_X1 U2944 ( .A(n3404), .ZN(n3398) );
  OR2_X1 U2945 ( .A1(n4462), .A2(n4715), .ZN(n4460) );
  INV_X1 U2946 ( .A(n2943), .ZN(n2319) );
  AND2_X1 U2947 ( .A1(n2912), .A2(n2917), .ZN(n4388) );
  NOR2_X1 U2948 ( .A1(IR_REG_2__SCAN_IN), .A2(IR_REG_4__SCAN_IN), .ZN(n2235)
         );
  AND2_X1 U2949 ( .A1(n3569), .A2(n3673), .ZN(n3565) );
  INV_X1 U2950 ( .A(n3024), .ZN(n3047) );
  NAND2_X1 U2951 ( .A1(n2735), .A2(n2732), .ZN(n2910) );
  INV_X1 U2952 ( .A(n2260), .ZN(n2442) );
  INV_X1 U2953 ( .A(n2415), .ZN(n2427) );
  AND4_X1 U2954 ( .A1(n2393), .A2(n2392), .A3(n2391), .A4(n2390), .ZN(n3387)
         );
  AND2_X1 U2955 ( .A1(n2997), .A2(n4621), .ZN(n2998) );
  INV_X1 U2956 ( .A(n3435), .ZN(n3429) );
  INV_X1 U2957 ( .A(n4661), .ZN(n4662) );
  OR2_X1 U2958 ( .A1(n3739), .A2(n3738), .ZN(n4211) );
  INV_X1 U2959 ( .A(n3482), .ZN(n4232) );
  INV_X1 U2960 ( .A(n4356), .ZN(n4349) );
  AND2_X1 U2961 ( .A1(n3816), .A2(n3817), .ZN(n3761) );
  INV_X1 U2962 ( .A(n4386), .ZN(n4434) );
  OR2_X1 U2963 ( .A1(n2975), .A2(D_REG_1__SCAN_IN), .ZN(n3125) );
  OR2_X1 U2964 ( .A1(n2975), .A2(D_REG_0__SCAN_IN), .ZN(n2697) );
  AND2_X1 U2965 ( .A1(n3722), .A2(DATAI_30_), .ZN(n4102) );
  AND2_X1 U2966 ( .A1(n4289), .A2(n4290), .ZN(n4323) );
  INV_X1 U2967 ( .A(n3746), .ZN(n4424) );
  INV_X1 U2968 ( .A(n4712), .ZN(n4703) );
  INV_X1 U2969 ( .A(IR_REG_11__SCAN_IN), .ZN(n2412) );
  AND2_X1 U2970 ( .A1(n3570), .A2(n3565), .ZN(n3566) );
  INV_X1 U2971 ( .A(n3707), .ZN(n3673) );
  NAND2_X1 U2972 ( .A1(n2895), .A2(n3044), .ZN(n3705) );
  OAI21_X1 U2973 ( .B1(n4303), .B2(n2646), .A(n2506), .ZN(n4271) );
  AND4_X1 U2974 ( .A1(n2446), .A2(n2445), .A3(n2444), .A4(n2443), .ZN(n4437)
         );
  INV_X1 U2975 ( .A(n3277), .ZN(n2616) );
  INV_X1 U2976 ( .A(n3150), .ZN(n3153) );
  INV_X1 U2977 ( .A(n4657), .ZN(n4654) );
  AND2_X1 U2978 ( .A1(n4682), .A2(n4088), .ZN(n4326) );
  INV_X1 U2979 ( .A(n4391), .ZN(n4439) );
  INV_X1 U2980 ( .A(REG1_REG_9__SCAN_IN), .ZN(n3952) );
  NAND2_X1 U2981 ( .A1(n3722), .A2(DATAI_26_), .ZN(n4172) );
  INV_X1 U2982 ( .A(n4270), .ZN(n4280) );
  INV_X1 U2983 ( .A(n4724), .ZN(n4715) );
  INV_X1 U2984 ( .A(n2725), .ZN(n4721) );
  INV_X1 U2985 ( .A(n3123), .ZN(n2974) );
  NAND2_X1 U2986 ( .A1(n2659), .A2(n2662), .ZN(n2976) );
  AND2_X1 U2987 ( .A1(n2921), .A2(n2920), .ZN(n4660) );
  INV_X1 U2988 ( .A(n3705), .ZN(n3689) );
  INV_X1 U2989 ( .A(DATAO_REG_30__SCAN_IN), .ZN(n3979) );
  INV_X1 U2990 ( .A(n4191), .ZN(n4238) );
  INV_X1 U2991 ( .A(n4295), .ZN(n4333) );
  INV_X1 U2992 ( .A(n3386), .ZN(n4014) );
  OR2_X1 U2993 ( .A1(n4626), .A2(n3866), .ZN(n3470) );
  OR2_X1 U2994 ( .A1(n4626), .A2(n4609), .ZN(n4673) );
  NAND2_X1 U2995 ( .A1(n4682), .A2(n3206), .ZN(n4344) );
  NAND2_X1 U2996 ( .A1(n4741), .A2(n4721), .ZN(n4540) );
  INV_X1 U2997 ( .A(REG0_REG_30__SCAN_IN), .ZN(n4549) );
  OR2_X1 U2998 ( .A1(n4208), .A2(n4242), .ZN(n4567) );
  OR2_X1 U2999 ( .A1(n4355), .A2(n4377), .ZN(n4590) );
  NAND2_X1 U3000 ( .A1(n4731), .A2(n4721), .ZN(n4606) );
  INV_X1 U3001 ( .A(n4731), .ZN(n4729) );
  NAND2_X1 U3002 ( .A1(n2975), .A2(n2974), .ZN(n4689) );
  AND2_X1 U3003 ( .A1(n2424), .A2(n2414), .ZN(n4616) );
  INV_X1 U3004 ( .A(n4017), .ZN(U4043) );
  OR4_X1 U3005 ( .A1(n2906), .A2(n2905), .A3(n2904), .A4(n2903), .ZN(U3220) );
  OAI21_X1 U3006 ( .B1(n2718), .B2(n2712), .A(n2711), .ZN(U3546) );
  NOR2_X1 U3007 ( .A1(IR_REG_3__SCAN_IN), .A2(IR_REG_5__SCAN_IN), .ZN(n2236)
         );
  NAND2_X1 U3008 ( .A1(n2376), .A2(n2247), .ZN(n2357) );
  NAND2_X1 U3009 ( .A1(n2358), .A2(n2385), .ZN(n2237) );
  INV_X1 U3010 ( .A(n2278), .ZN(n2238) );
  NAND2_X1 U3011 ( .A1(n2238), .A2(n2279), .ZN(n2411) );
  INV_X1 U3012 ( .A(n2435), .ZN(n2240) );
  NAND2_X1 U3013 ( .A1(n2240), .A2(n2239), .ZN(n2452) );
  NAND2_X1 U3014 ( .A1(n2452), .A2(IR_REG_31__SCAN_IN), .ZN(n2241) );
  XNOR2_X1 U3015 ( .A(n2241), .B(IR_REG_14__SCAN_IN), .ZN(n4614) );
  NOR2_X1 U3016 ( .A1(IR_REG_12__SCAN_IN), .A2(IR_REG_9__SCAN_IN), .ZN(n2245)
         );
  NAND4_X1 U3017 ( .A1(n2245), .A2(n2244), .A3(n2243), .A4(n2242), .ZN(n2480)
         );
  NAND4_X1 U3018 ( .A1(n2385), .A2(n2247), .A3(n2358), .A4(n2246), .ZN(n2248)
         );
  NOR2_X1 U3019 ( .A1(IR_REG_21__SCAN_IN), .A2(IR_REG_20__SCAN_IN), .ZN(n2252)
         );
  NOR2_X1 U3020 ( .A1(IR_REG_18__SCAN_IN), .A2(IR_REG_19__SCAN_IN), .ZN(n2251)
         );
  NOR2_X1 U3021 ( .A1(IR_REG_22__SCAN_IN), .A2(IR_REG_23__SCAN_IN), .ZN(n2250)
         );
  NAND2_X1 U3022 ( .A1(n2254), .A2(n2264), .ZN(n2652) );
  NAND2_X1 U3023 ( .A1(n2264), .A2(n2267), .ZN(n2253) );
  NAND2_X1 U3024 ( .A1(n2907), .A2(IR_REG_28__SCAN_IN), .ZN(n2256) );
  MUX2_X1 U3025 ( .A(n4614), .B(DATAI_14_), .S(n3722), .Z(n3592) );
  INV_X1 U3026 ( .A(n2347), .ZN(n2258) );
  INV_X1 U3027 ( .A(REG3_REG_7__SCAN_IN), .ZN(n2361) );
  INV_X1 U3028 ( .A(n2399), .ZN(n2259) );
  NAND2_X1 U3029 ( .A1(n2259), .A2(REG3_REG_10__SCAN_IN), .ZN(n2417) );
  NAND2_X1 U3030 ( .A1(n2415), .A2(REG3_REG_12__SCAN_IN), .ZN(n2440) );
  NAND2_X1 U3031 ( .A1(n2442), .A2(n2261), .ZN(n2262) );
  AND2_X1 U3032 ( .A1(n2448), .A2(n2262), .ZN(n4401) );
  XNOR2_X2 U3033 ( .A(n2268), .B(n3577), .ZN(n2273) );
  INV_X2 U3034 ( .A(n2273), .ZN(n4608) );
  NAND2_X1 U3035 ( .A1(n2269), .A2(IR_REG_31__SCAN_IN), .ZN(n2270) );
  INV_X1 U3036 ( .A(n2271), .ZN(n3580) );
  NAND2_X1 U3037 ( .A1(n4401), .A2(n2331), .ZN(n2277) );
  AND2_X2 U3038 ( .A1(n2965), .A2(n2273), .ZN(n2330) );
  AOI22_X1 U3039 ( .A1(n2008), .A2(REG0_REG_14__SCAN_IN), .B1(n2009), .B2(
        REG1_REG_14__SCAN_IN), .ZN(n2276) );
  NAND2_X4 U3040 ( .A1(n4608), .A2(n2274), .ZN(n2447) );
  NAND2_X1 U3041 ( .A1(n2329), .A2(REG2_REG_14__SCAN_IN), .ZN(n2275) );
  NAND2_X1 U3042 ( .A1(n2278), .A2(IR_REG_31__SCAN_IN), .ZN(n2280) );
  XNOR2_X1 U3043 ( .A(n2280), .B(n2279), .ZN(n3334) );
  INV_X1 U3044 ( .A(DATAI_10_), .ZN(n2281) );
  MUX2_X1 U3045 ( .A(n3334), .B(n2281), .S(n3722), .Z(n3404) );
  NAND2_X1 U3046 ( .A1(n2008), .A2(REG0_REG_10__SCAN_IN), .ZN(n2287) );
  NAND2_X1 U3047 ( .A1(n2329), .A2(REG2_REG_10__SCAN_IN), .ZN(n2286) );
  NAND2_X1 U3048 ( .A1(n2009), .A2(REG1_REG_10__SCAN_IN), .ZN(n2285) );
  INV_X1 U3049 ( .A(REG3_REG_10__SCAN_IN), .ZN(n2282) );
  NAND2_X1 U3050 ( .A1(n2399), .A2(n2282), .ZN(n2283) );
  AND2_X1 U3051 ( .A1(n2417), .A2(n2283), .ZN(n3406) );
  NAND2_X1 U3052 ( .A1(n2331), .A2(n3406), .ZN(n2284) );
  INV_X1 U3053 ( .A(n2317), .ZN(n2293) );
  NAND2_X1 U3054 ( .A1(n2288), .A2(IR_REG_1__SCAN_IN), .ZN(n2291) );
  NAND2_X1 U3055 ( .A1(n2291), .A2(n2290), .ZN(n2292) );
  NAND2_X2 U3056 ( .A1(n2293), .A2(n2292), .ZN(n2933) );
  NAND2_X1 U3057 ( .A1(n2009), .A2(REG1_REG_1__SCAN_IN), .ZN(n2298) );
  INV_X1 U3058 ( .A(REG0_REG_1__SCAN_IN), .ZN(n2295) );
  NAND2_X1 U3059 ( .A1(n2008), .A2(REG0_REG_0__SCAN_IN), .ZN(n2306) );
  INV_X1 U3060 ( .A(REG2_REG_0__SCAN_IN), .ZN(n2302) );
  NAND2_X1 U3061 ( .A1(n2009), .A2(REG1_REG_0__SCAN_IN), .ZN(n2303) );
  OAI21_X1 U3062 ( .B1(n3223), .B2(n3082), .A(n2233), .ZN(n2314) );
  NAND2_X1 U3063 ( .A1(n3223), .A2(n3082), .ZN(n3073) );
  INV_X1 U3064 ( .A(n2007), .ZN(n2308) );
  NAND2_X1 U3065 ( .A1(n2008), .A2(REG0_REG_2__SCAN_IN), .ZN(n2313) );
  INV_X1 U3066 ( .A(REG2_REG_2__SCAN_IN), .ZN(n2309) );
  NAND2_X1 U3067 ( .A1(n2009), .A2(REG1_REG_2__SCAN_IN), .ZN(n2311) );
  NAND2_X1 U3068 ( .A1(n2331), .A2(REG3_REG_2__SCAN_IN), .ZN(n2310) );
  NAND2_X1 U3069 ( .A1(n2742), .A2(n2315), .ZN(n3788) );
  NAND2_X1 U3070 ( .A1(n3791), .A2(n3788), .ZN(n3078) );
  NAND3_X1 U3071 ( .A1(n2314), .A2(n3073), .A3(n3078), .ZN(n3075) );
  NAND2_X1 U3072 ( .A1(n3087), .A2(n2315), .ZN(n2316) );
  NAND2_X1 U3073 ( .A1(n3075), .A2(n2316), .ZN(n3179) );
  NAND2_X1 U3074 ( .A1(n2317), .A2(n2092), .ZN(n2340) );
  NAND2_X1 U3075 ( .A1(n2340), .A2(IR_REG_31__SCAN_IN), .ZN(n2337) );
  XNOR2_X1 U3076 ( .A(n2337), .B(IR_REG_3__SCAN_IN), .ZN(n2943) );
  INV_X1 U3077 ( .A(REG3_REG_3__SCAN_IN), .ZN(n2320) );
  NAND2_X1 U3078 ( .A1(n2331), .A2(n2320), .ZN(n2325) );
  INV_X1 U3079 ( .A(REG2_REG_3__SCAN_IN), .ZN(n2321) );
  NAND2_X1 U3080 ( .A1(n2009), .A2(REG1_REG_3__SCAN_IN), .ZN(n2323) );
  NAND2_X1 U3081 ( .A1(n2008), .A2(REG0_REG_3__SCAN_IN), .ZN(n2322) );
  NAND2_X1 U3082 ( .A1(n3187), .A2(n4016), .ZN(n2326) );
  NAND2_X1 U3083 ( .A1(n3179), .A2(n2326), .ZN(n2328) );
  INV_X1 U3084 ( .A(n3187), .ZN(n3106) );
  NAND2_X1 U3085 ( .A1(n3106), .A2(n3168), .ZN(n2327) );
  NAND2_X1 U3086 ( .A1(n2328), .A2(n2327), .ZN(n3114) );
  NAND2_X1 U3087 ( .A1(n2008), .A2(REG0_REG_4__SCAN_IN), .ZN(n2335) );
  NAND2_X1 U3088 ( .A1(n2329), .A2(REG2_REG_4__SCAN_IN), .ZN(n2334) );
  NAND2_X1 U3089 ( .A1(n2009), .A2(REG1_REG_4__SCAN_IN), .ZN(n2333) );
  OAI21_X1 U3090 ( .B1(REG3_REG_3__SCAN_IN), .B2(REG3_REG_4__SCAN_IN), .A(
        n2347), .ZN(n3121) );
  INV_X1 U3091 ( .A(n3121), .ZN(n3177) );
  NAND2_X1 U3092 ( .A1(n2331), .A2(n3177), .ZN(n2332) );
  INV_X1 U3093 ( .A(IR_REG_3__SCAN_IN), .ZN(n2336) );
  NAND2_X1 U3094 ( .A1(n2337), .A2(n2336), .ZN(n2338) );
  NAND2_X1 U3095 ( .A1(n2338), .A2(IR_REG_31__SCAN_IN), .ZN(n2339) );
  XNOR2_X1 U3096 ( .A(n2339), .B(IR_REG_4__SCAN_IN), .ZN(n4621) );
  MUX2_X1 U3097 ( .A(n4621), .B(DATAI_4_), .S(n2378), .Z(n3165) );
  NAND2_X1 U3098 ( .A1(n3165), .A2(n3502), .ZN(n3794) );
  NAND2_X1 U3099 ( .A1(n2341), .A2(IR_REG_31__SCAN_IN), .ZN(n2343) );
  INV_X1 U3100 ( .A(IR_REG_5__SCAN_IN), .ZN(n2342) );
  XNOR2_X1 U3101 ( .A(n2343), .B(n2342), .ZN(n3019) );
  INV_X1 U3102 ( .A(DATAI_5_), .ZN(n2345) );
  MUX2_X1 U3103 ( .A(n3019), .B(n2345), .S(n2378), .Z(n2615) );
  NAND2_X1 U3104 ( .A1(n2008), .A2(REG0_REG_5__SCAN_IN), .ZN(n2352) );
  NAND2_X1 U3105 ( .A1(n2329), .A2(REG2_REG_5__SCAN_IN), .ZN(n2351) );
  NAND2_X1 U3106 ( .A1(n2009), .A2(REG1_REG_5__SCAN_IN), .ZN(n2350) );
  INV_X1 U3107 ( .A(REG3_REG_5__SCAN_IN), .ZN(n2346) );
  NAND2_X1 U3108 ( .A1(n2347), .A2(n2346), .ZN(n2348) );
  AND2_X1 U3109 ( .A1(n2369), .A2(n2348), .ZN(n3498) );
  NAND2_X1 U3110 ( .A1(n2331), .A2(n3498), .ZN(n2349) );
  AND2_X1 U3111 ( .A1(n2615), .A2(n3277), .ZN(n2354) );
  NAND2_X1 U3112 ( .A1(n3165), .A2(n2985), .ZN(n3239) );
  NAND2_X1 U3113 ( .A1(n3247), .A2(n2616), .ZN(n2353) );
  AND2_X1 U3114 ( .A1(n3239), .A2(n2353), .ZN(n2355) );
  NAND2_X1 U3115 ( .A1(n2357), .A2(IR_REG_31__SCAN_IN), .ZN(n2359) );
  NAND2_X1 U3116 ( .A1(n2359), .A2(n2358), .ZN(n2384) );
  OR2_X1 U3117 ( .A1(n2359), .A2(n2358), .ZN(n2360) );
  MUX2_X1 U3118 ( .A(n4618), .B(DATAI_7_), .S(n2378), .Z(n3213) );
  NAND2_X1 U3119 ( .A1(n2008), .A2(REG0_REG_7__SCAN_IN), .ZN(n2366) );
  NAND2_X1 U3120 ( .A1(n2329), .A2(REG2_REG_7__SCAN_IN), .ZN(n2365) );
  NAND2_X1 U3121 ( .A1(n2009), .A2(REG1_REG_7__SCAN_IN), .ZN(n2364) );
  NAND2_X1 U3122 ( .A1(n2371), .A2(n2361), .ZN(n2362) );
  AND2_X1 U3123 ( .A1(n2388), .A2(n2362), .ZN(n3217) );
  NAND2_X1 U3124 ( .A1(n2331), .A2(n3217), .ZN(n2363) );
  NAND2_X1 U3125 ( .A1(n3213), .A2(n3292), .ZN(n2618) );
  NAND2_X1 U3126 ( .A1(n2009), .A2(REG1_REG_6__SCAN_IN), .ZN(n2375) );
  INV_X1 U3127 ( .A(REG3_REG_6__SCAN_IN), .ZN(n2368) );
  NAND2_X1 U3128 ( .A1(n2369), .A2(n2368), .ZN(n2370) );
  AND2_X1 U3129 ( .A1(n2371), .A2(n2370), .ZN(n3286) );
  NAND2_X1 U3130 ( .A1(n2331), .A2(n3286), .ZN(n2374) );
  NAND2_X1 U3131 ( .A1(n2008), .A2(REG0_REG_6__SCAN_IN), .ZN(n2373) );
  NAND2_X1 U3132 ( .A1(n2329), .A2(REG2_REG_6__SCAN_IN), .ZN(n2372) );
  OR2_X1 U3133 ( .A1(n2376), .A2(n2267), .ZN(n2377) );
  XNOR2_X1 U3134 ( .A(n2377), .B(IR_REG_6__SCAN_IN), .ZN(n4619) );
  MUX2_X1 U3135 ( .A(n4619), .B(DATAI_6_), .S(n2378), .Z(n3282) );
  NAND2_X1 U3136 ( .A1(n3283), .A2(n2380), .ZN(n2383) );
  NAND3_X1 U3137 ( .A1(n3800), .A2(n3282), .A3(n4015), .ZN(n2382) );
  NAND2_X1 U3138 ( .A1(n3213), .A2(n2367), .ZN(n2381) );
  NAND2_X1 U3139 ( .A1(n2383), .A2(n2224), .ZN(n3296) );
  NAND2_X1 U3140 ( .A1(n2384), .A2(IR_REG_31__SCAN_IN), .ZN(n2386) );
  XNOR2_X1 U3141 ( .A(n2386), .B(n2385), .ZN(n3155) );
  INV_X1 U3142 ( .A(DATAI_8_), .ZN(n2955) );
  MUX2_X1 U3143 ( .A(n3155), .B(n2955), .S(n3722), .Z(n2787) );
  NAND2_X1 U3144 ( .A1(n2008), .A2(REG0_REG_8__SCAN_IN), .ZN(n2393) );
  NAND2_X1 U3145 ( .A1(n2329), .A2(REG2_REG_8__SCAN_IN), .ZN(n2392) );
  NAND2_X1 U3146 ( .A1(n2009), .A2(REG1_REG_8__SCAN_IN), .ZN(n2391) );
  NAND2_X1 U3147 ( .A1(n2388), .A2(n2387), .ZN(n2389) );
  AND2_X1 U31480 ( .A1(n2397), .A2(n2389), .ZN(n3299) );
  NAND2_X1 U31490 ( .A1(n2331), .A2(n3299), .ZN(n2390) );
  NAND2_X1 U3150 ( .A1(n2787), .A2(n3387), .ZN(n2395) );
  INV_X1 U3151 ( .A(n2787), .ZN(n3298) );
  NAND2_X1 U3152 ( .A1(n2008), .A2(REG0_REG_9__SCAN_IN), .ZN(n2403) );
  NAND2_X1 U3153 ( .A1(n2329), .A2(REG2_REG_9__SCAN_IN), .ZN(n2402) );
  NAND2_X1 U3154 ( .A1(n2009), .A2(REG1_REG_9__SCAN_IN), .ZN(n2401) );
  NAND2_X1 U3155 ( .A1(n2397), .A2(n2396), .ZN(n2398) );
  AND2_X1 U3156 ( .A1(n2399), .A2(n2398), .ZN(n3448) );
  NAND2_X1 U3157 ( .A1(n2331), .A2(n3448), .ZN(n2400) );
  NAND2_X1 U3158 ( .A1(n2481), .A2(IR_REG_31__SCAN_IN), .ZN(n2405) );
  XNOR2_X1 U3159 ( .A(n2405), .B(n2404), .ZN(n3268) );
  INV_X1 U3160 ( .A(DATAI_9_), .ZN(n2406) );
  NAND2_X1 U3161 ( .A1(n2411), .A2(IR_REG_31__SCAN_IN), .ZN(n2413) );
  NAND2_X1 U3162 ( .A1(n2413), .A2(n2412), .ZN(n2424) );
  OR2_X1 U3163 ( .A1(n2413), .A2(n2412), .ZN(n2414) );
  MUX2_X1 U3164 ( .A(n4616), .B(DATAI_11_), .S(n3722), .Z(n3310) );
  NAND2_X1 U3165 ( .A1(n2008), .A2(REG0_REG_11__SCAN_IN), .ZN(n2422) );
  NAND2_X1 U3166 ( .A1(n2329), .A2(REG2_REG_11__SCAN_IN), .ZN(n2421) );
  NAND2_X1 U3167 ( .A1(n2009), .A2(REG1_REG_11__SCAN_IN), .ZN(n2420) );
  NAND2_X1 U3168 ( .A1(n2417), .A2(n2416), .ZN(n2418) );
  AND2_X1 U3169 ( .A1(n2427), .A2(n2418), .ZN(n3422) );
  NAND2_X1 U3170 ( .A1(n2331), .A2(n3422), .ZN(n2419) );
  NAND2_X1 U3171 ( .A1(n3310), .A2(n4435), .ZN(n4406) );
  NAND2_X1 U3172 ( .A1(n3420), .A2(n4013), .ZN(n4408) );
  NAND2_X1 U3173 ( .A1(n4406), .A2(n4408), .ZN(n3753) );
  NAND2_X1 U3174 ( .A1(n3413), .A2(n3753), .ZN(n3412) );
  NAND2_X1 U3175 ( .A1(n3412), .A2(n2423), .ZN(n4445) );
  NAND2_X1 U3176 ( .A1(n2424), .A2(IR_REG_31__SCAN_IN), .ZN(n2425) );
  XNOR2_X1 U3177 ( .A(n2425), .B(IR_REG_12__SCAN_IN), .ZN(n3435) );
  MUX2_X1 U3178 ( .A(n3435), .B(DATAI_12_), .S(n3722), .Z(n4440) );
  NAND2_X1 U3179 ( .A1(n2009), .A2(REG1_REG_12__SCAN_IN), .ZN(n2432) );
  INV_X1 U3180 ( .A(REG3_REG_12__SCAN_IN), .ZN(n2426) );
  NAND2_X1 U3181 ( .A1(n2427), .A2(n2426), .ZN(n2428) );
  AND2_X1 U3182 ( .A1(n2440), .A2(n2428), .ZN(n4448) );
  NAND2_X1 U3183 ( .A1(n2331), .A2(n4448), .ZN(n2431) );
  NAND2_X1 U3184 ( .A1(n2008), .A2(REG0_REG_12__SCAN_IN), .ZN(n2430) );
  NAND2_X1 U3185 ( .A1(n2329), .A2(REG2_REG_12__SCAN_IN), .ZN(n2429) );
  NAND4_X1 U3186 ( .A1(n2432), .A2(n2431), .A3(n2430), .A4(n2429), .ZN(n4012)
         );
  NAND2_X1 U3187 ( .A1(n4440), .A2(n4012), .ZN(n2434) );
  INV_X1 U3188 ( .A(n4012), .ZN(n4413) );
  NAND2_X1 U3189 ( .A1(n2435), .A2(IR_REG_31__SCAN_IN), .ZN(n2436) );
  MUX2_X1 U3190 ( .A(IR_REG_31__SCAN_IN), .B(n2436), .S(IR_REG_13__SCAN_IN), 
        .Z(n2437) );
  NAND2_X1 U3191 ( .A1(n2437), .A2(n2452), .ZN(n4044) );
  INV_X1 U3192 ( .A(DATAI_13_), .ZN(n2438) );
  MUX2_X1 U3193 ( .A(n4044), .B(n2438), .S(n3722), .Z(n3746) );
  NAND2_X1 U3194 ( .A1(n2440), .A2(n2439), .ZN(n2441) );
  AND2_X1 U3195 ( .A1(n2442), .A2(n2441), .ZN(n4427) );
  NAND2_X1 U3196 ( .A1(n4427), .A2(n2331), .ZN(n2446) );
  NAND2_X1 U3197 ( .A1(n2008), .A2(REG0_REG_13__SCAN_IN), .ZN(n2445) );
  NAND2_X1 U3198 ( .A1(n2329), .A2(REG2_REG_13__SCAN_IN), .ZN(n2444) );
  NAND2_X1 U3199 ( .A1(n2009), .A2(REG1_REG_13__SCAN_IN), .ZN(n2443) );
  NAND2_X1 U3200 ( .A1(n4414), .A2(n3592), .ZN(n4368) );
  INV_X1 U3201 ( .A(n3592), .ZN(n4399) );
  NAND2_X1 U3202 ( .A1(n4011), .A2(n4399), .ZN(n3710) );
  NAND2_X1 U3203 ( .A1(n4368), .A2(n3710), .ZN(n4383) );
  INV_X1 U3204 ( .A(REG2_REG_15__SCAN_IN), .ZN(n4066) );
  NAND2_X1 U3205 ( .A1(n2448), .A2(n2056), .ZN(n2449) );
  NAND2_X1 U3206 ( .A1(n2458), .A2(n2449), .ZN(n3699) );
  OR2_X1 U3207 ( .A1(n3699), .A2(n2646), .ZN(n2451) );
  AOI22_X1 U3208 ( .A1(n2008), .A2(REG0_REG_15__SCAN_IN), .B1(n2009), .B2(
        REG1_REG_15__SCAN_IN), .ZN(n2450) );
  OAI211_X1 U3209 ( .C1(n2447), .C2(n4066), .A(n2451), .B(n2450), .ZN(n4389)
         );
  INV_X1 U32100 ( .A(n2452), .ZN(n2453) );
  NAND2_X1 U32110 ( .A1(n2453), .A2(n3884), .ZN(n2454) );
  NAND2_X1 U32120 ( .A1(n2454), .A2(IR_REG_31__SCAN_IN), .ZN(n2466) );
  XNOR2_X1 U32130 ( .A(n2466), .B(IR_REG_15__SCAN_IN), .ZN(n4613) );
  MUX2_X1 U32140 ( .A(DATAI_15_), .B(n4613), .S(n2344), .Z(n4373) );
  NAND2_X1 U32150 ( .A1(n4389), .A2(n4373), .ZN(n2456) );
  NOR2_X1 U32160 ( .A1(n4389), .A2(n4373), .ZN(n2455) );
  AOI21_X1 U32170 ( .B1(n4375), .B2(n2456), .A(n2455), .ZN(n4354) );
  NAND2_X1 U32180 ( .A1(n2458), .A2(n2457), .ZN(n2459) );
  AND2_X1 U32190 ( .A1(n2473), .A2(n2459), .ZN(n4359) );
  NAND2_X1 U32200 ( .A1(n4359), .A2(n2331), .ZN(n2464) );
  INV_X1 U32210 ( .A(REG2_REG_16__SCAN_IN), .ZN(n4362) );
  NAND2_X1 U32220 ( .A1(n2008), .A2(REG0_REG_16__SCAN_IN), .ZN(n2461) );
  NAND2_X1 U32230 ( .A1(n2009), .A2(REG1_REG_16__SCAN_IN), .ZN(n2460) );
  OAI211_X1 U32240 ( .C1(n4362), .C2(n2447), .A(n2461), .B(n2460), .ZN(n2462)
         );
  INV_X1 U32250 ( .A(n2462), .ZN(n2463) );
  INV_X1 U32260 ( .A(IR_REG_15__SCAN_IN), .ZN(n2465) );
  NAND2_X1 U32270 ( .A1(n2466), .A2(n2465), .ZN(n2467) );
  NAND2_X1 U32280 ( .A1(n2467), .A2(IR_REG_31__SCAN_IN), .ZN(n2468) );
  MUX2_X1 U32290 ( .A(DATAI_16_), .B(n4612), .S(n2344), .Z(n4356) );
  NAND2_X1 U32300 ( .A1(n4367), .A2(n4356), .ZN(n3832) );
  NAND2_X1 U32310 ( .A1(n2469), .A2(n4349), .ZN(n3828) );
  NAND2_X1 U32320 ( .A1(n3832), .A2(n3828), .ZN(n4353) );
  NAND2_X1 U32330 ( .A1(n4354), .A2(n4353), .ZN(n4352) );
  NAND2_X1 U32340 ( .A1(n4352), .A2(n2470), .ZN(n4329) );
  NAND2_X1 U32350 ( .A1(n2471), .A2(REG3_REG_17__SCAN_IN), .ZN(n2487) );
  INV_X1 U32360 ( .A(REG3_REG_17__SCAN_IN), .ZN(n2472) );
  NAND2_X1 U32370 ( .A1(n2473), .A2(n2472), .ZN(n2474) );
  NAND2_X1 U32380 ( .A1(n2487), .A2(n2474), .ZN(n4339) );
  OR2_X1 U32390 ( .A1(n4339), .A2(n2646), .ZN(n2479) );
  INV_X1 U32400 ( .A(REG2_REG_17__SCAN_IN), .ZN(n4340) );
  NAND2_X1 U32410 ( .A1(n2008), .A2(REG0_REG_17__SCAN_IN), .ZN(n2476) );
  NAND2_X1 U32420 ( .A1(n2009), .A2(REG1_REG_17__SCAN_IN), .ZN(n2475) );
  OAI211_X1 U32430 ( .C1(n4340), .C2(n2447), .A(n2476), .B(n2475), .ZN(n2477)
         );
  INV_X1 U32440 ( .A(n2477), .ZN(n2478) );
  OAI21_X1 U32450 ( .B1(n2481), .B2(n2480), .A(IR_REG_31__SCAN_IN), .ZN(n2482)
         );
  XNOR2_X1 U32460 ( .A(n2482), .B(IR_REG_17__SCAN_IN), .ZN(n4082) );
  MUX2_X1 U32470 ( .A(n4082), .B(DATAI_17_), .S(n3722), .Z(n4336) );
  NAND2_X1 U32480 ( .A1(n2487), .A2(n3675), .ZN(n2488) );
  NAND2_X1 U32490 ( .A1(n2501), .A2(n2488), .ZN(n4318) );
  OR2_X1 U32500 ( .A1(n4318), .A2(n2646), .ZN(n2494) );
  INV_X1 U32510 ( .A(n2009), .ZN(n2491) );
  INV_X1 U32520 ( .A(REG1_REG_18__SCAN_IN), .ZN(n4077) );
  NAND2_X1 U32530 ( .A1(n2329), .A2(REG2_REG_18__SCAN_IN), .ZN(n2490) );
  NAND2_X1 U32540 ( .A1(n2008), .A2(REG0_REG_18__SCAN_IN), .ZN(n2489) );
  OAI211_X1 U32550 ( .C1(n2491), .C2(n4077), .A(n2490), .B(n2489), .ZN(n2492)
         );
  INV_X1 U32560 ( .A(n2492), .ZN(n2493) );
  NAND2_X1 U32570 ( .A1(n2495), .A2(IR_REG_31__SCAN_IN), .ZN(n2496) );
  MUX2_X1 U32580 ( .A(IR_REG_31__SCAN_IN), .B(n2496), .S(IR_REG_18__SCAN_IN), 
        .Z(n2497) );
  INV_X1 U32590 ( .A(n2606), .ZN(n2507) );
  MUX2_X1 U32600 ( .A(n4083), .B(DATAI_18_), .S(n3722), .Z(n4315) );
  NAND2_X1 U32610 ( .A1(n4295), .A2(n4315), .ZN(n4289) );
  INV_X1 U32620 ( .A(n4315), .ZN(n3676) );
  NAND2_X1 U32630 ( .A1(n4333), .A2(n3676), .ZN(n4290) );
  NAND2_X1 U32640 ( .A1(n4295), .A2(n3676), .ZN(n2498) );
  NAND2_X1 U32650 ( .A1(n4321), .A2(n2498), .ZN(n4286) );
  NAND2_X1 U32660 ( .A1(n2501), .A2(n2500), .ZN(n2502) );
  NAND2_X1 U32670 ( .A1(n2514), .A2(n2502), .ZN(n4303) );
  INV_X1 U32680 ( .A(REG2_REG_19__SCAN_IN), .ZN(n4304) );
  NAND2_X1 U32690 ( .A1(n2008), .A2(REG0_REG_19__SCAN_IN), .ZN(n2504) );
  NAND2_X1 U32700 ( .A1(n2009), .A2(REG1_REG_19__SCAN_IN), .ZN(n2503) );
  OAI211_X1 U32710 ( .C1(n4304), .C2(n2447), .A(n2504), .B(n2503), .ZN(n2505)
         );
  INV_X1 U32720 ( .A(n2505), .ZN(n2506) );
  INV_X1 U32730 ( .A(n2510), .ZN(n2508) );
  NAND2_X1 U32740 ( .A1(n2508), .A2(IR_REG_19__SCAN_IN), .ZN(n2511) );
  MUX2_X1 U32750 ( .A(n4611), .B(DATAI_19_), .S(n3722), .Z(n3614) );
  NAND2_X1 U32760 ( .A1(n4271), .A2(n3614), .ZN(n2512) );
  NAND2_X1 U32770 ( .A1(n4286), .A2(n2512), .ZN(n4179) );
  INV_X1 U32780 ( .A(n4271), .ZN(n4311) );
  NAND2_X1 U32790 ( .A1(n4311), .A2(n4301), .ZN(n3479) );
  INV_X1 U32800 ( .A(n2514), .ZN(n2513) );
  NAND2_X1 U32810 ( .A1(n2514), .A2(n2058), .ZN(n2515) );
  AND2_X1 U32820 ( .A1(n2522), .A2(n2515), .ZN(n4281) );
  NAND2_X1 U32830 ( .A1(n4281), .A2(n2331), .ZN(n2521) );
  INV_X1 U32840 ( .A(REG2_REG_20__SCAN_IN), .ZN(n2518) );
  NAND2_X1 U32850 ( .A1(n2008), .A2(REG0_REG_20__SCAN_IN), .ZN(n2517) );
  NAND2_X1 U32860 ( .A1(n2009), .A2(REG1_REG_20__SCAN_IN), .ZN(n2516) );
  OAI211_X1 U32870 ( .C1(n2518), .C2(n2447), .A(n2517), .B(n2516), .ZN(n2519)
         );
  INV_X1 U32880 ( .A(n2519), .ZN(n2520) );
  OR2_X1 U32890 ( .A1(n4297), .A2(n4270), .ZN(n3745) );
  INV_X1 U32900 ( .A(REG3_REG_21__SCAN_IN), .ZN(n3978) );
  NAND2_X1 U32910 ( .A1(n2522), .A2(n3978), .ZN(n2523) );
  NAND2_X1 U32920 ( .A1(n2530), .A2(n2523), .ZN(n4260) );
  OR2_X1 U32930 ( .A1(n4260), .A2(n2646), .ZN(n2528) );
  INV_X1 U32940 ( .A(REG2_REG_21__SCAN_IN), .ZN(n4259) );
  NAND2_X1 U32950 ( .A1(n2008), .A2(REG0_REG_21__SCAN_IN), .ZN(n2525) );
  NAND2_X1 U32960 ( .A1(n2009), .A2(REG1_REG_21__SCAN_IN), .ZN(n2524) );
  OAI211_X1 U32970 ( .C1(n4259), .C2(n2447), .A(n2525), .B(n2524), .ZN(n2526)
         );
  INV_X1 U32980 ( .A(n2526), .ZN(n2527) );
  INV_X1 U32990 ( .A(n4257), .ZN(n4251) );
  NAND2_X1 U33000 ( .A1(n4273), .A2(n4251), .ZN(n3481) );
  NAND2_X1 U33010 ( .A1(n2530), .A2(n2529), .ZN(n2531) );
  AND2_X1 U33020 ( .A1(n2539), .A2(n2531), .ZN(n3492) );
  NAND2_X1 U33030 ( .A1(n3492), .A2(n2331), .ZN(n2536) );
  INV_X1 U33040 ( .A(REG2_REG_22__SCAN_IN), .ZN(n3493) );
  NAND2_X1 U33050 ( .A1(n2008), .A2(REG0_REG_22__SCAN_IN), .ZN(n2533) );
  NAND2_X1 U33060 ( .A1(n2009), .A2(REG1_REG_22__SCAN_IN), .ZN(n2532) );
  OAI211_X1 U33070 ( .C1(n3493), .C2(n2447), .A(n2533), .B(n2532), .ZN(n2534)
         );
  INV_X1 U33080 ( .A(n2534), .ZN(n2535) );
  NAND2_X1 U33090 ( .A1(n4254), .A2(n2702), .ZN(n2640) );
  NAND2_X1 U33100 ( .A1(n4236), .A2(n3491), .ZN(n4230) );
  NAND2_X1 U33110 ( .A1(n4254), .A2(n3491), .ZN(n2564) );
  INV_X1 U33120 ( .A(n2539), .ZN(n2537) );
  NAND2_X1 U33130 ( .A1(n2537), .A2(REG3_REG_23__SCAN_IN), .ZN(n2553) );
  INV_X1 U33140 ( .A(REG3_REG_23__SCAN_IN), .ZN(n2538) );
  NAND2_X1 U33150 ( .A1(n2539), .A2(n2538), .ZN(n2540) );
  NAND2_X1 U33160 ( .A1(n2553), .A2(n2540), .ZN(n4244) );
  OR2_X1 U33170 ( .A1(n4244), .A2(n2646), .ZN(n2545) );
  INV_X1 U33180 ( .A(REG2_REG_23__SCAN_IN), .ZN(n4243) );
  NAND2_X1 U33190 ( .A1(n2008), .A2(REG0_REG_23__SCAN_IN), .ZN(n2542) );
  NAND2_X1 U33200 ( .A1(n2009), .A2(REG1_REG_23__SCAN_IN), .ZN(n2541) );
  OAI211_X1 U33210 ( .C1(n4243), .C2(n2447), .A(n2542), .B(n2541), .ZN(n2543)
         );
  INV_X1 U33220 ( .A(n2543), .ZN(n2544) );
  NAND2_X1 U33230 ( .A1(n4215), .A2(n4241), .ZN(n2563) );
  AND2_X1 U33240 ( .A1(n4225), .A2(n2563), .ZN(n2569) );
  AND2_X1 U33250 ( .A1(n3479), .A2(n2569), .ZN(n4178) );
  NAND2_X1 U33260 ( .A1(n2555), .A2(n3967), .ZN(n2546) );
  NAND2_X1 U33270 ( .A1(n4200), .A2(n2331), .ZN(n2552) );
  INV_X1 U33280 ( .A(REG2_REG_25__SCAN_IN), .ZN(n2549) );
  NAND2_X1 U33290 ( .A1(n2008), .A2(REG0_REG_25__SCAN_IN), .ZN(n2548) );
  NAND2_X1 U33300 ( .A1(n2009), .A2(REG1_REG_25__SCAN_IN), .ZN(n2547) );
  OAI211_X1 U33310 ( .C1(n2549), .C2(n2447), .A(n2548), .B(n2547), .ZN(n2550)
         );
  INV_X1 U33320 ( .A(n2550), .ZN(n2551) );
  NAND2_X1 U33330 ( .A1(n2553), .A2(n3645), .ZN(n2554) );
  NAND2_X1 U33340 ( .A1(n4220), .A2(n2331), .ZN(n2560) );
  INV_X1 U33350 ( .A(REG1_REG_24__SCAN_IN), .ZN(n4485) );
  NAND2_X1 U33360 ( .A1(n2329), .A2(REG2_REG_24__SCAN_IN), .ZN(n2557) );
  NAND2_X1 U33370 ( .A1(n2008), .A2(REG0_REG_24__SCAN_IN), .ZN(n2556) );
  OAI211_X1 U33380 ( .C1(n2491), .C2(n4485), .A(n2557), .B(n2556), .ZN(n2558)
         );
  INV_X1 U33390 ( .A(n2558), .ZN(n2559) );
  NAND2_X1 U33400 ( .A1(n4191), .A2(n4214), .ZN(n4183) );
  AND2_X1 U33410 ( .A1(n2231), .A2(n4183), .ZN(n2562) );
  AND2_X1 U33420 ( .A1(n4178), .A2(n2562), .ZN(n2561) );
  NAND2_X1 U33430 ( .A1(n4179), .A2(n2561), .ZN(n4157) );
  INV_X1 U33440 ( .A(n4241), .ZN(n2643) );
  NAND2_X1 U33450 ( .A1(n3874), .A2(n2643), .ZN(n2568) );
  INV_X1 U33460 ( .A(n2563), .ZN(n2566) );
  NAND2_X1 U33470 ( .A1(n3663), .A2(n4257), .ZN(n3480) );
  OR2_X1 U33480 ( .A1(n2566), .A2(n4227), .ZN(n2567) );
  AND2_X1 U33490 ( .A1(n2568), .A2(n2567), .ZN(n4205) );
  AND2_X1 U33500 ( .A1(n4205), .A2(n2223), .ZN(n4182) );
  INV_X1 U33510 ( .A(n2569), .ZN(n2570) );
  NAND2_X1 U33520 ( .A1(n4297), .A2(n4270), .ZN(n3744) );
  OR2_X1 U3353 ( .A1(n2570), .A2(n3744), .ZN(n4180) );
  INV_X1 U33540 ( .A(n2573), .ZN(n2571) );
  NAND2_X1 U3355 ( .A1(n2571), .A2(REG3_REG_26__SCAN_IN), .ZN(n2584) );
  INV_X1 U3356 ( .A(REG3_REG_26__SCAN_IN), .ZN(n2572) );
  NAND2_X1 U3357 ( .A1(n2573), .A2(n2572), .ZN(n2574) );
  NAND2_X1 U3358 ( .A1(n2584), .A2(n2574), .ZN(n4169) );
  INV_X1 U3359 ( .A(REG2_REG_26__SCAN_IN), .ZN(n4168) );
  NAND2_X1 U3360 ( .A1(n2008), .A2(REG0_REG_26__SCAN_IN), .ZN(n2576) );
  NAND2_X1 U3361 ( .A1(n2009), .A2(REG1_REG_26__SCAN_IN), .ZN(n2575) );
  OAI211_X1 U3362 ( .C1(n4168), .C2(n2447), .A(n2576), .B(n2575), .ZN(n2577)
         );
  INV_X1 U3363 ( .A(n2577), .ZN(n2578) );
  OR2_X1 U3364 ( .A1(n4142), .A2(n4172), .ZN(n2580) );
  NAND2_X1 U3365 ( .A1(n4142), .A2(n4172), .ZN(n2582) );
  NAND2_X1 U3366 ( .A1(n2584), .A2(n2583), .ZN(n2585) );
  NAND2_X1 U3367 ( .A1(n4150), .A2(n2331), .ZN(n2591) );
  INV_X1 U3368 ( .A(REG2_REG_27__SCAN_IN), .ZN(n2588) );
  NAND2_X1 U3369 ( .A1(n2008), .A2(REG0_REG_27__SCAN_IN), .ZN(n2587) );
  NAND2_X1 U3370 ( .A1(n2009), .A2(REG1_REG_27__SCAN_IN), .ZN(n2586) );
  OAI211_X1 U3371 ( .C1(n2588), .C2(n2447), .A(n2587), .B(n2586), .ZN(n2589)
         );
  INV_X1 U3372 ( .A(n2589), .ZN(n2590) );
  NOR2_X1 U3373 ( .A1(n4165), .A2(n3845), .ZN(n2592) );
  INV_X1 U3374 ( .A(n2595), .ZN(n2593) );
  NAND2_X1 U3375 ( .A1(n2593), .A2(REG3_REG_28__SCAN_IN), .ZN(n4125) );
  INV_X1 U3376 ( .A(REG3_REG_28__SCAN_IN), .ZN(n2594) );
  NAND2_X1 U3377 ( .A1(n2595), .A2(n2594), .ZN(n2596) );
  NAND2_X1 U3378 ( .A1(n4125), .A2(n2596), .ZN(n4132) );
  INV_X1 U3379 ( .A(REG2_REG_28__SCAN_IN), .ZN(n4131) );
  NAND2_X1 U3380 ( .A1(n2008), .A2(REG0_REG_28__SCAN_IN), .ZN(n2598) );
  NAND2_X1 U3381 ( .A1(n2009), .A2(REG1_REG_28__SCAN_IN), .ZN(n2597) );
  OAI211_X1 U3382 ( .C1(n4131), .C2(n2447), .A(n2598), .B(n2597), .ZN(n2599)
         );
  INV_X1 U3383 ( .A(n2599), .ZN(n2600) );
  NAND2_X1 U3384 ( .A1(n4145), .A2(n4110), .ZN(n4115) );
  NAND2_X1 U3385 ( .A1(n4111), .A2(n3535), .ZN(n4114) );
  NAND2_X1 U3386 ( .A1(n2663), .A2(IR_REG_31__SCAN_IN), .ZN(n2607) );
  NAND2_X1 U3387 ( .A1(n2012), .A2(IR_REG_31__SCAN_IN), .ZN(n2609) );
  XNOR2_X1 U3388 ( .A(n3131), .B(n3868), .ZN(n2610) );
  NAND2_X1 U3389 ( .A1(n2698), .A2(n2720), .ZN(n3784) );
  NAND2_X1 U3390 ( .A1(n3784), .A2(n3787), .ZN(n3071) );
  INV_X1 U3391 ( .A(n3071), .ZN(n2612) );
  NAND2_X1 U3392 ( .A1(n3047), .A2(n3221), .ZN(n3025) );
  INV_X1 U3393 ( .A(n3025), .ZN(n3786) );
  NAND2_X1 U3394 ( .A1(n2612), .A2(n3786), .ZN(n3077) );
  NAND2_X1 U3395 ( .A1(n3077), .A2(n3787), .ZN(n2613) );
  NAND2_X1 U3396 ( .A1(n2613), .A2(n3750), .ZN(n3080) );
  NAND2_X1 U3397 ( .A1(n3080), .A2(n3788), .ZN(n3181) );
  NAND2_X1 U3398 ( .A1(n3187), .A2(n3168), .ZN(n3793) );
  NAND2_X1 U3399 ( .A1(n3106), .A2(n4016), .ZN(n3790) );
  NAND2_X1 U3400 ( .A1(n3181), .A2(n3754), .ZN(n3180) );
  NAND2_X1 U3401 ( .A1(n3180), .A2(n3793), .ZN(n3112) );
  INV_X1 U3402 ( .A(n3794), .ZN(n2614) );
  AND2_X1 U3403 ( .A1(n2615), .A2(n2616), .ZN(n3797) );
  NAND2_X1 U3404 ( .A1(n3247), .A2(n3277), .ZN(n3809) );
  INV_X1 U3405 ( .A(n3282), .ZN(n3285) );
  NAND2_X1 U3406 ( .A1(n3285), .A2(n4015), .ZN(n3810) );
  INV_X1 U3407 ( .A(n4015), .ZN(n2617) );
  NAND2_X1 U3408 ( .A1(n3282), .A2(n2617), .ZN(n3799) );
  INV_X1 U3409 ( .A(n2618), .ZN(n2619) );
  NAND2_X1 U3410 ( .A1(n3298), .A2(n3387), .ZN(n3805) );
  NAND2_X1 U3411 ( .A1(n3291), .A2(n3805), .ZN(n2620) );
  NAND2_X1 U3412 ( .A1(n2787), .A2(n3319), .ZN(n3803) );
  AND2_X1 U3413 ( .A1(n3382), .A2(n2409), .ZN(n3383) );
  NAND2_X1 U3414 ( .A1(n3389), .A2(n3396), .ZN(n3806) );
  NAND2_X1 U3415 ( .A1(n3404), .A2(n4014), .ZN(n3817) );
  NAND2_X1 U3416 ( .A1(n3395), .A2(n3817), .ZN(n2621) );
  NAND2_X1 U3417 ( .A1(n3398), .A2(n3386), .ZN(n3816) );
  NAND2_X1 U3418 ( .A1(n2621), .A2(n3816), .ZN(n3411) );
  NAND2_X1 U3419 ( .A1(n4446), .A2(n4012), .ZN(n4409) );
  NAND2_X1 U3420 ( .A1(n3746), .A2(n4387), .ZN(n2622) );
  NAND2_X1 U3421 ( .A1(n4409), .A2(n2622), .ZN(n2624) );
  INV_X1 U3422 ( .A(n4408), .ZN(n2623) );
  NOR2_X1 U3423 ( .A1(n2624), .A2(n2623), .ZN(n3818) );
  NAND2_X1 U3424 ( .A1(n3411), .A2(n3818), .ZN(n2628) );
  INV_X1 U3425 ( .A(n2624), .ZN(n2627) );
  NAND2_X1 U3426 ( .A1(n4440), .A2(n4413), .ZN(n4411) );
  NAND2_X1 U3427 ( .A1(n4406), .A2(n4411), .ZN(n2626) );
  NOR2_X1 U3428 ( .A1(n3746), .A2(n4387), .ZN(n2625) );
  AOI21_X1 U3429 ( .B1(n2627), .B2(n2626), .A(n2625), .ZN(n3826) );
  NAND2_X1 U3430 ( .A1(n2628), .A2(n3826), .ZN(n3709) );
  NAND2_X1 U3431 ( .A1(n3709), .A2(n2190), .ZN(n4385) );
  INV_X1 U3432 ( .A(n4389), .ZN(n2629) );
  NAND2_X1 U3433 ( .A1(n2629), .A2(n4373), .ZN(n3712) );
  NAND2_X1 U3434 ( .A1(n4389), .A2(n4376), .ZN(n3711) );
  NAND2_X1 U3435 ( .A1(n3712), .A2(n3711), .ZN(n4374) );
  INV_X1 U3436 ( .A(n4368), .ZN(n2630) );
  NOR2_X1 U3437 ( .A1(n4374), .A2(n2630), .ZN(n2631) );
  NAND2_X1 U3438 ( .A1(n4385), .A2(n2631), .ZN(n2632) );
  NAND2_X1 U3439 ( .A1(n2632), .A2(n3711), .ZN(n4346) );
  INV_X1 U3440 ( .A(n4353), .ZN(n3748) );
  NAND2_X1 U3441 ( .A1(n4271), .A2(n4301), .ZN(n2633) );
  NAND2_X1 U3442 ( .A1(n2633), .A2(n4290), .ZN(n2634) );
  AND2_X1 U3443 ( .A1(n4347), .A2(n2483), .ZN(n4288) );
  OR2_X1 U3444 ( .A1(n2634), .A2(n4288), .ZN(n3831) );
  INV_X1 U3445 ( .A(n2634), .ZN(n2637) );
  NAND2_X1 U3446 ( .A1(n2484), .A2(n4336), .ZN(n4287) );
  NAND2_X1 U3447 ( .A1(n4289), .A2(n4287), .ZN(n2636) );
  NOR2_X1 U3448 ( .A1(n4271), .A2(n4301), .ZN(n2635) );
  AOI21_X1 U3449 ( .B1(n2637), .B2(n2636), .A(n2635), .ZN(n4266) );
  OR2_X1 U3450 ( .A1(n4297), .A2(n4280), .ZN(n2638) );
  AND2_X1 U3451 ( .A1(n4266), .A2(n2638), .ZN(n3714) );
  NAND2_X1 U3452 ( .A1(n4297), .A2(n4280), .ZN(n3835) );
  NAND2_X1 U3453 ( .A1(n2639), .A2(n3835), .ZN(n3486) );
  NAND2_X1 U3454 ( .A1(n4273), .A2(n4257), .ZN(n3743) );
  AND2_X1 U3455 ( .A1(n4230), .A2(n3743), .ZN(n3839) );
  NAND2_X1 U3456 ( .A1(n3486), .A2(n3839), .ZN(n2642) );
  NAND2_X1 U3457 ( .A1(n3874), .A2(n4241), .ZN(n3740) );
  NAND2_X1 U34580 ( .A1(n3740), .A2(n2640), .ZN(n3838) );
  AND2_X1 U34590 ( .A1(n3663), .A2(n4251), .ZN(n3742) );
  AND2_X1 U3460 ( .A1(n4230), .A2(n3742), .ZN(n2641) );
  NOR2_X1 U3461 ( .A1(n3838), .A2(n2641), .ZN(n3716) );
  NAND2_X1 U3462 ( .A1(n4215), .A2(n2643), .ZN(n3741) );
  NOR2_X1 U3463 ( .A1(n4238), .A2(n4214), .ZN(n3738) );
  NAND2_X1 U3464 ( .A1(n4217), .A2(n4198), .ZN(n3778) );
  NAND2_X1 U3465 ( .A1(n4238), .A2(n4214), .ZN(n4187) );
  AND2_X1 U3466 ( .A1(n3778), .A2(n4187), .ZN(n3841) );
  NAND2_X1 U34670 ( .A1(n4186), .A2(n3841), .ZN(n4160) );
  NAND2_X1 U3468 ( .A1(n4142), .A2(n3686), .ZN(n3737) );
  OR2_X1 U34690 ( .A1(n4217), .A2(n4198), .ZN(n4159) );
  AND2_X1 U3470 ( .A1(n3737), .A2(n4159), .ZN(n3851) );
  AND2_X1 U34710 ( .A1(n4193), .A2(n4172), .ZN(n3731) );
  XNOR2_X1 U3472 ( .A(n4165), .B(n3845), .ZN(n4140) );
  INV_X1 U34730 ( .A(n3783), .ZN(n4108) );
  NAND2_X1 U3474 ( .A1(n3868), .A2(n4611), .ZN(n2645) );
  INV_X1 U34750 ( .A(n2611), .ZN(n2962) );
  NAND2_X1 U3476 ( .A1(n2644), .A2(n2962), .ZN(n3863) );
  OR2_X1 U34770 ( .A1(n4125), .A2(n2646), .ZN(n2651) );
  INV_X1 U3478 ( .A(REG0_REG_29__SCAN_IN), .ZN(n3934) );
  NAND2_X1 U34790 ( .A1(n2329), .A2(REG2_REG_29__SCAN_IN), .ZN(n2648) );
  NAND2_X1 U3480 ( .A1(n2009), .A2(REG1_REG_29__SCAN_IN), .ZN(n2647) );
  OAI211_X1 U34810 ( .C1(n2301), .C2(n3934), .A(n2648), .B(n2647), .ZN(n2649)
         );
  INV_X1 U3482 ( .A(n2649), .ZN(n2650) );
  NAND2_X1 U34830 ( .A1(n2651), .A2(n2650), .ZN(n3873) );
  NAND2_X1 U3484 ( .A1(n2652), .A2(IR_REG_31__SCAN_IN), .ZN(n2653) );
  MUX2_X1 U34850 ( .A(IR_REG_31__SCAN_IN), .B(n2653), .S(IR_REG_28__SCAN_IN), 
        .Z(n2654) );
  INV_X1 U3486 ( .A(n4609), .ZN(n2912) );
  NAND2_X1 U34870 ( .A1(n3873), .A2(n4388), .ZN(n2657) );
  NOR2_X1 U3488 ( .A1(n3535), .A2(n4391), .ZN(n2655) );
  AOI21_X1 U34890 ( .B1(n4165), .B2(n4386), .A(n2655), .ZN(n2656) );
  NAND2_X1 U3490 ( .A1(n2660), .A2(IR_REG_31__SCAN_IN), .ZN(n2661) );
  MUX2_X1 U34910 ( .A(IR_REG_31__SCAN_IN), .B(n2661), .S(IR_REG_25__SCAN_IN), 
        .Z(n2662) );
  NAND2_X1 U3492 ( .A1(n2976), .A2(B_REG_SCAN_IN), .ZN(n2671) );
  INV_X1 U34930 ( .A(n2663), .ZN(n2669) );
  MUX2_X1 U3494 ( .A(n2671), .B(B_REG_SCAN_IN), .S(n2677), .Z(n2675) );
  NAND2_X1 U34950 ( .A1(n2659), .A2(IR_REG_31__SCAN_IN), .ZN(n2672) );
  MUX2_X1 U3496 ( .A(IR_REG_31__SCAN_IN), .B(n2672), .S(IR_REG_26__SCAN_IN), 
        .Z(n2673) );
  NAND2_X1 U34970 ( .A1(n2674), .A2(n2673), .ZN(n2676) );
  NAND2_X1 U3498 ( .A1(n2676), .A2(n2976), .ZN(n2876) );
  NAND2_X1 U34990 ( .A1(n3125), .A2(n2876), .ZN(n2694) );
  NAND2_X1 U3500 ( .A1(n4712), .A2(n3766), .ZN(n2901) );
  NAND2_X1 U35010 ( .A1(n2611), .A2(n4088), .ZN(n2879) );
  NAND2_X1 U3502 ( .A1(n2917), .A2(n2879), .ZN(n3122) );
  NAND2_X1 U35030 ( .A1(n2901), .A2(n3122), .ZN(n2682) );
  OAI211_X1 U3504 ( .C1(n2012), .C2(IR_REG_22__SCAN_IN), .A(IR_REG_31__SCAN_IN), .B(IR_REG_23__SCAN_IN), .ZN(n2680) );
  NOR2_X1 U35050 ( .A1(n2682), .A2(n3123), .ZN(n2693) );
  NOR4_X1 U35060 ( .A1(D_REG_18__SCAN_IN), .A2(D_REG_19__SCAN_IN), .A3(
        D_REG_21__SCAN_IN), .A4(D_REG_22__SCAN_IN), .ZN(n2686) );
  NOR4_X1 U35070 ( .A1(D_REG_13__SCAN_IN), .A2(D_REG_17__SCAN_IN), .A3(
        D_REG_14__SCAN_IN), .A4(D_REG_16__SCAN_IN), .ZN(n2685) );
  NOR4_X1 U35080 ( .A1(D_REG_27__SCAN_IN), .A2(D_REG_28__SCAN_IN), .A3(
        D_REG_29__SCAN_IN), .A4(D_REG_30__SCAN_IN), .ZN(n2684) );
  NOR4_X1 U35090 ( .A1(D_REG_25__SCAN_IN), .A2(D_REG_23__SCAN_IN), .A3(
        D_REG_24__SCAN_IN), .A4(D_REG_26__SCAN_IN), .ZN(n2683) );
  NAND4_X1 U35100 ( .A1(n2686), .A2(n2685), .A3(n2684), .A4(n2683), .ZN(n2691)
         );
  NOR3_X1 U35110 ( .A1(D_REG_10__SCAN_IN), .A2(D_REG_15__SCAN_IN), .A3(
        D_REG_20__SCAN_IN), .ZN(n3880) );
  NOR3_X1 U35120 ( .A1(D_REG_2__SCAN_IN), .A2(D_REG_3__SCAN_IN), .A3(
        D_REG_31__SCAN_IN), .ZN(n2689) );
  NOR4_X1 U35130 ( .A1(D_REG_7__SCAN_IN), .A2(D_REG_9__SCAN_IN), .A3(
        D_REG_11__SCAN_IN), .A4(D_REG_12__SCAN_IN), .ZN(n2688) );
  NOR4_X1 U35140 ( .A1(D_REG_4__SCAN_IN), .A2(D_REG_5__SCAN_IN), .A3(
        D_REG_8__SCAN_IN), .A4(D_REG_6__SCAN_IN), .ZN(n2687) );
  NAND4_X1 U35150 ( .A1(n3880), .A2(n2689), .A3(n2688), .A4(n2687), .ZN(n2690)
         );
  NOR2_X1 U35160 ( .A1(n2691), .A2(n2690), .ZN(n2692) );
  INV_X1 U35170 ( .A(n2677), .ZN(n2695) );
  NAND2_X1 U35180 ( .A1(n2695), .A2(n2676), .ZN(n2696) );
  NAND2_X1 U35190 ( .A1(n3119), .A2(n3120), .ZN(n3246) );
  NAND2_X1 U35200 ( .A1(n2615), .A2(n3285), .ZN(n3196) );
  NAND2_X1 U35210 ( .A1(n2700), .A2(n2699), .ZN(n2701) );
  NAND2_X1 U35220 ( .A1(n4208), .A2(n4214), .ZN(n4196) );
  INV_X1 U35230 ( .A(n2703), .ZN(n2704) );
  NAND2_X1 U35240 ( .A1(n2704), .A2(n4110), .ZN(n2705) );
  NAND2_X1 U35250 ( .A1(n2033), .A2(n2705), .ZN(n4133) );
  INV_X1 U35260 ( .A(n4133), .ZN(n2708) );
  NAND2_X1 U35270 ( .A1(n2712), .A2(REG1_REG_28__SCAN_IN), .ZN(n2709) );
  INV_X1 U35280 ( .A(REG0_REG_28__SCAN_IN), .ZN(n2714) );
  OAI21_X1 U35290 ( .B1(n2718), .B2(n4729), .A(n2717), .ZN(U3514) );
  INV_X1 U35300 ( .A(n3131), .ZN(n2719) );
  AND2_X2 U35310 ( .A1(n2890), .A2(n2719), .ZN(n2741) );
  NAND2_X1 U35320 ( .A1(n2720), .A2(n2741), .ZN(n2722) );
  INV_X2 U35330 ( .A(n2729), .ZN(n2726) );
  NAND2_X1 U35340 ( .A1(n3223), .A2(n2726), .ZN(n2721) );
  NAND2_X1 U35350 ( .A1(n2722), .A2(n2721), .ZN(n2724) );
  AND2_X4 U35360 ( .A1(n2726), .A2(n2725), .ZN(n2754) );
  NAND2_X1 U35370 ( .A1(n2754), .A2(n3082), .ZN(n2728) );
  NAND2_X1 U35380 ( .A1(n3223), .A2(n3560), .ZN(n2727) );
  NAND2_X1 U35390 ( .A1(n2728), .A2(n2727), .ZN(n2738) );
  XNOR2_X1 U35400 ( .A(n2739), .B(n2738), .ZN(n3050) );
  INV_X1 U35410 ( .A(n3050), .ZN(n2737) );
  NAND2_X1 U35420 ( .A1(n3221), .A2(n2726), .ZN(n2731) );
  NAND2_X1 U35430 ( .A1(n3024), .A2(n2741), .ZN(n2730) );
  INV_X1 U35440 ( .A(REG1_REG_0__SCAN_IN), .ZN(n4023) );
  OR2_X1 U35450 ( .A1(n2890), .A2(n4023), .ZN(n2732) );
  NAND2_X1 U35460 ( .A1(n3221), .A2(n2741), .ZN(n2734) );
  NAND2_X1 U35470 ( .A1(n2754), .A2(n3024), .ZN(n2733) );
  OAI211_X1 U35480 ( .C1(n2890), .C2(n2300), .A(n2734), .B(n2733), .ZN(n2911)
         );
  AOI22_X1 U35490 ( .A1(n2910), .A2(n2911), .B1(n2735), .B2(n3533), .ZN(n3049)
         );
  INV_X1 U35500 ( .A(n3049), .ZN(n2736) );
  NAND2_X1 U35510 ( .A1(n2737), .A2(n2736), .ZN(n3051) );
  NAND2_X1 U35520 ( .A1(n2739), .A2(n2738), .ZN(n2740) );
  NAND2_X1 U35530 ( .A1(n2742), .A2(n2726), .ZN(n2743) );
  OAI21_X1 U35540 ( .B1(n2315), .B2(n3556), .A(n2743), .ZN(n2744) );
  XNOR2_X1 U35550 ( .A(n2744), .B(n3561), .ZN(n2748) );
  AOI22_X1 U35560 ( .A1(n2745), .A2(n2754), .B1(n2742), .B2(n3560), .ZN(n2749)
         );
  XNOR2_X1 U35570 ( .A(n2748), .B(n2749), .ZN(n3095) );
  NAND2_X1 U35580 ( .A1(n3094), .A2(n3095), .ZN(n3093) );
  NAND2_X1 U35590 ( .A1(n3165), .A2(n2726), .ZN(n2746) );
  OAI21_X1 U35600 ( .B1(n3502), .B2(n3556), .A(n2746), .ZN(n2747) );
  XNOR2_X1 U35610 ( .A(n2747), .B(n3533), .ZN(n2765) );
  AOI22_X1 U35620 ( .A1(n2985), .A2(n2754), .B1(n3165), .B2(n3560), .ZN(n2766)
         );
  XNOR2_X1 U35630 ( .A(n2765), .B(n2766), .ZN(n2762) );
  INV_X1 U35640 ( .A(n2748), .ZN(n2750) );
  NAND2_X1 U35650 ( .A1(n2750), .A2(n2749), .ZN(n3103) );
  NAND2_X1 U35660 ( .A1(n3187), .A2(n2726), .ZN(n2752) );
  NAND2_X1 U35670 ( .A1(n2741), .A2(n4016), .ZN(n2751) );
  NAND2_X1 U35680 ( .A1(n2752), .A2(n2751), .ZN(n2753) );
  NAND2_X1 U35690 ( .A1(n2754), .A2(n4016), .ZN(n2756) );
  NAND2_X1 U35700 ( .A1(n3187), .A2(n2741), .ZN(n2755) );
  NAND2_X1 U35710 ( .A1(n2756), .A2(n2755), .ZN(n2758) );
  INV_X1 U35720 ( .A(n2758), .ZN(n2757) );
  NAND2_X1 U35730 ( .A1(n2759), .A2(n2757), .ZN(n2760) );
  AND2_X1 U35740 ( .A1(n3103), .A2(n2760), .ZN(n3169) );
  NAND3_X1 U35750 ( .A1(n3093), .A2(n2763), .A3(n3169), .ZN(n3172) );
  XNOR2_X1 U35760 ( .A(n2759), .B(n2758), .ZN(n3102) );
  INV_X1 U35770 ( .A(n3102), .ZN(n2761) );
  NAND2_X1 U35780 ( .A1(n2761), .A2(n2760), .ZN(n3171) );
  INV_X1 U35790 ( .A(n3171), .ZN(n2764) );
  NAND2_X1 U35800 ( .A1(n2764), .A2(n2763), .ZN(n3173) );
  INV_X1 U35810 ( .A(n2765), .ZN(n2768) );
  INV_X1 U3582 ( .A(n2766), .ZN(n2767) );
  NAND2_X1 U3583 ( .A1(n2768), .A2(n2767), .ZN(n2769) );
  NAND2_X1 U3584 ( .A1(n3172), .A2(n2770), .ZN(n3499) );
  OAI22_X1 U3585 ( .A1(n2615), .A2(n3554), .B1(n3277), .B2(n3556), .ZN(n2771)
         );
  XNOR2_X1 U3586 ( .A(n2771), .B(n3533), .ZN(n2772) );
  OAI22_X1 U3587 ( .A1(n2615), .A2(n3556), .B1(n3277), .B2(n3557), .ZN(n2773)
         );
  XNOR2_X1 U3588 ( .A(n2772), .B(n2773), .ZN(n3501) );
  NAND2_X1 U3589 ( .A1(n3499), .A2(n3501), .ZN(n3500) );
  INV_X1 U3590 ( .A(n2772), .ZN(n2774) );
  NAND2_X1 U3591 ( .A1(n2774), .A2(n2773), .ZN(n2775) );
  NAND2_X1 U3592 ( .A1(n3282), .A2(n3560), .ZN(n2777) );
  NAND2_X1 U3593 ( .A1(n2754), .A2(n4015), .ZN(n2776) );
  NAND2_X1 U3594 ( .A1(n2777), .A2(n2776), .ZN(n3136) );
  NAND2_X1 U3595 ( .A1(n3282), .A2(n2726), .ZN(n2779) );
  NAND2_X1 U3596 ( .A1(n4015), .A2(n3560), .ZN(n2778) );
  NAND2_X1 U3597 ( .A1(n2779), .A2(n2778), .ZN(n2780) );
  XNOR2_X1 U3598 ( .A(n2780), .B(n3561), .ZN(n3135) );
  NAND2_X1 U3599 ( .A1(n3213), .A2(n2726), .ZN(n2781) );
  OAI21_X1 U3600 ( .B1(n3292), .B2(n3556), .A(n2781), .ZN(n2782) );
  XNOR2_X1 U3601 ( .A(n2782), .B(n3561), .ZN(n2785) );
  AOI22_X1 U3602 ( .A1(n2367), .A2(n2754), .B1(n3213), .B2(n3560), .ZN(n2783)
         );
  XNOR2_X1 U3603 ( .A(n2785), .B(n2783), .ZN(n3212) );
  INV_X1 U3604 ( .A(n2783), .ZN(n2784) );
  INV_X1 U3605 ( .A(n3256), .ZN(n2803) );
  OAI22_X1 U3606 ( .A1(n3554), .A2(n2787), .B1(n3387), .B2(n3556), .ZN(n2786)
         );
  XNOR2_X1 U3607 ( .A(n2786), .B(n3561), .ZN(n2800) );
  OAI22_X1 U3608 ( .A1(n3556), .A2(n2787), .B1(n3387), .B2(n3557), .ZN(n2799)
         );
  AND2_X1 U3609 ( .A1(n2800), .A2(n2799), .ZN(n3316) );
  OAI22_X1 U3610 ( .A1(n3396), .A2(n3556), .B1(n3554), .B2(n3382), .ZN(n2788)
         );
  XNOR2_X1 U3611 ( .A(n2788), .B(n3533), .ZN(n2791) );
  INV_X1 U3612 ( .A(n2791), .ZN(n2789) );
  OAI22_X1 U3613 ( .A1(n3382), .A2(n3556), .B1(n3396), .B2(n3557), .ZN(n2790)
         );
  OR2_X1 U3614 ( .A1(n2789), .A2(n2790), .ZN(n2801) );
  INV_X1 U3615 ( .A(n2801), .ZN(n2792) );
  XNOR2_X1 U3616 ( .A(n2791), .B(n2790), .ZN(n3315) );
  OR2_X1 U3617 ( .A1(n2792), .A2(n3315), .ZN(n3370) );
  INV_X1 U3618 ( .A(n3370), .ZN(n2795) );
  OAI22_X1 U3619 ( .A1(n3404), .A2(n3554), .B1(n3386), .B2(n3556), .ZN(n2793)
         );
  XNOR2_X1 U3620 ( .A(n2793), .B(n3561), .ZN(n2797) );
  OAI22_X1 U3621 ( .A1(n3404), .A2(n3556), .B1(n3386), .B2(n3557), .ZN(n2796)
         );
  XNOR2_X1 U3622 ( .A(n2797), .B(n2796), .ZN(n3377) );
  NAND2_X1 U3623 ( .A1(n2797), .A2(n2796), .ZN(n2798) );
  OR2_X1 U3624 ( .A1(n2800), .A2(n2799), .ZN(n3317) );
  AND2_X1 U3625 ( .A1(n3317), .A2(n2801), .ZN(n3369) );
  AND2_X1 U3626 ( .A1(n3369), .A2(n2794), .ZN(n3372) );
  AOI21_X2 U3627 ( .B1(n2803), .B2(n2226), .A(n2225), .ZN(n3309) );
  NAND2_X1 U3628 ( .A1(n3310), .A2(n3560), .ZN(n2804) );
  OAI21_X1 U3629 ( .B1(n4435), .B2(n3557), .A(n2804), .ZN(n3307) );
  NAND2_X1 U3630 ( .A1(n3310), .A2(n2726), .ZN(n2805) );
  OAI21_X1 U3631 ( .B1(n4435), .B2(n3556), .A(n2805), .ZN(n2806) );
  XNOR2_X1 U3632 ( .A(n2806), .B(n3561), .ZN(n3306) );
  NAND2_X1 U3633 ( .A1(n4440), .A2(n2726), .ZN(n2808) );
  NAND2_X1 U3634 ( .A1(n4012), .A2(n3560), .ZN(n2807) );
  NAND2_X1 U3635 ( .A1(n2808), .A2(n2807), .ZN(n2809) );
  XNOR2_X1 U3636 ( .A(n2809), .B(n3561), .ZN(n2812) );
  NAND2_X1 U3637 ( .A1(n4440), .A2(n3560), .ZN(n2811) );
  NAND2_X1 U3638 ( .A1(n2754), .A2(n4012), .ZN(n2810) );
  NAND2_X1 U3639 ( .A1(n2811), .A2(n2810), .ZN(n2813) );
  AND2_X1 U3640 ( .A1(n2812), .A2(n2813), .ZN(n3359) );
  INV_X1 U3641 ( .A(n2812), .ZN(n2815) );
  INV_X1 U3642 ( .A(n2813), .ZN(n2814) );
  NAND2_X1 U3643 ( .A1(n2815), .A2(n2814), .ZN(n3358) );
  OAI22_X1 U3644 ( .A1(n4437), .A2(n3556), .B1(n3746), .B2(n3554), .ZN(n2816)
         );
  XNOR2_X1 U3645 ( .A(n2816), .B(n3533), .ZN(n3440) );
  OAI22_X1 U3646 ( .A1(n4437), .A2(n3557), .B1(n3746), .B2(n3556), .ZN(n3441)
         );
  NAND2_X1 U3647 ( .A1(n2817), .A2(n3441), .ZN(n2820) );
  INV_X1 U3648 ( .A(n3443), .ZN(n2818) );
  NAND2_X1 U3649 ( .A1(n2818), .A2(n2172), .ZN(n2819) );
  NAND2_X1 U3650 ( .A1(n3592), .A2(n2726), .ZN(n2821) );
  OAI21_X1 U3651 ( .B1(n4414), .B2(n3556), .A(n2821), .ZN(n2822) );
  XNOR2_X1 U3652 ( .A(n2822), .B(n3561), .ZN(n2833) );
  OR2_X1 U3653 ( .A1(n4414), .A2(n3557), .ZN(n2824) );
  NAND2_X1 U3654 ( .A1(n3592), .A2(n3560), .ZN(n2823) );
  NAND2_X1 U3655 ( .A1(n2824), .A2(n2823), .ZN(n2834) );
  AND2_X1 U3656 ( .A1(n2833), .A2(n2834), .ZN(n3589) );
  NAND2_X1 U3657 ( .A1(n4389), .A2(n2754), .ZN(n2826) );
  NAND2_X1 U3658 ( .A1(n4373), .A2(n3560), .ZN(n2825) );
  NAND2_X1 U3659 ( .A1(n2826), .A2(n2825), .ZN(n3620) );
  NAND2_X1 U3660 ( .A1(n4389), .A2(n3560), .ZN(n2828) );
  NAND2_X1 U3661 ( .A1(n4373), .A2(n2726), .ZN(n2827) );
  NAND2_X1 U3662 ( .A1(n2828), .A2(n2827), .ZN(n2829) );
  XNOR2_X1 U3663 ( .A(n2829), .B(n3561), .ZN(n3622) );
  OAI22_X1 U3664 ( .A1(n4367), .A2(n3556), .B1(n4349), .B2(n3554), .ZN(n2830)
         );
  XNOR2_X1 U3665 ( .A(n2830), .B(n3561), .ZN(n2839) );
  INV_X1 U3666 ( .A(n2839), .ZN(n2832) );
  OAI22_X1 U3667 ( .A1(n4367), .A2(n3557), .B1(n4349), .B2(n3556), .ZN(n2838)
         );
  INV_X1 U3668 ( .A(n2838), .ZN(n2831) );
  NAND2_X1 U3669 ( .A1(n2832), .A2(n2831), .ZN(n2837) );
  INV_X1 U3670 ( .A(n2833), .ZN(n2836) );
  INV_X1 U3671 ( .A(n2834), .ZN(n2835) );
  NAND2_X1 U3672 ( .A1(n2836), .A2(n2835), .ZN(n3588) );
  OAI211_X1 U3673 ( .C1(n3620), .C2(n3622), .A(n2837), .B(n3588), .ZN(n2841)
         );
  INV_X1 U3674 ( .A(n2837), .ZN(n3625) );
  AND2_X1 U3675 ( .A1(n2839), .A2(n2838), .ZN(n3624) );
  AOI21_X1 U3676 ( .B1(n3620), .B2(n3622), .A(n3624), .ZN(n2840) );
  NAND2_X1 U3677 ( .A1(n4347), .A2(n3560), .ZN(n2843) );
  NAND2_X1 U3678 ( .A1(n4336), .A2(n2726), .ZN(n2842) );
  NAND2_X1 U3679 ( .A1(n2843), .A2(n2842), .ZN(n2844) );
  XNOR2_X1 U3680 ( .A(n2844), .B(n3533), .ZN(n2847) );
  AND2_X1 U3681 ( .A1(n4336), .A2(n2741), .ZN(n2845) );
  AOI21_X1 U3682 ( .B1(n4347), .B2(n2754), .A(n2845), .ZN(n2846) );
  NOR2_X1 U3683 ( .A1(n2847), .A2(n2846), .ZN(n3632) );
  NAND2_X1 U3684 ( .A1(n2847), .A2(n2846), .ZN(n3633) );
  OAI22_X1 U3685 ( .A1(n4295), .A2(n3557), .B1(n3556), .B2(n3676), .ZN(n3607)
         );
  OAI22_X1 U3686 ( .A1(n4295), .A2(n3556), .B1(n3554), .B2(n3676), .ZN(n2848)
         );
  XNOR2_X1 U3687 ( .A(n2848), .B(n3561), .ZN(n3670) );
  NAND2_X1 U3688 ( .A1(n4271), .A2(n3560), .ZN(n2850) );
  NAND2_X1 U3689 ( .A1(n3614), .A2(n2726), .ZN(n2849) );
  NAND2_X1 U3690 ( .A1(n2850), .A2(n2849), .ZN(n2851) );
  XNOR2_X1 U3691 ( .A(n2851), .B(n3533), .ZN(n2853) );
  AND2_X1 U3692 ( .A1(n3614), .A2(n3560), .ZN(n2852) );
  AOI21_X1 U3693 ( .B1(n4271), .B2(n2754), .A(n2852), .ZN(n2854) );
  NOR2_X1 U3694 ( .A1(n2853), .A2(n2854), .ZN(n3611) );
  AOI21_X1 U3695 ( .B1(n3607), .B2(n3670), .A(n3611), .ZN(n2859) );
  INV_X1 U3696 ( .A(n2853), .ZN(n2856) );
  INV_X1 U3697 ( .A(n2854), .ZN(n2855) );
  NOR2_X1 U3698 ( .A1(n2856), .A2(n2855), .ZN(n3610) );
  AOI21_X2 U3699 ( .B1(n3672), .B2(n2859), .A(n2858), .ZN(n3653) );
  NAND2_X1 U3700 ( .A1(n4297), .A2(n3560), .ZN(n2861) );
  NAND2_X1 U3701 ( .A1(n2726), .A2(n4270), .ZN(n2860) );
  NAND2_X1 U3702 ( .A1(n2861), .A2(n2860), .ZN(n2862) );
  XNOR2_X1 U3703 ( .A(n2862), .B(n3533), .ZN(n2865) );
  AND2_X1 U3704 ( .A1(n3560), .A2(n4270), .ZN(n2863) );
  AOI21_X1 U3705 ( .B1(n4297), .B2(n2754), .A(n2863), .ZN(n2864) );
  NOR2_X1 U3706 ( .A1(n2865), .A2(n2864), .ZN(n3651) );
  AND2_X1 U3707 ( .A1(n2865), .A2(n2864), .ZN(n2884) );
  NAND2_X1 U3708 ( .A1(n3663), .A2(n3560), .ZN(n2867) );
  NAND2_X1 U3709 ( .A1(n2726), .A2(n4257), .ZN(n2866) );
  NAND2_X1 U3710 ( .A1(n2867), .A2(n2866), .ZN(n2868) );
  XNOR2_X1 U3711 ( .A(n2868), .B(n3561), .ZN(n2874) );
  INV_X1 U3712 ( .A(n2874), .ZN(n2872) );
  NAND2_X1 U3713 ( .A1(n3663), .A2(n2754), .ZN(n2870) );
  NAND2_X1 U3714 ( .A1(n3560), .A2(n4257), .ZN(n2869) );
  NAND2_X1 U3715 ( .A1(n2870), .A2(n2869), .ZN(n2873) );
  INV_X1 U3716 ( .A(n2873), .ZN(n2871) );
  NAND2_X1 U3717 ( .A1(n2872), .A2(n2871), .ZN(n3509) );
  INV_X1 U3718 ( .A(n3509), .ZN(n2875) );
  AND2_X1 U3719 ( .A1(n2874), .A2(n2873), .ZN(n3508) );
  NOR2_X1 U3720 ( .A1(n2875), .A2(n3508), .ZN(n2886) );
  NAND3_X1 U3721 ( .A1(n3127), .A2(n2878), .A3(n3125), .ZN(n2894) );
  INV_X1 U3722 ( .A(n2917), .ZN(n2882) );
  INV_X1 U3723 ( .A(n2879), .ZN(n2880) );
  OR2_X1 U3724 ( .A1(n3026), .A2(n2880), .ZN(n2881) );
  NAND2_X1 U3725 ( .A1(n2882), .A2(n2881), .ZN(n2887) );
  NOR2_X1 U3726 ( .A1(n2887), .A2(n3123), .ZN(n2883) );
  AOI211_X1 U3727 ( .C1(n3653), .C2(n2184), .A(n3651), .B(n2886), .ZN(n2885)
         );
  AOI211_X1 U3728 ( .C1(n3510), .C2(n2886), .A(n3707), .B(n2885), .ZN(n2906)
         );
  NAND2_X1 U3729 ( .A1(n2887), .A2(n4391), .ZN(n2888) );
  NAND2_X1 U3730 ( .A1(n2894), .A2(n2888), .ZN(n2889) );
  NAND2_X1 U3731 ( .A1(n2889), .A2(n3122), .ZN(n3045) );
  NAND2_X1 U3732 ( .A1(n2890), .A2(n2916), .ZN(n2891) );
  OAI21_X1 U3733 ( .B1(n3045), .B2(n2891), .A(STATE_REG_SCAN_IN), .ZN(n2895)
         );
  NOR2_X1 U3734 ( .A1(n2892), .A2(n4690), .ZN(n2893) );
  NAND2_X1 U3735 ( .A1(n2894), .A2(n2896), .ZN(n3044) );
  NOR2_X1 U3736 ( .A1(n3689), .A2(n4260), .ZN(n2905) );
  INV_X1 U3737 ( .A(n4297), .ZN(n4252) );
  NOR2_X1 U3738 ( .A1(n3867), .A2(n2912), .ZN(n2897) );
  OAI22_X1 U3739 ( .A1(n4252), .A2(n3655), .B1(STATE_REG_SCAN_IN), .B2(n3978), 
        .ZN(n2904) );
  NOR2_X1 U3740 ( .A1(n3867), .A2(n4609), .ZN(n2898) );
  NOR2_X1 U3741 ( .A1(n3123), .A2(n4391), .ZN(n2899) );
  NAND2_X1 U3742 ( .A1(n2900), .A2(n2899), .ZN(n2902) );
  OAI22_X1 U3743 ( .A1(n4236), .A2(n3703), .B1(n3677), .B2(n4251), .ZN(n2903)
         );
  NAND2_X1 U3744 ( .A1(n2908), .A2(n2907), .ZN(n4095) );
  OR2_X1 U3745 ( .A1(n4095), .A2(REG2_REG_0__SCAN_IN), .ZN(n2909) );
  AND2_X1 U3746 ( .A1(n4609), .A2(n2909), .ZN(n4625) );
  XOR2_X1 U3747 ( .A(n2911), .B(n2910), .Z(n3056) );
  OR3_X1 U3748 ( .A1(n3056), .A2(n4624), .A3(n2912), .ZN(n2915) );
  NAND2_X1 U3749 ( .A1(n4609), .A2(n4624), .ZN(n3866) );
  INV_X1 U3750 ( .A(n3866), .ZN(n2913) );
  AND2_X1 U3751 ( .A1(IR_REG_0__SCAN_IN), .A2(REG2_REG_0__SCAN_IN), .ZN(n4020)
         );
  AOI21_X1 U3752 ( .B1(n2913), .B2(n4020), .A(n4017), .ZN(n2914) );
  OAI211_X1 U3753 ( .C1(IR_REG_0__SCAN_IN), .C2(n4625), .A(n2915), .B(n2914), 
        .ZN(n4043) );
  INV_X1 U3754 ( .A(n4043), .ZN(n2952) );
  INV_X1 U3755 ( .A(n4621), .ZN(n2947) );
  OR2_X1 U3756 ( .A1(n2916), .A2(U3149), .ZN(n3871) );
  NAND2_X1 U3757 ( .A1(n3123), .A2(n3871), .ZN(n2920) );
  NAND2_X1 U3758 ( .A1(n2917), .A2(n2916), .ZN(n2918) );
  INV_X1 U3759 ( .A(n2919), .ZN(n2921) );
  NAND2_X1 U3760 ( .A1(n4660), .A2(ADDR_REG_4__SCAN_IN), .ZN(n2922) );
  NAND2_X1 U3761 ( .A1(REG3_REG_4__SCAN_IN), .A2(U3149), .ZN(n3166) );
  OAI211_X1 U3762 ( .C1(n2947), .C2(n4673), .A(n2922), .B(n3166), .ZN(n2951)
         );
  NAND2_X1 U3763 ( .A1(n2940), .A2(REG2_REG_2__SCAN_IN), .ZN(n2927) );
  OAI21_X1 U3764 ( .B1(n2007), .B2(REG2_REG_2__SCAN_IN), .A(n2927), .ZN(n4034)
         );
  INV_X1 U3765 ( .A(n4034), .ZN(n2926) );
  INV_X1 U3766 ( .A(REG2_REG_1__SCAN_IN), .ZN(n2923) );
  NAND2_X1 U3767 ( .A1(n2933), .A2(REG2_REG_1__SCAN_IN), .ZN(n2924) );
  NAND2_X1 U3768 ( .A1(n4019), .A2(n4020), .ZN(n4018) );
  NAND2_X1 U3769 ( .A1(n2932), .A2(REG2_REG_1__SCAN_IN), .ZN(n4035) );
  NAND2_X1 U3770 ( .A1(n4018), .A2(n4035), .ZN(n2925) );
  NAND2_X1 U3771 ( .A1(n2991), .A2(REG2_REG_3__SCAN_IN), .ZN(n2930) );
  NAND2_X1 U3772 ( .A1(n2928), .A2(n2943), .ZN(n2929) );
  NAND2_X1 U3773 ( .A1(n2930), .A2(n2929), .ZN(n3001) );
  XNOR2_X1 U3774 ( .A(n3003), .B(REG2_REG_4__SCAN_IN), .ZN(n2949) );
  INV_X1 U3775 ( .A(n2933), .ZN(n2932) );
  INV_X1 U3776 ( .A(REG1_REG_1__SCAN_IN), .ZN(n2931) );
  NAND2_X1 U3777 ( .A1(n2932), .A2(n2931), .ZN(n2935) );
  NAND2_X1 U3778 ( .A1(n2933), .A2(REG1_REG_1__SCAN_IN), .ZN(n2934) );
  NAND2_X1 U3779 ( .A1(n2935), .A2(n2934), .ZN(n2937) );
  AND2_X1 U3780 ( .A1(IR_REG_0__SCAN_IN), .A2(REG1_REG_0__SCAN_IN), .ZN(n2936)
         );
  NAND2_X1 U3781 ( .A1(n2932), .A2(REG1_REG_1__SCAN_IN), .ZN(n4031) );
  NAND2_X1 U3782 ( .A1(n4021), .A2(n4031), .ZN(n2941) );
  INV_X1 U3783 ( .A(REG1_REG_2__SCAN_IN), .ZN(n2938) );
  OAI21_X1 U3784 ( .B1(n2007), .B2(n2938), .A(n2939), .ZN(n4029) );
  NAND2_X1 U3785 ( .A1(n2941), .A2(n4029), .ZN(n4033) );
  NAND2_X1 U3786 ( .A1(n2007), .A2(REG1_REG_2__SCAN_IN), .ZN(n2942) );
  NAND2_X1 U3787 ( .A1(n4033), .A2(n2942), .ZN(n2944) );
  XNOR2_X1 U3788 ( .A(n2944), .B(n2319), .ZN(n2990) );
  NAND2_X1 U3789 ( .A1(n2990), .A2(REG1_REG_3__SCAN_IN), .ZN(n2946) );
  NAND2_X1 U3790 ( .A1(n2944), .A2(n2943), .ZN(n2945) );
  XNOR2_X1 U3791 ( .A(n2999), .B(REG1_REG_4__SCAN_IN), .ZN(n2948) );
  OAI22_X1 U3792 ( .A1(n2949), .A2(n3470), .B1(n4657), .B2(n2948), .ZN(n2950)
         );
  OR3_X1 U3793 ( .A1(n2952), .A2(n2951), .A3(n2950), .ZN(U3244) );
  INV_X1 U3794 ( .A(DATAI_3_), .ZN(n2953) );
  MUX2_X1 U3795 ( .A(n2953), .B(n2319), .S(STATE_REG_SCAN_IN), .Z(n2954) );
  INV_X1 U3796 ( .A(n2954), .ZN(U3349) );
  MUX2_X1 U3797 ( .A(n2955), .B(n3155), .S(STATE_REG_SCAN_IN), .Z(n2956) );
  INV_X1 U3798 ( .A(n2956), .ZN(U3344) );
  MUX2_X1 U3799 ( .A(n3268), .B(n2406), .S(U3149), .Z(n2957) );
  INV_X1 U3800 ( .A(n2957), .ZN(U3343) );
  INV_X1 U3801 ( .A(DATAI_26_), .ZN(n2959) );
  NAND2_X1 U3802 ( .A1(n2979), .A2(STATE_REG_SCAN_IN), .ZN(n2958) );
  OAI21_X1 U3803 ( .B1(STATE_REG_SCAN_IN), .B2(n2959), .A(n2958), .ZN(U3326)
         );
  INV_X1 U3804 ( .A(DATAI_21_), .ZN(n2961) );
  NAND2_X1 U3805 ( .A1(n2644), .A2(STATE_REG_SCAN_IN), .ZN(n2960) );
  OAI21_X1 U3806 ( .B1(STATE_REG_SCAN_IN), .B2(n2961), .A(n2960), .ZN(U3331)
         );
  INV_X1 U3807 ( .A(DATAI_20_), .ZN(n2964) );
  NAND2_X1 U3808 ( .A1(n2962), .A2(STATE_REG_SCAN_IN), .ZN(n2963) );
  OAI21_X1 U3809 ( .B1(STATE_REG_SCAN_IN), .B2(n2964), .A(n2963), .ZN(U3332)
         );
  INV_X1 U3810 ( .A(DATAI_29_), .ZN(n2967) );
  NAND2_X1 U3811 ( .A1(n2965), .A2(STATE_REG_SCAN_IN), .ZN(n2966) );
  OAI21_X1 U3812 ( .B1(STATE_REG_SCAN_IN), .B2(n2967), .A(n2966), .ZN(U3323)
         );
  INV_X1 U3813 ( .A(DATAI_24_), .ZN(n2969) );
  NAND2_X1 U3814 ( .A1(n2677), .A2(STATE_REG_SCAN_IN), .ZN(n2968) );
  OAI21_X1 U3815 ( .B1(STATE_REG_SCAN_IN), .B2(n2969), .A(n2968), .ZN(U3328)
         );
  INV_X1 U3816 ( .A(DATAI_22_), .ZN(n2971) );
  NAND2_X1 U3817 ( .A1(n3868), .A2(STATE_REG_SCAN_IN), .ZN(n2970) );
  OAI21_X1 U3818 ( .B1(STATE_REG_SCAN_IN), .B2(n2971), .A(n2970), .ZN(U3330)
         );
  INV_X1 U3819 ( .A(DATAI_12_), .ZN(n2972) );
  MUX2_X1 U3820 ( .A(n2972), .B(n3429), .S(STATE_REG_SCAN_IN), .Z(n2973) );
  INV_X1 U3821 ( .A(n2973), .ZN(U3340) );
  INV_X1 U3822 ( .A(D_REG_1__SCAN_IN), .ZN(n2978) );
  INV_X1 U3823 ( .A(n2976), .ZN(n4610) );
  NOR3_X1 U3824 ( .A1(n4690), .A2(n2979), .A3(n4610), .ZN(n2977) );
  AOI21_X1 U3825 ( .B1(n4689), .B2(n2978), .A(n2977), .ZN(U3459) );
  INV_X1 U3826 ( .A(D_REG_0__SCAN_IN), .ZN(n2981) );
  NOR3_X1 U3827 ( .A1(n2677), .A2(n4690), .A3(n2979), .ZN(n2980) );
  AOI21_X1 U3828 ( .B1(n4689), .B2(n2981), .A(n2980), .ZN(U3458) );
  NOR2_X1 U3829 ( .A1(n4660), .A2(U4043), .ZN(U3148) );
  NAND2_X1 U3830 ( .A1(n2329), .A2(REG2_REG_30__SCAN_IN), .ZN(n2983) );
  NAND2_X1 U3831 ( .A1(n2009), .A2(REG1_REG_30__SCAN_IN), .ZN(n2982) );
  OAI211_X1 U3832 ( .C1(n2301), .C2(n4549), .A(n2983), .B(n2982), .ZN(n4120)
         );
  NAND2_X1 U3833 ( .A1(U4043), .A2(n4120), .ZN(n2984) );
  OAI21_X1 U3834 ( .B1(U4043), .B2(n3979), .A(n2984), .ZN(U3580) );
  INV_X1 U3835 ( .A(DATAO_REG_4__SCAN_IN), .ZN(n3936) );
  NAND2_X1 U3836 ( .A1(n2985), .A2(U4043), .ZN(n2986) );
  OAI21_X1 U3837 ( .B1(U4043), .B2(n3936), .A(n2986), .ZN(U3554) );
  INV_X1 U3838 ( .A(DATAO_REG_7__SCAN_IN), .ZN(n3937) );
  NAND2_X1 U3839 ( .A1(n2367), .A2(U4043), .ZN(n2987) );
  OAI21_X1 U3840 ( .B1(U4043), .B2(n3937), .A(n2987), .ZN(U3557) );
  INV_X1 U3841 ( .A(DATAO_REG_8__SCAN_IN), .ZN(n3986) );
  NAND2_X1 U3842 ( .A1(n3319), .A2(U4043), .ZN(n2988) );
  OAI21_X1 U3843 ( .B1(U4043), .B2(n3986), .A(n2988), .ZN(U3558) );
  INV_X1 U3844 ( .A(DATAO_REG_1__SCAN_IN), .ZN(n3941) );
  NAND2_X1 U3845 ( .A1(n3082), .A2(U4043), .ZN(n2989) );
  OAI21_X1 U3846 ( .B1(U4043), .B2(n3941), .A(n2989), .ZN(U3551) );
  XNOR2_X1 U3847 ( .A(n2990), .B(REG1_REG_3__SCAN_IN), .ZN(n2996) );
  XNOR2_X1 U3848 ( .A(n2991), .B(n2321), .ZN(n2994) );
  NOR2_X1 U3849 ( .A1(STATE_REG_SCAN_IN), .A2(n2320), .ZN(n3108) );
  AOI21_X1 U3850 ( .B1(n4660), .B2(ADDR_REG_3__SCAN_IN), .A(n3108), .ZN(n2992)
         );
  OAI21_X1 U3851 ( .B1(n2319), .B2(n4673), .A(n2992), .ZN(n2993) );
  AOI21_X1 U3852 ( .B1(n4670), .B2(n2994), .A(n2993), .ZN(n2995) );
  OAI21_X1 U3853 ( .B1(n2996), .B2(n4657), .A(n2995), .ZN(U3243) );
  MUX2_X1 U3854 ( .A(REG1_REG_5__SCAN_IN), .B(n4737), .S(n3019), .Z(n3016) );
  INV_X1 U3855 ( .A(n3019), .ZN(n4620) );
  XNOR2_X1 U3856 ( .A(n3032), .B(REG1_REG_6__SCAN_IN), .ZN(n3011) );
  INV_X1 U3857 ( .A(REG2_REG_5__SCAN_IN), .ZN(n3004) );
  MUX2_X1 U3858 ( .A(REG2_REG_5__SCAN_IN), .B(n3004), .S(n3019), .Z(n3013) );
  XNOR2_X1 U3859 ( .A(n3035), .B(n4619), .ZN(n3037) );
  XOR2_X1 U3860 ( .A(n3037), .B(REG2_REG_6__SCAN_IN), .Z(n3009) );
  INV_X1 U3861 ( .A(n4619), .ZN(n3007) );
  AND2_X1 U3862 ( .A1(U3149), .A2(REG3_REG_6__SCAN_IN), .ZN(n3140) );
  AOI21_X1 U3863 ( .B1(n4660), .B2(ADDR_REG_6__SCAN_IN), .A(n3140), .ZN(n3006)
         );
  OAI21_X1 U3864 ( .B1(n3007), .B2(n4673), .A(n3006), .ZN(n3008) );
  AOI21_X1 U3865 ( .B1(n3009), .B2(n4670), .A(n3008), .ZN(n3010) );
  OAI21_X1 U3866 ( .B1(n3011), .B2(n4657), .A(n3010), .ZN(U3246) );
  AOI211_X1 U3867 ( .C1(n3014), .C2(n3013), .A(n3470), .B(n3012), .ZN(n3022)
         );
  AOI211_X1 U3868 ( .C1(n3017), .C2(n3016), .A(n4657), .B(n3015), .ZN(n3021)
         );
  AND2_X1 U3869 ( .A1(U3149), .A2(REG3_REG_5__SCAN_IN), .ZN(n3504) );
  AOI21_X1 U3870 ( .B1(n4660), .B2(ADDR_REG_5__SCAN_IN), .A(n3504), .ZN(n3018)
         );
  OAI21_X1 U3871 ( .B1(n3019), .B2(n4673), .A(n3018), .ZN(n3020) );
  OR3_X1 U3872 ( .A1(n3022), .A2(n3021), .A3(n3020), .ZN(U3245) );
  NAND2_X1 U3873 ( .A1(n3023), .A2(n3024), .ZN(n3785) );
  AND2_X1 U3874 ( .A1(n3785), .A2(n3025), .ZN(n3763) );
  INV_X1 U3875 ( .A(n3763), .ZN(n4679) );
  NOR2_X1 U3876 ( .A1(n3023), .A2(n3026), .ZN(n4677) );
  INV_X1 U3877 ( .A(n4417), .ZN(n3416) );
  NOR2_X1 U3878 ( .A1(n3416), .A2(n4393), .ZN(n3028) );
  OAI22_X1 U3879 ( .A1(n3763), .A2(n3028), .B1(n3027), .B2(n4436), .ZN(n4675)
         );
  AOI211_X1 U3880 ( .C1(n4712), .C2(n4679), .A(n4677), .B(n4675), .ZN(n4698)
         );
  NAND2_X1 U3881 ( .A1(n2712), .A2(REG1_REG_0__SCAN_IN), .ZN(n3029) );
  OAI21_X1 U3882 ( .B1(n4698), .B2(n2712), .A(n3029), .ZN(U3518) );
  MUX2_X1 U3883 ( .A(n4739), .B(REG1_REG_7__SCAN_IN), .S(n4618), .Z(n3033) );
  INV_X1 U3884 ( .A(n3030), .ZN(n3031) );
  XOR2_X1 U3885 ( .A(n3033), .B(n3066), .Z(n3042) );
  INV_X1 U3886 ( .A(n4618), .ZN(n3064) );
  NAND2_X1 U3887 ( .A1(U3149), .A2(REG3_REG_7__SCAN_IN), .ZN(n3214) );
  NAND2_X1 U3888 ( .A1(n4660), .A2(ADDR_REG_7__SCAN_IN), .ZN(n3034) );
  OAI211_X1 U3889 ( .C1(n4673), .C2(n3064), .A(n3214), .B(n3034), .ZN(n3041)
         );
  NOR2_X1 U3890 ( .A1(n3035), .A2(n3007), .ZN(n3036) );
  INV_X1 U3891 ( .A(REG2_REG_7__SCAN_IN), .ZN(n3199) );
  MUX2_X1 U3892 ( .A(n3199), .B(REG2_REG_7__SCAN_IN), .S(n4618), .Z(n3038) );
  NOR2_X1 U3893 ( .A1(n3039), .A2(n3038), .ZN(n3060) );
  AOI211_X1 U3894 ( .C1(n3039), .C2(n3038), .A(n3470), .B(n3060), .ZN(n3040)
         );
  AOI211_X1 U3895 ( .C1(n3042), .C2(n4654), .A(n3041), .B(n3040), .ZN(n3043)
         );
  INV_X1 U3896 ( .A(n3043), .ZN(U3247) );
  INV_X1 U3897 ( .A(n3044), .ZN(n3046) );
  NOR3_X1 U3898 ( .A1(n3046), .A2(n3045), .A3(n3123), .ZN(n3101) );
  INV_X1 U3899 ( .A(REG3_REG_1__SCAN_IN), .ZN(n3233) );
  OAI22_X1 U3900 ( .A1(n3703), .A2(n2315), .B1(n3047), .B2(n3655), .ZN(n3048)
         );
  AOI21_X1 U3901 ( .B1(n3223), .B2(n3700), .A(n3048), .ZN(n3054) );
  AOI21_X1 U3902 ( .B1(n3050), .B2(n3049), .A(n3707), .ZN(n3052) );
  NAND2_X1 U3903 ( .A1(n3052), .A2(n3051), .ZN(n3053) );
  OAI211_X1 U3904 ( .C1(n3101), .C2(n3233), .A(n3054), .B(n3053), .ZN(U3219)
         );
  INV_X1 U3905 ( .A(REG3_REG_0__SCAN_IN), .ZN(n3058) );
  OAI22_X1 U3906 ( .A1(n3677), .A2(n3023), .B1(n3703), .B2(n3027), .ZN(n3055)
         );
  AOI21_X1 U3907 ( .B1(n3673), .B2(n3056), .A(n3055), .ZN(n3057) );
  OAI21_X1 U3908 ( .B1(n3101), .B2(n3058), .A(n3057), .ZN(U3229) );
  INV_X1 U3909 ( .A(n3155), .ZN(n3061) );
  XNOR2_X1 U3910 ( .A(n3144), .B(REG2_REG_8__SCAN_IN), .ZN(n3070) );
  NAND2_X1 U3911 ( .A1(REG3_REG_8__SCAN_IN), .A2(U3149), .ZN(n3259) );
  INV_X1 U3912 ( .A(n3259), .ZN(n3063) );
  NOR2_X1 U3913 ( .A1(n4673), .A2(n3155), .ZN(n3062) );
  AOI211_X1 U3914 ( .C1(n4660), .C2(ADDR_REG_8__SCAN_IN), .A(n3063), .B(n3062), 
        .ZN(n3069) );
  NAND2_X1 U3915 ( .A1(n4618), .A2(REG1_REG_7__SCAN_IN), .ZN(n3065) );
  OAI211_X1 U3916 ( .C1(n3067), .C2(REG1_REG_8__SCAN_IN), .A(n3157), .B(n4654), 
        .ZN(n3068) );
  OAI211_X1 U3917 ( .C1(n3070), .C2(n3470), .A(n3069), .B(n3068), .ZN(U3248)
         );
  NAND2_X1 U3918 ( .A1(n3072), .A2(n2233), .ZN(n3228) );
  NAND2_X1 U3919 ( .A1(n3228), .A2(n3073), .ZN(n3074) );
  NAND2_X1 U3920 ( .A1(n3074), .A2(n3750), .ZN(n3076) );
  NAND2_X1 U3921 ( .A1(n3076), .A2(n3075), .ZN(n3252) );
  NAND3_X1 U3922 ( .A1(n3077), .A2(n3078), .A3(n3787), .ZN(n3079) );
  NAND2_X1 U3923 ( .A1(n3080), .A2(n3079), .ZN(n3081) );
  NAND2_X1 U3924 ( .A1(n3081), .A2(n4393), .ZN(n3086) );
  NAND2_X1 U3925 ( .A1(n3252), .A2(n3416), .ZN(n3085) );
  AOI22_X1 U3926 ( .A1(n4388), .A2(n4016), .B1(n3082), .B2(n4386), .ZN(n3084)
         );
  NAND2_X1 U3927 ( .A1(n2742), .A2(n4439), .ZN(n3083) );
  NAND4_X1 U3928 ( .A1(n3086), .A2(n3085), .A3(n3084), .A4(n3083), .ZN(n3250)
         );
  AOI21_X1 U3929 ( .B1(n4712), .B2(n3252), .A(n3250), .ZN(n3092) );
  OAI21_X1 U3930 ( .B1(n3220), .B2(n3087), .A(n3186), .ZN(n3255) );
  OAI22_X1 U3931 ( .A1(n4540), .A2(n3255), .B1(n4741), .B2(n2938), .ZN(n3088)
         );
  INV_X1 U3932 ( .A(n3088), .ZN(n3089) );
  OAI21_X1 U3933 ( .B1(n3092), .B2(n2712), .A(n3089), .ZN(U3520) );
  INV_X1 U3934 ( .A(REG0_REG_2__SCAN_IN), .ZN(n3958) );
  OAI22_X1 U3935 ( .A1(n4606), .A2(n3255), .B1(n4731), .B2(n3958), .ZN(n3090)
         );
  INV_X1 U3936 ( .A(n3090), .ZN(n3091) );
  OAI21_X1 U3937 ( .B1(n3092), .B2(n4729), .A(n3091), .ZN(U3471) );
  INV_X1 U3938 ( .A(REG3_REG_2__SCAN_IN), .ZN(n3100) );
  OAI21_X1 U3939 ( .B1(n3095), .B2(n3094), .A(n3093), .ZN(n3096) );
  NAND2_X1 U3940 ( .A1(n3096), .A2(n3673), .ZN(n3099) );
  OAI22_X1 U3941 ( .A1(n3703), .A2(n3168), .B1(n3027), .B2(n3655), .ZN(n3097)
         );
  AOI21_X1 U3942 ( .B1(n2742), .B2(n3700), .A(n3097), .ZN(n3098) );
  OAI211_X1 U3943 ( .C1(n3101), .C2(n3100), .A(n3099), .B(n3098), .ZN(U3234)
         );
  NAND2_X1 U3944 ( .A1(n3093), .A2(n3103), .ZN(n3104) );
  XNOR2_X1 U3945 ( .A(n3102), .B(n3104), .ZN(n3105) );
  NAND2_X1 U3946 ( .A1(n3105), .A2(n3673), .ZN(n3110) );
  OAI22_X1 U3947 ( .A1(n3677), .A2(n3106), .B1(n3703), .B2(n3502), .ZN(n3107)
         );
  AOI211_X1 U3948 ( .C1(n3701), .C2(n2745), .A(n3108), .B(n3107), .ZN(n3109)
         );
  OAI211_X1 U3949 ( .C1(REG3_REG_3__SCAN_IN), .C2(n3689), .A(n3110), .B(n3109), 
        .ZN(U3215) );
  INV_X1 U3950 ( .A(DATAO_REG_21__SCAN_IN), .ZN(n3939) );
  NAND2_X1 U3951 ( .A1(n3663), .A2(U4043), .ZN(n3111) );
  OAI21_X1 U3952 ( .B1(U4043), .B2(n3939), .A(n3111), .ZN(U3571) );
  XOR2_X1 U3953 ( .A(n3755), .B(n3112), .Z(n3118) );
  OR2_X1 U3954 ( .A1(n3114), .A2(n3755), .ZN(n3240) );
  INV_X1 U3955 ( .A(n3240), .ZN(n3113) );
  AOI21_X1 U3956 ( .B1(n3755), .B2(n3114), .A(n3113), .ZN(n4713) );
  AOI22_X1 U3957 ( .A1(n2616), .A2(n4388), .B1(n4386), .B2(n4016), .ZN(n3115)
         );
  OAI21_X1 U3958 ( .B1(n3120), .B2(n4391), .A(n3115), .ZN(n3116) );
  AOI21_X1 U3959 ( .B1(n4713), .B2(n3416), .A(n3116), .ZN(n3117) );
  OAI21_X1 U3960 ( .B1(n4442), .B2(n3118), .A(n3117), .ZN(n4710) );
  OAI211_X1 U3961 ( .C1(n3119), .C2(n3120), .A(n3246), .B(n4721), .ZN(n4709)
         );
  OAI22_X1 U3962 ( .A1(n4709), .A2(n4611), .B1(n4360), .B2(n3121), .ZN(n3130)
         );
  INV_X1 U3963 ( .A(n3122), .ZN(n3124) );
  NOR2_X1 U3964 ( .A1(n3124), .A2(n3123), .ZN(n3126) );
  NAND4_X1 U3965 ( .A1(n3128), .A2(n3127), .A3(n3126), .A4(n3125), .ZN(n3129)
         );
  OAI21_X1 U3966 ( .B1(n4710), .B2(n3130), .A(n4682), .ZN(n3134) );
  OR2_X1 U3967 ( .A1(n3131), .A2(n4088), .ZN(n3205) );
  INV_X1 U3968 ( .A(n3205), .ZN(n3132) );
  AOI22_X1 U3969 ( .A1(n4713), .A2(n4680), .B1(REG2_REG_4__SCAN_IN), .B2(n4431), .ZN(n3133) );
  NAND2_X1 U3970 ( .A1(n3134), .A2(n3133), .ZN(U3286) );
  XOR2_X1 U3971 ( .A(n3136), .B(n3135), .Z(n3137) );
  XNOR2_X1 U3972 ( .A(n3138), .B(n3137), .ZN(n3143) );
  OAI22_X1 U3973 ( .A1(n3677), .A2(n3285), .B1(n3703), .B2(n3292), .ZN(n3139)
         );
  AOI211_X1 U3974 ( .C1(n3701), .C2(n2616), .A(n3140), .B(n3139), .ZN(n3142)
         );
  NAND2_X1 U3975 ( .A1(n3705), .A2(n3286), .ZN(n3141) );
  OAI211_X1 U3976 ( .C1(n3143), .C2(n3707), .A(n3142), .B(n3141), .ZN(U3236)
         );
  NAND2_X1 U3977 ( .A1(n3144), .A2(REG2_REG_8__SCAN_IN), .ZN(n3148) );
  INV_X1 U3978 ( .A(n3145), .ZN(n3146) );
  NAND2_X1 U3979 ( .A1(n3146), .A2(n3061), .ZN(n3147) );
  NAND2_X1 U3980 ( .A1(n3148), .A2(n3147), .ZN(n3150) );
  INV_X1 U3981 ( .A(REG2_REG_9__SCAN_IN), .ZN(n3264) );
  MUX2_X1 U3982 ( .A(REG2_REG_9__SCAN_IN), .B(n3264), .S(n3268), .Z(n3152) );
  NAND2_X1 U3983 ( .A1(n3150), .A2(n3149), .ZN(n3266) );
  INV_X1 U3984 ( .A(n3266), .ZN(n3151) );
  AOI211_X1 U3985 ( .C1(n3153), .C2(n3152), .A(n3470), .B(n3151), .ZN(n3164)
         );
  XNOR2_X1 U3986 ( .A(n3268), .B(REG1_REG_9__SCAN_IN), .ZN(n3158) );
  NAND2_X1 U3987 ( .A1(n3159), .A2(n3158), .ZN(n3270) );
  OAI211_X1 U3988 ( .C1(n3159), .C2(n3158), .A(n3270), .B(n4654), .ZN(n3162)
         );
  NAND2_X1 U3989 ( .A1(U3149), .A2(REG3_REG_9__SCAN_IN), .ZN(n3320) );
  INV_X1 U3990 ( .A(n3320), .ZN(n3160) );
  AOI21_X1 U3991 ( .B1(n4660), .B2(ADDR_REG_9__SCAN_IN), .A(n3160), .ZN(n3161)
         );
  OAI211_X1 U3992 ( .C1(n4673), .C2(n3268), .A(n3162), .B(n3161), .ZN(n3163)
         );
  OR2_X1 U3993 ( .A1(n3164), .A2(n3163), .ZN(U3249) );
  AOI22_X1 U3994 ( .A1(n3165), .A2(n3700), .B1(n3691), .B2(n2616), .ZN(n3167)
         );
  OAI211_X1 U3995 ( .C1(n3168), .C2(n3655), .A(n3167), .B(n3166), .ZN(n3176)
         );
  NAND2_X1 U3996 ( .A1(n3093), .A2(n3169), .ZN(n3170) );
  AND2_X1 U3997 ( .A1(n3171), .A2(n3170), .ZN(n3174) );
  AOI211_X1 U3998 ( .C1(n2762), .C2(n3174), .A(n3707), .B(n2042), .ZN(n3175)
         );
  AOI211_X1 U3999 ( .C1(n3177), .C2(n3705), .A(n3176), .B(n3175), .ZN(n3178)
         );
  INV_X1 U4000 ( .A(n3178), .ZN(U3227) );
  XNOR2_X1 U4001 ( .A(n3179), .B(n3754), .ZN(n4704) );
  INV_X1 U4002 ( .A(n4680), .ZN(n3234) );
  OAI21_X1 U4003 ( .B1(n3754), .B2(n3181), .A(n3180), .ZN(n3184) );
  AND2_X1 U4004 ( .A1(n3187), .A2(n4439), .ZN(n3183) );
  OAI22_X1 U4005 ( .A1(n2315), .A2(n4434), .B1(n3502), .B2(n4436), .ZN(n3182)
         );
  AOI211_X1 U4006 ( .C1(n3184), .C2(n4393), .A(n3183), .B(n3182), .ZN(n3185)
         );
  OAI21_X1 U4007 ( .B1(n4704), .B2(n4417), .A(n3185), .ZN(n4705) );
  NAND2_X1 U4008 ( .A1(n4705), .A2(n4682), .ZN(n3190) );
  AOI21_X1 U4009 ( .B1(n3187), .B2(n3186), .A(n3119), .ZN(n4707) );
  OAI22_X1 U4010 ( .A1(n4682), .A2(n2321), .B1(n4360), .B2(REG3_REG_3__SCAN_IN), .ZN(n3188) );
  AOI21_X1 U4011 ( .B1(n4358), .B2(n4707), .A(n3188), .ZN(n3189) );
  OAI211_X1 U4012 ( .C1(n4704), .C2(n3234), .A(n3190), .B(n3189), .ZN(U3287)
         );
  INV_X1 U4013 ( .A(n3800), .ZN(n3756) );
  XNOR2_X1 U4014 ( .A(n3191), .B(n3756), .ZN(n3194) );
  AOI22_X1 U4015 ( .A1(n3319), .A2(n4388), .B1(n4386), .B2(n4015), .ZN(n3192)
         );
  OAI21_X1 U4016 ( .B1(n2699), .B2(n4391), .A(n3192), .ZN(n3193) );
  AOI21_X1 U4017 ( .B1(n3194), .B2(n4393), .A(n3193), .ZN(n4728) );
  INV_X1 U4018 ( .A(n3195), .ZN(n3297) );
  OR2_X1 U4019 ( .A1(n3246), .A2(n3196), .ZN(n3284) );
  AOI21_X1 U4020 ( .B1(n3284), .B2(n3213), .A(n2725), .ZN(n3197) );
  NAND2_X1 U4021 ( .A1(n3297), .A2(n3197), .ZN(n4727) );
  INV_X1 U4022 ( .A(n4727), .ZN(n3201) );
  INV_X1 U4023 ( .A(n3217), .ZN(n3198) );
  OAI22_X1 U4024 ( .A1(n4682), .A2(n3199), .B1(n3198), .B2(n4360), .ZN(n3200)
         );
  AOI21_X1 U4025 ( .B1(n3201), .B2(n4326), .A(n3200), .ZN(n3210) );
  OR2_X1 U4026 ( .A1(n3283), .A2(n4015), .ZN(n3204) );
  NAND2_X1 U4027 ( .A1(n3283), .A2(n4015), .ZN(n3202) );
  NAND2_X1 U4028 ( .A1(n3202), .A2(n3285), .ZN(n3203) );
  AND2_X1 U4029 ( .A1(n3204), .A2(n3203), .ZN(n3207) );
  NAND2_X1 U4030 ( .A1(n3207), .A2(n3800), .ZN(n4725) );
  NAND2_X1 U4031 ( .A1(n4417), .A2(n3205), .ZN(n3206) );
  INV_X1 U4032 ( .A(n3207), .ZN(n3208) );
  NAND2_X1 U4033 ( .A1(n3208), .A2(n3756), .ZN(n4723) );
  NAND3_X1 U4034 ( .A1(n4725), .A2(n4452), .A3(n4723), .ZN(n3209) );
  OAI211_X1 U4035 ( .C1(n4728), .C2(n4431), .A(n3210), .B(n3209), .ZN(U3283)
         );
  XNOR2_X1 U4036 ( .A(n3211), .B(n3212), .ZN(n3219) );
  AOI22_X1 U4037 ( .A1(n3701), .A2(n4015), .B1(n3700), .B2(n3213), .ZN(n3215)
         );
  OAI211_X1 U4038 ( .C1(n3387), .C2(n3703), .A(n3215), .B(n3214), .ZN(n3216)
         );
  AOI21_X1 U4039 ( .B1(n3217), .B2(n3705), .A(n3216), .ZN(n3218) );
  OAI21_X1 U4040 ( .B1(n3219), .B2(n3707), .A(n3218), .ZN(U3210) );
  AOI21_X1 U4041 ( .B1(n3221), .B2(n3223), .A(n3220), .ZN(n4702) );
  NAND2_X1 U4042 ( .A1(n3072), .A2(n3025), .ZN(n3222) );
  NAND2_X1 U40430 ( .A1(n3077), .A2(n3222), .ZN(n3227) );
  NAND2_X1 U4044 ( .A1(n3223), .A2(n4439), .ZN(n3225) );
  NAND2_X1 U4045 ( .A1(n3024), .A2(n4386), .ZN(n3224) );
  OAI211_X1 U4046 ( .C1(n2315), .C2(n4436), .A(n3225), .B(n3224), .ZN(n3226)
         );
  AOI21_X1 U4047 ( .B1(n3227), .B2(n4393), .A(n3226), .ZN(n3231) );
  OR2_X1 U4048 ( .A1(n2233), .A2(n3072), .ZN(n3229) );
  AND2_X1 U4049 ( .A1(n3229), .A2(n3228), .ZN(n3232) );
  NAND2_X1 U4050 ( .A1(n3232), .A2(n3416), .ZN(n3230) );
  NAND2_X1 U4051 ( .A1(n3231), .A2(n3230), .ZN(n4701) );
  MUX2_X1 U4052 ( .A(n4701), .B(REG2_REG_1__SCAN_IN), .S(n4684), .Z(n3236) );
  INV_X1 U4053 ( .A(n3232), .ZN(n4699) );
  OAI22_X1 U4054 ( .A1(n3234), .A2(n4699), .B1(n3233), .B2(n4360), .ZN(n3235)
         );
  AOI211_X1 U4055 ( .C1(n4358), .C2(n4702), .A(n3236), .B(n3235), .ZN(n3237)
         );
  INV_X1 U4056 ( .A(n3237), .ZN(U3289) );
  INV_X1 U4057 ( .A(n3797), .ZN(n3238) );
  AND2_X1 U4058 ( .A1(n3238), .A2(n3809), .ZN(n3752) );
  NAND2_X1 U4059 ( .A1(n3240), .A2(n3239), .ZN(n3241) );
  XOR2_X1 U4060 ( .A(n3752), .B(n3241), .Z(n4716) );
  XOR2_X1 U4061 ( .A(n3242), .B(n3752), .Z(n3245) );
  AOI22_X1 U4062 ( .A1(n2985), .A2(n4386), .B1(n4388), .B2(n4015), .ZN(n3243)
         );
  OAI21_X1 U4063 ( .B1(n2615), .B2(n4391), .A(n3243), .ZN(n3244) );
  AOI21_X1 U4064 ( .B1(n3245), .B2(n4393), .A(n3244), .ZN(n4717) );
  MUX2_X1 U4065 ( .A(n4717), .B(n3004), .S(n4684), .Z(n3249) );
  AOI21_X1 U4066 ( .B1(n3247), .B2(n3246), .A(n2050), .ZN(n4720) );
  AOI22_X1 U4067 ( .A1(n4720), .A2(n4358), .B1(n3498), .B2(n4678), .ZN(n3248)
         );
  OAI211_X1 U4068 ( .C1(n4344), .C2(n4716), .A(n3249), .B(n3248), .ZN(U3285)
         );
  MUX2_X1 U4069 ( .A(n3250), .B(REG2_REG_2__SCAN_IN), .S(n4684), .Z(n3251) );
  INV_X1 U4070 ( .A(n3251), .ZN(n3254) );
  AOI22_X1 U4071 ( .A1(n4680), .A2(n3252), .B1(REG3_REG_2__SCAN_IN), .B2(n4678), .ZN(n3253) );
  OAI211_X1 U4072 ( .C1(n4450), .C2(n3255), .A(n3254), .B(n3253), .ZN(U3288)
         );
  INV_X1 U4073 ( .A(n3317), .ZN(n3257) );
  NOR2_X1 U4074 ( .A1(n3257), .A2(n3316), .ZN(n3258) );
  XNOR2_X1 U4075 ( .A(n3256), .B(n3258), .ZN(n3263) );
  AOI22_X1 U4076 ( .A1(n3701), .A2(n2367), .B1(n3700), .B2(n3298), .ZN(n3260)
         );
  OAI211_X1 U4077 ( .C1(n3396), .C2(n3703), .A(n3260), .B(n3259), .ZN(n3261)
         );
  AOI21_X1 U4078 ( .B1(n3299), .B2(n3705), .A(n3261), .ZN(n3262) );
  OAI21_X1 U4079 ( .B1(n3263), .B2(n3707), .A(n3262), .ZN(U3218) );
  XOR2_X1 U4080 ( .A(n3337), .B(REG2_REG_10__SCAN_IN), .Z(n3275) );
  NAND2_X1 U4081 ( .A1(U3149), .A2(REG3_REG_10__SCAN_IN), .ZN(n3367) );
  NAND2_X1 U4082 ( .A1(n4660), .A2(ADDR_REG_10__SCAN_IN), .ZN(n3267) );
  OAI211_X1 U4083 ( .C1(n4673), .C2(n3334), .A(n3367), .B(n3267), .ZN(n3274)
         );
  INV_X1 U4084 ( .A(n3271), .ZN(n3272) );
  AOI211_X1 U4085 ( .C1(n3272), .C2(n2115), .A(n4657), .B(n3343), .ZN(n3273)
         );
  AOI211_X1 U4086 ( .C1(n3275), .C2(n4670), .A(n3274), .B(n3273), .ZN(n3276)
         );
  INV_X1 U4087 ( .A(n3276), .ZN(U3250) );
  OAI22_X1 U4088 ( .A1(n3292), .A2(n4436), .B1(n3277), .B2(n4434), .ZN(n3281)
         );
  AND2_X1 U4089 ( .A1(n3799), .A2(n3810), .ZN(n3762) );
  XOR2_X1 U4090 ( .A(n3762), .B(n3278), .Z(n3279) );
  NOR2_X1 U4091 ( .A1(n3279), .A2(n4442), .ZN(n3280) );
  AOI211_X1 U4092 ( .C1(n4439), .C2(n3282), .A(n3281), .B(n3280), .ZN(n3325)
         );
  XOR2_X1 U4093 ( .A(n3283), .B(n3762), .Z(n3326) );
  INV_X1 U4094 ( .A(n3326), .ZN(n3289) );
  OAI21_X1 U4095 ( .B1(n2050), .B2(n3285), .A(n3284), .ZN(n3330) );
  AOI22_X1 U4096 ( .A1(n4431), .A2(REG2_REG_6__SCAN_IN), .B1(n3286), .B2(n4678), .ZN(n3287) );
  OAI21_X1 U4097 ( .B1(n3330), .B2(n4450), .A(n3287), .ZN(n3288) );
  AOI21_X1 U4098 ( .B1(n3289), .B2(n4452), .A(n3288), .ZN(n3290) );
  OAI21_X1 U4099 ( .B1(n3325), .B2(n4431), .A(n3290), .ZN(U3284) );
  AND2_X1 U4100 ( .A1(n3805), .A2(n3803), .ZN(n3749) );
  XNOR2_X1 U4101 ( .A(n3291), .B(n3749), .ZN(n3295) );
  OAI22_X1 U4102 ( .A1(n3292), .A2(n4434), .B1(n3396), .B2(n4436), .ZN(n3293)
         );
  AOI21_X1 U4103 ( .B1(n3298), .B2(n4439), .A(n3293), .ZN(n3294) );
  OAI21_X1 U4104 ( .B1(n3295), .B2(n4442), .A(n3294), .ZN(n3352) );
  INV_X1 U4105 ( .A(n3352), .ZN(n3304) );
  XNOR2_X1 U4106 ( .A(n3296), .B(n3749), .ZN(n3353) );
  AOI21_X1 U4107 ( .B1(n3298), .B2(n3297), .A(n2051), .ZN(n3355) );
  INV_X1 U4108 ( .A(n3355), .ZN(n3301) );
  AOI22_X1 U4109 ( .A1(n4431), .A2(REG2_REG_8__SCAN_IN), .B1(n3299), .B2(n4678), .ZN(n3300) );
  OAI21_X1 U4110 ( .B1(n3301), .B2(n4450), .A(n3300), .ZN(n3302) );
  AOI21_X1 U4111 ( .B1(n3353), .B2(n4452), .A(n3302), .ZN(n3303) );
  OAI21_X1 U4112 ( .B1(n3304), .B2(n4431), .A(n3303), .ZN(U3282) );
  INV_X1 U4113 ( .A(DATAO_REG_25__SCAN_IN), .ZN(n3980) );
  NAND2_X1 U4114 ( .A1(n4217), .A2(U4043), .ZN(n3305) );
  OAI21_X1 U4115 ( .B1(U4043), .B2(n3980), .A(n3305), .ZN(U3575) );
  XOR2_X1 U4116 ( .A(n3307), .B(n3306), .Z(n3308) );
  XNOR2_X1 U4117 ( .A(n3309), .B(n3308), .ZN(n3314) );
  AOI22_X1 U4118 ( .A1(n3310), .A2(n3700), .B1(n3691), .B2(n4012), .ZN(n3311)
         );
  NAND2_X1 U4119 ( .A1(U3149), .A2(REG3_REG_11__SCAN_IN), .ZN(n3347) );
  OAI211_X1 U4120 ( .C1(n3386), .C2(n3655), .A(n3311), .B(n3347), .ZN(n3312)
         );
  AOI21_X1 U4121 ( .B1(n3422), .B2(n3705), .A(n3312), .ZN(n3313) );
  OAI21_X1 U4122 ( .B1(n3314), .B2(n3707), .A(n3313), .ZN(U3233) );
  OR2_X1 U4123 ( .A1(n3256), .A2(n3316), .ZN(n3373) );
  NAND2_X1 U4124 ( .A1(n3373), .A2(n3317), .ZN(n3318) );
  XOR2_X1 U4125 ( .A(n3315), .B(n3318), .Z(n3324) );
  AOI22_X1 U4126 ( .A1(n3701), .A2(n3319), .B1(n3700), .B2(n3389), .ZN(n3321)
         );
  OAI211_X1 U4127 ( .C1(n3386), .C2(n3703), .A(n3321), .B(n3320), .ZN(n3322)
         );
  AOI21_X1 U4128 ( .B1(n3448), .B2(n3705), .A(n3322), .ZN(n3323) );
  OAI21_X1 U4129 ( .B1(n3324), .B2(n3707), .A(n3323), .ZN(U3228) );
  OAI21_X1 U4130 ( .B1(n4715), .B2(n3326), .A(n3325), .ZN(n3332) );
  INV_X1 U4131 ( .A(REG0_REG_6__SCAN_IN), .ZN(n3992) );
  OAI22_X1 U4132 ( .A1(n3330), .A2(n4606), .B1(n4731), .B2(n3992), .ZN(n3327)
         );
  AOI21_X1 U4133 ( .B1(n3332), .B2(n4731), .A(n3327), .ZN(n3328) );
  INV_X1 U4134 ( .A(n3328), .ZN(U3479) );
  INV_X1 U4135 ( .A(REG1_REG_6__SCAN_IN), .ZN(n3329) );
  OAI22_X1 U4136 ( .A1(n3330), .A2(n4540), .B1(n4741), .B2(n3329), .ZN(n3331)
         );
  AOI21_X1 U4137 ( .B1(n3332), .B2(n4741), .A(n3331), .ZN(n3333) );
  INV_X1 U4138 ( .A(n3333), .ZN(U3524) );
  INV_X1 U4139 ( .A(n3334), .ZN(n4617) );
  INV_X1 U4140 ( .A(REG2_REG_11__SCAN_IN), .ZN(n3338) );
  MUX2_X1 U4141 ( .A(n3338), .B(REG2_REG_11__SCAN_IN), .S(n4616), .Z(n3339) );
  AOI211_X1 U4142 ( .C1(n3340), .C2(n3339), .A(n3470), .B(n3428), .ZN(n3351)
         );
  AND2_X1 U4143 ( .A1(n3341), .A2(n4617), .ZN(n3342) );
  XNOR2_X1 U4144 ( .A(n4616), .B(REG1_REG_11__SCAN_IN), .ZN(n3344) );
  AOI211_X1 U4145 ( .C1(n3345), .C2(n3344), .A(n4657), .B(n3434), .ZN(n3350)
         );
  INV_X1 U4146 ( .A(n4616), .ZN(n3348) );
  NAND2_X1 U4147 ( .A1(n4660), .A2(ADDR_REG_11__SCAN_IN), .ZN(n3346) );
  OAI211_X1 U4148 ( .C1(n4673), .C2(n3348), .A(n3347), .B(n3346), .ZN(n3349)
         );
  OR3_X1 U4149 ( .A1(n3351), .A2(n3350), .A3(n3349), .ZN(U3251) );
  AOI21_X1 U4150 ( .B1(n3353), .B2(n4724), .A(n3352), .ZN(n3357) );
  AOI22_X1 U4151 ( .A1(n3355), .A2(n2716), .B1(REG0_REG_8__SCAN_IN), .B2(n4729), .ZN(n3354) );
  OAI21_X1 U4152 ( .B1(n3357), .B2(n4729), .A(n3354), .ZN(U3483) );
  AOI22_X1 U4153 ( .A1(n3355), .A2(n2707), .B1(REG1_REG_8__SCAN_IN), .B2(n2712), .ZN(n3356) );
  OAI21_X1 U4154 ( .B1(n3357), .B2(n2712), .A(n3356), .ZN(U3526) );
  INV_X1 U4155 ( .A(n3358), .ZN(n3360) );
  NOR2_X1 U4156 ( .A1(n3360), .A2(n3359), .ZN(n3361) );
  XNOR2_X1 U4157 ( .A(n3362), .B(n3361), .ZN(n3366) );
  AOI22_X1 U4158 ( .A1(n4440), .A2(n3700), .B1(n3691), .B2(n4387), .ZN(n3363)
         );
  NAND2_X1 U4159 ( .A1(U3149), .A2(REG3_REG_12__SCAN_IN), .ZN(n3431) );
  OAI211_X1 U4160 ( .C1(n4435), .C2(n3655), .A(n3363), .B(n3431), .ZN(n3364)
         );
  AOI21_X1 U4161 ( .B1(n4448), .B2(n3705), .A(n3364), .ZN(n3365) );
  OAI21_X1 U4162 ( .B1(n3366), .B2(n3707), .A(n3365), .ZN(U3221) );
  AOI22_X1 U4163 ( .A1(n3398), .A2(n3700), .B1(n3691), .B2(n4013), .ZN(n3368)
         );
  OAI211_X1 U4164 ( .C1(n3396), .C2(n3655), .A(n3368), .B(n3367), .ZN(n3379)
         );
  NAND2_X1 U4165 ( .A1(n3373), .A2(n3369), .ZN(n3371) );
  AND2_X1 U4166 ( .A1(n3371), .A2(n3370), .ZN(n3376) );
  NAND2_X1 U4167 ( .A1(n3373), .A2(n3372), .ZN(n3375) );
  AOI211_X1 U4168 ( .C1(n3377), .C2(n3376), .A(n3707), .B(n2043), .ZN(n3378)
         );
  AOI211_X1 U4169 ( .C1(n3406), .C2(n3705), .A(n3379), .B(n3378), .ZN(n3380)
         );
  INV_X1 U4170 ( .A(n3380), .ZN(U3214) );
  OAI21_X1 U4171 ( .B1(n2051), .B2(n3382), .A(n3381), .ZN(n3450) );
  INV_X1 U4172 ( .A(n3383), .ZN(n3819) );
  XOR2_X1 U4173 ( .A(n3384), .B(n3751), .Z(n3454) );
  XNOR2_X1 U4174 ( .A(n3385), .B(n3751), .ZN(n3391) );
  OAI22_X1 U4175 ( .A1(n3387), .A2(n4434), .B1(n3386), .B2(n4436), .ZN(n3388)
         );
  AOI21_X1 U4176 ( .B1(n3389), .B2(n4439), .A(n3388), .ZN(n3390) );
  OAI21_X1 U4177 ( .B1(n3391), .B2(n4442), .A(n3390), .ZN(n3451) );
  AOI21_X1 U4178 ( .B1(n3454), .B2(n4724), .A(n3451), .ZN(n3393) );
  MUX2_X1 U4179 ( .A(n3952), .B(n3393), .S(n4741), .Z(n3392) );
  OAI21_X1 U4180 ( .B1(n4540), .B2(n3450), .A(n3392), .ZN(U3527) );
  INV_X1 U4181 ( .A(REG0_REG_9__SCAN_IN), .ZN(n3885) );
  MUX2_X1 U4182 ( .A(n3885), .B(n3393), .S(n4731), .Z(n3394) );
  OAI21_X1 U4183 ( .B1(n3450), .B2(n4606), .A(n3394), .ZN(U3485) );
  XOR2_X1 U4184 ( .A(n3395), .B(n3761), .Z(n3400) );
  OAI22_X1 U4185 ( .A1(n3396), .A2(n4434), .B1(n4435), .B2(n4436), .ZN(n3397)
         );
  AOI21_X1 U4186 ( .B1(n3398), .B2(n4439), .A(n3397), .ZN(n3399) );
  OAI21_X1 U4187 ( .B1(n3400), .B2(n4442), .A(n3399), .ZN(n3472) );
  INV_X1 U4188 ( .A(n3472), .ZN(n3410) );
  XOR2_X1 U4189 ( .A(n3761), .B(n3401), .Z(n3473) );
  INV_X1 U4190 ( .A(n3381), .ZN(n3405) );
  INV_X1 U4191 ( .A(n3402), .ZN(n3403) );
  OAI21_X1 U4192 ( .B1(n3405), .B2(n3404), .A(n3403), .ZN(n3478) );
  AOI22_X1 U4193 ( .A1(n4431), .A2(REG2_REG_10__SCAN_IN), .B1(n3406), .B2(
        n4678), .ZN(n3407) );
  OAI21_X1 U4194 ( .B1(n3478), .B2(n4450), .A(n3407), .ZN(n3408) );
  AOI21_X1 U4195 ( .B1(n3473), .B2(n4452), .A(n3408), .ZN(n3409) );
  OAI21_X1 U4196 ( .B1(n3410), .B2(n4431), .A(n3409), .ZN(U3280) );
  XNOR2_X1 U4197 ( .A(n3411), .B(n3753), .ZN(n3418) );
  OAI21_X1 U4198 ( .B1(n3413), .B2(n3753), .A(n3412), .ZN(n4537) );
  AOI22_X1 U4199 ( .A1(n4014), .A2(n4386), .B1(n4388), .B2(n4012), .ZN(n3414)
         );
  OAI21_X1 U4200 ( .B1(n3420), .B2(n4391), .A(n3414), .ZN(n3415) );
  AOI21_X1 U4201 ( .B1(n4537), .B2(n3416), .A(n3415), .ZN(n3417) );
  OAI21_X1 U4202 ( .B1(n4442), .B2(n3418), .A(n3417), .ZN(n4536) );
  INV_X1 U4203 ( .A(n4536), .ZN(n3426) );
  NOR2_X1 U4204 ( .A1(n3402), .A2(n3420), .ZN(n3421) );
  OR2_X1 U4205 ( .A1(n3419), .A2(n3421), .ZN(n4607) );
  AOI22_X1 U4206 ( .A1(n4431), .A2(REG2_REG_11__SCAN_IN), .B1(n3422), .B2(
        n4678), .ZN(n3423) );
  OAI21_X1 U4207 ( .B1(n4607), .B2(n4450), .A(n3423), .ZN(n3424) );
  AOI21_X1 U4208 ( .B1(n4537), .B2(n4680), .A(n3424), .ZN(n3425) );
  OAI21_X1 U4209 ( .B1(n3426), .B2(n4431), .A(n3425), .ZN(U3279) );
  XOR2_X1 U4210 ( .A(REG2_REG_12__SCAN_IN), .B(n3457), .Z(n3439) );
  NAND2_X1 U4211 ( .A1(n4660), .A2(ADDR_REG_12__SCAN_IN), .ZN(n3430) );
  OAI211_X1 U4212 ( .C1(n4673), .C2(n3429), .A(n3431), .B(n3430), .ZN(n3432)
         );
  INV_X1 U4213 ( .A(n3432), .ZN(n3438) );
  XNOR2_X1 U4214 ( .A(n3464), .B(n3435), .ZN(n3436) );
  NAND2_X1 U4215 ( .A1(n3436), .A2(REG1_REG_12__SCAN_IN), .ZN(n3463) );
  OAI211_X1 U4216 ( .C1(n3436), .C2(REG1_REG_12__SCAN_IN), .A(n3463), .B(n4654), .ZN(n3437) );
  OAI211_X1 U4217 ( .C1(n3439), .C2(n3470), .A(n3438), .B(n3437), .ZN(U3252)
         );
  XOR2_X1 U4218 ( .A(n3441), .B(n3440), .Z(n3442) );
  XNOR2_X1 U4219 ( .A(n3443), .B(n3442), .ZN(n3447) );
  AOI22_X1 U4220 ( .A1(n4424), .A2(n3700), .B1(n3691), .B2(n4011), .ZN(n3444)
         );
  NAND2_X1 U4221 ( .A1(U3149), .A2(REG3_REG_13__SCAN_IN), .ZN(n3460) );
  OAI211_X1 U4222 ( .C1(n4413), .C2(n3655), .A(n3444), .B(n3460), .ZN(n3445)
         );
  AOI21_X1 U4223 ( .B1(n4427), .B2(n3705), .A(n3445), .ZN(n3446) );
  OAI21_X1 U4224 ( .B1(n3447), .B2(n3707), .A(n3446), .ZN(U3231) );
  INV_X1 U4225 ( .A(n3448), .ZN(n3449) );
  OAI22_X1 U4226 ( .A1(n3450), .A2(n4450), .B1(n3449), .B2(n4360), .ZN(n3453)
         );
  MUX2_X1 U4227 ( .A(REG2_REG_9__SCAN_IN), .B(n3451), .S(n4682), .Z(n3452) );
  AOI211_X1 U4228 ( .C1(n3454), .C2(n4452), .A(n3453), .B(n3452), .ZN(n3455)
         );
  INV_X1 U4229 ( .A(n3455), .ZN(U3281) );
  INV_X1 U4230 ( .A(REG2_REG_12__SCAN_IN), .ZN(n3456) );
  INV_X1 U4231 ( .A(REG2_REG_13__SCAN_IN), .ZN(n3458) );
  NOR2_X1 U4232 ( .A1(n4044), .A2(n3458), .ZN(n4045) );
  AOI21_X1 U4233 ( .B1(n3458), .B2(n4044), .A(n4045), .ZN(n3459) );
  XNOR2_X1 U4234 ( .A(n4046), .B(n3459), .ZN(n3471) );
  INV_X1 U4235 ( .A(n3460), .ZN(n3462) );
  NOR2_X1 U4236 ( .A1(n4673), .A2(n4044), .ZN(n3461) );
  AOI211_X1 U4237 ( .C1(n4660), .C2(ADDR_REG_13__SCAN_IN), .A(n3462), .B(n3461), .ZN(n3469) );
  XNOR2_X1 U4238 ( .A(n4044), .B(REG1_REG_13__SCAN_IN), .ZN(n3467) );
  OAI21_X1 U4239 ( .B1(n3464), .B2(n3429), .A(n3463), .ZN(n3466) );
  INV_X1 U4240 ( .A(n4051), .ZN(n3465) );
  OAI211_X1 U4241 ( .C1(n3467), .C2(n3466), .A(n3465), .B(n4654), .ZN(n3468)
         );
  OAI211_X1 U4242 ( .C1(n3471), .C2(n3470), .A(n3469), .B(n3468), .ZN(U3253)
         );
  INV_X1 U4243 ( .A(REG0_REG_10__SCAN_IN), .ZN(n3474) );
  AOI21_X1 U4244 ( .B1(n4724), .B2(n3473), .A(n3472), .ZN(n3476) );
  MUX2_X1 U4245 ( .A(n3474), .B(n3476), .S(n4731), .Z(n3475) );
  OAI21_X1 U4246 ( .B1(n3478), .B2(n4606), .A(n3475), .ZN(U3487) );
  MUX2_X1 U4247 ( .A(n2115), .B(n3476), .S(n4741), .Z(n3477) );
  OAI21_X1 U4248 ( .B1(n4540), .B2(n3478), .A(n3477), .ZN(U3528) );
  NAND2_X1 U4249 ( .A1(n4179), .A2(n3479), .ZN(n4265) );
  NAND2_X1 U4250 ( .A1(n4265), .A2(n3744), .ZN(n4226) );
  NAND2_X1 U4251 ( .A1(n4249), .A2(n3480), .ZN(n3484) );
  NAND2_X1 U4252 ( .A1(n3484), .A2(n3483), .ZN(n3485) );
  OAI21_X1 U4253 ( .B1(n3486), .B2(n3742), .A(n3743), .ZN(n4233) );
  XNOR2_X1 U4254 ( .A(n4233), .B(n4232), .ZN(n3489) );
  AOI22_X1 U4255 ( .A1(n3663), .A2(n4386), .B1(n3491), .B2(n4439), .ZN(n3487)
         );
  OAI21_X1 U4256 ( .B1(n4215), .B2(n4436), .A(n3487), .ZN(n3488) );
  AOI21_X1 U4257 ( .B1(n3489), .B2(n4393), .A(n3488), .ZN(n4494) );
  INV_X1 U4258 ( .A(n4494), .ZN(n3496) );
  INV_X1 U4259 ( .A(n3490), .ZN(n4492) );
  NAND2_X1 U4260 ( .A1(n2041), .A2(n3491), .ZN(n4491) );
  AND3_X1 U4261 ( .A1(n4492), .A2(n4358), .A3(n4491), .ZN(n3495) );
  INV_X1 U4262 ( .A(n3492), .ZN(n3668) );
  OAI22_X1 U4263 ( .A1(n3668), .A2(n4360), .B1(n3493), .B2(n4682), .ZN(n3494)
         );
  AOI211_X1 U4264 ( .C1(n3496), .C2(n4682), .A(n3495), .B(n3494), .ZN(n3497)
         );
  OAI21_X1 U4265 ( .B1(n4495), .B2(n4344), .A(n3497), .ZN(U3268) );
  INV_X1 U4266 ( .A(n3498), .ZN(n3507) );
  OAI211_X1 U4267 ( .C1(n3499), .C2(n3501), .A(n3500), .B(n3673), .ZN(n3506)
         );
  OAI22_X1 U4268 ( .A1(n3677), .A2(n2615), .B1(n3502), .B2(n3655), .ZN(n3503)
         );
  AOI211_X1 U4269 ( .C1(n3691), .C2(n4015), .A(n3504), .B(n3503), .ZN(n3505)
         );
  OAI211_X1 U4270 ( .C1(n3689), .C2(n3507), .A(n3506), .B(n3505), .ZN(U3224)
         );
  OAI22_X1 U4271 ( .A1(n4236), .A2(n3557), .B1(n3556), .B2(n2702), .ZN(n3513)
         );
  OAI22_X1 U4272 ( .A1(n4236), .A2(n3556), .B1(n3554), .B2(n2702), .ZN(n3511)
         );
  XNOR2_X1 U4273 ( .A(n3511), .B(n3561), .ZN(n3514) );
  XOR2_X1 U4274 ( .A(n3513), .B(n3514), .Z(n3661) );
  OAI22_X1 U4275 ( .A1(n4215), .A2(n3556), .B1(n3554), .B2(n4241), .ZN(n3512)
         );
  XNOR2_X1 U4276 ( .A(n3512), .B(n3533), .ZN(n3516) );
  OAI22_X1 U4277 ( .A1(n4215), .A2(n3557), .B1(n3556), .B2(n4241), .ZN(n3517)
         );
  XNOR2_X1 U4278 ( .A(n3516), .B(n3517), .ZN(n3599) );
  OR2_X1 U4279 ( .A1(n3514), .A2(n3513), .ZN(n3600) );
  INV_X1 U4280 ( .A(n3516), .ZN(n3518) );
  NAND2_X1 U4281 ( .A1(n3518), .A2(n3517), .ZN(n3539) );
  NOR2_X1 U4282 ( .A1(n4214), .A2(n3556), .ZN(n3519) );
  AOI21_X1 U4283 ( .B1(n4238), .B2(n2754), .A(n3519), .ZN(n3549) );
  NAND2_X1 U4284 ( .A1(n3539), .A2(n3549), .ZN(n3540) );
  INV_X1 U4285 ( .A(n3540), .ZN(n3520) );
  NAND2_X1 U4286 ( .A1(n3597), .A2(n3520), .ZN(n3640) );
  OAI22_X1 U4287 ( .A1(n4191), .A2(n3556), .B1(n3554), .B2(n4214), .ZN(n3521)
         );
  XNOR2_X1 U4288 ( .A(n3521), .B(n3561), .ZN(n3643) );
  NAND2_X1 U4289 ( .A1(n4217), .A2(n2741), .ZN(n3523) );
  NAND2_X1 U4290 ( .A1(n2726), .A2(n3527), .ZN(n3522) );
  NAND2_X1 U4291 ( .A1(n3523), .A2(n3522), .ZN(n3524) );
  XNOR2_X1 U4292 ( .A(n3524), .B(n3561), .ZN(n3546) );
  INV_X1 U4293 ( .A(n4217), .ZN(n4163) );
  OAI22_X1 U4294 ( .A1(n4163), .A2(n3557), .B1(n3556), .B2(n4198), .ZN(n3545)
         );
  NAND2_X1 U4295 ( .A1(n3546), .A2(n3545), .ZN(n3543) );
  OAI21_X1 U4296 ( .B1(n3546), .B2(n3545), .A(n3543), .ZN(n3525) );
  XNOR2_X1 U4297 ( .A(n3526), .B(n3525), .ZN(n3532) );
  AOI22_X1 U4298 ( .A1(n3700), .A2(n3527), .B1(REG3_REG_25__SCAN_IN), .B2(
        U3149), .ZN(n3529) );
  NAND2_X1 U4299 ( .A1(n4200), .A2(n3705), .ZN(n3528) );
  OAI211_X1 U4300 ( .C1(n4191), .C2(n3655), .A(n3529), .B(n3528), .ZN(n3530)
         );
  AOI21_X1 U4301 ( .B1(n4193), .B2(n3691), .A(n3530), .ZN(n3531) );
  OAI21_X1 U4302 ( .B1(n3532), .B2(n3707), .A(n3531), .ZN(U3222) );
  OAI22_X1 U4303 ( .A1(n4145), .A2(n3556), .B1(n3554), .B2(n3535), .ZN(n3534)
         );
  XNOR2_X1 U4304 ( .A(n3534), .B(n3533), .ZN(n3537) );
  OAI22_X1 U4305 ( .A1(n4145), .A2(n3557), .B1(n3556), .B2(n3535), .ZN(n3536)
         );
  XNOR2_X1 U4306 ( .A(n3537), .B(n3536), .ZN(n3570) );
  INV_X1 U4307 ( .A(n3570), .ZN(n3538) );
  NAND2_X1 U4308 ( .A1(n3538), .A2(n3673), .ZN(n3576) );
  INV_X1 U4309 ( .A(n3539), .ZN(n3541) );
  OAI21_X1 U4310 ( .B1(n3643), .B2(n3541), .A(n3540), .ZN(n3542) );
  NAND2_X1 U4311 ( .A1(n3597), .A2(n3544), .ZN(n3553) );
  INV_X1 U4312 ( .A(n3643), .ZN(n3550) );
  INV_X1 U4313 ( .A(n3545), .ZN(n3548) );
  AOI21_X1 U4314 ( .B1(n3550), .B2(n3549), .A(n3548), .ZN(n3547) );
  NAND3_X1 U4315 ( .A1(n3550), .A2(n3549), .A3(n3548), .ZN(n3551) );
  OAI22_X1 U4316 ( .A1(n4142), .A2(n3556), .B1(n3554), .B2(n4172), .ZN(n3555)
         );
  XNOR2_X1 U4317 ( .A(n3555), .B(n3561), .ZN(n3559) );
  OAI22_X1 U4318 ( .A1(n4142), .A2(n3557), .B1(n3556), .B2(n4172), .ZN(n3558)
         );
  NAND2_X1 U4319 ( .A1(n3559), .A2(n3558), .ZN(n3682) );
  NOR2_X1 U4320 ( .A1(n3559), .A2(n3558), .ZN(n3681) );
  AOI21_X2 U4321 ( .B1(n3685), .B2(n3682), .A(n3681), .ZN(n3582) );
  AOI22_X1 U4322 ( .A1(n4165), .A2(n2754), .B1(n3560), .B2(n3845), .ZN(n3563)
         );
  AOI22_X1 U4323 ( .A1(n4165), .A2(n3560), .B1(n2726), .B2(n3845), .ZN(n3562)
         );
  XNOR2_X1 U4324 ( .A(n3562), .B(n3561), .ZN(n3564) );
  NAND2_X1 U4325 ( .A1(n3582), .A2(n3581), .ZN(n3575) );
  OR2_X1 U4326 ( .A1(n3564), .A2(n3563), .ZN(n3569) );
  NAND2_X1 U4327 ( .A1(n3575), .A2(n3566), .ZN(n3574) );
  NAND2_X1 U4328 ( .A1(n3873), .A2(n3691), .ZN(n3568) );
  AOI22_X1 U4329 ( .A1(n3700), .A2(n4110), .B1(REG3_REG_28__SCAN_IN), .B2(
        U3149), .ZN(n3567) );
  OAI211_X1 U4330 ( .C1(n3689), .C2(n4132), .A(n3568), .B(n3567), .ZN(n3572)
         );
  NOR3_X1 U4331 ( .A1(n3570), .A2(n3707), .A3(n3569), .ZN(n3571) );
  AOI211_X1 U4332 ( .C1(n3701), .C2(n4165), .A(n3572), .B(n3571), .ZN(n3573)
         );
  OAI211_X1 U4333 ( .C1(n3576), .C2(n3575), .A(n3574), .B(n3573), .ZN(U3217)
         );
  NAND3_X1 U4334 ( .A1(n3577), .A2(IR_REG_31__SCAN_IN), .A3(STATE_REG_SCAN_IN), 
        .ZN(n3579) );
  INV_X1 U4335 ( .A(DATAI_31_), .ZN(n3578) );
  OAI22_X1 U4336 ( .A1(n3580), .A2(n3579), .B1(STATE_REG_SCAN_IN), .B2(n3578), 
        .ZN(U3321) );
  XNOR2_X1 U4337 ( .A(n3582), .B(n3581), .ZN(n3587) );
  AOI22_X1 U4338 ( .A1(n3700), .A2(n3845), .B1(REG3_REG_27__SCAN_IN), .B2(
        U3149), .ZN(n3584) );
  NAND2_X1 U4339 ( .A1(n4150), .A2(n3705), .ZN(n3583) );
  OAI211_X1 U4340 ( .C1(n4142), .C2(n3655), .A(n3584), .B(n3583), .ZN(n3585)
         );
  AOI21_X1 U4341 ( .B1(n4111), .B2(n3691), .A(n3585), .ZN(n3586) );
  OAI21_X1 U4342 ( .B1(n3587), .B2(n3707), .A(n3586), .ZN(U3211) );
  INV_X1 U4343 ( .A(n3588), .ZN(n3621) );
  NOR2_X1 U4344 ( .A1(n3621), .A2(n3589), .ZN(n3590) );
  XNOR2_X1 U4345 ( .A(n3591), .B(n3590), .ZN(n3596) );
  AOI22_X1 U4346 ( .A1(n3592), .A2(n3700), .B1(n3691), .B2(n4389), .ZN(n3593)
         );
  NAND2_X1 U4347 ( .A1(U3149), .A2(REG3_REG_14__SCAN_IN), .ZN(n4048) );
  OAI211_X1 U4348 ( .C1(n4437), .C2(n3655), .A(n3593), .B(n4048), .ZN(n3594)
         );
  AOI21_X1 U4349 ( .B1(n4401), .B2(n3705), .A(n3594), .ZN(n3595) );
  OAI21_X1 U4350 ( .B1(n3596), .B2(n3707), .A(n3595), .ZN(U3212) );
  INV_X1 U4351 ( .A(n3597), .ZN(n3602) );
  AOI21_X1 U4352 ( .B1(n3598), .B2(n3600), .A(n3599), .ZN(n3601) );
  OR3_X1 U4353 ( .A1(n3602), .A2(n3601), .A3(n3707), .ZN(n3606) );
  AOI22_X1 U4354 ( .A1(n4254), .A2(n3701), .B1(REG3_REG_23__SCAN_IN), .B2(
        U3149), .ZN(n3603) );
  OAI21_X1 U4355 ( .B1(n3677), .B2(n4241), .A(n3603), .ZN(n3604) );
  AOI21_X1 U4356 ( .B1(n3691), .B2(n4238), .A(n3604), .ZN(n3605) );
  OAI211_X1 U4357 ( .C1(n3689), .C2(n4244), .A(n3606), .B(n3605), .ZN(U3213)
         );
  INV_X1 U4358 ( .A(n3607), .ZN(n3669) );
  INV_X1 U4359 ( .A(n3672), .ZN(n3608) );
  OAI21_X1 U4360 ( .B1(n3608), .B2(n3607), .A(n3670), .ZN(n3609) );
  OAI21_X1 U4361 ( .B1(n3669), .B2(n3672), .A(n3609), .ZN(n3613) );
  NOR2_X1 U4362 ( .A1(n3611), .A2(n3610), .ZN(n3612) );
  XNOR2_X1 U4363 ( .A(n3613), .B(n3612), .ZN(n3619) );
  INV_X1 U4364 ( .A(n4303), .ZN(n3617) );
  AOI22_X1 U4365 ( .A1(n4333), .A2(n3701), .B1(n3700), .B2(n3614), .ZN(n3615)
         );
  NAND2_X1 U4366 ( .A1(U3149), .A2(REG3_REG_19__SCAN_IN), .ZN(n4087) );
  OAI211_X1 U4367 ( .C1(n4252), .C2(n3703), .A(n3615), .B(n4087), .ZN(n3616)
         );
  AOI21_X1 U4368 ( .B1(n3617), .B2(n3705), .A(n3616), .ZN(n3618) );
  OAI21_X1 U4369 ( .B1(n3619), .B2(n3707), .A(n3618), .ZN(U3216) );
  INV_X1 U4370 ( .A(n3620), .ZN(n3697) );
  NOR2_X1 U4371 ( .A1(n2027), .A2(n3621), .ZN(n3623) );
  NAND2_X1 U4372 ( .A1(n3623), .A2(n3622), .ZN(n3695) );
  NOR2_X1 U4373 ( .A1(n3623), .A2(n3622), .ZN(n3694) );
  AOI21_X1 U4374 ( .B1(n3697), .B2(n3695), .A(n3694), .ZN(n3627) );
  NOR2_X1 U4375 ( .A1(n3625), .A2(n3624), .ZN(n3626) );
  XNOR2_X1 U4376 ( .A(n3627), .B(n3626), .ZN(n3631) );
  AOI22_X1 U4377 ( .A1(n3701), .A2(n4389), .B1(n3700), .B2(n4356), .ZN(n3628)
         );
  NAND2_X1 U4378 ( .A1(U3149), .A2(REG3_REG_16__SCAN_IN), .ZN(n4068) );
  OAI211_X1 U4379 ( .C1(n2484), .C2(n3703), .A(n3628), .B(n4068), .ZN(n3629)
         );
  AOI21_X1 U4380 ( .B1(n4359), .B2(n3705), .A(n3629), .ZN(n3630) );
  OAI21_X1 U4381 ( .B1(n3631), .B2(n3707), .A(n3630), .ZN(U3223) );
  NAND2_X1 U4382 ( .A1(n2155), .A2(n3633), .ZN(n3634) );
  XNOR2_X1 U4383 ( .A(n3635), .B(n3634), .ZN(n3636) );
  NAND2_X1 U4384 ( .A1(n3636), .A2(n3673), .ZN(n3639) );
  AND2_X1 U4385 ( .A1(U3149), .A2(REG3_REG_17__SCAN_IN), .ZN(n4645) );
  OAI22_X1 U4386 ( .A1(n3677), .A2(n2483), .B1(n3703), .B2(n4295), .ZN(n3637)
         );
  AOI211_X1 U4387 ( .C1(n3701), .C2(n2469), .A(n4645), .B(n3637), .ZN(n3638)
         );
  OAI211_X1 U4388 ( .C1(n3689), .C2(n4339), .A(n3639), .B(n3638), .ZN(U3225)
         );
  INV_X1 U4389 ( .A(n3640), .ZN(n3642) );
  NOR2_X1 U4390 ( .A1(n3642), .A2(n3641), .ZN(n3644) );
  XNOR2_X1 U4391 ( .A(n3644), .B(n3643), .ZN(n3650) );
  OAI22_X1 U4392 ( .A1(n3677), .A2(n4214), .B1(STATE_REG_SCAN_IN), .B2(n3645), 
        .ZN(n3647) );
  NOR2_X1 U4393 ( .A1(n4215), .A2(n3655), .ZN(n3646) );
  AOI211_X1 U4394 ( .C1(n3691), .C2(n4217), .A(n3647), .B(n3646), .ZN(n3649)
         );
  NAND2_X1 U4395 ( .A1(n4220), .A2(n3705), .ZN(n3648) );
  OAI211_X1 U4396 ( .C1(n3650), .C2(n3707), .A(n3649), .B(n3648), .ZN(U3226)
         );
  NAND2_X1 U4397 ( .A1(n2182), .A2(n2184), .ZN(n3652) );
  AOI22_X1 U4398 ( .A1(n3654), .A2(n2184), .B1(n3653), .B2(n3652), .ZN(n3659)
         );
  OAI22_X1 U4399 ( .A1(n4311), .A2(n3655), .B1(STATE_REG_SCAN_IN), .B2(n2058), 
        .ZN(n3657) );
  OAI22_X1 U4400 ( .A1(n4273), .A2(n3703), .B1(n3677), .B2(n4280), .ZN(n3656)
         );
  AOI211_X1 U4401 ( .C1(n4281), .C2(n3705), .A(n3657), .B(n3656), .ZN(n3658)
         );
  OAI21_X1 U4402 ( .B1(n3659), .B2(n3707), .A(n3658), .ZN(U3230) );
  OAI21_X1 U4403 ( .B1(n3661), .B2(n3660), .A(n3598), .ZN(n3662) );
  NAND2_X1 U4404 ( .A1(n3662), .A2(n3673), .ZN(n3667) );
  AOI22_X1 U4405 ( .A1(n3663), .A2(n3701), .B1(REG3_REG_22__SCAN_IN), .B2(
        U3149), .ZN(n3664) );
  OAI21_X1 U4406 ( .B1(n3677), .B2(n2702), .A(n3664), .ZN(n3665) );
  AOI21_X1 U4407 ( .B1(n3874), .B2(n3691), .A(n3665), .ZN(n3666) );
  OAI211_X1 U4408 ( .C1(n3689), .C2(n3668), .A(n3667), .B(n3666), .ZN(U3232)
         );
  XNOR2_X1 U4409 ( .A(n3670), .B(n3669), .ZN(n3671) );
  XNOR2_X1 U4410 ( .A(n3672), .B(n3671), .ZN(n3674) );
  NAND2_X1 U4411 ( .A1(n3674), .A2(n3673), .ZN(n3680) );
  NOR2_X1 U4412 ( .A1(n3675), .A2(STATE_REG_SCAN_IN), .ZN(n4661) );
  OAI22_X1 U4413 ( .A1(n4311), .A2(n3703), .B1(n3677), .B2(n3676), .ZN(n3678)
         );
  AOI211_X1 U4414 ( .C1(n3701), .C2(n4347), .A(n4661), .B(n3678), .ZN(n3679)
         );
  OAI211_X1 U4415 ( .C1(n3689), .C2(n4318), .A(n3680), .B(n3679), .ZN(U3235)
         );
  INV_X1 U4416 ( .A(n3681), .ZN(n3683) );
  NAND2_X1 U4417 ( .A1(n3683), .A2(n3682), .ZN(n3684) );
  XNOR2_X1 U4418 ( .A(n3685), .B(n3684), .ZN(n3693) );
  NAND2_X1 U4419 ( .A1(n4217), .A2(n3701), .ZN(n3688) );
  AOI22_X1 U4420 ( .A1(n3700), .A2(n3686), .B1(REG3_REG_26__SCAN_IN), .B2(
        U3149), .ZN(n3687) );
  OAI211_X1 U4421 ( .C1(n3689), .C2(n4169), .A(n3688), .B(n3687), .ZN(n3690)
         );
  AOI21_X1 U4422 ( .B1(n4165), .B2(n3691), .A(n3690), .ZN(n3692) );
  OAI21_X1 U4423 ( .B1(n3693), .B2(n3707), .A(n3692), .ZN(U3237) );
  INV_X1 U4424 ( .A(n3694), .ZN(n3696) );
  NAND2_X1 U4425 ( .A1(n3696), .A2(n3695), .ZN(n3698) );
  XNOR2_X1 U4426 ( .A(n3698), .B(n3697), .ZN(n3708) );
  INV_X1 U4427 ( .A(n3699), .ZN(n4378) );
  AOI22_X1 U4428 ( .A1(n3701), .A2(n4011), .B1(n3700), .B2(n4373), .ZN(n3702)
         );
  NAND2_X1 U4429 ( .A1(U3149), .A2(REG3_REG_15__SCAN_IN), .ZN(n4641) );
  OAI211_X1 U4430 ( .C1(n4367), .C2(n3703), .A(n3702), .B(n4641), .ZN(n3704)
         );
  AOI21_X1 U4431 ( .B1(n4378), .B2(n3705), .A(n3704), .ZN(n3706) );
  OAI21_X1 U4432 ( .B1(n3708), .B2(n3707), .A(n3706), .ZN(U3238) );
  NAND2_X1 U4433 ( .A1(n3712), .A2(n4368), .ZN(n3823) );
  NAND2_X1 U4434 ( .A1(n3711), .A2(n3710), .ZN(n3808) );
  NAND2_X1 U4435 ( .A1(n3808), .A2(n3712), .ZN(n3824) );
  OAI21_X1 U4436 ( .B1(n3709), .B2(n3823), .A(n3824), .ZN(n3713) );
  AOI211_X1 U4437 ( .C1(n3713), .C2(n3832), .A(n2090), .B(n3831), .ZN(n3715)
         );
  INV_X1 U4438 ( .A(n3714), .ZN(n3836) );
  OAI21_X1 U4439 ( .B1(n3715), .B2(n3836), .A(n3835), .ZN(n3718) );
  INV_X1 U4440 ( .A(n3716), .ZN(n3717) );
  AOI21_X1 U4441 ( .B1(n3718), .B2(n3839), .A(n3717), .ZN(n3719) );
  OR2_X1 U4442 ( .A1(n3738), .A2(n2084), .ZN(n3842) );
  OAI21_X1 U4443 ( .B1(n3719), .B2(n3842), .A(n3841), .ZN(n3725) );
  AND2_X1 U4444 ( .A1(n2024), .A2(n4115), .ZN(n3726) );
  NAND2_X1 U4445 ( .A1(n3722), .A2(DATAI_29_), .ZN(n4093) );
  OR2_X1 U4446 ( .A1(n3873), .A2(n4093), .ZN(n3724) );
  INV_X1 U4447 ( .A(REG2_REG_31__SCAN_IN), .ZN(n3900) );
  NAND2_X1 U4448 ( .A1(n2008), .A2(REG0_REG_31__SCAN_IN), .ZN(n3721) );
  NAND2_X1 U4449 ( .A1(n2009), .A2(REG1_REG_31__SCAN_IN), .ZN(n3720) );
  OAI211_X1 U4450 ( .C1(n2447), .C2(n3900), .A(n3721), .B(n3720), .ZN(n4097)
         );
  NAND2_X1 U4451 ( .A1(n3722), .A2(DATAI_31_), .ZN(n4098) );
  NAND2_X1 U4452 ( .A1(n4097), .A2(n4098), .ZN(n3854) );
  INV_X1 U4453 ( .A(n4120), .ZN(n3723) );
  NAND2_X1 U4454 ( .A1(n3723), .A2(n4102), .ZN(n3765) );
  AND3_X1 U4455 ( .A1(n3724), .A2(n3854), .A3(n3765), .ZN(n3728) );
  NAND4_X1 U4456 ( .A1(n3725), .A2(n3851), .A3(n3726), .A4(n3728), .ZN(n3736)
         );
  INV_X1 U4457 ( .A(n3726), .ZN(n3730) );
  NAND2_X1 U4458 ( .A1(n3873), .A2(n4093), .ZN(n3727) );
  AND2_X1 U4459 ( .A1(n4114), .A2(n3727), .ZN(n3847) );
  INV_X1 U4460 ( .A(n3728), .ZN(n3729) );
  AOI21_X1 U4461 ( .B1(n3730), .B2(n3847), .A(n3729), .ZN(n3852) );
  INV_X1 U4462 ( .A(n3731), .ZN(n3844) );
  NAND3_X1 U4463 ( .A1(n3847), .A2(n4140), .A3(n3844), .ZN(n3734) );
  NOR2_X1 U4464 ( .A1(n4097), .A2(n4098), .ZN(n3856) );
  INV_X1 U4465 ( .A(n4102), .ZN(n3732) );
  NAND2_X1 U4466 ( .A1(n3732), .A2(n4120), .ZN(n3853) );
  NOR2_X1 U4467 ( .A1(n3853), .A2(n4098), .ZN(n3733) );
  AOI211_X1 U4468 ( .C1(n3852), .C2(n3734), .A(n3856), .B(n3733), .ZN(n3735)
         );
  AOI22_X1 U4469 ( .A1(n3736), .A2(n3735), .B1(n4102), .B2(n4098), .ZN(n3864)
         );
  XNOR2_X1 U4470 ( .A(n3873), .B(n4093), .ZN(n4462) );
  INV_X1 U4471 ( .A(n4462), .ZN(n4118) );
  NAND2_X1 U4472 ( .A1(n3844), .A2(n3737), .ZN(n4161) );
  INV_X1 U4473 ( .A(n4187), .ZN(n3739) );
  NAND2_X1 U4474 ( .A1(n3741), .A2(n3740), .ZN(n4235) );
  INV_X1 U4475 ( .A(n4235), .ZN(n3776) );
  INV_X1 U4476 ( .A(n3742), .ZN(n3834) );
  NAND2_X1 U4477 ( .A1(n3834), .A2(n3743), .ZN(n4250) );
  XNOR2_X1 U4478 ( .A(n4271), .B(n4301), .ZN(n4292) );
  NAND2_X1 U4479 ( .A1(n3745), .A2(n3744), .ZN(n4268) );
  INV_X1 U4480 ( .A(n4374), .ZN(n3747) );
  XNOR2_X1 U4481 ( .A(n3746), .B(n4437), .ZN(n4416) );
  AND4_X1 U4482 ( .A1(n4323), .A2(n3748), .A3(n3747), .A4(n4416), .ZN(n3773)
         );
  NAND4_X1 U4483 ( .A1(n3752), .A2(n3751), .A3(n3750), .A4(n3749), .ZN(n3759)
         );
  INV_X1 U4484 ( .A(n3753), .ZN(n3757) );
  NAND4_X1 U4485 ( .A1(n3757), .A2(n3756), .A3(n3755), .A4(n3754), .ZN(n3758)
         );
  NOR2_X1 U4486 ( .A1(n3759), .A2(n3758), .ZN(n3772) );
  INV_X1 U4487 ( .A(n4288), .ZN(n3760) );
  NAND2_X1 U4488 ( .A1(n3760), .A2(n4287), .ZN(n4331) );
  NAND4_X1 U4489 ( .A1(n3763), .A2(n2612), .A3(n3762), .A4(n3761), .ZN(n3770)
         );
  AND2_X1 U4490 ( .A1(n3853), .A2(n3854), .ZN(n3767) );
  INV_X1 U4491 ( .A(n3856), .ZN(n3764) );
  NAND4_X1 U4492 ( .A1(n3767), .A2(n3766), .A3(n3765), .A4(n3764), .ZN(n3769)
         );
  NAND2_X1 U4493 ( .A1(n4411), .A2(n4409), .ZN(n4444) );
  OR2_X1 U4494 ( .A1(n4383), .A2(n4444), .ZN(n3768) );
  NOR4_X1 U4495 ( .A1(n4331), .A2(n3770), .A3(n3769), .A4(n3768), .ZN(n3771)
         );
  NAND4_X1 U4496 ( .A1(n4268), .A2(n3773), .A3(n3772), .A4(n3771), .ZN(n3774)
         );
  NOR3_X1 U4497 ( .A1(n4250), .A2(n4292), .A3(n3774), .ZN(n3775) );
  NAND3_X1 U4498 ( .A1(n3776), .A2(n4232), .A3(n3775), .ZN(n3777) );
  NOR2_X1 U4499 ( .A1(n4211), .A2(n3777), .ZN(n3780) );
  NAND2_X1 U4500 ( .A1(n4159), .A2(n3778), .ZN(n4188) );
  INV_X1 U4501 ( .A(n4188), .ZN(n3779) );
  NAND2_X1 U4502 ( .A1(n3780), .A2(n3779), .ZN(n3781) );
  NOR2_X1 U4503 ( .A1(n4161), .A2(n3781), .ZN(n3782) );
  NAND4_X1 U4504 ( .A1(n3783), .A2(n4140), .A3(n4118), .A4(n3782), .ZN(n3861)
         );
  OAI211_X1 U4505 ( .C1(n3786), .C2(n2644), .A(n3785), .B(n3784), .ZN(n3789)
         );
  NAND3_X1 U4506 ( .A1(n3789), .A2(n3788), .A3(n3787), .ZN(n3792) );
  NAND3_X1 U4507 ( .A1(n3792), .A2(n3791), .A3(n3790), .ZN(n3795) );
  NAND3_X1 U4508 ( .A1(n3795), .A2(n3794), .A3(n3793), .ZN(n3802) );
  INV_X1 U4509 ( .A(n3796), .ZN(n3798) );
  NOR3_X1 U4510 ( .A1(n2072), .A2(n3798), .A3(n3797), .ZN(n3801) );
  AOI211_X1 U4511 ( .C1(n3802), .C2(n3801), .A(n2068), .B(n3800), .ZN(n3807)
         );
  NAND2_X1 U4512 ( .A1(n3804), .A2(n3803), .ZN(n3811) );
  OAI211_X1 U4513 ( .C1(n3807), .C2(n3811), .A(n3806), .B(n3805), .ZN(n3815)
         );
  INV_X1 U4514 ( .A(n3808), .ZN(n3814) );
  NAND2_X1 U4515 ( .A1(n2069), .A2(n3810), .ZN(n3812) );
  OAI21_X1 U4516 ( .B1(n3812), .B2(n3811), .A(n3816), .ZN(n3813) );
  AOI22_X1 U4517 ( .A1(n3815), .A2(n3814), .B1(n3824), .B2(n3813), .ZN(n3822)
         );
  INV_X1 U4518 ( .A(n3816), .ZN(n3820) );
  OAI211_X1 U4519 ( .C1(n3820), .C2(n3819), .A(n3818), .B(n3817), .ZN(n3821)
         );
  NOR2_X1 U4520 ( .A1(n3822), .A2(n3821), .ZN(n3830) );
  INV_X1 U4521 ( .A(n3823), .ZN(n3827) );
  INV_X1 U4522 ( .A(n3824), .ZN(n3825) );
  AOI21_X1 U4523 ( .B1(n3827), .B2(n3826), .A(n3825), .ZN(n3829) );
  OAI21_X1 U4524 ( .B1(n3830), .B2(n3829), .A(n3828), .ZN(n3833) );
  AOI21_X1 U4525 ( .B1(n3833), .B2(n3832), .A(n3831), .ZN(n3837) );
  OAI211_X1 U4526 ( .C1(n3837), .C2(n3836), .A(n3835), .B(n3834), .ZN(n3840)
         );
  AOI21_X1 U4527 ( .B1(n3840), .B2(n3839), .A(n3838), .ZN(n3843) );
  OAI21_X1 U4528 ( .B1(n3843), .B2(n3842), .A(n3841), .ZN(n3850) );
  INV_X1 U4529 ( .A(n4165), .ZN(n3846) );
  OAI21_X1 U4530 ( .B1(n3846), .B2(n3845), .A(n3844), .ZN(n3849) );
  INV_X1 U4531 ( .A(n3847), .ZN(n3848) );
  AOI211_X1 U4532 ( .C1(n3851), .C2(n3850), .A(n3849), .B(n3848), .ZN(n3859)
         );
  INV_X1 U4533 ( .A(n3852), .ZN(n3858) );
  INV_X1 U4534 ( .A(n3853), .ZN(n3855) );
  OAI21_X1 U4535 ( .B1(n3856), .B2(n3855), .A(n3854), .ZN(n3857) );
  OAI21_X1 U4536 ( .B1(n3859), .B2(n3858), .A(n3857), .ZN(n3860) );
  MUX2_X1 U4537 ( .A(n3861), .B(n3860), .S(n2611), .Z(n3862) );
  OAI21_X1 U4538 ( .B1(n3864), .B2(n3863), .A(n3862), .ZN(n3865) );
  XNOR2_X1 U4539 ( .A(n3865), .B(n4611), .ZN(n3872) );
  NOR2_X1 U4540 ( .A1(n3867), .A2(n3866), .ZN(n3870) );
  OAI21_X1 U4541 ( .B1(n3868), .B2(n3871), .A(B_REG_SCAN_IN), .ZN(n3869) );
  OAI22_X1 U4542 ( .A1(n3872), .A2(n3871), .B1(n3870), .B2(n3869), .ZN(U3239)
         );
  MUX2_X1 U4543 ( .A(n4097), .B(DATAO_REG_31__SCAN_IN), .S(n4017), .Z(U3581)
         );
  MUX2_X1 U4544 ( .A(n3873), .B(DATAO_REG_29__SCAN_IN), .S(n4017), .Z(U3579)
         );
  MUX2_X1 U4545 ( .A(n4111), .B(DATAO_REG_28__SCAN_IN), .S(n4017), .Z(U3578)
         );
  MUX2_X1 U4546 ( .A(n4165), .B(DATAO_REG_27__SCAN_IN), .S(n4017), .Z(U3577)
         );
  MUX2_X1 U4547 ( .A(n4193), .B(DATAO_REG_26__SCAN_IN), .S(n4017), .Z(U3576)
         );
  MUX2_X1 U4548 ( .A(n4238), .B(DATAO_REG_24__SCAN_IN), .S(n4017), .Z(U3574)
         );
  MUX2_X1 U4549 ( .A(n3874), .B(DATAO_REG_23__SCAN_IN), .S(n4017), .Z(U3573)
         );
  MUX2_X1 U4550 ( .A(n4254), .B(DATAO_REG_22__SCAN_IN), .S(n4017), .Z(U3572)
         );
  MUX2_X1 U4551 ( .A(n4297), .B(DATAO_REG_20__SCAN_IN), .S(n4017), .Z(U3570)
         );
  MUX2_X1 U4552 ( .A(n4271), .B(DATAO_REG_19__SCAN_IN), .S(n4017), .Z(n4010)
         );
  INV_X1 U4553 ( .A(DATAI_19_), .ZN(n3908) );
  NOR3_X1 U4554 ( .A1(REG1_REG_17__SCAN_IN), .A2(ADDR_REG_16__SCAN_IN), .A3(
        n3908), .ZN(n3878) );
  INV_X1 U4555 ( .A(REG0_REG_3__SCAN_IN), .ZN(n4708) );
  NOR4_X1 U4556 ( .A1(n4066), .A2(n4739), .A3(n4708), .A4(n2295), .ZN(n3877)
         );
  INV_X1 U4557 ( .A(REG2_REG_29__SCAN_IN), .ZN(n3903) );
  NAND4_X1 U4558 ( .A1(DATAI_27_), .A2(REG2_REG_20__SCAN_IN), .A3(DATAI_4_), 
        .A4(n3903), .ZN(n3875) );
  NOR4_X1 U4559 ( .A1(REG3_REG_21__SCAN_IN), .A2(REG2_REG_22__SCAN_IN), .A3(
        n3900), .A4(n3875), .ZN(n3876) );
  NAND4_X1 U4560 ( .A1(ADDR_REG_11__SCAN_IN), .A2(n3878), .A3(n3877), .A4(
        n3876), .ZN(n3898) );
  INV_X1 U4561 ( .A(ADDR_REG_15__SCAN_IN), .ZN(n4643) );
  NOR4_X1 U4562 ( .A1(DATAO_REG_8__SCAN_IN), .A2(ADDR_REG_14__SCAN_IN), .A3(
        DATAO_REG_25__SCAN_IN), .A4(n4643), .ZN(n3879) );
  NAND4_X1 U4563 ( .A1(n3880), .A2(IR_REG_26__SCAN_IN), .A3(n3879), .A4(n3979), 
        .ZN(n3897) );
  OR4_X1 U4564 ( .A1(REG1_REG_22__SCAN_IN), .A2(REG1_REG_18__SCAN_IN), .A3(
        DATAI_1_), .A4(B_REG_SCAN_IN), .ZN(n3894) );
  NOR4_X1 U4565 ( .A1(ADDR_REG_19__SCAN_IN), .A2(REG2_REG_4__SCAN_IN), .A3(
        DATAO_REG_1__SCAN_IN), .A4(n3967), .ZN(n3883) );
  INV_X1 U4566 ( .A(REG2_REG_10__SCAN_IN), .ZN(n3953) );
  INV_X1 U4567 ( .A(REG1_REG_4__SCAN_IN), .ZN(n4735) );
  NOR3_X1 U4568 ( .A1(REG2_REG_6__SCAN_IN), .A2(n3953), .A3(n4735), .ZN(n3882)
         );
  INV_X1 U4569 ( .A(REG1_REG_12__SCAN_IN), .ZN(n4534) );
  NOR4_X1 U4570 ( .A1(IR_REG_16__SCAN_IN), .A2(REG1_REG_5__SCAN_IN), .A3(n4534), .A4(n3952), .ZN(n3881) );
  NAND4_X1 U4571 ( .A1(n3883), .A2(ADDR_REG_8__SCAN_IN), .A3(n3882), .A4(n3881), .ZN(n3893) );
  NOR4_X1 U4572 ( .A1(n3884), .A2(IR_REG_22__SCAN_IN), .A3(IR_REG_11__SCAN_IN), 
        .A4(IR_REG_19__SCAN_IN), .ZN(n3890) );
  INV_X1 U4573 ( .A(DATAI_7_), .ZN(n3923) );
  NAND4_X1 U4574 ( .A1(DATAI_6_), .A2(DATAI_2_), .A3(n3885), .A4(n3923), .ZN(
        n3888) );
  NOR4_X1 U4575 ( .A1(REG0_REG_29__SCAN_IN), .A2(REG1_REG_20__SCAN_IN), .A3(
        REG1_REG_24__SCAN_IN), .A4(REG0_REG_30__SCAN_IN), .ZN(n3886) );
  NAND3_X1 U4576 ( .A1(n3992), .A2(n3958), .A3(n3886), .ZN(n3887) );
  NOR4_X1 U4577 ( .A1(REG3_REG_11__SCAN_IN), .A2(n3888), .A3(DATAI_11_), .A4(
        n3887), .ZN(n3889) );
  NAND3_X1 U4578 ( .A1(n3890), .A2(DATAO_REG_7__SCAN_IN), .A3(n3889), .ZN(
        n3892) );
  NAND4_X1 U4579 ( .A1(REG1_REG_16__SCAN_IN), .A2(REG2_REG_3__SCAN_IN), .A3(
        IR_REG_7__SCAN_IN), .A4(DATAI_8_), .ZN(n3891) );
  OR4_X1 U4580 ( .A1(n3894), .A2(n3893), .A3(n3892), .A4(n3891), .ZN(n3896) );
  OR3_X1 U4581 ( .A1(DATAO_REG_21__SCAN_IN), .A2(ADDR_REG_5__SCAN_IN), .A3(
        n3936), .ZN(n3895) );
  NOR4_X1 U4582 ( .A1(n3898), .A2(n3897), .A3(n3896), .A4(n3895), .ZN(n4008)
         );
  AOI22_X1 U4583 ( .A1(n3900), .A2(keyinput9), .B1(n3493), .B2(keyinput11), 
        .ZN(n3899) );
  OAI221_X1 U4584 ( .B1(n3900), .B2(keyinput9), .C1(n3493), .C2(keyinput11), 
        .A(n3899), .ZN(n3912) );
  INV_X1 U4585 ( .A(DATAI_4_), .ZN(n3902) );
  AOI22_X1 U4586 ( .A1(n3903), .A2(keyinput21), .B1(keyinput16), .B2(n3902), 
        .ZN(n3901) );
  OAI221_X1 U4587 ( .B1(n3903), .B2(keyinput21), .C1(n3902), .C2(keyinput16), 
        .A(n3901), .ZN(n3911) );
  INV_X1 U4588 ( .A(DATAI_27_), .ZN(n3905) );
  AOI22_X1 U4589 ( .A1(n2518), .A2(keyinput14), .B1(n3905), .B2(keyinput7), 
        .ZN(n3904) );
  OAI221_X1 U4590 ( .B1(n2518), .B2(keyinput14), .C1(n3905), .C2(keyinput7), 
        .A(n3904), .ZN(n3910) );
  INV_X1 U4591 ( .A(ADDR_REG_11__SCAN_IN), .ZN(n3907) );
  AOI22_X1 U4592 ( .A1(n3908), .A2(keyinput27), .B1(keyinput47), .B2(n3907), 
        .ZN(n3906) );
  OAI221_X1 U4593 ( .B1(n3908), .B2(keyinput27), .C1(n3907), .C2(keyinput47), 
        .A(n3906), .ZN(n3909) );
  NOR4_X1 U4594 ( .A1(n3912), .A2(n3911), .A3(n3910), .A4(n3909), .ZN(n3950)
         );
  AOI22_X1 U4595 ( .A1(n2295), .A2(keyinput19), .B1(n4708), .B2(keyinput15), 
        .ZN(n3913) );
  OAI221_X1 U4596 ( .B1(n2295), .B2(keyinput19), .C1(n4708), .C2(keyinput15), 
        .A(n3913), .ZN(n3921) );
  AOI22_X1 U4597 ( .A1(n4739), .A2(keyinput0), .B1(n4066), .B2(keyinput10), 
        .ZN(n3914) );
  OAI221_X1 U4598 ( .B1(n4739), .B2(keyinput0), .C1(n4066), .C2(keyinput10), 
        .A(n3914), .ZN(n3920) );
  INV_X1 U4599 ( .A(ADDR_REG_16__SCAN_IN), .ZN(n4070) );
  INV_X1 U4600 ( .A(REG1_REG_17__SCAN_IN), .ZN(n4513) );
  AOI22_X1 U4601 ( .A1(n4070), .A2(keyinput2), .B1(n4513), .B2(keyinput55), 
        .ZN(n3915) );
  OAI221_X1 U4602 ( .B1(n4070), .B2(keyinput2), .C1(n4513), .C2(keyinput55), 
        .A(n3915), .ZN(n3919) );
  XNOR2_X1 U4603 ( .A(REG0_REG_9__SCAN_IN), .B(keyinput5), .ZN(n3917) );
  XNOR2_X1 U4604 ( .A(DATAI_2_), .B(keyinput13), .ZN(n3916) );
  NAND2_X1 U4605 ( .A1(n3917), .A2(n3916), .ZN(n3918) );
  NOR4_X1 U4606 ( .A1(n3921), .A2(n3920), .A3(n3919), .A4(n3918), .ZN(n3949)
         );
  INV_X1 U4607 ( .A(DATAI_6_), .ZN(n3924) );
  AOI22_X1 U4608 ( .A1(n3924), .A2(keyinput1), .B1(n3923), .B2(keyinput35), 
        .ZN(n3922) );
  OAI221_X1 U4609 ( .B1(n3924), .B2(keyinput1), .C1(n3923), .C2(keyinput35), 
        .A(n3922), .ZN(n3932) );
  INV_X1 U4610 ( .A(REG1_REG_20__SCAN_IN), .ZN(n4502) );
  AOI22_X1 U4611 ( .A1(n4502), .A2(keyinput4), .B1(keyinput3), .B2(n4485), 
        .ZN(n3925) );
  OAI221_X1 U4612 ( .B1(n4502), .B2(keyinput4), .C1(n4485), .C2(keyinput3), 
        .A(n3925), .ZN(n3931) );
  XNOR2_X1 U4613 ( .A(IR_REG_11__SCAN_IN), .B(keyinput6), .ZN(n3929) );
  XNOR2_X1 U4614 ( .A(IR_REG_14__SCAN_IN), .B(keyinput18), .ZN(n3928) );
  XNOR2_X1 U4615 ( .A(REG1_REG_16__SCAN_IN), .B(keyinput63), .ZN(n3927) );
  XNOR2_X1 U4616 ( .A(IR_REG_19__SCAN_IN), .B(keyinput8), .ZN(n3926) );
  NAND4_X1 U4617 ( .A1(n3929), .A2(n3928), .A3(n3927), .A4(n3926), .ZN(n3930)
         );
  NOR3_X1 U4618 ( .A1(n3932), .A2(n3931), .A3(n3930), .ZN(n3948) );
  AOI22_X1 U4619 ( .A1(n3934), .A2(keyinput39), .B1(keyinput23), .B2(n4549), 
        .ZN(n3933) );
  OAI221_X1 U4620 ( .B1(n3934), .B2(keyinput39), .C1(n4549), .C2(keyinput23), 
        .A(n3933), .ZN(n3946) );
  AOI22_X1 U4621 ( .A1(n3937), .A2(keyinput17), .B1(keyinput12), .B2(n3936), 
        .ZN(n3935) );
  OAI221_X1 U4622 ( .B1(n3937), .B2(keyinput17), .C1(n3936), .C2(keyinput12), 
        .A(n3935), .ZN(n3945) );
  INV_X1 U4623 ( .A(D_REG_10__SCAN_IN), .ZN(n4687) );
  AOI22_X1 U4624 ( .A1(n4687), .A2(keyinput31), .B1(keyinput51), .B2(n3939), 
        .ZN(n3938) );
  OAI221_X1 U4625 ( .B1(n4687), .B2(keyinput31), .C1(n3939), .C2(keyinput51), 
        .A(n3938), .ZN(n3944) );
  INV_X1 U4626 ( .A(ADDR_REG_5__SCAN_IN), .ZN(n3942) );
  AOI22_X1 U4627 ( .A1(n3942), .A2(keyinput59), .B1(keyinput43), .B2(n3941), 
        .ZN(n3940) );
  OAI221_X1 U4628 ( .B1(n3942), .B2(keyinput59), .C1(n3941), .C2(keyinput43), 
        .A(n3940), .ZN(n3943) );
  NOR4_X1 U4629 ( .A1(n3946), .A2(n3945), .A3(n3944), .A4(n3943), .ZN(n3947)
         );
  NAND4_X1 U4630 ( .A1(n3950), .A2(n3949), .A3(n3948), .A4(n3947), .ZN(n4007)
         );
  AOI22_X1 U4631 ( .A1(n3953), .A2(keyinput50), .B1(keyinput45), .B2(n3952), 
        .ZN(n3951) );
  OAI221_X1 U4632 ( .B1(n3953), .B2(keyinput50), .C1(n3952), .C2(keyinput45), 
        .A(n3951), .ZN(n3964) );
  INV_X1 U4633 ( .A(REG2_REG_6__SCAN_IN), .ZN(n3956) );
  INV_X1 U4634 ( .A(ADDR_REG_8__SCAN_IN), .ZN(n3955) );
  AOI22_X1 U4635 ( .A1(n3956), .A2(keyinput37), .B1(keyinput26), .B2(n3955), 
        .ZN(n3954) );
  OAI221_X1 U4636 ( .B1(n3956), .B2(keyinput37), .C1(n3955), .C2(keyinput26), 
        .A(n3954), .ZN(n3963) );
  AOI22_X1 U4637 ( .A1(n4534), .A2(keyinput48), .B1(keyinput36), .B2(n3958), 
        .ZN(n3957) );
  OAI221_X1 U4638 ( .B1(n4534), .B2(keyinput48), .C1(n3958), .C2(keyinput36), 
        .A(n3957), .ZN(n3962) );
  INV_X1 U4639 ( .A(IR_REG_16__SCAN_IN), .ZN(n3960) );
  AOI22_X1 U4640 ( .A1(n4737), .A2(keyinput58), .B1(n3960), .B2(keyinput25), 
        .ZN(n3959) );
  OAI221_X1 U4641 ( .B1(n4737), .B2(keyinput58), .C1(n3960), .C2(keyinput25), 
        .A(n3959), .ZN(n3961) );
  NOR4_X1 U4642 ( .A1(n3964), .A2(n3963), .A3(n3962), .A4(n3961), .ZN(n4005)
         );
  INV_X1 U4643 ( .A(B_REG_SCAN_IN), .ZN(n4094) );
  AOI22_X1 U4644 ( .A1(n2321), .A2(keyinput28), .B1(n4094), .B2(keyinput33), 
        .ZN(n3965) );
  OAI221_X1 U4645 ( .B1(n2321), .B2(keyinput28), .C1(n4094), .C2(keyinput33), 
        .A(n3965), .ZN(n3976) );
  INV_X1 U4646 ( .A(REG2_REG_4__SCAN_IN), .ZN(n3968) );
  AOI22_X1 U4647 ( .A1(n3968), .A2(keyinput34), .B1(n3967), .B2(keyinput40), 
        .ZN(n3966) );
  OAI221_X1 U4648 ( .B1(n3968), .B2(keyinput34), .C1(n3967), .C2(keyinput40), 
        .A(n3966), .ZN(n3975) );
  INV_X1 U4649 ( .A(ADDR_REG_19__SCAN_IN), .ZN(n3970) );
  AOI22_X1 U4650 ( .A1(n3970), .A2(keyinput44), .B1(n4077), .B2(keyinput62), 
        .ZN(n3969) );
  OAI221_X1 U4651 ( .B1(n3970), .B2(keyinput44), .C1(n4077), .C2(keyinput62), 
        .A(n3969), .ZN(n3974) );
  XOR2_X1 U4652 ( .A(n4735), .B(keyinput54), .Z(n3972) );
  XNOR2_X1 U4653 ( .A(REG3_REG_11__SCAN_IN), .B(keyinput53), .ZN(n3971) );
  NAND2_X1 U4654 ( .A1(n3972), .A2(n3971), .ZN(n3973) );
  NOR4_X1 U4655 ( .A1(n3976), .A2(n3975), .A3(n3974), .A4(n3973), .ZN(n4004)
         );
  AOI22_X1 U4656 ( .A1(n3979), .A2(keyinput24), .B1(n3978), .B2(keyinput41), 
        .ZN(n3977) );
  OAI221_X1 U4657 ( .B1(n3979), .B2(keyinput24), .C1(n3978), .C2(keyinput41), 
        .A(n3977), .ZN(n3983) );
  XNOR2_X1 U4658 ( .A(n2186), .B(keyinput22), .ZN(n3982) );
  XNOR2_X1 U4659 ( .A(n3980), .B(keyinput30), .ZN(n3981) );
  OR3_X1 U4660 ( .A1(n3983), .A2(n3982), .A3(n3981), .ZN(n3989) );
  INV_X1 U4661 ( .A(D_REG_20__SCAN_IN), .ZN(n4685) );
  AOI22_X1 U4662 ( .A1(n4685), .A2(keyinput42), .B1(keyinput60), .B2(n4643), 
        .ZN(n3984) );
  OAI221_X1 U4663 ( .B1(n4685), .B2(keyinput42), .C1(n4643), .C2(keyinput60), 
        .A(n3984), .ZN(n3988) );
  INV_X1 U4664 ( .A(ADDR_REG_14__SCAN_IN), .ZN(n4049) );
  AOI22_X1 U4665 ( .A1(n3986), .A2(keyinput52), .B1(n4049), .B2(keyinput56), 
        .ZN(n3985) );
  OAI221_X1 U4666 ( .B1(n3986), .B2(keyinput52), .C1(n4049), .C2(keyinput56), 
        .A(n3985), .ZN(n3987) );
  NOR3_X1 U4667 ( .A1(n3989), .A2(n3988), .A3(n3987), .ZN(n4003) );
  INV_X1 U4668 ( .A(REG1_REG_22__SCAN_IN), .ZN(n3991) );
  INV_X1 U4669 ( .A(D_REG_15__SCAN_IN), .ZN(n4686) );
  AOI22_X1 U4670 ( .A1(n3991), .A2(keyinput32), .B1(n4686), .B2(keyinput49), 
        .ZN(n3990) );
  OAI221_X1 U4671 ( .B1(n3991), .B2(keyinput32), .C1(n4686), .C2(keyinput49), 
        .A(n3990), .ZN(n4001) );
  XNOR2_X1 U4672 ( .A(keyinput20), .B(n3992), .ZN(n4000) );
  INV_X1 U4673 ( .A(DATAI_11_), .ZN(n3993) );
  XNOR2_X1 U4674 ( .A(keyinput29), .B(n3993), .ZN(n3999) );
  XNOR2_X1 U4675 ( .A(IR_REG_7__SCAN_IN), .B(keyinput46), .ZN(n3997) );
  XNOR2_X1 U4676 ( .A(DATAI_8_), .B(keyinput57), .ZN(n3996) );
  XNOR2_X1 U4677 ( .A(IR_REG_22__SCAN_IN), .B(keyinput61), .ZN(n3995) );
  XNOR2_X1 U4678 ( .A(DATAI_1_), .B(keyinput38), .ZN(n3994) );
  NAND4_X1 U4679 ( .A1(n3997), .A2(n3996), .A3(n3995), .A4(n3994), .ZN(n3998)
         );
  NOR4_X1 U4680 ( .A1(n4001), .A2(n4000), .A3(n3999), .A4(n3998), .ZN(n4002)
         );
  NAND4_X1 U4681 ( .A1(n4005), .A2(n4004), .A3(n4003), .A4(n4002), .ZN(n4006)
         );
  NOR3_X1 U4682 ( .A1(n4008), .A2(n4007), .A3(n4006), .ZN(n4009) );
  XOR2_X1 U4683 ( .A(n4010), .B(n4009), .Z(U3569) );
  MUX2_X1 U4684 ( .A(n4333), .B(DATAO_REG_18__SCAN_IN), .S(n4017), .Z(U3568)
         );
  MUX2_X1 U4685 ( .A(n4347), .B(DATAO_REG_17__SCAN_IN), .S(n4017), .Z(U3567)
         );
  MUX2_X1 U4686 ( .A(DATAO_REG_16__SCAN_IN), .B(n2469), .S(U4043), .Z(U3566)
         );
  MUX2_X1 U4687 ( .A(n4389), .B(DATAO_REG_15__SCAN_IN), .S(n4017), .Z(U3565)
         );
  MUX2_X1 U4688 ( .A(DATAO_REG_14__SCAN_IN), .B(n4011), .S(U4043), .Z(U3564)
         );
  MUX2_X1 U4689 ( .A(n4387), .B(DATAO_REG_13__SCAN_IN), .S(n4017), .Z(U3563)
         );
  MUX2_X1 U4690 ( .A(n4012), .B(DATAO_REG_12__SCAN_IN), .S(n4017), .Z(U3562)
         );
  MUX2_X1 U4691 ( .A(DATAO_REG_11__SCAN_IN), .B(n4013), .S(U4043), .Z(U3561)
         );
  MUX2_X1 U4692 ( .A(DATAO_REG_10__SCAN_IN), .B(n4014), .S(U4043), .Z(U3560)
         );
  MUX2_X1 U4693 ( .A(n2409), .B(DATAO_REG_9__SCAN_IN), .S(n4017), .Z(U3559) );
  MUX2_X1 U4694 ( .A(n4015), .B(DATAO_REG_6__SCAN_IN), .S(n4017), .Z(U3556) );
  MUX2_X1 U4695 ( .A(DATAO_REG_5__SCAN_IN), .B(n2616), .S(U4043), .Z(U3555) );
  MUX2_X1 U4696 ( .A(n4016), .B(DATAO_REG_3__SCAN_IN), .S(n4017), .Z(U3553) );
  MUX2_X1 U4697 ( .A(DATAO_REG_2__SCAN_IN), .B(n2745), .S(U4043), .Z(U3552) );
  MUX2_X1 U4698 ( .A(n3024), .B(DATAO_REG_0__SCAN_IN), .S(n4017), .Z(U3550) );
  OAI211_X1 U4699 ( .C1(n4020), .C2(n4019), .A(n4670), .B(n4018), .ZN(n4028)
         );
  MUX2_X1 U4700 ( .A(REG1_REG_1__SCAN_IN), .B(n2931), .S(n2933), .Z(n4022) );
  OAI21_X1 U4701 ( .B1(n2300), .B2(n4023), .A(n4022), .ZN(n4024) );
  NAND3_X1 U4702 ( .A1(n4654), .A2(n4021), .A3(n4024), .ZN(n4027) );
  INV_X1 U4703 ( .A(n4673), .ZN(n4067) );
  NAND2_X1 U4704 ( .A1(n4067), .A2(n2932), .ZN(n4026) );
  AOI22_X1 U4705 ( .A1(n4660), .A2(ADDR_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(U3149), .ZN(n4025) );
  NAND4_X1 U4706 ( .A1(n4028), .A2(n4027), .A3(n4026), .A4(n4025), .ZN(U3241)
         );
  AOI22_X1 U4707 ( .A1(ADDR_REG_2__SCAN_IN), .A2(n4660), .B1(
        REG3_REG_2__SCAN_IN), .B2(U3149), .ZN(n4042) );
  INV_X1 U4708 ( .A(n4029), .ZN(n4030) );
  NAND3_X1 U4709 ( .A1(n4021), .A2(n4031), .A3(n4030), .ZN(n4032) );
  NAND3_X1 U4710 ( .A1(n4654), .A2(n4033), .A3(n4032), .ZN(n4039) );
  NAND3_X1 U4711 ( .A1(n4018), .A2(n4035), .A3(n4034), .ZN(n4036) );
  NAND3_X1 U4712 ( .A1(n4670), .A2(n4037), .A3(n4036), .ZN(n4038) );
  OAI211_X1 U4713 ( .C1(n4673), .C2(n2308), .A(n4039), .B(n4038), .ZN(n4040)
         );
  INV_X1 U4714 ( .A(n4040), .ZN(n4041) );
  NAND3_X1 U4715 ( .A1(n4043), .A2(n4042), .A3(n4041), .ZN(U3242) );
  INV_X1 U4716 ( .A(n4044), .ZN(n4615) );
  XNOR2_X1 U4717 ( .A(n4063), .B(n4614), .ZN(n4047) );
  NAND2_X1 U4718 ( .A1(n4047), .A2(REG2_REG_14__SCAN_IN), .ZN(n4065) );
  OAI211_X1 U4719 ( .C1(n4047), .C2(REG2_REG_14__SCAN_IN), .A(n4065), .B(n4670), .ZN(n4055) );
  INV_X1 U4720 ( .A(n4660), .ZN(n4644) );
  OAI21_X1 U4721 ( .B1(n4644), .B2(n4049), .A(n4048), .ZN(n4050) );
  AOI21_X1 U4722 ( .B1(n4614), .B2(n4067), .A(n4050), .ZN(n4054) );
  XNOR2_X1 U4723 ( .A(n4056), .B(n4614), .ZN(n4052) );
  NAND2_X1 U4724 ( .A1(n4052), .A2(REG1_REG_14__SCAN_IN), .ZN(n4059) );
  OAI211_X1 U4725 ( .C1(n4052), .C2(REG1_REG_14__SCAN_IN), .A(n4059), .B(n4654), .ZN(n4053) );
  NAND3_X1 U4726 ( .A1(n4055), .A2(n4054), .A3(n4053), .ZN(U3254) );
  INV_X1 U4727 ( .A(n4614), .ZN(n4062) );
  XOR2_X1 U4728 ( .A(REG1_REG_15__SCAN_IN), .B(n4613), .Z(n4635) );
  INV_X1 U4729 ( .A(n4613), .ZN(n4639) );
  INV_X1 U4730 ( .A(REG1_REG_15__SCAN_IN), .ZN(n4522) );
  NOR2_X1 U4731 ( .A1(n4639), .A2(n4522), .ZN(n4060) );
  XOR2_X1 U4732 ( .A(REG1_REG_16__SCAN_IN), .B(n4075), .Z(n4074) );
  OR2_X1 U4733 ( .A1(n4063), .A2(n4062), .ZN(n4064) );
  NAND2_X1 U4734 ( .A1(n4065), .A2(n4064), .ZN(n4633) );
  MUX2_X1 U4735 ( .A(REG2_REG_15__SCAN_IN), .B(n4066), .S(n4613), .Z(n4632) );
  XOR2_X1 U4736 ( .A(n4362), .B(n4080), .Z(n4072) );
  NAND2_X1 U4737 ( .A1(n4067), .A2(n4612), .ZN(n4069) );
  OAI211_X1 U4738 ( .C1(n4070), .C2(n4644), .A(n4069), .B(n4068), .ZN(n4071)
         );
  AOI21_X1 U4739 ( .B1(n4072), .B2(n4670), .A(n4071), .ZN(n4073) );
  OAI21_X1 U4740 ( .B1(n4074), .B2(n4657), .A(n4073), .ZN(U3256) );
  INV_X1 U4741 ( .A(n4082), .ZN(n4695) );
  AOI22_X1 U4742 ( .A1(n4082), .A2(REG1_REG_17__SCAN_IN), .B1(n4513), .B2(
        n4695), .ZN(n4648) );
  OR2_X1 U4743 ( .A1(n4082), .A2(REG1_REG_17__SCAN_IN), .ZN(n4076) );
  INV_X1 U4744 ( .A(n4083), .ZN(n4693) );
  AOI22_X1 U4745 ( .A1(REG1_REG_18__SCAN_IN), .A2(n4693), .B1(n4083), .B2(
        n4077), .ZN(n4658) );
  NAND2_X1 U4746 ( .A1(REG2_REG_18__SCAN_IN), .A2(n4083), .ZN(n4078) );
  OAI21_X1 U4747 ( .B1(REG2_REG_18__SCAN_IN), .B2(n4083), .A(n4078), .ZN(n4668) );
  NOR2_X1 U4748 ( .A1(n4082), .A2(REG2_REG_17__SCAN_IN), .ZN(n4081) );
  AOI21_X1 U4749 ( .B1(REG2_REG_17__SCAN_IN), .B2(n4082), .A(n4081), .ZN(n4651) );
  NOR2_X1 U4750 ( .A1(n4668), .A2(n4667), .ZN(n4666) );
  AOI21_X1 U4751 ( .B1(n4083), .B2(REG2_REG_18__SCAN_IN), .A(n4666), .ZN(n4085) );
  MUX2_X1 U4752 ( .A(REG2_REG_19__SCAN_IN), .B(n4304), .S(n4611), .Z(n4084) );
  XNOR2_X1 U4753 ( .A(n4085), .B(n4084), .ZN(n4090) );
  NAND2_X1 U4754 ( .A1(n4660), .A2(ADDR_REG_19__SCAN_IN), .ZN(n4086) );
  OAI211_X1 U4755 ( .C1(n4673), .C2(n4088), .A(n4087), .B(n4086), .ZN(n4089)
         );
  AOI21_X1 U4756 ( .B1(n4090), .B2(n4670), .A(n4089), .ZN(n4091) );
  OAI21_X1 U4757 ( .B1(n4092), .B2(n4657), .A(n4091), .ZN(U3259) );
  XNOR2_X1 U4758 ( .A(n4101), .B(n4098), .ZN(n4544) );
  OR2_X1 U4759 ( .A1(n4095), .A2(n4094), .ZN(n4096) );
  AND2_X1 U4760 ( .A1(n4388), .A2(n4096), .ZN(n4121) );
  NAND2_X1 U4761 ( .A1(n4121), .A2(n4097), .ZN(n4104) );
  OAI21_X1 U4762 ( .B1(n4098), .B2(n4391), .A(n4104), .ZN(n4541) );
  NAND2_X1 U4763 ( .A1(n4682), .A2(n4541), .ZN(n4100) );
  NAND2_X1 U4764 ( .A1(n4431), .A2(REG2_REG_31__SCAN_IN), .ZN(n4099) );
  OAI211_X1 U4765 ( .C1(n4544), .C2(n4450), .A(n4100), .B(n4099), .ZN(U3260)
         );
  INV_X1 U4766 ( .A(REG2_REG_30__SCAN_IN), .ZN(n4107) );
  AOI21_X1 U4767 ( .B1(n4102), .B2(n2019), .A(n4101), .ZN(n4545) );
  NAND2_X1 U4768 ( .A1(n4545), .A2(n4358), .ZN(n4106) );
  NAND2_X1 U4769 ( .A1(n4102), .A2(n4439), .ZN(n4103) );
  NAND2_X1 U4770 ( .A1(n4104), .A2(n4103), .ZN(n4546) );
  NAND2_X1 U4771 ( .A1(n4682), .A2(n4546), .ZN(n4105) );
  OAI211_X1 U4772 ( .C1(n4682), .C2(n4107), .A(n4106), .B(n4105), .ZN(U3261)
         );
  NAND2_X1 U4773 ( .A1(n4111), .A2(n4110), .ZN(n4463) );
  NAND2_X1 U4774 ( .A1(n4461), .A2(n4463), .ZN(n4112) );
  XNOR2_X1 U4775 ( .A(n4112), .B(n4462), .ZN(n4129) );
  NAND2_X1 U4776 ( .A1(n2033), .A2(n4119), .ZN(n4113) );
  AOI22_X1 U4777 ( .A1(n4465), .A2(n4358), .B1(REG2_REG_29__SCAN_IN), .B2(
        n4431), .ZN(n4128) );
  INV_X1 U4778 ( .A(n4114), .ZN(n4116) );
  AOI22_X1 U4779 ( .A1(n4121), .A2(n4120), .B1(n4439), .B2(n4119), .ZN(n4122)
         );
  OAI21_X1 U4780 ( .B1(n4145), .B2(n4434), .A(n4122), .ZN(n4123) );
  OAI21_X1 U4781 ( .B1(n4125), .B2(n4360), .A(n4469), .ZN(n4126) );
  NAND2_X1 U4782 ( .A1(n4126), .A2(n4682), .ZN(n4127) );
  OAI211_X1 U4783 ( .C1(n4129), .C2(n4344), .A(n4128), .B(n4127), .ZN(U3354)
         );
  INV_X1 U4784 ( .A(n4130), .ZN(n4138) );
  OAI22_X1 U4785 ( .A1(n4132), .A2(n4360), .B1(n4131), .B2(n4682), .ZN(n4135)
         );
  NOR2_X1 U4786 ( .A1(n4133), .A2(n4450), .ZN(n4134) );
  AOI211_X1 U4787 ( .C1(n4136), .C2(n4682), .A(n4135), .B(n4134), .ZN(n4137)
         );
  OAI21_X1 U4788 ( .B1(n4138), .B2(n4344), .A(n4137), .ZN(U3262) );
  XOR2_X1 U4789 ( .A(n4140), .B(n4139), .Z(n4471) );
  INV_X1 U4790 ( .A(n4471), .ZN(n4155) );
  XNOR2_X1 U4791 ( .A(n4141), .B(n4140), .ZN(n4147) );
  OAI22_X1 U4792 ( .A1(n4142), .A2(n4434), .B1(n4148), .B2(n4391), .ZN(n4143)
         );
  INV_X1 U4793 ( .A(n4143), .ZN(n4144) );
  OAI21_X1 U4794 ( .B1(n4145), .B2(n4436), .A(n4144), .ZN(n4146) );
  AOI21_X1 U4795 ( .B1(n4147), .B2(n4393), .A(n4146), .ZN(n4472) );
  INV_X1 U4796 ( .A(n4472), .ZN(n4153) );
  NOR2_X1 U4797 ( .A1(n4170), .A2(n4148), .ZN(n4149) );
  OR2_X1 U4798 ( .A1(n2703), .A2(n4149), .ZN(n4474) );
  AOI22_X1 U4799 ( .A1(n4150), .A2(n4678), .B1(REG2_REG_27__SCAN_IN), .B2(
        n4431), .ZN(n4151) );
  OAI21_X1 U4800 ( .B1(n4474), .B2(n4450), .A(n4151), .ZN(n4152) );
  AOI21_X1 U4801 ( .B1(n4153), .B2(n4682), .A(n4152), .ZN(n4154) );
  OAI21_X1 U4802 ( .B1(n4155), .B2(n4344), .A(n4154), .ZN(U3263) );
  NAND2_X1 U4803 ( .A1(n4157), .A2(n4156), .ZN(n4158) );
  XOR2_X1 U4804 ( .A(n4161), .B(n4158), .Z(n4476) );
  INV_X1 U4805 ( .A(n4476), .ZN(n4177) );
  NAND2_X1 U4806 ( .A1(n4160), .A2(n4159), .ZN(n4162) );
  XNOR2_X1 U4807 ( .A(n4162), .B(n4161), .ZN(n4167) );
  OAI22_X1 U4808 ( .A1(n4163), .A2(n4434), .B1(n4172), .B2(n4391), .ZN(n4164)
         );
  AOI21_X1 U4809 ( .B1(n4388), .B2(n4165), .A(n4164), .ZN(n4166) );
  OAI22_X1 U4810 ( .A1(n4169), .A2(n4360), .B1(n4168), .B2(n4682), .ZN(n4175)
         );
  INV_X1 U4811 ( .A(n4197), .ZN(n4173) );
  INV_X1 U4812 ( .A(n4170), .ZN(n4171) );
  OAI21_X1 U4813 ( .B1(n4173), .B2(n4172), .A(n4171), .ZN(n4555) );
  NOR2_X1 U4814 ( .A1(n4555), .A2(n4450), .ZN(n4174) );
  AOI211_X1 U4815 ( .C1(n4475), .C2(n4682), .A(n4175), .B(n4174), .ZN(n4176)
         );
  OAI21_X1 U4816 ( .B1(n4177), .B2(n4344), .A(n4176), .ZN(U3264) );
  NAND2_X1 U4817 ( .A1(n4179), .A2(n4178), .ZN(n4181) );
  NAND2_X1 U4818 ( .A1(n4206), .A2(n4182), .ZN(n4184) );
  NAND2_X1 U4819 ( .A1(n4184), .A2(n4183), .ZN(n4185) );
  XNOR2_X1 U4820 ( .A(n4185), .B(n4188), .ZN(n4480) );
  INV_X1 U4821 ( .A(n4480), .ZN(n4204) );
  NAND2_X1 U4822 ( .A1(n4186), .A2(n4187), .ZN(n4189) );
  XNOR2_X1 U4823 ( .A(n4189), .B(n4188), .ZN(n4190) );
  NAND2_X1 U4824 ( .A1(n4190), .A2(n4393), .ZN(n4195) );
  OAI22_X1 U4825 ( .A1(n4191), .A2(n4434), .B1(n4198), .B2(n4391), .ZN(n4192)
         );
  AOI21_X1 U4826 ( .B1(n4193), .B2(n4388), .A(n4192), .ZN(n4194) );
  NAND2_X1 U4827 ( .A1(n4195), .A2(n4194), .ZN(n4479) );
  INV_X1 U4828 ( .A(n4196), .ZN(n4199) );
  OAI21_X1 U4829 ( .B1(n4199), .B2(n4198), .A(n4197), .ZN(n4559) );
  AOI22_X1 U4830 ( .A1(n4200), .A2(n4678), .B1(REG2_REG_25__SCAN_IN), .B2(
        n4431), .ZN(n4201) );
  OAI21_X1 U4831 ( .B1(n4559), .B2(n4450), .A(n4201), .ZN(n4202) );
  AOI21_X1 U4832 ( .B1(n4682), .B2(n4479), .A(n4202), .ZN(n4203) );
  OAI21_X1 U4833 ( .B1(n4204), .B2(n4344), .A(n4203), .ZN(U3265) );
  NAND2_X1 U4834 ( .A1(n4206), .A2(n4205), .ZN(n4207) );
  XOR2_X1 U4835 ( .A(n4211), .B(n4207), .Z(n4484) );
  OR2_X1 U4836 ( .A1(n4208), .A2(n4214), .ZN(n4209) );
  NAND2_X1 U4837 ( .A1(n4196), .A2(n4209), .ZN(n4563) );
  INV_X1 U4838 ( .A(n4211), .ZN(n4212) );
  XNOR2_X1 U4839 ( .A(n4210), .B(n4212), .ZN(n4213) );
  NAND2_X1 U4840 ( .A1(n4213), .A2(n4393), .ZN(n4219) );
  OAI22_X1 U4841 ( .A1(n4215), .A2(n4434), .B1(n4214), .B2(n4391), .ZN(n4216)
         );
  AOI21_X1 U4842 ( .B1(n4217), .B2(n4388), .A(n4216), .ZN(n4218) );
  NAND2_X1 U4843 ( .A1(n4219), .A2(n4218), .ZN(n4483) );
  NAND2_X1 U4844 ( .A1(n4483), .A2(n4682), .ZN(n4222) );
  AOI22_X1 U4845 ( .A1(n4220), .A2(n4678), .B1(REG2_REG_24__SCAN_IN), .B2(
        n4431), .ZN(n4221) );
  OAI211_X1 U4846 ( .C1(n4563), .C2(n4450), .A(n4222), .B(n4221), .ZN(n4223)
         );
  AOI21_X1 U4847 ( .B1(n4484), .B2(n4452), .A(n4223), .ZN(n4224) );
  INV_X1 U4848 ( .A(n4224), .ZN(U3266) );
  NAND2_X1 U4849 ( .A1(n4226), .A2(n4225), .ZN(n4228) );
  NAND2_X1 U4850 ( .A1(n4228), .A2(n4227), .ZN(n4229) );
  XOR2_X1 U4851 ( .A(n4235), .B(n4229), .Z(n4488) );
  INV_X1 U4852 ( .A(n4488), .ZN(n4248) );
  INV_X1 U4853 ( .A(n4230), .ZN(n4231) );
  AOI21_X1 U4854 ( .B1(n4233), .B2(n4232), .A(n4231), .ZN(n4234) );
  XOR2_X1 U4855 ( .A(n4235), .B(n4234), .Z(n4240) );
  OAI22_X1 U4856 ( .A1(n4236), .A2(n4434), .B1(n4391), .B2(n4241), .ZN(n4237)
         );
  AOI21_X1 U4857 ( .B1(n4238), .B2(n4388), .A(n4237), .ZN(n4239) );
  OAI21_X1 U4858 ( .B1(n4240), .B2(n4442), .A(n4239), .ZN(n4487) );
  NOR2_X1 U4859 ( .A1(n3490), .A2(n4241), .ZN(n4242) );
  NOR2_X1 U4860 ( .A1(n4567), .A2(n4450), .ZN(n4246) );
  OAI22_X1 U4861 ( .A1(n4244), .A2(n4360), .B1(n4243), .B2(n4682), .ZN(n4245)
         );
  AOI211_X1 U4862 ( .C1(n4487), .C2(n4682), .A(n4246), .B(n4245), .ZN(n4247)
         );
  OAI21_X1 U4863 ( .B1(n4248), .B2(n4344), .A(n4247), .ZN(U3267) );
  XNOR2_X1 U4864 ( .A(n4249), .B(n4250), .ZN(n4497) );
  INV_X1 U4865 ( .A(n4497), .ZN(n4264) );
  XOR2_X1 U4866 ( .A(n4250), .B(n3486), .Z(n4256) );
  OAI22_X1 U4867 ( .A1(n4252), .A2(n4434), .B1(n4391), .B2(n4251), .ZN(n4253)
         );
  AOI21_X1 U4868 ( .B1(n4254), .B2(n4388), .A(n4253), .ZN(n4255) );
  OAI21_X1 U4869 ( .B1(n4256), .B2(n4442), .A(n4255), .ZN(n4496) );
  NAND2_X1 U4870 ( .A1(n4279), .A2(n4257), .ZN(n4258) );
  NAND2_X1 U4871 ( .A1(n2041), .A2(n4258), .ZN(n4572) );
  NOR2_X1 U4872 ( .A1(n4572), .A2(n4450), .ZN(n4262) );
  OAI22_X1 U4873 ( .A1(n4260), .A2(n4360), .B1(n4259), .B2(n4682), .ZN(n4261)
         );
  AOI211_X1 U4874 ( .C1(n4496), .C2(n4682), .A(n4262), .B(n4261), .ZN(n4263)
         );
  OAI21_X1 U4875 ( .B1(n4264), .B2(n4344), .A(n4263), .ZN(U3269) );
  XNOR2_X1 U4876 ( .A(n4265), .B(n4268), .ZN(n4277) );
  NAND2_X1 U4877 ( .A1(n4267), .A2(n4266), .ZN(n4269) );
  XNOR2_X1 U4878 ( .A(n4269), .B(n4268), .ZN(n4275) );
  AOI22_X1 U4879 ( .A1(n4271), .A2(n4386), .B1(n4270), .B2(n4439), .ZN(n4272)
         );
  OAI21_X1 U4880 ( .B1(n4273), .B2(n4436), .A(n4272), .ZN(n4274) );
  AOI21_X1 U4881 ( .B1(n4275), .B2(n4393), .A(n4274), .ZN(n4276) );
  OAI21_X1 U4882 ( .B1(n4277), .B2(n4417), .A(n4276), .ZN(n4500) );
  INV_X1 U4883 ( .A(n4500), .ZN(n4285) );
  INV_X1 U4884 ( .A(n4277), .ZN(n4501) );
  OAI21_X1 U4885 ( .B1(n4278), .B2(n4280), .A(n4279), .ZN(n4576) );
  AOI22_X1 U4886 ( .A1(n4281), .A2(n4678), .B1(REG2_REG_20__SCAN_IN), .B2(
        n4431), .ZN(n4282) );
  OAI21_X1 U4887 ( .B1(n4576), .B2(n4450), .A(n4282), .ZN(n4283) );
  AOI21_X1 U4888 ( .B1(n4501), .B2(n4680), .A(n4283), .ZN(n4284) );
  OAI21_X1 U4889 ( .B1(n4285), .B2(n4431), .A(n4284), .ZN(U3270) );
  XNOR2_X1 U4890 ( .A(n4286), .B(n4292), .ZN(n4505) );
  INV_X1 U4891 ( .A(n4505), .ZN(n4308) );
  OAI21_X1 U4892 ( .B1(n4330), .B2(n4288), .A(n4287), .ZN(n4309) );
  INV_X1 U4893 ( .A(n4289), .ZN(n4291) );
  OAI21_X1 U4894 ( .B1(n4309), .B2(n4291), .A(n4290), .ZN(n4294) );
  INV_X1 U4895 ( .A(n4292), .ZN(n4293) );
  XNOR2_X1 U4896 ( .A(n4294), .B(n4293), .ZN(n4299) );
  OAI22_X1 U4897 ( .A1(n4295), .A2(n4434), .B1(n4391), .B2(n4301), .ZN(n4296)
         );
  AOI21_X1 U4898 ( .B1(n4297), .B2(n4388), .A(n4296), .ZN(n4298) );
  OAI21_X1 U4899 ( .B1(n4299), .B2(n4442), .A(n4298), .ZN(n4504) );
  INV_X1 U4900 ( .A(n4316), .ZN(n4302) );
  INV_X1 U4901 ( .A(n4278), .ZN(n4300) );
  OAI21_X1 U4902 ( .B1(n4302), .B2(n4301), .A(n4300), .ZN(n4580) );
  NOR2_X1 U4903 ( .A1(n4580), .A2(n4450), .ZN(n4306) );
  OAI22_X1 U4904 ( .A1(n4682), .A2(n4304), .B1(n4303), .B2(n4360), .ZN(n4305)
         );
  AOI211_X1 U4905 ( .C1(n4504), .C2(n4682), .A(n4306), .B(n4305), .ZN(n4307)
         );
  OAI21_X1 U4906 ( .B1(n4308), .B2(n4344), .A(n4307), .ZN(U3271) );
  XNOR2_X1 U4907 ( .A(n4309), .B(n4323), .ZN(n4313) );
  AOI22_X1 U4908 ( .A1(n4347), .A2(n4386), .B1(n4315), .B2(n4439), .ZN(n4310)
         );
  OAI21_X1 U4909 ( .B1(n4311), .B2(n4436), .A(n4310), .ZN(n4312) );
  AOI21_X1 U4910 ( .B1(n4313), .B2(n4393), .A(n4312), .ZN(n4509) );
  AOI21_X1 U4911 ( .B1(n4338), .B2(n4315), .A(n2725), .ZN(n4317) );
  NAND2_X1 U4912 ( .A1(n4317), .A2(n4316), .ZN(n4508) );
  INV_X1 U4913 ( .A(n4508), .ZN(n4327) );
  INV_X1 U4914 ( .A(REG2_REG_18__SCAN_IN), .ZN(n4319) );
  OAI22_X1 U4915 ( .A1(n4682), .A2(n4319), .B1(n4318), .B2(n4360), .ZN(n4325)
         );
  INV_X1 U4916 ( .A(n4321), .ZN(n4322) );
  AOI21_X1 U4917 ( .B1(n4323), .B2(n4320), .A(n4322), .ZN(n4510) );
  NOR2_X1 U4918 ( .A1(n4510), .A2(n4344), .ZN(n4324) );
  AOI211_X1 U4919 ( .C1(n4327), .C2(n4326), .A(n4325), .B(n4324), .ZN(n4328)
         );
  OAI21_X1 U4920 ( .B1(n4684), .B2(n4509), .A(n4328), .ZN(U3272) );
  XOR2_X1 U4921 ( .A(n4331), .B(n4329), .Z(n4512) );
  INV_X1 U4922 ( .A(n4512), .ZN(n4345) );
  XOR2_X1 U4923 ( .A(n4331), .B(n4330), .Z(n4335) );
  OAI22_X1 U4924 ( .A1(n4367), .A2(n4434), .B1(n4391), .B2(n2483), .ZN(n4332)
         );
  AOI21_X1 U4925 ( .B1(n4333), .B2(n4388), .A(n4332), .ZN(n4334) );
  OAI21_X1 U4926 ( .B1(n4335), .B2(n4442), .A(n4334), .ZN(n4511) );
  NAND2_X1 U4927 ( .A1(n2049), .A2(n4336), .ZN(n4337) );
  NAND2_X1 U4928 ( .A1(n4338), .A2(n4337), .ZN(n4585) );
  NOR2_X1 U4929 ( .A1(n4585), .A2(n4450), .ZN(n4342) );
  OAI22_X1 U4930 ( .A1(n4682), .A2(n4340), .B1(n4339), .B2(n4360), .ZN(n4341)
         );
  AOI211_X1 U4931 ( .C1(n4511), .C2(n4682), .A(n4342), .B(n4341), .ZN(n4343)
         );
  OAI21_X1 U4932 ( .B1(n4345), .B2(n4344), .A(n4343), .ZN(U3273) );
  XNOR2_X1 U4933 ( .A(n4346), .B(n4353), .ZN(n4351) );
  AOI22_X1 U4934 ( .A1(n4347), .A2(n4388), .B1(n4386), .B2(n4389), .ZN(n4348)
         );
  OAI21_X1 U4935 ( .B1(n4349), .B2(n4391), .A(n4348), .ZN(n4350) );
  AOI21_X1 U4936 ( .B1(n4351), .B2(n4393), .A(n4350), .ZN(n4517) );
  OAI21_X1 U4937 ( .B1(n4354), .B2(n4353), .A(n4352), .ZN(n4518) );
  INV_X1 U4938 ( .A(n4518), .ZN(n4365) );
  INV_X1 U4939 ( .A(n4355), .ZN(n4357) );
  NAND2_X1 U4940 ( .A1(n4357), .A2(n4356), .ZN(n4515) );
  AND3_X1 U4941 ( .A1(n4515), .A2(n4358), .A3(n2049), .ZN(n4364) );
  INV_X1 U4942 ( .A(n4359), .ZN(n4361) );
  OAI22_X1 U4943 ( .A1(n4682), .A2(n4362), .B1(n4361), .B2(n4360), .ZN(n4363)
         );
  AOI211_X1 U4944 ( .C1(n4365), .C2(n4452), .A(n4364), .B(n4363), .ZN(n4366)
         );
  OAI21_X1 U4945 ( .B1(n4684), .B2(n4517), .A(n4366), .ZN(U3274) );
  OAI22_X1 U4946 ( .A1(n4367), .A2(n4436), .B1(n4414), .B2(n4434), .ZN(n4372)
         );
  NAND2_X1 U4947 ( .A1(n4385), .A2(n4368), .ZN(n4369) );
  XNOR2_X1 U4948 ( .A(n4369), .B(n4374), .ZN(n4370) );
  NOR2_X1 U4949 ( .A1(n4370), .A2(n4442), .ZN(n4371) );
  AOI211_X1 U4950 ( .C1(n4439), .C2(n4373), .A(n4372), .B(n4371), .ZN(n4519)
         );
  XNOR2_X1 U4951 ( .A(n4375), .B(n4374), .ZN(n4521) );
  NOR2_X1 U4952 ( .A1(n4397), .A2(n4376), .ZN(n4377) );
  AOI22_X1 U4953 ( .A1(n4431), .A2(REG2_REG_15__SCAN_IN), .B1(n4378), .B2(
        n4678), .ZN(n4379) );
  OAI21_X1 U4954 ( .B1(n4590), .B2(n4450), .A(n4379), .ZN(n4380) );
  AOI21_X1 U4955 ( .B1(n4521), .B2(n4452), .A(n4380), .ZN(n4381) );
  OAI21_X1 U4956 ( .B1(n4684), .B2(n4519), .A(n4381), .ZN(U3275) );
  OAI21_X1 U4957 ( .B1(n4384), .B2(n4383), .A(n4382), .ZN(n4525) );
  INV_X1 U4958 ( .A(n4525), .ZN(n4396) );
  OAI21_X1 U4959 ( .B1(n2190), .B2(n3709), .A(n4385), .ZN(n4394) );
  AOI22_X1 U4960 ( .A1(n4389), .A2(n4388), .B1(n4387), .B2(n4386), .ZN(n4390)
         );
  OAI21_X1 U4961 ( .B1(n4399), .B2(n4391), .A(n4390), .ZN(n4392) );
  AOI21_X1 U4962 ( .B1(n4394), .B2(n4393), .A(n4392), .ZN(n4395) );
  OAI21_X1 U4963 ( .B1(n4396), .B2(n4417), .A(n4395), .ZN(n4524) );
  INV_X1 U4964 ( .A(n4524), .ZN(n4405) );
  INV_X1 U4965 ( .A(n4426), .ZN(n4400) );
  INV_X1 U4966 ( .A(n4397), .ZN(n4398) );
  OAI21_X1 U4967 ( .B1(n4400), .B2(n4399), .A(n4398), .ZN(n4594) );
  AOI22_X1 U4968 ( .A1(n4431), .A2(REG2_REG_14__SCAN_IN), .B1(n4401), .B2(
        n4678), .ZN(n4402) );
  OAI21_X1 U4969 ( .B1(n4594), .B2(n4450), .A(n4402), .ZN(n4403) );
  AOI21_X1 U4970 ( .B1(n4525), .B2(n4680), .A(n4403), .ZN(n4404) );
  OAI21_X1 U4971 ( .B1(n4405), .B2(n4431), .A(n4404), .ZN(U3276) );
  INV_X1 U4972 ( .A(n4406), .ZN(n4407) );
  AOI21_X1 U4973 ( .B1(n3411), .B2(n4408), .A(n4407), .ZN(n4433) );
  INV_X1 U4974 ( .A(n4409), .ZN(n4410) );
  AOI21_X1 U4975 ( .B1(n4433), .B2(n4411), .A(n4410), .ZN(n4412) );
  XOR2_X1 U4976 ( .A(n4416), .B(n4412), .Z(n4421) );
  OAI22_X1 U4977 ( .A1(n4414), .A2(n4436), .B1(n4413), .B2(n4434), .ZN(n4419)
         );
  XOR2_X1 U4978 ( .A(n4416), .B(n4415), .Z(n4422) );
  NOR2_X1 U4979 ( .A1(n4422), .A2(n4417), .ZN(n4418) );
  AOI211_X1 U4980 ( .C1(n4439), .C2(n4424), .A(n4419), .B(n4418), .ZN(n4420)
         );
  OAI21_X1 U4981 ( .B1(n4442), .B2(n4421), .A(n4420), .ZN(n4528) );
  INV_X1 U4982 ( .A(n4528), .ZN(n4432) );
  INV_X1 U4983 ( .A(n4422), .ZN(n4529) );
  NAND2_X1 U4984 ( .A1(n4423), .A2(n4424), .ZN(n4425) );
  NAND2_X1 U4985 ( .A1(n4426), .A2(n4425), .ZN(n4598) );
  AOI22_X1 U4986 ( .A1(n4431), .A2(REG2_REG_13__SCAN_IN), .B1(n4427), .B2(
        n4678), .ZN(n4428) );
  OAI21_X1 U4987 ( .B1(n4598), .B2(n4450), .A(n4428), .ZN(n4429) );
  AOI21_X1 U4988 ( .B1(n4529), .B2(n4680), .A(n4429), .ZN(n4430) );
  OAI21_X1 U4989 ( .B1(n4432), .B2(n4431), .A(n4430), .ZN(U3277) );
  XOR2_X1 U4990 ( .A(n4444), .B(n4433), .Z(n4443) );
  OAI22_X1 U4991 ( .A1(n4437), .A2(n4436), .B1(n4435), .B2(n4434), .ZN(n4438)
         );
  AOI21_X1 U4992 ( .B1(n4440), .B2(n4439), .A(n4438), .ZN(n4441) );
  OAI21_X1 U4993 ( .B1(n4443), .B2(n4442), .A(n4441), .ZN(n4532) );
  INV_X1 U4994 ( .A(n4532), .ZN(n4454) );
  XNOR2_X1 U4995 ( .A(n4445), .B(n4444), .ZN(n4533) );
  OR2_X1 U4996 ( .A1(n3419), .A2(n4446), .ZN(n4447) );
  NAND2_X1 U4997 ( .A1(n4423), .A2(n4447), .ZN(n4602) );
  AOI22_X1 U4998 ( .A1(n4431), .A2(REG2_REG_12__SCAN_IN), .B1(n4448), .B2(
        n4678), .ZN(n4449) );
  OAI21_X1 U4999 ( .B1(n4602), .B2(n4450), .A(n4449), .ZN(n4451) );
  AOI21_X1 U5000 ( .B1(n4533), .B2(n4452), .A(n4451), .ZN(n4453) );
  OAI21_X1 U5001 ( .B1(n4454), .B2(n4431), .A(n4453), .ZN(U3278) );
  NAND2_X1 U5002 ( .A1(n4741), .A2(n4541), .ZN(n4456) );
  NAND2_X1 U5003 ( .A1(n2712), .A2(REG1_REG_31__SCAN_IN), .ZN(n4455) );
  OAI211_X1 U5004 ( .C1(n4544), .C2(n4540), .A(n4456), .B(n4455), .ZN(U3549)
         );
  INV_X1 U5005 ( .A(REG1_REG_30__SCAN_IN), .ZN(n4459) );
  NAND2_X1 U5006 ( .A1(n4545), .A2(n2707), .ZN(n4458) );
  NAND2_X1 U5007 ( .A1(n4741), .A2(n4546), .ZN(n4457) );
  OAI211_X1 U5008 ( .C1(n4741), .C2(n4459), .A(n4458), .B(n4457), .ZN(U3548)
         );
  NAND4_X1 U5009 ( .A1(n4461), .A2(n4724), .A3(n4462), .A4(n4463), .ZN(n4467)
         );
  NOR3_X1 U5010 ( .A1(n4463), .A2(n4462), .A3(n4715), .ZN(n4464) );
  NAND2_X1 U5011 ( .A1(n4470), .A2(n4469), .ZN(n4550) );
  MUX2_X1 U5012 ( .A(REG1_REG_29__SCAN_IN), .B(n4550), .S(n4741), .Z(U3547) );
  NAND2_X1 U5013 ( .A1(n4471), .A2(n4724), .ZN(n4473) );
  OAI211_X1 U5014 ( .C1(n2725), .C2(n4474), .A(n4473), .B(n4472), .ZN(n4551)
         );
  MUX2_X1 U5015 ( .A(REG1_REG_27__SCAN_IN), .B(n4551), .S(n4741), .Z(U3545) );
  INV_X1 U5016 ( .A(REG1_REG_26__SCAN_IN), .ZN(n4477) );
  AOI21_X1 U5017 ( .B1(n4476), .B2(n4724), .A(n4475), .ZN(n4552) );
  MUX2_X1 U5018 ( .A(n4477), .B(n4552), .S(n4741), .Z(n4478) );
  OAI21_X1 U5019 ( .B1(n4540), .B2(n4555), .A(n4478), .ZN(U3544) );
  INV_X1 U5020 ( .A(REG1_REG_25__SCAN_IN), .ZN(n4481) );
  AOI21_X1 U5021 ( .B1(n4480), .B2(n4724), .A(n4479), .ZN(n4556) );
  OAI21_X1 U5022 ( .B1(n4540), .B2(n4559), .A(n4482), .ZN(U3543) );
  AOI21_X1 U5023 ( .B1(n4484), .B2(n4724), .A(n4483), .ZN(n4560) );
  MUX2_X1 U5024 ( .A(n4485), .B(n4560), .S(n4741), .Z(n4486) );
  OAI21_X1 U5025 ( .B1(n4540), .B2(n4563), .A(n4486), .ZN(U3542) );
  INV_X1 U5026 ( .A(REG1_REG_23__SCAN_IN), .ZN(n4489) );
  AOI21_X1 U5027 ( .B1(n4488), .B2(n4724), .A(n4487), .ZN(n4564) );
  MUX2_X1 U5028 ( .A(n4489), .B(n4564), .S(n4741), .Z(n4490) );
  OAI21_X1 U5029 ( .B1(n4540), .B2(n4567), .A(n4490), .ZN(U3541) );
  NAND3_X1 U5030 ( .A1(n4492), .A2(n4721), .A3(n4491), .ZN(n4493) );
  OAI211_X1 U5031 ( .C1(n4495), .C2(n4715), .A(n4494), .B(n4493), .ZN(n4568)
         );
  MUX2_X1 U5032 ( .A(REG1_REG_22__SCAN_IN), .B(n4568), .S(n4741), .Z(U3540) );
  INV_X1 U5033 ( .A(REG1_REG_21__SCAN_IN), .ZN(n4498) );
  AOI21_X1 U5034 ( .B1(n4497), .B2(n4724), .A(n4496), .ZN(n4569) );
  MUX2_X1 U5035 ( .A(n4498), .B(n4569), .S(n4741), .Z(n4499) );
  OAI21_X1 U5036 ( .B1(n4540), .B2(n4572), .A(n4499), .ZN(U3539) );
  AOI21_X1 U5037 ( .B1(n4712), .B2(n4501), .A(n4500), .ZN(n4573) );
  MUX2_X1 U5038 ( .A(n4502), .B(n4573), .S(n4741), .Z(n4503) );
  OAI21_X1 U5039 ( .B1(n4540), .B2(n4576), .A(n4503), .ZN(U3538) );
  INV_X1 U5040 ( .A(REG1_REG_19__SCAN_IN), .ZN(n4506) );
  AOI21_X1 U5041 ( .B1(n4505), .B2(n4724), .A(n4504), .ZN(n4577) );
  MUX2_X1 U5042 ( .A(n4506), .B(n4577), .S(n4741), .Z(n4507) );
  OAI21_X1 U5043 ( .B1(n4540), .B2(n4580), .A(n4507), .ZN(U3537) );
  OAI211_X1 U5044 ( .C1(n4510), .C2(n4715), .A(n4509), .B(n4508), .ZN(n4581)
         );
  MUX2_X1 U5045 ( .A(REG1_REG_18__SCAN_IN), .B(n4581), .S(n4741), .Z(U3536) );
  AOI21_X1 U5046 ( .B1(n4512), .B2(n4724), .A(n4511), .ZN(n4582) );
  MUX2_X1 U5047 ( .A(n4513), .B(n4582), .S(n4741), .Z(n4514) );
  OAI21_X1 U5048 ( .B1(n4540), .B2(n4585), .A(n4514), .ZN(U3535) );
  NAND3_X1 U5049 ( .A1(n4515), .A2(n4721), .A3(n2049), .ZN(n4516) );
  OAI211_X1 U5050 ( .C1(n4518), .C2(n4715), .A(n4517), .B(n4516), .ZN(n4586)
         );
  MUX2_X1 U5051 ( .A(REG1_REG_16__SCAN_IN), .B(n4586), .S(n4741), .Z(U3534) );
  INV_X1 U5052 ( .A(n4519), .ZN(n4520) );
  AOI21_X1 U5053 ( .B1(n4521), .B2(n4724), .A(n4520), .ZN(n4587) );
  MUX2_X1 U5054 ( .A(n4522), .B(n4587), .S(n4741), .Z(n4523) );
  OAI21_X1 U5055 ( .B1(n4540), .B2(n4590), .A(n4523), .ZN(U3533) );
  INV_X1 U5056 ( .A(REG1_REG_14__SCAN_IN), .ZN(n4526) );
  AOI21_X1 U5057 ( .B1(n4712), .B2(n4525), .A(n4524), .ZN(n4591) );
  MUX2_X1 U5058 ( .A(n4526), .B(n4591), .S(n4741), .Z(n4527) );
  OAI21_X1 U5059 ( .B1(n4540), .B2(n4594), .A(n4527), .ZN(U3532) );
  INV_X1 U5060 ( .A(REG1_REG_13__SCAN_IN), .ZN(n4530) );
  AOI21_X1 U5061 ( .B1(n4712), .B2(n4529), .A(n4528), .ZN(n4595) );
  MUX2_X1 U5062 ( .A(n4530), .B(n4595), .S(n4741), .Z(n4531) );
  OAI21_X1 U5063 ( .B1(n4540), .B2(n4598), .A(n4531), .ZN(U3531) );
  AOI21_X1 U5064 ( .B1(n4724), .B2(n4533), .A(n4532), .ZN(n4599) );
  MUX2_X1 U5065 ( .A(n4534), .B(n4599), .S(n4741), .Z(n4535) );
  OAI21_X1 U5066 ( .B1(n4540), .B2(n4602), .A(n4535), .ZN(U3530) );
  INV_X1 U5067 ( .A(REG1_REG_11__SCAN_IN), .ZN(n4538) );
  AOI21_X1 U5068 ( .B1(n4712), .B2(n4537), .A(n4536), .ZN(n4603) );
  MUX2_X1 U5069 ( .A(n4538), .B(n4603), .S(n4741), .Z(n4539) );
  OAI21_X1 U5070 ( .B1(n4540), .B2(n4607), .A(n4539), .ZN(U3529) );
  NAND2_X1 U5071 ( .A1(n4731), .A2(n4541), .ZN(n4543) );
  NAND2_X1 U5072 ( .A1(n4729), .A2(REG0_REG_31__SCAN_IN), .ZN(n4542) );
  OAI211_X1 U5073 ( .C1(n4544), .C2(n4606), .A(n4543), .B(n4542), .ZN(U3517)
         );
  NAND2_X1 U5074 ( .A1(n4545), .A2(n2716), .ZN(n4548) );
  NAND2_X1 U5075 ( .A1(n4731), .A2(n4546), .ZN(n4547) );
  OAI211_X1 U5076 ( .C1(n4731), .C2(n4549), .A(n4548), .B(n4547), .ZN(U3516)
         );
  MUX2_X1 U5077 ( .A(REG0_REG_29__SCAN_IN), .B(n4550), .S(n4731), .Z(U3515) );
  MUX2_X1 U5078 ( .A(REG0_REG_27__SCAN_IN), .B(n4551), .S(n4731), .Z(U3513) );
  INV_X1 U5079 ( .A(REG0_REG_26__SCAN_IN), .ZN(n4553) );
  MUX2_X1 U5080 ( .A(n4553), .B(n4552), .S(n4731), .Z(n4554) );
  OAI21_X1 U5081 ( .B1(n4555), .B2(n4606), .A(n4554), .ZN(U3512) );
  INV_X1 U5082 ( .A(REG0_REG_25__SCAN_IN), .ZN(n4557) );
  OAI21_X1 U5083 ( .B1(n4559), .B2(n4606), .A(n4558), .ZN(U3511) );
  INV_X1 U5084 ( .A(REG0_REG_24__SCAN_IN), .ZN(n4561) );
  MUX2_X1 U5085 ( .A(n4561), .B(n4560), .S(n4731), .Z(n4562) );
  OAI21_X1 U5086 ( .B1(n4563), .B2(n4606), .A(n4562), .ZN(U3510) );
  INV_X1 U5087 ( .A(REG0_REG_23__SCAN_IN), .ZN(n4565) );
  MUX2_X1 U5088 ( .A(n4565), .B(n4564), .S(n4731), .Z(n4566) );
  OAI21_X1 U5089 ( .B1(n4567), .B2(n4606), .A(n4566), .ZN(U3509) );
  MUX2_X1 U5090 ( .A(REG0_REG_22__SCAN_IN), .B(n4568), .S(n4731), .Z(U3508) );
  INV_X1 U5091 ( .A(REG0_REG_21__SCAN_IN), .ZN(n4570) );
  MUX2_X1 U5092 ( .A(n4570), .B(n4569), .S(n4731), .Z(n4571) );
  OAI21_X1 U5093 ( .B1(n4572), .B2(n4606), .A(n4571), .ZN(U3507) );
  INV_X1 U5094 ( .A(REG0_REG_20__SCAN_IN), .ZN(n4574) );
  MUX2_X1 U5095 ( .A(n4574), .B(n4573), .S(n4731), .Z(n4575) );
  OAI21_X1 U5096 ( .B1(n4576), .B2(n4606), .A(n4575), .ZN(U3506) );
  INV_X1 U5097 ( .A(REG0_REG_19__SCAN_IN), .ZN(n4578) );
  MUX2_X1 U5098 ( .A(n4578), .B(n4577), .S(n4731), .Z(n4579) );
  OAI21_X1 U5099 ( .B1(n4580), .B2(n4606), .A(n4579), .ZN(U3505) );
  MUX2_X1 U5100 ( .A(REG0_REG_18__SCAN_IN), .B(n4581), .S(n4731), .Z(U3503) );
  INV_X1 U5101 ( .A(REG0_REG_17__SCAN_IN), .ZN(n4583) );
  MUX2_X1 U5102 ( .A(n4583), .B(n4582), .S(n4731), .Z(n4584) );
  OAI21_X1 U5103 ( .B1(n4585), .B2(n4606), .A(n4584), .ZN(U3501) );
  MUX2_X1 U5104 ( .A(REG0_REG_16__SCAN_IN), .B(n4586), .S(n4731), .Z(U3499) );
  INV_X1 U5105 ( .A(REG0_REG_15__SCAN_IN), .ZN(n4588) );
  MUX2_X1 U5106 ( .A(n4588), .B(n4587), .S(n4731), .Z(n4589) );
  OAI21_X1 U5107 ( .B1(n4590), .B2(n4606), .A(n4589), .ZN(U3497) );
  INV_X1 U5108 ( .A(REG0_REG_14__SCAN_IN), .ZN(n4592) );
  MUX2_X1 U5109 ( .A(n4592), .B(n4591), .S(n4731), .Z(n4593) );
  OAI21_X1 U5110 ( .B1(n4594), .B2(n4606), .A(n4593), .ZN(U3495) );
  INV_X1 U5111 ( .A(REG0_REG_13__SCAN_IN), .ZN(n4596) );
  MUX2_X1 U5112 ( .A(n4596), .B(n4595), .S(n4731), .Z(n4597) );
  OAI21_X1 U5113 ( .B1(n4598), .B2(n4606), .A(n4597), .ZN(U3493) );
  INV_X1 U5114 ( .A(REG0_REG_12__SCAN_IN), .ZN(n4600) );
  MUX2_X1 U5115 ( .A(n4600), .B(n4599), .S(n4731), .Z(n4601) );
  OAI21_X1 U5116 ( .B1(n4602), .B2(n4606), .A(n4601), .ZN(U3491) );
  INV_X1 U5117 ( .A(REG0_REG_11__SCAN_IN), .ZN(n4604) );
  MUX2_X1 U5118 ( .A(n4604), .B(n4603), .S(n4731), .Z(n4605) );
  OAI21_X1 U5119 ( .B1(n4607), .B2(n4606), .A(n4605), .ZN(U3489) );
  MUX2_X1 U5120 ( .A(DATAI_30_), .B(n4608), .S(STATE_REG_SCAN_IN), .Z(U3322)
         );
  MUX2_X1 U5121 ( .A(n4609), .B(DATAI_28_), .S(U3149), .Z(U3324) );
  MUX2_X1 U5122 ( .A(DATAI_27_), .B(n4624), .S(STATE_REG_SCAN_IN), .Z(U3325)
         );
  MUX2_X1 U5123 ( .A(n4610), .B(DATAI_25_), .S(U3149), .Z(U3327) );
  MUX2_X1 U5124 ( .A(n4611), .B(DATAI_19_), .S(U3149), .Z(U3333) );
  MUX2_X1 U5125 ( .A(DATAI_16_), .B(n4612), .S(STATE_REG_SCAN_IN), .Z(U3336)
         );
  MUX2_X1 U5126 ( .A(DATAI_15_), .B(n4613), .S(STATE_REG_SCAN_IN), .Z(U3337)
         );
  MUX2_X1 U5127 ( .A(n4614), .B(DATAI_14_), .S(U3149), .Z(U3338) );
  MUX2_X1 U5128 ( .A(n4615), .B(DATAI_13_), .S(U3149), .Z(U3339) );
  MUX2_X1 U5129 ( .A(n4616), .B(DATAI_11_), .S(U3149), .Z(U3341) );
  MUX2_X1 U5130 ( .A(n4617), .B(DATAI_10_), .S(U3149), .Z(U3342) );
  MUX2_X1 U5131 ( .A(n4618), .B(DATAI_7_), .S(U3149), .Z(U3345) );
  MUX2_X1 U5132 ( .A(n4619), .B(DATAI_6_), .S(U3149), .Z(U3346) );
  MUX2_X1 U5133 ( .A(n4620), .B(DATAI_5_), .S(U3149), .Z(U3347) );
  MUX2_X1 U5134 ( .A(DATAI_4_), .B(n4621), .S(STATE_REG_SCAN_IN), .Z(U3348) );
  MUX2_X1 U5135 ( .A(n2007), .B(DATAI_2_), .S(U3149), .Z(U3350) );
  MUX2_X1 U5136 ( .A(n2932), .B(DATAI_1_), .S(U3149), .Z(U3351) );
  INV_X1 U5137 ( .A(n4626), .ZN(n4623) );
  OAI211_X1 U5138 ( .C1(REG1_REG_0__SCAN_IN), .C2(n4624), .A(n4623), .B(n4625), 
        .ZN(n4630) );
  OAI22_X1 U5139 ( .A1(n4626), .A2(n4625), .B1(n4657), .B2(REG1_REG_0__SCAN_IN), .ZN(n4627) );
  INV_X1 U5140 ( .A(n4627), .ZN(n4629) );
  AOI22_X1 U5141 ( .A1(ADDR_REG_0__SCAN_IN), .A2(n4660), .B1(
        REG3_REG_0__SCAN_IN), .B2(U3149), .ZN(n4628) );
  OAI221_X1 U5142 ( .B1(IR_REG_0__SCAN_IN), .B2(n4630), .C1(n2300), .C2(n4629), 
        .A(n4628), .ZN(U3240) );
  OAI211_X1 U5143 ( .C1(n4633), .C2(n4632), .A(n4631), .B(n4670), .ZN(n4638)
         );
  OAI211_X1 U5144 ( .C1(n4636), .C2(n4635), .A(n4634), .B(n4654), .ZN(n4637)
         );
  OAI211_X1 U5145 ( .C1(n4673), .C2(n4639), .A(n4638), .B(n4637), .ZN(n4640)
         );
  INV_X1 U5146 ( .A(n4640), .ZN(n4642) );
  OAI211_X1 U5147 ( .C1(n4644), .C2(n4643), .A(n4642), .B(n4641), .ZN(U3255)
         );
  AOI21_X1 U5148 ( .B1(n4660), .B2(ADDR_REG_17__SCAN_IN), .A(n4645), .ZN(n4656) );
  OAI21_X1 U5149 ( .B1(n4648), .B2(n4647), .A(n4646), .ZN(n4653) );
  OAI21_X1 U5150 ( .B1(n4651), .B2(n4650), .A(n4649), .ZN(n4652) );
  AOI22_X1 U5151 ( .A1(n4654), .A2(n4653), .B1(n4670), .B2(n4652), .ZN(n4655)
         );
  OAI211_X1 U5152 ( .C1(n4695), .C2(n4673), .A(n4656), .B(n4655), .ZN(U3257)
         );
  NAND2_X1 U5153 ( .A1(n4660), .A2(ADDR_REG_18__SCAN_IN), .ZN(n4663) );
  NAND2_X1 U5154 ( .A1(n4663), .A2(n4662), .ZN(n4664) );
  AOI21_X1 U5155 ( .B1(n4668), .B2(n4667), .A(n4666), .ZN(n4669) );
  NAND2_X1 U5156 ( .A1(n4670), .A2(n4669), .ZN(n4671) );
  OAI211_X1 U5157 ( .C1(n4673), .C2(n4693), .A(n4672), .B(n4671), .ZN(U3258)
         );
  INV_X1 U5158 ( .A(n4674), .ZN(n4676) );
  AOI21_X1 U5159 ( .B1(n4677), .B2(n4676), .A(n4675), .ZN(n4683) );
  AOI22_X1 U5160 ( .A1(n4680), .A2(n4679), .B1(REG3_REG_0__SCAN_IN), .B2(n4678), .ZN(n4681) );
  OAI221_X1 U5161 ( .B1(n4684), .B2(n4683), .C1(n4682), .C2(n2302), .A(n4681), 
        .ZN(U3290) );
  AND2_X1 U5162 ( .A1(D_REG_31__SCAN_IN), .A2(n4689), .ZN(U3291) );
  AND2_X1 U5163 ( .A1(D_REG_30__SCAN_IN), .A2(n4689), .ZN(U3292) );
  AND2_X1 U5164 ( .A1(D_REG_29__SCAN_IN), .A2(n4689), .ZN(U3293) );
  AND2_X1 U5165 ( .A1(D_REG_28__SCAN_IN), .A2(n4689), .ZN(U3294) );
  AND2_X1 U5166 ( .A1(D_REG_27__SCAN_IN), .A2(n4689), .ZN(U3295) );
  AND2_X1 U5167 ( .A1(D_REG_26__SCAN_IN), .A2(n4689), .ZN(U3296) );
  AND2_X1 U5168 ( .A1(D_REG_25__SCAN_IN), .A2(n4689), .ZN(U3297) );
  AND2_X1 U5169 ( .A1(D_REG_24__SCAN_IN), .A2(n4689), .ZN(U3298) );
  AND2_X1 U5170 ( .A1(D_REG_23__SCAN_IN), .A2(n4689), .ZN(U3299) );
  AND2_X1 U5171 ( .A1(D_REG_22__SCAN_IN), .A2(n4689), .ZN(U3300) );
  AND2_X1 U5172 ( .A1(D_REG_21__SCAN_IN), .A2(n4689), .ZN(U3301) );
  INV_X1 U5173 ( .A(n4689), .ZN(n4688) );
  NOR2_X1 U5174 ( .A1(n4688), .A2(n4685), .ZN(U3302) );
  AND2_X1 U5175 ( .A1(D_REG_19__SCAN_IN), .A2(n4689), .ZN(U3303) );
  AND2_X1 U5176 ( .A1(D_REG_18__SCAN_IN), .A2(n4689), .ZN(U3304) );
  AND2_X1 U5177 ( .A1(D_REG_17__SCAN_IN), .A2(n4689), .ZN(U3305) );
  AND2_X1 U5178 ( .A1(D_REG_16__SCAN_IN), .A2(n4689), .ZN(U3306) );
  NOR2_X1 U5179 ( .A1(n4688), .A2(n4686), .ZN(U3307) );
  AND2_X1 U5180 ( .A1(D_REG_14__SCAN_IN), .A2(n4689), .ZN(U3308) );
  AND2_X1 U5181 ( .A1(D_REG_13__SCAN_IN), .A2(n4689), .ZN(U3309) );
  AND2_X1 U5182 ( .A1(D_REG_12__SCAN_IN), .A2(n4689), .ZN(U3310) );
  AND2_X1 U5183 ( .A1(D_REG_11__SCAN_IN), .A2(n4689), .ZN(U3311) );
  NOR2_X1 U5184 ( .A1(n4688), .A2(n4687), .ZN(U3312) );
  AND2_X1 U5185 ( .A1(D_REG_9__SCAN_IN), .A2(n4689), .ZN(U3313) );
  AND2_X1 U5186 ( .A1(D_REG_8__SCAN_IN), .A2(n4689), .ZN(U3314) );
  AND2_X1 U5187 ( .A1(D_REG_7__SCAN_IN), .A2(n4689), .ZN(U3315) );
  AND2_X1 U5188 ( .A1(D_REG_6__SCAN_IN), .A2(n4689), .ZN(U3316) );
  AND2_X1 U5189 ( .A1(D_REG_5__SCAN_IN), .A2(n4689), .ZN(U3317) );
  AND2_X1 U5190 ( .A1(D_REG_4__SCAN_IN), .A2(n4689), .ZN(U3318) );
  AND2_X1 U5191 ( .A1(D_REG_3__SCAN_IN), .A2(n4689), .ZN(U3319) );
  AND2_X1 U5192 ( .A1(D_REG_2__SCAN_IN), .A2(n4689), .ZN(U3320) );
  OAI21_X1 U5193 ( .B1(STATE_REG_SCAN_IN), .B2(DATAI_23_), .A(n4690), .ZN(
        n4691) );
  INV_X1 U5194 ( .A(n4691), .ZN(U3329) );
  INV_X1 U5195 ( .A(DATAI_18_), .ZN(n4692) );
  AOI22_X1 U5196 ( .A1(STATE_REG_SCAN_IN), .A2(n4693), .B1(n4692), .B2(U3149), 
        .ZN(U3334) );
  INV_X1 U5197 ( .A(DATAI_17_), .ZN(n4694) );
  AOI22_X1 U5198 ( .A1(STATE_REG_SCAN_IN), .A2(n4695), .B1(n4694), .B2(U3149), 
        .ZN(U3335) );
  OAI22_X1 U5199 ( .A1(U3149), .A2(IR_REG_0__SCAN_IN), .B1(DATAI_0_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4696) );
  INV_X1 U5200 ( .A(n4696), .ZN(U3352) );
  INV_X1 U5201 ( .A(REG0_REG_0__SCAN_IN), .ZN(n4697) );
  AOI22_X1 U5202 ( .A1(n4731), .A2(n4698), .B1(n4697), .B2(n4729), .ZN(U3467)
         );
  NOR2_X1 U5203 ( .A1(n4699), .A2(n4703), .ZN(n4700) );
  AOI211_X1 U5204 ( .C1(n4721), .C2(n4702), .A(n4701), .B(n4700), .ZN(n4732)
         );
  AOI22_X1 U5205 ( .A1(n4731), .A2(n4732), .B1(n2295), .B2(n4729), .ZN(U3469)
         );
  NOR2_X1 U5206 ( .A1(n4704), .A2(n4703), .ZN(n4706) );
  AOI211_X1 U5207 ( .C1(n4721), .C2(n4707), .A(n4706), .B(n4705), .ZN(n4734)
         );
  AOI22_X1 U5208 ( .A1(n4731), .A2(n4734), .B1(n4708), .B2(n4729), .ZN(U3473)
         );
  INV_X1 U5209 ( .A(n4709), .ZN(n4711) );
  AOI211_X1 U5210 ( .C1(n4713), .C2(n4712), .A(n4711), .B(n4710), .ZN(n4736)
         );
  INV_X1 U5211 ( .A(REG0_REG_4__SCAN_IN), .ZN(n4714) );
  AOI22_X1 U5212 ( .A1(n4731), .A2(n4736), .B1(n4714), .B2(n4729), .ZN(U3475)
         );
  NOR2_X1 U5213 ( .A1(n4716), .A2(n4715), .ZN(n4719) );
  INV_X1 U5214 ( .A(n4717), .ZN(n4718) );
  AOI211_X1 U5215 ( .C1(n4721), .C2(n4720), .A(n4719), .B(n4718), .ZN(n4738)
         );
  INV_X1 U5216 ( .A(REG0_REG_5__SCAN_IN), .ZN(n4722) );
  AOI22_X1 U5217 ( .A1(n4731), .A2(n4738), .B1(n4722), .B2(n4729), .ZN(U3477)
         );
  NAND3_X1 U5218 ( .A1(n4725), .A2(n4724), .A3(n4723), .ZN(n4726) );
  AND3_X1 U5219 ( .A1(n4728), .A2(n4727), .A3(n4726), .ZN(n4740) );
  INV_X1 U5220 ( .A(REG0_REG_7__SCAN_IN), .ZN(n4730) );
  AOI22_X1 U5221 ( .A1(n4731), .A2(n4740), .B1(n4730), .B2(n4729), .ZN(U3481)
         );
  AOI22_X1 U5222 ( .A1(n4741), .A2(n4732), .B1(n2931), .B2(n2712), .ZN(U3519)
         );
  INV_X1 U5223 ( .A(REG1_REG_3__SCAN_IN), .ZN(n4733) );
  AOI22_X1 U5224 ( .A1(n4741), .A2(n4734), .B1(n4733), .B2(n2712), .ZN(U3521)
         );
  AOI22_X1 U5225 ( .A1(n4741), .A2(n4736), .B1(n4735), .B2(n2712), .ZN(U3522)
         );
  AOI22_X1 U5226 ( .A1(n4741), .A2(n4738), .B1(n4737), .B2(n2712), .ZN(U3523)
         );
  AOI22_X1 U5227 ( .A1(n4741), .A2(n4740), .B1(n4739), .B2(n2712), .ZN(U3525)
         );
endmodule

