

module b20_C_gen_AntiSAT_k_128_3 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, keyinput_f0, 
        keyinput_f1, keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5, 
        keyinput_f6, keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10, 
        keyinput_f11, keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15, 
        keyinput_f16, keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20, 
        keyinput_f21, keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25, 
        keyinput_f26, keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30, 
        keyinput_f31, keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35, 
        keyinput_f36, keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40, 
        keyinput_f41, keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45, 
        keyinput_f46, keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50, 
        keyinput_f51, keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55, 
        keyinput_f56, keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60, 
        keyinput_f61, keyinput_f62, keyinput_f63, keyinput_g0, keyinput_g1, 
        keyinput_g2, keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, 
        keyinput_g7, keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, 
        keyinput_g12, keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, 
        keyinput_g17, keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, 
        keyinput_g22, keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, 
        keyinput_g27, keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, 
        keyinput_g32, keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, 
        keyinput_g37, keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, 
        keyinput_g42, keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, 
        keyinput_g47, keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, 
        keyinput_g52, keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, 
        keyinput_g57, keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, 
        keyinput_g62, keyinput_g63, ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, 
        ADD_1068_U57, ADD_1068_U58, ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, 
        ADD_1068_U62, ADD_1068_U63, ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, 
        ADD_1068_U50, ADD_1068_U51, ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, 
        ADD_1068_U5, ADD_1068_U46, U126, U123, P1_U3355, P1_U3354, P1_U3353, 
        P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, 
        P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, 
        P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, 
        P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, 
        P1_U3324, P1_U3439, P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, 
        P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, 
        P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, 
        P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, 
        P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, 
        P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, 
        P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, 
        P1_U3501, P1_U3504, P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, 
        P1_U3513, P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, 
        P1_U3520, P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, 
        P1_U3527, P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, 
        P1_U3534, P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, 
        P1_U3541, P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, 
        P1_U3548, P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, 
        P1_U3292, P1_U3291, P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, 
        P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, 
        P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, 
        P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, 
        P1_U3356, P1_U3264, P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, 
        P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, 
        P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, 
        P1_U3244, P1_U3243, P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, 
        P1_U3559, P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, 
        P1_U3566, P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, 
        P1_U3573, P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, 
        P1_U3580, P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, 
        P1_U3241, P1_U3240, P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, 
        P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, 
        P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, 
        P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, 
        P1_U3213, P1_U3086, P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, 
        P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, 
        P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, 
        P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, 
        P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, 
        P2_U3264, P2_U3376, P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, 
        P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, 
        P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, 
        P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, 
        P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, 
        P2_U3396, P2_U3399, P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, 
        P2_U3417, P2_U3420, P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, 
        P2_U3438, P2_U3441, P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, 
        P2_U3450, P2_U3451, P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, 
        P2_U3457, P2_U3458, P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, 
        P2_U3464, P2_U3465, P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, 
        P2_U3471, P2_U3472, P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, 
        P2_U3478, P2_U3479, P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, 
        P2_U3485, P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, 
        P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, 
        P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, 
        P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, 
        P2_U3211, P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, 
        P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, 
        P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, 
        P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, 
        P2_U3183, P2_U3182, P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, 
        P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, 
        P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, 
        P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, 
        P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, 
        P2_U3181, P2_U3180, P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, 
        P2_U3174, P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, 
        P2_U3167, P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, 
        P2_U3160, P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, 
        P2_U3153, P2_U3151, P2_U3150, P2_U3893 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, keyinput_f0, keyinput_f1, keyinput_f2,
         keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, keyinput_f7,
         keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, keyinput_f12,
         keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, keyinput_f17,
         keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, keyinput_f22,
         keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, keyinput_f27,
         keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, keyinput_f32,
         keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, keyinput_f37,
         keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, keyinput_f42,
         keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, keyinput_f47,
         keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, keyinput_f52,
         keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, keyinput_f57,
         keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, keyinput_f62,
         keyinput_f63, keyinput_g0, keyinput_g1, keyinput_g2, keyinput_g3,
         keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7, keyinput_g8,
         keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12, keyinput_g13,
         keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17, keyinput_g18,
         keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22, keyinput_g23,
         keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27, keyinput_g28,
         keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32, keyinput_g33,
         keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37, keyinput_g38,
         keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42, keyinput_g43,
         keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47, keyinput_g48,
         keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52, keyinput_g53,
         keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57, keyinput_g58,
         keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62, keyinput_g63;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4351, n4352, n4353, n4354, n4355, n4357, n4358, n4359, n4360, n4361,
         n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371,
         n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381,
         n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391,
         n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401,
         n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411,
         n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421,
         n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431,
         n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441,
         n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451,
         n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461,
         n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471,
         n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481,
         n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491,
         n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501,
         n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511,
         n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521,
         n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531,
         n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541,
         n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551,
         n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561,
         n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571,
         n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581,
         n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591,
         n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601,
         n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611,
         n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621,
         n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631,
         n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641,
         n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651,
         n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661,
         n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671,
         n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681,
         n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691,
         n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701,
         n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711,
         n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721,
         n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731,
         n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741,
         n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751,
         n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761,
         n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771,
         n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781,
         n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791,
         n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801,
         n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811,
         n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821,
         n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831,
         n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841,
         n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851,
         n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861,
         n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871,
         n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881,
         n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891,
         n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901,
         n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911,
         n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921,
         n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931,
         n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941,
         n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951,
         n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961,
         n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971,
         n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981,
         n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991,
         n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001,
         n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011,
         n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021,
         n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031,
         n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041,
         n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051,
         n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061,
         n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071,
         n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081,
         n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091,
         n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101,
         n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111,
         n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121,
         n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131,
         n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141,
         n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151,
         n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161,
         n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171,
         n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181,
         n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191,
         n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201,
         n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211,
         n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221,
         n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231,
         n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241,
         n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251,
         n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261,
         n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271,
         n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281,
         n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291,
         n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301,
         n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311,
         n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321,
         n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331,
         n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341,
         n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351,
         n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361,
         n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371,
         n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381,
         n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391,
         n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401,
         n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411,
         n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421,
         n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431,
         n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441,
         n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451,
         n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461,
         n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471,
         n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481,
         n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491,
         n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501,
         n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511,
         n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521,
         n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531,
         n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541,
         n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551,
         n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561,
         n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571,
         n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581,
         n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591,
         n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601,
         n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611,
         n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621,
         n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631,
         n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641,
         n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651,
         n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661,
         n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671,
         n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681,
         n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691,
         n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701,
         n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711,
         n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721,
         n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731,
         n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741,
         n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751,
         n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761,
         n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771,
         n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781,
         n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791,
         n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801,
         n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811,
         n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821,
         n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831,
         n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841,
         n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851,
         n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861,
         n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871,
         n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881,
         n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891,
         n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901,
         n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911,
         n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921,
         n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931,
         n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941,
         n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951,
         n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961,
         n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971,
         n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981,
         n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991,
         n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001,
         n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011,
         n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021,
         n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031,
         n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041,
         n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051,
         n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061,
         n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071,
         n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081,
         n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091,
         n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101,
         n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111,
         n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121,
         n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131,
         n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141,
         n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151,
         n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161,
         n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171,
         n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181,
         n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191,
         n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201,
         n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211,
         n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221,
         n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231,
         n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241,
         n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251,
         n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261,
         n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271,
         n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281,
         n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291,
         n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301,
         n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311,
         n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321,
         n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331,
         n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341,
         n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351,
         n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361,
         n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371,
         n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381,
         n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391,
         n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401,
         n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411,
         n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421,
         n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431,
         n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441,
         n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451,
         n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461,
         n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471,
         n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481,
         n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491,
         n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501,
         n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511,
         n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521,
         n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531,
         n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541,
         n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551,
         n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561,
         n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571,
         n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581,
         n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591,
         n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601,
         n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611,
         n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621,
         n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631,
         n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641,
         n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651,
         n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661,
         n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671,
         n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681,
         n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691,
         n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701,
         n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711,
         n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721,
         n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731,
         n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741,
         n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751,
         n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761,
         n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771,
         n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781,
         n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791,
         n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801,
         n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811,
         n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821,
         n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831,
         n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841,
         n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851,
         n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861,
         n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871,
         n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881,
         n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891,
         n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901,
         n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911,
         n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921,
         n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931,
         n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941,
         n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951,
         n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961,
         n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971,
         n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981,
         n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991,
         n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001,
         n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011,
         n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021,
         n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031,
         n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041,
         n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051,
         n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061,
         n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071,
         n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081,
         n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091,
         n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101,
         n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111,
         n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121,
         n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131,
         n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141,
         n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151,
         n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161,
         n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171,
         n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181,
         n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191,
         n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201,
         n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211,
         n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221,
         n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231,
         n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241,
         n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251,
         n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261,
         n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271,
         n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281,
         n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291,
         n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301,
         n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311,
         n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321,
         n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331,
         n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341,
         n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351,
         n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361,
         n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371,
         n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381,
         n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391,
         n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401,
         n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411,
         n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421,
         n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431,
         n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441,
         n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451,
         n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461,
         n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471,
         n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481,
         n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491,
         n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501,
         n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511,
         n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521,
         n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531,
         n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541,
         n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551,
         n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561,
         n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571,
         n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581,
         n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591,
         n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601,
         n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611,
         n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621,
         n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631,
         n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641,
         n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651,
         n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661,
         n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671,
         n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681,
         n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691,
         n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701,
         n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711,
         n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721,
         n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731,
         n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741,
         n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751,
         n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761,
         n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771,
         n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781,
         n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791,
         n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801,
         n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811,
         n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821,
         n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831,
         n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841,
         n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851,
         n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861,
         n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871,
         n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881,
         n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891,
         n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901,
         n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911,
         n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921,
         n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931,
         n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941,
         n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951,
         n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961,
         n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971,
         n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981,
         n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991,
         n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001,
         n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011,
         n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021,
         n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031,
         n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041,
         n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051,
         n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061,
         n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071,
         n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081,
         n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091,
         n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101,
         n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111,
         n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121,
         n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131,
         n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141,
         n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151,
         n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161,
         n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171,
         n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181,
         n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191,
         n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201,
         n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211,
         n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221,
         n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231,
         n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241,
         n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251,
         n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261,
         n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271,
         n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281,
         n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291,
         n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301,
         n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311,
         n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321,
         n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331,
         n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341,
         n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351,
         n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361,
         n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371,
         n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381,
         n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391,
         n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401,
         n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411,
         n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421,
         n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431,
         n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441,
         n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451,
         n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461,
         n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471,
         n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481,
         n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491,
         n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501,
         n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511,
         n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521,
         n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531,
         n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541,
         n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551,
         n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561,
         n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571,
         n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581,
         n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591,
         n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601,
         n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611,
         n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621,
         n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631,
         n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641,
         n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651,
         n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661,
         n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671,
         n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681,
         n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691,
         n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701,
         n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711,
         n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721,
         n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731,
         n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741,
         n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751,
         n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761,
         n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771,
         n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781,
         n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791,
         n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801,
         n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811,
         n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821,
         n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831,
         n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841,
         n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851,
         n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861,
         n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871,
         n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881,
         n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891,
         n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901,
         n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911,
         n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921,
         n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931,
         n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941,
         n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951,
         n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961,
         n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971,
         n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981,
         n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991,
         n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001,
         n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011,
         n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021,
         n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031,
         n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041,
         n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051,
         n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061,
         n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071,
         n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081,
         n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091,
         n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101,
         n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111,
         n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121,
         n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131,
         n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141,
         n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151,
         n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161,
         n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171,
         n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181,
         n9182, n9183, n9184, n9185, n9187, n9188, n9189, n9190, n9191, n9192,
         n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202,
         n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212,
         n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222,
         n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232,
         n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242,
         n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252,
         n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262,
         n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272,
         n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282,
         n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292,
         n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302,
         n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312,
         n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322,
         n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332,
         n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342,
         n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352,
         n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362,
         n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372,
         n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382,
         n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392,
         n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402,
         n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412,
         n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422,
         n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432,
         n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442,
         n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452,
         n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462,
         n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472,
         n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482,
         n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492,
         n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502,
         n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512,
         n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522,
         n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532,
         n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542,
         n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552,
         n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562,
         n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572,
         n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582,
         n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
         n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602,
         n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
         n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
         n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
         n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
         n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
         n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
         n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
         n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
         n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
         n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
         n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
         n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
         n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
         n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
         n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
         n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
         n10122, n10123, n10124, n10125, n10126, n10127;

  INV_X1 U4854 ( .A(P2_STATE_REG_SCAN_IN), .ZN(n9917) );
  CLKBUF_X2 U4855 ( .A(n4917), .Z(n4354) );
  INV_X1 U4856 ( .A(n5188), .ZN(n5265) );
  AND2_X1 U4857 ( .A1(n8658), .A2(n8731), .ZN(n8734) );
  CLKBUF_X2 U4858 ( .A(n5933), .Z(n8578) );
  INV_X1 U4859 ( .A(n5552), .ZN(n7751) );
  CLKBUF_X3 U4860 ( .A(n5858), .Z(n4353) );
  XNOR2_X1 U4861 ( .A(n4355), .B(n6669), .ZN(n5778) );
  CLKBUF_X2 U4862 ( .A(n5416), .Z(n5677) );
  NAND4_X1 U4863 ( .A1(n5909), .A2(n5908), .A3(n5907), .A4(n5906), .ZN(n8756)
         );
  CLKBUF_X2 U4864 ( .A(n5992), .Z(n4362) );
  CLKBUF_X2 U4865 ( .A(n5992), .Z(n4363) );
  INV_X1 U4868 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  INV_X1 U4870 ( .A(n5334), .ZN(n5340) );
  INV_X1 U4871 ( .A(n7732), .ZN(n7747) );
  INV_X1 U4872 ( .A(n8745), .ZN(n9010) );
  INV_X1 U4873 ( .A(n6978), .ZN(n9541) );
  BUF_X1 U4874 ( .A(n5163), .Z(n4358) );
  NAND2_X1 U4875 ( .A1(n4960), .A2(n4959), .ZN(n5108) );
  AND2_X1 U4876 ( .A1(n8187), .A2(n7701), .ZN(n8200) );
  XNOR2_X1 U4877 ( .A(n5108), .B(n5109), .ZN(n6481) );
  INV_X1 U4878 ( .A(n8486), .ZN(n9567) );
  INV_X1 U4879 ( .A(n8490), .ZN(n8752) );
  INV_X2 U4880 ( .A(n9510), .ZN(n9485) );
  AND4_X1 U4881 ( .A1(n5030), .A2(n5029), .A3(n5028), .A4(n5027), .ZN(n4351)
         );
  INV_X1 U4882 ( .A(n6436), .ZN(n4352) );
  AOI21_X2 U4883 ( .B1(n7897), .B2(n7898), .A(n6374), .ZN(n7901) );
  OAI21_X2 U4884 ( .B1(n5564), .B2(P2_IR_REG_18__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5565) );
  XNOR2_X2 U4885 ( .A(n5279), .B(P1_IR_REG_30__SCAN_IN), .ZN(n5903) );
  OR2_X2 U4886 ( .A1(n9185), .A2(n5278), .ZN(n5279) );
  XNOR2_X2 U4887 ( .A(n5733), .B(P2_IR_REG_25__SCAN_IN), .ZN(n7228) );
  NOR2_X2 U4888 ( .A1(n4467), .A2(n5688), .ZN(n5734) );
  NAND2_X1 U4889 ( .A1(n5793), .A2(n5792), .ZN(n6780) );
  AND2_X1 U4890 ( .A1(n5132), .A2(n5131), .ZN(n9601) );
  NAND2_X1 U4891 ( .A1(n5117), .A2(n5116), .ZN(n7475) );
  NAND2_X1 U4892 ( .A1(n8678), .A2(n8478), .ZN(n7154) );
  NAND2_X1 U4893 ( .A1(n8752), .A2(n9567), .ZN(n8475) );
  INV_X1 U4894 ( .A(n7054), .ZN(n9548) );
  NAND2_X1 U4895 ( .A1(n7613), .A2(n7617), .ZN(n6661) );
  INV_X1 U4896 ( .A(n6872), .ZN(n9747) );
  NAND4_X1 U4897 ( .A1(n5384), .A2(n5383), .A3(n5382), .A4(n5381), .ZN(n9745)
         );
  INV_X1 U4898 ( .A(n6970), .ZN(n6969) );
  NAND2_X4 U4899 ( .A1(n6285), .A2(n6325), .ZN(n6307) );
  BUF_X2 U4900 ( .A(n5426), .Z(n7752) );
  INV_X4 U4901 ( .A(n6436), .ZN(n4923) );
  NOR3_X1 U4902 ( .A1(n7935), .A2(n7900), .A3(n7899), .ZN(n7902) );
  AND2_X1 U4903 ( .A1(n6380), .A2(n6379), .ZN(n6381) );
  NAND2_X1 U4904 ( .A1(n4704), .A2(n7932), .ZN(n5854) );
  OR2_X1 U4905 ( .A1(n7746), .A2(n7745), .ZN(n7750) );
  NAND2_X1 U4906 ( .A1(n4637), .A2(n9493), .ZN(n4644) );
  NAND2_X1 U4907 ( .A1(n5839), .A2(n5838), .ZN(n7889) );
  AOI21_X1 U4908 ( .B1(n8925), .B2(n9493), .A(n8924), .ZN(n9111) );
  NAND2_X1 U4909 ( .A1(n4493), .A2(n4723), .ZN(n4724) );
  NOR2_X1 U4910 ( .A1(n8419), .A2(n8421), .ZN(n8423) );
  NAND2_X1 U4911 ( .A1(n8148), .A2(n5605), .ZN(n8137) );
  AOI21_X1 U4912 ( .B1(n4621), .B2(n4623), .A(n4619), .ZN(n4618) );
  AOI21_X1 U4913 ( .B1(n9591), .B2(n9109), .A(n9108), .ZN(n9110) );
  NAND2_X1 U4914 ( .A1(n7448), .A2(n7447), .ZN(n7446) );
  NAND2_X1 U4915 ( .A1(n4657), .A2(n4656), .ZN(n6120) );
  NAND2_X1 U4916 ( .A1(n5555), .A2(n5554), .ZN(n8310) );
  AND2_X1 U4917 ( .A1(n5212), .A2(n5211), .ZN(n9017) );
  NAND2_X1 U4918 ( .A1(n5217), .A2(n5216), .ZN(n9140) );
  NAND2_X1 U4919 ( .A1(n7401), .A2(n7400), .ZN(n7567) );
  INV_X1 U4920 ( .A(n9068), .ZN(n7829) );
  XNOR2_X1 U4921 ( .A(n5210), .B(n5209), .ZN(n6832) );
  NAND2_X1 U4922 ( .A1(n5543), .A2(n5542), .ZN(n8317) );
  AOI21_X1 U4923 ( .B1(n5178), .B2(n5177), .A(n4979), .ZN(n5184) );
  OAI21_X1 U4924 ( .B1(n6575), .B2(n6574), .A(n5779), .ZN(n6585) );
  NOR2_X1 U4925 ( .A1(n7157), .A2(n7156), .ZN(n7158) );
  NAND2_X1 U4926 ( .A1(n5107), .A2(n5106), .ZN(n7343) );
  OAI21_X2 U4927 ( .B1(n6459), .B2(n5188), .A(n4477), .ZN(n8491) );
  NAND2_X1 U4928 ( .A1(n7640), .A2(n7632), .ZN(n6790) );
  CLKBUF_X1 U4929 ( .A(n8430), .Z(n8460) );
  OAI21_X1 U4930 ( .B1(n6341), .B2(n9500), .A(n9499), .ZN(n8430) );
  NOR2_X1 U4931 ( .A1(n4568), .A2(n4573), .ZN(n4478) );
  NOR2_X1 U4932 ( .A1(n4569), .A2(n4390), .ZN(n4568) );
  OAI211_X1 U4933 ( .C1(n5052), .C2(n6447), .A(n5073), .B(n5072), .ZN(n6978)
         );
  INV_X1 U4934 ( .A(n9761), .ZN(n8004) );
  NAND2_X1 U4935 ( .A1(n5776), .A2(n5775), .ZN(n5858) );
  INV_X2 U4936 ( .A(n6463), .ZN(n6493) );
  NAND3_X1 U4937 ( .A1(n4571), .A2(n4951), .A3(n4570), .ZN(n5099) );
  AND4_X1 U4938 ( .A1(n5405), .A2(n5404), .A3(n5403), .A4(n5402), .ZN(n6872)
         );
  AND3_X1 U4939 ( .A1(n5954), .A2(n5953), .A3(n5952), .ZN(n6896) );
  INV_X2 U4940 ( .A(n6285), .ZN(n6321) );
  NOR2_X1 U4941 ( .A1(n8005), .A2(n7814), .ZN(n9729) );
  AND3_X1 U4942 ( .A1(n5936), .A2(n5935), .A3(n5934), .ZN(n5938) );
  NAND4_X2 U4943 ( .A1(n5926), .A2(n5925), .A3(n5924), .A4(n5923), .ZN(n6898)
         );
  AND4_X1 U4944 ( .A1(n5983), .A2(n5982), .A3(n5981), .A4(n5980), .ZN(n7160)
         );
  OR2_X1 U4945 ( .A1(n4573), .A2(n4572), .ZN(n4571) );
  AND2_X2 U4946 ( .A1(n5340), .A2(n7495), .ZN(n5599) );
  AND3_X2 U4947 ( .A1(n5045), .A2(n5044), .A3(n5043), .ZN(n6897) );
  INV_X2 U4948 ( .A(n5904), .ZN(n5958) );
  INV_X1 U4949 ( .A(n4949), .ZN(n4573) );
  INV_X1 U4950 ( .A(n5753), .ZN(n7259) );
  NAND2_X1 U4951 ( .A1(n5379), .A2(n6436), .ZN(n5552) );
  OR2_X1 U4952 ( .A1(n4948), .A2(n5086), .ZN(n4949) );
  AND2_X1 U4953 ( .A1(n9308), .A2(n8793), .ZN(n9309) );
  NAND2_X2 U4954 ( .A1(n5304), .A2(n5295), .ZN(n6408) );
  OR2_X1 U4955 ( .A1(n8020), .A2(n7807), .ZN(n5774) );
  NAND2_X1 U4956 ( .A1(n9503), .A2(n6854), .ZN(n6892) );
  AND2_X1 U4957 ( .A1(n5301), .A2(n5315), .ZN(n5295) );
  XNOR2_X1 U4958 ( .A(n5202), .B(n5201), .ZN(n9503) );
  XNOR2_X1 U4959 ( .A(n5332), .B(P2_IR_REG_29__SCAN_IN), .ZN(n7495) );
  NAND2_X1 U4960 ( .A1(n5345), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5347) );
  OR2_X1 U4961 ( .A1(n5331), .A2(n5330), .ZN(n5332) );
  NAND2_X4 U4962 ( .A1(n5286), .A2(n5287), .ZN(n5052) );
  XNOR2_X1 U4963 ( .A(n5687), .B(P2_IR_REG_21__SCAN_IN), .ZN(n7808) );
  NAND2_X1 U4964 ( .A1(n5200), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5202) );
  XNOR2_X1 U4965 ( .A(n5274), .B(n4894), .ZN(n6854) );
  OR2_X1 U4966 ( .A1(n5277), .A2(n5278), .ZN(n5034) );
  XNOR2_X1 U4967 ( .A(n5272), .B(P1_IR_REG_21__SCAN_IN), .ZN(n8735) );
  AND2_X1 U4968 ( .A1(n4351), .A2(n4893), .ZN(n4476) );
  AND2_X1 U4969 ( .A1(n4895), .A2(n4894), .ZN(n4893) );
  AND3_X1 U4970 ( .A1(n4709), .A2(n4708), .A3(n5318), .ZN(n5393) );
  AND2_X1 U4971 ( .A1(n5025), .A2(n5026), .ZN(n4895) );
  INV_X4 U4972 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X1 U4973 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n4918) );
  NOR2_X2 U4974 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .ZN(
        n4896) );
  INV_X1 U4975 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5024) );
  NOR2_X1 U4976 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_9__SCAN_IN), .ZN(
        n4705) );
  NOR2_X1 U4977 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(P2_IR_REG_6__SCAN_IN), .ZN(
        n4706) );
  NOR2_X1 U4978 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .ZN(
        n4707) );
  NOR3_X1 U4979 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .A3(
        P2_IR_REG_10__SCAN_IN), .ZN(n5319) );
  NOR2_X2 U4980 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n5061) );
  NOR2_X1 U4981 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n5025) );
  NOR2_X1 U4982 ( .A1(P1_IR_REG_23__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), .ZN(
        n5031) );
  NOR3_X1 U4983 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_16__SCAN_IN), .A3(
        P1_IR_REG_18__SCAN_IN), .ZN(n5030) );
  XNOR2_X2 U4984 ( .A(n5804), .B(n7389), .ZN(n7277) );
  INV_X4 U4985 ( .A(n6307), .ZN(n6284) );
  NOR3_X2 U4986 ( .A1(n8989), .A2(n4490), .A3(n9119), .ZN(n4492) );
  INV_X1 U4987 ( .A(n6669), .ZN(n9779) );
  NAND2_X1 U4988 ( .A1(n6669), .A2(n9763), .ZN(n7613) );
  INV_X1 U4991 ( .A(n4355), .ZN(n5801) );
  INV_X2 U4992 ( .A(n9534), .ZN(n6974) );
  OAI211_X2 U4993 ( .C1(n5052), .C2(n8776), .A(n5060), .B(n5059), .ZN(n9534)
         );
  OAI21_X2 U4994 ( .B1(n5738), .B2(n7228), .A(n7259), .ZN(n5739) );
  AND2_X4 U4995 ( .A1(n5903), .A2(n5282), .ZN(n5959) );
  NAND2_X1 U4996 ( .A1(n6408), .A2(n5910), .ZN(n4917) );
  INV_X1 U4997 ( .A(n5904), .ZN(n4359) );
  INV_X1 U4998 ( .A(n5904), .ZN(n4360) );
  CLKBUF_X1 U4999 ( .A(n5992), .Z(n4361) );
  AND2_X1 U5000 ( .A1(n5903), .A2(n5902), .ZN(n5992) );
  INV_X1 U5001 ( .A(n5649), .ZN(n4797) );
  OR2_X1 U5002 ( .A1(n8267), .A2(n7938), .ZN(n7729) );
  INV_X1 U5003 ( .A(n8367), .ZN(n4688) );
  NAND2_X1 U5004 ( .A1(n9083), .A2(n9061), .ZN(n8465) );
  OR2_X1 U5005 ( .A1(n9083), .A2(n9061), .ZN(n8528) );
  OR2_X1 U5006 ( .A1(n6276), .A2(n6275), .ZN(n6311) );
  AOI21_X1 U5007 ( .B1(n4866), .B2(n4868), .A(n4412), .ZN(n4864) );
  AOI21_X1 U5008 ( .B1(n8525), .B2(n8524), .A(n8701), .ZN(n4586) );
  NAND2_X1 U5009 ( .A1(n7717), .A2(n4525), .ZN(n4524) );
  AND2_X1 U5010 ( .A1(n7716), .A2(n7747), .ZN(n4525) );
  AND2_X1 U5011 ( .A1(n9904), .A2(n5206), .ZN(n4990) );
  AND2_X1 U5012 ( .A1(n8304), .A2(n7947), .ZN(n7711) );
  AOI21_X1 U5013 ( .B1(P2_REG2_REG_6__SCAN_IN), .B2(n6920), .A(n6919), .ZN(
        n6921) );
  NAND2_X1 U5014 ( .A1(n6984), .A2(n5466), .ZN(n4542) );
  NAND2_X1 U5015 ( .A1(n5434), .A2(n6863), .ZN(n5435) );
  AOI21_X1 U5016 ( .B1(n4796), .B2(n4794), .A(n4439), .ZN(n4793) );
  INV_X1 U5017 ( .A(n5648), .ZN(n4794) );
  NOR2_X1 U5018 ( .A1(n4913), .A2(n4787), .ZN(n4786) );
  INV_X1 U5019 ( .A(n5616), .ZN(n4787) );
  OR2_X1 U5020 ( .A1(n7916), .A2(n7985), .ZN(n7609) );
  AND2_X1 U5021 ( .A1(n6255), .A2(n6254), .ZN(n6257) );
  OAI21_X1 U5022 ( .B1(n6284), .B2(n6897), .A(n5927), .ZN(n4661) );
  AOI22_X1 U5023 ( .A1(n6898), .A2(n6287), .B1(n7030), .B2(n6323), .ZN(n5930)
         );
  NOR2_X1 U5024 ( .A1(n9075), .A2(n4891), .ZN(n4890) );
  INV_X1 U5025 ( .A(n7826), .ZN(n4891) );
  OR2_X1 U5026 ( .A1(n9590), .A2(n7472), .ZN(n8511) );
  OR2_X1 U5027 ( .A1(n6067), .A2(n6066), .ZN(n6069) );
  OAI21_X1 U5028 ( .B1(n5215), .B2(n4995), .A(n4994), .ZN(n5219) );
  NOR2_X1 U5029 ( .A1(n4977), .A2(n4976), .ZN(n5178) );
  NOR2_X1 U5030 ( .A1(n4975), .A2(n4974), .ZN(n4976) );
  AND2_X1 U5031 ( .A1(n4941), .A2(n5077), .ZN(n4732) );
  NAND4_X2 U5032 ( .A1(n4896), .A2(n5061), .A3(n5048), .A4(n5024), .ZN(n5082)
         );
  AND2_X1 U5033 ( .A1(n5774), .A2(n5773), .ZN(n5775) );
  NAND2_X1 U5034 ( .A1(n5772), .A2(n5771), .ZN(n5776) );
  OR2_X1 U5035 ( .A1(n5868), .A2(n6379), .ZN(n5871) );
  NAND2_X1 U5036 ( .A1(n6618), .A2(n4401), .ZN(n6675) );
  AND2_X1 U5037 ( .A1(n5635), .A2(n5634), .ZN(n7938) );
  NAND2_X1 U5038 ( .A1(n6808), .A2(n6807), .ZN(n6916) );
  XNOR2_X1 U5039 ( .A(n8031), .B(n8030), .ZN(n9734) );
  NOR2_X1 U5040 ( .A1(n5501), .A2(n5500), .ZN(n5502) );
  NAND2_X1 U5041 ( .A1(n4539), .A2(n4905), .ZN(n7346) );
  OR2_X1 U5042 ( .A1(n7394), .A2(n7451), .ZN(n4905) );
  NAND2_X1 U5043 ( .A1(n7219), .A2(n4800), .ZN(n4539) );
  OR2_X1 U5044 ( .A1(n9825), .A2(n7999), .ZN(n4800) );
  AND2_X1 U5045 ( .A1(n5379), .A2(n4923), .ZN(n5426) );
  AOI21_X1 U5046 ( .B1(n8099), .B2(n7728), .A(n5720), .ZN(n8091) );
  INV_X1 U5047 ( .A(n4786), .ZN(n4783) );
  AND2_X1 U5048 ( .A1(n4781), .A2(n4784), .ZN(n4780) );
  NAND2_X1 U5049 ( .A1(n4786), .A2(n4782), .ZN(n4781) );
  OAI21_X1 U5050 ( .B1(n5615), .B2(n4406), .A(n4785), .ZN(n4784) );
  INV_X1 U5051 ( .A(n5605), .ZN(n4782) );
  OR2_X1 U5052 ( .A1(n8317), .A2(n7994), .ZN(n8187) );
  INV_X1 U5053 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5447) );
  NAND2_X1 U5054 ( .A1(n4679), .A2(n4678), .ZN(n7596) );
  NAND2_X1 U5055 ( .A1(n4374), .A2(n4684), .ZN(n4678) );
  AND2_X1 U5056 ( .A1(n4374), .A2(n8399), .ZN(n4680) );
  NAND2_X1 U5057 ( .A1(n6008), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n6027) );
  OR2_X1 U5058 ( .A1(n6233), .A2(n6232), .ZN(n6248) );
  AND2_X1 U5059 ( .A1(n6283), .A2(n6282), .ZN(n8876) );
  INV_X1 U5060 ( .A(n5959), .ZN(n6337) );
  NAND2_X1 U5061 ( .A1(n4604), .A2(n4603), .ZN(n4602) );
  NAND2_X1 U5062 ( .A1(n9318), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n4603) );
  NAND2_X1 U5063 ( .A1(n5269), .A2(n5268), .ZN(n8587) );
  OAI21_X1 U5064 ( .B1(n4881), .B2(n4880), .A(n4393), .ZN(n4879) );
  NAND2_X1 U5065 ( .A1(n5176), .A2(n5175), .ZN(n9083) );
  INV_X1 U5066 ( .A(n5267), .ZN(n5203) );
  NAND2_X1 U5067 ( .A1(n7160), .A2(n7054), .ZN(n8478) );
  NAND2_X1 U5068 ( .A1(n6934), .A2(n6897), .ZN(n6899) );
  XNOR2_X1 U5069 ( .A(n5281), .B(P1_IR_REG_29__SCAN_IN), .ZN(n5902) );
  INV_X1 U5070 ( .A(n6402), .ZN(n4692) );
  AND2_X1 U5071 ( .A1(n4791), .A2(n4789), .ZN(n5684) );
  OAI21_X1 U5072 ( .B1(n7616), .B2(n4520), .A(n4518), .ZN(n7618) );
  NAND2_X1 U5073 ( .A1(n4519), .A2(n7747), .ZN(n4518) );
  NAND2_X1 U5074 ( .A1(n7617), .A2(n7817), .ZN(n4520) );
  NAND2_X1 U5075 ( .A1(n8693), .A2(n8509), .ZN(n4450) );
  NAND2_X1 U5076 ( .A1(n4582), .A2(n9052), .ZN(n8543) );
  INV_X1 U5077 ( .A(n4584), .ZN(n4583) );
  OAI21_X1 U5078 ( .B1(n8529), .B2(n4586), .A(n8734), .ZN(n4585) );
  AND2_X1 U5079 ( .A1(n8200), .A2(n7698), .ZN(n4513) );
  AOI21_X1 U5080 ( .B1(n8555), .B2(n8977), .A(n4565), .ZN(n4564) );
  NAND2_X1 U5081 ( .A1(n4508), .A2(n4506), .ZN(n7703) );
  NAND2_X1 U5082 ( .A1(n8464), .A2(n8465), .ZN(n8527) );
  NAND2_X1 U5083 ( .A1(n4522), .A2(n4521), .ZN(n7722) );
  AND2_X1 U5084 ( .A1(n7721), .A2(n7770), .ZN(n4521) );
  OAI21_X1 U5085 ( .B1(n8568), .B2(n8567), .A(n8566), .ZN(n8569) );
  AND2_X1 U5086 ( .A1(n4852), .A2(n7762), .ZN(n4849) );
  OAI21_X1 U5087 ( .B1(n4499), .B2(n4498), .A(n4495), .ZN(n4494) );
  NAND2_X1 U5088 ( .A1(n7725), .A2(n8117), .ZN(n4498) );
  NOR2_X1 U5089 ( .A1(n4497), .A2(n4496), .ZN(n4495) );
  NOR2_X1 U5090 ( .A1(n7726), .A2(n4835), .ZN(n4499) );
  NAND2_X1 U5091 ( .A1(n4724), .A2(n4720), .ZN(n4722) );
  NAND2_X1 U5092 ( .A1(n7737), .A2(n7743), .ZN(n4720) );
  NAND2_X1 U5093 ( .A1(n6969), .A2(n9541), .ZN(n8466) );
  NOR2_X1 U5094 ( .A1(n9130), .A2(n9135), .ZN(n4491) );
  OAI21_X1 U5095 ( .B1(n4676), .B2(n5278), .A(n5189), .ZN(n4675) );
  INV_X1 U5096 ( .A(n4968), .ZN(n4737) );
  NOR2_X1 U5097 ( .A1(n4596), .A2(n4593), .ZN(n4592) );
  INV_X1 U5098 ( .A(n4594), .ZN(n4593) );
  INV_X1 U5099 ( .A(n4738), .ZN(n4596) );
  INV_X1 U5100 ( .A(SI_9_), .ZN(n10065) );
  AOI21_X1 U5101 ( .B1(n4850), .B2(n4848), .A(n4846), .ZN(n7767) );
  NOR2_X1 U5102 ( .A1(n4847), .A2(n4856), .ZN(n4846) );
  AND2_X1 U5103 ( .A1(n4854), .A2(n4849), .ZN(n4848) );
  INV_X1 U5104 ( .A(n4854), .ZN(n4847) );
  NOR2_X1 U5105 ( .A1(n6921), .A2(n7007), .ZN(n7014) );
  XNOR2_X1 U5106 ( .A(n4764), .B(n7289), .ZN(n4767) );
  NAND2_X1 U5107 ( .A1(n7318), .A2(n4536), .ZN(n7426) );
  NAND2_X1 U5108 ( .A1(n8009), .A2(n8010), .ZN(n8011) );
  NAND2_X1 U5109 ( .A1(n9667), .A2(n8013), .ZN(n8014) );
  OR2_X1 U5110 ( .A1(n9711), .A2(n8028), .ZN(n8031) );
  AND2_X1 U5111 ( .A1(n4371), .A2(n4420), .ZN(n4559) );
  AND2_X1 U5112 ( .A1(n4815), .A2(n5712), .ZN(n4814) );
  NAND2_X1 U5113 ( .A1(n4816), .A2(n7663), .ZN(n4815) );
  NAND2_X1 U5114 ( .A1(n5711), .A2(n5477), .ZN(n4799) );
  NAND2_X1 U5115 ( .A1(n4550), .A2(n6869), .ZN(n4809) );
  NAND2_X1 U5116 ( .A1(n9801), .A2(n5437), .ZN(n4550) );
  OR2_X1 U5117 ( .A1(n8261), .A2(n7904), .ZN(n7728) );
  AOI21_X1 U5118 ( .B1(n4839), .B2(n4843), .A(n7723), .ZN(n4837) );
  OR2_X1 U5119 ( .A1(n8298), .A2(n7893), .ZN(n7710) );
  NAND2_X1 U5120 ( .A1(n4547), .A2(n8200), .ZN(n4546) );
  NAND2_X1 U5121 ( .A1(n4466), .A2(n5356), .ZN(n5489) );
  AND2_X1 U5122 ( .A1(n6200), .A2(n6199), .ZN(n6202) );
  INV_X1 U5123 ( .A(n6229), .ZN(n4666) );
  INV_X1 U5124 ( .A(n6204), .ZN(n4668) );
  NAND2_X1 U5125 ( .A1(n6217), .A2(n6216), .ZN(n4669) );
  NAND2_X1 U5126 ( .A1(n4576), .A2(n4575), .ZN(n4574) );
  AOI21_X1 U5127 ( .B1(n8610), .B2(n8734), .A(n8573), .ZN(n4575) );
  OR2_X1 U5128 ( .A1(n9103), .A2(n8867), .ZN(n8624) );
  NAND2_X1 U5129 ( .A1(n4491), .A2(n8957), .ZN(n4490) );
  OR2_X1 U5130 ( .A1(n9125), .A2(n8964), .ZN(n8596) );
  INV_X1 U5131 ( .A(n4867), .ZN(n4866) );
  OAI21_X1 U5132 ( .B1(n4389), .B2(n4868), .A(n7837), .ZN(n4867) );
  OR2_X1 U5133 ( .A1(n9130), .A2(n8980), .ZN(n8558) );
  OR2_X1 U5134 ( .A1(n6098), .A2(n6097), .ZN(n6110) );
  INV_X1 U5135 ( .A(n6042), .ZN(n6040) );
  AND2_X1 U5136 ( .A1(n7163), .A2(n8478), .ZN(n4632) );
  NAND2_X1 U5137 ( .A1(n6970), .A2(n6978), .ZN(n8477) );
  INV_X1 U5138 ( .A(n8673), .ZN(n6907) );
  NAND2_X1 U5139 ( .A1(n9491), .A2(n6974), .ZN(n8468) );
  OR2_X1 U5140 ( .A1(n8890), .A2(n8898), .ZN(n8591) );
  NOR2_X1 U5141 ( .A1(n8989), .A2(n9135), .ZN(n8981) );
  NAND2_X1 U5142 ( .A1(n5252), .A2(n5251), .ZN(n5261) );
  OR2_X1 U5143 ( .A1(n5250), .A2(n5249), .ZN(n5251) );
  OR2_X1 U5144 ( .A1(n5248), .A2(n10043), .ZN(n5252) );
  XNOR2_X1 U5145 ( .A(n5250), .B(n5249), .ZN(n5248) );
  NOR2_X2 U5146 ( .A1(n5082), .A2(n4647), .ZN(n4646) );
  NAND2_X1 U5147 ( .A1(n4649), .A2(n4648), .ZN(n4647) );
  INV_X1 U5148 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n4649) );
  INV_X1 U5149 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n4648) );
  INV_X1 U5150 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n4888) );
  INV_X1 U5151 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n4887) );
  AOI21_X1 U5152 ( .B1(n4731), .B2(n4728), .A(n4408), .ZN(n4726) );
  NAND2_X1 U5153 ( .A1(n5119), .A2(n4454), .ZN(n4741) );
  OAI21_X1 U5154 ( .B1(n4967), .B2(SI_12_), .A(n4968), .ZN(n5126) );
  AND2_X1 U5155 ( .A1(n4740), .A2(n4965), .ZN(n4738) );
  INV_X1 U5156 ( .A(n5126), .ZN(n4740) );
  NAND2_X1 U5157 ( .A1(n4956), .A2(n10065), .ZN(n4959) );
  NOR2_X1 U5158 ( .A1(n5827), .A2(n7964), .ZN(n4904) );
  NAND2_X1 U5159 ( .A1(n6780), .A2(n4702), .ZN(n6939) );
  AND2_X1 U5160 ( .A1(n6375), .A2(n5865), .ZN(n7899) );
  INV_X1 U5161 ( .A(n7911), .ZN(n5822) );
  INV_X1 U5162 ( .A(n5798), .ZN(n4701) );
  AND2_X1 U5163 ( .A1(n6940), .A2(n5796), .ZN(n4702) );
  NAND2_X1 U5164 ( .A1(n4695), .A2(n7389), .ZN(n4694) );
  INV_X1 U5165 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n4696) );
  AND2_X1 U5166 ( .A1(n7817), .A2(n7808), .ZN(n7732) );
  AND2_X1 U5167 ( .A1(n5334), .A2(n7495), .ZN(n5335) );
  NAND2_X1 U5168 ( .A1(n4459), .A2(n4458), .ZN(n4457) );
  OR2_X1 U5169 ( .A1(n8046), .A2(n4460), .ZN(n4459) );
  NAND2_X1 U5170 ( .A1(n8046), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n4458) );
  AND2_X1 U5171 ( .A1(n6653), .A2(n6652), .ZN(n6741) );
  NAND2_X1 U5172 ( .A1(n4753), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n4752) );
  NAND2_X1 U5173 ( .A1(n6746), .A2(n6805), .ZN(n6813) );
  NOR2_X1 U5174 ( .A1(n6741), .A2(n4535), .ZN(n6799) );
  NOR2_X1 U5175 ( .A1(n6742), .A2(n6651), .ZN(n4535) );
  NOR2_X1 U5176 ( .A1(n6918), .A2(n4533), .ZN(n7000) );
  AND2_X1 U5177 ( .A1(n6920), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n4533) );
  AND2_X1 U5178 ( .A1(n4764), .A2(n7295), .ZN(n4769) );
  XNOR2_X1 U5179 ( .A(n7426), .B(n7418), .ZN(n7321) );
  NAND2_X1 U5180 ( .A1(n7430), .A2(n7431), .ZN(n8009) );
  XNOR2_X1 U5181 ( .A(n8011), .B(n8050), .ZN(n9650) );
  NOR2_X1 U5182 ( .A1(n8024), .A2(n9656), .ZN(n9677) );
  NOR2_X1 U5183 ( .A1(n9677), .A2(n9676), .ZN(n9675) );
  NAND2_X1 U5184 ( .A1(n9668), .A2(n9669), .ZN(n9667) );
  NAND2_X1 U5185 ( .A1(n9671), .A2(n9672), .ZN(n9670) );
  OR2_X1 U5186 ( .A1(n9675), .A2(n4760), .ZN(n4757) );
  NAND2_X1 U5187 ( .A1(n4763), .A2(n8042), .ZN(n4760) );
  NAND2_X1 U5188 ( .A1(n9675), .A2(n4759), .ZN(n4756) );
  XNOR2_X1 U5189 ( .A(n8014), .B(n8042), .ZN(n9686) );
  NAND2_X1 U5190 ( .A1(n9687), .A2(n8054), .ZN(n9707) );
  XNOR2_X1 U5191 ( .A(n8017), .B(n8039), .ZN(n9724) );
  OR2_X1 U5192 ( .A1(n5518), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5531) );
  NAND2_X1 U5193 ( .A1(n6990), .A2(n5710), .ZN(n4818) );
  NAND2_X1 U5194 ( .A1(n4818), .A2(n4816), .ZN(n7189) );
  NAND2_X1 U5195 ( .A1(n7192), .A2(n7783), .ZN(n7191) );
  INV_X1 U5196 ( .A(n4542), .ZN(n7192) );
  AOI21_X1 U5197 ( .B1(n7089), .B2(n5455), .A(n5454), .ZN(n6985) );
  NAND2_X1 U5198 ( .A1(n6545), .A2(n6598), .ZN(n7612) );
  AND2_X1 U5199 ( .A1(n5741), .A2(n5740), .ZN(n6602) );
  NAND2_X1 U5200 ( .A1(n4798), .A2(n5649), .ZN(n8093) );
  AOI21_X1 U5201 ( .B1(n8116), .B2(n7730), .A(n5719), .ZN(n8099) );
  AOI21_X1 U5202 ( .B1(n8148), .B2(n4780), .A(n4778), .ZN(n4777) );
  NAND2_X1 U5203 ( .A1(n4779), .A2(n5636), .ZN(n4778) );
  NAND2_X1 U5204 ( .A1(n4780), .A2(n4783), .ZN(n4779) );
  AND2_X1 U5205 ( .A1(n7729), .A2(n7730), .ZN(n8117) );
  AND2_X1 U5206 ( .A1(n4841), .A2(n7770), .ZN(n4839) );
  AOI21_X1 U5207 ( .B1(n4842), .B2(n4845), .A(n7718), .ZN(n4841) );
  NAND2_X1 U5208 ( .A1(n8155), .A2(n4842), .ZN(n4840) );
  INV_X1 U5209 ( .A(n7716), .ZN(n4845) );
  NAND2_X1 U5210 ( .A1(n7793), .A2(n4804), .ZN(n4803) );
  INV_X1 U5211 ( .A(n7506), .ZN(n4804) );
  NAND2_X1 U5212 ( .A1(n4821), .A2(n4825), .ZN(n4820) );
  AND2_X1 U5213 ( .A1(n4823), .A2(n7610), .ZN(n4821) );
  OR2_X1 U5214 ( .A1(n5885), .A2(n7747), .ZN(n9760) );
  NAND2_X1 U5215 ( .A1(n4824), .A2(n7695), .ZN(n4823) );
  INV_X1 U5216 ( .A(n4827), .ZN(n4824) );
  AOI21_X1 U5217 ( .B1(n4830), .B2(n4829), .A(n4828), .ZN(n4827) );
  INV_X1 U5218 ( .A(n7694), .ZN(n4828) );
  NAND2_X1 U5219 ( .A1(n4830), .A2(n7695), .ZN(n4825) );
  NAND2_X1 U5220 ( .A1(n4538), .A2(n4907), .ZN(n7544) );
  OR2_X1 U5221 ( .A1(n7478), .A2(n7376), .ZN(n4907) );
  NAND2_X1 U5222 ( .A1(n7441), .A2(n5524), .ZN(n4538) );
  OR2_X1 U5223 ( .A1(n7872), .A2(n7996), .ZN(n5524) );
  NOR2_X1 U5224 ( .A1(n5716), .A2(n7686), .ZN(n4831) );
  AND2_X1 U5225 ( .A1(n7695), .A2(n7694), .ZN(n7692) );
  INV_X1 U5226 ( .A(n9762), .ZN(n9744) );
  INV_X1 U5227 ( .A(n9760), .ZN(n9746) );
  INV_X1 U5228 ( .A(n7685), .ZN(n4832) );
  NAND2_X1 U5229 ( .A1(n5492), .A2(n5491), .ZN(n9834) );
  NAND2_X1 U5230 ( .A1(n5692), .A2(n5691), .ZN(n9765) );
  AND2_X1 U5231 ( .A1(n5734), .A2(n4422), .ZN(n5331) );
  AND2_X1 U5232 ( .A1(n5324), .A2(n4861), .ZN(n4860) );
  INV_X1 U5233 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n5324) );
  INV_X1 U5234 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n4861) );
  NOR2_X1 U5235 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n5322) );
  OR2_X1 U5236 ( .A1(n5330), .A2(n5385), .ZN(n5386) );
  AOI21_X1 U5237 ( .B1(n4373), .B2(n4660), .A(n4405), .ZN(n4656) );
  OR2_X1 U5238 ( .A1(n6174), .A2(n6173), .ZN(n6176) );
  OR2_X1 U5239 ( .A1(n6027), .A2(n6026), .ZN(n6042) );
  AOI21_X1 U5240 ( .B1(n8756), .B2(n6323), .A(n5915), .ZN(n5920) );
  NAND2_X1 U5241 ( .A1(n4688), .A2(n6262), .ZN(n4683) );
  INV_X1 U5242 ( .A(n6248), .ZN(n6246) );
  AND2_X1 U5243 ( .A1(n6486), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6406) );
  NAND2_X1 U5244 ( .A1(n9312), .A2(n8821), .ZN(n4604) );
  NAND2_X1 U5245 ( .A1(n4602), .A2(n4601), .ZN(n4600) );
  INV_X1 U5246 ( .A(n9324), .ZN(n4601) );
  NOR2_X1 U5247 ( .A1(n9248), .A2(n4438), .ZN(n9264) );
  NAND2_X1 U5248 ( .A1(n8910), .A2(n8878), .ZN(n4884) );
  NAND2_X1 U5249 ( .A1(n8930), .A2(n4479), .ZN(n4484) );
  INV_X1 U5250 ( .A(n4481), .ZN(n4479) );
  AND2_X1 U5251 ( .A1(n8624), .A2(n8864), .ZN(n8900) );
  AND2_X1 U5252 ( .A1(n6297), .A2(n6296), .ZN(n8897) );
  INV_X1 U5253 ( .A(n8938), .ZN(n8950) );
  NOR2_X1 U5254 ( .A1(n8976), .A2(n7847), .ZN(n8962) );
  NAND2_X1 U5255 ( .A1(n4375), .A2(n4394), .ZN(n4869) );
  NAND2_X1 U5256 ( .A1(n9045), .A2(n7845), .ZN(n9028) );
  NAND2_X1 U5257 ( .A1(n8537), .A2(n4433), .ZN(n4634) );
  NAND2_X1 U5258 ( .A1(n4635), .A2(n4433), .ZN(n4633) );
  OAI21_X1 U5259 ( .B1(n7845), .B2(n4636), .A(n8996), .ZN(n4635) );
  NAND2_X1 U5260 ( .A1(n4392), .A2(n4882), .ZN(n4881) );
  OR2_X1 U5261 ( .A1(n4418), .A2(n4911), .ZN(n4882) );
  INV_X1 U5262 ( .A(n9039), .ZN(n4883) );
  NOR2_X1 U5263 ( .A1(n9078), .A2(n7829), .ZN(n5182) );
  NOR2_X1 U5264 ( .A1(n9078), .A2(n4485), .ZN(n9040) );
  INV_X1 U5265 ( .A(n4487), .ZN(n4485) );
  AND4_X1 U5266 ( .A1(n6127), .A2(n6126), .A3(n6125), .A4(n6124), .ZN(n9061)
         );
  NAND2_X1 U5267 ( .A1(n9074), .A2(n9075), .ZN(n4625) );
  AND2_X1 U5268 ( .A1(n8528), .A2(n8465), .ZN(n9075) );
  AND2_X1 U5269 ( .A1(n8338), .A2(n8519), .ZN(n7563) );
  AOI21_X1 U5270 ( .B1(n4874), .B2(n4365), .A(n4381), .ZN(n4873) );
  INV_X1 U5271 ( .A(n8635), .ZN(n4874) );
  NOR2_X1 U5272 ( .A1(n8635), .A2(n4628), .ZN(n4875) );
  NAND2_X1 U5273 ( .A1(n8681), .A2(n4627), .ZN(n8683) );
  NAND2_X1 U5274 ( .A1(n7261), .A2(n4631), .ZN(n4627) );
  AND2_X1 U5275 ( .A1(n8471), .A2(n8474), .ZN(n4631) );
  AND2_X1 U5276 ( .A1(n8506), .A2(n8501), .ZN(n7273) );
  NAND2_X1 U5277 ( .A1(n7163), .A2(n8471), .ZN(n9475) );
  AND2_X1 U5278 ( .A1(n5286), .A2(n8622), .ZN(n9490) );
  OR2_X1 U5279 ( .A1(n5267), .A2(n6433), .ZN(n5045) );
  INV_X1 U5280 ( .A(n9490), .ZN(n9060) );
  AND2_X1 U5281 ( .A1(n8591), .A2(n8618), .ZN(n8882) );
  NAND2_X1 U5282 ( .A1(n8886), .A2(n4483), .ZN(n9098) );
  NAND2_X1 U5283 ( .A1(n4484), .A2(n8890), .ZN(n4483) );
  INV_X1 U5284 ( .A(n8957), .ZN(n9125) );
  AND2_X1 U5285 ( .A1(n5166), .A2(n5165), .ZN(n9295) );
  OR2_X1 U5286 ( .A1(n9513), .A2(n8730), .ZN(n9568) );
  AND2_X1 U5287 ( .A1(n8734), .A2(n6854), .ZN(n9565) );
  INV_X1 U5288 ( .A(n6897), .ZN(n7030) );
  XNOR2_X1 U5289 ( .A(n5248), .B(SI_29_), .ZN(n5673) );
  XNOR2_X1 U5290 ( .A(n5291), .B(P1_IR_REG_26__SCAN_IN), .ZN(n5304) );
  INV_X1 U5291 ( .A(n4713), .ZN(n5233) );
  AOI21_X1 U5292 ( .B1(n4718), .B2(n4716), .A(n4434), .ZN(n4713) );
  XNOR2_X1 U5293 ( .A(n5229), .B(n5228), .ZN(n7117) );
  AND2_X1 U5294 ( .A1(n4718), .A2(n4719), .ZN(n5229) );
  XNOR2_X1 U5295 ( .A(n5297), .B(P1_IR_REG_22__SCAN_IN), .ZN(n8589) );
  NAND2_X1 U5296 ( .A1(n5184), .A2(n4991), .ZN(n5207) );
  XNOR2_X1 U5297 ( .A(n5199), .B(n5198), .ZN(n6848) );
  XNOR2_X1 U5298 ( .A(n5173), .B(n5172), .ZN(n6720) );
  NAND2_X1 U5299 ( .A1(n4591), .A2(n4590), .ZN(n5144) );
  XNOR2_X1 U5300 ( .A(n4944), .B(n4943), .ZN(n5077) );
  NAND2_X1 U5301 ( .A1(n4733), .A2(n4938), .ZN(n4941) );
  INV_X1 U5302 ( .A(n5070), .ZN(n4733) );
  NAND2_X1 U5303 ( .A1(n5875), .A2(n5874), .ZN(n5879) );
  AOI21_X1 U5304 ( .B1(n7897), .B2(n5873), .A(n5872), .ZN(n5875) );
  AND4_X1 U5305 ( .A1(n5537), .A2(n5536), .A3(n5535), .A4(n5534), .ZN(n7912)
         );
  AND4_X1 U5306 ( .A1(n5476), .A2(n5475), .A3(n5474), .A4(n5473), .ZN(n7282)
         );
  AOI21_X1 U5307 ( .B1(n6585), .B2(n6584), .A(n5783), .ZN(n6620) );
  AND4_X1 U5308 ( .A1(n5561), .A2(n5560), .A3(n5559), .A4(n5558), .ZN(n7885)
         );
  NAND2_X1 U5309 ( .A1(n5870), .A2(n5869), .ZN(n6402) );
  AND4_X1 U5310 ( .A1(n5365), .A2(n5364), .A3(n5363), .A4(n5362), .ZN(n7451)
         );
  AND2_X1 U5311 ( .A1(n5625), .A2(n5624), .ZN(n7903) );
  NAND2_X1 U5312 ( .A1(n7980), .A2(n5821), .ZN(n7910) );
  NAND2_X1 U5313 ( .A1(n6620), .A2(n6619), .ZN(n6618) );
  AND4_X1 U5314 ( .A1(n5462), .A2(n5461), .A3(n5460), .A4(n5459), .ZN(n7090)
         );
  AND3_X1 U5315 ( .A1(n5572), .A2(n5571), .A3(n5570), .ZN(n7947) );
  NAND2_X1 U5316 ( .A1(n5505), .A2(n5504), .ZN(n9286) );
  AND3_X1 U5317 ( .A1(n5594), .A2(n5593), .A3(n5592), .ZN(n7957) );
  AND4_X1 U5318 ( .A1(n5551), .A2(n5550), .A3(n5549), .A4(n5548), .ZN(n7994)
         );
  INV_X1 U5319 ( .A(n8003), .ZN(n5437) );
  AOI21_X1 U5320 ( .B1(n4517), .B2(n4516), .A(n4515), .ZN(n7813) );
  AOI21_X1 U5321 ( .B1(n7750), .B2(n7749), .A(n4379), .ZN(n4517) );
  OR2_X1 U5322 ( .A1(n7812), .A2(n4423), .ZN(n4515) );
  NAND2_X1 U5323 ( .A1(n7748), .A2(n7732), .ZN(n4516) );
  NAND2_X1 U5324 ( .A1(n5658), .A2(n5657), .ZN(n8102) );
  INV_X1 U5325 ( .A(n7903), .ZN(n8138) );
  NOR2_X1 U5326 ( .A1(n6409), .A2(n6515), .ZN(n6522) );
  OR2_X1 U5327 ( .A1(n6525), .A2(n6526), .ZN(n4456) );
  NOR2_X1 U5328 ( .A1(n6522), .A2(n4461), .ZN(n6525) );
  NOR2_X1 U5329 ( .A1(n4462), .A2(n6421), .ZN(n4461) );
  INV_X1 U5330 ( .A(n6524), .ZN(n4462) );
  XNOR2_X1 U5331 ( .A(n4457), .B(n6562), .ZN(n6526) );
  XNOR2_X1 U5332 ( .A(n6799), .B(n6805), .ZN(n6801) );
  XNOR2_X1 U5333 ( .A(n7000), .B(n4532), .ZN(n7002) );
  NAND2_X1 U5334 ( .A1(n6916), .A2(n4436), .ZN(n7009) );
  NOR2_X1 U5335 ( .A1(n7003), .A2(n7004), .ZN(n7121) );
  OAI21_X1 U5336 ( .B1(n8067), .B2(n8066), .A(n4470), .ZN(n4469) );
  NOR2_X1 U5337 ( .A1(n4471), .A2(n8065), .ZN(n4470) );
  XNOR2_X1 U5338 ( .A(n8035), .B(n8038), .ZN(n4774) );
  INV_X1 U5339 ( .A(n8208), .ZN(n9753) );
  NAND2_X1 U5340 ( .A1(n5651), .A2(n5650), .ZN(n8257) );
  NAND2_X1 U5341 ( .A1(n5427), .A2(n4806), .ZN(n6863) );
  NOR2_X1 U5342 ( .A1(n4398), .A2(n4807), .ZN(n4806) );
  NOR2_X1 U5343 ( .A1(n5379), .A2(n6920), .ZN(n4807) );
  OR2_X1 U5344 ( .A1(n7861), .A2(n9796), .ZN(n5725) );
  NOR2_X1 U5345 ( .A1(n9836), .A2(n8256), .ZN(n4552) );
  AOI21_X1 U5346 ( .B1(n4557), .B2(n9765), .A(n4554), .ZN(n8255) );
  NAND2_X1 U5347 ( .A1(n4556), .A2(n4555), .ZN(n4554) );
  XNOR2_X1 U5348 ( .A(n8093), .B(n8092), .ZN(n4557) );
  NAND2_X1 U5349 ( .A1(n8111), .A2(n9744), .ZN(n4555) );
  NAND2_X1 U5350 ( .A1(n5607), .A2(n5606), .ZN(n8280) );
  INV_X1 U5351 ( .A(n8753), .ZN(n7164) );
  NAND2_X1 U5352 ( .A1(n8445), .A2(n7598), .ZN(n7600) );
  NAND2_X1 U5353 ( .A1(n5243), .A2(n5242), .ZN(n9109) );
  NOR2_X1 U5354 ( .A1(n8407), .A2(n6897), .ZN(n6729) );
  NAND2_X1 U5355 ( .A1(n5195), .A2(n5194), .ZN(n9154) );
  AND4_X1 U5356 ( .A1(n6015), .A2(n6014), .A3(n6013), .A4(n6012), .ZN(n8483)
         );
  INV_X1 U5357 ( .A(n8462), .ZN(n8444) );
  INV_X1 U5358 ( .A(n8934), .ZN(n9114) );
  INV_X1 U5359 ( .A(n7471), .ZN(n8751) );
  AND2_X1 U5360 ( .A1(n5067), .A2(n5074), .ZN(n9318) );
  NAND2_X1 U5361 ( .A1(n4673), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5190) );
  NAND2_X1 U5362 ( .A1(n4358), .A2(n4676), .ZN(n4673) );
  NOR2_X1 U5363 ( .A1(n9426), .A2(n4598), .ZN(n9440) );
  AND2_X1 U5364 ( .A1(n9435), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n4598) );
  OR2_X1 U5365 ( .A1(n9453), .A2(n9452), .ZN(n9462) );
  NAND2_X1 U5366 ( .A1(n8845), .A2(n4613), .ZN(n4612) );
  INV_X1 U5367 ( .A(n4614), .ZN(n4613) );
  OAI21_X1 U5368 ( .B1(n8846), .B2(n9413), .A(n9460), .ZN(n4614) );
  NAND2_X1 U5369 ( .A1(n8923), .A2(n8922), .ZN(n8924) );
  INV_X1 U5370 ( .A(n9109), .ZN(n8916) );
  AND2_X1 U5371 ( .A1(n5093), .A2(n4424), .ZN(n4477) );
  INV_X1 U5372 ( .A(n9472), .ZN(n9067) );
  OR2_X1 U5373 ( .A1(n8660), .A2(n6343), .ZN(n9499) );
  OAI211_X1 U5374 ( .C1(n6897), .C2(n7029), .A(n9496), .B(n9494), .ZN(n9521)
         );
  NAND2_X1 U5375 ( .A1(n8854), .A2(n5290), .ZN(n9091) );
  OAI21_X1 U5376 ( .B1(n8851), .B2(n9613), .A(n9093), .ZN(n5289) );
  INV_X1 U5377 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n4645) );
  NAND2_X1 U5378 ( .A1(n4641), .A2(n4386), .ZN(n4639) );
  INV_X1 U5379 ( .A(n4642), .ZN(n4641) );
  INV_X1 U5380 ( .A(n8735), .ZN(n8738) );
  CLKBUF_X1 U5381 ( .A(n9503), .Z(n4453) );
  INV_X1 U5382 ( .A(n7617), .ZN(n4519) );
  NAND2_X1 U5383 ( .A1(n7611), .A2(n7808), .ZN(n7616) );
  NAND2_X1 U5384 ( .A1(n4513), .A2(n4514), .ZN(n4507) );
  NAND2_X1 U5385 ( .A1(n7696), .A2(n7697), .ZN(n4514) );
  AOI21_X1 U5386 ( .B1(n8539), .B2(n8514), .A(n8538), .ZN(n8546) );
  NAND2_X1 U5387 ( .A1(n4509), .A2(n7693), .ZN(n4508) );
  AND2_X1 U5388 ( .A1(n4513), .A2(n4425), .ZN(n4509) );
  AND2_X1 U5389 ( .A1(n4507), .A2(n4510), .ZN(n4506) );
  NOR2_X1 U5390 ( .A1(n4512), .A2(n4511), .ZN(n4510) );
  INV_X1 U5391 ( .A(n7701), .ZN(n4511) );
  OAI21_X1 U5392 ( .B1(n8553), .B2(n4566), .A(n4564), .ZN(n4563) );
  INV_X1 U5393 ( .A(n8555), .ZN(n4566) );
  NAND2_X1 U5394 ( .A1(n6898), .A2(n6897), .ZN(n8668) );
  NAND2_X1 U5395 ( .A1(n7708), .A2(n4527), .ZN(n4526) );
  NOR2_X1 U5396 ( .A1(n4528), .A2(n7747), .ZN(n4527) );
  INV_X1 U5397 ( .A(n7714), .ZN(n4528) );
  INV_X1 U5398 ( .A(n8145), .ZN(n4523) );
  INV_X1 U5399 ( .A(n7731), .ZN(n4497) );
  INV_X1 U5400 ( .A(n8101), .ZN(n4496) );
  INV_X1 U5401 ( .A(n8526), .ZN(n4561) );
  INV_X1 U5402 ( .A(n8527), .ZN(n4562) );
  INV_X1 U5403 ( .A(n5171), .ZN(n4972) );
  NAND2_X1 U5404 ( .A1(n4855), .A2(n9279), .ZN(n4854) );
  AND2_X1 U5405 ( .A1(n7764), .A2(n7763), .ZN(n4856) );
  AND2_X1 U5406 ( .A1(n5439), .A2(n9940), .ZN(n5456) );
  NOR2_X1 U5407 ( .A1(n5440), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5439) );
  NAND2_X1 U5408 ( .A1(n4580), .A2(n8734), .ZN(n4579) );
  OR2_X1 U5409 ( .A1(n8570), .A2(n8734), .ZN(n4581) );
  INV_X1 U5410 ( .A(n8610), .ZN(n4577) );
  NAND2_X1 U5411 ( .A1(n7261), .A2(n8474), .ZN(n8631) );
  NAND2_X1 U5412 ( .A1(n5022), .A2(n5021), .ZN(n5250) );
  NOR2_X1 U5413 ( .A1(n4712), .A2(n4434), .ZN(n4711) );
  INV_X1 U5414 ( .A(n5004), .ZN(n4712) );
  INV_X1 U5415 ( .A(n4715), .ZN(n4714) );
  OAI21_X1 U5416 ( .B1(n4716), .B2(n4434), .A(n5232), .ZN(n4715) );
  AND2_X1 U5417 ( .A1(n5222), .A2(n5000), .ZN(n5004) );
  OR2_X1 U5418 ( .A1(n4728), .A2(n4992), .ZN(n4727) );
  AND2_X1 U5419 ( .A1(n4991), .A2(SI_20_), .ZN(n4992) );
  AOI21_X1 U5420 ( .B1(n4990), .B2(n4730), .A(n4729), .ZN(n4728) );
  INV_X1 U5421 ( .A(n5208), .ZN(n4729) );
  INV_X1 U5422 ( .A(n4991), .ZN(n4730) );
  INV_X1 U5423 ( .A(n4990), .ZN(n4731) );
  OR2_X1 U5424 ( .A1(n5167), .A2(n4975), .ZN(n4971) );
  AND2_X1 U5425 ( .A1(n4972), .A2(n10069), .ZN(n4975) );
  INV_X1 U5426 ( .A(n5142), .ZN(n4969) );
  NOR2_X1 U5427 ( .A1(n4961), .A2(n4595), .ZN(n4594) );
  INV_X1 U5428 ( .A(n4959), .ZN(n4595) );
  INV_X1 U5429 ( .A(n5109), .ZN(n4961) );
  NAND2_X1 U5430 ( .A1(n4473), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n4920) );
  INV_X1 U5431 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4473) );
  NAND2_X1 U5432 ( .A1(n4475), .A2(n4474), .ZN(n4919) );
  INV_X1 U5433 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n4475) );
  INV_X1 U5434 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4474) );
  NOR2_X1 U5435 ( .A1(n7800), .A2(n7735), .ZN(n4723) );
  NAND2_X1 U5436 ( .A1(n4494), .A2(n7736), .ZN(n4493) );
  NAND2_X1 U5437 ( .A1(n6558), .A2(n6559), .ZN(n6648) );
  AND3_X1 U5438 ( .A1(n4748), .A2(n8021), .A3(n4747), .ZN(n8023) );
  NAND2_X1 U5439 ( .A1(n9703), .A2(n4534), .ZN(n8017) );
  OR2_X1 U5440 ( .A1(n8040), .A2(n8016), .ZN(n4534) );
  NAND2_X1 U5441 ( .A1(n9725), .A2(n4446), .ZN(n8058) );
  NOR2_X1 U5442 ( .A1(n5619), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n5628) );
  AND2_X1 U5443 ( .A1(n5579), .A2(n10021), .ZN(n5589) );
  AND2_X1 U5444 ( .A1(n5338), .A2(n10066), .ZN(n5545) );
  NOR2_X1 U5445 ( .A1(n5531), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5338) );
  NAND2_X1 U5446 ( .A1(n5456), .A2(n5336), .ZN(n5482) );
  INV_X1 U5447 ( .A(n6790), .ZN(n7773) );
  NAND2_X1 U5448 ( .A1(n8006), .A2(n6614), .ZN(n7611) );
  INV_X1 U5449 ( .A(n4913), .ZN(n4785) );
  INV_X1 U5450 ( .A(n4831), .ZN(n4829) );
  NOR2_X1 U5451 ( .A1(P2_IR_REG_26__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), .ZN(
        n4862) );
  INV_X1 U5452 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5756) );
  NAND2_X1 U5453 ( .A1(n4859), .A2(n4371), .ZN(n5726) );
  NOR2_X1 U5454 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n5320) );
  NOR2_X1 U5455 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), .ZN(
        n5321) );
  OR2_X1 U5456 ( .A1(n5411), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n5422) );
  INV_X1 U5457 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n4708) );
  INV_X1 U5458 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n5318) );
  NOR2_X1 U5459 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5385) );
  OR2_X1 U5460 ( .A1(n7460), .A2(n4660), .ZN(n4659) );
  INV_X1 U5461 ( .A(n6096), .ZN(n4660) );
  INV_X1 U5462 ( .A(n8442), .ZN(n4687) );
  INV_X1 U5463 ( .A(n8441), .ZN(n4686) );
  AND2_X1 U5464 ( .A1(n6240), .A2(n6239), .ZN(n6242) );
  NOR2_X1 U5465 ( .A1(n4655), .A2(n4654), .ZN(n4653) );
  INV_X1 U5466 ( .A(n6110), .ZN(n6108) );
  OR2_X1 U5467 ( .A1(n9109), .A2(n8897), .ZN(n8706) );
  NAND2_X1 U5468 ( .A1(n4482), .A2(n8916), .ZN(n4481) );
  OR2_X1 U5469 ( .A1(n9114), .A2(n8876), .ZN(n8625) );
  INV_X1 U5470 ( .A(n4869), .ZN(n4868) );
  INV_X1 U5471 ( .A(n7833), .ZN(n4880) );
  NOR2_X1 U5472 ( .A1(n9154), .A2(n7829), .ZN(n4487) );
  OR2_X1 U5473 ( .A1(n7823), .A2(n8384), .ZN(n7843) );
  OR2_X1 U5474 ( .A1(n6086), .A2(n6085), .ZN(n6098) );
  NOR2_X1 U5475 ( .A1(n7268), .A2(n7475), .ZN(n7269) );
  NAND2_X1 U5476 ( .A1(n6054), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n6086) );
  INV_X1 U5477 ( .A(n6069), .ZN(n6054) );
  NAND2_X1 U5478 ( .A1(n7068), .A2(n9548), .ZN(n8678) );
  NAND2_X1 U5479 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n5978) );
  NOR2_X1 U5480 ( .A1(n8989), .A2(n4489), .ZN(n8965) );
  INV_X1 U5481 ( .A(n4491), .ZN(n4489) );
  OR2_X1 U5482 ( .A1(n7239), .A2(n7343), .ZN(n7268) );
  NOR2_X1 U5483 ( .A1(n4899), .A2(n4717), .ZN(n4716) );
  INV_X1 U5484 ( .A(n5228), .ZN(n4717) );
  AND2_X1 U5485 ( .A1(n5196), .A2(n4987), .ZN(n4988) );
  AND2_X1 U5486 ( .A1(n5183), .A2(n4985), .ZN(n4991) );
  NAND2_X1 U5487 ( .A1(n4672), .A2(n4671), .ZN(n5192) );
  AOI21_X1 U5488 ( .B1(n4674), .B2(n5278), .A(n5278), .ZN(n4671) );
  INV_X1 U5489 ( .A(n4675), .ZN(n4674) );
  NOR2_X1 U5490 ( .A1(n5167), .A2(n4588), .ZN(n4587) );
  INV_X1 U5491 ( .A(n4970), .ZN(n4588) );
  NAND2_X1 U5492 ( .A1(n4739), .A2(n5133), .ZN(n4590) );
  NAND2_X1 U5493 ( .A1(n4735), .A2(n4396), .ZN(n4739) );
  XNOR2_X1 U5494 ( .A(n4962), .B(n10040), .ZN(n5109) );
  OAI21_X1 U5495 ( .B1(n5099), .B2(n4742), .A(n4955), .ZN(n5102) );
  INV_X1 U5496 ( .A(n4414), .ZN(n4742) );
  AND2_X1 U5497 ( .A1(n4959), .A2(n4958), .ZN(n4910) );
  NAND2_X1 U5498 ( .A1(n4952), .A2(n10092), .ZN(n4955) );
  NAND2_X1 U5499 ( .A1(n4390), .A2(n5092), .ZN(n4572) );
  AND2_X1 U5500 ( .A1(n4732), .A2(n5092), .ZN(n4567) );
  OAI21_X1 U5501 ( .B1(n6431), .B2(n4931), .A(n4930), .ZN(n4932) );
  AND2_X1 U5502 ( .A1(n7898), .A2(n5853), .ZN(n7933) );
  AND2_X1 U5503 ( .A1(n5694), .A2(n5379), .ZN(n5885) );
  OR2_X1 U5504 ( .A1(n5428), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5440) );
  OR2_X1 U5505 ( .A1(n5867), .A2(n5866), .ZN(n6379) );
  AND2_X1 U5506 ( .A1(n7761), .A2(n7760), .ZN(n8069) );
  AND2_X1 U5507 ( .A1(n5604), .A2(n5603), .ZN(n5844) );
  OAI21_X1 U5508 ( .B1(n6535), .B2(P2_REG1_REG_2__SCAN_IN), .A(n4529), .ZN(
        n6533) );
  NAND2_X1 U5509 ( .A1(n6535), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n4529) );
  NAND2_X1 U5510 ( .A1(n6533), .A2(n6532), .ZN(n6559) );
  XNOR2_X1 U5511 ( .A(n6648), .B(n6560), .ZN(n6646) );
  AND2_X1 U5512 ( .A1(n4914), .A2(n6642), .ZN(n6566) );
  NAND2_X1 U5513 ( .A1(n6566), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n6644) );
  NOR2_X1 U5514 ( .A1(n6804), .A2(n4464), .ZN(n6808) );
  NOR2_X1 U5515 ( .A1(n4465), .A2(n6753), .ZN(n4464) );
  INV_X1 U5516 ( .A(n6806), .ZN(n4465) );
  NAND2_X1 U5517 ( .A1(n4755), .A2(n4447), .ZN(n6815) );
  AND2_X1 U5518 ( .A1(n6921), .A2(n7007), .ZN(n6922) );
  AOI21_X1 U5519 ( .B1(n7009), .B2(n7008), .A(n4463), .ZN(n7125) );
  AND2_X1 U5520 ( .A1(n7006), .A2(n7007), .ZN(n4463) );
  AOI21_X1 U5521 ( .B1(n7018), .B2(n7016), .A(n7017), .ZN(n7136) );
  NAND2_X1 U5522 ( .A1(n6924), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n7018) );
  INV_X1 U5523 ( .A(n8057), .ZN(n6419) );
  OR2_X1 U5524 ( .A1(n5450), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n5467) );
  INV_X1 U5525 ( .A(n4767), .ZN(n7138) );
  INV_X1 U5526 ( .A(n4769), .ZN(n4768) );
  NOR2_X1 U5527 ( .A1(n7297), .A2(n7198), .ZN(n4766) );
  NOR2_X1 U5528 ( .A1(n7138), .A2(n7198), .ZN(n7294) );
  NAND2_X1 U5529 ( .A1(n7428), .A2(n7429), .ZN(n7430) );
  OR2_X1 U5530 ( .A1(n7326), .A2(n4749), .ZN(n4747) );
  NAND2_X1 U5531 ( .A1(n4750), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n4749) );
  INV_X1 U5532 ( .A(n7414), .ZN(n4750) );
  OR2_X1 U5533 ( .A1(n4387), .A2(n7414), .ZN(n4748) );
  OR2_X1 U5534 ( .A1(n7326), .A2(n7327), .ZN(n4751) );
  NAND2_X1 U5535 ( .A1(n9649), .A2(n8012), .ZN(n9668) );
  NAND2_X1 U5536 ( .A1(n4761), .A2(n4759), .ZN(n4758) );
  NAND2_X1 U5537 ( .A1(n9670), .A2(n8053), .ZN(n9688) );
  NAND2_X1 U5538 ( .A1(n9688), .A2(n9689), .ZN(n9687) );
  NAND2_X1 U5539 ( .A1(n9685), .A2(n8015), .ZN(n9704) );
  NAND2_X1 U5540 ( .A1(n9704), .A2(n9705), .ZN(n9703) );
  AND2_X1 U5541 ( .A1(n4762), .A2(n4391), .ZN(n9713) );
  NAND2_X1 U5542 ( .A1(n9706), .A2(n8055), .ZN(n9726) );
  NAND2_X1 U5543 ( .A1(n9726), .A2(n9727), .ZN(n9725) );
  NAND2_X1 U5544 ( .A1(n8058), .A2(n8059), .ZN(n9203) );
  AND2_X1 U5545 ( .A1(n4559), .A2(n5327), .ZN(n4558) );
  INV_X1 U5546 ( .A(n4773), .ZN(n4471) );
  AOI21_X1 U5547 ( .B1(n9200), .B2(P2_ADDR_REG_19__SCAN_IN), .A(n4449), .ZN(
        n4773) );
  OAI21_X1 U5548 ( .B1(n9734), .B2(n4771), .A(n4770), .ZN(n9211) );
  NAND2_X1 U5549 ( .A1(n4772), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n4771) );
  INV_X1 U5550 ( .A(n9212), .ZN(n4772) );
  INV_X1 U5551 ( .A(n4853), .ZN(n4852) );
  OAI21_X1 U5552 ( .B1(n8077), .B2(n4857), .A(n4404), .ZN(n4853) );
  NOR2_X1 U5553 ( .A1(n8077), .A2(n8092), .ZN(n4851) );
  NAND2_X1 U5554 ( .A1(n7762), .A2(n7740), .ZN(n7800) );
  NAND2_X1 U5555 ( .A1(n4796), .A2(n8077), .ZN(n4792) );
  AOI21_X1 U5556 ( .B1(n8077), .B2(n4790), .A(n5672), .ZN(n4789) );
  INV_X1 U5557 ( .A(n4793), .ZN(n4790) );
  OR2_X1 U5558 ( .A1(n5608), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5619) );
  NAND2_X1 U5559 ( .A1(n5589), .A2(n10019), .ZN(n5597) );
  OR2_X1 U5560 ( .A1(n5556), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5568) );
  NAND2_X1 U5561 ( .A1(n5493), .A2(n5337), .ZN(n5518) );
  AND4_X1 U5562 ( .A1(n5523), .A2(n5522), .A3(n5521), .A4(n5520), .ZN(n7376)
         );
  OR2_X1 U5563 ( .A1(n5482), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5484) );
  AOI21_X1 U5564 ( .B1(n4814), .B2(n4817), .A(n4812), .ZN(n4811) );
  INV_X1 U5565 ( .A(n7671), .ZN(n4812) );
  NAND2_X1 U5566 ( .A1(n4541), .A2(n4540), .ZN(n7219) );
  NAND2_X1 U5567 ( .A1(n4416), .A2(n4364), .ZN(n4540) );
  NAND2_X1 U5568 ( .A1(n4542), .A2(n4378), .ZN(n4541) );
  AND2_X1 U5569 ( .A1(n7673), .A2(n7672), .ZN(n7782) );
  OR2_X1 U5570 ( .A1(n9823), .A2(n7282), .ZN(n7649) );
  AND2_X1 U5571 ( .A1(n7653), .A2(n6991), .ZN(n7779) );
  NAND2_X1 U5572 ( .A1(n5436), .A2(n4809), .ZN(n4808) );
  INV_X1 U5573 ( .A(n4809), .ZN(n6836) );
  AND2_X1 U5574 ( .A1(n6841), .A2(n7639), .ZN(n7775) );
  NAND2_X1 U5575 ( .A1(n9758), .A2(n9759), .ZN(n9757) );
  INV_X1 U5576 ( .A(n7612), .ZN(n5703) );
  OR2_X1 U5577 ( .A1(n8069), .A2(n8068), .ZN(n9280) );
  NAND2_X1 U5578 ( .A1(n4788), .A2(n4793), .ZN(n8079) );
  NAND2_X1 U5579 ( .A1(n8094), .A2(n9746), .ZN(n4556) );
  AND2_X1 U5580 ( .A1(n7728), .A2(n7727), .ZN(n8101) );
  NAND2_X1 U5581 ( .A1(n4836), .A2(n4834), .ZN(n8116) );
  AOI21_X1 U5582 ( .B1(n4837), .B2(n4838), .A(n4835), .ZN(n4834) );
  INV_X1 U5583 ( .A(n4839), .ZN(n4838) );
  INV_X1 U5584 ( .A(n7797), .ZN(n8158) );
  NAND2_X1 U5585 ( .A1(n8170), .A2(n8169), .ZN(n8168) );
  INV_X1 U5586 ( .A(n4545), .ZN(n4544) );
  OAI22_X1 U5587 ( .A1(n4546), .A2(n5563), .B1(n8203), .B2(n8310), .ZN(n4545)
         );
  OAI21_X1 U5588 ( .B1(n7374), .B2(n5512), .A(n7372), .ZN(n7441) );
  INV_X1 U5589 ( .A(n9807), .ZN(n9835) );
  AND3_X1 U5590 ( .A1(n4452), .A2(n5760), .A3(n6357), .ZN(n5882) );
  AND2_X1 U5591 ( .A1(n9768), .A2(n9819), .ZN(n9796) );
  AND2_X1 U5592 ( .A1(n6417), .A2(n6548), .ZN(n6439) );
  INV_X1 U5593 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5728) );
  INV_X1 U5594 ( .A(n4859), .ZN(n5688) );
  NAND2_X1 U5595 ( .A1(n5539), .A2(n5538), .ZN(n4697) );
  XNOR2_X1 U5596 ( .A(n4776), .B(n4775), .ZN(n6560) );
  NOR2_X1 U5597 ( .A1(n5393), .A2(n5330), .ZN(n4776) );
  AND2_X1 U5598 ( .A1(n6305), .A2(n6304), .ZN(n7597) );
  INV_X1 U5599 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n6026) );
  NAND2_X1 U5600 ( .A1(n6122), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n6136) );
  INV_X1 U5601 ( .A(n6134), .ZN(n6122) );
  NAND2_X1 U5602 ( .A1(n4690), .A2(n4689), .ZN(n4685) );
  NAND2_X1 U5603 ( .A1(n4663), .A2(n4662), .ZN(n8419) );
  OR2_X1 U5604 ( .A1(n4370), .A2(n4665), .ZN(n4662) );
  NAND2_X1 U5605 ( .A1(n4670), .A2(n4370), .ZN(n4667) );
  INV_X1 U5606 ( .A(n5987), .ZN(n5990) );
  OR2_X1 U5607 ( .A1(n6344), .A2(n8660), .ZN(n6341) );
  AOI21_X1 U5608 ( .B1(n8576), .B2(n8882), .A(n8575), .ZN(n8582) );
  AND2_X1 U5609 ( .A1(n8589), .A2(n8735), .ZN(n8622) );
  AND4_X1 U5610 ( .A1(n6115), .A2(n6114), .A3(n6113), .A4(n6112), .ZN(n7568)
         );
  NAND2_X1 U5611 ( .A1(n8823), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n4599) );
  NOR2_X1 U5612 ( .A1(n9233), .A2(n4605), .ZN(n9249) );
  AND2_X1 U5613 ( .A1(n8826), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n4605) );
  NOR2_X1 U5614 ( .A1(n9249), .A2(n9250), .ZN(n9248) );
  NAND2_X1 U5615 ( .A1(n9264), .A2(n9265), .ZN(n9263) );
  NOR2_X1 U5616 ( .A1(n9218), .A2(n4607), .ZN(n9353) );
  AND2_X1 U5617 ( .A1(n8830), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n4607) );
  NOR2_X1 U5618 ( .A1(n9353), .A2(n9354), .ZN(n9352) );
  NOR2_X1 U5619 ( .A1(n9352), .A2(n4606), .ZN(n9368) );
  AND2_X1 U5620 ( .A1(n9351), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n4606) );
  NAND2_X1 U5621 ( .A1(n9368), .A2(n9369), .ZN(n9367) );
  NOR2_X1 U5622 ( .A1(n9382), .A2(n4609), .ZN(n9399) );
  AND2_X1 U5623 ( .A1(n8833), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n4609) );
  NOR2_X1 U5624 ( .A1(n9399), .A2(n9400), .ZN(n9398) );
  NOR2_X1 U5625 ( .A1(n9398), .A2(n4608), .ZN(n8835) );
  AND2_X1 U5626 ( .A1(n9397), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n4608) );
  AND2_X1 U5627 ( .A1(n5162), .A2(n4677), .ZN(n4676) );
  INV_X1 U5628 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n4677) );
  NAND2_X1 U5629 ( .A1(n8930), .A2(n4480), .ZN(n8886) );
  NOR2_X1 U5630 ( .A1(n8890), .A2(n4481), .ZN(n4480) );
  NAND2_X1 U5631 ( .A1(n5258), .A2(n5257), .ZN(n8856) );
  AND2_X1 U5632 ( .A1(n8885), .A2(n6312), .ZN(n8904) );
  NAND2_X1 U5633 ( .A1(n8917), .A2(n8863), .ZN(n8894) );
  NAND2_X1 U5634 ( .A1(n8920), .A2(n9490), .ZN(n8923) );
  AND2_X1 U5635 ( .A1(n8625), .A2(n8862), .ZN(n8937) );
  AND2_X1 U5636 ( .A1(n8599), .A2(n8860), .ZN(n8647) );
  AND3_X1 U5637 ( .A1(n6252), .A2(n6251), .A3(n6250), .ZN(n8964) );
  NOR2_X1 U5638 ( .A1(n8962), .A2(n8961), .ZN(n8946) );
  AND3_X1 U5639 ( .A1(n6237), .A2(n6236), .A3(n6235), .ZN(n8980) );
  NOR2_X1 U5640 ( .A1(n8998), .A2(n7846), .ZN(n8978) );
  NOR2_X1 U5641 ( .A1(n8978), .A2(n8977), .ZN(n8976) );
  NAND2_X1 U5642 ( .A1(n9021), .A2(n9017), .ZN(n9011) );
  OR2_X1 U5643 ( .A1(n9011), .A2(n9140), .ZN(n8989) );
  NAND2_X1 U5644 ( .A1(n6161), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n6192) );
  NOR2_X1 U5645 ( .A1(n9078), .A2(n4486), .ZN(n9021) );
  NAND2_X1 U5646 ( .A1(n9025), .A2(n4487), .ZN(n4486) );
  AND2_X1 U5647 ( .A1(n8541), .A2(n9027), .ZN(n9046) );
  NAND2_X1 U5648 ( .A1(n6150), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n6174) );
  INV_X1 U5649 ( .A(n6152), .ZN(n6150) );
  OR2_X1 U5650 ( .A1(n6136), .A2(n8382), .ZN(n6152) );
  NOR2_X1 U5651 ( .A1(n7585), .A2(n7823), .ZN(n9079) );
  OR2_X1 U5652 ( .A1(n7406), .A2(n7560), .ZN(n7584) );
  OR2_X1 U5653 ( .A1(n7584), .A2(n8338), .ZN(n7585) );
  OAI21_X1 U5654 ( .B1(n4873), .B2(n4872), .A(n4380), .ZN(n4871) );
  NAND2_X1 U5655 ( .A1(n4415), .A2(n7150), .ZN(n4629) );
  INV_X1 U5656 ( .A(n8632), .ZN(n4630) );
  AND2_X1 U5657 ( .A1(n9477), .A2(n9561), .ZN(n7211) );
  NAND2_X1 U5658 ( .A1(n7211), .A2(n9567), .ZN(n7239) );
  NAND2_X1 U5659 ( .A1(n8481), .A2(n8474), .ZN(n7205) );
  NOR2_X1 U5660 ( .A1(n9476), .A2(n9473), .ZN(n9477) );
  NAND2_X1 U5661 ( .A1(n5993), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n6010) );
  OR2_X1 U5662 ( .A1(n6976), .A2(n7054), .ZN(n9476) );
  INV_X1 U5663 ( .A(n5951), .ZN(n5954) );
  NAND2_X1 U5664 ( .A1(n8589), .A2(n9503), .ZN(n6893) );
  NAND2_X1 U5665 ( .A1(n6897), .A2(n7029), .ZN(n9494) );
  INV_X1 U5666 ( .A(n6898), .ZN(n6934) );
  INV_X1 U5667 ( .A(n8864), .ZN(n4619) );
  INV_X1 U5668 ( .A(n4622), .ZN(n4621) );
  OAI21_X1 U5669 ( .B1(n8919), .B2(n4623), .A(n8900), .ZN(n4622) );
  INV_X1 U5670 ( .A(n8863), .ZN(n4623) );
  INV_X1 U5671 ( .A(n9568), .ZN(n9496) );
  AND2_X1 U5672 ( .A1(n5156), .A2(n5155), .ZN(n9614) );
  AND2_X1 U5673 ( .A1(n5141), .A2(n5140), .ZN(n9607) );
  OR2_X1 U5674 ( .A1(n5267), .A2(n6449), .ZN(n5060) );
  NAND2_X1 U5675 ( .A1(n6408), .A2(n6406), .ZN(n8660) );
  XNOR2_X1 U5676 ( .A(n5264), .B(n5263), .ZN(n8322) );
  OAI21_X1 U5677 ( .B1(n5261), .B2(n5260), .A(n5259), .ZN(n5264) );
  XNOR2_X1 U5678 ( .A(n5261), .B(n5260), .ZN(n7855) );
  AND2_X1 U5679 ( .A1(n4376), .A2(n4421), .ZN(n4885) );
  INV_X1 U5680 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5276) );
  AND2_X1 U5681 ( .A1(n5031), .A2(n4887), .ZN(n4886) );
  NOR2_X1 U5682 ( .A1(n4978), .A2(SI_17_), .ZN(n4979) );
  NAND2_X1 U5683 ( .A1(n4358), .A2(n5162), .ZN(n5179) );
  AND2_X1 U5684 ( .A1(n5129), .A2(n5128), .ZN(n6511) );
  NAND2_X1 U5685 ( .A1(n4741), .A2(n4738), .ZN(n5129) );
  NAND2_X1 U5686 ( .A1(n4741), .A2(n4965), .ZN(n5127) );
  AND2_X1 U5687 ( .A1(n5098), .A2(n5104), .ZN(n8828) );
  XNOR2_X1 U5688 ( .A(n4947), .B(SI_6_), .ZN(n5086) );
  AND2_X1 U5689 ( .A1(n6780), .A2(n5796), .ZN(n6941) );
  INV_X1 U5690 ( .A(n4704), .ZN(n4703) );
  NAND2_X1 U5691 ( .A1(n7932), .A2(n5850), .ZN(n7875) );
  NOR2_X1 U5692 ( .A1(n4904), .A2(n4908), .ZN(n5830) );
  INV_X1 U5693 ( .A(n8102), .ZN(n8080) );
  AND4_X1 U5694 ( .A1(n5445), .A2(n5444), .A3(n5443), .A4(n5442), .ZN(n6986)
         );
  NAND2_X1 U5695 ( .A1(n6939), .A2(n5798), .ZN(n6953) );
  AND3_X1 U5696 ( .A1(n5584), .A2(n5583), .A3(n5582), .ZN(n7893) );
  INV_X1 U5697 ( .A(n4699), .ZN(n4698) );
  OAI21_X1 U5698 ( .B1(n4700), .B2(n4702), .A(n6950), .ZN(n4699) );
  OR2_X1 U5699 ( .A1(n6949), .A2(n4701), .ZN(n4700) );
  INV_X1 U5700 ( .A(n7984), .ZN(n7968) );
  NAND2_X1 U5701 ( .A1(n7446), .A2(n5809), .ZN(n7522) );
  NAND2_X1 U5702 ( .A1(n4693), .A2(n4402), .ZN(n7385) );
  AND2_X1 U5703 ( .A1(n4693), .A2(n4694), .ZN(n7386) );
  NAND2_X1 U5704 ( .A1(n5818), .A2(n5817), .ZN(n7980) );
  INV_X1 U5705 ( .A(n7978), .ZN(n5817) );
  INV_X1 U5706 ( .A(n6419), .ZN(n8046) );
  AND2_X1 U5707 ( .A1(n7761), .A2(n5682), .ZN(n8081) );
  INV_X1 U5708 ( .A(n5844), .ZN(n8161) );
  INV_X1 U5709 ( .A(n6986), .ZN(n6783) );
  NAND4_X1 U5710 ( .A1(n5421), .A2(n5420), .A3(n5419), .A4(n5418), .ZN(n8003)
         );
  AND2_X1 U5711 ( .A1(n4456), .A2(n4455), .ZN(n6557) );
  NAND2_X1 U5712 ( .A1(n4457), .A2(n6562), .ZN(n4455) );
  AOI22_X1 U5713 ( .A1(n6801), .A2(P2_REG1_REG_5__SCAN_IN), .B1(n6805), .B2(
        n6800), .ZN(n6802) );
  AND2_X1 U5714 ( .A1(n4531), .A2(n4530), .ZN(n7003) );
  NAND2_X1 U5715 ( .A1(n7001), .A2(n4532), .ZN(n4530) );
  NAND2_X1 U5716 ( .A1(n7002), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n4531) );
  OAI21_X1 U5717 ( .B1(n7287), .B2(n7288), .A(n4537), .ZN(n7292) );
  NAND2_X1 U5718 ( .A1(n7122), .A2(n7295), .ZN(n4537) );
  NAND2_X1 U5719 ( .A1(n4748), .A2(n4747), .ZN(n8022) );
  NAND2_X1 U5720 ( .A1(n5675), .A2(n5674), .ZN(n5683) );
  NAND2_X1 U5721 ( .A1(n5673), .A2(n7751), .ZN(n5675) );
  INV_X1 U5722 ( .A(n9834), .ZN(n5501) );
  NAND2_X1 U5723 ( .A1(n7191), .A2(n5477), .ZN(n7174) );
  AND2_X1 U5724 ( .A1(n4818), .A2(n7654), .ZN(n7190) );
  NAND2_X1 U5725 ( .A1(n9775), .A2(n6665), .ZN(n8208) );
  INV_X1 U5726 ( .A(n9854), .ZN(n9852) );
  NAND2_X1 U5727 ( .A1(n8091), .A2(n8090), .ZN(n4858) );
  NAND2_X1 U5728 ( .A1(n5639), .A2(n5638), .ZN(n8261) );
  NAND2_X1 U5729 ( .A1(n5627), .A2(n5626), .ZN(n8267) );
  OAI21_X1 U5730 ( .B1(n8148), .B2(n4783), .A(n4780), .ZN(n8110) );
  NAND2_X1 U5731 ( .A1(n5618), .A2(n5617), .ZN(n8273) );
  AOI21_X1 U5732 ( .B1(n8137), .B2(n5616), .A(n5615), .ZN(n8122) );
  AND2_X1 U5733 ( .A1(n4840), .A2(n4839), .ZN(n8130) );
  NAND2_X1 U5734 ( .A1(n4840), .A2(n4841), .ZN(n8135) );
  NAND2_X1 U5735 ( .A1(n5596), .A2(n5595), .ZN(n8286) );
  AOI21_X1 U5736 ( .B1(n8155), .B2(n7714), .A(n4845), .ZN(n8144) );
  NAND2_X1 U5737 ( .A1(n5588), .A2(n5587), .ZN(n8292) );
  NAND2_X1 U5738 ( .A1(n5578), .A2(n5577), .ZN(n8298) );
  NAND2_X1 U5739 ( .A1(n5567), .A2(n5566), .ZN(n8304) );
  OAI21_X1 U5740 ( .B1(n4802), .B2(n8200), .A(n4547), .ZN(n8191) );
  NOR2_X1 U5741 ( .A1(n4543), .A2(n4549), .ZN(n8201) );
  NAND2_X1 U5742 ( .A1(n5355), .A2(n5354), .ZN(n7916) );
  NAND2_X1 U5743 ( .A1(n4822), .A2(n4823), .ZN(n7504) );
  OR2_X1 U5744 ( .A1(n7381), .A2(n4825), .ZN(n4822) );
  NAND2_X1 U5745 ( .A1(n5530), .A2(n5529), .ZN(n7976) );
  NAND2_X1 U5746 ( .A1(n4826), .A2(n4830), .ZN(n7543) );
  NAND2_X1 U5747 ( .A1(n7381), .A2(n4831), .ZN(n4826) );
  INV_X1 U5748 ( .A(n8254), .ZN(n8316) );
  NAND2_X1 U5749 ( .A1(n5517), .A2(n5516), .ZN(n7872) );
  AND2_X1 U5750 ( .A1(n4833), .A2(n4832), .ZN(n7443) );
  NAND2_X1 U5751 ( .A1(n7381), .A2(n5715), .ZN(n4833) );
  INV_X1 U5752 ( .A(n6863), .ZN(n6860) );
  OR2_X1 U5753 ( .A1(n9838), .A2(n9807), .ZN(n8254) );
  AND2_X1 U5754 ( .A1(n6403), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6548) );
  NAND2_X1 U5755 ( .A1(n8323), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5329) );
  NAND2_X1 U5756 ( .A1(n4859), .A2(n4860), .ZN(n5685) );
  INV_X1 U5757 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6460) );
  INV_X1 U5758 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6438) );
  XNOR2_X1 U5759 ( .A(n5425), .B(n5447), .ZN(n6920) );
  INV_X1 U5760 ( .A(n9614), .ZN(n8338) );
  AND4_X1 U5761 ( .A1(n6047), .A2(n6046), .A3(n6045), .A4(n6044), .ZN(n7471)
         );
  AND4_X1 U5762 ( .A1(n6103), .A2(n6102), .A3(n6101), .A4(n6100), .ZN(n7559)
         );
  NAND2_X1 U5763 ( .A1(n4681), .A2(n4683), .ZN(n8366) );
  NAND2_X1 U5764 ( .A1(n4690), .A2(n4682), .ZN(n4681) );
  NAND2_X1 U5765 ( .A1(n5235), .A2(n5234), .ZN(n9119) );
  INV_X1 U5766 ( .A(n4685), .ZN(n8402) );
  CLKBUF_X1 U5767 ( .A(n6768), .Z(n6769) );
  OR2_X1 U5768 ( .A1(n5267), .A2(n6448), .ZN(n5072) );
  AND4_X1 U5769 ( .A1(n6032), .A2(n6031), .A3(n6030), .A4(n6029), .ZN(n8490)
         );
  INV_X1 U5770 ( .A(n9017), .ZN(n9145) );
  NAND2_X1 U5771 ( .A1(n7459), .A2(n7460), .ZN(n4658) );
  AND4_X1 U5772 ( .A1(n6073), .A2(n6072), .A3(n6071), .A4(n6070), .ZN(n8750)
         );
  INV_X1 U5773 ( .A(n8748), .ZN(n7538) );
  INV_X1 U5774 ( .A(n4651), .ZN(n4650) );
  INV_X1 U5775 ( .A(n9501), .ZN(n9527) );
  INV_X1 U5776 ( .A(n8426), .ZN(n8455) );
  AND2_X1 U5777 ( .A1(n6311), .A2(n6277), .ZN(n8932) );
  INV_X1 U5778 ( .A(n9295), .ZN(n7823) );
  AND3_X1 U5779 ( .A1(n5285), .A2(n5284), .A3(n5283), .ZN(n8619) );
  INV_X1 U5780 ( .A(n8876), .ZN(n8921) );
  NAND2_X1 U5781 ( .A1(n6271), .A2(n6270), .ZN(n8938) );
  OR2_X1 U5782 ( .A1(n8369), .A2(n6265), .ZN(n6271) );
  INV_X1 U5783 ( .A(n7568), .ZN(n8519) );
  NAND2_X1 U5784 ( .A1(n4901), .A2(n5999), .ZN(n8753) );
  NAND2_X1 U5785 ( .A1(n5959), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5937) );
  OR2_X1 U5786 ( .A1(n5904), .A2(n5905), .ZN(n5906) );
  OR2_X1 U5787 ( .A1(n6408), .A2(n6407), .ZN(n8755) );
  NAND2_X1 U5788 ( .A1(n8759), .A2(n8758), .ZN(n8757) );
  INV_X1 U5789 ( .A(n4604), .ZN(n9313) );
  INV_X1 U5790 ( .A(n4602), .ZN(n9323) );
  INV_X1 U5791 ( .A(n4600), .ZN(n9322) );
  XNOR2_X1 U5792 ( .A(n8835), .B(n8836), .ZN(n9419) );
  INV_X1 U5793 ( .A(n9451), .ZN(n9446) );
  NAND2_X1 U5794 ( .A1(n4597), .A2(n8841), .ZN(n9453) );
  NAND2_X1 U5795 ( .A1(n9440), .A2(n9439), .ZN(n4597) );
  NAND2_X1 U5796 ( .A1(n4884), .A2(n8879), .ZN(n8899) );
  INV_X1 U5797 ( .A(n4484), .ZN(n8903) );
  AND2_X1 U5798 ( .A1(n5239), .A2(n5238), .ZN(n8934) );
  INV_X1 U5799 ( .A(n9119), .ZN(n8873) );
  AND2_X1 U5800 ( .A1(n5231), .A2(n5230), .ZN(n8957) );
  NAND2_X1 U5801 ( .A1(n4865), .A2(n4869), .ZN(n8960) );
  NAND2_X1 U5802 ( .A1(n7836), .A2(n4389), .ZN(n4865) );
  NAND2_X1 U5803 ( .A1(n5221), .A2(n5220), .ZN(n9135) );
  NAND2_X1 U5804 ( .A1(n7836), .A2(n7835), .ZN(n8975) );
  NAND2_X1 U5805 ( .A1(n9028), .A2(n8537), .ZN(n8999) );
  NAND2_X1 U5806 ( .A1(n4878), .A2(n4881), .ZN(n9005) );
  NAND2_X1 U5807 ( .A1(n4883), .A2(n4372), .ZN(n4878) );
  INV_X1 U5808 ( .A(n5182), .ZN(n9063) );
  AND2_X1 U5809 ( .A1(n5181), .A2(n5180), .ZN(n9068) );
  NAND2_X1 U5810 ( .A1(n4625), .A2(n8699), .ZN(n9056) );
  AND2_X1 U5811 ( .A1(n4889), .A2(n4435), .ZN(n9053) );
  NAND2_X1 U5812 ( .A1(n7827), .A2(n7826), .ZN(n9073) );
  INV_X1 U5813 ( .A(n9607), .ZN(n7560) );
  INV_X1 U5814 ( .A(n9601), .ZN(n7464) );
  NAND2_X1 U5815 ( .A1(n4870), .A2(n4873), .ZN(n7487) );
  NAND2_X1 U5816 ( .A1(n7361), .A2(n4875), .ZN(n4870) );
  AOI21_X1 U5817 ( .B1(n7361), .B2(n7360), .A(n4365), .ZN(n7409) );
  NAND2_X1 U5818 ( .A1(n7150), .A2(n8478), .ZN(n9467) );
  NAND2_X1 U5819 ( .A1(n7217), .A2(n6895), .ZN(n9482) );
  NAND2_X1 U5820 ( .A1(n9100), .A2(n8871), .ZN(n4642) );
  INV_X1 U5821 ( .A(n8872), .ZN(n4637) );
  NAND2_X1 U5822 ( .A1(n9521), .A2(n4626), .ZN(n9523) );
  NAND2_X1 U5823 ( .A1(n7030), .A2(n9591), .ZN(n4626) );
  XNOR2_X1 U5824 ( .A(n5225), .B(n5224), .ZN(n7076) );
  INV_X1 U5825 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n6462) );
  XNOR2_X1 U5826 ( .A(n4478), .B(n5092), .ZN(n6459) );
  INV_X1 U5827 ( .A(n5085), .ZN(n4569) );
  INV_X1 U5828 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6453) );
  AND2_X1 U5829 ( .A1(n4942), .A2(n4941), .ZN(n5076) );
  NAND2_X1 U5830 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n4610) );
  NAND2_X1 U5831 ( .A1(n4691), .A2(n4897), .ZN(P2_U3154) );
  NAND2_X1 U5832 ( .A1(n6618), .A2(n5785), .ZN(n6677) );
  INV_X1 U5833 ( .A(n4456), .ZN(n6555) );
  OAI21_X1 U5834 ( .B1(n4377), .B2(n4472), .A(n4468), .ZN(P2_U3201) );
  AOI21_X1 U5835 ( .B1(n4774), .B2(n6749), .A(n4469), .ZN(n4468) );
  NOR2_X1 U5836 ( .A1(n6370), .A2(n6371), .ZN(n6372) );
  NAND2_X1 U5837 ( .A1(n6368), .A2(n9836), .ZN(n5770) );
  OAI21_X1 U5838 ( .B1(n8255), .B2(n9838), .A(n4413), .ZN(P2_U3454) );
  NOR2_X1 U5839 ( .A1(n4437), .A2(n4552), .ZN(n4551) );
  OR2_X1 U5840 ( .A1(n8258), .A2(n8320), .ZN(n4553) );
  AOI21_X1 U5841 ( .B1(n7601), .B2(n7600), .A(n7599), .ZN(n7607) );
  OR2_X1 U5842 ( .A1(n7599), .A2(n6333), .ZN(n6355) );
  NAND2_X1 U5843 ( .A1(n5922), .A2(n5921), .ZN(n6726) );
  NAND2_X1 U5844 ( .A1(n8729), .A2(n8728), .ZN(n4451) );
  AOI21_X1 U5845 ( .B1(n9431), .B2(P1_ADDR_REG_19__SCAN_IN), .A(n8850), .ZN(
        n4615) );
  NAND2_X1 U5846 ( .A1(n4612), .A2(n8731), .ZN(n4611) );
  NAND2_X1 U5847 ( .A1(n8849), .A2(n4453), .ZN(n4616) );
  NOR2_X1 U5848 ( .A1(n9111), .A2(n9485), .ZN(n8926) );
  NAND2_X1 U5849 ( .A1(n9091), .A2(n9546), .ZN(n5317) );
  NAND2_X1 U5850 ( .A1(n4442), .A2(n9493), .ZN(n4640) );
  OR2_X1 U5851 ( .A1(n7284), .A2(n8000), .ZN(n4364) );
  NOR2_X1 U5852 ( .A1(n7475), .A2(n7359), .ZN(n4365) );
  NAND2_X1 U5853 ( .A1(n6053), .A2(n6052), .ZN(n4366) );
  NAND2_X1 U5854 ( .A1(n5223), .A2(n5004), .ZN(n4718) );
  INV_X2 U5855 ( .A(n5052), .ZN(n5103) );
  NAND2_X1 U5856 ( .A1(n4624), .A2(n8670), .ZN(n4367) );
  OR2_X1 U5857 ( .A1(n8292), .A2(n7957), .ZN(n7716) );
  INV_X1 U5858 ( .A(n8593), .ZN(n4565) );
  OR2_X1 U5859 ( .A1(n5688), .A2(P2_IR_REG_20__SCAN_IN), .ZN(n4368) );
  AND4_X1 U5860 ( .A1(n6974), .A2(n7029), .A3(n6897), .A4(n9501), .ZN(n4369)
         );
  NOR2_X1 U5861 ( .A1(n8360), .A2(n4668), .ZN(n4370) );
  AND2_X1 U5862 ( .A1(n4860), .A2(n5325), .ZN(n4371) );
  AND2_X1 U5863 ( .A1(n4392), .A2(n4912), .ZN(n4372) );
  AND2_X1 U5864 ( .A1(n4659), .A2(n7498), .ZN(n4373) );
  AND2_X1 U5865 ( .A1(n4683), .A2(n4403), .ZN(n4374) );
  OR2_X1 U5866 ( .A1(n9135), .A2(n8744), .ZN(n4375) );
  OR2_X1 U5867 ( .A1(n5903), .A2(n5902), .ZN(n5904) );
  AND3_X1 U5868 ( .A1(n5031), .A2(n4888), .A3(n4887), .ZN(n4376) );
  XNOR2_X1 U5869 ( .A(n8063), .B(n8062), .ZN(n4377) );
  INV_X1 U5870 ( .A(n7803), .ZN(n4855) );
  AND2_X1 U5871 ( .A1(n5477), .A2(n4364), .ZN(n4378) );
  OR2_X1 U5872 ( .A1(n7801), .A2(n7807), .ZN(n4379) );
  NAND2_X1 U5873 ( .A1(n9601), .A2(n7538), .ZN(n4380) );
  AND4_X1 U5874 ( .A1(n6060), .A2(n6059), .A3(n6058), .A4(n6057), .ZN(n7472)
         );
  INV_X1 U5875 ( .A(n8537), .ZN(n4636) );
  AND2_X1 U5876 ( .A1(n7472), .A2(n4876), .ZN(n4381) );
  NAND2_X1 U5877 ( .A1(n4417), .A2(n7689), .ZN(n4830) );
  OR2_X1 U5878 ( .A1(n4548), .A2(n5563), .ZN(n4382) );
  AND2_X1 U5879 ( .A1(n4875), .A2(n8634), .ZN(n4383) );
  AND2_X1 U5880 ( .A1(n4685), .A2(n6261), .ZN(n4384) );
  AND2_X1 U5881 ( .A1(n7830), .A2(n4435), .ZN(n4385) );
  INV_X1 U5882 ( .A(n7338), .ZN(n4655) );
  INV_X1 U5883 ( .A(n7360), .ZN(n4628) );
  OR2_X1 U5884 ( .A1(n9546), .A2(n4645), .ZN(n4386) );
  INV_X1 U5885 ( .A(n9516), .ZN(n9493) );
  INV_X1 U5886 ( .A(n5335), .ZN(n5399) );
  OR2_X1 U5887 ( .A1(n7418), .A2(n7412), .ZN(n4387) );
  AND2_X1 U5888 ( .A1(n5094), .A2(n4895), .ZN(n5113) );
  AND2_X1 U5889 ( .A1(n4703), .A2(n7932), .ZN(n4388) );
  OR2_X1 U5890 ( .A1(n7976), .A2(n7912), .ZN(n7695) );
  INV_X1 U5891 ( .A(n8890), .ZN(n9097) );
  NAND2_X1 U5892 ( .A1(n5036), .A2(n5035), .ZN(n8890) );
  INV_X1 U5893 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n5278) );
  INV_X1 U5894 ( .A(n9148), .ZN(n9025) );
  NAND2_X1 U5895 ( .A1(n5205), .A2(n5204), .ZN(n9148) );
  AND2_X1 U5896 ( .A1(n4375), .A2(n7835), .ZN(n4389) );
  NAND2_X1 U5897 ( .A1(n5084), .A2(n4946), .ZN(n4390) );
  OR2_X1 U5898 ( .A1(n8042), .A2(n8026), .ZN(n4391) );
  OR2_X1 U5899 ( .A1(n9148), .A2(n9047), .ZN(n4392) );
  XNOR2_X1 U5900 ( .A(n8257), .B(n8102), .ZN(n8090) );
  AND4_X1 U5901 ( .A1(n5433), .A2(n5432), .A3(n5431), .A4(n5430), .ZN(n7091)
         );
  NAND2_X1 U5902 ( .A1(n4670), .A2(n6204), .ZN(n8359) );
  INV_X1 U5903 ( .A(n7771), .ZN(n4512) );
  NOR2_X1 U5904 ( .A1(n5082), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n5094) );
  XNOR2_X1 U5905 ( .A(n5329), .B(P2_IR_REG_30__SCAN_IN), .ZN(n5334) );
  AND2_X1 U5906 ( .A1(n5094), .A2(n5025), .ZN(n5110) );
  OR2_X1 U5907 ( .A1(n9017), .A2(n9026), .ZN(n4393) );
  AND2_X1 U5908 ( .A1(n9135), .A2(n8744), .ZN(n4394) );
  AND2_X1 U5909 ( .A1(n4476), .A2(n4646), .ZN(n5270) );
  AND2_X1 U5910 ( .A1(n4600), .A2(n4599), .ZN(n4395) );
  AND2_X1 U5911 ( .A1(n4736), .A2(n4734), .ZN(n4396) );
  NOR2_X1 U5912 ( .A1(n9732), .A2(n8032), .ZN(n4397) );
  NAND2_X1 U5913 ( .A1(n5270), .A2(n5031), .ZN(n5293) );
  INV_X1 U5914 ( .A(n4843), .ZN(n4842) );
  OAI21_X1 U5915 ( .B1(n4845), .B2(n7714), .A(n4844), .ZN(n4843) );
  INV_X1 U5916 ( .A(n4548), .ZN(n4547) );
  OAI22_X1 U5917 ( .A1(n8200), .A2(n4801), .B1(n7994), .B2(n7931), .ZN(n4548)
         );
  AND2_X1 U5918 ( .A1(n5426), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n4398) );
  AND2_X1 U5919 ( .A1(n5227), .A2(n5226), .ZN(n8971) );
  INV_X1 U5920 ( .A(n8971), .ZN(n9130) );
  AND2_X1 U5921 ( .A1(n4644), .A2(n8871), .ZN(n4399) );
  AND2_X1 U5922 ( .A1(n8504), .A2(n8503), .ZN(n4400) );
  INV_X1 U5923 ( .A(n4817), .ZN(n4816) );
  NAND2_X1 U5924 ( .A1(n5711), .A2(n7654), .ZN(n4817) );
  INV_X1 U5925 ( .A(n8878), .ZN(n8919) );
  NAND2_X1 U5926 ( .A1(n7754), .A2(n7753), .ZN(n9279) );
  INV_X1 U5927 ( .A(n4488), .ZN(n8951) );
  NOR2_X1 U5928 ( .A1(n8989), .A2(n4490), .ZN(n4488) );
  AND2_X1 U5929 ( .A1(n5786), .A2(n5785), .ZN(n4401) );
  AND2_X1 U5930 ( .A1(n4694), .A2(n5805), .ZN(n4402) );
  AND2_X1 U5931 ( .A1(n4687), .A2(n4686), .ZN(n4403) );
  OR2_X1 U5932 ( .A1(n8273), .A2(n7903), .ZN(n7769) );
  INV_X1 U5933 ( .A(n7769), .ZN(n4835) );
  OR2_X1 U5934 ( .A1(n8086), .A2(n5722), .ZN(n4404) );
  NOR2_X1 U5935 ( .A1(n6107), .A2(n6106), .ZN(n4405) );
  AND2_X1 U5936 ( .A1(n8121), .A2(n7903), .ZN(n4406) );
  INV_X1 U5937 ( .A(n4684), .ZN(n4682) );
  NAND2_X1 U5938 ( .A1(n4688), .A2(n4689), .ZN(n4684) );
  AND4_X1 U5939 ( .A1(n8727), .A2(n8726), .A3(n8725), .A4(n8724), .ZN(n4407)
         );
  INV_X1 U5940 ( .A(n4801), .ZN(n4549) );
  NAND2_X1 U5941 ( .A1(n7916), .A2(n8202), .ZN(n4801) );
  NOR2_X1 U5942 ( .A1(n9904), .A2(n5206), .ZN(n4408) );
  NAND3_X1 U5943 ( .A1(n4351), .A2(n4893), .A3(n5094), .ZN(n4409) );
  NAND2_X1 U5944 ( .A1(n5270), .A2(n4886), .ZN(n4410) );
  AND4_X1 U5945 ( .A1(n5323), .A2(n5322), .A3(n5321), .A4(n5320), .ZN(n4411)
         );
  AND2_X1 U5946 ( .A1(n8286), .A2(n5844), .ZN(n7719) );
  INV_X1 U5947 ( .A(n7719), .ZN(n4844) );
  AND2_X1 U5948 ( .A1(n9130), .A2(n8743), .ZN(n4412) );
  AND2_X1 U5949 ( .A1(n4553), .A2(n4551), .ZN(n4413) );
  AND2_X1 U5950 ( .A1(n4955), .A2(n4954), .ZN(n4414) );
  AND2_X1 U5951 ( .A1(n7609), .A2(n7610), .ZN(n7697) );
  INV_X1 U5952 ( .A(n4796), .ZN(n4795) );
  NOR2_X1 U5953 ( .A1(n5659), .A2(n4797), .ZN(n4796) );
  INV_X1 U5954 ( .A(n9801), .ZN(n6879) );
  AND3_X1 U5955 ( .A1(n5415), .A2(n5414), .A3(n5413), .ZN(n9801) );
  AND2_X1 U5956 ( .A1(n4632), .A2(n4630), .ZN(n4415) );
  NAND2_X1 U5957 ( .A1(n4562), .A2(n4561), .ZN(n8701) );
  NAND2_X1 U5958 ( .A1(n7784), .A2(n4799), .ZN(n4416) );
  NAND2_X1 U5959 ( .A1(n7690), .A2(n4832), .ZN(n4417) );
  NAND2_X1 U5960 ( .A1(n5671), .A2(n5670), .ZN(n8094) );
  INV_X1 U5961 ( .A(n8094), .ZN(n5722) );
  AND2_X1 U5962 ( .A1(n9148), .A2(n9047), .ZN(n4418) );
  AND2_X1 U5963 ( .A1(n4858), .A2(n4857), .ZN(n4419) );
  AND3_X1 U5964 ( .A1(n5728), .A2(n5756), .A3(n5326), .ZN(n4420) );
  NOR2_X1 U5965 ( .A1(P1_IR_REG_27__SCAN_IN), .A2(P1_IR_REG_26__SCAN_IN), .ZN(
        n4421) );
  AND2_X1 U5966 ( .A1(n4862), .A2(n5346), .ZN(n4422) );
  AND2_X1 U5967 ( .A1(n9279), .A2(n8069), .ZN(n4423) );
  OR2_X1 U5968 ( .A1(n5052), .A2(n9243), .ZN(n4424) );
  AND2_X1 U5969 ( .A1(n7692), .A2(n7691), .ZN(n4425) );
  AND2_X1 U5970 ( .A1(n5538), .A2(n4696), .ZN(n4426) );
  AND2_X1 U5971 ( .A1(n8468), .A2(n8670), .ZN(n4427) );
  AND2_X1 U5972 ( .A1(n9052), .A2(n8699), .ZN(n4428) );
  AND2_X1 U5973 ( .A1(n5810), .A2(n5809), .ZN(n4429) );
  AND2_X1 U5974 ( .A1(n8880), .A2(n8879), .ZN(n4430) );
  INV_X1 U5975 ( .A(n6814), .ZN(n4753) );
  AND2_X1 U5976 ( .A1(n4664), .A2(n6201), .ZN(n4431) );
  OR2_X1 U5977 ( .A1(n8280), .A2(n7958), .ZN(n7770) );
  OR2_X1 U5978 ( .A1(n5683), .A2(n8081), .ZN(n7762) );
  NAND2_X1 U5979 ( .A1(n4372), .A2(n7833), .ZN(n4432) );
  INV_X1 U5980 ( .A(n4665), .ZN(n4664) );
  NAND2_X1 U5981 ( .A1(n4669), .A2(n4666), .ZN(n4665) );
  NAND2_X1 U5982 ( .A1(n7164), .A2(n9473), .ZN(n7163) );
  INV_X1 U5983 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n4775) );
  INV_X1 U5984 ( .A(n7007), .ZN(n4532) );
  AND2_X1 U5985 ( .A1(n8601), .A2(n8550), .ZN(n4433) );
  NOR2_X1 U5986 ( .A1(n5082), .A2(n5152), .ZN(n5163) );
  AND2_X1 U5987 ( .A1(n5006), .A2(n9938), .ZN(n4434) );
  INV_X1 U5988 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n4894) );
  NAND2_X1 U5989 ( .A1(n7033), .A2(n6906), .ZN(n8666) );
  XNOR2_X1 U5990 ( .A(n5386), .B(P2_IR_REG_2__SCAN_IN), .ZN(n6535) );
  NAND2_X1 U5991 ( .A1(n5125), .A2(n5124), .ZN(n9590) );
  INV_X1 U5992 ( .A(n9590), .ZN(n4876) );
  NOR2_X1 U5993 ( .A1(n8756), .A2(n7029), .ZN(n6932) );
  NAND2_X1 U5994 ( .A1(n9083), .A2(n8746), .ZN(n4435) );
  NAND2_X1 U5995 ( .A1(n7250), .A2(n6039), .ZN(n7337) );
  AOI21_X1 U5996 ( .B1(n4883), .B2(n4912), .A(n4911), .ZN(n9020) );
  NAND2_X1 U5997 ( .A1(n4658), .A2(n6096), .ZN(n7497) );
  OR2_X1 U5998 ( .A1(n6917), .A2(n6920), .ZN(n4436) );
  NAND2_X1 U5999 ( .A1(n5247), .A2(n5246), .ZN(n9103) );
  INV_X1 U6000 ( .A(n9103), .ZN(n4482) );
  AND3_X1 U6001 ( .A1(n4707), .A2(n4706), .A3(n4705), .ZN(n5356) );
  XNOR2_X1 U6002 ( .A(n5366), .B(P2_IR_REG_1__SCAN_IN), .ZN(n6421) );
  NAND2_X1 U6003 ( .A1(n8512), .A2(n8693), .ZN(n8634) );
  INV_X1 U6004 ( .A(n8634), .ZN(n4872) );
  AND4_X1 U6005 ( .A1(n5488), .A2(n5487), .A3(n5486), .A4(n5485), .ZN(n7389)
         );
  AND2_X1 U6006 ( .A1(n8257), .A2(n8316), .ZN(n4437) );
  AND2_X1 U6007 ( .A1(n8828), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n4438) );
  NAND2_X1 U6008 ( .A1(n5661), .A2(n5660), .ZN(n8086) );
  INV_X1 U6009 ( .A(n8086), .ZN(n4721) );
  AND2_X1 U6010 ( .A1(n8257), .A2(n8102), .ZN(n4439) );
  OR2_X1 U6011 ( .A1(n7545), .A2(n4803), .ZN(n4802) );
  OR2_X1 U6012 ( .A1(n4969), .A2(n10026), .ZN(n4440) );
  INV_X1 U6013 ( .A(n7958), .ZN(n8149) );
  AND2_X1 U6014 ( .A1(n5614), .A2(n5613), .ZN(n7958) );
  AND2_X1 U6015 ( .A1(n5822), .A2(n5821), .ZN(n4441) );
  INV_X1 U6016 ( .A(n4899), .ZN(n4719) );
  INV_X1 U6017 ( .A(n7049), .ZN(n7042) );
  AND2_X1 U6018 ( .A1(n7269), .A2(n4876), .ZN(n7366) );
  INV_X1 U6019 ( .A(n6753), .ZN(n6805) );
  NAND2_X1 U6020 ( .A1(n5726), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5755) );
  NAND2_X1 U6021 ( .A1(n4813), .A2(n4811), .ZN(n7223) );
  NAND2_X1 U6022 ( .A1(n4386), .A2(n9618), .ZN(n4442) );
  INV_X1 U6023 ( .A(n4452), .ZN(n5772) );
  NOR2_X1 U6024 ( .A1(n7294), .A2(n4769), .ZN(n4443) );
  AND2_X1 U6025 ( .A1(n4629), .A2(n8683), .ZN(n4444) );
  INV_X1 U6026 ( .A(n4763), .ZN(n4761) );
  NAND2_X1 U6027 ( .A1(n9665), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n4763) );
  AND2_X1 U6028 ( .A1(n4751), .A2(n4387), .ZN(n4445) );
  INV_X1 U6029 ( .A(n8042), .ZN(n4759) );
  INV_X1 U6030 ( .A(n9729), .ZN(n4472) );
  NAND2_X1 U6031 ( .A1(n4650), .A2(n6708), .ZN(n6711) );
  OR2_X1 U6032 ( .A1(n9513), .A2(n8722), .ZN(n9613) );
  INV_X1 U6033 ( .A(n7160), .ZN(n7068) );
  NAND2_X1 U6034 ( .A1(n5932), .A2(n6708), .ZN(n6724) );
  OR2_X1 U6035 ( .A1(n8056), .A2(n8030), .ZN(n4446) );
  AND2_X1 U6036 ( .A1(n6813), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n4447) );
  AND2_X1 U6037 ( .A1(n4755), .A2(n6813), .ZN(n4448) );
  INV_X1 U6038 ( .A(SI_13_), .ZN(n4734) );
  AND2_X1 U6039 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(P2_U3151), .ZN(n4449) );
  INV_X1 U6040 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n4746) );
  INV_X1 U6041 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n4460) );
  INV_X1 U6042 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n4754) );
  AOI21_X1 U6043 ( .B1(n4738), .B2(n4966), .A(n4737), .ZN(n4736) );
  INV_X1 U6044 ( .A(n4966), .ZN(n4454) );
  OAI21_X1 U6045 ( .B1(n7951), .B2(n5847), .A(n5846), .ZN(n5849) );
  NOR3_X1 U6046 ( .A1(n7901), .A2(n6377), .A3(n6376), .ZN(n6382) );
  OAI21_X1 U6047 ( .B1(n5739), .B2(P2_D_REG_0__SCAN_IN), .A(n6443), .ZN(n4452)
         );
  AND3_X2 U6048 ( .A1(n4466), .A2(n4411), .A3(n5356), .ZN(n4859) );
  OAI21_X1 U6049 ( .B1(n4400), .B2(n4450), .A(n8512), .ZN(n8505) );
  NAND3_X1 U6050 ( .A1(n4451), .A2(n8740), .A3(n4407), .ZN(P1_U3242) );
  MUX2_X1 U6051 ( .A(n8470), .B(n8469), .S(n8514), .Z(n8480) );
  NAND4_X1 U6052 ( .A1(n4646), .A2(n4351), .A3(n4893), .A4(n4376), .ZN(n5033)
         );
  NAND2_X1 U6053 ( .A1(n4574), .A2(n8572), .ZN(n8576) );
  AND2_X1 U6054 ( .A1(n8569), .A2(n8625), .ZN(n4580) );
  NAND2_X1 U6055 ( .A1(n4578), .A2(n4577), .ZN(n4576) );
  NAND2_X1 U6056 ( .A1(n4585), .A2(n4583), .ZN(n4582) );
  XNOR2_X1 U6057 ( .A(n5778), .B(n9763), .ZN(n6575) );
  NAND2_X1 U6058 ( .A1(n6767), .A2(n5976), .ZN(n5987) );
  NAND2_X1 U6059 ( .A1(n4667), .A2(n4669), .ZN(n6230) );
  NAND2_X1 U6060 ( .A1(n5920), .A2(n5916), .ZN(n6628) );
  NAND2_X1 U6061 ( .A1(n6893), .A2(n5913), .ZN(n5914) );
  NAND2_X1 U6062 ( .A1(n5947), .A2(n6710), .ZN(n6712) );
  NOR2_X1 U6063 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n5151) );
  NAND2_X1 U6064 ( .A1(n6824), .A2(n6825), .ZN(n6768) );
  OAI21_X1 U6065 ( .B1(n8392), .B2(n8389), .A(n8388), .ZN(n8348) );
  OAI21_X1 U6066 ( .B1(n8875), .B2(n8874), .A(n4903), .ZN(n8929) );
  NOR2_X1 U6067 ( .A1(n9039), .A2(n4432), .ZN(n4877) );
  AOI21_X1 U6068 ( .B1(n7361), .B2(n4383), .A(n4871), .ZN(n7562) );
  NAND2_X1 U6069 ( .A1(n4643), .A2(n4644), .ZN(n9169) );
  NAND2_X2 U6070 ( .A1(n7079), .A2(n5803), .ZN(n5804) );
  INV_X1 U6071 ( .A(n4559), .ZN(n4467) );
  AND2_X2 U6072 ( .A1(n5319), .A2(n5393), .ZN(n4466) );
  NAND2_X4 U6073 ( .A1(n4805), .A2(n4560), .ZN(n6436) );
  NAND2_X2 U6074 ( .A1(n4920), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n4560) );
  NAND2_X2 U6075 ( .A1(n4919), .A2(n4918), .ZN(n4805) );
  AND3_X2 U6076 ( .A1(n4476), .A2(n4646), .A3(n4885), .ZN(n5277) );
  NAND2_X1 U6077 ( .A1(n8930), .A2(n8916), .ZN(n8911) );
  INV_X1 U6078 ( .A(n4492), .ZN(n8931) );
  NAND3_X1 U6079 ( .A1(n6897), .A2(n9501), .A3(n7029), .ZN(n9497) );
  NAND2_X1 U6080 ( .A1(n4503), .A2(n4500), .ZN(n7746) );
  NAND2_X1 U6081 ( .A1(n4501), .A2(n7747), .ZN(n4500) );
  NAND2_X1 U6082 ( .A1(n4502), .A2(n7764), .ZN(n4501) );
  NAND2_X1 U6083 ( .A1(n4722), .A2(n5722), .ZN(n4502) );
  NAND2_X1 U6084 ( .A1(n4504), .A2(n7732), .ZN(n4503) );
  NAND2_X1 U6085 ( .A1(n4505), .A2(n7742), .ZN(n4504) );
  NAND2_X1 U6086 ( .A1(n4722), .A2(n4721), .ZN(n4505) );
  AND2_X1 U6087 ( .A1(n4508), .A2(n4507), .ZN(n7702) );
  NAND3_X1 U6088 ( .A1(n4526), .A2(n4524), .A3(n4523), .ZN(n4522) );
  OR2_X1 U6089 ( .A1(n7320), .A2(n7319), .ZN(n4536) );
  NAND2_X1 U6090 ( .A1(n7292), .A2(n7291), .ZN(n7318) );
  INV_X2 U6091 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n4709) );
  NOR2_X2 U6092 ( .A1(n7544), .A2(n7692), .ZN(n7545) );
  NAND2_X2 U6093 ( .A1(n5693), .A2(n8057), .ZN(n5379) );
  NAND2_X1 U6094 ( .A1(n5410), .A2(n7751), .ZN(n5415) );
  INV_X1 U6095 ( .A(n4802), .ZN(n4543) );
  OAI21_X1 U6096 ( .B1(n4543), .B2(n4382), .A(n4544), .ZN(n8180) );
  INV_X1 U6097 ( .A(n8180), .ZN(n5576) );
  OAI21_X2 U6098 ( .B1(n8156), .B2(n8146), .A(n8145), .ZN(n8148) );
  AOI21_X2 U6099 ( .B1(n8168), .B2(n8157), .A(n8158), .ZN(n8156) );
  NAND2_X1 U6100 ( .A1(n4859), .A2(n4558), .ZN(n5348) );
  NAND2_X1 U6101 ( .A1(n5348), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5349) );
  NAND3_X1 U6102 ( .A1(n4805), .A2(P2_DATAO_REG_1__SCAN_IN), .A3(n4560), .ZN(
        n4921) );
  NAND3_X1 U6103 ( .A1(n4805), .A2(P2_DATAO_REG_4__SCAN_IN), .A3(n4560), .ZN(
        n4745) );
  NAND2_X1 U6104 ( .A1(n4563), .A2(n8557), .ZN(n8561) );
  NAND3_X1 U6105 ( .A1(n4949), .A2(n4567), .A3(n4942), .ZN(n4570) );
  NAND2_X1 U6106 ( .A1(n4942), .A2(n4732), .ZN(n5085) );
  NAND3_X1 U6107 ( .A1(n4581), .A2(n4579), .A3(n8706), .ZN(n4578) );
  OAI22_X1 U6108 ( .A1(n8530), .A2(n8734), .B1(n8532), .B2(n8531), .ZN(n4584)
         );
  NAND2_X1 U6109 ( .A1(n5135), .A2(SI_13_), .ZN(n4591) );
  NAND2_X1 U6110 ( .A1(n4589), .A2(n4587), .ZN(n5170) );
  NAND3_X1 U6111 ( .A1(n4591), .A2(n4590), .A3(n4440), .ZN(n4589) );
  NAND2_X1 U6112 ( .A1(n4589), .A2(n4970), .ZN(n5168) );
  NAND2_X1 U6113 ( .A1(n4960), .A2(n4594), .ZN(n5119) );
  NAND2_X1 U6114 ( .A1(n4960), .A2(n4592), .ZN(n4735) );
  MUX2_X1 U6115 ( .A(P1_REG2_REG_1__SCAN_IN), .B(n6690), .S(n8763), .Z(n8759)
         );
  XNOR2_X1 U6116 ( .A(n4610), .B(P1_IR_REG_1__SCAN_IN), .ZN(n8763) );
  NAND3_X1 U6117 ( .A1(n4616), .A2(n4615), .A3(n4611), .ZN(P1_U3262) );
  NAND2_X4 U6118 ( .A1(n5052), .A2(n6436), .ZN(n5267) );
  XNOR2_X2 U6119 ( .A(n4617), .B(P1_IR_REG_27__SCAN_IN), .ZN(n5287) );
  NAND2_X1 U6120 ( .A1(n5291), .A2(n5032), .ZN(n4617) );
  NAND2_X1 U6121 ( .A1(n8918), .A2(n8919), .ZN(n8917) );
  OAI21_X1 U6122 ( .B1(n8918), .B2(n4623), .A(n4621), .ZN(n8893) );
  NAND2_X1 U6123 ( .A1(n4620), .A2(n4618), .ZN(n8866) );
  NAND2_X1 U6124 ( .A1(n8918), .A2(n4621), .ZN(n4620) );
  NAND2_X1 U6125 ( .A1(n4624), .A2(n4427), .ZN(n6971) );
  NAND3_X1 U6126 ( .A1(n7033), .A2(n6906), .A3(n6907), .ZN(n4624) );
  NAND2_X1 U6127 ( .A1(n4625), .A2(n4428), .ZN(n9054) );
  NAND3_X1 U6128 ( .A1(n4629), .A2(n4628), .A3(n8683), .ZN(n7362) );
  NAND2_X1 U6129 ( .A1(n7150), .A2(n4632), .ZN(n7264) );
  OAI21_X2 U6130 ( .B1(n9045), .B2(n4634), .A(n4633), .ZN(n8998) );
  OAI21_X1 U6131 ( .B1(n4639), .B2(n9099), .A(n4442), .ZN(n4638) );
  NOR2_X1 U6132 ( .A1(n9099), .A2(n4642), .ZN(n4643) );
  OAI21_X1 U6133 ( .B1(n8872), .B2(n4640), .A(n4638), .ZN(P1_U3519) );
  NAND2_X1 U6134 ( .A1(n4651), .A2(n6708), .ZN(n5947) );
  NAND3_X1 U6135 ( .A1(n5922), .A2(n5921), .A3(n5932), .ZN(n4651) );
  NAND2_X1 U6136 ( .A1(n7249), .A2(n7251), .ZN(n7250) );
  OAI211_X1 U6137 ( .C1(n6039), .C2(n4655), .A(n4652), .B(n4366), .ZN(n7467)
         );
  NAND2_X1 U6138 ( .A1(n7249), .A2(n4653), .ZN(n4652) );
  INV_X1 U6139 ( .A(n7251), .ZN(n4654) );
  NAND2_X1 U6140 ( .A1(n7459), .A2(n4373), .ZN(n4657) );
  XNOR2_X1 U6141 ( .A(n4661), .B(n6321), .ZN(n5931) );
  NAND2_X1 U6142 ( .A1(n8411), .A2(n4431), .ZN(n4663) );
  NAND2_X1 U6143 ( .A1(n8411), .A2(n6201), .ZN(n4670) );
  NAND2_X1 U6144 ( .A1(n4358), .A2(n4674), .ZN(n4672) );
  NAND2_X1 U6145 ( .A1(n8400), .A2(n4680), .ZN(n4679) );
  NAND2_X1 U6146 ( .A1(n8400), .A2(n8399), .ZN(n4690) );
  INV_X1 U6147 ( .A(n8398), .ZN(n4689) );
  NAND3_X1 U6148 ( .A1(n5879), .A2(n4692), .A3(n7954), .ZN(n4691) );
  NAND2_X1 U6149 ( .A1(n7277), .A2(n7278), .ZN(n4693) );
  INV_X1 U6150 ( .A(n5804), .ZN(n4695) );
  NAND2_X1 U6151 ( .A1(n5539), .A2(n4426), .ZN(n5564) );
  NAND2_X1 U6152 ( .A1(n4697), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5540) );
  NAND2_X1 U6153 ( .A1(n7446), .A2(n4429), .ZN(n7520) );
  NAND2_X1 U6154 ( .A1(n7980), .A2(n4441), .ZN(n7909) );
  OAI21_X2 U6155 ( .B1(n6780), .B2(n4700), .A(n4698), .ZN(n7081) );
  NAND2_X1 U6156 ( .A1(n5850), .A2(n7958), .ZN(n4704) );
  NAND2_X1 U6157 ( .A1(n4710), .A2(n4714), .ZN(n5010) );
  NAND2_X1 U6158 ( .A1(n5223), .A2(n4711), .ZN(n4710) );
  INV_X1 U6159 ( .A(n4724), .ZN(n7744) );
  NAND2_X1 U6160 ( .A1(n5184), .A2(n4727), .ZN(n4725) );
  NAND2_X1 U6161 ( .A1(n4725), .A2(n4726), .ZN(n5215) );
  NAND2_X1 U6162 ( .A1(n4735), .A2(n4736), .ZN(n5135) );
  NAND3_X1 U6163 ( .A1(n4745), .A2(n4744), .A3(n4743), .ZN(n4940) );
  NAND3_X1 U6164 ( .A1(n4920), .A2(P2_ADDR_REG_19__SCAN_IN), .A3(
        P1_DATAO_REG_4__SCAN_IN), .ZN(n4743) );
  NAND3_X1 U6165 ( .A1(n4919), .A2(n4918), .A3(P1_DATAO_REG_4__SCAN_IN), .ZN(
        n4744) );
  INV_X4 U6166 ( .A(n6436), .ZN(n6431) );
  INV_X1 U6167 ( .A(n4751), .ZN(n7413) );
  OAI22_X1 U6168 ( .A1(n6745), .A2(n4752), .B1(n6814), .B2(n6813), .ZN(n6919)
         );
  INV_X1 U6169 ( .A(n6745), .ZN(n4755) );
  NOR2_X1 U6170 ( .A1(n9675), .A2(n4761), .ZN(n8026) );
  NAND3_X1 U6171 ( .A1(n4757), .A2(n4758), .A3(n4756), .ZN(n9694) );
  NAND4_X1 U6172 ( .A1(n4757), .A2(n4758), .A3(n4756), .A4(
        P2_REG2_REG_15__SCAN_IN), .ZN(n4762) );
  INV_X1 U6173 ( .A(n4762), .ZN(n9692) );
  INV_X1 U6174 ( .A(n7293), .ZN(n4764) );
  NAND2_X1 U6175 ( .A1(n4767), .A2(n4766), .ZN(n4765) );
  OAI21_X1 U6176 ( .B1(n4768), .B2(n7297), .A(n4765), .ZN(n7325) );
  NAND2_X1 U6177 ( .A1(n8032), .A2(n4772), .ZN(n4770) );
  NOR2_X1 U6178 ( .A1(n9734), .A2(n9733), .ZN(n9732) );
  INV_X1 U6179 ( .A(n4777), .ZN(n8109) );
  OR2_X1 U6180 ( .A1(n8100), .A2(n4795), .ZN(n4788) );
  NAND2_X1 U6181 ( .A1(n8100), .A2(n5648), .ZN(n4798) );
  OR2_X1 U6182 ( .A1(n8100), .A2(n4792), .ZN(n4791) );
  NAND3_X1 U6183 ( .A1(n4810), .A2(n4808), .A3(n5438), .ZN(n7089) );
  NAND3_X1 U6184 ( .A1(n5436), .A2(n4916), .A3(n6835), .ZN(n4810) );
  NAND2_X1 U6185 ( .A1(n6990), .A2(n4814), .ZN(n4813) );
  NAND2_X1 U6186 ( .A1(n4821), .A2(n7381), .ZN(n4819) );
  NAND3_X1 U6187 ( .A1(n4820), .A2(n4819), .A3(n7609), .ZN(n8199) );
  NAND2_X1 U6188 ( .A1(n8155), .A2(n4837), .ZN(n4836) );
  NAND2_X1 U6189 ( .A1(n8091), .A2(n4851), .ZN(n4850) );
  NAND2_X1 U6190 ( .A1(n4850), .A2(n4852), .ZN(n7765) );
  NAND2_X1 U6191 ( .A1(n5721), .A2(n8102), .ZN(n4857) );
  NAND2_X1 U6192 ( .A1(n5734), .A2(n4862), .ZN(n5345) );
  NAND2_X1 U6193 ( .A1(n7049), .A2(n7050), .ZN(n7155) );
  AND2_X1 U6194 ( .A1(n8466), .A2(n8477), .ZN(n7049) );
  NAND2_X1 U6195 ( .A1(n7836), .A2(n4866), .ZN(n4863) );
  NAND2_X1 U6196 ( .A1(n4863), .A2(n4864), .ZN(n8945) );
  OAI22_X4 U6197 ( .A1(n7274), .A2(n7273), .B1(n8751), .B2(n7343), .ZN(n7361)
         );
  NOR2_X1 U6198 ( .A1(n4877), .A2(n4879), .ZN(n8988) );
  NAND2_X1 U6199 ( .A1(n4884), .A2(n4430), .ZN(n8902) );
  NAND2_X1 U6200 ( .A1(n7827), .A2(n4890), .ZN(n4892) );
  NAND2_X1 U6201 ( .A1(n4892), .A2(n4385), .ZN(n7832) );
  CLKBUF_X1 U6202 ( .A(n4892), .Z(n4889) );
  INV_X1 U6203 ( .A(n4889), .ZN(n9072) );
  NAND3_X1 U6204 ( .A1(n5094), .A2(n4351), .A3(n4895), .ZN(n5273) );
  NOR2_X4 U6205 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5048) );
  NAND3_X1 U6206 ( .A1(n5048), .A2(n5061), .A3(n4896), .ZN(n5080) );
  AND2_X1 U6207 ( .A1(n8902), .A2(n8901), .ZN(n9102) );
  NAND2_X1 U6208 ( .A1(n5933), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n5953) );
  AND2_X4 U6209 ( .A1(n5340), .A2(n5333), .ZN(n5398) );
  NAND2_X1 U6210 ( .A1(n5280), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5281) );
  NOR2_X1 U6211 ( .A1(n7596), .A2(n6306), .ZN(n7599) );
  AND2_X2 U6212 ( .A1(n5965), .A2(n5964), .ZN(n6970) );
  NAND2_X1 U6213 ( .A1(n5933), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5909) );
  INV_X1 U6214 ( .A(n7783), .ZN(n5711) );
  AND2_X1 U6215 ( .A1(n5901), .A2(n5900), .ZN(n4897) );
  NOR2_X1 U6216 ( .A1(n7110), .A2(n7104), .ZN(n4898) );
  NOR2_X1 U6217 ( .A1(n5003), .A2(n5224), .ZN(n4899) );
  AND2_X1 U6218 ( .A1(n5959), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n4900) );
  AND2_X1 U6219 ( .A1(n5998), .A2(n5997), .ZN(n4901) );
  AND2_X1 U6220 ( .A1(n4363), .A2(n9470), .ZN(n4902) );
  OR2_X1 U6221 ( .A1(n8873), .A2(n8950), .ZN(n4903) );
  INV_X1 U6222 ( .A(n8750), .ZN(n7359) );
  AND2_X1 U6223 ( .A1(n6318), .A2(n6317), .ZN(n8867) );
  XNOR2_X1 U6224 ( .A(n4927), .B(n4924), .ZN(n5041) );
  AND3_X1 U6225 ( .A1(n8475), .A2(n8474), .A3(n8734), .ZN(n4906) );
  AND2_X1 U6226 ( .A1(n5829), .A2(n7885), .ZN(n4908) );
  OR2_X1 U6227 ( .A1(n9546), .A2(n5316), .ZN(n4909) );
  INV_X1 U6228 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n4931) );
  NAND2_X1 U6229 ( .A1(n8657), .A2(n8622), .ZN(n9062) );
  INV_X1 U6230 ( .A(n9062), .ZN(n9489) );
  INV_X1 U6231 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n4922) );
  INV_X1 U6232 ( .A(n9047), .ZN(n9009) );
  INV_X1 U6233 ( .A(n8384), .ZN(n9076) );
  NAND2_X1 U6234 ( .A1(n7366), .A2(n9601), .ZN(n7406) );
  AND2_X1 U6235 ( .A1(n9154), .A2(n9034), .ZN(n4911) );
  OR2_X1 U6236 ( .A1(n9154), .A2(n9034), .ZN(n4912) );
  AND2_X1 U6237 ( .A1(n8273), .A2(n8138), .ZN(n4913) );
  OR2_X1 U6238 ( .A1(n6565), .A2(n6647), .ZN(n4914) );
  INV_X1 U6239 ( .A(n7384), .ZN(n5805) );
  AND3_X1 U6240 ( .A1(n8707), .A2(n9006), .A3(n8706), .ZN(n4915) );
  AND2_X1 U6241 ( .A1(n6789), .A2(n6790), .ZN(n4916) );
  OR2_X1 U6242 ( .A1(n9090), .A2(n9089), .ZN(n9644) );
  OR2_X1 U6243 ( .A1(n9090), .A2(n6330), .ZN(n9618) );
  AND2_X1 U6244 ( .A1(n8511), .A2(n8684), .ZN(n8503) );
  INV_X1 U6245 ( .A(n8734), .ZN(n8514) );
  NAND2_X1 U6246 ( .A1(n8515), .A2(n8514), .ZN(n8516) );
  INV_X1 U6247 ( .A(n7091), .ZN(n5434) );
  NOR2_X1 U6248 ( .A1(n4855), .A2(n7732), .ZN(n7749) );
  INV_X1 U6249 ( .A(n8383), .ZN(n7828) );
  INV_X1 U6250 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5026) );
  INV_X1 U6251 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5336) );
  INV_X1 U6252 ( .A(n7998), .ZN(n5500) );
  INV_X1 U6253 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n5327) );
  OR2_X1 U6254 ( .A1(n8957), .A2(n4354), .ZN(n6255) );
  INV_X1 U6255 ( .A(n8696), .ZN(n7565) );
  INV_X1 U6256 ( .A(n7806), .ZN(n7807) );
  NOR2_X1 U6257 ( .A1(n7320), .A2(n7296), .ZN(n7324) );
  INV_X1 U6258 ( .A(n8117), .ZN(n5636) );
  AND2_X1 U6259 ( .A1(n8304), .A2(n8193), .ZN(n5574) );
  XNOR2_X1 U6260 ( .A(n9745), .B(n5780), .ZN(n7619) );
  NAND2_X1 U6261 ( .A1(n6108), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n6134) );
  INV_X1 U6262 ( .A(n6010), .ZN(n6008) );
  INV_X1 U6263 ( .A(n6208), .ZN(n6207) );
  NAND2_X1 U6264 ( .A1(n6040), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n6067) );
  INV_X1 U6265 ( .A(n5213), .ZN(n4993) );
  AND2_X1 U6266 ( .A1(n4973), .A2(n5169), .ZN(n4974) );
  NAND2_X1 U6267 ( .A1(n4963), .A2(n5118), .ZN(n4966) );
  INV_X1 U6268 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n9940) );
  INV_X1 U6269 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n10058) );
  INV_X1 U6270 ( .A(n5871), .ZN(n5872) );
  NOR2_X1 U6271 ( .A1(n5494), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5493) );
  INV_X1 U6272 ( .A(n7523), .ZN(n5810) );
  OAI21_X1 U6273 ( .B1(n7809), .B2(n7808), .A(n7807), .ZN(n7810) );
  INV_X1 U6274 ( .A(n5599), .ZN(n7757) );
  NOR2_X1 U6275 ( .A1(n6922), .A2(n7014), .ZN(n6924) );
  INV_X1 U6276 ( .A(n8039), .ZN(n8030) );
  INV_X1 U6277 ( .A(n7800), .ZN(n7737) );
  NOR2_X1 U6278 ( .A1(n5652), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n5663) );
  NOR2_X1 U6279 ( .A1(n5568), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n5579) );
  NOR2_X1 U6280 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n5400) );
  NOR2_X1 U6281 ( .A1(n9854), .A2(n5680), .ZN(n6371) );
  INV_X1 U6282 ( .A(n7787), .ZN(n7350) );
  INV_X1 U6283 ( .A(n8334), .ZN(n6117) );
  INV_X1 U6284 ( .A(n6176), .ZN(n6161) );
  NAND2_X1 U6285 ( .A1(n6246), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n6263) );
  OR2_X1 U6286 ( .A1(n6036), .A2(n6038), .ZN(n6039) );
  INV_X1 U6287 ( .A(n6325), .ZN(n6287) );
  OR2_X1 U6288 ( .A1(n6263), .A2(n8368), .ZN(n6276) );
  OR2_X1 U6289 ( .A1(n6192), .A2(n8412), .ZN(n6208) );
  NOR2_X1 U6290 ( .A1(n8869), .A2(n8868), .ZN(n8870) );
  NAND2_X1 U6291 ( .A1(n6207), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n6233) );
  NOR2_X1 U6292 ( .A1(n7849), .A2(n7848), .ZN(n7850) );
  INV_X1 U6293 ( .A(n4453), .ZN(n8731) );
  OR2_X1 U6294 ( .A1(n4989), .A2(n4988), .ZN(n5206) );
  NAND2_X1 U6295 ( .A1(n4967), .A2(SI_12_), .ZN(n4968) );
  INV_X1 U6296 ( .A(SI_10_), .ZN(n10040) );
  NAND2_X1 U6297 ( .A1(n6431), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n4930) );
  INV_X1 U6298 ( .A(n7899), .ZN(n6374) );
  OR2_X1 U6299 ( .A1(n5484), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5494) );
  OR2_X1 U6300 ( .A1(n5894), .A2(n5884), .ZN(n7971) );
  OR2_X1 U6301 ( .A1(n5894), .A2(n5887), .ZN(n7984) );
  AND2_X1 U6302 ( .A1(n5663), .A2(n5662), .ZN(n7859) );
  NOR2_X1 U6303 ( .A1(n9721), .A2(n8064), .ZN(n8065) );
  OR2_X1 U6304 ( .A1(n5640), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n5652) );
  OR2_X1 U6305 ( .A1(n5597), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n5608) );
  NAND2_X1 U6306 ( .A1(n5545), .A2(n5544), .ZN(n5556) );
  INV_X1 U6307 ( .A(n7780), .ZN(n6992) );
  AND2_X1 U6308 ( .A1(n5772), .A2(n6602), .ZN(n6359) );
  INV_X1 U6309 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n5767) );
  AND2_X1 U6310 ( .A1(n7769), .A2(n7768), .ZN(n8132) );
  INV_X1 U6311 ( .A(n7711), .ZN(n7706) );
  INV_X1 U6312 ( .A(n7997), .ZN(n7348) );
  OR2_X1 U6313 ( .A1(n9771), .A2(n7817), .ZN(n9819) );
  AND2_X1 U6314 ( .A1(n8399), .A2(n6245), .ZN(n8341) );
  OR2_X1 U6315 ( .A1(n7601), .A2(n7597), .ZN(n6306) );
  NAND2_X1 U6316 ( .A1(n6346), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8458) );
  NAND2_X1 U6317 ( .A1(n5933), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5925) );
  OR2_X1 U6318 ( .A1(n9305), .A2(n8657), .ZN(n9460) );
  OR2_X1 U6319 ( .A1(n9305), .A2(n6694), .ZN(n9451) );
  AOI21_X1 U6320 ( .B1(n8920), .B2(n9489), .A(n8870), .ZN(n8871) );
  NAND2_X1 U6321 ( .A1(n8706), .A2(n8863), .ZN(n8878) );
  AND2_X1 U6322 ( .A1(n9103), .A2(n9591), .ZN(n9104) );
  INV_X1 U6323 ( .A(n9613), .ZN(n9591) );
  INV_X1 U6324 ( .A(n8491), .ZN(n9561) );
  AND2_X1 U6325 ( .A1(n6904), .A2(n8588), .ZN(n9516) );
  XNOR2_X1 U6326 ( .A(n4978), .B(n9926), .ZN(n5177) );
  INV_X1 U6327 ( .A(n5113), .ZN(n5114) );
  INV_X1 U6328 ( .A(SI_7_), .ZN(n10023) );
  INV_X1 U6329 ( .A(SI_8_), .ZN(n10092) );
  OAI21_X1 U6330 ( .B1(n6386), .B2(n7991), .A(n6385), .ZN(n6387) );
  AND2_X1 U6331 ( .A1(n5647), .A2(n5646), .ZN(n7904) );
  AND4_X1 U6332 ( .A1(n5344), .A2(n5343), .A3(n5342), .A4(n5341), .ZN(n7985)
         );
  OR2_X1 U6333 ( .A1(P2_U3150), .A2(n6418), .ZN(n9720) );
  INV_X1 U6334 ( .A(n7377), .ZN(n9770) );
  INV_X1 U6335 ( .A(n8212), .ZN(n8245) );
  OR2_X1 U6336 ( .A1(n7817), .A2(n7808), .ZN(n9807) );
  AND2_X1 U6337 ( .A1(n5451), .A2(n5467), .ZN(n7007) );
  AND4_X1 U6338 ( .A1(n6157), .A2(n6156), .A3(n6155), .A4(n6154), .ZN(n8383)
         );
  AND4_X1 U6339 ( .A1(n6140), .A2(n6139), .A3(n6138), .A4(n6137), .ZN(n8384)
         );
  INV_X1 U6340 ( .A(n9413), .ZN(n9454) );
  AND2_X1 U6341 ( .A1(n8511), .A2(n8509), .ZN(n8635) );
  AND2_X1 U6342 ( .A1(n9510), .A2(n4453), .ZN(n9480) );
  AND2_X1 U6343 ( .A1(n9510), .A2(n6910), .ZN(n9472) );
  NOR2_X1 U6344 ( .A1(n9105), .A2(n9104), .ZN(n9106) );
  INV_X1 U6345 ( .A(n9617), .ZN(n9538) );
  NAND2_X1 U6346 ( .A1(n9505), .A2(n9593), .ZN(n9617) );
  NAND2_X1 U6347 ( .A1(n5303), .A2(n5304), .ZN(n6883) );
  AND2_X1 U6348 ( .A1(n5154), .A2(n5153), .ZN(n9397) );
  XNOR2_X1 U6349 ( .A(n4950), .B(n10023), .ZN(n5092) );
  INV_X1 U6350 ( .A(n7954), .ZN(n7977) );
  INV_X1 U6351 ( .A(n7973), .ZN(n7991) );
  INV_X1 U6352 ( .A(n7904), .ZN(n8111) );
  INV_X1 U6353 ( .A(n9775), .ZN(n9777) );
  INV_X1 U6354 ( .A(n8223), .ZN(n8248) );
  NOR2_X1 U6355 ( .A1(n5766), .A2(n5768), .ZN(n5769) );
  OR2_X1 U6356 ( .A1(n9838), .A2(n9796), .ZN(n8320) );
  AND2_X1 U6357 ( .A1(n5765), .A2(n5764), .ZN(n9838) );
  INV_X1 U6358 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6478) );
  INV_X1 U6359 ( .A(n6560), .ZN(n6647) );
  NAND2_X1 U6360 ( .A1(n6332), .A2(n6331), .ZN(n8462) );
  INV_X1 U6361 ( .A(n8897), .ZN(n8939) );
  AND4_X1 U6362 ( .A1(n6197), .A2(n6196), .A3(n6195), .A4(n6194), .ZN(n9026)
         );
  INV_X1 U6363 ( .A(n7559), .ZN(n8747) );
  INV_X1 U6364 ( .A(n9431), .ZN(n9466) );
  INV_X1 U6365 ( .A(n9480), .ZN(n9085) );
  INV_X1 U6366 ( .A(n9482), .ZN(n9071) );
  INV_X1 U6367 ( .A(n8589), .ZN(n8658) );
  INV_X1 U6368 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n6480) );
  INV_X1 U6369 ( .A(n8005), .ZN(P2_U3893) );
  NAND2_X1 U6370 ( .A1(n5317), .A2(n4909), .ZN(P1_U3521) );
  OAI21_X2 U6371 ( .B1(n4352), .B2(n4922), .A(n4921), .ZN(n4927) );
  INV_X1 U6372 ( .A(SI_1_), .ZN(n4924) );
  NAND2_X1 U6373 ( .A1(n6436), .A2(SI_0_), .ZN(n5378) );
  INV_X1 U6374 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n4926) );
  AND2_X1 U6375 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n4925) );
  NAND2_X1 U6376 ( .A1(n4923), .A2(n4925), .ZN(n5039) );
  OAI21_X1 U6377 ( .B1(n5378), .B2(n4926), .A(n5039), .ZN(n5042) );
  NAND2_X1 U6378 ( .A1(n5041), .A2(n5042), .ZN(n4929) );
  NAND2_X1 U6379 ( .A1(n4927), .A2(SI_1_), .ZN(n4928) );
  NAND2_X1 U6380 ( .A1(n4929), .A2(n4928), .ZN(n5046) );
  INV_X1 U6381 ( .A(SI_2_), .ZN(n9903) );
  XNOR2_X1 U6382 ( .A(n4932), .B(n9903), .ZN(n5047) );
  NAND2_X1 U6383 ( .A1(n5046), .A2(n5047), .ZN(n4934) );
  NAND2_X1 U6384 ( .A1(n4932), .A2(SI_2_), .ZN(n4933) );
  NAND2_X1 U6385 ( .A1(n4934), .A2(n4933), .ZN(n5058) );
  MUX2_X1 U6386 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .S(n4923), .Z(n4936) );
  INV_X1 U6387 ( .A(SI_3_), .ZN(n4935) );
  XNOR2_X1 U6388 ( .A(n4936), .B(n4935), .ZN(n5057) );
  NAND2_X1 U6389 ( .A1(n5058), .A2(n5057), .ZN(n5069) );
  NAND2_X1 U6390 ( .A1(n4936), .A2(SI_3_), .ZN(n5068) );
  NAND2_X1 U6391 ( .A1(n4940), .A2(SI_4_), .ZN(n4938) );
  AND2_X1 U6392 ( .A1(n5068), .A2(n4938), .ZN(n4937) );
  NAND2_X1 U6393 ( .A1(n5069), .A2(n4937), .ZN(n4942) );
  INV_X1 U6394 ( .A(SI_4_), .ZN(n4939) );
  XNOR2_X1 U6395 ( .A(n4940), .B(n4939), .ZN(n5070) );
  MUX2_X1 U6396 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n4923), .Z(n4944) );
  INV_X1 U6397 ( .A(SI_5_), .ZN(n4943) );
  NAND2_X1 U6398 ( .A1(n4944), .A2(SI_5_), .ZN(n5084) );
  MUX2_X1 U6399 ( .A(n6438), .B(n6453), .S(n4352), .Z(n4947) );
  INV_X1 U6400 ( .A(n4947), .ZN(n4945) );
  NAND2_X1 U6401 ( .A1(n4945), .A2(SI_6_), .ZN(n4946) );
  INV_X1 U6402 ( .A(n4946), .ZN(n4948) );
  MUX2_X1 U6403 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n6431), .Z(n4950) );
  NAND2_X1 U6404 ( .A1(n4950), .A2(SI_7_), .ZN(n4951) );
  MUX2_X1 U6405 ( .A(n6460), .B(n6462), .S(n6431), .Z(n4952) );
  INV_X1 U6406 ( .A(n4952), .ZN(n4953) );
  NAND2_X1 U6407 ( .A1(n4953), .A2(SI_8_), .ZN(n4954) );
  MUX2_X1 U6408 ( .A(n6478), .B(n6480), .S(n6431), .Z(n4956) );
  INV_X1 U6409 ( .A(n4956), .ZN(n4957) );
  NAND2_X1 U6410 ( .A1(n4957), .A2(SI_9_), .ZN(n4958) );
  NAND2_X1 U6411 ( .A1(n5102), .A2(n4910), .ZN(n4960) );
  MUX2_X1 U6412 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .S(n4923), .Z(n4962) );
  MUX2_X1 U6413 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .S(n4923), .Z(n5120) );
  NAND2_X1 U6414 ( .A1(n5120), .A2(SI_11_), .ZN(n4963) );
  NAND2_X1 U6415 ( .A1(n4962), .A2(SI_10_), .ZN(n5118) );
  INV_X1 U6416 ( .A(n5120), .ZN(n4964) );
  INV_X1 U6417 ( .A(SI_11_), .ZN(n9932) );
  NAND2_X1 U6418 ( .A1(n4964), .A2(n9932), .ZN(n4965) );
  MUX2_X1 U6419 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .S(n4923), .Z(n4967) );
  MUX2_X1 U6420 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n6431), .Z(n5133) );
  MUX2_X1 U6421 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n4923), .Z(n5142) );
  INV_X1 U6422 ( .A(SI_14_), .ZN(n10026) );
  NAND2_X1 U6423 ( .A1(n4969), .A2(n10026), .ZN(n4970) );
  MUX2_X1 U6424 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .S(n4923), .Z(n5158) );
  NOR2_X1 U6425 ( .A1(n5158), .A2(SI_15_), .ZN(n5167) );
  MUX2_X1 U6426 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(P2_DATAO_REG_16__SCAN_IN), 
        .S(n4923), .Z(n5171) );
  INV_X1 U6427 ( .A(SI_16_), .ZN(n10069) );
  NOR2_X1 U6428 ( .A1(n5168), .A2(n4971), .ZN(n4977) );
  OR2_X1 U6429 ( .A1(n4972), .A2(n10069), .ZN(n4973) );
  NAND2_X1 U6430 ( .A1(n5158), .A2(SI_15_), .ZN(n5169) );
  MUX2_X1 U6431 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(P2_DATAO_REG_17__SCAN_IN), 
        .S(n6431), .Z(n4978) );
  INV_X1 U6432 ( .A(SI_17_), .ZN(n9926) );
  MUX2_X1 U6433 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n4923), .Z(n4980) );
  NAND2_X1 U6434 ( .A1(n4980), .A2(SI_18_), .ZN(n5196) );
  INV_X1 U6435 ( .A(n4980), .ZN(n4981) );
  INV_X1 U6436 ( .A(SI_18_), .ZN(n10052) );
  NAND2_X1 U6437 ( .A1(n4981), .A2(n10052), .ZN(n4982) );
  NAND2_X1 U6438 ( .A1(n5196), .A2(n4982), .ZN(n5185) );
  INV_X1 U6439 ( .A(n5185), .ZN(n5183) );
  MUX2_X1 U6440 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(P2_DATAO_REG_19__SCAN_IN), 
        .S(n6431), .Z(n4986) );
  INV_X1 U6441 ( .A(n4986), .ZN(n4984) );
  INV_X1 U6442 ( .A(SI_19_), .ZN(n4983) );
  NAND2_X1 U6443 ( .A1(n4984), .A2(n4983), .ZN(n4985) );
  INV_X1 U6444 ( .A(n4985), .ZN(n4989) );
  XNOR2_X1 U6445 ( .A(n4986), .B(SI_19_), .ZN(n5198) );
  INV_X1 U6446 ( .A(n5198), .ZN(n4987) );
  MUX2_X1 U6447 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(P2_DATAO_REG_20__SCAN_IN), 
        .S(n4923), .Z(n5208) );
  MUX2_X1 U6448 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(P2_DATAO_REG_21__SCAN_IN), 
        .S(n6431), .Z(n5213) );
  INV_X1 U6449 ( .A(SI_21_), .ZN(n10055) );
  NOR2_X1 U6450 ( .A1(n4993), .A2(n10055), .ZN(n4995) );
  NAND2_X1 U6451 ( .A1(n4993), .A2(n10055), .ZN(n4994) );
  MUX2_X1 U6452 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(P2_DATAO_REG_22__SCAN_IN), 
        .S(n6431), .Z(n4996) );
  INV_X1 U6453 ( .A(SI_22_), .ZN(n4997) );
  XNOR2_X1 U6454 ( .A(n4996), .B(n4997), .ZN(n5218) );
  NAND2_X1 U6455 ( .A1(n5219), .A2(n5218), .ZN(n5223) );
  INV_X1 U6456 ( .A(n4996), .ZN(n4998) );
  NAND2_X1 U6457 ( .A1(n4998), .A2(n4997), .ZN(n5222) );
  MUX2_X1 U6458 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(P2_DATAO_REG_23__SCAN_IN), 
        .S(n6431), .Z(n5002) );
  INV_X1 U6459 ( .A(n5002), .ZN(n4999) );
  INV_X1 U6460 ( .A(SI_23_), .ZN(n5001) );
  NAND2_X1 U6461 ( .A1(n4999), .A2(n5001), .ZN(n5000) );
  INV_X1 U6462 ( .A(n5000), .ZN(n5003) );
  XNOR2_X1 U6463 ( .A(n5002), .B(n5001), .ZN(n5224) );
  MUX2_X1 U6464 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(P2_DATAO_REG_24__SCAN_IN), 
        .S(n4923), .Z(n5005) );
  INV_X1 U6465 ( .A(SI_24_), .ZN(n9938) );
  XNOR2_X1 U6466 ( .A(n5005), .B(n9938), .ZN(n5228) );
  INV_X1 U6467 ( .A(n5005), .ZN(n5006) );
  MUX2_X1 U6468 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(P2_DATAO_REG_25__SCAN_IN), 
        .S(n4923), .Z(n5007) );
  INV_X1 U6469 ( .A(SI_25_), .ZN(n9944) );
  XNOR2_X1 U6470 ( .A(n5007), .B(n9944), .ZN(n5232) );
  INV_X1 U6471 ( .A(n5007), .ZN(n5008) );
  NAND2_X1 U6472 ( .A1(n5008), .A2(n9944), .ZN(n5009) );
  NAND2_X1 U6473 ( .A1(n5010), .A2(n5009), .ZN(n5237) );
  MUX2_X1 U6474 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(P2_DATAO_REG_26__SCAN_IN), 
        .S(n4923), .Z(n5011) );
  INV_X1 U6475 ( .A(SI_26_), .ZN(n9945) );
  XNOR2_X1 U6476 ( .A(n5011), .B(n9945), .ZN(n5236) );
  NAND2_X1 U6477 ( .A1(n5237), .A2(n5236), .ZN(n5014) );
  INV_X1 U6478 ( .A(n5011), .ZN(n5012) );
  NAND2_X1 U6479 ( .A1(n5012), .A2(n9945), .ZN(n5013) );
  NAND2_X1 U6480 ( .A1(n5014), .A2(n5013), .ZN(n5240) );
  MUX2_X1 U6481 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(P2_DATAO_REG_27__SCAN_IN), 
        .S(n6431), .Z(n5015) );
  INV_X1 U6482 ( .A(SI_27_), .ZN(n10025) );
  XNOR2_X1 U6483 ( .A(n5015), .B(n10025), .ZN(n5241) );
  NAND2_X1 U6484 ( .A1(n5240), .A2(n5241), .ZN(n5018) );
  INV_X1 U6485 ( .A(n5015), .ZN(n5016) );
  NAND2_X1 U6486 ( .A1(n5016), .A2(n10025), .ZN(n5017) );
  NAND2_X1 U6487 ( .A1(n5018), .A2(n5017), .ZN(n5245) );
  MUX2_X1 U6488 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(P2_DATAO_REG_28__SCAN_IN), 
        .S(n6431), .Z(n5019) );
  INV_X1 U6489 ( .A(SI_28_), .ZN(n10068) );
  XNOR2_X1 U6490 ( .A(n5019), .B(n10068), .ZN(n5244) );
  NAND2_X1 U6491 ( .A1(n5245), .A2(n5244), .ZN(n5022) );
  INV_X1 U6492 ( .A(n5019), .ZN(n5020) );
  NAND2_X1 U6493 ( .A1(n5020), .A2(n10068), .ZN(n5021) );
  INV_X1 U6494 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n5023) );
  INV_X1 U6495 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n9194) );
  MUX2_X1 U6496 ( .A(n5023), .B(n9194), .S(n6431), .Z(n5249) );
  NOR2_X1 U6497 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n5029) );
  NOR2_X1 U6498 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n5028) );
  NOR2_X1 U6499 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n5027) );
  NAND2_X1 U6500 ( .A1(n5033), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5291) );
  NAND2_X1 U6501 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_26__SCAN_IN), 
        .ZN(n5032) );
  XNOR2_X2 U6502 ( .A(n5034), .B(n5276), .ZN(n5286) );
  NAND2_X2 U6503 ( .A1(n5052), .A2(n6431), .ZN(n5188) );
  NAND2_X1 U6504 ( .A1(n5673), .A2(n5265), .ZN(n5036) );
  OR2_X1 U6505 ( .A1(n5267), .A2(n9194), .ZN(n5035) );
  INV_X1 U6506 ( .A(SI_0_), .ZN(n5038) );
  INV_X1 U6507 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5037) );
  OAI21_X1 U6508 ( .B1(n6436), .B2(n5038), .A(n5037), .ZN(n5040) );
  AND2_X1 U6509 ( .A1(n5040), .A2(n5039), .ZN(n9196) );
  MUX2_X1 U6510 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9196), .S(n5052), .Z(n9519) );
  INV_X1 U6511 ( .A(n9519), .ZN(n7029) );
  INV_X1 U6512 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6433) );
  XNOR2_X1 U6513 ( .A(n5041), .B(n5042), .ZN(n6454) );
  OR2_X1 U6514 ( .A1(n5188), .A2(n6454), .ZN(n5044) );
  NAND2_X1 U6515 ( .A1(n5103), .A2(n8763), .ZN(n5043) );
  INV_X1 U6516 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6435) );
  OR2_X1 U6517 ( .A1(n5267), .A2(n6435), .ZN(n5051) );
  XNOR2_X1 U6518 ( .A(n5047), .B(n5046), .ZN(n6456) );
  OR2_X1 U6519 ( .A1(n5188), .A2(n6456), .ZN(n5050) );
  OR2_X1 U6520 ( .A1(n5048), .A2(n5278), .ZN(n5063) );
  XNOR2_X1 U6521 ( .A(n5063), .B(P1_IR_REG_2__SCAN_IN), .ZN(n8777) );
  NAND2_X1 U6522 ( .A1(n5103), .A2(n8777), .ZN(n5049) );
  AND3_X2 U6523 ( .A1(n5051), .A2(n5050), .A3(n5049), .ZN(n9501) );
  INV_X1 U6524 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5053) );
  NAND2_X1 U6525 ( .A1(n5063), .A2(n5053), .ZN(n5054) );
  NAND2_X1 U6526 ( .A1(n5054), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5056) );
  INV_X1 U6527 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n5055) );
  XNOR2_X1 U6528 ( .A(n5056), .B(n5055), .ZN(n8776) );
  INV_X1 U6529 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6449) );
  XNOR2_X1 U6530 ( .A(n5058), .B(n5057), .ZN(n6457) );
  OR2_X1 U6531 ( .A1(n5188), .A2(n6457), .ZN(n5059) );
  OR2_X1 U6532 ( .A1(n5061), .A2(n5278), .ZN(n5062) );
  AND2_X1 U6533 ( .A1(n5063), .A2(n5062), .ZN(n5066) );
  INV_X1 U6534 ( .A(n5066), .ZN(n5064) );
  NAND2_X1 U6535 ( .A1(n5064), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n5067) );
  INV_X1 U6536 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5065) );
  NAND2_X1 U6537 ( .A1(n5066), .A2(n5065), .ZN(n5074) );
  INV_X1 U6538 ( .A(n9318), .ZN(n6447) );
  NAND2_X1 U6539 ( .A1(n5069), .A2(n5068), .ZN(n5071) );
  XNOR2_X1 U6540 ( .A(n5071), .B(n5070), .ZN(n6455) );
  OR2_X1 U6541 ( .A1(n5188), .A2(n6455), .ZN(n5073) );
  INV_X1 U6542 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6448) );
  NAND2_X1 U6543 ( .A1(n4369), .A2(n9541), .ZN(n6976) );
  NAND2_X1 U6544 ( .A1(n5074), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5075) );
  XNOR2_X1 U6545 ( .A(n5075), .B(P1_IR_REG_5__SCAN_IN), .ZN(n8823) );
  INV_X1 U6546 ( .A(n8823), .ZN(n9332) );
  INV_X1 U6547 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6451) );
  OR2_X1 U6548 ( .A1(n5267), .A2(n6451), .ZN(n5079) );
  XNOR2_X1 U6549 ( .A(n5076), .B(n5077), .ZN(n6450) );
  OR2_X1 U6550 ( .A1(n5188), .A2(n6450), .ZN(n5078) );
  OAI211_X1 U6551 ( .C1(n5052), .C2(n9332), .A(n5079), .B(n5078), .ZN(n7054)
         );
  NAND2_X1 U6552 ( .A1(n5080), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5081) );
  MUX2_X1 U6553 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5081), .S(
        P1_IR_REG_6__SCAN_IN), .Z(n5083) );
  AND2_X1 U6554 ( .A1(n5083), .A2(n5082), .ZN(n8825) );
  INV_X1 U6555 ( .A(n8825), .ZN(n9346) );
  NAND2_X1 U6556 ( .A1(n5085), .A2(n5084), .ZN(n5087) );
  XNOR2_X1 U6557 ( .A(n5087), .B(n5086), .ZN(n6452) );
  OR2_X1 U6558 ( .A1(n5188), .A2(n6452), .ZN(n5089) );
  OR2_X1 U6559 ( .A1(n5267), .A2(n6453), .ZN(n5088) );
  OAI211_X1 U6560 ( .C1(n5052), .C2(n9346), .A(n5089), .B(n5088), .ZN(n9473)
         );
  NAND2_X1 U6561 ( .A1(n5082), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5090) );
  XNOR2_X1 U6562 ( .A(n5090), .B(P1_IR_REG_7__SCAN_IN), .ZN(n8826) );
  INV_X1 U6563 ( .A(n8826), .ZN(n9243) );
  INV_X1 U6564 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n5091) );
  OR2_X1 U6565 ( .A1(n5267), .A2(n5091), .ZN(n5093) );
  NOR2_X1 U6566 ( .A1(n5094), .A2(n5278), .ZN(n5095) );
  NAND2_X1 U6567 ( .A1(n5095), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n5098) );
  INV_X1 U6568 ( .A(n5095), .ZN(n5097) );
  INV_X1 U6569 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n5096) );
  NAND2_X1 U6570 ( .A1(n5097), .A2(n5096), .ZN(n5104) );
  INV_X1 U6571 ( .A(n8828), .ZN(n9258) );
  XNOR2_X1 U6572 ( .A(n5099), .B(n4414), .ZN(n6461) );
  OR2_X1 U6573 ( .A1(n6461), .A2(n5188), .ZN(n5101) );
  OR2_X1 U6574 ( .A1(n5267), .A2(n6462), .ZN(n5100) );
  OAI211_X1 U6575 ( .C1(n5052), .C2(n9258), .A(n5101), .B(n5100), .ZN(n8486)
         );
  XNOR2_X1 U6576 ( .A(n5102), .B(n4910), .ZN(n6477) );
  NAND2_X1 U6577 ( .A1(n6477), .A2(n5265), .ZN(n5107) );
  NAND2_X1 U6578 ( .A1(n5104), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5105) );
  XNOR2_X1 U6579 ( .A(n5105), .B(P1_IR_REG_9__SCAN_IN), .ZN(n8829) );
  AOI22_X1 U6580 ( .A1(n5203), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n5103), .B2(
        n8829), .ZN(n5106) );
  NAND2_X1 U6581 ( .A1(n6481), .A2(n5265), .ZN(n5117) );
  NOR2_X1 U6582 ( .A1(n5110), .A2(n5278), .ZN(n5111) );
  MUX2_X1 U6583 ( .A(n5278), .B(n5111), .S(P1_IR_REG_10__SCAN_IN), .Z(n5112)
         );
  INV_X1 U6584 ( .A(n5112), .ZN(n5115) );
  AND2_X1 U6585 ( .A1(n5115), .A2(n5114), .ZN(n8830) );
  AOI22_X1 U6586 ( .A1(n5203), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n5103), .B2(
        n8830), .ZN(n5116) );
  NAND2_X1 U6587 ( .A1(n5119), .A2(n5118), .ZN(n5122) );
  XNOR2_X1 U6588 ( .A(n5120), .B(SI_11_), .ZN(n5121) );
  XNOR2_X1 U6589 ( .A(n5122), .B(n5121), .ZN(n6488) );
  NAND2_X1 U6590 ( .A1(n6488), .A2(n5265), .ZN(n5125) );
  OR2_X1 U6591 ( .A1(n5113), .A2(n5278), .ZN(n5123) );
  XNOR2_X1 U6592 ( .A(n5123), .B(P1_IR_REG_11__SCAN_IN), .ZN(n9351) );
  AOI22_X1 U6593 ( .A1(n5203), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n5103), .B2(
        n9351), .ZN(n5124) );
  NAND2_X1 U6594 ( .A1(n5127), .A2(n5126), .ZN(n5128) );
  NAND2_X1 U6595 ( .A1(n6511), .A2(n5265), .ZN(n5132) );
  INV_X1 U6596 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n5130) );
  NAND2_X1 U6597 ( .A1(n5113), .A2(n5130), .ZN(n5146) );
  NAND2_X1 U6598 ( .A1(n5146), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5137) );
  XNOR2_X1 U6599 ( .A(n5137), .B(P1_IR_REG_12__SCAN_IN), .ZN(n8832) );
  AOI22_X1 U6600 ( .A1(n5203), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n5103), .B2(
        n8832), .ZN(n5131) );
  XNOR2_X1 U6601 ( .A(n5133), .B(SI_13_), .ZN(n5134) );
  XNOR2_X1 U6602 ( .A(n5135), .B(n5134), .ZN(n6580) );
  NAND2_X1 U6603 ( .A1(n6580), .A2(n5265), .ZN(n5141) );
  INV_X1 U6604 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n5136) );
  NAND2_X1 U6605 ( .A1(n5137), .A2(n5136), .ZN(n5138) );
  NAND2_X1 U6606 ( .A1(n5138), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5139) );
  XNOR2_X1 U6607 ( .A(n5139), .B(P1_IR_REG_13__SCAN_IN), .ZN(n8833) );
  AOI22_X1 U6608 ( .A1(n5203), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n5103), .B2(
        n8833), .ZN(n5140) );
  XNOR2_X1 U6609 ( .A(n5142), .B(SI_14_), .ZN(n5143) );
  XNOR2_X1 U6610 ( .A(n5144), .B(n5143), .ZN(n6591) );
  NAND2_X1 U6611 ( .A1(n6591), .A2(n5265), .ZN(n5156) );
  INV_X1 U6612 ( .A(n5151), .ZN(n5145) );
  OAI21_X1 U6613 ( .B1(n5146), .B2(n5145), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n5147) );
  MUX2_X1 U6614 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5147), .S(
        P1_IR_REG_14__SCAN_IN), .Z(n5154) );
  NOR2_X1 U6615 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n5150) );
  NOR2_X1 U6616 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n5149) );
  NOR2_X1 U6617 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n5148) );
  NAND4_X1 U6618 ( .A1(n5151), .A2(n5150), .A3(n5149), .A4(n5148), .ZN(n5152)
         );
  INV_X1 U6619 ( .A(n4358), .ZN(n5153) );
  AOI22_X1 U6620 ( .A1(n5203), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n5103), .B2(
        n9397), .ZN(n5155) );
  INV_X1 U6621 ( .A(SI_15_), .ZN(n5157) );
  XNOR2_X1 U6622 ( .A(n5158), .B(n5157), .ZN(n5159) );
  XNOR2_X1 U6623 ( .A(n5168), .B(n5159), .ZN(n6633) );
  NAND2_X1 U6624 ( .A1(n6633), .A2(n5265), .ZN(n5166) );
  NOR2_X1 U6625 ( .A1(n4358), .A2(n5278), .ZN(n5160) );
  MUX2_X1 U6626 ( .A(n5278), .B(n5160), .S(P1_IR_REG_15__SCAN_IN), .Z(n5161)
         );
  INV_X1 U6627 ( .A(n5161), .ZN(n5164) );
  INV_X1 U6628 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n5162) );
  NAND2_X1 U6629 ( .A1(n5164), .A2(n5179), .ZN(n8836) );
  INV_X1 U6630 ( .A(n8836), .ZN(n9422) );
  AOI22_X1 U6631 ( .A1(n5203), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n5103), .B2(
        n9422), .ZN(n5165) );
  NAND2_X1 U6632 ( .A1(n5170), .A2(n5169), .ZN(n5173) );
  XNOR2_X1 U6633 ( .A(n5171), .B(SI_16_), .ZN(n5172) );
  NAND2_X1 U6634 ( .A1(n6720), .A2(n5265), .ZN(n5176) );
  NAND2_X1 U6635 ( .A1(n5179), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5174) );
  XNOR2_X1 U6636 ( .A(n5174), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9435) );
  AOI22_X1 U6637 ( .A1(n5203), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n5103), .B2(
        n9435), .ZN(n5175) );
  INV_X1 U6638 ( .A(n9083), .ZN(n9164) );
  NAND2_X1 U6639 ( .A1(n9079), .A2(n9164), .ZN(n9078) );
  XNOR2_X1 U6640 ( .A(n5178), .B(n5177), .ZN(n6706) );
  NAND2_X1 U6641 ( .A1(n6706), .A2(n5265), .ZN(n5181) );
  XNOR2_X1 U6642 ( .A(n5190), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9444) );
  AOI22_X1 U6643 ( .A1(n5203), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n5103), .B2(
        n9444), .ZN(n5180) );
  NAND2_X1 U6644 ( .A1(n5184), .A2(n5183), .ZN(n5197) );
  INV_X1 U6645 ( .A(n5184), .ZN(n5186) );
  NAND2_X1 U6646 ( .A1(n5186), .A2(n5185), .ZN(n5187) );
  NAND2_X1 U6647 ( .A1(n5197), .A2(n5187), .ZN(n6764) );
  OR2_X1 U6648 ( .A1(n6764), .A2(n5188), .ZN(n5195) );
  INV_X1 U6649 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5189) );
  INV_X1 U6650 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n5191) );
  NAND2_X1 U6651 ( .A1(n5192), .A2(n5191), .ZN(n5200) );
  OR2_X1 U6652 ( .A1(n5192), .A2(n5191), .ZN(n5193) );
  AND2_X1 U6653 ( .A1(n5200), .A2(n5193), .ZN(n8842) );
  AOI22_X1 U6654 ( .A1(n5203), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n5103), .B2(
        n8842), .ZN(n5194) );
  NAND2_X1 U6655 ( .A1(n5197), .A2(n5196), .ZN(n5199) );
  NAND2_X1 U6656 ( .A1(n6848), .A2(n5265), .ZN(n5205) );
  INV_X1 U6657 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5201) );
  AOI22_X1 U6658 ( .A1(n5203), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n5103), .B2(
        n8731), .ZN(n5204) );
  AND2_X1 U6659 ( .A1(n5207), .A2(n5206), .ZN(n5210) );
  XNOR2_X1 U6660 ( .A(n5208), .B(n9904), .ZN(n5209) );
  NAND2_X1 U6661 ( .A1(n6832), .A2(n5265), .ZN(n5212) );
  INV_X1 U6662 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n6852) );
  OR2_X1 U6663 ( .A1(n5267), .A2(n6852), .ZN(n5211) );
  XNOR2_X1 U6664 ( .A(n5213), .B(SI_21_), .ZN(n5214) );
  XNOR2_X1 U6665 ( .A(n5215), .B(n5214), .ZN(n6855) );
  NAND2_X1 U6666 ( .A1(n6855), .A2(n5265), .ZN(n5217) );
  INV_X1 U6667 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n6915) );
  OR2_X1 U6668 ( .A1(n5267), .A2(n6915), .ZN(n5216) );
  XNOR2_X1 U6669 ( .A(n5219), .B(n5218), .ZN(n7060) );
  NAND2_X1 U6670 ( .A1(n7060), .A2(n5265), .ZN(n5221) );
  INV_X1 U6671 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7063) );
  OR2_X1 U6672 ( .A1(n5267), .A2(n7063), .ZN(n5220) );
  NAND2_X1 U6673 ( .A1(n5223), .A2(n5222), .ZN(n5225) );
  NAND2_X1 U6674 ( .A1(n7076), .A2(n5265), .ZN(n5227) );
  INV_X1 U6675 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n7078) );
  OR2_X1 U6676 ( .A1(n5267), .A2(n7078), .ZN(n5226) );
  NAND2_X1 U6677 ( .A1(n7117), .A2(n5265), .ZN(n5231) );
  INV_X1 U6678 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7146) );
  OR2_X1 U6679 ( .A1(n5267), .A2(n7146), .ZN(n5230) );
  XNOR2_X1 U6680 ( .A(n5233), .B(n5232), .ZN(n7227) );
  NAND2_X1 U6681 ( .A1(n7227), .A2(n5265), .ZN(n5235) );
  INV_X1 U6682 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7246) );
  OR2_X1 U6683 ( .A1(n5267), .A2(n7246), .ZN(n5234) );
  XNOR2_X1 U6684 ( .A(n5237), .B(n5236), .ZN(n7258) );
  NAND2_X1 U6685 ( .A1(n7258), .A2(n5265), .ZN(n5239) );
  INV_X1 U6686 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n7334) );
  OR2_X1 U6687 ( .A1(n5267), .A2(n7334), .ZN(n5238) );
  NOR2_X4 U6688 ( .A1(n8931), .A2(n9114), .ZN(n8930) );
  XNOR2_X1 U6689 ( .A(n5240), .B(n5241), .ZN(n7356) );
  NAND2_X1 U6690 ( .A1(n7356), .A2(n5265), .ZN(n5243) );
  INV_X1 U6691 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n7822) );
  OR2_X1 U6692 ( .A1(n5267), .A2(n7822), .ZN(n5242) );
  XNOR2_X1 U6693 ( .A(n5245), .B(n5244), .ZN(n7395) );
  NAND2_X1 U6694 ( .A1(n7395), .A2(n5265), .ZN(n5247) );
  INV_X1 U6695 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n7440) );
  OR2_X1 U6696 ( .A1(n5267), .A2(n7440), .ZN(n5246) );
  INV_X1 U6697 ( .A(SI_29_), .ZN(n10043) );
  INV_X1 U6698 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n7857) );
  INV_X1 U6699 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n5253) );
  MUX2_X1 U6700 ( .A(n7857), .B(n5253), .S(n6436), .Z(n5254) );
  NAND2_X1 U6701 ( .A1(n5254), .A2(n10027), .ZN(n5259) );
  INV_X1 U6702 ( .A(n5254), .ZN(n5255) );
  NAND2_X1 U6703 ( .A1(n5255), .A2(SI_30_), .ZN(n5256) );
  NAND2_X1 U6704 ( .A1(n5259), .A2(n5256), .ZN(n5260) );
  NAND2_X1 U6705 ( .A1(n7855), .A2(n5265), .ZN(n5258) );
  OR2_X1 U6706 ( .A1(n5267), .A2(n7857), .ZN(n5257) );
  NOR2_X2 U6707 ( .A1(n8886), .A2(n8856), .ZN(n8855) );
  MUX2_X1 U6708 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n6436), .Z(n5262) );
  INV_X1 U6709 ( .A(SI_31_), .ZN(n10056) );
  XNOR2_X1 U6710 ( .A(n5262), .B(n10056), .ZN(n5263) );
  NAND2_X1 U6711 ( .A1(n8322), .A2(n5265), .ZN(n5269) );
  INV_X1 U6712 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n5266) );
  OR2_X1 U6713 ( .A1(n5267), .A2(n5266), .ZN(n5268) );
  XNOR2_X1 U6714 ( .A(n8855), .B(n8587), .ZN(n5275) );
  INV_X1 U6715 ( .A(n5270), .ZN(n5271) );
  NAND2_X1 U6716 ( .A1(n5271), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5297) );
  NAND2_X1 U6717 ( .A1(n4409), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5272) );
  NAND2_X1 U6718 ( .A1(n8658), .A2(n8738), .ZN(n9513) );
  NAND2_X1 U6719 ( .A1(n5273), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5274) );
  INV_X1 U6720 ( .A(n6854), .ZN(n8730) );
  NAND2_X1 U6721 ( .A1(n5275), .A2(n9496), .ZN(n8854) );
  INV_X1 U6722 ( .A(n8587), .ZN(n8851) );
  INV_X1 U6723 ( .A(n6892), .ZN(n8722) );
  NAND2_X1 U6724 ( .A1(n5277), .A2(n5276), .ZN(n5280) );
  NOR2_X2 U6725 ( .A1(n5280), .A2(P1_IR_REG_29__SCAN_IN), .ZN(n9185) );
  INV_X1 U6726 ( .A(n5902), .ZN(n5282) );
  NOR2_X2 U6727 ( .A1(n5903), .A2(n5282), .ZN(n5933) );
  NAND2_X1 U6728 ( .A1(n8578), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n5285) );
  NAND2_X1 U6729 ( .A1(n5959), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n5284) );
  NAND2_X1 U6730 ( .A1(n4360), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n5283) );
  INV_X1 U6731 ( .A(n5286), .ZN(n8657) );
  INV_X1 U6732 ( .A(n5287), .ZN(n9302) );
  NAND2_X1 U6733 ( .A1(n9302), .A2(P1_B_REG_SCAN_IN), .ZN(n5288) );
  NAND2_X1 U6734 ( .A1(n9490), .A2(n5288), .ZN(n8868) );
  OR2_X1 U6735 ( .A1(n8619), .A2(n8868), .ZN(n9093) );
  INV_X1 U6736 ( .A(n5289), .ZN(n5290) );
  NAND2_X1 U6737 ( .A1(n4410), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5292) );
  XNOR2_X1 U6738 ( .A(n5292), .B(P1_IR_REG_25__SCAN_IN), .ZN(n5301) );
  NAND2_X1 U6739 ( .A1(n5293), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5294) );
  XNOR2_X1 U6740 ( .A(n5294), .B(P1_IR_REG_24__SCAN_IN), .ZN(n5315) );
  INV_X1 U6741 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5296) );
  NAND2_X1 U6742 ( .A1(n5297), .A2(n5296), .ZN(n5298) );
  NAND2_X1 U6743 ( .A1(n5298), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5300) );
  INV_X1 U6744 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n5299) );
  XNOR2_X1 U6745 ( .A(n5300), .B(n5299), .ZN(n6486) );
  AND2_X1 U6746 ( .A1(n8622), .A2(n6892), .ZN(n6345) );
  NOR2_X1 U6747 ( .A1(n8660), .A2(n6345), .ZN(n6629) );
  INV_X1 U6748 ( .A(n5301), .ZN(n7248) );
  NAND2_X1 U6749 ( .A1(n7248), .A2(P1_B_REG_SCAN_IN), .ZN(n5302) );
  MUX2_X1 U6750 ( .A(n5302), .B(P1_B_REG_SCAN_IN), .S(n5315), .Z(n5303) );
  INV_X1 U6751 ( .A(n5304), .ZN(n7336) );
  NAND2_X1 U6752 ( .A1(n7336), .A2(n7248), .ZN(n9183) );
  OAI21_X1 U6753 ( .B1(n6883), .B2(P1_D_REG_1__SCAN_IN), .A(n9183), .ZN(n6328)
         );
  INV_X1 U6754 ( .A(n6883), .ZN(n5314) );
  NOR4_X1 U6755 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n5313) );
  NOR4_X1 U6756 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n5312) );
  OR4_X1 U6757 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n5310) );
  NOR4_X1 U6758 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n5308) );
  NOR4_X1 U6759 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n5307) );
  NOR4_X1 U6760 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n5306) );
  NOR4_X1 U6761 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n5305) );
  NAND4_X1 U6762 ( .A1(n5308), .A2(n5307), .A3(n5306), .A4(n5305), .ZN(n5309)
         );
  NOR4_X1 U6763 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        n5310), .A4(n5309), .ZN(n5311) );
  NAND3_X1 U6764 ( .A1(n5313), .A2(n5312), .A3(n5311), .ZN(n6885) );
  NAND2_X1 U6765 ( .A1(n5314), .A2(n6885), .ZN(n6329) );
  NAND2_X1 U6766 ( .A1(n9565), .A2(n8738), .ZN(n6343) );
  NAND4_X1 U6767 ( .A1(n6629), .A2(n6328), .A3(n6329), .A4(n6343), .ZN(n9090)
         );
  INV_X1 U6768 ( .A(n5315), .ZN(n7148) );
  NAND2_X1 U6769 ( .A1(n7336), .A2(n7148), .ZN(n9184) );
  OAI21_X1 U6770 ( .B1(n6883), .B2(P1_D_REG_0__SCAN_IN), .A(n9184), .ZN(n9089)
         );
  INV_X1 U6771 ( .A(n9089), .ZN(n6330) );
  INV_X2 U6772 ( .A(n9618), .ZN(n9546) );
  INV_X1 U6773 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n5316) );
  NOR2_X1 U6774 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n5323) );
  INV_X1 U6775 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5325) );
  INV_X1 U6776 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n5326) );
  INV_X1 U6777 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5328) );
  NAND2_X1 U6778 ( .A1(n5331), .A2(n5328), .ZN(n8323) );
  INV_X1 U6779 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n5330) );
  INV_X1 U6780 ( .A(n7495), .ZN(n5333) );
  AND2_X2 U6781 ( .A1(n5334), .A2(n5333), .ZN(n5416) );
  NAND2_X1 U6782 ( .A1(n5677), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n5344) );
  NAND2_X1 U6783 ( .A1(n5398), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n5343) );
  INV_X2 U6784 ( .A(n5399), .ZN(n5676) );
  NAND2_X1 U6785 ( .A1(n5400), .A2(n10058), .ZN(n5428) );
  INV_X1 U6786 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n5337) );
  INV_X1 U6787 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n10066) );
  INV_X1 U6788 ( .A(n5545), .ZN(n5546) );
  INV_X1 U6789 ( .A(n5338), .ZN(n5533) );
  NAND2_X1 U6790 ( .A1(n5533), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5339) );
  NAND2_X1 U6791 ( .A1(n5546), .A2(n5339), .ZN(n7915) );
  NAND2_X1 U6792 ( .A1(n5676), .A2(n7915), .ZN(n5342) );
  NAND2_X1 U6793 ( .A1(n5599), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n5341) );
  INV_X1 U6794 ( .A(n7985), .ZN(n8202) );
  INV_X1 U6795 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5346) );
  XNOR2_X2 U6796 ( .A(n5347), .B(n5346), .ZN(n5693) );
  MUX2_X1 U6797 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5349), .S(
        P2_IR_REG_27__SCAN_IN), .Z(n5350) );
  NAND2_X2 U6798 ( .A1(n5345), .A2(n5350), .ZN(n8057) );
  NAND2_X1 U6799 ( .A1(n6720), .A2(n7751), .ZN(n5355) );
  INV_X4 U6800 ( .A(n5379), .ZN(n5407) );
  OR2_X1 U6801 ( .A1(n5489), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n5503) );
  INV_X1 U6802 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5525) );
  INV_X1 U6803 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5513) );
  INV_X1 U6804 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n5351) );
  NAND3_X1 U6805 ( .A1(n5525), .A2(n5513), .A3(n5351), .ZN(n5352) );
  NOR2_X1 U6806 ( .A1(n5503), .A2(n5352), .ZN(n5539) );
  OR2_X1 U6807 ( .A1(n5539), .A2(n5330), .ZN(n5353) );
  XNOR2_X1 U6808 ( .A(n5353), .B(P2_IR_REG_16__SCAN_IN), .ZN(n8040) );
  AOI22_X1 U6809 ( .A1(n7752), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n5407), .B2(
        n8040), .ZN(n5354) );
  NAND2_X1 U6810 ( .A1(n6488), .A2(n7751), .ZN(n5360) );
  NAND2_X1 U6811 ( .A1(n5393), .A2(n4775), .ZN(n5411) );
  INV_X1 U6812 ( .A(n5356), .ZN(n5357) );
  OR2_X1 U6813 ( .A1(n5411), .A2(n5357), .ZN(n5478) );
  OAI21_X1 U6814 ( .B1(n5478), .B2(P2_IR_REG_10__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5358) );
  XNOR2_X1 U6815 ( .A(n5358), .B(P2_IR_REG_11__SCAN_IN), .ZN(n7418) );
  AOI22_X1 U6816 ( .A1(n7752), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n5407), .B2(
        n7418), .ZN(n5359) );
  NAND2_X1 U6817 ( .A1(n5360), .A2(n5359), .ZN(n9825) );
  NAND2_X1 U6818 ( .A1(n5677), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n5365) );
  NAND2_X1 U6819 ( .A1(n5599), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n5364) );
  INV_X2 U6820 ( .A(n5399), .ZN(n5642) );
  NAND2_X1 U6821 ( .A1(n5484), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5361) );
  NAND2_X1 U6822 ( .A1(n5494), .A2(n5361), .ZN(n7391) );
  NAND2_X1 U6823 ( .A1(n5642), .A2(n7391), .ZN(n5363) );
  NAND2_X1 U6824 ( .A1(n5398), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5362) );
  INV_X1 U6825 ( .A(n7451), .ZN(n7999) );
  NAND2_X1 U6826 ( .A1(n5426), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n5368) );
  NAND2_X1 U6827 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5366) );
  NAND2_X1 U6828 ( .A1(n5407), .A2(n6421), .ZN(n5367) );
  OAI211_X2 U6829 ( .C1(n5552), .C2(n6454), .A(n5368), .B(n5367), .ZN(n6669)
         );
  NAND2_X1 U6830 ( .A1(n5599), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5372) );
  NAND2_X1 U6831 ( .A1(n5398), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n5371) );
  NAND2_X1 U6832 ( .A1(n5416), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n5370) );
  NAND2_X1 U6833 ( .A1(n5335), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n5369) );
  NAND4_X2 U6834 ( .A1(n5372), .A2(n5371), .A3(n5370), .A4(n5369), .ZN(n5373)
         );
  INV_X2 U6835 ( .A(n5373), .ZN(n9763) );
  NAND2_X1 U6836 ( .A1(n9779), .A2(n5373), .ZN(n7617) );
  NAND2_X1 U6837 ( .A1(n5398), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5377) );
  NAND2_X1 U6838 ( .A1(n5416), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5376) );
  NAND2_X1 U6839 ( .A1(n5676), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n5375) );
  NAND2_X1 U6840 ( .A1(n5599), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5374) );
  AND4_X1 U6841 ( .A1(n5377), .A2(n5376), .A3(n5375), .A4(n5374), .ZN(n6545)
         );
  XNOR2_X1 U6842 ( .A(n5378), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n8330) );
  MUX2_X1 U6843 ( .A(P2_IR_REG_0__SCAN_IN), .B(n8330), .S(n5379), .Z(n6598) );
  INV_X1 U6844 ( .A(n6598), .ZN(n6614) );
  OR2_X1 U6845 ( .A1(n6545), .A2(n6614), .ZN(n6667) );
  NAND2_X1 U6846 ( .A1(n6661), .A2(n6667), .ZN(n6666) );
  NAND2_X1 U6847 ( .A1(n9763), .A2(n9779), .ZN(n5380) );
  NAND2_X1 U6848 ( .A1(n6666), .A2(n5380), .ZN(n9758) );
  NAND2_X1 U6849 ( .A1(n5416), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n5384) );
  NAND2_X1 U6850 ( .A1(n5599), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5383) );
  NAND2_X1 U6851 ( .A1(n5676), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n5382) );
  NAND2_X1 U6852 ( .A1(n5398), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5381) );
  NAND2_X1 U6853 ( .A1(n5426), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n5388) );
  NAND2_X1 U6854 ( .A1(n5407), .A2(n6535), .ZN(n5387) );
  OAI211_X1 U6855 ( .C1(n5552), .C2(n6456), .A(n5388), .B(n5387), .ZN(n5780)
         );
  INV_X1 U6856 ( .A(n7619), .ZN(n9759) );
  INV_X1 U6857 ( .A(n9745), .ZN(n5781) );
  INV_X1 U6858 ( .A(n5780), .ZN(n9769) );
  NAND2_X1 U6859 ( .A1(n5781), .A2(n9769), .ZN(n9741) );
  NAND2_X1 U6860 ( .A1(n5398), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5392) );
  NAND2_X1 U6861 ( .A1(n5677), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n5391) );
  INV_X1 U6862 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n9752) );
  NAND2_X1 U6863 ( .A1(n5642), .A2(n9752), .ZN(n5390) );
  NAND2_X1 U6864 ( .A1(n5599), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5389) );
  AND4_X2 U6865 ( .A1(n5392), .A2(n5391), .A3(n5390), .A4(n5389), .ZN(n9761)
         );
  NAND2_X1 U6866 ( .A1(n5426), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n5395) );
  NAND2_X1 U6867 ( .A1(n5407), .A2(n6560), .ZN(n5394) );
  OAI211_X1 U6868 ( .C1(n5552), .C2(n6457), .A(n5395), .B(n5394), .ZN(n9789)
         );
  INV_X1 U6869 ( .A(n9789), .ZN(n7622) );
  NAND2_X1 U6870 ( .A1(n9761), .A2(n7622), .ZN(n5396) );
  AND2_X1 U6871 ( .A1(n9741), .A2(n5396), .ZN(n5397) );
  NAND2_X1 U6872 ( .A1(n9757), .A2(n5397), .ZN(n6835) );
  OR2_X1 U6873 ( .A1(n9761), .A2(n7622), .ZN(n6789) );
  NAND2_X1 U6874 ( .A1(n5398), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n5405) );
  NAND2_X1 U6875 ( .A1(n5416), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5404) );
  INV_X1 U6876 ( .A(n5400), .ZN(n5417) );
  NAND2_X1 U6877 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n5401) );
  NAND2_X1 U6878 ( .A1(n5417), .A2(n5401), .ZN(n6794) );
  NAND2_X1 U6879 ( .A1(n5642), .A2(n6794), .ZN(n5403) );
  NAND2_X1 U6880 ( .A1(n5599), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5402) );
  NAND2_X1 U6881 ( .A1(n5426), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n5409) );
  NAND2_X1 U6882 ( .A1(n5411), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5406) );
  XNOR2_X1 U6883 ( .A(n5406), .B(P2_IR_REG_4__SCAN_IN), .ZN(n6742) );
  NAND2_X1 U6884 ( .A1(n5407), .A2(n6742), .ZN(n5408) );
  OAI211_X1 U6885 ( .C1(n5552), .C2(n6455), .A(n5409), .B(n5408), .ZN(n6795)
         );
  INV_X1 U6886 ( .A(n6795), .ZN(n9795) );
  NAND2_X1 U6887 ( .A1(n9747), .A2(n9795), .ZN(n7640) );
  NAND2_X1 U6888 ( .A1(n6872), .A2(n6795), .ZN(n7632) );
  INV_X1 U6889 ( .A(n6450), .ZN(n5410) );
  NAND2_X1 U6890 ( .A1(n7752), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n5414) );
  NAND2_X1 U6891 ( .A1(n5422), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5412) );
  XNOR2_X1 U6892 ( .A(n5412), .B(P2_IR_REG_5__SCAN_IN), .ZN(n6753) );
  NAND2_X1 U6893 ( .A1(n5407), .A2(n6753), .ZN(n5413) );
  NAND2_X1 U6894 ( .A1(n5398), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5421) );
  NAND2_X1 U6895 ( .A1(n5677), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n5420) );
  XNOR2_X1 U6896 ( .A(n5417), .B(P2_REG3_REG_5__SCAN_IN), .ZN(n6876) );
  NAND2_X1 U6897 ( .A1(n5642), .A2(n6876), .ZN(n5419) );
  NAND2_X1 U6898 ( .A1(n5599), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n5418) );
  NAND2_X1 U6899 ( .A1(n6879), .A2(n8003), .ZN(n6837) );
  INV_X1 U6900 ( .A(n5422), .ZN(n5424) );
  INV_X1 U6901 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5423) );
  NAND2_X1 U6902 ( .A1(n5424), .A2(n5423), .ZN(n5446) );
  NAND2_X1 U6903 ( .A1(n5446), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5425) );
  OR2_X1 U6904 ( .A1(n5552), .A2(n6452), .ZN(n5427) );
  NAND2_X1 U6905 ( .A1(n5398), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5433) );
  NAND2_X1 U6906 ( .A1(n5677), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n5432) );
  NAND2_X1 U6907 ( .A1(n5428), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5429) );
  NAND2_X1 U6908 ( .A1(n5440), .A2(n5429), .ZN(n6843) );
  NAND2_X1 U6909 ( .A1(n5642), .A2(n6843), .ZN(n5431) );
  NAND2_X1 U6910 ( .A1(n5599), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5430) );
  AND2_X1 U6911 ( .A1(n6837), .A2(n5435), .ZN(n5436) );
  NAND2_X1 U6912 ( .A1(n7091), .A2(n6860), .ZN(n5438) );
  NAND2_X1 U6913 ( .A1(n6872), .A2(n9795), .ZN(n6869) );
  NAND2_X1 U6914 ( .A1(n5398), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5445) );
  NAND2_X1 U6915 ( .A1(n5677), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n5444) );
  INV_X1 U6916 ( .A(n5439), .ZN(n5457) );
  NAND2_X1 U6917 ( .A1(n5440), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5441) );
  NAND2_X1 U6918 ( .A1(n5457), .A2(n5441), .ZN(n7097) );
  NAND2_X1 U6919 ( .A1(n5642), .A2(n7097), .ZN(n5443) );
  NAND2_X1 U6920 ( .A1(n5599), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n5442) );
  OR2_X1 U6921 ( .A1(n6459), .A2(n5552), .ZN(n5453) );
  INV_X1 U6922 ( .A(n5446), .ZN(n5448) );
  NAND2_X1 U6923 ( .A1(n5448), .A2(n5447), .ZN(n5450) );
  NAND2_X1 U6924 ( .A1(n5450), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5449) );
  MUX2_X1 U6925 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5449), .S(
        P2_IR_REG_7__SCAN_IN), .Z(n5451) );
  AOI22_X1 U6926 ( .A1(n7752), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n5407), .B2(
        n7007), .ZN(n5452) );
  NAND2_X1 U6927 ( .A1(n5453), .A2(n5452), .ZN(n7101) );
  NAND2_X1 U6928 ( .A1(n6986), .A2(n7101), .ZN(n7653) );
  INV_X1 U6929 ( .A(n7101), .ZN(n9808) );
  NAND2_X1 U6930 ( .A1(n9808), .A2(n6783), .ZN(n6991) );
  INV_X1 U6931 ( .A(n7779), .ZN(n5455) );
  AND2_X1 U6932 ( .A1(n6986), .A2(n9808), .ZN(n5454) );
  NAND2_X1 U6933 ( .A1(n5398), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n5462) );
  NAND2_X1 U6934 ( .A1(n5677), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n5461) );
  INV_X1 U6935 ( .A(n5456), .ZN(n5471) );
  NAND2_X1 U6936 ( .A1(n5457), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5458) );
  NAND2_X1 U6937 ( .A1(n5471), .A2(n5458), .ZN(n6994) );
  NAND2_X1 U6938 ( .A1(n5676), .A2(n6994), .ZN(n5460) );
  NAND2_X1 U6939 ( .A1(n5599), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5459) );
  OR2_X1 U6940 ( .A1(n6461), .A2(n5552), .ZN(n5465) );
  NAND2_X1 U6941 ( .A1(n5467), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5463) );
  XNOR2_X1 U6942 ( .A(n5463), .B(P2_IR_REG_8__SCAN_IN), .ZN(n7023) );
  AOI22_X1 U6943 ( .A1(n7752), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n5407), .B2(
        n7023), .ZN(n5464) );
  NAND2_X1 U6944 ( .A1(n5465), .A2(n5464), .ZN(n9814) );
  OR2_X1 U6945 ( .A1(n7090), .A2(n9814), .ZN(n7648) );
  NAND2_X1 U6946 ( .A1(n9814), .A2(n7090), .ZN(n7654) );
  AND2_X1 U6947 ( .A1(n7648), .A2(n7654), .ZN(n7780) );
  NAND2_X1 U6948 ( .A1(n6985), .A2(n6992), .ZN(n6984) );
  INV_X1 U6949 ( .A(n7090), .ZN(n8002) );
  NAND2_X1 U6950 ( .A1(n8002), .A2(n9814), .ZN(n5466) );
  NAND2_X1 U6951 ( .A1(n6477), .A2(n7751), .ZN(n5470) );
  OAI21_X1 U6952 ( .B1(n5467), .B2(P2_IR_REG_8__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5468) );
  XNOR2_X1 U6953 ( .A(n5468), .B(P2_IR_REG_9__SCAN_IN), .ZN(n7289) );
  AOI22_X1 U6954 ( .A1(n7752), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n5407), .B2(
        n7289), .ZN(n5469) );
  NAND2_X1 U6955 ( .A1(n5470), .A2(n5469), .ZN(n9823) );
  NAND2_X1 U6956 ( .A1(n5398), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5476) );
  NAND2_X1 U6957 ( .A1(n5677), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n5475) );
  NAND2_X1 U6958 ( .A1(n5471), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n5472) );
  NAND2_X1 U6959 ( .A1(n5482), .A2(n5472), .ZN(n7196) );
  NAND2_X1 U6960 ( .A1(n5642), .A2(n7196), .ZN(n5474) );
  NAND2_X1 U6961 ( .A1(n5599), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n5473) );
  NAND2_X1 U6962 ( .A1(n9823), .A2(n7282), .ZN(n7657) );
  NAND2_X1 U6963 ( .A1(n7649), .A2(n7657), .ZN(n7783) );
  INV_X1 U6964 ( .A(n7282), .ZN(n8001) );
  OR2_X1 U6965 ( .A1(n9823), .A2(n8001), .ZN(n5477) );
  NAND2_X1 U6966 ( .A1(n6481), .A2(n7751), .ZN(n5481) );
  NAND2_X1 U6967 ( .A1(n5478), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5479) );
  XNOR2_X1 U6968 ( .A(n5479), .B(P2_IR_REG_10__SCAN_IN), .ZN(n7320) );
  AOI22_X1 U6969 ( .A1(n7752), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n5407), .B2(
        n7320), .ZN(n5480) );
  NAND2_X1 U6970 ( .A1(n5481), .A2(n5480), .ZN(n7284) );
  NAND2_X1 U6971 ( .A1(n5398), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5488) );
  NAND2_X1 U6972 ( .A1(n5677), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n5487) );
  NAND2_X1 U6973 ( .A1(n5482), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5483) );
  NAND2_X1 U6974 ( .A1(n5484), .A2(n5483), .ZN(n7279) );
  NAND2_X1 U6975 ( .A1(n5642), .A2(n7279), .ZN(n5486) );
  NAND2_X1 U6976 ( .A1(n5599), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n5485) );
  OR2_X1 U6977 ( .A1(n7284), .A2(n7389), .ZN(n7668) );
  NAND2_X1 U6978 ( .A1(n7284), .A2(n7389), .ZN(n7671) );
  NAND2_X1 U6979 ( .A1(n7668), .A2(n7671), .ZN(n7784) );
  INV_X1 U6980 ( .A(n7389), .ZN(n8000) );
  INV_X1 U6981 ( .A(n9825), .ZN(n7394) );
  NAND2_X1 U6982 ( .A1(n6511), .A2(n7751), .ZN(n5492) );
  NAND2_X1 U6983 ( .A1(n5489), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5490) );
  XNOR2_X1 U6984 ( .A(n5490), .B(P2_IR_REG_12__SCAN_IN), .ZN(n7425) );
  AOI22_X1 U6985 ( .A1(n7752), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n5407), .B2(
        n7425), .ZN(n5491) );
  NAND2_X1 U6986 ( .A1(n5398), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5499) );
  NAND2_X1 U6987 ( .A1(n5677), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n5498) );
  INV_X1 U6988 ( .A(n5493), .ZN(n5506) );
  NAND2_X1 U6989 ( .A1(n5494), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5495) );
  NAND2_X1 U6990 ( .A1(n5506), .A2(n5495), .ZN(n7453) );
  NAND2_X1 U6991 ( .A1(n5642), .A2(n7453), .ZN(n5497) );
  NAND2_X1 U6992 ( .A1(n5599), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n5496) );
  NAND4_X1 U6993 ( .A1(n5499), .A2(n5498), .A3(n5497), .A4(n5496), .ZN(n7998)
         );
  XNOR2_X1 U6994 ( .A(n9834), .B(n7998), .ZN(n7787) );
  AOI21_X1 U6995 ( .B1(n7346), .B2(n7350), .A(n5502), .ZN(n7374) );
  NAND2_X1 U6996 ( .A1(n6580), .A2(n7751), .ZN(n5505) );
  NAND2_X1 U6997 ( .A1(n5503), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5514) );
  XNOR2_X1 U6998 ( .A(n5514), .B(P2_IR_REG_13__SCAN_IN), .ZN(n8050) );
  AOI22_X1 U6999 ( .A1(n7752), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n5407), .B2(
        n8050), .ZN(n5504) );
  NAND2_X1 U7000 ( .A1(n5398), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5511) );
  NAND2_X1 U7001 ( .A1(n5677), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n5510) );
  NAND2_X1 U7002 ( .A1(n5506), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n5507) );
  NAND2_X1 U7003 ( .A1(n5518), .A2(n5507), .ZN(n7524) );
  NAND2_X1 U7004 ( .A1(n5676), .A2(n7524), .ZN(n5509) );
  NAND2_X1 U7005 ( .A1(n5599), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n5508) );
  NAND4_X1 U7006 ( .A1(n5511), .A2(n5510), .A3(n5509), .A4(n5508), .ZN(n7997)
         );
  OR2_X1 U7007 ( .A1(n9286), .A2(n7997), .ZN(n7373) );
  INV_X1 U7008 ( .A(n7373), .ZN(n5512) );
  NAND2_X1 U7009 ( .A1(n9286), .A2(n7997), .ZN(n7372) );
  NAND2_X1 U7010 ( .A1(n6591), .A2(n7751), .ZN(n5517) );
  NAND2_X1 U7011 ( .A1(n5514), .A2(n5513), .ZN(n5515) );
  NAND2_X1 U7012 ( .A1(n5515), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5526) );
  XNOR2_X1 U7013 ( .A(n5526), .B(P2_IR_REG_14__SCAN_IN), .ZN(n8044) );
  AOI22_X1 U7014 ( .A1(n7752), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n5407), .B2(
        n8044), .ZN(n5516) );
  NAND2_X1 U7015 ( .A1(n5398), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5523) );
  NAND2_X1 U7016 ( .A1(n5677), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n5522) );
  NAND2_X1 U7017 ( .A1(n5518), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5519) );
  NAND2_X1 U7018 ( .A1(n5531), .A2(n5519), .ZN(n7868) );
  NAND2_X1 U7019 ( .A1(n5642), .A2(n7868), .ZN(n5521) );
  NAND2_X1 U7020 ( .A1(n5599), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n5520) );
  INV_X1 U7021 ( .A(n7376), .ZN(n7996) );
  INV_X1 U7022 ( .A(n7872), .ZN(n7478) );
  NAND2_X1 U7023 ( .A1(n6633), .A2(n7751), .ZN(n5530) );
  NAND2_X1 U7024 ( .A1(n5526), .A2(n5525), .ZN(n5527) );
  NAND2_X1 U7025 ( .A1(n5527), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5528) );
  XNOR2_X1 U7026 ( .A(n5528), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8042) );
  AOI22_X1 U7027 ( .A1(n7752), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n5407), .B2(
        n8042), .ZN(n5529) );
  NAND2_X1 U7028 ( .A1(n5398), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n5537) );
  NAND2_X1 U7029 ( .A1(n5677), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n5536) );
  NAND2_X1 U7030 ( .A1(n5531), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5532) );
  NAND2_X1 U7031 ( .A1(n5533), .A2(n5532), .ZN(n7988) );
  NAND2_X1 U7032 ( .A1(n5642), .A2(n7988), .ZN(n5535) );
  NAND2_X1 U7033 ( .A1(n5599), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n5534) );
  NAND2_X1 U7034 ( .A1(n7976), .A2(n7912), .ZN(n7694) );
  NAND2_X1 U7035 ( .A1(n7916), .A2(n7985), .ZN(n7610) );
  INV_X1 U7036 ( .A(n7912), .ZN(n7995) );
  NOR2_X1 U7037 ( .A1(n7976), .A2(n7995), .ZN(n7506) );
  NAND2_X1 U7038 ( .A1(n6706), .A2(n7751), .ZN(n5543) );
  INV_X1 U7039 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5538) );
  MUX2_X1 U7040 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5540), .S(
        P2_IR_REG_17__SCAN_IN), .Z(n5541) );
  AND2_X1 U7041 ( .A1(n5541), .A2(n5564), .ZN(n8039) );
  AOI22_X1 U7042 ( .A1(n7752), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n5407), .B2(
        n8039), .ZN(n5542) );
  NAND2_X1 U7043 ( .A1(n5398), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n5551) );
  NAND2_X1 U7044 ( .A1(n5677), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n5550) );
  INV_X1 U7045 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n5544) );
  NAND2_X1 U7046 ( .A1(n5546), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n5547) );
  NAND2_X1 U7047 ( .A1(n5556), .A2(n5547), .ZN(n8205) );
  NAND2_X1 U7048 ( .A1(n5642), .A2(n8205), .ZN(n5549) );
  NAND2_X1 U7049 ( .A1(n5599), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n5548) );
  NAND2_X1 U7050 ( .A1(n8317), .A2(n7994), .ZN(n7701) );
  INV_X1 U7051 ( .A(n8317), .ZN(n7931) );
  OR2_X1 U7052 ( .A1(n6764), .A2(n5552), .ZN(n5555) );
  NAND2_X1 U7053 ( .A1(n5564), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5553) );
  XNOR2_X1 U7054 ( .A(n5553), .B(P2_IR_REG_18__SCAN_IN), .ZN(n9204) );
  AOI22_X1 U7055 ( .A1(n7752), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n5407), .B2(
        n9204), .ZN(n5554) );
  INV_X1 U7056 ( .A(n8310), .ZN(n5562) );
  NAND2_X1 U7057 ( .A1(n5556), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5557) );
  NAND2_X1 U7058 ( .A1(n5568), .A2(n5557), .ZN(n8196) );
  NAND2_X1 U7059 ( .A1(n8196), .A2(n5642), .ZN(n5561) );
  NAND2_X1 U7060 ( .A1(n5398), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n5560) );
  NAND2_X1 U7061 ( .A1(n5677), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n5559) );
  NAND2_X1 U7062 ( .A1(n5599), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n5558) );
  NOR2_X1 U7063 ( .A1(n5562), .A2(n7885), .ZN(n5563) );
  INV_X1 U7064 ( .A(n7885), .ZN(n8203) );
  NAND2_X1 U7065 ( .A1(n6848), .A2(n7751), .ZN(n5567) );
  XNOR2_X2 U7066 ( .A(n5565), .B(P2_IR_REG_19__SCAN_IN), .ZN(n8020) );
  AOI22_X1 U7067 ( .A1(n7752), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n8020), .B2(
        n5407), .ZN(n5566) );
  INV_X1 U7068 ( .A(n8304), .ZN(n5573) );
  INV_X1 U7069 ( .A(n5579), .ZN(n5580) );
  NAND2_X1 U7070 ( .A1(n5568), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n5569) );
  NAND2_X1 U7071 ( .A1(n5580), .A2(n5569), .ZN(n8184) );
  NAND2_X1 U7072 ( .A1(n8184), .A2(n5642), .ZN(n5572) );
  AOI22_X1 U7073 ( .A1(n5398), .A2(P2_REG0_REG_19__SCAN_IN), .B1(n5677), .B2(
        P2_REG2_REG_19__SCAN_IN), .ZN(n5571) );
  NAND2_X1 U7074 ( .A1(n5599), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n5570) );
  NAND2_X1 U7075 ( .A1(n5573), .A2(n7947), .ZN(n5575) );
  INV_X1 U7076 ( .A(n7947), .ZN(n8193) );
  AOI21_X1 U7077 ( .B1(n5576), .B2(n5575), .A(n5574), .ZN(n8170) );
  NAND2_X1 U7078 ( .A1(n6832), .A2(n7751), .ZN(n5578) );
  NAND2_X1 U7079 ( .A1(n7752), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n5577) );
  INV_X1 U7080 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n10021) );
  INV_X1 U7081 ( .A(n5589), .ZN(n5590) );
  NAND2_X1 U7082 ( .A1(n5580), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n5581) );
  NAND2_X1 U7083 ( .A1(n5590), .A2(n5581), .ZN(n8174) );
  NAND2_X1 U7084 ( .A1(n8174), .A2(n5676), .ZN(n5584) );
  AOI22_X1 U7085 ( .A1(n5398), .A2(P2_REG0_REG_20__SCAN_IN), .B1(n5416), .B2(
        P2_REG2_REG_20__SCAN_IN), .ZN(n5583) );
  NAND2_X1 U7086 ( .A1(n5599), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n5582) );
  INV_X1 U7087 ( .A(n7710), .ZN(n5585) );
  NAND2_X1 U7088 ( .A1(n8298), .A2(n7893), .ZN(n7713) );
  INV_X1 U7089 ( .A(n7713), .ZN(n5717) );
  NOR2_X1 U7090 ( .A1(n5585), .A2(n5717), .ZN(n7795) );
  INV_X1 U7091 ( .A(n7795), .ZN(n8169) );
  INV_X1 U7092 ( .A(n8298), .ZN(n5586) );
  NAND2_X1 U7093 ( .A1(n5586), .A2(n7893), .ZN(n8157) );
  NAND2_X1 U7094 ( .A1(n6855), .A2(n7751), .ZN(n5588) );
  NAND2_X1 U7095 ( .A1(n7752), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n5587) );
  INV_X1 U7096 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n10019) );
  NAND2_X1 U7097 ( .A1(n5590), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n5591) );
  NAND2_X1 U7098 ( .A1(n5597), .A2(n5591), .ZN(n8164) );
  NAND2_X1 U7099 ( .A1(n8164), .A2(n5642), .ZN(n5594) );
  AOI22_X1 U7100 ( .A1(n5398), .A2(P2_REG0_REG_21__SCAN_IN), .B1(n5677), .B2(
        P2_REG2_REG_21__SCAN_IN), .ZN(n5593) );
  NAND2_X1 U7101 ( .A1(n5599), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n5592) );
  NAND2_X1 U7102 ( .A1(n8292), .A2(n7957), .ZN(n7714) );
  NAND2_X1 U7103 ( .A1(n7716), .A2(n7714), .ZN(n7797) );
  INV_X1 U7104 ( .A(n7957), .ZN(n8171) );
  NOR2_X1 U7105 ( .A1(n8292), .A2(n8171), .ZN(n8146) );
  NAND2_X1 U7106 ( .A1(n7060), .A2(n7751), .ZN(n5596) );
  NAND2_X1 U7107 ( .A1(n7752), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n5595) );
  NAND2_X1 U7108 ( .A1(n5597), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n5598) );
  NAND2_X1 U7109 ( .A1(n5608), .A2(n5598), .ZN(n8152) );
  NAND2_X1 U7110 ( .A1(n8152), .A2(n5642), .ZN(n5604) );
  INV_X1 U7111 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n8229) );
  NAND2_X1 U7112 ( .A1(n5398), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n5601) );
  NAND2_X1 U7113 ( .A1(n5677), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n5600) );
  OAI211_X1 U7114 ( .C1(n8229), .C2(n7757), .A(n5601), .B(n5600), .ZN(n5602)
         );
  INV_X1 U7115 ( .A(n5602), .ZN(n5603) );
  NOR2_X1 U7116 ( .A1(n8286), .A2(n5844), .ZN(n7718) );
  INV_X1 U7117 ( .A(n7718), .ZN(n5718) );
  NAND2_X1 U7118 ( .A1(n5718), .A2(n4844), .ZN(n8145) );
  INV_X1 U7119 ( .A(n8286), .ZN(n7963) );
  NAND2_X1 U7120 ( .A1(n7963), .A2(n5844), .ZN(n5605) );
  NAND2_X1 U7121 ( .A1(n7076), .A2(n7751), .ZN(n5607) );
  NAND2_X1 U7122 ( .A1(n7752), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n5606) );
  NAND2_X1 U7123 ( .A1(n5608), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5609) );
  NAND2_X1 U7124 ( .A1(n5619), .A2(n5609), .ZN(n8141) );
  NAND2_X1 U7125 ( .A1(n8141), .A2(n5676), .ZN(n5614) );
  INV_X1 U7126 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n8226) );
  NAND2_X1 U7127 ( .A1(n5677), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n5611) );
  NAND2_X1 U7128 ( .A1(n5398), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n5610) );
  OAI211_X1 U7129 ( .C1(n8226), .C2(n7757), .A(n5611), .B(n5610), .ZN(n5612)
         );
  INV_X1 U7130 ( .A(n5612), .ZN(n5613) );
  NAND2_X1 U7131 ( .A1(n8280), .A2(n8149), .ZN(n5616) );
  NOR2_X1 U7132 ( .A1(n8280), .A2(n8149), .ZN(n5615) );
  NAND2_X1 U7133 ( .A1(n7117), .A2(n7751), .ZN(n5618) );
  NAND2_X1 U7134 ( .A1(n7752), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n5617) );
  INV_X1 U7135 ( .A(n8273), .ZN(n8121) );
  INV_X1 U7136 ( .A(n5628), .ZN(n5629) );
  NAND2_X1 U7137 ( .A1(n5619), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n5620) );
  NAND2_X1 U7138 ( .A1(n5629), .A2(n5620), .ZN(n8127) );
  NAND2_X1 U7139 ( .A1(n8127), .A2(n5642), .ZN(n5625) );
  INV_X1 U7140 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n8222) );
  NAND2_X1 U7141 ( .A1(n5677), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n5622) );
  NAND2_X1 U7142 ( .A1(n5398), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n5621) );
  OAI211_X1 U7143 ( .C1(n8222), .C2(n7757), .A(n5622), .B(n5621), .ZN(n5623)
         );
  INV_X1 U7144 ( .A(n5623), .ZN(n5624) );
  NAND2_X1 U7145 ( .A1(n7227), .A2(n7751), .ZN(n5627) );
  NAND2_X1 U7146 ( .A1(n7752), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n5626) );
  INV_X1 U7147 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n10050) );
  NAND2_X1 U7148 ( .A1(n5628), .A2(n10050), .ZN(n5640) );
  NAND2_X1 U7149 ( .A1(n5629), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n5630) );
  NAND2_X1 U7150 ( .A1(n5640), .A2(n5630), .ZN(n8115) );
  NAND2_X1 U7151 ( .A1(n8115), .A2(n5642), .ZN(n5635) );
  INV_X1 U7152 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n8219) );
  NAND2_X1 U7153 ( .A1(n5398), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n5632) );
  NAND2_X1 U7154 ( .A1(n5416), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n5631) );
  OAI211_X1 U7155 ( .C1(n8219), .C2(n7757), .A(n5632), .B(n5631), .ZN(n5633)
         );
  INV_X1 U7156 ( .A(n5633), .ZN(n5634) );
  NAND2_X1 U7157 ( .A1(n8267), .A2(n7938), .ZN(n7730) );
  INV_X1 U7158 ( .A(n8267), .ZN(n8108) );
  NAND2_X1 U7159 ( .A1(n8108), .A2(n7938), .ZN(n5637) );
  NAND2_X1 U7160 ( .A1(n8109), .A2(n5637), .ZN(n8100) );
  NAND2_X1 U7161 ( .A1(n7258), .A2(n7751), .ZN(n5639) );
  NAND2_X1 U7162 ( .A1(n7752), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n5638) );
  NAND2_X1 U7163 ( .A1(n5640), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n5641) );
  NAND2_X1 U7164 ( .A1(n5652), .A2(n5641), .ZN(n8105) );
  NAND2_X1 U7165 ( .A1(n8105), .A2(n5642), .ZN(n5647) );
  INV_X1 U7166 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n8216) );
  NAND2_X1 U7167 ( .A1(n5398), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n5644) );
  NAND2_X1 U7168 ( .A1(n5416), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n5643) );
  OAI211_X1 U7169 ( .C1(n8216), .C2(n7757), .A(n5644), .B(n5643), .ZN(n5645)
         );
  INV_X1 U7170 ( .A(n5645), .ZN(n5646) );
  NAND2_X1 U7171 ( .A1(n8261), .A2(n8111), .ZN(n5648) );
  INV_X1 U7172 ( .A(n8261), .ZN(n6386) );
  NAND2_X1 U7173 ( .A1(n6386), .A2(n7904), .ZN(n5649) );
  NAND2_X1 U7174 ( .A1(n7356), .A2(n7751), .ZN(n5651) );
  NAND2_X1 U7175 ( .A1(n7752), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n5650) );
  INV_X1 U7176 ( .A(n5663), .ZN(n5664) );
  NAND2_X1 U7177 ( .A1(n5652), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n5653) );
  NAND2_X1 U7178 ( .A1(n5664), .A2(n5653), .ZN(n8096) );
  NAND2_X1 U7179 ( .A1(n8096), .A2(n5642), .ZN(n5658) );
  INV_X1 U7180 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n8213) );
  NAND2_X1 U7181 ( .A1(n5398), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n5655) );
  NAND2_X1 U7182 ( .A1(n5416), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n5654) );
  OAI211_X1 U7183 ( .C1(n8213), .C2(n7757), .A(n5655), .B(n5654), .ZN(n5656)
         );
  INV_X1 U7184 ( .A(n5656), .ZN(n5657) );
  NOR2_X1 U7185 ( .A1(n8257), .A2(n8102), .ZN(n5659) );
  NAND2_X1 U7186 ( .A1(n7395), .A2(n7751), .ZN(n5661) );
  NAND2_X1 U7187 ( .A1(n7752), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n5660) );
  INV_X1 U7188 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n5662) );
  INV_X1 U7189 ( .A(n7859), .ZN(n5666) );
  NAND2_X1 U7190 ( .A1(n5664), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n5665) );
  NAND2_X1 U7191 ( .A1(n5666), .A2(n5665), .ZN(n8085) );
  NAND2_X1 U7192 ( .A1(n8085), .A2(n5642), .ZN(n5671) );
  INV_X1 U7193 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n8209) );
  NAND2_X1 U7194 ( .A1(n5398), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n5668) );
  NAND2_X1 U7195 ( .A1(n5677), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n5667) );
  OAI211_X1 U7196 ( .C1(n8209), .C2(n7757), .A(n5668), .B(n5667), .ZN(n5669)
         );
  INV_X1 U7197 ( .A(n5669), .ZN(n5670) );
  XNOR2_X2 U7198 ( .A(n8086), .B(n5722), .ZN(n8077) );
  NOR2_X1 U7199 ( .A1(n4721), .A2(n5722), .ZN(n5672) );
  NAND2_X1 U7200 ( .A1(n7752), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n5674) );
  NAND2_X1 U7201 ( .A1(n7859), .A2(n5676), .ZN(n7761) );
  INV_X1 U7202 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n5680) );
  NAND2_X1 U7203 ( .A1(n5398), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n5679) );
  NAND2_X1 U7204 ( .A1(n5677), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n5678) );
  OAI211_X1 U7205 ( .C1(n5680), .C2(n7757), .A(n5679), .B(n5678), .ZN(n5681)
         );
  INV_X1 U7206 ( .A(n5681), .ZN(n5682) );
  NAND2_X1 U7207 ( .A1(n5683), .A2(n8081), .ZN(n7740) );
  XNOR2_X1 U7208 ( .A(n5684), .B(n7800), .ZN(n5702) );
  NAND2_X1 U7209 ( .A1(n5685), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5686) );
  XNOR2_X1 U7210 ( .A(n5686), .B(P2_IR_REG_22__SCAN_IN), .ZN(n7817) );
  NAND2_X1 U7211 ( .A1(n8020), .A2(n7817), .ZN(n5692) );
  NAND2_X1 U7212 ( .A1(n4368), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5687) );
  NAND2_X1 U7213 ( .A1(n5688), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5689) );
  MUX2_X1 U7214 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5689), .S(
        P2_IR_REG_20__SCAN_IN), .Z(n5690) );
  NAND2_X1 U7215 ( .A1(n5690), .A2(n4368), .ZN(n7806) );
  NAND2_X1 U7216 ( .A1(n7808), .A2(n7807), .ZN(n5691) );
  INV_X1 U7217 ( .A(n5693), .ZN(n7814) );
  NAND2_X1 U7218 ( .A1(n7814), .A2(n6419), .ZN(n5694) );
  NAND2_X1 U7219 ( .A1(n5885), .A2(n7732), .ZN(n9762) );
  INV_X1 U7220 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n5697) );
  NAND2_X1 U7221 ( .A1(n5398), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n5696) );
  NAND2_X1 U7222 ( .A1(n5416), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n5695) );
  OAI211_X1 U7223 ( .C1(n5697), .C2(n7757), .A(n5696), .B(n5695), .ZN(n5698)
         );
  INV_X1 U7224 ( .A(n5698), .ZN(n5699) );
  AND2_X1 U7225 ( .A1(n7761), .A2(n5699), .ZN(n7741) );
  NAND2_X1 U7226 ( .A1(n5379), .A2(P2_B_REG_SCAN_IN), .ZN(n5700) );
  NAND2_X1 U7227 ( .A1(n9746), .A2(n5700), .ZN(n8068) );
  OAI22_X1 U7228 ( .A1(n5722), .A2(n9762), .B1(n7741), .B2(n8068), .ZN(n5701)
         );
  AOI21_X1 U7229 ( .B1(n5702), .B2(n9765), .A(n5701), .ZN(n7865) );
  INV_X1 U7230 ( .A(n6661), .ZN(n5704) );
  NAND2_X1 U7231 ( .A1(n5704), .A2(n5703), .ZN(n6662) );
  NAND2_X1 U7232 ( .A1(n6662), .A2(n7613), .ZN(n9756) );
  NAND2_X1 U7233 ( .A1(n9756), .A2(n7619), .ZN(n5705) );
  NAND2_X1 U7234 ( .A1(n5781), .A2(n5780), .ZN(n7624) );
  NAND2_X1 U7235 ( .A1(n5705), .A2(n7624), .ZN(n9749) );
  XNOR2_X1 U7236 ( .A(n8004), .B(n9789), .ZN(n9750) );
  NAND2_X1 U7237 ( .A1(n9749), .A2(n9750), .ZN(n5706) );
  NAND2_X1 U7238 ( .A1(n9761), .A2(n9789), .ZN(n7638) );
  NAND2_X1 U7239 ( .A1(n5706), .A2(n7638), .ZN(n6788) );
  NAND2_X1 U7240 ( .A1(n6788), .A2(n7773), .ZN(n5707) );
  NAND2_X1 U7241 ( .A1(n5707), .A2(n7632), .ZN(n6867) );
  NAND2_X1 U7242 ( .A1(n5437), .A2(n6879), .ZN(n6841) );
  NAND2_X1 U7243 ( .A1(n8003), .A2(n9801), .ZN(n7639) );
  NAND2_X1 U7244 ( .A1(n6867), .A2(n7775), .ZN(n6866) );
  NAND2_X1 U7245 ( .A1(n7091), .A2(n6863), .ZN(n7635) );
  AND2_X1 U7246 ( .A1(n6841), .A2(n7635), .ZN(n7644) );
  NAND2_X1 U7247 ( .A1(n6866), .A2(n7644), .ZN(n5709) );
  AND2_X1 U7248 ( .A1(n5434), .A2(n6860), .ZN(n7643) );
  INV_X1 U7249 ( .A(n7643), .ZN(n5708) );
  NAND2_X1 U7250 ( .A1(n5709), .A2(n5708), .ZN(n7087) );
  NAND2_X1 U7251 ( .A1(n7087), .A2(n7779), .ZN(n6990) );
  NAND2_X1 U7252 ( .A1(n7648), .A2(n6991), .ZN(n7663) );
  INV_X1 U7253 ( .A(n7663), .ZN(n5710) );
  NAND2_X1 U7254 ( .A1(n7668), .A2(n7649), .ZN(n7660) );
  INV_X1 U7255 ( .A(n7660), .ZN(n5712) );
  OR2_X1 U7256 ( .A1(n9825), .A2(n7451), .ZN(n7673) );
  NAND2_X1 U7257 ( .A1(n9825), .A2(n7451), .ZN(n7672) );
  NAND2_X1 U7258 ( .A1(n7223), .A2(n7782), .ZN(n5713) );
  NAND2_X1 U7259 ( .A1(n5713), .A2(n7672), .ZN(n7351) );
  INV_X1 U7260 ( .A(n7351), .ZN(n5714) );
  NAND2_X1 U7261 ( .A1(n5714), .A2(n7787), .ZN(n7349) );
  NAND2_X1 U7262 ( .A1(n5501), .A2(n7998), .ZN(n7681) );
  NAND2_X1 U7263 ( .A1(n7349), .A2(n7681), .ZN(n7381) );
  AND2_X1 U7264 ( .A1(n9286), .A2(n7348), .ZN(n7686) );
  INV_X1 U7265 ( .A(n7686), .ZN(n5715) );
  NOR2_X1 U7266 ( .A1(n9286), .A2(n7348), .ZN(n7685) );
  OR2_X1 U7267 ( .A1(n7872), .A2(n7376), .ZN(n7690) );
  NAND2_X1 U7268 ( .A1(n7872), .A2(n7376), .ZN(n7689) );
  INV_X1 U7269 ( .A(n7689), .ZN(n5716) );
  NAND2_X1 U7270 ( .A1(n8199), .A2(n7701), .ZN(n8188) );
  OR2_X1 U7271 ( .A1(n8310), .A2(n7885), .ZN(n7772) );
  AND2_X1 U7272 ( .A1(n7772), .A2(n8187), .ZN(n7699) );
  NAND2_X1 U7273 ( .A1(n8310), .A2(n7885), .ZN(n7771) );
  AOI21_X1 U7274 ( .B1(n8188), .B2(n7699), .A(n4512), .ZN(n8178) );
  OR2_X1 U7275 ( .A1(n8304), .A2(n7947), .ZN(n7709) );
  NAND2_X1 U7276 ( .A1(n7709), .A2(n7706), .ZN(n8179) );
  OAI21_X1 U7277 ( .B1(n8178), .B2(n8179), .A(n7706), .ZN(n8167) );
  AOI21_X1 U7278 ( .B1(n8167), .B2(n7710), .A(n5717), .ZN(n8155) );
  NAND2_X1 U7279 ( .A1(n8273), .A2(n7903), .ZN(n7768) );
  NAND2_X1 U7280 ( .A1(n8280), .A2(n7958), .ZN(n8128) );
  NAND2_X1 U7281 ( .A1(n7768), .A2(n8128), .ZN(n7723) );
  INV_X1 U7282 ( .A(n7729), .ZN(n5719) );
  NAND2_X1 U7283 ( .A1(n8261), .A2(n7904), .ZN(n7727) );
  INV_X1 U7284 ( .A(n7727), .ZN(n5720) );
  INV_X1 U7285 ( .A(n8257), .ZN(n5721) );
  XNOR2_X1 U7286 ( .A(n7765), .B(n7737), .ZN(n7861) );
  INV_X1 U7287 ( .A(n8020), .ZN(n8064) );
  AND2_X1 U7288 ( .A1(n8064), .A2(n7817), .ZN(n6361) );
  AND2_X1 U7289 ( .A1(n7808), .A2(n7806), .ZN(n6664) );
  AND2_X1 U7290 ( .A1(n6361), .A2(n6664), .ZN(n5883) );
  NOR2_X1 U7291 ( .A1(n5883), .A2(n9835), .ZN(n6608) );
  INV_X1 U7292 ( .A(n6361), .ZN(n5723) );
  NAND2_X1 U7293 ( .A1(n5723), .A2(n5774), .ZN(n5724) );
  NAND2_X1 U7294 ( .A1(n6608), .A2(n5724), .ZN(n9768) );
  NAND2_X1 U7295 ( .A1(n8020), .A2(n7806), .ZN(n9771) );
  NAND2_X1 U7296 ( .A1(n7865), .A2(n5725), .ZN(n6368) );
  NAND2_X1 U7297 ( .A1(n5755), .A2(n5756), .ZN(n5727) );
  NAND2_X1 U7298 ( .A1(n5727), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5729) );
  NAND2_X1 U7299 ( .A1(n5729), .A2(n5728), .ZN(n5732) );
  OR2_X1 U7300 ( .A1(n5729), .A2(n5728), .ZN(n5730) );
  NAND2_X1 U7301 ( .A1(n5732), .A2(n5730), .ZN(n7120) );
  INV_X1 U7302 ( .A(P2_B_REG_SCAN_IN), .ZN(n5731) );
  XNOR2_X1 U7303 ( .A(n7120), .B(n5731), .ZN(n5738) );
  NAND2_X1 U7304 ( .A1(n5732), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5733) );
  INV_X1 U7305 ( .A(n5734), .ZN(n5735) );
  NAND2_X1 U7306 ( .A1(n5735), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5736) );
  MUX2_X1 U7307 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5736), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n5737) );
  NAND2_X1 U7308 ( .A1(n5737), .A2(n5348), .ZN(n5753) );
  NAND2_X1 U7309 ( .A1(n5753), .A2(n7120), .ZN(n6443) );
  OR2_X1 U7310 ( .A1(n5739), .A2(P2_D_REG_1__SCAN_IN), .ZN(n5741) );
  OR2_X1 U7311 ( .A1(n7259), .A2(n7228), .ZN(n5740) );
  NOR2_X1 U7312 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .ZN(
        n5745) );
  NOR4_X1 U7313 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_22__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n5744) );
  NOR4_X1 U7314 ( .A1(P2_D_REG_12__SCAN_IN), .A2(P2_D_REG_25__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_23__SCAN_IN), .ZN(n5743) );
  NOR4_X1 U7315 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_28__SCAN_IN), .A3(
        P2_D_REG_27__SCAN_IN), .A4(P2_D_REG_26__SCAN_IN), .ZN(n5742) );
  NAND4_X1 U7316 ( .A1(n5745), .A2(n5744), .A3(n5743), .A4(n5742), .ZN(n5751)
         );
  NOR4_X1 U7317 ( .A1(P2_D_REG_14__SCAN_IN), .A2(P2_D_REG_13__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n5749) );
  NOR4_X1 U7318 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_9__SCAN_IN), .A3(
        P2_D_REG_17__SCAN_IN), .A4(P2_D_REG_15__SCAN_IN), .ZN(n5748) );
  NOR4_X1 U7319 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n5747) );
  NOR4_X1 U7320 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_19__SCAN_IN), .ZN(n5746) );
  NAND4_X1 U7321 ( .A1(n5749), .A2(n5748), .A3(n5747), .A4(n5746), .ZN(n5750)
         );
  NOR2_X1 U7322 ( .A1(n5751), .A2(n5750), .ZN(n5752) );
  OR2_X1 U7323 ( .A1(n5739), .A2(n5752), .ZN(n6357) );
  NAND2_X1 U7324 ( .A1(n6359), .A2(n6357), .ZN(n5889) );
  NOR2_X1 U7325 ( .A1(n5753), .A2(n7120), .ZN(n5754) );
  NAND2_X1 U7326 ( .A1(n7228), .A2(n5754), .ZN(n6417) );
  XNOR2_X1 U7327 ( .A(n5755), .B(n5756), .ZN(n6403) );
  INV_X1 U7328 ( .A(n6439), .ZN(n5757) );
  NOR2_X1 U7329 ( .A1(n5889), .A2(n5757), .ZN(n5880) );
  NOR2_X1 U7330 ( .A1(n7808), .A2(n7806), .ZN(n5771) );
  AND2_X1 U7331 ( .A1(n5771), .A2(n7817), .ZN(n5758) );
  NAND2_X1 U7332 ( .A1(n8020), .A2(n5758), .ZN(n5761) );
  INV_X1 U7333 ( .A(n5761), .ZN(n5891) );
  OR2_X1 U7334 ( .A1(n5883), .A2(n5891), .ZN(n5759) );
  NAND2_X1 U7335 ( .A1(n5880), .A2(n5759), .ZN(n5765) );
  INV_X1 U7336 ( .A(n6602), .ZN(n5760) );
  NOR2_X1 U7337 ( .A1(n9835), .A2(n7732), .ZN(n5762) );
  AND2_X1 U7338 ( .A1(n5762), .A2(n5761), .ZN(n5876) );
  INV_X1 U7339 ( .A(n5876), .ZN(n5763) );
  NAND2_X1 U7340 ( .A1(n9771), .A2(n9835), .ZN(n8120) );
  NAND2_X1 U7341 ( .A1(n5763), .A2(n8120), .ZN(n5888) );
  NAND3_X1 U7342 ( .A1(n5882), .A2(n6439), .A3(n5888), .ZN(n5764) );
  INV_X2 U7343 ( .A(n9838), .ZN(n9836) );
  INV_X1 U7344 ( .A(n5683), .ZN(n6369) );
  NOR2_X1 U7345 ( .A1(n6369), .A2(n8254), .ZN(n5766) );
  NOR2_X1 U7346 ( .A1(n9836), .A2(n5767), .ZN(n5768) );
  NAND2_X1 U7347 ( .A1(n5770), .A2(n5769), .ZN(P2_U3456) );
  INV_X1 U7348 ( .A(n6664), .ZN(n5773) );
  NAND2_X1 U7349 ( .A1(n5801), .A2(n6614), .ZN(n5777) );
  AND2_X1 U7350 ( .A1(n7612), .A2(n5777), .ZN(n6574) );
  NAND2_X1 U7351 ( .A1(n5778), .A2(n9763), .ZN(n5779) );
  XNOR2_X1 U7352 ( .A(n4353), .B(n5780), .ZN(n5782) );
  XNOR2_X1 U7353 ( .A(n5782), .B(n9745), .ZN(n6584) );
  AND2_X1 U7354 ( .A1(n5782), .A2(n5781), .ZN(n5783) );
  XNOR2_X1 U7355 ( .A(n7622), .B(n4353), .ZN(n5784) );
  XNOR2_X1 U7356 ( .A(n5784), .B(n9761), .ZN(n6619) );
  NAND2_X1 U7357 ( .A1(n5784), .A2(n8004), .ZN(n5785) );
  XNOR2_X1 U7358 ( .A(n4353), .B(n6795), .ZN(n5787) );
  XNOR2_X1 U7359 ( .A(n5787), .B(n6872), .ZN(n6678) );
  INV_X1 U7360 ( .A(n6678), .ZN(n5786) );
  NAND2_X1 U7361 ( .A1(n5787), .A2(n6872), .ZN(n5788) );
  NAND2_X1 U7362 ( .A1(n6675), .A2(n5788), .ZN(n6733) );
  XNOR2_X1 U7363 ( .A(n4353), .B(n9801), .ZN(n5789) );
  XNOR2_X1 U7364 ( .A(n5789), .B(n5437), .ZN(n6734) );
  NAND2_X1 U7365 ( .A1(n6733), .A2(n6734), .ZN(n5791) );
  OR2_X1 U7366 ( .A1(n5789), .A2(n8003), .ZN(n5790) );
  NAND2_X1 U7367 ( .A1(n5791), .A2(n5790), .ZN(n6779) );
  INV_X1 U7368 ( .A(n6779), .ZN(n5793) );
  XNOR2_X1 U7369 ( .A(n4353), .B(n6863), .ZN(n5794) );
  XNOR2_X1 U7370 ( .A(n5794), .B(n7091), .ZN(n6778) );
  INV_X1 U7371 ( .A(n6778), .ZN(n5792) );
  INV_X1 U7372 ( .A(n5794), .ZN(n5795) );
  NAND2_X1 U7373 ( .A1(n5795), .A2(n5434), .ZN(n5796) );
  XNOR2_X1 U7374 ( .A(n7101), .B(n4353), .ZN(n5797) );
  XNOR2_X1 U7375 ( .A(n5797), .B(n6783), .ZN(n6940) );
  NAND2_X1 U7376 ( .A1(n5797), .A2(n6986), .ZN(n5798) );
  XNOR2_X1 U7377 ( .A(n9814), .B(n4353), .ZN(n5799) );
  AND2_X1 U7378 ( .A1(n5799), .A2(n7090), .ZN(n6949) );
  INV_X1 U7379 ( .A(n5799), .ZN(n5800) );
  NAND2_X1 U7380 ( .A1(n5800), .A2(n8002), .ZN(n6950) );
  XNOR2_X1 U7381 ( .A(n9823), .B(n4357), .ZN(n5802) );
  XNOR2_X1 U7382 ( .A(n5802), .B(n7282), .ZN(n7080) );
  NAND2_X1 U7383 ( .A1(n7081), .A2(n7080), .ZN(n7079) );
  NAND2_X1 U7384 ( .A1(n5802), .A2(n8001), .ZN(n5803) );
  XNOR2_X1 U7385 ( .A(n7284), .B(n4353), .ZN(n7278) );
  XNOR2_X1 U7386 ( .A(n7782), .B(n4357), .ZN(n7384) );
  NAND2_X1 U7387 ( .A1(n7384), .A2(n7999), .ZN(n5806) );
  NAND2_X1 U7388 ( .A1(n7385), .A2(n5806), .ZN(n7448) );
  XNOR2_X1 U7389 ( .A(n9834), .B(n4353), .ZN(n5807) );
  XNOR2_X1 U7390 ( .A(n5807), .B(n7998), .ZN(n7447) );
  INV_X1 U7391 ( .A(n5807), .ZN(n5808) );
  NAND2_X1 U7392 ( .A1(n5808), .A2(n7998), .ZN(n5809) );
  XNOR2_X1 U7393 ( .A(n9286), .B(n4353), .ZN(n5811) );
  XNOR2_X1 U7394 ( .A(n5811), .B(n7348), .ZN(n7523) );
  NAND2_X1 U7395 ( .A1(n5811), .A2(n7348), .ZN(n5812) );
  NAND2_X1 U7396 ( .A1(n7520), .A2(n5812), .ZN(n7867) );
  XNOR2_X1 U7397 ( .A(n7872), .B(n4357), .ZN(n5813) );
  XNOR2_X1 U7398 ( .A(n5813), .B(n7376), .ZN(n7866) );
  NAND2_X1 U7399 ( .A1(n7867), .A2(n7866), .ZN(n5816) );
  INV_X1 U7400 ( .A(n5813), .ZN(n5814) );
  NAND2_X1 U7401 ( .A1(n5814), .A2(n7376), .ZN(n5815) );
  NAND2_X1 U7402 ( .A1(n5816), .A2(n5815), .ZN(n7979) );
  INV_X1 U7403 ( .A(n7979), .ZN(n5818) );
  XNOR2_X1 U7404 ( .A(n7976), .B(n4353), .ZN(n5819) );
  XNOR2_X1 U7405 ( .A(n5819), .B(n7912), .ZN(n7978) );
  INV_X1 U7406 ( .A(n5819), .ZN(n5820) );
  NAND2_X1 U7407 ( .A1(n5820), .A2(n7995), .ZN(n5821) );
  XNOR2_X1 U7408 ( .A(n7916), .B(n4353), .ZN(n5823) );
  XNOR2_X1 U7409 ( .A(n5823), .B(n7985), .ZN(n7911) );
  NAND2_X1 U7410 ( .A1(n5823), .A2(n7985), .ZN(n7920) );
  NAND2_X1 U7411 ( .A1(n7909), .A2(n7920), .ZN(n7924) );
  XNOR2_X1 U7412 ( .A(n8317), .B(n4357), .ZN(n5825) );
  XNOR2_X1 U7413 ( .A(n5825), .B(n7994), .ZN(n7923) );
  XNOR2_X1 U7414 ( .A(n8310), .B(n4357), .ZN(n5828) );
  XNOR2_X1 U7415 ( .A(n5828), .B(n7885), .ZN(n7967) );
  AND2_X1 U7416 ( .A1(n7923), .A2(n7967), .ZN(n5824) );
  NAND2_X1 U7417 ( .A1(n7924), .A2(n5824), .ZN(n5831) );
  INV_X1 U7418 ( .A(n7967), .ZN(n5827) );
  INV_X1 U7419 ( .A(n5825), .ZN(n5826) );
  NAND2_X1 U7420 ( .A1(n5826), .A2(n7994), .ZN(n7964) );
  INV_X1 U7421 ( .A(n5828), .ZN(n5829) );
  NAND2_X1 U7422 ( .A1(n5831), .A2(n5830), .ZN(n7881) );
  XNOR2_X1 U7423 ( .A(n8304), .B(n4357), .ZN(n5832) );
  XNOR2_X1 U7424 ( .A(n5832), .B(n7947), .ZN(n7882) );
  NAND2_X1 U7425 ( .A1(n7881), .A2(n7882), .ZN(n5835) );
  INV_X1 U7426 ( .A(n5832), .ZN(n5833) );
  NAND2_X1 U7427 ( .A1(n5833), .A2(n7947), .ZN(n5834) );
  NAND2_X1 U7428 ( .A1(n5835), .A2(n5834), .ZN(n7943) );
  XNOR2_X1 U7429 ( .A(n8298), .B(n4357), .ZN(n5836) );
  XNOR2_X1 U7430 ( .A(n5836), .B(n7893), .ZN(n7944) );
  NAND2_X1 U7431 ( .A1(n7943), .A2(n7944), .ZN(n5839) );
  INV_X1 U7432 ( .A(n5836), .ZN(n5837) );
  NAND2_X1 U7433 ( .A1(n5837), .A2(n7893), .ZN(n5838) );
  XNOR2_X1 U7434 ( .A(n8292), .B(n4357), .ZN(n5840) );
  XNOR2_X1 U7435 ( .A(n5840), .B(n7957), .ZN(n7890) );
  NAND2_X1 U7436 ( .A1(n7889), .A2(n7890), .ZN(n5843) );
  INV_X1 U7437 ( .A(n5840), .ZN(n5841) );
  NAND2_X1 U7438 ( .A1(n5841), .A2(n7957), .ZN(n5842) );
  NAND2_X1 U7439 ( .A1(n5843), .A2(n5842), .ZN(n7951) );
  XNOR2_X1 U7440 ( .A(n8286), .B(n4353), .ZN(n7952) );
  AND2_X1 U7441 ( .A1(n7952), .A2(n5844), .ZN(n5847) );
  INV_X1 U7442 ( .A(n7952), .ZN(n5845) );
  NAND2_X1 U7443 ( .A1(n5845), .A2(n8161), .ZN(n5846) );
  XNOR2_X1 U7444 ( .A(n8280), .B(n4357), .ZN(n5848) );
  OR2_X2 U7445 ( .A1(n5849), .A2(n5848), .ZN(n7932) );
  NAND2_X1 U7446 ( .A1(n5849), .A2(n5848), .ZN(n5850) );
  XNOR2_X1 U7447 ( .A(n8273), .B(n4353), .ZN(n5851) );
  NAND2_X1 U7448 ( .A1(n5851), .A2(n7903), .ZN(n7898) );
  INV_X1 U7449 ( .A(n5851), .ZN(n5852) );
  NAND2_X1 U7450 ( .A1(n5852), .A2(n8138), .ZN(n5853) );
  NAND2_X2 U7451 ( .A1(n5854), .A2(n7933), .ZN(n7897) );
  XNOR2_X1 U7452 ( .A(n8261), .B(n4357), .ZN(n5856) );
  XNOR2_X1 U7453 ( .A(n5856), .B(n7904), .ZN(n6376) );
  INV_X1 U7454 ( .A(n6376), .ZN(n5855) );
  XNOR2_X1 U7455 ( .A(n8267), .B(n4353), .ZN(n5863) );
  NAND2_X1 U7456 ( .A1(n5863), .A2(n7938), .ZN(n6375) );
  OR2_X1 U7457 ( .A1(n5855), .A2(n6375), .ZN(n5862) );
  AND2_X1 U7458 ( .A1(n7898), .A2(n5862), .ZN(n6378) );
  INV_X1 U7459 ( .A(n5856), .ZN(n5857) );
  NAND2_X1 U7460 ( .A1(n5857), .A2(n7904), .ZN(n5861) );
  AND2_X1 U7461 ( .A1(n6378), .A2(n5861), .ZN(n5873) );
  XNOR2_X1 U7462 ( .A(n8257), .B(n4353), .ZN(n6395) );
  XNOR2_X1 U7463 ( .A(n6395), .B(n8080), .ZN(n5874) );
  INV_X1 U7464 ( .A(n5874), .ZN(n5859) );
  AND2_X1 U7465 ( .A1(n5873), .A2(n5859), .ZN(n5860) );
  NAND2_X1 U7466 ( .A1(n7897), .A2(n5860), .ZN(n5870) );
  INV_X1 U7467 ( .A(n5861), .ZN(n5868) );
  INV_X1 U7468 ( .A(n5862), .ZN(n5867) );
  INV_X1 U7469 ( .A(n5863), .ZN(n5864) );
  INV_X1 U7470 ( .A(n7938), .ZN(n8123) );
  NAND2_X1 U7471 ( .A1(n5864), .A2(n8123), .ZN(n5865) );
  AND2_X1 U7472 ( .A1(n7899), .A2(n6376), .ZN(n5866) );
  OR2_X1 U7473 ( .A1(n5874), .A2(n5871), .ZN(n5869) );
  NAND2_X1 U7474 ( .A1(n5880), .A2(n5876), .ZN(n5878) );
  NAND3_X1 U7475 ( .A1(n5882), .A2(n6439), .A3(n5891), .ZN(n5877) );
  NAND2_X1 U7476 ( .A1(n5878), .A2(n5877), .ZN(n7954) );
  NAND2_X1 U7477 ( .A1(n5880), .A2(n9835), .ZN(n5881) );
  NOR2_X1 U7478 ( .A1(n9819), .A2(n7808), .ZN(n6360) );
  NAND2_X1 U7479 ( .A1(n6439), .A2(n6360), .ZN(n7377) );
  NAND2_X1 U7480 ( .A1(n5881), .A2(n7377), .ZN(n7973) );
  NAND2_X1 U7481 ( .A1(n8257), .A2(n7973), .ZN(n5901) );
  INV_X1 U7482 ( .A(n5882), .ZN(n5894) );
  AND2_X1 U7483 ( .A1(n6439), .A2(n5883), .ZN(n7815) );
  NAND2_X1 U7484 ( .A1(n7815), .A2(n5885), .ZN(n5884) );
  INV_X1 U7485 ( .A(n5885), .ZN(n5886) );
  NAND2_X1 U7486 ( .A1(n7815), .A2(n5886), .ZN(n5887) );
  NAND2_X1 U7487 ( .A1(n8094), .A2(n7968), .ZN(n5898) );
  NAND2_X1 U7488 ( .A1(n5889), .A2(n5888), .ZN(n5893) );
  NAND2_X1 U7489 ( .A1(n5774), .A2(n7732), .ZN(n6356) );
  NAND2_X1 U7490 ( .A1(n6417), .A2(n6356), .ZN(n5890) );
  AOI21_X1 U7491 ( .B1(n5894), .B2(n5891), .A(n5890), .ZN(n5892) );
  NAND2_X1 U7492 ( .A1(n5893), .A2(n5892), .ZN(n6546) );
  NAND2_X1 U7493 ( .A1(n6546), .A2(P2_STATE_REG_SCAN_IN), .ZN(n5896) );
  NAND2_X1 U7494 ( .A1(n5894), .A2(n7815), .ZN(n6547) );
  INV_X1 U7495 ( .A(n6403), .ZN(n6416) );
  NAND2_X1 U7496 ( .A1(n6416), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7819) );
  AND2_X1 U7497 ( .A1(n6547), .A2(n7819), .ZN(n5895) );
  NAND2_X2 U7498 ( .A1(n5896), .A2(n5895), .ZN(n7987) );
  AOI22_X1 U7499 ( .A1(n8096), .A2(n7987), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        n9917), .ZN(n5897) );
  OAI211_X1 U7500 ( .C1(n7904), .C2(n7971), .A(n5898), .B(n5897), .ZN(n5899)
         );
  INV_X1 U7501 ( .A(n5899), .ZN(n5900) );
  NAND2_X1 U7502 ( .A1(n5959), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n5908) );
  NAND2_X1 U7503 ( .A1(n4362), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n5907) );
  INV_X1 U7504 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n5905) );
  NAND2_X1 U7505 ( .A1(n8735), .A2(n6854), .ZN(n6890) );
  INV_X1 U7506 ( .A(n6890), .ZN(n5910) );
  NAND2_X1 U7507 ( .A1(n6893), .A2(n8738), .ZN(n5911) );
  NAND2_X1 U7508 ( .A1(n8735), .A2(n8730), .ZN(n8588) );
  NAND2_X1 U7509 ( .A1(n5911), .A2(n8588), .ZN(n5912) );
  NAND2_X4 U7510 ( .A1(n6408), .A2(n5912), .ZN(n6285) );
  NAND2_X1 U7511 ( .A1(n6892), .A2(n6890), .ZN(n5913) );
  NAND2_X4 U7512 ( .A1(n6408), .A2(n5914), .ZN(n6325) );
  AND2_X1 U7513 ( .A1(n9519), .A2(n6307), .ZN(n5915) );
  INV_X1 U7514 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n9620) );
  OR2_X1 U7515 ( .A1(n6408), .A2(n9620), .ZN(n5916) );
  NAND2_X1 U7516 ( .A1(n8756), .A2(n6287), .ZN(n5919) );
  INV_X1 U7517 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n6686) );
  NOR2_X1 U7518 ( .A1(n6408), .A2(n6686), .ZN(n5917) );
  AOI21_X1 U7519 ( .B1(n9519), .B2(n6323), .A(n5917), .ZN(n5918) );
  NAND2_X1 U7520 ( .A1(n5919), .A2(n5918), .ZN(n6627) );
  NAND2_X1 U7521 ( .A1(n6628), .A2(n6627), .ZN(n5922) );
  NAND2_X1 U7522 ( .A1(n5920), .A2(n6321), .ZN(n5921) );
  NAND2_X1 U7523 ( .A1(n4359), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n5926) );
  NAND2_X1 U7524 ( .A1(n5959), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5924) );
  NAND2_X1 U7525 ( .A1(n4361), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n5923) );
  INV_X2 U7526 ( .A(n4917), .ZN(n6323) );
  NAND2_X1 U7527 ( .A1(n6898), .A2(n6323), .ZN(n5927) );
  INV_X1 U7528 ( .A(n5931), .ZN(n5929) );
  INV_X1 U7529 ( .A(n5930), .ZN(n5928) );
  NAND2_X1 U7530 ( .A1(n5929), .A2(n5928), .ZN(n5932) );
  NAND2_X1 U7531 ( .A1(n5931), .A2(n5930), .ZN(n6708) );
  NAND2_X1 U7532 ( .A1(n4360), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5936) );
  NAND2_X1 U7533 ( .A1(n5933), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5935) );
  NAND2_X1 U7534 ( .A1(n4363), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n5934) );
  NAND2_X2 U7535 ( .A1(n5938), .A2(n5937), .ZN(n8754) );
  NAND2_X1 U7536 ( .A1(n8754), .A2(n6323), .ZN(n5940) );
  NAND2_X1 U7537 ( .A1(n9527), .A2(n6307), .ZN(n5939) );
  NAND2_X1 U7538 ( .A1(n5940), .A2(n5939), .ZN(n5941) );
  XNOR2_X1 U7539 ( .A(n5941), .B(n6321), .ZN(n5942) );
  AOI22_X1 U7540 ( .A1(n8754), .A2(n6287), .B1(n9527), .B2(n6323), .ZN(n5943)
         );
  NAND2_X1 U7541 ( .A1(n5942), .A2(n5943), .ZN(n5948) );
  INV_X1 U7542 ( .A(n5942), .ZN(n5945) );
  INV_X1 U7543 ( .A(n5943), .ZN(n5944) );
  NAND2_X1 U7544 ( .A1(n5945), .A2(n5944), .ZN(n5946) );
  AND2_X1 U7545 ( .A1(n5948), .A2(n5946), .ZN(n6710) );
  NAND2_X1 U7546 ( .A1(n6712), .A2(n5948), .ZN(n6824) );
  INV_X1 U7547 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n5950) );
  NAND2_X1 U7548 ( .A1(n5959), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5949) );
  OAI21_X1 U7549 ( .B1(n5904), .B2(n5950), .A(n5949), .ZN(n5951) );
  INV_X1 U7550 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n6826) );
  NAND2_X1 U7551 ( .A1(n4363), .A2(n6826), .ZN(n5952) );
  OAI22_X1 U7552 ( .A1(n6896), .A2(n4354), .B1(n6974), .B2(n6284), .ZN(n5955)
         );
  XNOR2_X1 U7553 ( .A(n5955), .B(n6321), .ZN(n5971) );
  OR2_X1 U7554 ( .A1(n6896), .A2(n6325), .ZN(n5957) );
  NAND2_X1 U7555 ( .A1(n9534), .A2(n6323), .ZN(n5956) );
  NAND2_X1 U7556 ( .A1(n5957), .A2(n5956), .ZN(n5969) );
  XNOR2_X1 U7557 ( .A(n5971), .B(n5969), .ZN(n6825) );
  NAND2_X1 U7558 ( .A1(n5933), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5965) );
  NAND2_X1 U7559 ( .A1(n5958), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5963) );
  NAND2_X1 U7560 ( .A1(n5959), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n5962) );
  INV_X1 U7561 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n6772) );
  NAND2_X1 U7562 ( .A1(n6826), .A2(n6772), .ZN(n5960) );
  AND2_X1 U7563 ( .A1(n5960), .A2(n5978), .ZN(n6977) );
  NAND2_X1 U7564 ( .A1(n4362), .A2(n6977), .ZN(n5961) );
  AND3_X1 U7565 ( .A1(n5963), .A2(n5962), .A3(n5961), .ZN(n5964) );
  OAI22_X1 U7566 ( .A1(n6970), .A2(n4354), .B1(n9541), .B2(n6284), .ZN(n5966)
         );
  XNOR2_X1 U7567 ( .A(n5966), .B(n6321), .ZN(n5973) );
  OR2_X1 U7568 ( .A1(n6970), .A2(n6325), .ZN(n5968) );
  NAND2_X1 U7569 ( .A1(n6978), .A2(n6323), .ZN(n5967) );
  NAND2_X1 U7570 ( .A1(n5968), .A2(n5967), .ZN(n5974) );
  XNOR2_X1 U7571 ( .A(n5973), .B(n5974), .ZN(n6770) );
  INV_X1 U7572 ( .A(n5969), .ZN(n5970) );
  NAND2_X1 U7573 ( .A1(n5971), .A2(n5970), .ZN(n6771) );
  AND2_X1 U7574 ( .A1(n6770), .A2(n6771), .ZN(n5972) );
  NAND2_X1 U7575 ( .A1(n6768), .A2(n5972), .ZN(n6767) );
  INV_X1 U7576 ( .A(n5973), .ZN(n5975) );
  NAND2_X1 U7577 ( .A1(n5975), .A2(n5974), .ZN(n5976) );
  NAND2_X1 U7578 ( .A1(n5933), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5983) );
  NAND2_X1 U7579 ( .A1(n5958), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n5982) );
  INV_X1 U7580 ( .A(n5978), .ZN(n5977) );
  NAND2_X1 U7581 ( .A1(n5977), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n5995) );
  INV_X1 U7582 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n6963) );
  NAND2_X1 U7583 ( .A1(n5978), .A2(n6963), .ZN(n5979) );
  AND2_X1 U7584 ( .A1(n5995), .A2(n5979), .ZN(n7053) );
  NAND2_X1 U7585 ( .A1(n4362), .A2(n7053), .ZN(n5981) );
  NAND2_X1 U7586 ( .A1(n5959), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n5980) );
  OAI22_X1 U7587 ( .A1(n7160), .A2(n4354), .B1(n9548), .B2(n6284), .ZN(n5984)
         );
  XNOR2_X1 U7588 ( .A(n5984), .B(n6285), .ZN(n5988) );
  NAND2_X1 U7589 ( .A1(n5987), .A2(n5988), .ZN(n6959) );
  OR2_X1 U7590 ( .A1(n7160), .A2(n6325), .ZN(n5986) );
  NAND2_X1 U7591 ( .A1(n7054), .A2(n6323), .ZN(n5985) );
  AND2_X1 U7592 ( .A1(n5986), .A2(n5985), .ZN(n6961) );
  NAND2_X1 U7593 ( .A1(n6959), .A2(n6961), .ZN(n5991) );
  INV_X1 U7594 ( .A(n5988), .ZN(n5989) );
  NAND2_X1 U7595 ( .A1(n5990), .A2(n5989), .ZN(n6960) );
  NAND2_X1 U7596 ( .A1(n5991), .A2(n6960), .ZN(n7066) );
  NAND2_X1 U7597 ( .A1(n5958), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5998) );
  INV_X1 U7598 ( .A(n5995), .ZN(n5993) );
  INV_X1 U7599 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n5994) );
  NAND2_X1 U7600 ( .A1(n5995), .A2(n5994), .ZN(n5996) );
  AND2_X1 U7601 ( .A1(n6010), .A2(n5996), .ZN(n9470) );
  NOR2_X1 U7602 ( .A1(n4900), .A2(n4902), .ZN(n5997) );
  NAND2_X1 U7603 ( .A1(n8578), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n5999) );
  INV_X1 U7604 ( .A(n9473), .ZN(n9554) );
  OAI22_X1 U7605 ( .A1(n7164), .A2(n4354), .B1(n9554), .B2(n6284), .ZN(n6000)
         );
  XNOR2_X1 U7606 ( .A(n6000), .B(n6321), .ZN(n6003) );
  OR2_X1 U7607 ( .A1(n7164), .A2(n6325), .ZN(n6002) );
  NAND2_X1 U7608 ( .A1(n9473), .A2(n6323), .ZN(n6001) );
  AND2_X1 U7609 ( .A1(n6002), .A2(n6001), .ZN(n6004) );
  NAND2_X1 U7610 ( .A1(n6003), .A2(n6004), .ZN(n7105) );
  INV_X1 U7611 ( .A(n6003), .ZN(n6006) );
  INV_X1 U7612 ( .A(n6004), .ZN(n6005) );
  NAND2_X1 U7613 ( .A1(n6006), .A2(n6005), .ZN(n6007) );
  AND2_X1 U7614 ( .A1(n7105), .A2(n6007), .ZN(n7067) );
  NAND2_X1 U7615 ( .A1(n8578), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6015) );
  NAND2_X1 U7616 ( .A1(n5958), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n6014) );
  INV_X1 U7617 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n6009) );
  NAND2_X1 U7618 ( .A1(n6010), .A2(n6009), .ZN(n6011) );
  AND2_X1 U7619 ( .A1(n6027), .A2(n6011), .ZN(n7112) );
  NAND2_X1 U7620 ( .A1(n4362), .A2(n7112), .ZN(n6013) );
  NAND2_X1 U7621 ( .A1(n5959), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n6012) );
  OAI22_X1 U7622 ( .A1(n8483), .A2(n4354), .B1(n9561), .B2(n6284), .ZN(n6016)
         );
  XNOR2_X1 U7623 ( .A(n6016), .B(n6321), .ZN(n6023) );
  INV_X1 U7624 ( .A(n6023), .ZN(n6020) );
  OR2_X1 U7625 ( .A1(n8483), .A2(n6325), .ZN(n6018) );
  NAND2_X1 U7626 ( .A1(n8491), .A2(n6323), .ZN(n6017) );
  AND2_X1 U7627 ( .A1(n6018), .A2(n6017), .ZN(n6022) );
  INV_X1 U7628 ( .A(n6022), .ZN(n6019) );
  NAND2_X1 U7629 ( .A1(n6020), .A2(n6019), .ZN(n6021) );
  AND2_X1 U7630 ( .A1(n7067), .A2(n6021), .ZN(n6025) );
  INV_X1 U7631 ( .A(n6021), .ZN(n7110) );
  AND2_X1 U7632 ( .A1(n6023), .A2(n6022), .ZN(n7108) );
  INV_X1 U7633 ( .A(n7108), .ZN(n6024) );
  AND2_X1 U7634 ( .A1(n6024), .A2(n7105), .ZN(n7104) );
  AOI21_X2 U7635 ( .B1(n7066), .B2(n6025), .A(n4898), .ZN(n6036) );
  NAND2_X1 U7636 ( .A1(n5958), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n6032) );
  NAND2_X1 U7637 ( .A1(n5959), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6031) );
  NAND2_X1 U7638 ( .A1(n6027), .A2(n6026), .ZN(n6028) );
  AND2_X1 U7639 ( .A1(n6042), .A2(n6028), .ZN(n7255) );
  NAND2_X1 U7640 ( .A1(n4363), .A2(n7255), .ZN(n6030) );
  NAND2_X1 U7641 ( .A1(n8578), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6029) );
  OAI22_X1 U7642 ( .A1(n8490), .A2(n4354), .B1(n9567), .B2(n6284), .ZN(n6033)
         );
  XNOR2_X1 U7643 ( .A(n6033), .B(n6321), .ZN(n6037) );
  XNOR2_X1 U7644 ( .A(n6036), .B(n6037), .ZN(n7249) );
  OR2_X1 U7645 ( .A1(n8490), .A2(n6325), .ZN(n6035) );
  NAND2_X1 U7646 ( .A1(n8486), .A2(n6323), .ZN(n6034) );
  AND2_X1 U7647 ( .A1(n6035), .A2(n6034), .ZN(n7251) );
  INV_X1 U7648 ( .A(n6037), .ZN(n6038) );
  NAND2_X1 U7649 ( .A1(n5958), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n6047) );
  NAND2_X1 U7650 ( .A1(n8578), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6046) );
  INV_X1 U7651 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n6041) );
  NAND2_X1 U7652 ( .A1(n6042), .A2(n6041), .ZN(n6043) );
  AND2_X1 U7653 ( .A1(n6067), .A2(n6043), .ZN(n7339) );
  NAND2_X1 U7654 ( .A1(n4363), .A2(n7339), .ZN(n6045) );
  NAND2_X1 U7655 ( .A1(n5959), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6044) );
  INV_X1 U7656 ( .A(n7343), .ZN(n9576) );
  OAI22_X1 U7657 ( .A1(n7471), .A2(n4354), .B1(n9576), .B2(n6284), .ZN(n6048)
         );
  XNOR2_X1 U7658 ( .A(n6048), .B(n6321), .ZN(n6053) );
  OR2_X1 U7659 ( .A1(n7471), .A2(n6325), .ZN(n6050) );
  NAND2_X1 U7660 ( .A1(n7343), .A2(n6323), .ZN(n6049) );
  NAND2_X1 U7661 ( .A1(n6050), .A2(n6049), .ZN(n6051) );
  XNOR2_X1 U7662 ( .A(n6053), .B(n6051), .ZN(n7338) );
  INV_X1 U7663 ( .A(n6051), .ZN(n6052) );
  NAND2_X1 U7664 ( .A1(n9590), .A2(n6307), .ZN(n6062) );
  NAND2_X1 U7665 ( .A1(n5958), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n6060) );
  NAND2_X1 U7666 ( .A1(n5959), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6059) );
  INV_X1 U7667 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n6066) );
  INV_X1 U7668 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n6055) );
  NAND2_X1 U7669 ( .A1(n6069), .A2(n6055), .ZN(n6056) );
  AND2_X1 U7670 ( .A1(n6086), .A2(n6056), .ZN(n7536) );
  NAND2_X1 U7671 ( .A1(n4363), .A2(n7536), .ZN(n6058) );
  NAND2_X1 U7672 ( .A1(n8578), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n6057) );
  OR2_X1 U7673 ( .A1(n7472), .A2(n4354), .ZN(n6061) );
  NAND2_X1 U7674 ( .A1(n6062), .A2(n6061), .ZN(n6063) );
  XNOR2_X1 U7675 ( .A(n6063), .B(n6285), .ZN(n6079) );
  NAND2_X1 U7676 ( .A1(n9590), .A2(n6323), .ZN(n6065) );
  OR2_X1 U7677 ( .A1(n7472), .A2(n6325), .ZN(n6064) );
  NAND2_X1 U7678 ( .A1(n6065), .A2(n6064), .ZN(n7532) );
  NAND2_X1 U7679 ( .A1(n5958), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n6073) );
  NAND2_X1 U7680 ( .A1(n5959), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6072) );
  NAND2_X1 U7681 ( .A1(n6067), .A2(n6066), .ZN(n6068) );
  AND2_X1 U7682 ( .A1(n6069), .A2(n6068), .ZN(n7266) );
  NAND2_X1 U7683 ( .A1(n4362), .A2(n7266), .ZN(n6071) );
  NAND2_X1 U7684 ( .A1(n8578), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n6070) );
  OR2_X1 U7685 ( .A1(n8750), .A2(n6325), .ZN(n6075) );
  NAND2_X1 U7686 ( .A1(n7475), .A2(n6323), .ZN(n6074) );
  NAND2_X1 U7687 ( .A1(n6075), .A2(n6074), .ZN(n7468) );
  NAND2_X1 U7688 ( .A1(n7475), .A2(n6307), .ZN(n6076) );
  OAI21_X1 U7689 ( .B1(n8750), .B2(n4354), .A(n6076), .ZN(n6077) );
  XNOR2_X1 U7690 ( .A(n6077), .B(n6285), .ZN(n6080) );
  AOI22_X1 U7691 ( .A1(n6079), .A2(n7532), .B1(n7468), .B2(n6080), .ZN(n6078)
         );
  NAND2_X1 U7692 ( .A1(n7467), .A2(n6078), .ZN(n6084) );
  OAI21_X1 U7693 ( .B1(n6080), .B2(n7468), .A(n7532), .ZN(n6082) );
  INV_X1 U7694 ( .A(n6079), .ZN(n7533) );
  INV_X1 U7695 ( .A(n6080), .ZN(n7531) );
  NOR2_X1 U7696 ( .A1(n7532), .A2(n7468), .ZN(n6081) );
  AOI22_X1 U7697 ( .A1(n6082), .A2(n7533), .B1(n7531), .B2(n6081), .ZN(n6083)
         );
  NAND2_X1 U7698 ( .A1(n6084), .A2(n6083), .ZN(n7459) );
  NAND2_X1 U7699 ( .A1(n8578), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n6091) );
  NAND2_X1 U7700 ( .A1(n5958), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n6090) );
  INV_X1 U7701 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n6085) );
  NAND2_X1 U7702 ( .A1(n6086), .A2(n6085), .ZN(n6087) );
  AND2_X1 U7703 ( .A1(n6098), .A2(n6087), .ZN(n7404) );
  NAND2_X1 U7704 ( .A1(n4362), .A2(n7404), .ZN(n6089) );
  NAND2_X1 U7705 ( .A1(n5959), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n6088) );
  NAND4_X1 U7706 ( .A1(n6091), .A2(n6090), .A3(n6089), .A4(n6088), .ZN(n8748)
         );
  OAI22_X1 U7707 ( .A1(n9601), .A2(n6284), .B1(n7538), .B2(n4354), .ZN(n6092)
         );
  XNOR2_X1 U7708 ( .A(n6092), .B(n6321), .ZN(n6095) );
  OAI22_X1 U7709 ( .A1(n9601), .A2(n4354), .B1(n7538), .B2(n6325), .ZN(n6093)
         );
  XNOR2_X1 U7710 ( .A(n6095), .B(n6093), .ZN(n7460) );
  INV_X1 U7711 ( .A(n6093), .ZN(n6094) );
  NAND2_X1 U7712 ( .A1(n6095), .A2(n6094), .ZN(n6096) );
  NAND2_X1 U7713 ( .A1(n8578), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n6103) );
  NAND2_X1 U7714 ( .A1(n5958), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n6102) );
  INV_X1 U7715 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n6097) );
  NAND2_X1 U7716 ( .A1(n6098), .A2(n6097), .ZN(n6099) );
  AND2_X1 U7717 ( .A1(n6110), .A2(n6099), .ZN(n7488) );
  NAND2_X1 U7718 ( .A1(n4363), .A2(n7488), .ZN(n6101) );
  NAND2_X1 U7719 ( .A1(n5959), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n6100) );
  OAI22_X1 U7720 ( .A1(n9607), .A2(n6284), .B1(n7559), .B2(n4354), .ZN(n6104)
         );
  XNOR2_X1 U7721 ( .A(n6104), .B(n6321), .ZN(n6105) );
  OAI22_X1 U7722 ( .A1(n9607), .A2(n4354), .B1(n7559), .B2(n6325), .ZN(n6106)
         );
  XNOR2_X1 U7723 ( .A(n6105), .B(n6106), .ZN(n7498) );
  INV_X1 U7724 ( .A(n6105), .ZN(n6107) );
  NAND2_X1 U7725 ( .A1(n5958), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n6115) );
  NAND2_X1 U7726 ( .A1(n5959), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n6114) );
  INV_X1 U7727 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n6109) );
  NAND2_X1 U7728 ( .A1(n6110), .A2(n6109), .ZN(n6111) );
  AND2_X1 U7729 ( .A1(n6134), .A2(n6111), .ZN(n7587) );
  NAND2_X1 U7730 ( .A1(n4363), .A2(n7587), .ZN(n6113) );
  NAND2_X1 U7731 ( .A1(n8578), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n6112) );
  OAI22_X1 U7732 ( .A1(n9614), .A2(n6284), .B1(n7568), .B2(n4354), .ZN(n6116)
         );
  XNOR2_X1 U7733 ( .A(n6116), .B(n6321), .ZN(n6119) );
  XNOR2_X1 U7734 ( .A(n6120), .B(n6119), .ZN(n8331) );
  INV_X1 U7735 ( .A(n8331), .ZN(n6118) );
  OAI22_X1 U7736 ( .A1(n9614), .A2(n4354), .B1(n7568), .B2(n6325), .ZN(n8334)
         );
  NAND2_X1 U7737 ( .A1(n6118), .A2(n6117), .ZN(n8332) );
  NAND2_X1 U7738 ( .A1(n6120), .A2(n6119), .ZN(n6121) );
  NAND2_X1 U7739 ( .A1(n8332), .A2(n6121), .ZN(n8374) );
  NAND2_X1 U7740 ( .A1(n9083), .A2(n6307), .ZN(n6129) );
  NAND2_X1 U7741 ( .A1(n8578), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n6127) );
  NAND2_X1 U7742 ( .A1(n5958), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n6126) );
  INV_X1 U7743 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n8382) );
  NAND2_X1 U7744 ( .A1(n6136), .A2(n8382), .ZN(n6123) );
  AND2_X1 U7745 ( .A1(n6152), .A2(n6123), .ZN(n9080) );
  NAND2_X1 U7746 ( .A1(n4362), .A2(n9080), .ZN(n6125) );
  NAND2_X1 U7747 ( .A1(n5959), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n6124) );
  OR2_X1 U7748 ( .A1(n9061), .A2(n4354), .ZN(n6128) );
  NAND2_X1 U7749 ( .A1(n6129), .A2(n6128), .ZN(n6130) );
  XNOR2_X1 U7750 ( .A(n6130), .B(n6285), .ZN(n8378) );
  NAND2_X1 U7751 ( .A1(n9083), .A2(n6323), .ZN(n6132) );
  OR2_X1 U7752 ( .A1(n9061), .A2(n6325), .ZN(n6131) );
  NAND2_X1 U7753 ( .A1(n6132), .A2(n6131), .ZN(n8377) );
  OR2_X1 U7754 ( .A1(n9295), .A2(n4354), .ZN(n6142) );
  INV_X1 U7755 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n6133) );
  NAND2_X1 U7756 ( .A1(n6134), .A2(n6133), .ZN(n6135) );
  AND2_X1 U7757 ( .A1(n6136), .A2(n6135), .ZN(n7577) );
  NAND2_X1 U7758 ( .A1(n4363), .A2(n7577), .ZN(n6140) );
  NAND2_X1 U7759 ( .A1(n5958), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n6139) );
  NAND2_X1 U7760 ( .A1(n5959), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n6138) );
  NAND2_X1 U7761 ( .A1(n8578), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n6137) );
  OR2_X1 U7762 ( .A1(n8384), .A2(n6325), .ZN(n6141) );
  NAND2_X1 U7763 ( .A1(n6142), .A2(n6141), .ZN(n8452) );
  OAI22_X1 U7764 ( .A1(n9295), .A2(n6284), .B1(n8384), .B2(n4354), .ZN(n6143)
         );
  XNOR2_X1 U7765 ( .A(n6143), .B(n6285), .ZN(n8375) );
  OAI22_X1 U7766 ( .A1(n8378), .A2(n8377), .B1(n8452), .B2(n8375), .ZN(n6149)
         );
  NAND2_X1 U7767 ( .A1(n8375), .A2(n8452), .ZN(n6145) );
  INV_X1 U7768 ( .A(n8377), .ZN(n6144) );
  NAND2_X1 U7769 ( .A1(n6145), .A2(n6144), .ZN(n6147) );
  INV_X1 U7770 ( .A(n6145), .ZN(n6146) );
  AOI22_X1 U7771 ( .A1(n8378), .A2(n6147), .B1(n6146), .B2(n8377), .ZN(n6148)
         );
  OAI21_X2 U7772 ( .B1(n8374), .B2(n6149), .A(n6148), .ZN(n8392) );
  NAND2_X1 U7773 ( .A1(n5958), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n6157) );
  NAND2_X1 U7774 ( .A1(n5959), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n6156) );
  INV_X1 U7775 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n6151) );
  NAND2_X1 U7776 ( .A1(n6152), .A2(n6151), .ZN(n6153) );
  AND2_X1 U7777 ( .A1(n6174), .A2(n6153), .ZN(n9064) );
  NAND2_X1 U7778 ( .A1(n4362), .A2(n9064), .ZN(n6155) );
  NAND2_X1 U7779 ( .A1(n8578), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n6154) );
  OAI22_X1 U7780 ( .A1(n9068), .A2(n6284), .B1(n8383), .B2(n4354), .ZN(n6158)
         );
  XNOR2_X1 U7781 ( .A(n6158), .B(n6285), .ZN(n6160) );
  OAI22_X1 U7782 ( .A1(n9068), .A2(n4354), .B1(n8383), .B2(n6325), .ZN(n6159)
         );
  AND2_X1 U7783 ( .A1(n6160), .A2(n6159), .ZN(n8389) );
  OR2_X1 U7784 ( .A1(n6160), .A2(n6159), .ZN(n8388) );
  NAND2_X1 U7785 ( .A1(n9148), .A2(n6307), .ZN(n6169) );
  NAND2_X1 U7786 ( .A1(n8578), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n6167) );
  NAND2_X1 U7787 ( .A1(n5958), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n6166) );
  INV_X1 U7788 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n6173) );
  INV_X1 U7789 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n6162) );
  NAND2_X1 U7790 ( .A1(n6176), .A2(n6162), .ZN(n6163) );
  AND2_X1 U7791 ( .A1(n6192), .A2(n6163), .ZN(n9023) );
  NAND2_X1 U7792 ( .A1(n4362), .A2(n9023), .ZN(n6165) );
  NAND2_X1 U7793 ( .A1(n5959), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n6164) );
  NAND4_X1 U7794 ( .A1(n6167), .A2(n6166), .A3(n6165), .A4(n6164), .ZN(n9047)
         );
  NAND2_X1 U7795 ( .A1(n9047), .A2(n6323), .ZN(n6168) );
  NAND2_X1 U7796 ( .A1(n6169), .A2(n6168), .ZN(n6170) );
  XNOR2_X1 U7797 ( .A(n6170), .B(n6285), .ZN(n8352) );
  NAND2_X1 U7798 ( .A1(n9148), .A2(n6323), .ZN(n6172) );
  NAND2_X1 U7799 ( .A1(n9047), .A2(n6287), .ZN(n6171) );
  NAND2_X1 U7800 ( .A1(n6172), .A2(n6171), .ZN(n8351) );
  NAND2_X1 U7801 ( .A1(n9154), .A2(n6323), .ZN(n6182) );
  NAND2_X1 U7802 ( .A1(n8578), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n6180) );
  NAND2_X1 U7803 ( .A1(n5958), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n6179) );
  NAND2_X1 U7804 ( .A1(n6174), .A2(n6173), .ZN(n6175) );
  AND2_X1 U7805 ( .A1(n6176), .A2(n6175), .ZN(n9041) );
  NAND2_X1 U7806 ( .A1(n4363), .A2(n9041), .ZN(n6178) );
  NAND2_X1 U7807 ( .A1(n5959), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n6177) );
  NAND4_X1 U7808 ( .A1(n6180), .A2(n6179), .A3(n6178), .A4(n6177), .ZN(n9034)
         );
  NAND2_X1 U7809 ( .A1(n9034), .A2(n6287), .ZN(n6181) );
  NAND2_X1 U7810 ( .A1(n6182), .A2(n6181), .ZN(n8434) );
  NAND2_X1 U7811 ( .A1(n9154), .A2(n6307), .ZN(n6184) );
  NAND2_X1 U7812 ( .A1(n9034), .A2(n6323), .ZN(n6183) );
  NAND2_X1 U7813 ( .A1(n6184), .A2(n6183), .ZN(n6185) );
  XNOR2_X1 U7814 ( .A(n6185), .B(n6285), .ZN(n8349) );
  OAI22_X1 U7815 ( .A1(n8352), .A2(n8351), .B1(n8434), .B2(n8349), .ZN(n6191)
         );
  NAND2_X1 U7816 ( .A1(n8349), .A2(n8434), .ZN(n6187) );
  INV_X1 U7817 ( .A(n8351), .ZN(n6186) );
  NAND2_X1 U7818 ( .A1(n6187), .A2(n6186), .ZN(n6189) );
  INV_X1 U7819 ( .A(n6187), .ZN(n6188) );
  AOI22_X1 U7820 ( .A1(n8352), .A2(n6189), .B1(n6188), .B2(n8351), .ZN(n6190)
         );
  OAI21_X2 U7821 ( .B1(n8348), .B2(n6191), .A(n6190), .ZN(n8411) );
  NAND2_X1 U7822 ( .A1(n5958), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n6197) );
  NAND2_X1 U7823 ( .A1(n5959), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n6196) );
  INV_X1 U7824 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n8412) );
  NAND2_X1 U7825 ( .A1(n6192), .A2(n8412), .ZN(n6193) );
  AND2_X1 U7826 ( .A1(n6208), .A2(n6193), .ZN(n9014) );
  NAND2_X1 U7827 ( .A1(n4362), .A2(n9014), .ZN(n6195) );
  NAND2_X1 U7828 ( .A1(n8578), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n6194) );
  OAI22_X1 U7829 ( .A1(n9017), .A2(n6284), .B1(n9026), .B2(n4354), .ZN(n6198)
         );
  XNOR2_X1 U7830 ( .A(n6198), .B(n6321), .ZN(n8409) );
  OR2_X1 U7831 ( .A1(n9017), .A2(n4354), .ZN(n6200) );
  OR2_X1 U7832 ( .A1(n9026), .A2(n6325), .ZN(n6199) );
  NAND2_X1 U7833 ( .A1(n8409), .A2(n6202), .ZN(n6201) );
  INV_X1 U7834 ( .A(n8409), .ZN(n6203) );
  INV_X1 U7835 ( .A(n6202), .ZN(n8408) );
  NAND2_X1 U7836 ( .A1(n6203), .A2(n8408), .ZN(n6204) );
  NAND2_X1 U7837 ( .A1(n9140), .A2(n6307), .ZN(n6213) );
  INV_X1 U7838 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n8993) );
  NAND2_X1 U7839 ( .A1(n5958), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n6206) );
  NAND2_X1 U7840 ( .A1(n8578), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n6205) );
  AND2_X1 U7841 ( .A1(n6206), .A2(n6205), .ZN(n6211) );
  INV_X1 U7842 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n8361) );
  NAND2_X1 U7843 ( .A1(n6208), .A2(n8361), .ZN(n6209) );
  NAND2_X1 U7844 ( .A1(n6233), .A2(n6209), .ZN(n8992) );
  INV_X1 U7845 ( .A(n4363), .ZN(n6265) );
  OR2_X1 U7846 ( .A1(n8992), .A2(n6265), .ZN(n6210) );
  OAI211_X1 U7847 ( .C1(n6337), .C2(n8993), .A(n6211), .B(n6210), .ZN(n8745)
         );
  NAND2_X1 U7848 ( .A1(n8745), .A2(n6323), .ZN(n6212) );
  NAND2_X1 U7849 ( .A1(n6213), .A2(n6212), .ZN(n6214) );
  XNOR2_X1 U7850 ( .A(n6214), .B(n6321), .ZN(n6217) );
  AND2_X1 U7851 ( .A1(n8745), .A2(n6287), .ZN(n6215) );
  AOI21_X1 U7852 ( .B1(n9140), .B2(n6323), .A(n6215), .ZN(n6216) );
  XNOR2_X1 U7853 ( .A(n6217), .B(n6216), .ZN(n8360) );
  NAND2_X1 U7854 ( .A1(n9135), .A2(n6307), .ZN(n6225) );
  XNOR2_X1 U7855 ( .A(n6233), .B(P1_REG3_REG_22__SCAN_IN), .ZN(n8982) );
  NAND2_X1 U7856 ( .A1(n8982), .A2(n4362), .ZN(n6223) );
  INV_X1 U7857 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n6220) );
  NAND2_X1 U7858 ( .A1(n8578), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n6219) );
  NAND2_X1 U7859 ( .A1(n4360), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n6218) );
  OAI211_X1 U7860 ( .C1(n6220), .C2(n6337), .A(n6219), .B(n6218), .ZN(n6221)
         );
  INV_X1 U7861 ( .A(n6221), .ZN(n6222) );
  NAND2_X1 U7862 ( .A1(n6223), .A2(n6222), .ZN(n8744) );
  NAND2_X1 U7863 ( .A1(n8744), .A2(n6323), .ZN(n6224) );
  NAND2_X1 U7864 ( .A1(n6225), .A2(n6224), .ZN(n6226) );
  XNOR2_X1 U7865 ( .A(n6226), .B(n6321), .ZN(n6229) );
  NAND2_X1 U7866 ( .A1(n9135), .A2(n6323), .ZN(n6228) );
  NAND2_X1 U7867 ( .A1(n8744), .A2(n6287), .ZN(n6227) );
  NAND2_X1 U7868 ( .A1(n6228), .A2(n6227), .ZN(n8421) );
  AND2_X2 U7869 ( .A1(n6230), .A2(n6229), .ZN(n8418) );
  INV_X1 U7870 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n8424) );
  INV_X1 U7871 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n6231) );
  OAI21_X1 U7872 ( .B1(n6233), .B2(n8424), .A(n6231), .ZN(n6234) );
  NAND2_X1 U7873 ( .A1(P1_REG3_REG_22__SCAN_IN), .A2(P1_REG3_REG_23__SCAN_IN), 
        .ZN(n6232) );
  NAND2_X1 U7874 ( .A1(n6234), .A2(n6248), .ZN(n8967) );
  OR2_X1 U7875 ( .A1(n8967), .A2(n6265), .ZN(n6237) );
  AOI22_X1 U7876 ( .A1(n8578), .A2(P1_REG1_REG_23__SCAN_IN), .B1(n5958), .B2(
        P1_REG0_REG_23__SCAN_IN), .ZN(n6236) );
  NAND2_X1 U7877 ( .A1(n5959), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n6235) );
  OAI22_X1 U7878 ( .A1(n8971), .A2(n6284), .B1(n8980), .B2(n4354), .ZN(n6238)
         );
  XNOR2_X1 U7879 ( .A(n6238), .B(n6321), .ZN(n6241) );
  OR2_X1 U7880 ( .A1(n8971), .A2(n4354), .ZN(n6240) );
  INV_X1 U7881 ( .A(n8980), .ZN(n8743) );
  NAND2_X1 U7882 ( .A1(n8743), .A2(n6287), .ZN(n6239) );
  NAND2_X1 U7883 ( .A1(n6241), .A2(n6242), .ZN(n8399) );
  INV_X1 U7884 ( .A(n6241), .ZN(n6244) );
  INV_X1 U7885 ( .A(n6242), .ZN(n6243) );
  NAND2_X1 U7886 ( .A1(n6244), .A2(n6243), .ZN(n6245) );
  OAI21_X2 U7887 ( .B1(n8423), .B2(n8418), .A(n8341), .ZN(n8400) );
  INV_X1 U7888 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n6247) );
  NAND2_X1 U7889 ( .A1(n6248), .A2(n6247), .ZN(n6249) );
  NAND2_X1 U7890 ( .A1(n6263), .A2(n6249), .ZN(n8953) );
  OR2_X1 U7891 ( .A1(n8953), .A2(n6265), .ZN(n6252) );
  AOI22_X1 U7892 ( .A1(n8578), .A2(P1_REG1_REG_24__SCAN_IN), .B1(n5958), .B2(
        P1_REG0_REG_24__SCAN_IN), .ZN(n6251) );
  NAND2_X1 U7893 ( .A1(n5959), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n6250) );
  OAI22_X1 U7894 ( .A1(n8957), .A2(n6284), .B1(n8964), .B2(n4354), .ZN(n6253)
         );
  XNOR2_X1 U7895 ( .A(n6253), .B(n6321), .ZN(n6256) );
  INV_X1 U7896 ( .A(n8964), .ZN(n8742) );
  NAND2_X1 U7897 ( .A1(n8742), .A2(n6287), .ZN(n6254) );
  NAND2_X1 U7898 ( .A1(n6256), .A2(n6257), .ZN(n6261) );
  INV_X1 U7899 ( .A(n6256), .ZN(n6259) );
  INV_X1 U7900 ( .A(n6257), .ZN(n6258) );
  NAND2_X1 U7901 ( .A1(n6259), .A2(n6258), .ZN(n6260) );
  NAND2_X1 U7902 ( .A1(n6261), .A2(n6260), .ZN(n8398) );
  INV_X1 U7903 ( .A(n6261), .ZN(n6262) );
  NAND2_X1 U7904 ( .A1(n9119), .A2(n6307), .ZN(n6273) );
  INV_X1 U7905 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n8368) );
  NAND2_X1 U7906 ( .A1(n6263), .A2(n8368), .ZN(n6264) );
  NAND2_X1 U7907 ( .A1(n6276), .A2(n6264), .ZN(n8369) );
  INV_X1 U7908 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n6268) );
  NAND2_X1 U7909 ( .A1(n8578), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n6267) );
  NAND2_X1 U7910 ( .A1(n4360), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n6266) );
  OAI211_X1 U7911 ( .C1(n6268), .C2(n6337), .A(n6267), .B(n6266), .ZN(n6269)
         );
  INV_X1 U7912 ( .A(n6269), .ZN(n6270) );
  NAND2_X1 U7913 ( .A1(n8938), .A2(n6323), .ZN(n6272) );
  NAND2_X1 U7914 ( .A1(n6273), .A2(n6272), .ZN(n6274) );
  XNOR2_X1 U7915 ( .A(n6274), .B(n6285), .ZN(n6291) );
  OAI22_X1 U7916 ( .A1(n8873), .A2(n4354), .B1(n8950), .B2(n6325), .ZN(n6290)
         );
  XNOR2_X1 U7917 ( .A(n6291), .B(n6290), .ZN(n8367) );
  INV_X1 U7918 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n6275) );
  NAND2_X1 U7919 ( .A1(n6276), .A2(n6275), .ZN(n6277) );
  NAND2_X1 U7920 ( .A1(n8932), .A2(n4362), .ZN(n6283) );
  INV_X1 U7921 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n6280) );
  NAND2_X1 U7922 ( .A1(n4360), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n6279) );
  NAND2_X1 U7923 ( .A1(n8578), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n6278) );
  OAI211_X1 U7924 ( .C1(n6280), .C2(n6337), .A(n6279), .B(n6278), .ZN(n6281)
         );
  INV_X1 U7925 ( .A(n6281), .ZN(n6282) );
  OAI22_X1 U7926 ( .A1(n8934), .A2(n6284), .B1(n8876), .B2(n4354), .ZN(n6286)
         );
  XNOR2_X1 U7927 ( .A(n6286), .B(n6285), .ZN(n6305) );
  OR2_X1 U7928 ( .A1(n8934), .A2(n4354), .ZN(n6289) );
  NAND2_X1 U7929 ( .A1(n8921), .A2(n6287), .ZN(n6288) );
  NAND2_X1 U7930 ( .A1(n6289), .A2(n6288), .ZN(n6304) );
  XNOR2_X1 U7931 ( .A(n6305), .B(n6304), .ZN(n8441) );
  NOR2_X1 U7932 ( .A1(n6291), .A2(n6290), .ZN(n8442) );
  NAND2_X1 U7933 ( .A1(n9109), .A2(n6307), .ZN(n6299) );
  XNOR2_X1 U7934 ( .A(n6311), .B(P1_REG3_REG_27__SCAN_IN), .ZN(n8914) );
  NAND2_X1 U7935 ( .A1(n8914), .A2(n4363), .ZN(n6297) );
  INV_X1 U7936 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n6294) );
  NAND2_X1 U7937 ( .A1(n4360), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n6293) );
  NAND2_X1 U7938 ( .A1(n8578), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n6292) );
  OAI211_X1 U7939 ( .C1(n6294), .C2(n6337), .A(n6293), .B(n6292), .ZN(n6295)
         );
  INV_X1 U7940 ( .A(n6295), .ZN(n6296) );
  NAND2_X1 U7941 ( .A1(n8939), .A2(n6323), .ZN(n6298) );
  NAND2_X1 U7942 ( .A1(n6299), .A2(n6298), .ZN(n6300) );
  XNOR2_X1 U7943 ( .A(n6300), .B(n6321), .ZN(n6303) );
  NOR2_X1 U7944 ( .A1(n8897), .A2(n6325), .ZN(n6301) );
  AOI21_X1 U7945 ( .B1(n9109), .B2(n6323), .A(n6301), .ZN(n6302) );
  NAND2_X1 U7946 ( .A1(n6303), .A2(n6302), .ZN(n6349) );
  OAI21_X1 U7947 ( .B1(n6303), .B2(n6302), .A(n6349), .ZN(n7601) );
  NAND2_X1 U7948 ( .A1(n9103), .A2(n6307), .ZN(n6320) );
  INV_X1 U7949 ( .A(n6311), .ZN(n6309) );
  AND2_X1 U7950 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .ZN(n6308) );
  NAND2_X1 U7951 ( .A1(n6309), .A2(n6308), .ZN(n8885) );
  INV_X1 U7952 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n7602) );
  INV_X1 U7953 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n6310) );
  OAI21_X1 U7954 ( .B1(n6311), .B2(n7602), .A(n6310), .ZN(n6312) );
  NAND2_X1 U7955 ( .A1(n8904), .A2(n4363), .ZN(n6318) );
  INV_X1 U7956 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n6315) );
  NAND2_X1 U7957 ( .A1(n5958), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n6314) );
  NAND2_X1 U7958 ( .A1(n8578), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n6313) );
  OAI211_X1 U7959 ( .C1(n6315), .C2(n6337), .A(n6314), .B(n6313), .ZN(n6316)
         );
  INV_X1 U7960 ( .A(n6316), .ZN(n6317) );
  OR2_X1 U7961 ( .A1(n8867), .A2(n4354), .ZN(n6319) );
  NAND2_X1 U7962 ( .A1(n6320), .A2(n6319), .ZN(n6322) );
  XNOR2_X1 U7963 ( .A(n6322), .B(n6321), .ZN(n6327) );
  NAND2_X1 U7964 ( .A1(n9103), .A2(n6323), .ZN(n6324) );
  OAI21_X1 U7965 ( .B1(n8867), .B2(n6325), .A(n6324), .ZN(n6326) );
  XNOR2_X1 U7966 ( .A(n6327), .B(n6326), .ZN(n6334) );
  INV_X1 U7967 ( .A(n6334), .ZN(n6350) );
  INV_X1 U7968 ( .A(n6328), .ZN(n6887) );
  NAND3_X1 U7969 ( .A1(n6330), .A2(n6887), .A3(n6329), .ZN(n6344) );
  INV_X1 U7970 ( .A(n6341), .ZN(n6332) );
  INV_X1 U7971 ( .A(n8622), .ZN(n6340) );
  AND2_X1 U7972 ( .A1(n6340), .A2(n9613), .ZN(n6331) );
  NAND3_X1 U7973 ( .A1(n6350), .A2(n8444), .A3(n6349), .ZN(n6333) );
  NAND3_X1 U7974 ( .A1(n7599), .A2(n6334), .A3(n8444), .ZN(n6354) );
  NOR2_X1 U7975 ( .A1(n9513), .A2(n6854), .ZN(n6910) );
  INV_X1 U7976 ( .A(n6910), .ZN(n9500) );
  INV_X1 U7977 ( .A(n8885), .ZN(n6339) );
  INV_X1 U7978 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n8884) );
  NAND2_X1 U7979 ( .A1(n8578), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n6336) );
  NAND2_X1 U7980 ( .A1(n4360), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n6335) );
  OAI211_X1 U7981 ( .C1(n8884), .C2(n6337), .A(n6336), .B(n6335), .ZN(n6338)
         );
  AOI21_X1 U7982 ( .B1(n6339), .B2(n4362), .A(n6338), .ZN(n8898) );
  OR2_X1 U7983 ( .A1(n6340), .A2(n6892), .ZN(n8655) );
  NOR2_X1 U7984 ( .A1(n6341), .A2(n8655), .ZN(n6342) );
  NAND2_X1 U7985 ( .A1(n6342), .A2(n5286), .ZN(n8427) );
  NAND2_X1 U7986 ( .A1(n6342), .A2(n8657), .ZN(n8426) );
  NAND2_X1 U7987 ( .A1(n8939), .A2(n8455), .ZN(n6348) );
  NAND2_X1 U7988 ( .A1(n6344), .A2(n6343), .ZN(n6630) );
  INV_X1 U7989 ( .A(n6345), .ZN(n6886) );
  NAND4_X1 U7990 ( .A1(n6630), .A2(n6486), .A3(n6408), .A4(n6886), .ZN(n6346)
         );
  INV_X1 U7991 ( .A(n8458), .ZN(n8446) );
  AOI22_X1 U7992 ( .A1(n8904), .A2(n8446), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3086), .ZN(n6347) );
  OAI211_X1 U7993 ( .C1(n8898), .C2(n8427), .A(n6348), .B(n6347), .ZN(n6352)
         );
  NOR3_X1 U7994 ( .A1(n6350), .A2(n8462), .A3(n6349), .ZN(n6351) );
  AOI211_X1 U7995 ( .C1(n9103), .C2(n8430), .A(n6352), .B(n6351), .ZN(n6353)
         );
  NAND3_X1 U7996 ( .A1(n6355), .A2(n6354), .A3(n6353), .ZN(P1_U3220) );
  NAND3_X1 U7997 ( .A1(n6357), .A2(n6439), .A3(n6356), .ZN(n6358) );
  NOR2_X1 U7998 ( .A1(n6359), .A2(n6358), .ZN(n6604) );
  INV_X1 U7999 ( .A(n6360), .ZN(n6363) );
  NAND2_X1 U8000 ( .A1(n6361), .A2(n7807), .ZN(n6362) );
  NAND2_X1 U8001 ( .A1(n6362), .A2(n7747), .ZN(n6364) );
  AOI21_X1 U8002 ( .B1(n5772), .B2(n6363), .A(n6364), .ZN(n6366) );
  INV_X1 U8003 ( .A(n6364), .ZN(n6601) );
  NOR2_X1 U8004 ( .A1(n6602), .A2(n6601), .ZN(n6365) );
  NOR2_X1 U8005 ( .A1(n6366), .A2(n6365), .ZN(n6367) );
  AND2_X2 U8006 ( .A1(n6604), .A2(n6367), .ZN(n9854) );
  NAND2_X1 U8007 ( .A1(n6368), .A2(n9854), .ZN(n6373) );
  NAND2_X1 U8008 ( .A1(n9854), .A2(n9835), .ZN(n8212) );
  NOR2_X1 U8009 ( .A1(n6369), .A2(n8212), .ZN(n6370) );
  NAND2_X1 U8010 ( .A1(n6373), .A2(n6372), .ZN(P2_U3488) );
  INV_X1 U8011 ( .A(n6375), .ZN(n6377) );
  NAND2_X1 U8012 ( .A1(n7897), .A2(n6378), .ZN(n6380) );
  OAI21_X1 U8013 ( .B1(n6382), .B2(n6381), .A(n7954), .ZN(n6389) );
  INV_X1 U8014 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n9942) );
  OAI22_X1 U8015 ( .A1(n7938), .A2(n7971), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9942), .ZN(n6384) );
  NOR2_X1 U8016 ( .A1(n8080), .A2(n7984), .ZN(n6383) );
  AOI211_X1 U8017 ( .C1(n8105), .C2(n7987), .A(n6384), .B(n6383), .ZN(n6385)
         );
  INV_X1 U8018 ( .A(n6387), .ZN(n6388) );
  NAND2_X1 U8019 ( .A1(n6389), .A2(n6388), .ZN(P2_U3180) );
  XNOR2_X1 U8020 ( .A(n8094), .B(n4357), .ZN(n6390) );
  XNOR2_X1 U8021 ( .A(n8086), .B(n6390), .ZN(n6391) );
  INV_X1 U8022 ( .A(n6391), .ZN(n6396) );
  OAI211_X1 U8023 ( .C1(n8080), .C2(n6395), .A(n6396), .B(n7954), .ZN(n6401)
         );
  AND2_X1 U8024 ( .A1(n6391), .A2(n7954), .ZN(n6392) );
  NAND2_X1 U8025 ( .A1(n6402), .A2(n6392), .ZN(n6400) );
  AOI22_X1 U8026 ( .A1(n8085), .A2(n7987), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        n9917), .ZN(n6394) );
  INV_X1 U8027 ( .A(n7971), .ZN(n7982) );
  NAND2_X1 U8028 ( .A1(n8102), .A2(n7982), .ZN(n6393) );
  OAI211_X1 U8029 ( .C1(n8081), .C2(n7984), .A(n6394), .B(n6393), .ZN(n6398)
         );
  NOR4_X1 U8030 ( .A1(n6396), .A2(n6395), .A3(n8080), .A4(n7977), .ZN(n6397)
         );
  AOI211_X1 U8031 ( .C1(n8086), .C2(n7973), .A(n6398), .B(n6397), .ZN(n6399)
         );
  OAI211_X1 U8032 ( .C1(n6402), .C2(n6401), .A(n6400), .B(n6399), .ZN(P2_U3160) );
  INV_X1 U8033 ( .A(n6548), .ZN(n6440) );
  OR2_X2 U8034 ( .A1(n6417), .A2(n6440), .ZN(n8005) );
  NAND2_X1 U8035 ( .A1(n6417), .A2(n7747), .ZN(n6404) );
  NAND2_X1 U8036 ( .A1(n6404), .A2(n6403), .ZN(n6411) );
  NAND2_X1 U8037 ( .A1(n6411), .A2(n5379), .ZN(n6405) );
  NAND2_X1 U8038 ( .A1(n6405), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3150) );
  INV_X1 U8039 ( .A(n6406), .ZN(n6407) );
  INV_X2 U8040 ( .A(n8755), .ZN(P1_U3973) );
  MUX2_X1 U8041 ( .A(P2_REG2_REG_1__SCAN_IN), .B(P2_REG1_REG_1__SCAN_IN), .S(
        n8057), .Z(n6524) );
  XOR2_X1 U8042 ( .A(n6421), .B(n6524), .Z(n6409) );
  MUX2_X1 U8043 ( .A(P2_REG2_REG_0__SCAN_IN), .B(P2_REG1_REG_0__SCAN_IN), .S(
        n8057), .Z(n6516) );
  NOR2_X1 U8044 ( .A1(n6516), .A2(n4709), .ZN(n6515) );
  AOI211_X1 U8045 ( .C1(n6409), .C2(n6515), .A(n4472), .B(n6522), .ZN(n6430)
         );
  NOR2_X1 U8046 ( .A1(n8057), .A2(n9917), .ZN(n7357) );
  NAND2_X1 U8047 ( .A1(n6411), .A2(n7357), .ZN(n6410) );
  MUX2_X1 U8048 ( .A(n8005), .B(n6410), .S(n5693), .Z(n9721) );
  INV_X1 U8049 ( .A(n6421), .ZN(n6523) );
  NOR2_X1 U8050 ( .A1(n9721), .A2(n6523), .ZN(n6429) );
  NOR2_X1 U8051 ( .A1(n5693), .A2(P2_U3151), .ZN(n7396) );
  NAND2_X1 U8052 ( .A1(n7396), .A2(n6411), .ZN(n6518) );
  OR2_X1 U8053 ( .A1(n6518), .A2(n6419), .ZN(n8066) );
  AND2_X1 U8054 ( .A1(n5385), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6529) );
  NAND2_X1 U8055 ( .A1(n4709), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6412) );
  OAI22_X1 U8056 ( .A1(n6529), .A2(n6421), .B1(n5385), .B2(n6412), .ZN(n6528)
         );
  INV_X1 U8057 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n6413) );
  XNOR2_X1 U8058 ( .A(n6528), .B(n6413), .ZN(n6415) );
  INV_X1 U8059 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n6414) );
  OAI22_X1 U8060 ( .A1(n8066), .A2(n6415), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6414), .ZN(n6428) );
  NOR2_X1 U8061 ( .A1(n6417), .A2(n6416), .ZN(n6418) );
  INV_X1 U8062 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n9858) );
  OR2_X1 U8063 ( .A1(n6518), .A2(n8046), .ZN(n9736) );
  INV_X1 U8064 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n6425) );
  NAND2_X1 U8065 ( .A1(n4709), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6420) );
  NAND2_X1 U8066 ( .A1(n6421), .A2(n6420), .ZN(n6422) );
  NAND2_X1 U8067 ( .A1(n5385), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6536) );
  NAND2_X1 U8068 ( .A1(n6422), .A2(n6536), .ZN(n6424) );
  OR2_X1 U8069 ( .A1(n6424), .A2(n6425), .ZN(n6537) );
  INV_X1 U8070 ( .A(n6537), .ZN(n6423) );
  AOI21_X1 U8071 ( .B1(n6425), .B2(n6424), .A(n6423), .ZN(n6426) );
  OAI22_X1 U8072 ( .A1(n9720), .A2(n9858), .B1(n9736), .B2(n6426), .ZN(n6427)
         );
  OR4_X1 U8073 ( .A1(n6430), .A2(n6429), .A3(n6428), .A4(n6427), .ZN(P2_U3183)
         );
  NAND2_X1 U8074 ( .A1(n6436), .A2(P1_U3086), .ZN(n7858) );
  AND2_X1 U8075 ( .A1(n4923), .A2(P1_U3086), .ZN(n7075) );
  INV_X2 U8076 ( .A(n7075), .ZN(n9193) );
  INV_X1 U8077 ( .A(n8763), .ZN(n6432) );
  OAI222_X1 U8078 ( .A1(n7858), .A2(n6433), .B1(n9193), .B2(n6454), .C1(
        P1_U3086), .C2(n6432), .ZN(P1_U3354) );
  INV_X1 U8079 ( .A(n8777), .ZN(n6434) );
  OAI222_X1 U8080 ( .A1(n7858), .A2(n6435), .B1(n9193), .B2(n6456), .C1(
        P1_U3086), .C2(n6434), .ZN(P1_U3353) );
  NOR2_X1 U8081 ( .A1(n6436), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8326) );
  INV_X1 U8082 ( .A(n8326), .ZN(n7118) );
  INV_X1 U8083 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6437) );
  NAND2_X1 U8084 ( .A1(n6436), .A2(n9917), .ZN(n6834) );
  OAI222_X1 U8085 ( .A1(n7118), .A2(n6437), .B1(n6834), .B2(n6450), .C1(
        P2_U3151), .C2(n6805), .ZN(P2_U3290) );
  OAI222_X1 U8086 ( .A1(n7118), .A2(n6438), .B1(n6834), .B2(n6452), .C1(n9917), 
        .C2(n6920), .ZN(P2_U3289) );
  NAND2_X1 U8087 ( .A1(n6439), .A2(n5739), .ZN(n6463) );
  INV_X1 U8088 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n6442) );
  NOR3_X1 U8089 ( .A1(n7228), .A2(n7259), .A3(n6440), .ZN(n6441) );
  AOI21_X1 U8090 ( .B1(n6463), .B2(n6442), .A(n6441), .ZN(P2_U3377) );
  INV_X1 U8091 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n6445) );
  INV_X1 U8092 ( .A(n6443), .ZN(n6444) );
  AOI22_X1 U8093 ( .A1(n6463), .A2(n6445), .B1(n6548), .B2(n6444), .ZN(
        P2_U3376) );
  INV_X1 U8094 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6446) );
  OAI222_X1 U8095 ( .A1(n7118), .A2(n6446), .B1(n6834), .B2(n6459), .C1(
        P2_U3151), .C2(n4532), .ZN(P2_U3288) );
  INV_X1 U8096 ( .A(n7858), .ZN(n9189) );
  INV_X1 U8097 ( .A(n9189), .ZN(n9195) );
  OAI222_X1 U8098 ( .A1(n9195), .A2(n6448), .B1(n9193), .B2(n6455), .C1(
        P1_U3086), .C2(n6447), .ZN(P1_U3351) );
  OAI222_X1 U8099 ( .A1(n9195), .A2(n6449), .B1(n9193), .B2(n6457), .C1(
        P1_U3086), .C2(n8776), .ZN(P1_U3352) );
  OAI222_X1 U8100 ( .A1(n9195), .A2(n6451), .B1(n9193), .B2(n6450), .C1(
        P1_U3086), .C2(n9332), .ZN(P1_U3350) );
  OAI222_X1 U8101 ( .A1(n9195), .A2(n6453), .B1(n9193), .B2(n6452), .C1(
        P1_U3086), .C2(n9346), .ZN(P1_U3349) );
  CLKBUF_X1 U8102 ( .A(n6834), .Z(n8328) );
  OAI222_X1 U8103 ( .A1(n7118), .A2(n4922), .B1(n8328), .B2(n6454), .C1(n9917), 
        .C2(n6523), .ZN(P2_U3294) );
  INV_X1 U8104 ( .A(n6742), .ZN(n6755) );
  OAI222_X1 U8105 ( .A1(n6755), .A2(P2_U3151), .B1(n8328), .B2(n6455), .C1(
        n7118), .C2(n4746), .ZN(P2_U3291) );
  INV_X1 U8106 ( .A(n6535), .ZN(n6562) );
  OAI222_X1 U8107 ( .A1(n7118), .A2(n4931), .B1(n8328), .B2(n6456), .C1(n9917), 
        .C2(n6562), .ZN(P2_U3293) );
  INV_X1 U8108 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6458) );
  OAI222_X1 U8109 ( .A1(n7118), .A2(n6458), .B1(n8328), .B2(n6457), .C1(
        P2_U3151), .C2(n6647), .ZN(P2_U3292) );
  OAI222_X1 U8110 ( .A1(P1_U3086), .A2(n9243), .B1(n9193), .B2(n6459), .C1(
        n9195), .C2(n5091), .ZN(P1_U3348) );
  INV_X1 U8111 ( .A(n7023), .ZN(n7137) );
  OAI222_X1 U8112 ( .A1(n7118), .A2(n6460), .B1(n6834), .B2(n6461), .C1(n9917), 
        .C2(n7137), .ZN(P2_U3287) );
  OAI222_X1 U8113 ( .A1(n7858), .A2(n6462), .B1(n9193), .B2(n6461), .C1(
        P1_U3086), .C2(n9258), .ZN(P1_U3347) );
  INV_X1 U8114 ( .A(P2_D_REG_3__SCAN_IN), .ZN(n6464) );
  NOR2_X1 U8115 ( .A1(n6493), .A2(n6464), .ZN(P2_U3262) );
  INV_X1 U8116 ( .A(P2_D_REG_5__SCAN_IN), .ZN(n6465) );
  NOR2_X1 U8117 ( .A1(n6493), .A2(n6465), .ZN(P2_U3260) );
  INV_X1 U8118 ( .A(P2_D_REG_14__SCAN_IN), .ZN(n6466) );
  NOR2_X1 U8119 ( .A1(n6493), .A2(n6466), .ZN(P2_U3251) );
  INV_X1 U8120 ( .A(P2_D_REG_12__SCAN_IN), .ZN(n6467) );
  NOR2_X1 U8121 ( .A1(n6493), .A2(n6467), .ZN(P2_U3253) );
  INV_X1 U8122 ( .A(P2_D_REG_7__SCAN_IN), .ZN(n6468) );
  NOR2_X1 U8123 ( .A1(n6493), .A2(n6468), .ZN(P2_U3258) );
  INV_X1 U8124 ( .A(P2_D_REG_6__SCAN_IN), .ZN(n6469) );
  NOR2_X1 U8125 ( .A1(n6493), .A2(n6469), .ZN(P2_U3259) );
  INV_X1 U8126 ( .A(P2_D_REG_15__SCAN_IN), .ZN(n6470) );
  NOR2_X1 U8127 ( .A1(n6493), .A2(n6470), .ZN(P2_U3250) );
  INV_X1 U8128 ( .A(P2_D_REG_4__SCAN_IN), .ZN(n6471) );
  NOR2_X1 U8129 ( .A1(n6493), .A2(n6471), .ZN(P2_U3261) );
  INV_X1 U8130 ( .A(P2_D_REG_19__SCAN_IN), .ZN(n6472) );
  NOR2_X1 U8131 ( .A1(n6493), .A2(n6472), .ZN(P2_U3246) );
  INV_X1 U8132 ( .A(P2_D_REG_18__SCAN_IN), .ZN(n6473) );
  NOR2_X1 U8133 ( .A1(n6493), .A2(n6473), .ZN(P2_U3247) );
  INV_X1 U8134 ( .A(P2_D_REG_17__SCAN_IN), .ZN(n6474) );
  NOR2_X1 U8135 ( .A1(n6493), .A2(n6474), .ZN(P2_U3248) );
  INV_X1 U8136 ( .A(P2_D_REG_16__SCAN_IN), .ZN(n6475) );
  NOR2_X1 U8137 ( .A1(n6493), .A2(n6475), .ZN(P2_U3249) );
  INV_X1 U8138 ( .A(P2_D_REG_13__SCAN_IN), .ZN(n6476) );
  NOR2_X1 U8139 ( .A1(n6493), .A2(n6476), .ZN(P2_U3252) );
  INV_X1 U8140 ( .A(n6477), .ZN(n6479) );
  INV_X1 U8141 ( .A(n7289), .ZN(n7295) );
  OAI222_X1 U8142 ( .A1(n8328), .A2(n6479), .B1(n7295), .B2(P2_U3151), .C1(
        n6478), .C2(n7118), .ZN(P2_U3286) );
  INV_X1 U8143 ( .A(n8829), .ZN(n9273) );
  OAI222_X1 U8144 ( .A1(n7858), .A2(n6480), .B1(n9193), .B2(n6479), .C1(n9273), 
        .C2(P1_U3086), .ZN(P1_U3346) );
  INV_X1 U8145 ( .A(n6481), .ZN(n6483) );
  INV_X1 U8146 ( .A(n7320), .ZN(n7323) );
  INV_X1 U8147 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6482) );
  OAI222_X1 U8148 ( .A1(n6834), .A2(n6483), .B1(n7323), .B2(n9917), .C1(n6482), 
        .C2(n7118), .ZN(P2_U3285) );
  INV_X1 U8149 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n6484) );
  INV_X1 U8150 ( .A(n8830), .ZN(n9228) );
  OAI222_X1 U8151 ( .A1(n9195), .A2(n6484), .B1(n9193), .B2(n6483), .C1(n9228), 
        .C2(P1_U3086), .ZN(P1_U3345) );
  NAND2_X1 U8152 ( .A1(n8622), .A2(n6486), .ZN(n6485) );
  AND2_X1 U8153 ( .A1(n5052), .A2(n6485), .ZN(n6693) );
  INV_X1 U8154 ( .A(n6693), .ZN(n6487) );
  OR2_X1 U8155 ( .A1(n6486), .A2(P1_U3086), .ZN(n8732) );
  NAND2_X1 U8156 ( .A1(n8660), .A2(n8732), .ZN(n6692) );
  AND2_X1 U8157 ( .A1(n6487), .A2(n6692), .ZN(n9431) );
  NOR2_X1 U8158 ( .A1(n9431), .A2(P1_U3973), .ZN(P1_U3085) );
  INV_X1 U8159 ( .A(n6488), .ZN(n6491) );
  AOI22_X1 U8160 ( .A1(n9351), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n9189), .ZN(n6489) );
  OAI21_X1 U8161 ( .B1(n6491), .B2(n9193), .A(n6489), .ZN(P1_U3344) );
  NAND2_X1 U8162 ( .A1(n6783), .A2(P2_U3893), .ZN(n6490) );
  OAI21_X1 U8163 ( .B1(P2_U3893), .B2(n5091), .A(n6490), .ZN(P2_U3498) );
  INV_X1 U8164 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6492) );
  INV_X1 U8165 ( .A(n7418), .ZN(n7427) );
  OAI222_X1 U8166 ( .A1(n7118), .A2(n6492), .B1(n6834), .B2(n6491), .C1(
        P2_U3151), .C2(n7427), .ZN(P2_U3284) );
  INV_X1 U8167 ( .A(P2_D_REG_23__SCAN_IN), .ZN(n6494) );
  NOR2_X1 U8168 ( .A1(n6493), .A2(n6494), .ZN(P2_U3242) );
  INV_X1 U8169 ( .A(P2_D_REG_10__SCAN_IN), .ZN(n6495) );
  NOR2_X1 U8170 ( .A1(n6493), .A2(n6495), .ZN(P2_U3255) );
  INV_X1 U8171 ( .A(P2_D_REG_2__SCAN_IN), .ZN(n6496) );
  NOR2_X1 U8172 ( .A1(n6493), .A2(n6496), .ZN(P2_U3263) );
  INV_X1 U8173 ( .A(P2_D_REG_21__SCAN_IN), .ZN(n6497) );
  NOR2_X1 U8174 ( .A1(n6493), .A2(n6497), .ZN(P2_U3244) );
  INV_X1 U8175 ( .A(P2_D_REG_26__SCAN_IN), .ZN(n6498) );
  NOR2_X1 U8176 ( .A1(n6493), .A2(n6498), .ZN(P2_U3239) );
  INV_X1 U8177 ( .A(P2_D_REG_25__SCAN_IN), .ZN(n6499) );
  NOR2_X1 U8178 ( .A1(n6493), .A2(n6499), .ZN(P2_U3240) );
  INV_X1 U8179 ( .A(P2_D_REG_31__SCAN_IN), .ZN(n6500) );
  NOR2_X1 U8180 ( .A1(n6493), .A2(n6500), .ZN(P2_U3234) );
  INV_X1 U8181 ( .A(P2_D_REG_24__SCAN_IN), .ZN(n6501) );
  NOR2_X1 U8182 ( .A1(n6493), .A2(n6501), .ZN(P2_U3241) );
  INV_X1 U8183 ( .A(P2_D_REG_20__SCAN_IN), .ZN(n6502) );
  NOR2_X1 U8184 ( .A1(n6493), .A2(n6502), .ZN(P2_U3245) );
  INV_X1 U8185 ( .A(P2_D_REG_8__SCAN_IN), .ZN(n6503) );
  NOR2_X1 U8186 ( .A1(n6493), .A2(n6503), .ZN(P2_U3257) );
  INV_X1 U8187 ( .A(P2_D_REG_9__SCAN_IN), .ZN(n6504) );
  NOR2_X1 U8188 ( .A1(n6493), .A2(n6504), .ZN(P2_U3256) );
  INV_X1 U8189 ( .A(P2_D_REG_29__SCAN_IN), .ZN(n6505) );
  NOR2_X1 U8190 ( .A1(n6493), .A2(n6505), .ZN(P2_U3236) );
  INV_X1 U8191 ( .A(P2_D_REG_11__SCAN_IN), .ZN(n6506) );
  NOR2_X1 U8192 ( .A1(n6493), .A2(n6506), .ZN(P2_U3254) );
  INV_X1 U8193 ( .A(P2_D_REG_28__SCAN_IN), .ZN(n6507) );
  NOR2_X1 U8194 ( .A1(n6493), .A2(n6507), .ZN(P2_U3237) );
  INV_X1 U8195 ( .A(P2_D_REG_27__SCAN_IN), .ZN(n6508) );
  NOR2_X1 U8196 ( .A1(n6493), .A2(n6508), .ZN(P2_U3238) );
  INV_X1 U8197 ( .A(P2_D_REG_30__SCAN_IN), .ZN(n6509) );
  NOR2_X1 U8198 ( .A1(n6493), .A2(n6509), .ZN(P2_U3235) );
  INV_X1 U8199 ( .A(P2_D_REG_22__SCAN_IN), .ZN(n6510) );
  NOR2_X1 U8200 ( .A1(n6493), .A2(n6510), .ZN(P2_U3243) );
  INV_X1 U8201 ( .A(n6511), .ZN(n6513) );
  INV_X1 U8202 ( .A(n7425), .ZN(n8008) );
  INV_X1 U8203 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6512) );
  OAI222_X1 U8204 ( .A1(n6834), .A2(n6513), .B1(n8008), .B2(P2_U3151), .C1(
        n6512), .C2(n7118), .ZN(P2_U3283) );
  INV_X1 U8205 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n6514) );
  INV_X1 U8206 ( .A(n8832), .ZN(n9377) );
  OAI222_X1 U8207 ( .A1(n7858), .A2(n6514), .B1(n9193), .B2(n6513), .C1(n9377), 
        .C2(P1_U3086), .ZN(P1_U3343) );
  INV_X1 U8208 ( .A(n9720), .ZN(n9200) );
  INV_X1 U8209 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n6606) );
  NOR2_X1 U8210 ( .A1(n6606), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6520) );
  AOI21_X1 U8211 ( .B1(n6516), .B2(n4709), .A(n6515), .ZN(n6517) );
  AOI21_X1 U8212 ( .B1(n6518), .B2(n4472), .A(n6517), .ZN(n6519) );
  AOI211_X1 U8213 ( .C1(P2_ADDR_REG_0__SCAN_IN), .C2(n9200), .A(n6520), .B(
        n6519), .ZN(n6521) );
  OAI21_X1 U8214 ( .B1(n4709), .B2(n9721), .A(n6521), .ZN(P2_U3182) );
  AOI211_X1 U8215 ( .C1(n6526), .C2(n6525), .A(n4472), .B(n6555), .ZN(n6544)
         );
  INV_X1 U8216 ( .A(n8066), .ZN(n9730) );
  INV_X1 U8217 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n6527) );
  NAND2_X1 U8218 ( .A1(n6528), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n6531) );
  INV_X1 U8219 ( .A(n6529), .ZN(n6530) );
  NAND2_X1 U8220 ( .A1(n6531), .A2(n6530), .ZN(n6532) );
  OAI21_X1 U8221 ( .B1(n6533), .B2(n6532), .A(n6559), .ZN(n6534) );
  AOI22_X1 U8222 ( .A1(n9200), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(n9730), .B2(
        n6534), .ZN(n6542) );
  INV_X1 U8223 ( .A(n9736), .ZN(n6749) );
  XNOR2_X1 U8224 ( .A(n6535), .B(P2_REG2_REG_2__SCAN_IN), .ZN(n6539) );
  NAND2_X1 U8225 ( .A1(n6537), .A2(n6536), .ZN(n6538) );
  NAND2_X1 U8226 ( .A1(n6539), .A2(n6538), .ZN(n6564) );
  OAI21_X1 U8227 ( .B1(n6539), .B2(n6538), .A(n6564), .ZN(n6540) );
  AOI22_X1 U8228 ( .A1(n6749), .A2(n6540), .B1(P2_REG3_REG_2__SCAN_IN), .B2(
        P2_U3151), .ZN(n6541) );
  OAI211_X1 U8229 ( .C1(n6562), .C2(n9721), .A(n6542), .B(n6541), .ZN(n6543)
         );
  OR2_X1 U8230 ( .A1(n6544), .A2(n6543), .ZN(P2_U3184) );
  INV_X1 U8231 ( .A(n6545), .ZN(n8006) );
  AND2_X1 U8232 ( .A1(n7612), .A2(n7611), .ZN(n7774) );
  INV_X1 U8233 ( .A(n7774), .ZN(n6609) );
  INV_X1 U8234 ( .A(n6546), .ZN(n6549) );
  NAND3_X1 U8235 ( .A1(n6549), .A2(n6548), .A3(n6547), .ZN(n6588) );
  AOI22_X1 U8236 ( .A1(n6609), .A2(n7954), .B1(n6588), .B2(
        P2_REG3_REG_0__SCAN_IN), .ZN(n6551) );
  AOI22_X1 U8237 ( .A1(n7973), .A2(n6598), .B1(n7968), .B2(n5373), .ZN(n6550)
         );
  NAND2_X1 U8238 ( .A1(n6551), .A2(n6550), .ZN(P2_U3172) );
  NAND2_X1 U8239 ( .A1(n6969), .A2(P1_U3973), .ZN(n6552) );
  OAI21_X1 U8240 ( .B1(P1_U3973), .B2(n4746), .A(n6552), .ZN(P1_U3558) );
  NAND2_X1 U8241 ( .A1(n8755), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n6553) );
  OAI21_X1 U8242 ( .B1(n8619), .B2(n8755), .A(n6553), .ZN(P1_U3585) );
  NAND2_X1 U8243 ( .A1(n8755), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n6554) );
  OAI21_X1 U8244 ( .B1(n9026), .B2(n8755), .A(n6554), .ZN(P1_U3574) );
  MUX2_X1 U8245 ( .A(P2_REG2_REG_3__SCAN_IN), .B(P2_REG1_REG_3__SCAN_IN), .S(
        n8046), .Z(n6636) );
  XNOR2_X1 U8246 ( .A(n6560), .B(n6636), .ZN(n6556) );
  NAND2_X1 U8247 ( .A1(n6557), .A2(n6556), .ZN(n6635) );
  OAI21_X1 U8248 ( .B1(n6557), .B2(n6556), .A(n6635), .ZN(n6572) );
  NOR2_X1 U8249 ( .A1(n9721), .A2(n6647), .ZN(n6571) );
  NAND2_X1 U8250 ( .A1(n6562), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6558) );
  INV_X1 U8251 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n6561) );
  XNOR2_X1 U8252 ( .A(n6646), .B(n6561), .ZN(n6569) );
  NAND2_X1 U8253 ( .A1(n6562), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6563) );
  NAND2_X1 U8254 ( .A1(n6564), .A2(n6563), .ZN(n6565) );
  NAND2_X1 U8255 ( .A1(n6565), .A2(n6647), .ZN(n6642) );
  OAI21_X1 U8256 ( .B1(n6566), .B2(P2_REG2_REG_3__SCAN_IN), .A(n6644), .ZN(
        n6567) );
  AOI22_X1 U8257 ( .A1(n9200), .A2(P2_ADDR_REG_3__SCAN_IN), .B1(n6749), .B2(
        n6567), .ZN(n6568) );
  NAND2_X1 U8258 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_U3151), .ZN(n6622) );
  OAI211_X1 U8259 ( .C1(n6569), .C2(n8066), .A(n6568), .B(n6622), .ZN(n6570)
         );
  AOI211_X1 U8260 ( .C1(n6572), .C2(n9729), .A(n6571), .B(n6570), .ZN(n6573)
         );
  INV_X1 U8261 ( .A(n6573), .ZN(P2_U3185) );
  XOR2_X1 U8262 ( .A(n6575), .B(n6574), .Z(n6579) );
  AOI22_X1 U8263 ( .A1(n8006), .A2(n7982), .B1(n7968), .B2(n9745), .ZN(n6576)
         );
  OAI21_X1 U8264 ( .B1(n7991), .B2(n9779), .A(n6576), .ZN(n6577) );
  AOI21_X1 U8265 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(n6588), .A(n6577), .ZN(
        n6578) );
  OAI21_X1 U8266 ( .B1(n7977), .B2(n6579), .A(n6578), .ZN(P2_U3162) );
  INV_X1 U8267 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n6581) );
  INV_X1 U8268 ( .A(n6580), .ZN(n6582) );
  INV_X1 U8269 ( .A(n8833), .ZN(n9392) );
  OAI222_X1 U8270 ( .A1(n7858), .A2(n6581), .B1(n9193), .B2(n6582), .C1(
        P1_U3086), .C2(n9392), .ZN(P1_U3342) );
  INV_X1 U8271 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6583) );
  INV_X1 U8272 ( .A(n8050), .ZN(n9647) );
  OAI222_X1 U8273 ( .A1(n7118), .A2(n6583), .B1(n6834), .B2(n6582), .C1(n9917), 
        .C2(n9647), .ZN(P2_U3282) );
  XOR2_X1 U8274 ( .A(n6585), .B(n6584), .Z(n6590) );
  AOI22_X1 U8275 ( .A1(n7982), .A2(n5373), .B1(n8004), .B2(n7968), .ZN(n6586)
         );
  OAI21_X1 U8276 ( .B1(n7991), .B2(n9769), .A(n6586), .ZN(n6587) );
  AOI21_X1 U8277 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(n6588), .A(n6587), .ZN(
        n6589) );
  OAI21_X1 U8278 ( .B1(n6590), .B2(n7977), .A(n6589), .ZN(P2_U3177) );
  INV_X1 U8279 ( .A(n6591), .ZN(n6617) );
  AOI22_X1 U8280 ( .A1(n9397), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n9189), .ZN(n6592) );
  OAI21_X1 U8281 ( .B1(n6617), .B2(n9193), .A(n6592), .ZN(P1_U3341) );
  INV_X1 U8282 ( .A(n9796), .ZN(n9831) );
  OAI21_X1 U8283 ( .B1(n9831), .B2(n9765), .A(n6609), .ZN(n6593) );
  OR2_X1 U8284 ( .A1(n9763), .A2(n9760), .ZN(n6605) );
  NAND2_X1 U8285 ( .A1(n6593), .A2(n6605), .ZN(n6597) );
  INV_X1 U8286 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n6594) );
  NOR2_X1 U8287 ( .A1(n9836), .A2(n6594), .ZN(n6595) );
  AOI21_X1 U8288 ( .B1(n9836), .B2(n6597), .A(n6595), .ZN(n6596) );
  OAI21_X1 U8289 ( .B1(n6614), .B2(n8254), .A(n6596), .ZN(P2_U3390) );
  INV_X1 U8290 ( .A(n6597), .ZN(n6600) );
  AOI22_X1 U8291 ( .A1(n8245), .A2(n6598), .B1(n9852), .B2(
        P2_REG1_REG_0__SCAN_IN), .ZN(n6599) );
  OAI21_X1 U8292 ( .B1(n6600), .B2(n9852), .A(n6599), .ZN(P2_U3459) );
  MUX2_X1 U8293 ( .A(n5772), .B(n6602), .S(n6601), .Z(n6603) );
  NAND2_X1 U8294 ( .A1(n6604), .A2(n6603), .ZN(n6610) );
  NOR2_X2 U8295 ( .A1(n6610), .A2(n8120), .ZN(n9751) );
  INV_X1 U8296 ( .A(n9751), .ZN(n8076) );
  INV_X1 U8297 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n6612) );
  OAI21_X1 U8298 ( .B1(n7377), .B2(n6606), .A(n6605), .ZN(n6607) );
  AOI21_X1 U8299 ( .B1(n6609), .B2(n6608), .A(n6607), .ZN(n6611) );
  NAND2_X2 U8300 ( .A1(n6610), .A2(n7377), .ZN(n9775) );
  MUX2_X1 U8301 ( .A(n6612), .B(n6611), .S(n9775), .Z(n6613) );
  OAI21_X1 U8302 ( .B1(n8076), .B2(n6614), .A(n6613), .ZN(P2_U3233) );
  INV_X1 U8303 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6616) );
  NAND2_X1 U8304 ( .A1(n8519), .A2(P1_U3973), .ZN(n6615) );
  OAI21_X1 U8305 ( .B1(n6616), .B2(P1_U3973), .A(n6615), .ZN(P1_U3568) );
  INV_X1 U8306 ( .A(n8044), .ZN(n9665) );
  OAI222_X1 U8307 ( .A1(n9665), .A2(n9917), .B1(n8328), .B2(n6617), .C1(n7118), 
        .C2(n6616), .ZN(P2_U3281) );
  INV_X1 U8308 ( .A(n7987), .ZN(n6626) );
  OAI211_X1 U8309 ( .C1(n6620), .C2(n6619), .A(n6618), .B(n7954), .ZN(n6625)
         );
  NAND2_X1 U8310 ( .A1(n7982), .A2(n9745), .ZN(n6621) );
  OAI211_X1 U8311 ( .C1(n6872), .C2(n7984), .A(n6622), .B(n6621), .ZN(n6623)
         );
  AOI21_X1 U8312 ( .B1(n7973), .B2(n9789), .A(n6623), .ZN(n6624) );
  OAI211_X1 U8313 ( .C1(n6626), .C2(P2_REG3_REG_3__SCAN_IN), .A(n6625), .B(
        n6624), .ZN(P2_U3158) );
  XNOR2_X1 U8314 ( .A(n6628), .B(n6627), .ZN(n6687) );
  NAND2_X1 U8315 ( .A1(n6630), .A2(n6629), .ZN(n6730) );
  AOI22_X1 U8316 ( .A1(n8430), .A2(n9519), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        n6730), .ZN(n6632) );
  INV_X1 U8317 ( .A(n8427), .ZN(n8454) );
  NAND2_X1 U8318 ( .A1(n8454), .A2(n6898), .ZN(n6631) );
  OAI211_X1 U8319 ( .C1(n6687), .C2(n8462), .A(n6632), .B(n6631), .ZN(P1_U3232) );
  INV_X1 U8320 ( .A(n6633), .ZN(n6672) );
  INV_X1 U8321 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n6634) );
  OAI222_X1 U8322 ( .A1(n6834), .A2(n6672), .B1(n4759), .B2(n9917), .C1(n6634), 
        .C2(n7118), .ZN(P2_U3280) );
  MUX2_X1 U8323 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n8046), .Z(n6756) );
  XOR2_X1 U8324 ( .A(n6742), .B(n6756), .Z(n6638) );
  OAI21_X1 U8325 ( .B1(n6636), .B2(n6647), .A(n6635), .ZN(n6637) );
  NOR2_X1 U8326 ( .A1(n6637), .A2(n6638), .ZN(n6754) );
  AOI211_X1 U8327 ( .C1(n6638), .C2(n6637), .A(n4472), .B(n6754), .ZN(n6639)
         );
  INV_X1 U8328 ( .A(n6639), .ZN(n6660) );
  NAND2_X1 U8329 ( .A1(n6644), .A2(n6642), .ZN(n6640) );
  XNOR2_X1 U8330 ( .A(n6742), .B(P2_REG2_REG_4__SCAN_IN), .ZN(n6641) );
  NAND2_X1 U8331 ( .A1(n6640), .A2(n6641), .ZN(n6744) );
  INV_X1 U8332 ( .A(n6641), .ZN(n6643) );
  NAND3_X1 U8333 ( .A1(n6644), .A2(n6643), .A3(n6642), .ZN(n6645) );
  AOI21_X1 U8334 ( .B1(n6744), .B2(n6645), .A(n9736), .ZN(n6658) );
  INV_X1 U8335 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n6656) );
  NAND2_X1 U8336 ( .A1(n6646), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6650) );
  NAND2_X1 U8337 ( .A1(n6648), .A2(n6647), .ZN(n6649) );
  NAND2_X1 U8338 ( .A1(n6650), .A2(n6649), .ZN(n6653) );
  INV_X1 U8339 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6651) );
  MUX2_X1 U8340 ( .A(n6651), .B(P2_REG1_REG_4__SCAN_IN), .S(n6742), .Z(n6652)
         );
  NOR2_X1 U8341 ( .A1(n6653), .A2(n6652), .ZN(n6654) );
  NOR2_X1 U8342 ( .A1(n6741), .A2(n6654), .ZN(n6655) );
  OAI22_X1 U8343 ( .A1(n9720), .A2(n6656), .B1(n8066), .B2(n6655), .ZN(n6657)
         );
  INV_X1 U8344 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n9929) );
  NOR2_X1 U8345 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9929), .ZN(n6680) );
  NOR3_X1 U8346 ( .A1(n6658), .A2(n6657), .A3(n6680), .ZN(n6659) );
  OAI211_X1 U8347 ( .C1(n9721), .C2(n6755), .A(n6660), .B(n6659), .ZN(P2_U3186) );
  INV_X1 U8348 ( .A(n6662), .ZN(n6663) );
  AOI21_X1 U8349 ( .B1(n7612), .B2(n6661), .A(n6663), .ZN(n9780) );
  NAND2_X1 U8350 ( .A1(n8020), .A2(n6664), .ZN(n9773) );
  NAND2_X1 U8351 ( .A1(n9768), .A2(n9773), .ZN(n6665) );
  OAI21_X1 U8352 ( .B1(n6667), .B2(n6661), .A(n6666), .ZN(n6668) );
  AOI222_X1 U8353 ( .A1(n9765), .A2(n6668), .B1(n9745), .B2(n9746), .C1(n8006), 
        .C2(n9744), .ZN(n9778) );
  MUX2_X1 U8354 ( .A(n6425), .B(n9778), .S(n9775), .Z(n6671) );
  AOI22_X1 U8355 ( .A1(n9751), .A2(n6669), .B1(n9770), .B2(
        P2_REG3_REG_1__SCAN_IN), .ZN(n6670) );
  OAI211_X1 U8356 ( .C1(n9780), .C2(n8208), .A(n6671), .B(n6670), .ZN(P2_U3232) );
  INV_X1 U8357 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n6673) );
  OAI222_X1 U8358 ( .A1(n9195), .A2(n6673), .B1(n9193), .B2(n6672), .C1(n8836), 
        .C2(P1_U3086), .ZN(P1_U3340) );
  NAND2_X1 U8359 ( .A1(n8755), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n6674) );
  OAI21_X1 U8360 ( .B1(n8898), .B2(n8755), .A(n6674), .ZN(P1_U3583) );
  INV_X1 U8361 ( .A(n6675), .ZN(n6676) );
  AOI21_X1 U8362 ( .B1(n6678), .B2(n6677), .A(n6676), .ZN(n6684) );
  NOR2_X1 U8363 ( .A1(n9761), .A2(n7971), .ZN(n6679) );
  AOI211_X1 U8364 ( .C1(n7968), .C2(n8003), .A(n6680), .B(n6679), .ZN(n6681)
         );
  OAI21_X1 U8365 ( .B1(n9795), .B2(n7991), .A(n6681), .ZN(n6682) );
  AOI21_X1 U8366 ( .B1(n6794), .B2(n7987), .A(n6682), .ZN(n6683) );
  OAI21_X1 U8367 ( .B1(n6684), .B2(n7977), .A(n6683), .ZN(P2_U3170) );
  INV_X1 U8368 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n6685) );
  AOI21_X1 U8369 ( .B1(n9302), .B2(n6685), .A(n5286), .ZN(n9301) );
  NOR2_X1 U8370 ( .A1(n6686), .A2(n6685), .ZN(n8758) );
  MUX2_X1 U8371 ( .A(n8758), .B(n6687), .S(n5287), .Z(n6688) );
  NAND2_X1 U8372 ( .A1(n6688), .A2(n8657), .ZN(n6689) );
  OAI211_X1 U8373 ( .C1(P1_IR_REG_0__SCAN_IN), .C2(n9301), .A(n6689), .B(
        P1_U3973), .ZN(n9319) );
  INV_X1 U8374 ( .A(n9319), .ZN(n6705) );
  INV_X1 U8375 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n9511) );
  MUX2_X1 U8376 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n9511), .S(n8777), .Z(n6696)
         );
  INV_X1 U8377 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n6690) );
  NAND2_X1 U8378 ( .A1(n8763), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6691) );
  NAND2_X1 U8379 ( .A1(n8757), .A2(n6691), .ZN(n6695) );
  NAND2_X1 U8380 ( .A1(n6693), .A2(n6692), .ZN(n9305) );
  OR2_X1 U8381 ( .A1(n5286), .A2(n5287), .ZN(n6694) );
  NAND2_X1 U8382 ( .A1(n6696), .A2(n6695), .ZN(n8773) );
  OAI211_X1 U8383 ( .C1(n6696), .C2(n6695), .A(n9446), .B(n8773), .ZN(n6703)
         );
  AOI22_X1 U8384 ( .A1(n9431), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n6702) );
  INV_X1 U8385 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n9624) );
  MUX2_X1 U8386 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n9624), .S(n8777), .Z(n6699)
         );
  INV_X1 U8387 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n9622) );
  MUX2_X1 U8388 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n9622), .S(n8763), .Z(n8762)
         );
  AND2_X1 U8389 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n8761) );
  NAND2_X1 U8390 ( .A1(n8762), .A2(n8761), .ZN(n8760) );
  NAND2_X1 U8391 ( .A1(n8763), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6697) );
  NAND2_X1 U8392 ( .A1(n8760), .A2(n6697), .ZN(n6698) );
  OR2_X1 U8393 ( .A1(n9305), .A2(n9302), .ZN(n9413) );
  NAND2_X1 U8394 ( .A1(n6699), .A2(n6698), .ZN(n8779) );
  OAI211_X1 U8395 ( .C1(n6699), .C2(n6698), .A(n9454), .B(n8779), .ZN(n6701)
         );
  INV_X1 U8396 ( .A(n9460), .ZN(n9443) );
  NAND2_X1 U8397 ( .A1(n9443), .A2(n8777), .ZN(n6700) );
  NAND4_X1 U8398 ( .A1(n6703), .A2(n6702), .A3(n6701), .A4(n6700), .ZN(n6704)
         );
  OR2_X1 U8399 ( .A1(n6705), .A2(n6704), .ZN(P1_U3245) );
  INV_X1 U8400 ( .A(n6706), .ZN(n6719) );
  INV_X1 U8401 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n6707) );
  OAI222_X1 U8402 ( .A1(n6834), .A2(n6719), .B1(n8030), .B2(P2_U3151), .C1(
        n6707), .C2(n7118), .ZN(P2_U3278) );
  INV_X1 U8403 ( .A(n6708), .ZN(n6709) );
  NOR2_X1 U8404 ( .A1(n6710), .A2(n6709), .ZN(n6714) );
  INV_X1 U8405 ( .A(n6712), .ZN(n6713) );
  AOI21_X1 U8406 ( .B1(n6714), .B2(n6711), .A(n6713), .ZN(n6717) );
  AOI22_X1 U8407 ( .A1(n8430), .A2(n9527), .B1(P1_REG3_REG_2__SCAN_IN), .B2(
        n6730), .ZN(n6716) );
  INV_X1 U8408 ( .A(n6896), .ZN(n9491) );
  AOI22_X1 U8409 ( .A1(n8455), .A2(n6898), .B1(n8454), .B2(n9491), .ZN(n6715)
         );
  OAI211_X1 U8410 ( .C1(n6717), .C2(n8462), .A(n6716), .B(n6715), .ZN(P1_U3237) );
  INV_X1 U8411 ( .A(n9444), .ZN(n8809) );
  INV_X1 U8412 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n6718) );
  OAI222_X1 U8413 ( .A1(P1_U3086), .A2(n8809), .B1(n9193), .B2(n6719), .C1(
        n6718), .C2(n7858), .ZN(P1_U3338) );
  INV_X1 U8414 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n6721) );
  INV_X1 U8415 ( .A(n6720), .ZN(n6722) );
  INV_X1 U8416 ( .A(n8040), .ZN(n9701) );
  OAI222_X1 U8417 ( .A1(n7118), .A2(n6721), .B1(n8328), .B2(n6722), .C1(
        P2_U3151), .C2(n9701), .ZN(P2_U3279) );
  INV_X1 U8418 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n6723) );
  INV_X1 U8419 ( .A(n9435), .ZN(n8838) );
  OAI222_X1 U8420 ( .A1(n9195), .A2(n6723), .B1(n9193), .B2(n6722), .C1(
        P1_U3086), .C2(n8838), .ZN(P1_U3339) );
  INV_X1 U8421 ( .A(n6711), .ZN(n6725) );
  AOI21_X1 U8422 ( .B1(n6726), .B2(n6724), .A(n6725), .ZN(n6732) );
  INV_X1 U8423 ( .A(n8430), .ZN(n8407) );
  INV_X1 U8424 ( .A(n8756), .ZN(n6727) );
  INV_X1 U8425 ( .A(n8754), .ZN(n6901) );
  OAI22_X1 U8426 ( .A1(n6727), .A2(n8426), .B1(n8427), .B2(n6901), .ZN(n6728)
         );
  AOI211_X1 U8427 ( .C1(P1_REG3_REG_1__SCAN_IN), .C2(n6730), .A(n6729), .B(
        n6728), .ZN(n6731) );
  OAI21_X1 U8428 ( .B1(n6732), .B2(n8462), .A(n6731), .ZN(P1_U3222) );
  XOR2_X1 U8429 ( .A(n6733), .B(n6734), .Z(n6739) );
  NOR2_X1 U8430 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10058), .ZN(n6747) );
  NOR2_X1 U8431 ( .A1(n7091), .A2(n7984), .ZN(n6735) );
  AOI211_X1 U8432 ( .C1(n7982), .C2(n9747), .A(n6747), .B(n6735), .ZN(n6736)
         );
  OAI21_X1 U8433 ( .B1(n9801), .B2(n7991), .A(n6736), .ZN(n6737) );
  AOI21_X1 U8434 ( .B1(n6876), .B2(n7987), .A(n6737), .ZN(n6738) );
  OAI21_X1 U8435 ( .B1(n6739), .B2(n7977), .A(n6738), .ZN(P2_U3167) );
  INV_X1 U8436 ( .A(n9204), .ZN(n9206) );
  INV_X1 U8437 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n6740) );
  OAI222_X1 U8438 ( .A1(n8328), .A2(n6764), .B1(n9206), .B2(n9917), .C1(n6740), 
        .C2(n7118), .ZN(P2_U3277) );
  XNOR2_X1 U8439 ( .A(n6801), .B(P2_REG1_REG_5__SCAN_IN), .ZN(n6761) );
  INV_X1 U8440 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n6752) );
  INV_X1 U8441 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n6793) );
  OR2_X1 U8442 ( .A1(n6742), .A2(n6793), .ZN(n6743) );
  NAND2_X1 U8443 ( .A1(n6744), .A2(n6743), .ZN(n6746) );
  NOR2_X1 U8444 ( .A1(n6746), .A2(n6805), .ZN(n6745) );
  OAI21_X1 U8445 ( .B1(n4448), .B2(P2_REG2_REG_5__SCAN_IN), .A(n6815), .ZN(
        n6748) );
  AOI21_X1 U8446 ( .B1(n6749), .B2(n6748), .A(n6747), .ZN(n6751) );
  INV_X1 U8447 ( .A(n9721), .ZN(n7142) );
  NAND2_X1 U8448 ( .A1(n7142), .A2(n6753), .ZN(n6750) );
  OAI211_X1 U8449 ( .C1(n6752), .C2(n9720), .A(n6751), .B(n6750), .ZN(n6760)
         );
  MUX2_X1 U8450 ( .A(P2_REG2_REG_5__SCAN_IN), .B(P2_REG1_REG_5__SCAN_IN), .S(
        n8046), .Z(n6806) );
  XOR2_X1 U8451 ( .A(n6753), .B(n6806), .Z(n6758) );
  AOI21_X1 U8452 ( .B1(n6756), .B2(n6755), .A(n6754), .ZN(n6757) );
  NOR2_X1 U8453 ( .A1(n6757), .A2(n6758), .ZN(n6804) );
  AOI211_X1 U8454 ( .C1(n6758), .C2(n6757), .A(n4472), .B(n6804), .ZN(n6759)
         );
  AOI211_X1 U8455 ( .C1(n9730), .C2(n6761), .A(n6760), .B(n6759), .ZN(n6762)
         );
  INV_X1 U8456 ( .A(n6762), .ZN(P2_U3187) );
  INV_X1 U8457 ( .A(n8842), .ZN(n9459) );
  INV_X1 U8458 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n6763) );
  OAI222_X1 U8459 ( .A1(P1_U3086), .A2(n9459), .B1(n9193), .B2(n6764), .C1(
        n6763), .C2(n9195), .ZN(P1_U3337) );
  NAND2_X1 U8460 ( .A1(n8005), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n6765) );
  OAI21_X1 U8461 ( .B1(n7741), .B2(n8005), .A(n6765), .ZN(P2_U3521) );
  NAND2_X1 U8462 ( .A1(n8005), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n6766) );
  OAI21_X1 U8463 ( .B1(n8081), .B2(n8005), .A(n6766), .ZN(P2_U3520) );
  NAND2_X1 U8464 ( .A1(n6767), .A2(n8444), .ZN(n6777) );
  AOI21_X1 U8465 ( .B1(n6769), .B2(n6771), .A(n6770), .ZN(n6776) );
  AOI22_X1 U8466 ( .A1(n8455), .A2(n9491), .B1(n6978), .B2(n8430), .ZN(n6775)
         );
  NOR2_X1 U8467 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6772), .ZN(n9307) );
  NOR2_X1 U8468 ( .A1(n8427), .A2(n7160), .ZN(n6773) );
  AOI211_X1 U8469 ( .C1(n8446), .C2(n6977), .A(n9307), .B(n6773), .ZN(n6774)
         );
  OAI211_X1 U8470 ( .C1(n6777), .C2(n6776), .A(n6775), .B(n6774), .ZN(P1_U3230) );
  AOI21_X1 U8471 ( .B1(n6779), .B2(n6778), .A(n7977), .ZN(n6781) );
  NAND2_X1 U8472 ( .A1(n6781), .A2(n6780), .ZN(n6787) );
  NAND2_X1 U8473 ( .A1(P2_U3151), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n6810) );
  INV_X1 U8474 ( .A(n6810), .ZN(n6782) );
  AOI21_X1 U8475 ( .B1(n6783), .B2(n7968), .A(n6782), .ZN(n6784) );
  OAI21_X1 U8476 ( .B1(n5437), .B2(n7971), .A(n6784), .ZN(n6785) );
  AOI21_X1 U8477 ( .B1(n6843), .B2(n7987), .A(n6785), .ZN(n6786) );
  OAI211_X1 U8478 ( .C1(n6860), .C2(n7991), .A(n6787), .B(n6786), .ZN(P2_U3179) );
  XNOR2_X1 U8479 ( .A(n6788), .B(n6790), .ZN(n9797) );
  AND2_X1 U8480 ( .A1(n6835), .A2(n6789), .ZN(n6791) );
  XNOR2_X1 U8481 ( .A(n6791), .B(n6790), .ZN(n6792) );
  AOI222_X1 U8482 ( .A1(n9765), .A2(n6792), .B1(n8004), .B2(n9744), .C1(n8003), 
        .C2(n9746), .ZN(n9794) );
  MUX2_X1 U8483 ( .A(n6793), .B(n9794), .S(n9775), .Z(n6797) );
  AOI22_X1 U8484 ( .A1(n9751), .A2(n6795), .B1(n9770), .B2(n6794), .ZN(n6796)
         );
  OAI211_X1 U8485 ( .C1(n8208), .C2(n9797), .A(n6797), .B(n6796), .ZN(P2_U3229) );
  INV_X1 U8486 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n6798) );
  MUX2_X1 U8487 ( .A(n6798), .B(P2_REG1_REG_6__SCAN_IN), .S(n6920), .Z(n6803)
         );
  INV_X1 U8488 ( .A(n6799), .ZN(n6800) );
  NOR2_X1 U8489 ( .A1(n6802), .A2(n6803), .ZN(n6918) );
  AOI21_X1 U8490 ( .B1(n6803), .B2(n6802), .A(n6918), .ZN(n6823) );
  MUX2_X1 U8491 ( .A(P2_REG2_REG_6__SCAN_IN), .B(P2_REG1_REG_6__SCAN_IN), .S(
        n8046), .Z(n6917) );
  XOR2_X1 U8492 ( .A(n6920), .B(n6917), .Z(n6807) );
  OAI21_X1 U8493 ( .B1(n6808), .B2(n6807), .A(n6916), .ZN(n6809) );
  NAND2_X1 U8494 ( .A1(n6809), .A2(n9729), .ZN(n6822) );
  INV_X1 U8495 ( .A(n6920), .ZN(n6820) );
  INV_X1 U8496 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n6811) );
  OAI21_X1 U8497 ( .B1(n9720), .B2(n6811), .A(n6810), .ZN(n6819) );
  INV_X1 U8498 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n6812) );
  MUX2_X1 U8499 ( .A(n6812), .B(P2_REG2_REG_6__SCAN_IN), .S(n6920), .Z(n6814)
         );
  INV_X1 U8500 ( .A(n6919), .ZN(n6817) );
  NAND3_X1 U8501 ( .A1(n6815), .A2(n6814), .A3(n6813), .ZN(n6816) );
  AOI21_X1 U8502 ( .B1(n6817), .B2(n6816), .A(n9736), .ZN(n6818) );
  AOI211_X1 U8503 ( .C1(n7142), .C2(n6820), .A(n6819), .B(n6818), .ZN(n6821)
         );
  OAI211_X1 U8504 ( .C1(n6823), .C2(n8066), .A(n6822), .B(n6821), .ZN(P2_U3188) );
  OAI21_X1 U8505 ( .B1(n6825), .B2(n6824), .A(n6769), .ZN(n6830) );
  AOI22_X1 U8506 ( .A1(n8455), .A2(n8754), .B1(n9534), .B2(n8460), .ZN(n6828)
         );
  NOR2_X1 U8507 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6826), .ZN(n8768) );
  AOI21_X1 U8508 ( .B1(n8446), .B2(n6826), .A(n8768), .ZN(n6827) );
  OAI211_X1 U8509 ( .C1(n6970), .C2(n8427), .A(n6828), .B(n6827), .ZN(n6829)
         );
  AOI21_X1 U8510 ( .B1(n6830), .B2(n8444), .A(n6829), .ZN(n6831) );
  INV_X1 U8511 ( .A(n6831), .ZN(P1_U3218) );
  INV_X1 U8512 ( .A(n6832), .ZN(n6853) );
  INV_X1 U8513 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n6833) );
  OAI222_X1 U8514 ( .A1(n6834), .A2(n6853), .B1(P2_U3151), .B2(n7806), .C1(
        n6833), .C2(n7118), .ZN(P2_U3275) );
  INV_X1 U8515 ( .A(n9765), .ZN(n7505) );
  XNOR2_X1 U8516 ( .A(n5434), .B(n6863), .ZN(n7778) );
  NAND2_X1 U8517 ( .A1(n6835), .A2(n4916), .ZN(n6870) );
  NAND2_X1 U8518 ( .A1(n6870), .A2(n6836), .ZN(n6838) );
  NAND2_X1 U8519 ( .A1(n6838), .A2(n6837), .ZN(n6839) );
  XOR2_X1 U8520 ( .A(n7778), .B(n6839), .Z(n6840) );
  OAI222_X1 U8521 ( .A1(n9760), .A2(n6986), .B1(n9762), .B2(n5437), .C1(n7505), 
        .C2(n6840), .ZN(n6857) );
  INV_X1 U8522 ( .A(n6857), .ZN(n6847) );
  NAND2_X1 U8523 ( .A1(n6866), .A2(n6841), .ZN(n6842) );
  XNOR2_X1 U8524 ( .A(n6842), .B(n7778), .ZN(n6858) );
  AOI22_X1 U8525 ( .A1(n9777), .A2(P2_REG2_REG_6__SCAN_IN), .B1(n9770), .B2(
        n6843), .ZN(n6844) );
  OAI21_X1 U8526 ( .B1(n6860), .B2(n8076), .A(n6844), .ZN(n6845) );
  AOI21_X1 U8527 ( .B1(n6858), .B2(n9753), .A(n6845), .ZN(n6846) );
  OAI21_X1 U8528 ( .B1(n6847), .B2(n9777), .A(n6846), .ZN(P2_U3227) );
  INV_X1 U8529 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n6849) );
  INV_X1 U8530 ( .A(n6848), .ZN(n6850) );
  OAI222_X1 U8531 ( .A1(n7118), .A2(n6849), .B1(n8328), .B2(n6850), .C1(n8064), 
        .C2(P2_U3151), .ZN(P2_U3276) );
  INV_X1 U8532 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n6851) );
  OAI222_X1 U8533 ( .A1(n9195), .A2(n6851), .B1(n9193), .B2(n6850), .C1(
        P1_U3086), .C2(n4453), .ZN(P1_U3336) );
  OAI222_X1 U8534 ( .A1(n6854), .A2(P1_U3086), .B1(n9193), .B2(n6853), .C1(
        n6852), .C2(n9195), .ZN(P1_U3335) );
  INV_X1 U8535 ( .A(n6855), .ZN(n6914) );
  AOI22_X1 U8536 ( .A1(n7808), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_21__SCAN_IN), .B2(n8326), .ZN(n6856) );
  OAI21_X1 U8537 ( .B1(n6914), .B2(n8328), .A(n6856), .ZN(P2_U3274) );
  AOI21_X1 U8538 ( .B1(n9831), .B2(n6858), .A(n6857), .ZN(n6865) );
  INV_X1 U8539 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n6859) );
  OAI22_X1 U8540 ( .A1(n6860), .A2(n8254), .B1(n9836), .B2(n6859), .ZN(n6861)
         );
  INV_X1 U8541 ( .A(n6861), .ZN(n6862) );
  OAI21_X1 U8542 ( .B1(n6865), .B2(n9838), .A(n6862), .ZN(P2_U3408) );
  AOI22_X1 U8543 ( .A1(n8245), .A2(n6863), .B1(n9852), .B2(
        P2_REG1_REG_6__SCAN_IN), .ZN(n6864) );
  OAI21_X1 U8544 ( .B1(n6865), .B2(n9852), .A(n6864), .ZN(P2_U3465) );
  OAI21_X1 U8545 ( .B1(n6867), .B2(n7775), .A(n6866), .ZN(n9804) );
  INV_X1 U8546 ( .A(n9804), .ZN(n6882) );
  INV_X1 U8547 ( .A(n9773), .ZN(n6868) );
  NAND2_X1 U8548 ( .A1(n9775), .A2(n6868), .ZN(n7202) );
  NAND2_X1 U8549 ( .A1(n6870), .A2(n6869), .ZN(n6871) );
  XNOR2_X1 U8550 ( .A(n6871), .B(n7775), .ZN(n6875) );
  INV_X1 U8551 ( .A(n9768), .ZN(n7093) );
  OAI22_X1 U8552 ( .A1(n7091), .A2(n9760), .B1(n6872), .B2(n9762), .ZN(n6873)
         );
  AOI21_X1 U8553 ( .B1(n9804), .B2(n7093), .A(n6873), .ZN(n6874) );
  OAI21_X1 U8554 ( .B1(n7505), .B2(n6875), .A(n6874), .ZN(n9802) );
  NAND2_X1 U8555 ( .A1(n9802), .A2(n9775), .ZN(n6881) );
  INV_X1 U8556 ( .A(n6876), .ZN(n6877) );
  OAI22_X1 U8557 ( .A1(n9775), .A2(n4754), .B1(n6877), .B2(n7377), .ZN(n6878)
         );
  AOI21_X1 U8558 ( .B1(n9751), .B2(n6879), .A(n6878), .ZN(n6880) );
  OAI211_X1 U8559 ( .C1(n6882), .C2(n7202), .A(n6881), .B(n6880), .ZN(P2_U3228) );
  INV_X1 U8560 ( .A(n8660), .ZN(n6884) );
  NAND2_X2 U8561 ( .A1(n6884), .A2(n6883), .ZN(n9512) );
  OAI21_X1 U8562 ( .B1(n6885), .B2(n8660), .A(n9512), .ZN(n6888) );
  NAND4_X1 U8563 ( .A1(n6888), .A2(n6887), .A3(n9089), .A4(n6886), .ZN(n6889)
         );
  NAND2_X2 U8564 ( .A1(n6889), .A2(n9499), .ZN(n9510) );
  NOR2_X1 U8565 ( .A1(n6890), .A2(n4453), .ZN(n6891) );
  NAND2_X1 U8566 ( .A1(n9510), .A2(n6891), .ZN(n7217) );
  NAND2_X1 U8567 ( .A1(n8655), .A2(n9513), .ZN(n6933) );
  AND2_X1 U8568 ( .A1(n6893), .A2(n6892), .ZN(n6894) );
  OR2_X1 U8569 ( .A1(n6933), .A2(n6894), .ZN(n9505) );
  INV_X1 U8570 ( .A(n9505), .ZN(n9597) );
  NAND2_X1 U8571 ( .A1(n9510), .A2(n9597), .ZN(n6895) );
  NAND2_X1 U8572 ( .A1(n6896), .A2(n9534), .ZN(n8672) );
  NAND2_X1 U8573 ( .A1(n8672), .A2(n8468), .ZN(n8627) );
  NAND2_X1 U8574 ( .A1(n8756), .A2(n9519), .ZN(n7027) );
  XNOR2_X2 U8575 ( .A(n6898), .B(n6897), .ZN(n7028) );
  NAND2_X1 U8576 ( .A1(n7027), .A2(n7028), .ZN(n6900) );
  NAND2_X1 U8577 ( .A1(n6900), .A2(n6899), .ZN(n9486) );
  XNOR2_X1 U8578 ( .A(n8754), .B(n9501), .ZN(n9488) );
  NAND2_X1 U8579 ( .A1(n9486), .A2(n9488), .ZN(n6903) );
  NAND2_X1 U8580 ( .A1(n6901), .A2(n9501), .ZN(n6902) );
  NAND2_X1 U8581 ( .A1(n6903), .A2(n6902), .ZN(n6973) );
  XOR2_X1 U8582 ( .A(n8627), .B(n6973), .Z(n9537) );
  INV_X1 U8583 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n6909) );
  NAND2_X1 U8584 ( .A1(n8589), .A2(n8731), .ZN(n6904) );
  INV_X1 U8585 ( .A(n7028), .ZN(n6905) );
  NAND2_X1 U8586 ( .A1(n6905), .A2(n6932), .ZN(n7033) );
  NAND2_X1 U8587 ( .A1(n6934), .A2(n7030), .ZN(n6906) );
  NOR2_X1 U8588 ( .A1(n8754), .A2(n9501), .ZN(n8673) );
  NAND2_X1 U8589 ( .A1(n8754), .A2(n9501), .ZN(n8670) );
  XNOR2_X1 U8590 ( .A(n8627), .B(n4367), .ZN(n6908) );
  AOI222_X1 U8591 ( .A1(n9493), .A2(n6908), .B1(n8754), .B2(n9489), .C1(n6969), 
        .C2(n9490), .ZN(n9536) );
  MUX2_X1 U8592 ( .A(n6909), .B(n9536), .S(n9510), .Z(n6913) );
  AOI211_X1 U8593 ( .C1(n9534), .C2(n9497), .A(n9568), .B(n4369), .ZN(n9533)
         );
  OAI22_X1 U8594 ( .A1(n9067), .A2(n6974), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        n9499), .ZN(n6911) );
  AOI21_X1 U8595 ( .B1(n9533), .B2(n9480), .A(n6911), .ZN(n6912) );
  OAI211_X1 U8596 ( .C1(n9071), .C2(n9537), .A(n6913), .B(n6912), .ZN(P1_U3290) );
  OAI222_X1 U8597 ( .A1(n9195), .A2(n6915), .B1(n9193), .B2(n6914), .C1(
        P1_U3086), .C2(n8738), .ZN(P1_U3334) );
  MUX2_X1 U8598 ( .A(P2_REG2_REG_7__SCAN_IN), .B(P2_REG1_REG_7__SCAN_IN), .S(
        n8046), .Z(n7005) );
  XNOR2_X1 U8599 ( .A(n7005), .B(n7007), .ZN(n7008) );
  XOR2_X1 U8600 ( .A(n7008), .B(n7009), .Z(n6931) );
  XNOR2_X1 U8601 ( .A(n7002), .B(P2_REG1_REG_7__SCAN_IN), .ZN(n6929) );
  INV_X1 U8602 ( .A(n6924), .ZN(n6923) );
  INV_X1 U8603 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n7099) );
  NAND2_X1 U8604 ( .A1(n6923), .A2(n7099), .ZN(n6925) );
  AOI21_X1 U8605 ( .B1(n6925), .B2(n7018), .A(n9736), .ZN(n6928) );
  INV_X1 U8606 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n10042) );
  NOR2_X1 U8607 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10042), .ZN(n6942) );
  AOI21_X1 U8608 ( .B1(n9200), .B2(P2_ADDR_REG_7__SCAN_IN), .A(n6942), .ZN(
        n6926) );
  OAI21_X1 U8609 ( .B1(n4532), .B2(n9721), .A(n6926), .ZN(n6927) );
  AOI211_X1 U8610 ( .C1(n6929), .C2(n9730), .A(n6928), .B(n6927), .ZN(n6930)
         );
  OAI21_X1 U8611 ( .B1(n6931), .B2(n4472), .A(n6930), .ZN(P2_U3189) );
  AND2_X1 U8612 ( .A1(n8756), .A2(n7029), .ZN(n8667) );
  OR2_X1 U8613 ( .A1(n8667), .A2(n6932), .ZN(n9514) );
  INV_X1 U8614 ( .A(n6933), .ZN(n6935) );
  NOR2_X1 U8615 ( .A1(n6934), .A2(n9060), .ZN(n9518) );
  AOI21_X1 U8616 ( .B1(n9514), .B2(n6935), .A(n9518), .ZN(n6938) );
  INV_X1 U8617 ( .A(n9499), .ZN(n9471) );
  AOI22_X1 U8618 ( .A1(n9485), .A2(P1_REG2_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(n9471), .ZN(n6937) );
  NAND2_X1 U8619 ( .A1(n9480), .A2(n9496), .ZN(n8887) );
  INV_X1 U8620 ( .A(n8887), .ZN(n9037) );
  OAI21_X1 U8621 ( .B1(n9037), .B2(n9472), .A(n9519), .ZN(n6936) );
  OAI211_X1 U8622 ( .C1(n6938), .C2(n9485), .A(n6937), .B(n6936), .ZN(P1_U3293) );
  OAI21_X1 U8623 ( .B1(n6941), .B2(n6940), .A(n6939), .ZN(n6947) );
  NOR2_X1 U8624 ( .A1(n7991), .A2(n9808), .ZN(n6946) );
  NAND2_X1 U8625 ( .A1(n7987), .A2(n7097), .ZN(n6944) );
  AOI21_X1 U8626 ( .B1(n8002), .B2(n7968), .A(n6942), .ZN(n6943) );
  OAI211_X1 U8627 ( .C1(n7091), .C2(n7971), .A(n6944), .B(n6943), .ZN(n6945)
         );
  AOI211_X1 U8628 ( .C1(n6947), .C2(n7954), .A(n6946), .B(n6945), .ZN(n6948)
         );
  INV_X1 U8629 ( .A(n6948), .ZN(P2_U3153) );
  INV_X1 U8630 ( .A(n6949), .ZN(n6951) );
  NAND2_X1 U8631 ( .A1(n6951), .A2(n6950), .ZN(n6952) );
  XNOR2_X1 U8632 ( .A(n6953), .B(n6952), .ZN(n6958) );
  NAND2_X1 U8633 ( .A1(n7987), .A2(n6994), .ZN(n6955) );
  NOR2_X1 U8634 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9940), .ZN(n7011) );
  AOI21_X1 U8635 ( .B1(n8001), .B2(n7968), .A(n7011), .ZN(n6954) );
  OAI211_X1 U8636 ( .C1(n6986), .C2(n7971), .A(n6955), .B(n6954), .ZN(n6956)
         );
  AOI21_X1 U8637 ( .B1(n9814), .B2(n7973), .A(n6956), .ZN(n6957) );
  OAI21_X1 U8638 ( .B1(n6958), .B2(n7977), .A(n6957), .ZN(P2_U3161) );
  NAND2_X1 U8639 ( .A1(n6960), .A2(n6959), .ZN(n6962) );
  XNOR2_X1 U8640 ( .A(n6962), .B(n6961), .ZN(n6968) );
  INV_X1 U8641 ( .A(n7053), .ZN(n6964) );
  OR2_X1 U8642 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6963), .ZN(n9334) );
  OAI21_X1 U8643 ( .B1(n8458), .B2(n6964), .A(n9334), .ZN(n6966) );
  OAI22_X1 U8644 ( .A1(n8407), .A2(n9548), .B1(n8426), .B2(n6970), .ZN(n6965)
         );
  AOI211_X1 U8645 ( .C1(n8454), .C2(n8753), .A(n6966), .B(n6965), .ZN(n6967)
         );
  OAI21_X1 U8646 ( .B1(n6968), .B2(n8462), .A(n6967), .ZN(P1_U3227) );
  NAND2_X1 U8647 ( .A1(n6971), .A2(n8672), .ZN(n7043) );
  XNOR2_X1 U8648 ( .A(n7042), .B(n7043), .ZN(n6972) );
  OAI222_X1 U8649 ( .A1(n9060), .A2(n7160), .B1(n9062), .B2(n6896), .C1(n6972), 
        .C2(n9516), .ZN(n9542) );
  INV_X1 U8650 ( .A(n9542), .ZN(n6983) );
  NAND2_X1 U8651 ( .A1(n6973), .A2(n8627), .ZN(n7048) );
  NAND2_X1 U8652 ( .A1(n6896), .A2(n6974), .ZN(n7046) );
  NAND2_X1 U8653 ( .A1(n7048), .A2(n7046), .ZN(n6975) );
  XNOR2_X1 U8654 ( .A(n7042), .B(n6975), .ZN(n9544) );
  OAI211_X1 U8655 ( .C1(n4369), .C2(n9541), .A(n6976), .B(n9496), .ZN(n9540)
         );
  AOI22_X1 U8656 ( .A1(n9485), .A2(P1_REG2_REG_4__SCAN_IN), .B1(n6977), .B2(
        n9471), .ZN(n6980) );
  NAND2_X1 U8657 ( .A1(n9472), .A2(n6978), .ZN(n6979) );
  OAI211_X1 U8658 ( .C1(n9540), .C2(n9085), .A(n6980), .B(n6979), .ZN(n6981)
         );
  AOI21_X1 U8659 ( .B1(n9544), .B2(n9482), .A(n6981), .ZN(n6982) );
  OAI21_X1 U8660 ( .B1(n6983), .B2(n9485), .A(n6982), .ZN(P1_U3289) );
  OAI211_X1 U8661 ( .C1(n6985), .C2(n6992), .A(n6984), .B(n9765), .ZN(n6989)
         );
  OAI22_X1 U8662 ( .A1(n6986), .A2(n9762), .B1(n7282), .B2(n9760), .ZN(n6987)
         );
  INV_X1 U8663 ( .A(n6987), .ZN(n6988) );
  NAND2_X1 U8664 ( .A1(n6989), .A2(n6988), .ZN(n9817) );
  INV_X1 U8665 ( .A(n9817), .ZN(n6999) );
  NAND2_X1 U8666 ( .A1(n6990), .A2(n6991), .ZN(n6993) );
  XNOR2_X1 U8667 ( .A(n6993), .B(n6992), .ZN(n9813) );
  INV_X1 U8668 ( .A(n9814), .ZN(n6996) );
  AOI22_X1 U8669 ( .A1(n9777), .A2(P2_REG2_REG_8__SCAN_IN), .B1(n9770), .B2(
        n6994), .ZN(n6995) );
  OAI21_X1 U8670 ( .B1(n6996), .B2(n8076), .A(n6995), .ZN(n6997) );
  AOI21_X1 U8671 ( .B1(n9813), .B2(n9753), .A(n6997), .ZN(n6998) );
  OAI21_X1 U8672 ( .B1(n6999), .B2(n9777), .A(n6998), .ZN(P2_U3225) );
  INV_X1 U8673 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n9847) );
  MUX2_X1 U8674 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n9847), .S(n7023), .Z(n7004)
         );
  INV_X1 U8675 ( .A(n7000), .ZN(n7001) );
  AOI21_X1 U8676 ( .B1(n7004), .B2(n7003), .A(n7121), .ZN(n7026) );
  INV_X1 U8677 ( .A(n7005), .ZN(n7006) );
  MUX2_X1 U8678 ( .A(P2_REG2_REG_8__SCAN_IN), .B(P2_REG1_REG_8__SCAN_IN), .S(
        n8046), .Z(n7123) );
  XOR2_X1 U8679 ( .A(n7023), .B(n7123), .Z(n7124) );
  XNOR2_X1 U8680 ( .A(n7125), .B(n7124), .ZN(n7010) );
  NAND2_X1 U8681 ( .A1(n7010), .A2(n9729), .ZN(n7025) );
  INV_X1 U8682 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n7013) );
  INV_X1 U8683 ( .A(n7011), .ZN(n7012) );
  OAI21_X1 U8684 ( .B1(n9720), .B2(n7013), .A(n7012), .ZN(n7022) );
  INV_X1 U8685 ( .A(n7014), .ZN(n7016) );
  INV_X1 U8686 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7015) );
  MUX2_X1 U8687 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n7015), .S(n7023), .Z(n7017)
         );
  INV_X1 U8688 ( .A(n7136), .ZN(n7020) );
  NAND3_X1 U8689 ( .A1(n7018), .A2(n7017), .A3(n7016), .ZN(n7019) );
  AOI21_X1 U8690 ( .B1(n7020), .B2(n7019), .A(n9736), .ZN(n7021) );
  AOI211_X1 U8691 ( .C1(n7142), .C2(n7023), .A(n7022), .B(n7021), .ZN(n7024)
         );
  OAI211_X1 U8692 ( .C1(n7026), .C2(n8066), .A(n7025), .B(n7024), .ZN(P2_U3190) );
  XNOR2_X1 U8693 ( .A(n7027), .B(n7028), .ZN(n9524) );
  INV_X1 U8694 ( .A(n7217), .ZN(n9506) );
  AOI22_X1 U8695 ( .A1(n9472), .A2(n7030), .B1(n9471), .B2(
        P1_REG3_REG_1__SCAN_IN), .ZN(n7031) );
  OAI21_X1 U8696 ( .B1(n9085), .B2(n9521), .A(n7031), .ZN(n7040) );
  NAND2_X1 U8697 ( .A1(n9524), .A2(n9597), .ZN(n7038) );
  AOI22_X1 U8698 ( .A1(n9489), .A2(n8756), .B1(n8754), .B2(n9490), .ZN(n7037)
         );
  INV_X1 U8699 ( .A(n6932), .ZN(n7032) );
  NAND2_X1 U8700 ( .A1(n7032), .A2(n7028), .ZN(n7034) );
  NAND2_X1 U8701 ( .A1(n7034), .A2(n7033), .ZN(n7035) );
  NAND2_X1 U8702 ( .A1(n7035), .A2(n9493), .ZN(n7036) );
  NAND3_X1 U8703 ( .A1(n7038), .A2(n7037), .A3(n7036), .ZN(n9522) );
  MUX2_X1 U8704 ( .A(n9522), .B(P1_REG2_REG_1__SCAN_IN), .S(n9485), .Z(n7039)
         );
  AOI211_X1 U8705 ( .C1(n9524), .C2(n9506), .A(n7040), .B(n7039), .ZN(n7041)
         );
  INV_X1 U8706 ( .A(n7041), .ZN(P1_U3292) );
  NAND2_X1 U8707 ( .A1(n7043), .A2(n7049), .ZN(n7044) );
  NAND2_X1 U8708 ( .A1(n7044), .A2(n8477), .ZN(n7149) );
  XNOR2_X1 U8709 ( .A(n7154), .B(n7149), .ZN(n7045) );
  OAI222_X1 U8710 ( .A1(n9060), .A2(n7164), .B1(n9062), .B2(n6970), .C1(n7045), 
        .C2(n9516), .ZN(n9549) );
  INV_X1 U8711 ( .A(n9549), .ZN(n7059) );
  NAND2_X1 U8712 ( .A1(n6970), .A2(n9541), .ZN(n7050) );
  AND2_X1 U8713 ( .A1(n7046), .A2(n7050), .ZN(n7047) );
  NAND2_X1 U8714 ( .A1(n7048), .A2(n7047), .ZN(n7159) );
  AND2_X1 U8715 ( .A1(n7159), .A2(n7155), .ZN(n7051) );
  XNOR2_X1 U8716 ( .A(n7154), .B(n7051), .ZN(n9551) );
  INV_X1 U8717 ( .A(n6976), .ZN(n7052) );
  OAI211_X1 U8718 ( .C1(n7052), .C2(n9548), .A(n9496), .B(n9476), .ZN(n9547)
         );
  AOI22_X1 U8719 ( .A1(n9485), .A2(P1_REG2_REG_5__SCAN_IN), .B1(n7053), .B2(
        n9471), .ZN(n7056) );
  NAND2_X1 U8720 ( .A1(n9472), .A2(n7054), .ZN(n7055) );
  OAI211_X1 U8721 ( .C1(n9547), .C2(n9085), .A(n7056), .B(n7055), .ZN(n7057)
         );
  AOI21_X1 U8722 ( .B1(n9551), .B2(n9482), .A(n7057), .ZN(n7058) );
  OAI21_X1 U8723 ( .B1(n7059), .B2(n9485), .A(n7058), .ZN(P1_U3288) );
  INV_X1 U8724 ( .A(n7060), .ZN(n7062) );
  INV_X1 U8725 ( .A(n7817), .ZN(n7615) );
  INV_X1 U8726 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7061) );
  OAI222_X1 U8727 ( .A1(n8328), .A2(n7062), .B1(n9917), .B2(n7615), .C1(n7061), 
        .C2(n7118), .ZN(P2_U3273) );
  OAI222_X1 U8728 ( .A1(n9195), .A2(n7063), .B1(n9193), .B2(n7062), .C1(n8658), 
        .C2(P1_U3086), .ZN(P1_U3333) );
  INV_X1 U8729 ( .A(n7076), .ZN(n7065) );
  NAND2_X1 U8730 ( .A1(n8326), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n7064) );
  OAI211_X1 U8731 ( .C1(n7065), .C2(n8328), .A(n7819), .B(n7064), .ZN(P2_U3272) );
  NAND2_X1 U8732 ( .A1(n7066), .A2(n7067), .ZN(n7106) );
  OAI21_X1 U8733 ( .B1(n7067), .B2(n7066), .A(n7106), .ZN(n7073) );
  AOI22_X1 U8734 ( .A1(n8455), .A2(n7068), .B1(n9473), .B2(n8460), .ZN(n7071)
         );
  NAND2_X1 U8735 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n9348) );
  INV_X1 U8736 ( .A(n9348), .ZN(n7069) );
  AOI21_X1 U8737 ( .B1(n8446), .B2(n9470), .A(n7069), .ZN(n7070) );
  OAI211_X1 U8738 ( .C1(n8483), .C2(n8427), .A(n7071), .B(n7070), .ZN(n7072)
         );
  AOI21_X1 U8739 ( .B1(n7073), .B2(n8444), .A(n7072), .ZN(n7074) );
  INV_X1 U8740 ( .A(n7074), .ZN(P1_U3239) );
  NAND2_X1 U8741 ( .A1(n7076), .A2(n7075), .ZN(n7077) );
  OAI211_X1 U8742 ( .C1(n7078), .C2(n7858), .A(n7077), .B(n8732), .ZN(P1_U3332) );
  OAI211_X1 U8743 ( .C1(n7081), .C2(n7080), .A(n7079), .B(n7954), .ZN(n7086)
         );
  NAND2_X1 U8744 ( .A1(n7987), .A2(n7196), .ZN(n7083) );
  NOR2_X1 U8745 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5336), .ZN(n7133) );
  AOI21_X1 U8746 ( .B1(n8000), .B2(n7968), .A(n7133), .ZN(n7082) );
  OAI211_X1 U8747 ( .C1(n7090), .C2(n7971), .A(n7083), .B(n7082), .ZN(n7084)
         );
  AOI21_X1 U8748 ( .B1(n9823), .B2(n7973), .A(n7084), .ZN(n7085) );
  NAND2_X1 U8749 ( .A1(n7086), .A2(n7085), .ZN(P2_U3171) );
  OR2_X1 U8750 ( .A1(n7087), .A2(n7779), .ZN(n7088) );
  AND2_X1 U8751 ( .A1(n6990), .A2(n7088), .ZN(n7094) );
  INV_X1 U8752 ( .A(n7094), .ZN(n9809) );
  XNOR2_X1 U8753 ( .A(n7089), .B(n7779), .ZN(n7096) );
  OAI22_X1 U8754 ( .A1(n7091), .A2(n9762), .B1(n7090), .B2(n9760), .ZN(n7092)
         );
  AOI21_X1 U8755 ( .B1(n7094), .B2(n7093), .A(n7092), .ZN(n7095) );
  OAI21_X1 U8756 ( .B1(n7096), .B2(n7505), .A(n7095), .ZN(n9811) );
  NAND2_X1 U8757 ( .A1(n9811), .A2(n9775), .ZN(n7103) );
  INV_X1 U8758 ( .A(n7097), .ZN(n7098) );
  OAI22_X1 U8759 ( .A1(n9775), .A2(n7099), .B1(n7098), .B2(n7377), .ZN(n7100)
         );
  AOI21_X1 U8760 ( .B1(n9751), .B2(n7101), .A(n7100), .ZN(n7102) );
  OAI211_X1 U8761 ( .C1(n9809), .C2(n7202), .A(n7103), .B(n7102), .ZN(P2_U3226) );
  NAND2_X1 U8762 ( .A1(n7106), .A2(n7104), .ZN(n7111) );
  NAND2_X1 U8763 ( .A1(n7106), .A2(n7105), .ZN(n7107) );
  OAI21_X1 U8764 ( .B1(n7110), .B2(n7108), .A(n7107), .ZN(n7109) );
  OAI211_X1 U8765 ( .C1(n7111), .C2(n7110), .A(n8444), .B(n7109), .ZN(n7116)
         );
  INV_X1 U8766 ( .A(n7112), .ZN(n7209) );
  NAND2_X1 U8767 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3086), .ZN(n9245) );
  OAI21_X1 U8768 ( .B1(n8458), .B2(n7209), .A(n9245), .ZN(n7114) );
  OAI22_X1 U8769 ( .A1(n8490), .A2(n8427), .B1(n8426), .B2(n7164), .ZN(n7113)
         );
  AOI211_X1 U8770 ( .C1(n8491), .C2(n8430), .A(n7114), .B(n7113), .ZN(n7115)
         );
  NAND2_X1 U8771 ( .A1(n7116), .A2(n7115), .ZN(P1_U3213) );
  INV_X1 U8772 ( .A(n7117), .ZN(n7147) );
  INV_X1 U8773 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7119) );
  OAI222_X1 U8774 ( .A1(n8328), .A2(n7147), .B1(P2_U3151), .B2(n7120), .C1(
        n7119), .C2(n7118), .ZN(P2_U3271) );
  AOI21_X1 U8775 ( .B1(n7137), .B2(P2_REG1_REG_8__SCAN_IN), .A(n7121), .ZN(
        n7290) );
  INV_X1 U8776 ( .A(n7290), .ZN(n7122) );
  XNOR2_X1 U8777 ( .A(n7122), .B(n7295), .ZN(n7287) );
  XNOR2_X1 U8778 ( .A(n7287), .B(P2_REG1_REG_9__SCAN_IN), .ZN(n7145) );
  OAI22_X1 U8779 ( .A1(n7125), .A2(n7124), .B1(n7123), .B2(n7137), .ZN(n7129)
         );
  MUX2_X1 U8780 ( .A(P2_REG2_REG_9__SCAN_IN), .B(P2_REG1_REG_9__SCAN_IN), .S(
        n8057), .Z(n7126) );
  NAND2_X1 U8781 ( .A1(n7126), .A2(n7295), .ZN(n7130) );
  NAND2_X1 U8782 ( .A1(n7129), .A2(n7130), .ZN(n7303) );
  INV_X1 U8783 ( .A(n7126), .ZN(n7127) );
  NAND2_X1 U8784 ( .A1(n7127), .A2(n7289), .ZN(n7302) );
  INV_X1 U8785 ( .A(n7302), .ZN(n7128) );
  NOR2_X1 U8786 ( .A1(n7303), .A2(n7128), .ZN(n7132) );
  AOI21_X1 U8787 ( .B1(n7130), .B2(n7302), .A(n7129), .ZN(n7131) );
  OAI21_X1 U8788 ( .B1(n7132), .B2(n7131), .A(n9729), .ZN(n7144) );
  INV_X1 U8789 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n7135) );
  INV_X1 U8790 ( .A(n7133), .ZN(n7134) );
  OAI21_X1 U8791 ( .B1(n9720), .B2(n7135), .A(n7134), .ZN(n7141) );
  INV_X1 U8792 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7198) );
  AOI21_X1 U8793 ( .B1(P2_REG2_REG_8__SCAN_IN), .B2(n7137), .A(n7136), .ZN(
        n7293) );
  AOI21_X1 U8794 ( .B1(n7198), .B2(n7138), .A(n7294), .ZN(n7139) );
  NOR2_X1 U8795 ( .A1(n7139), .A2(n9736), .ZN(n7140) );
  AOI211_X1 U8796 ( .C1(n7142), .C2(n7289), .A(n7141), .B(n7140), .ZN(n7143)
         );
  OAI211_X1 U8797 ( .C1(n7145), .C2(n8066), .A(n7144), .B(n7143), .ZN(P2_U3191) );
  OAI222_X1 U8798 ( .A1(n7148), .A2(P1_U3086), .B1(n9193), .B2(n7147), .C1(
        n7146), .C2(n7858), .ZN(P1_U3331) );
  NAND2_X1 U8799 ( .A1(n7149), .A2(n7157), .ZN(n7150) );
  NAND2_X1 U8800 ( .A1(n8753), .A2(n9554), .ZN(n8471) );
  NAND2_X1 U8801 ( .A1(n7264), .A2(n8471), .ZN(n7204) );
  NAND2_X1 U8802 ( .A1(n8483), .A2(n8491), .ZN(n8481) );
  INV_X1 U8803 ( .A(n8483), .ZN(n9468) );
  NAND2_X1 U8804 ( .A1(n9468), .A2(n9561), .ZN(n8474) );
  OAI21_X1 U8805 ( .B1(n7204), .B2(n7205), .A(n8481), .ZN(n7231) );
  NAND2_X1 U8806 ( .A1(n8490), .A2(n8486), .ZN(n8482) );
  NAND2_X1 U8807 ( .A1(n8482), .A2(n8475), .ZN(n7237) );
  INV_X1 U8808 ( .A(n7237), .ZN(n7151) );
  XNOR2_X1 U8809 ( .A(n7231), .B(n7151), .ZN(n7153) );
  OAI22_X1 U8810 ( .A1(n8483), .A2(n9062), .B1(n7471), .B2(n9060), .ZN(n7152)
         );
  AOI21_X1 U8811 ( .B1(n7153), .B2(n9493), .A(n7152), .ZN(n9573) );
  INV_X1 U8812 ( .A(n7154), .ZN(n7157) );
  INV_X1 U8813 ( .A(n7155), .ZN(n7156) );
  NAND2_X1 U8814 ( .A1(n7159), .A2(n7158), .ZN(n7162) );
  NAND2_X1 U8815 ( .A1(n7160), .A2(n9548), .ZN(n7161) );
  NAND2_X1 U8816 ( .A1(n7162), .A2(n7161), .ZN(n9474) );
  NAND2_X1 U8817 ( .A1(n9474), .A2(n9475), .ZN(n7166) );
  NAND2_X1 U8818 ( .A1(n7164), .A2(n9554), .ZN(n7165) );
  NAND2_X1 U8819 ( .A1(n7166), .A2(n7165), .ZN(n7203) );
  NAND2_X1 U8820 ( .A1(n7203), .A2(n7205), .ZN(n7168) );
  NAND2_X1 U8821 ( .A1(n8483), .A2(n9561), .ZN(n7167) );
  NAND2_X1 U8822 ( .A1(n7168), .A2(n7167), .ZN(n7238) );
  XNOR2_X1 U8823 ( .A(n7238), .B(n7237), .ZN(n9571) );
  OR2_X1 U8824 ( .A1(n7211), .A2(n9567), .ZN(n7169) );
  NAND2_X1 U8825 ( .A1(n7239), .A2(n7169), .ZN(n9569) );
  AOI22_X1 U8826 ( .A1(n9485), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n7255), .B2(
        n9471), .ZN(n7171) );
  NAND2_X1 U8827 ( .A1(n9472), .A2(n8486), .ZN(n7170) );
  OAI211_X1 U8828 ( .C1(n9569), .C2(n8887), .A(n7171), .B(n7170), .ZN(n7172)
         );
  AOI21_X1 U8829 ( .B1(n9571), .B2(n9482), .A(n7172), .ZN(n7173) );
  OAI21_X1 U8830 ( .B1(n9573), .B2(n9485), .A(n7173), .ZN(P1_U3285) );
  XOR2_X1 U8831 ( .A(n7784), .B(n7174), .Z(n7175) );
  OAI222_X1 U8832 ( .A1(n9762), .A2(n7282), .B1(n9760), .B2(n7451), .C1(n7505), 
        .C2(n7175), .ZN(n7181) );
  INV_X1 U8833 ( .A(n7181), .ZN(n7180) );
  NAND2_X1 U8834 ( .A1(n7189), .A2(n7649), .ZN(n7176) );
  XNOR2_X1 U8835 ( .A(n7176), .B(n7784), .ZN(n7182) );
  INV_X1 U8836 ( .A(n7284), .ZN(n7185) );
  AOI22_X1 U8837 ( .A1(n9777), .A2(P2_REG2_REG_10__SCAN_IN), .B1(n9770), .B2(
        n7279), .ZN(n7177) );
  OAI21_X1 U8838 ( .B1(n7185), .B2(n8076), .A(n7177), .ZN(n7178) );
  AOI21_X1 U8839 ( .B1(n7182), .B2(n9753), .A(n7178), .ZN(n7179) );
  OAI21_X1 U8840 ( .B1(n7180), .B2(n9777), .A(n7179), .ZN(P2_U3223) );
  AOI21_X1 U8841 ( .B1(n9831), .B2(n7182), .A(n7181), .ZN(n7188) );
  AOI22_X1 U8842 ( .A1(n7284), .A2(n8245), .B1(n9852), .B2(
        P2_REG1_REG_10__SCAN_IN), .ZN(n7183) );
  OAI21_X1 U8843 ( .B1(n7188), .B2(n9852), .A(n7183), .ZN(P2_U3469) );
  INV_X1 U8844 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n7184) );
  OAI22_X1 U8845 ( .A1(n7185), .A2(n8254), .B1(n9836), .B2(n7184), .ZN(n7186)
         );
  INV_X1 U8846 ( .A(n7186), .ZN(n7187) );
  OAI21_X1 U8847 ( .B1(n7188), .B2(n9838), .A(n7187), .ZN(P2_U3420) );
  OAI21_X1 U8848 ( .B1(n7190), .B2(n5711), .A(n7189), .ZN(n9820) );
  OAI21_X1 U8849 ( .B1(n7192), .B2(n7783), .A(n7191), .ZN(n7193) );
  NAND2_X1 U8850 ( .A1(n7193), .A2(n9765), .ZN(n7195) );
  AOI22_X1 U8851 ( .A1(n9744), .A2(n8002), .B1(n8000), .B2(n9746), .ZN(n7194)
         );
  OAI211_X1 U8852 ( .C1(n9768), .C2(n9820), .A(n7195), .B(n7194), .ZN(n9821)
         );
  NAND2_X1 U8853 ( .A1(n9821), .A2(n9775), .ZN(n7201) );
  INV_X1 U8854 ( .A(n7196), .ZN(n7197) );
  OAI22_X1 U8855 ( .A1(n9775), .A2(n7198), .B1(n7197), .B2(n7377), .ZN(n7199)
         );
  AOI21_X1 U8856 ( .B1(n9751), .B2(n9823), .A(n7199), .ZN(n7200) );
  OAI211_X1 U8857 ( .C1(n9820), .C2(n7202), .A(n7201), .B(n7200), .ZN(P2_U3224) );
  XNOR2_X1 U8858 ( .A(n7203), .B(n7205), .ZN(n9564) );
  INV_X1 U8859 ( .A(n9564), .ZN(n7218) );
  XOR2_X1 U8860 ( .A(n7205), .B(n7204), .Z(n7208) );
  AOI22_X1 U8861 ( .A1(n9490), .A2(n8752), .B1(n8753), .B2(n9489), .ZN(n7207)
         );
  NAND2_X1 U8862 ( .A1(n9564), .A2(n9597), .ZN(n7206) );
  OAI211_X1 U8863 ( .C1(n7208), .C2(n9516), .A(n7207), .B(n7206), .ZN(n9562)
         );
  NAND2_X1 U8864 ( .A1(n9562), .A2(n9510), .ZN(n7216) );
  INV_X1 U8865 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n7210) );
  OAI22_X1 U8866 ( .A1(n9510), .A2(n7210), .B1(n7209), .B2(n9499), .ZN(n7214)
         );
  INV_X1 U8867 ( .A(n7211), .ZN(n7212) );
  OAI211_X1 U8868 ( .C1(n9561), .C2(n9477), .A(n7212), .B(n9496), .ZN(n9560)
         );
  NOR2_X1 U8869 ( .A1(n9560), .A2(n9085), .ZN(n7213) );
  AOI211_X1 U8870 ( .C1(n9472), .C2(n8491), .A(n7214), .B(n7213), .ZN(n7215)
         );
  OAI211_X1 U8871 ( .C1(n7218), .C2(n7217), .A(n7216), .B(n7215), .ZN(P1_U3286) );
  XNOR2_X1 U8872 ( .A(n7219), .B(n7782), .ZN(n7222) );
  NAND2_X1 U8873 ( .A1(n7998), .A2(n9746), .ZN(n7220) );
  OAI21_X1 U8874 ( .B1(n7389), .B2(n9762), .A(n7220), .ZN(n7221) );
  AOI21_X1 U8875 ( .B1(n7222), .B2(n9765), .A(n7221), .ZN(n9828) );
  XNOR2_X1 U8876 ( .A(n7223), .B(n7782), .ZN(n9826) );
  AOI22_X1 U8877 ( .A1(n9777), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n9770), .B2(
        n7391), .ZN(n7224) );
  OAI21_X1 U8878 ( .B1(n7394), .B2(n8076), .A(n7224), .ZN(n7225) );
  AOI21_X1 U8879 ( .B1(n9826), .B2(n9753), .A(n7225), .ZN(n7226) );
  OAI21_X1 U8880 ( .B1(n9828), .B2(n9777), .A(n7226), .ZN(P2_U3222) );
  INV_X1 U8881 ( .A(n7227), .ZN(n7247) );
  AOI22_X1 U8882 ( .A1(n7228), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_25__SCAN_IN), .B2(n8326), .ZN(n7229) );
  OAI21_X1 U8883 ( .B1(n7247), .B2(n8328), .A(n7229), .ZN(P2_U3270) );
  INV_X1 U8884 ( .A(n8482), .ZN(n7230) );
  OAI21_X1 U8885 ( .B1(n7231), .B2(n7230), .A(n8475), .ZN(n7233) );
  NAND2_X1 U8886 ( .A1(n7471), .A2(n7343), .ZN(n8506) );
  NAND2_X1 U8887 ( .A1(n8751), .A2(n9576), .ZN(n8501) );
  INV_X1 U8888 ( .A(n7273), .ZN(n7232) );
  XNOR2_X1 U8889 ( .A(n7233), .B(n7232), .ZN(n7235) );
  NOR2_X1 U8890 ( .A1(n8490), .A2(n9062), .ZN(n7234) );
  AOI21_X1 U8891 ( .B1(n7235), .B2(n9493), .A(n7234), .ZN(n9580) );
  NOR2_X1 U8892 ( .A1(n8752), .A2(n8486), .ZN(n7236) );
  AOI21_X2 U8893 ( .B1(n7238), .B2(n7237), .A(n7236), .ZN(n7274) );
  XNOR2_X1 U8894 ( .A(n7274), .B(n7273), .ZN(n9578) );
  XNOR2_X1 U8895 ( .A(n7239), .B(n9576), .ZN(n7241) );
  NOR2_X1 U8896 ( .A1(n8750), .A2(n9060), .ZN(n7240) );
  AOI21_X1 U8897 ( .B1(n7241), .B2(n9496), .A(n7240), .ZN(n9575) );
  AOI22_X1 U8898 ( .A1(n9485), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n7339), .B2(
        n9471), .ZN(n7243) );
  NAND2_X1 U8899 ( .A1(n9472), .A2(n7343), .ZN(n7242) );
  OAI211_X1 U8900 ( .C1(n9575), .C2(n9085), .A(n7243), .B(n7242), .ZN(n7244)
         );
  AOI21_X1 U8901 ( .B1(n9578), .B2(n9482), .A(n7244), .ZN(n7245) );
  OAI21_X1 U8902 ( .B1(n9580), .B2(n9485), .A(n7245), .ZN(P1_U3284) );
  OAI222_X1 U8903 ( .A1(n7248), .A2(P1_U3086), .B1(n9193), .B2(n7247), .C1(
        n7246), .C2(n7858), .ZN(P1_U3330) );
  OAI21_X1 U8904 ( .B1(n7249), .B2(n7251), .A(n7250), .ZN(n7252) );
  NAND2_X1 U8905 ( .A1(n7252), .A2(n8444), .ZN(n7257) );
  NAND2_X1 U8906 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_U3086), .ZN(n9260) );
  INV_X1 U8907 ( .A(n9260), .ZN(n7254) );
  OAI22_X1 U8908 ( .A1(n8483), .A2(n8426), .B1(n8427), .B2(n7471), .ZN(n7253)
         );
  AOI211_X1 U8909 ( .C1(n7255), .C2(n8446), .A(n7254), .B(n7253), .ZN(n7256)
         );
  OAI211_X1 U8910 ( .C1(n9567), .C2(n8407), .A(n7257), .B(n7256), .ZN(P1_U3221) );
  INV_X1 U8911 ( .A(n7258), .ZN(n7335) );
  AOI22_X1 U8912 ( .A1(n7259), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_26__SCAN_IN), .B2(n8326), .ZN(n7260) );
  OAI21_X1 U8913 ( .B1(n7335), .B2(n8328), .A(n7260), .ZN(P2_U3269) );
  NAND3_X1 U8914 ( .A1(n8506), .A2(n8482), .A3(n8481), .ZN(n8632) );
  NAND2_X1 U8915 ( .A1(n8501), .A2(n8475), .ZN(n7262) );
  INV_X1 U8916 ( .A(n7262), .ZN(n7261) );
  NAND2_X1 U8917 ( .A1(n7262), .A2(n8506), .ZN(n7263) );
  NAND2_X1 U8918 ( .A1(n8632), .A2(n7263), .ZN(n8681) );
  OR2_X1 U8919 ( .A1(n8750), .A2(n7475), .ZN(n8684) );
  NAND2_X1 U8920 ( .A1(n7475), .A2(n8750), .ZN(n8508) );
  NAND2_X1 U8921 ( .A1(n8684), .A2(n8508), .ZN(n7360) );
  OAI21_X1 U8922 ( .B1(n4444), .B2(n4628), .A(n7362), .ZN(n7265) );
  INV_X1 U8923 ( .A(n7472), .ZN(n8749) );
  AOI222_X1 U8924 ( .A1(n9493), .A2(n7265), .B1(n8751), .B2(n9489), .C1(n8749), 
        .C2(n9490), .ZN(n9583) );
  INV_X1 U8925 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n7267) );
  INV_X1 U8926 ( .A(n7266), .ZN(n7470) );
  OAI22_X1 U8927 ( .A1(n9510), .A2(n7267), .B1(n7470), .B2(n9499), .ZN(n7272)
         );
  INV_X1 U8928 ( .A(n7475), .ZN(n9584) );
  INV_X1 U8929 ( .A(n7268), .ZN(n7270) );
  INV_X1 U8930 ( .A(n7269), .ZN(n7367) );
  OAI211_X1 U8931 ( .C1(n9584), .C2(n7270), .A(n7367), .B(n9496), .ZN(n9582)
         );
  NOR2_X1 U8932 ( .A1(n9582), .A2(n9085), .ZN(n7271) );
  AOI211_X1 U8933 ( .C1(n9472), .C2(n7475), .A(n7272), .B(n7271), .ZN(n7276)
         );
  XNOR2_X1 U8934 ( .A(n7361), .B(n7360), .ZN(n9586) );
  NAND2_X1 U8935 ( .A1(n9586), .A2(n9482), .ZN(n7275) );
  OAI211_X1 U8936 ( .C1(n9583), .C2(n9485), .A(n7276), .B(n7275), .ZN(P1_U3283) );
  XOR2_X1 U8937 ( .A(n7277), .B(n7278), .Z(n7286) );
  NAND2_X1 U8938 ( .A1(n7987), .A2(n7279), .ZN(n7281) );
  INV_X1 U8939 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n10036) );
  NOR2_X1 U8940 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10036), .ZN(n7306) );
  AOI21_X1 U8941 ( .B1(n7999), .B2(n7968), .A(n7306), .ZN(n7280) );
  OAI211_X1 U8942 ( .C1(n7282), .C2(n7971), .A(n7281), .B(n7280), .ZN(n7283)
         );
  AOI21_X1 U8943 ( .B1(n7284), .B2(n7973), .A(n7283), .ZN(n7285) );
  OAI21_X1 U8944 ( .B1(n7286), .B2(n7977), .A(n7285), .ZN(P2_U3157) );
  INV_X1 U8945 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n7288) );
  INV_X1 U8946 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n7319) );
  AOI22_X1 U8947 ( .A1(n7320), .A2(n7319), .B1(P2_REG1_REG_10__SCAN_IN), .B2(
        n7323), .ZN(n7291) );
  OAI21_X1 U8948 ( .B1(n7292), .B2(n7291), .A(n7318), .ZN(n7311) );
  INV_X1 U8949 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7296) );
  AOI22_X1 U8950 ( .A1(n7320), .A2(P2_REG2_REG_10__SCAN_IN), .B1(n7296), .B2(
        n7323), .ZN(n7297) );
  AOI21_X1 U8951 ( .B1(n4443), .B2(n7297), .A(n7325), .ZN(n7309) );
  MUX2_X1 U8952 ( .A(n7296), .B(n7319), .S(n8046), .Z(n7298) );
  NAND2_X1 U8953 ( .A1(n7298), .A2(n7320), .ZN(n7313) );
  INV_X1 U8954 ( .A(n7298), .ZN(n7299) );
  NAND2_X1 U8955 ( .A1(n7299), .A2(n7323), .ZN(n7300) );
  NAND2_X1 U8956 ( .A1(n7313), .A2(n7300), .ZN(n7301) );
  AOI21_X1 U8957 ( .B1(n7303), .B2(n7302), .A(n7301), .ZN(n7315) );
  AND3_X1 U8958 ( .A1(n7303), .A2(n7302), .A3(n7301), .ZN(n7304) );
  OAI21_X1 U8959 ( .B1(n7315), .B2(n7304), .A(n9729), .ZN(n7308) );
  NOR2_X1 U8960 ( .A1(n9721), .A2(n7323), .ZN(n7305) );
  AOI211_X1 U8961 ( .C1(n9200), .C2(P2_ADDR_REG_10__SCAN_IN), .A(n7306), .B(
        n7305), .ZN(n7307) );
  OAI211_X1 U8962 ( .C1(n7309), .C2(n9736), .A(n7308), .B(n7307), .ZN(n7310)
         );
  AOI21_X1 U8963 ( .B1(n9730), .B2(n7311), .A(n7310), .ZN(n7312) );
  INV_X1 U8964 ( .A(n7312), .ZN(P2_U3192) );
  INV_X1 U8965 ( .A(n7313), .ZN(n7314) );
  NOR2_X1 U8966 ( .A1(n7315), .A2(n7314), .ZN(n7317) );
  MUX2_X1 U8967 ( .A(P2_REG2_REG_11__SCAN_IN), .B(P2_REG1_REG_11__SCAN_IN), 
        .S(n8057), .Z(n7415) );
  XNOR2_X1 U8968 ( .A(n7415), .B(n7427), .ZN(n7316) );
  NOR2_X1 U8969 ( .A1(n7317), .A2(n7316), .ZN(n7416) );
  AOI21_X1 U8970 ( .B1(n7317), .B2(n7316), .A(n7416), .ZN(n7333) );
  NAND2_X1 U8971 ( .A1(P2_REG1_REG_11__SCAN_IN), .A2(n7321), .ZN(n7428) );
  OAI21_X1 U8972 ( .B1(P2_REG1_REG_11__SCAN_IN), .B2(n7321), .A(n7428), .ZN(
        n7331) );
  INV_X1 U8973 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n9920) );
  NOR2_X1 U8974 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9920), .ZN(n7387) );
  AOI21_X1 U8975 ( .B1(n9200), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n7387), .ZN(
        n7322) );
  OAI21_X1 U8976 ( .B1(n7427), .B2(n9721), .A(n7322), .ZN(n7330) );
  INV_X1 U8977 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n7327) );
  NOR2_X1 U8978 ( .A1(n7325), .A2(n7324), .ZN(n7412) );
  XNOR2_X1 U8979 ( .A(n7412), .B(n7418), .ZN(n7326) );
  AOI21_X1 U8980 ( .B1(n7327), .B2(n7326), .A(n7413), .ZN(n7328) );
  NOR2_X1 U8981 ( .A1(n7328), .A2(n9736), .ZN(n7329) );
  AOI211_X1 U8982 ( .C1(n9730), .C2(n7331), .A(n7330), .B(n7329), .ZN(n7332)
         );
  OAI21_X1 U8983 ( .B1(n7333), .B2(n4472), .A(n7332), .ZN(P2_U3193) );
  OAI222_X1 U8984 ( .A1(n7336), .A2(P1_U3086), .B1(n9193), .B2(n7335), .C1(
        n7334), .C2(n7858), .ZN(P1_U3329) );
  XOR2_X1 U8985 ( .A(n7337), .B(n7338), .Z(n7345) );
  INV_X1 U8986 ( .A(n7339), .ZN(n7340) );
  NAND2_X1 U8987 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_U3086), .ZN(n9275) );
  OAI21_X1 U8988 ( .B1(n8458), .B2(n7340), .A(n9275), .ZN(n7342) );
  OAI22_X1 U8989 ( .A1(n8490), .A2(n8426), .B1(n8427), .B2(n8750), .ZN(n7341)
         );
  AOI211_X1 U8990 ( .C1(n7343), .C2(n8430), .A(n7342), .B(n7341), .ZN(n7344)
         );
  OAI21_X1 U8991 ( .B1(n7345), .B2(n8462), .A(n7344), .ZN(P1_U3231) );
  XNOR2_X1 U8992 ( .A(n7346), .B(n7350), .ZN(n7347) );
  OAI222_X1 U8993 ( .A1(n9760), .A2(n7348), .B1(n9762), .B2(n7451), .C1(n7505), 
        .C2(n7347), .ZN(n9832) );
  NAND2_X1 U8994 ( .A1(n7351), .A2(n7350), .ZN(n9830) );
  NAND3_X1 U8995 ( .A1(n7349), .A2(n9830), .A3(n9753), .ZN(n7353) );
  AOI22_X1 U8996 ( .A1(n9777), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n9770), .B2(
        n7453), .ZN(n7352) );
  OAI211_X1 U8997 ( .C1(n5501), .C2(n8076), .A(n7353), .B(n7352), .ZN(n7354)
         );
  AOI21_X1 U8998 ( .B1(n9832), .B2(n9775), .A(n7354), .ZN(n7355) );
  INV_X1 U8999 ( .A(n7355), .ZN(P2_U3221) );
  INV_X1 U9000 ( .A(n7356), .ZN(n7821) );
  AOI21_X1 U9001 ( .B1(n8326), .B2(P1_DATAO_REG_27__SCAN_IN), .A(n7357), .ZN(
        n7358) );
  OAI21_X1 U9002 ( .B1(n7821), .B2(n8328), .A(n7358), .ZN(P2_U3268) );
  NAND2_X1 U9003 ( .A1(n9590), .A2(n7472), .ZN(n8509) );
  XOR2_X1 U9004 ( .A(n8635), .B(n7409), .Z(n9594) );
  AND2_X1 U9005 ( .A1(n7362), .A2(n8508), .ZN(n7363) );
  NAND2_X1 U9006 ( .A1(n7363), .A2(n8635), .ZN(n7401) );
  OAI211_X1 U9007 ( .C1(n8635), .C2(n7363), .A(n7401), .B(n9493), .ZN(n7365)
         );
  NAND2_X1 U9008 ( .A1(n8748), .A2(n9490), .ZN(n7364) );
  OAI211_X1 U9009 ( .C1(n8750), .C2(n9062), .A(n7365), .B(n7364), .ZN(n9588)
         );
  AOI211_X1 U9010 ( .C1(n9590), .C2(n7367), .A(n9568), .B(n7366), .ZN(n9589)
         );
  NAND2_X1 U9011 ( .A1(n9589), .A2(n9480), .ZN(n7369) );
  AOI22_X1 U9012 ( .A1(n9485), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n7536), .B2(
        n9471), .ZN(n7368) );
  OAI211_X1 U9013 ( .C1(n4876), .C2(n9067), .A(n7369), .B(n7368), .ZN(n7370)
         );
  AOI21_X1 U9014 ( .B1(n9510), .B2(n9588), .A(n7370), .ZN(n7371) );
  OAI21_X1 U9015 ( .B1(n9594), .B2(n9071), .A(n7371), .ZN(P1_U3282) );
  INV_X1 U9016 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n9657) );
  AND2_X1 U9017 ( .A1(n7373), .A2(n7372), .ZN(n7682) );
  INV_X1 U9018 ( .A(n7682), .ZN(n7788) );
  XNOR2_X1 U9019 ( .A(n7374), .B(n7788), .ZN(n7375) );
  OAI222_X1 U9020 ( .A1(n9762), .A2(n5500), .B1(n9760), .B2(n7376), .C1(n7505), 
        .C2(n7375), .ZN(n9284) );
  INV_X1 U9021 ( .A(n9286), .ZN(n7379) );
  INV_X1 U9022 ( .A(n7524), .ZN(n7378) );
  OAI22_X1 U9023 ( .A1(n7379), .A2(n8120), .B1(n7378), .B2(n7377), .ZN(n7380)
         );
  OAI21_X1 U9024 ( .B1(n9284), .B2(n7380), .A(n9775), .ZN(n7383) );
  XNOR2_X1 U9025 ( .A(n7381), .B(n7682), .ZN(n9283) );
  NAND2_X1 U9026 ( .A1(n9283), .A2(n9753), .ZN(n7382) );
  OAI211_X1 U9027 ( .C1(n9657), .C2(n9775), .A(n7383), .B(n7382), .ZN(P2_U3220) );
  OAI211_X1 U9028 ( .C1(n7386), .C2(n5805), .A(n7954), .B(n7385), .ZN(n7393)
         );
  AOI21_X1 U9029 ( .B1(n7968), .B2(n7998), .A(n7387), .ZN(n7388) );
  OAI21_X1 U9030 ( .B1(n7389), .B2(n7971), .A(n7388), .ZN(n7390) );
  AOI21_X1 U9031 ( .B1(n7391), .B2(n7987), .A(n7390), .ZN(n7392) );
  OAI211_X1 U9032 ( .C1(n7394), .C2(n7991), .A(n7393), .B(n7392), .ZN(P2_U3176) );
  INV_X1 U9033 ( .A(n7395), .ZN(n7439) );
  AOI21_X1 U9034 ( .B1(n8326), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n7396), .ZN(
        n7397) );
  OAI21_X1 U9035 ( .B1(n7439), .B2(n8328), .A(n7397), .ZN(P2_U3267) );
  INV_X1 U9036 ( .A(n7401), .ZN(n7398) );
  INV_X1 U9037 ( .A(n8511), .ZN(n7399) );
  NAND2_X1 U9038 ( .A1(n9601), .A2(n8748), .ZN(n8512) );
  NAND2_X1 U9039 ( .A1(n7464), .A2(n7538), .ZN(n8693) );
  OAI21_X1 U9040 ( .B1(n7398), .B2(n7399), .A(n8634), .ZN(n7402) );
  NOR2_X1 U9041 ( .A1(n8634), .A2(n7399), .ZN(n7400) );
  NAND2_X1 U9042 ( .A1(n7402), .A2(n7567), .ZN(n7403) );
  AOI222_X1 U9043 ( .A1(n9493), .A2(n7403), .B1(n8749), .B2(n9489), .C1(n8747), 
        .C2(n9490), .ZN(n9600) );
  INV_X1 U9044 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n7405) );
  INV_X1 U9045 ( .A(n7404), .ZN(n7461) );
  OAI22_X1 U9046 ( .A1(n9510), .A2(n7405), .B1(n7461), .B2(n9499), .ZN(n7408)
         );
  OAI211_X1 U9047 ( .C1(n7366), .C2(n9601), .A(n9496), .B(n7406), .ZN(n9599)
         );
  NOR2_X1 U9048 ( .A1(n9599), .A2(n9085), .ZN(n7407) );
  AOI211_X1 U9049 ( .C1(n9472), .C2(n7464), .A(n7408), .B(n7407), .ZN(n7411)
         );
  XNOR2_X1 U9050 ( .A(n7487), .B(n8634), .ZN(n9603) );
  NAND2_X1 U9051 ( .A1(n9603), .A2(n9482), .ZN(n7410) );
  OAI211_X1 U9052 ( .C1(n9600), .C2(n9485), .A(n7411), .B(n7410), .ZN(P1_U3281) );
  NAND2_X1 U9053 ( .A1(P2_REG2_REG_12__SCAN_IN), .A2(n8008), .ZN(n8021) );
  OAI21_X1 U9054 ( .B1(P2_REG2_REG_12__SCAN_IN), .B2(n8008), .A(n8021), .ZN(
        n7414) );
  AOI21_X1 U9055 ( .B1(n4445), .B2(n7414), .A(n8022), .ZN(n7438) );
  INV_X1 U9056 ( .A(n7415), .ZN(n7417) );
  AOI21_X1 U9057 ( .B1(n7418), .B2(n7417), .A(n7416), .ZN(n8049) );
  INV_X1 U9058 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n7420) );
  INV_X1 U9059 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n7419) );
  MUX2_X1 U9060 ( .A(n7420), .B(n7419), .S(n8057), .Z(n7421) );
  NOR2_X1 U9061 ( .A1(n7421), .A2(n7425), .ZN(n8047) );
  NAND2_X1 U9062 ( .A1(n7421), .A2(n7425), .ZN(n8048) );
  INV_X1 U9063 ( .A(n8048), .ZN(n7422) );
  NOR2_X1 U9064 ( .A1(n8047), .A2(n7422), .ZN(n7424) );
  NAND2_X1 U9065 ( .A1(n8049), .A2(n7424), .ZN(n7423) );
  OAI211_X1 U9066 ( .C1(n8049), .C2(n7424), .A(n9729), .B(n7423), .ZN(n7437)
         );
  AOI22_X1 U9067 ( .A1(P2_REG1_REG_12__SCAN_IN), .A2(n8008), .B1(n7425), .B2(
        n7419), .ZN(n7431) );
  NAND2_X1 U9068 ( .A1(n7427), .A2(n7426), .ZN(n7429) );
  OAI21_X1 U9069 ( .B1(n7431), .B2(n7430), .A(n8009), .ZN(n7435) );
  INV_X1 U9070 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n7432) );
  NOR2_X1 U9071 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7432), .ZN(n7449) );
  AOI21_X1 U9072 ( .B1(n9200), .B2(P2_ADDR_REG_12__SCAN_IN), .A(n7449), .ZN(
        n7433) );
  OAI21_X1 U9073 ( .B1(n8008), .B2(n9721), .A(n7433), .ZN(n7434) );
  AOI21_X1 U9074 ( .B1(n7435), .B2(n9730), .A(n7434), .ZN(n7436) );
  OAI211_X1 U9075 ( .C1(n7438), .C2(n9736), .A(n7437), .B(n7436), .ZN(P2_U3194) );
  OAI222_X1 U9076 ( .A1(n9195), .A2(n7440), .B1(n9193), .B2(n7439), .C1(n5286), 
        .C2(P1_U3086), .ZN(P1_U3327) );
  INV_X1 U9077 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n8007) );
  AND2_X1 U9078 ( .A1(n7690), .A2(n7689), .ZN(n7790) );
  XNOR2_X1 U9079 ( .A(n7441), .B(n7790), .ZN(n7442) );
  AOI222_X1 U9080 ( .A1(n9765), .A2(n7442), .B1(n7995), .B2(n9746), .C1(n7997), 
        .C2(n9744), .ZN(n7479) );
  MUX2_X1 U9081 ( .A(n8007), .B(n7479), .S(n9854), .Z(n7445) );
  XNOR2_X1 U9082 ( .A(n7443), .B(n7790), .ZN(n7482) );
  NOR2_X1 U9083 ( .A1(n9852), .A2(n9796), .ZN(n8223) );
  AOI22_X1 U9084 ( .A1(n7482), .A2(n8223), .B1(n8245), .B2(n7872), .ZN(n7444)
         );
  NAND2_X1 U9085 ( .A1(n7445), .A2(n7444), .ZN(P2_U3473) );
  OAI211_X1 U9086 ( .C1(n7448), .C2(n7447), .A(n7446), .B(n7954), .ZN(n7455)
         );
  AOI21_X1 U9087 ( .B1(n7968), .B2(n7997), .A(n7449), .ZN(n7450) );
  OAI21_X1 U9088 ( .B1(n7451), .B2(n7971), .A(n7450), .ZN(n7452) );
  AOI21_X1 U9089 ( .B1(n7453), .B2(n7987), .A(n7452), .ZN(n7454) );
  OAI211_X1 U9090 ( .C1(n5501), .C2(n7991), .A(n7455), .B(n7454), .ZN(P2_U3164) );
  INV_X1 U9091 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n7456) );
  MUX2_X1 U9092 ( .A(n7456), .B(n7479), .S(n9836), .Z(n7458) );
  INV_X1 U9093 ( .A(n8320), .ZN(n8274) );
  AOI22_X1 U9094 ( .A1(n7482), .A2(n8274), .B1(n8316), .B2(n7872), .ZN(n7457)
         );
  NAND2_X1 U9095 ( .A1(n7458), .A2(n7457), .ZN(P2_U3432) );
  XOR2_X1 U9096 ( .A(n7459), .B(n7460), .Z(n7466) );
  NAND2_X1 U9097 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n9379) );
  OAI21_X1 U9098 ( .B1(n8458), .B2(n7461), .A(n9379), .ZN(n7463) );
  OAI22_X1 U9099 ( .A1(n7559), .A2(n8427), .B1(n8426), .B2(n7472), .ZN(n7462)
         );
  AOI211_X1 U9100 ( .C1(n7464), .C2(n8430), .A(n7463), .B(n7462), .ZN(n7465)
         );
  OAI21_X1 U9101 ( .B1(n7466), .B2(n8462), .A(n7465), .ZN(P1_U3224) );
  XNOR2_X1 U9102 ( .A(n7467), .B(n7531), .ZN(n7469) );
  NOR2_X1 U9103 ( .A1(n7469), .A2(n7468), .ZN(n7530) );
  AOI21_X1 U9104 ( .B1(n7469), .B2(n7468), .A(n7530), .ZN(n7477) );
  NAND2_X1 U9105 ( .A1(P1_REG3_REG_10__SCAN_IN), .A2(P1_U3086), .ZN(n9230) );
  OAI21_X1 U9106 ( .B1(n8458), .B2(n7470), .A(n9230), .ZN(n7474) );
  OAI22_X1 U9107 ( .A1(n7472), .A2(n8427), .B1(n8426), .B2(n7471), .ZN(n7473)
         );
  AOI211_X1 U9108 ( .C1(n7475), .C2(n8460), .A(n7474), .B(n7473), .ZN(n7476)
         );
  OAI21_X1 U9109 ( .B1(n7477), .B2(n8462), .A(n7476), .ZN(P1_U3217) );
  NOR2_X1 U9110 ( .A1(n7478), .A2(n8120), .ZN(n7481) );
  INV_X1 U9111 ( .A(n7479), .ZN(n7480) );
  AOI211_X1 U9112 ( .C1(n9770), .C2(n7868), .A(n7481), .B(n7480), .ZN(n7484)
         );
  AOI22_X1 U9113 ( .A1(n7482), .A2(n9753), .B1(P2_REG2_REG_14__SCAN_IN), .B2(
        n9777), .ZN(n7483) );
  OAI21_X1 U9114 ( .B1(n7484), .B2(n9777), .A(n7483), .ZN(P2_U3219) );
  NAND2_X1 U9115 ( .A1(n7560), .A2(n7559), .ZN(n8692) );
  OR2_X1 U9116 ( .A1(n7560), .A2(n7559), .ZN(n8696) );
  NAND2_X1 U9117 ( .A1(n8692), .A2(n8696), .ZN(n8638) );
  NAND2_X1 U9118 ( .A1(n7567), .A2(n8693), .ZN(n7485) );
  XOR2_X1 U9119 ( .A(n8638), .B(n7485), .Z(n7486) );
  AOI222_X1 U9120 ( .A1(n9493), .A2(n7486), .B1(n8748), .B2(n9489), .C1(n8519), 
        .C2(n9490), .ZN(n9606) );
  XOR2_X1 U9121 ( .A(n8638), .B(n7562), .Z(n9609) );
  NAND2_X1 U9122 ( .A1(n9609), .A2(n9482), .ZN(n7494) );
  INV_X1 U9123 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n7489) );
  INV_X1 U9124 ( .A(n7488), .ZN(n7500) );
  OAI22_X1 U9125 ( .A1(n9510), .A2(n7489), .B1(n7500), .B2(n9499), .ZN(n7492)
         );
  INV_X1 U9126 ( .A(n7406), .ZN(n7490) );
  OAI211_X1 U9127 ( .C1(n7490), .C2(n9607), .A(n9496), .B(n7584), .ZN(n9605)
         );
  NOR2_X1 U9128 ( .A1(n9605), .A2(n9085), .ZN(n7491) );
  AOI211_X1 U9129 ( .C1(n9472), .C2(n7560), .A(n7492), .B(n7491), .ZN(n7493)
         );
  OAI211_X1 U9130 ( .C1(n9485), .C2(n9606), .A(n7494), .B(n7493), .ZN(P1_U3280) );
  INV_X1 U9131 ( .A(n5673), .ZN(n9192) );
  AOI22_X1 U9132 ( .A1(n7495), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_29__SCAN_IN), .B2(n8326), .ZN(n7496) );
  OAI21_X1 U9133 ( .B1(n9192), .B2(n8328), .A(n7496), .ZN(P2_U3266) );
  XOR2_X1 U9134 ( .A(n7497), .B(n7498), .Z(n7503) );
  AOI22_X1 U9135 ( .A1(n8454), .A2(n8519), .B1(n8455), .B2(n8748), .ZN(n7499)
         );
  NAND2_X1 U9136 ( .A1(P1_U3086), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n9394) );
  OAI211_X1 U9137 ( .C1(n8458), .C2(n7500), .A(n7499), .B(n9394), .ZN(n7501)
         );
  AOI21_X1 U9138 ( .B1(n7560), .B2(n8460), .A(n7501), .ZN(n7502) );
  OAI21_X1 U9139 ( .B1(n7503), .B2(n8462), .A(n7502), .ZN(P1_U3234) );
  INV_X1 U9140 ( .A(n7697), .ZN(n7793) );
  XNOR2_X1 U9141 ( .A(n7504), .B(n7793), .ZN(n7519) );
  INV_X1 U9142 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n7510) );
  NOR2_X1 U9143 ( .A1(n4543), .A2(n7505), .ZN(n7509) );
  OAI21_X1 U9144 ( .B1(n7545), .B2(n7506), .A(n7697), .ZN(n7508) );
  OAI22_X1 U9145 ( .A1(n7912), .A2(n9762), .B1(n7994), .B2(n9760), .ZN(n7507)
         );
  AOI21_X1 U9146 ( .B1(n7509), .B2(n7508), .A(n7507), .ZN(n7515) );
  MUX2_X1 U9147 ( .A(n7510), .B(n7515), .S(n9775), .Z(n7512) );
  AOI22_X1 U9148 ( .A1(n7916), .A2(n9751), .B1(n9770), .B2(n7915), .ZN(n7511)
         );
  OAI211_X1 U9149 ( .C1(n7519), .C2(n8208), .A(n7512), .B(n7511), .ZN(P2_U3217) );
  INV_X1 U9150 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8016) );
  MUX2_X1 U9151 ( .A(n8016), .B(n7515), .S(n9854), .Z(n7514) );
  NAND2_X1 U9152 ( .A1(n7916), .A2(n8245), .ZN(n7513) );
  OAI211_X1 U9153 ( .C1(n7519), .C2(n8248), .A(n7514), .B(n7513), .ZN(P2_U3475) );
  INV_X1 U9154 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n7516) );
  MUX2_X1 U9155 ( .A(n7516), .B(n7515), .S(n9836), .Z(n7518) );
  NAND2_X1 U9156 ( .A1(n7916), .A2(n8316), .ZN(n7517) );
  OAI211_X1 U9157 ( .C1(n7519), .C2(n8320), .A(n7518), .B(n7517), .ZN(P2_U3438) );
  INV_X1 U9158 ( .A(n7520), .ZN(n7521) );
  AOI21_X1 U9159 ( .B1(n7523), .B2(n7522), .A(n7521), .ZN(n7529) );
  NAND2_X1 U9160 ( .A1(n7987), .A2(n7524), .ZN(n7526) );
  AOI22_X1 U9161 ( .A1(n7996), .A2(n7968), .B1(P2_REG3_REG_13__SCAN_IN), .B2(
        n9917), .ZN(n7525) );
  OAI211_X1 U9162 ( .C1(n5500), .C2(n7971), .A(n7526), .B(n7525), .ZN(n7527)
         );
  AOI21_X1 U9163 ( .B1(n9286), .B2(n7973), .A(n7527), .ZN(n7528) );
  OAI21_X1 U9164 ( .B1(n7529), .B2(n7977), .A(n7528), .ZN(P2_U3174) );
  AOI21_X1 U9165 ( .B1(n7531), .B2(n7467), .A(n7530), .ZN(n7535) );
  XNOR2_X1 U9166 ( .A(n7533), .B(n7532), .ZN(n7534) );
  XNOR2_X1 U9167 ( .A(n7535), .B(n7534), .ZN(n7542) );
  INV_X1 U9168 ( .A(n7536), .ZN(n7537) );
  NAND2_X1 U9169 ( .A1(P1_U3086), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n9364) );
  OAI21_X1 U9170 ( .B1(n8458), .B2(n7537), .A(n9364), .ZN(n7540) );
  OAI22_X1 U9171 ( .A1(n8750), .A2(n8426), .B1(n8427), .B2(n7538), .ZN(n7539)
         );
  AOI211_X1 U9172 ( .C1(n9590), .C2(n8430), .A(n7540), .B(n7539), .ZN(n7541)
         );
  OAI21_X1 U9173 ( .B1(n7542), .B2(n8462), .A(n7541), .ZN(P1_U3236) );
  XNOR2_X1 U9174 ( .A(n7543), .B(n7692), .ZN(n7558) );
  INV_X1 U9175 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n7549) );
  INV_X1 U9176 ( .A(n7544), .ZN(n7547) );
  INV_X1 U9177 ( .A(n7692), .ZN(n7792) );
  INV_X1 U9178 ( .A(n7545), .ZN(n7546) );
  OAI21_X1 U9179 ( .B1(n7547), .B2(n7792), .A(n7546), .ZN(n7548) );
  AOI222_X1 U9180 ( .A1(n9765), .A2(n7548), .B1(n8202), .B2(n9746), .C1(n7996), 
        .C2(n9744), .ZN(n7555) );
  MUX2_X1 U9181 ( .A(n7549), .B(n7555), .S(n9836), .Z(n7551) );
  NAND2_X1 U9182 ( .A1(n7976), .A2(n8316), .ZN(n7550) );
  OAI211_X1 U9183 ( .C1(n7558), .C2(n8320), .A(n7551), .B(n7550), .ZN(P2_U3435) );
  INV_X1 U9184 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n7552) );
  MUX2_X1 U9185 ( .A(n7552), .B(n7555), .S(n9854), .Z(n7554) );
  NAND2_X1 U9186 ( .A1(n7976), .A2(n8245), .ZN(n7553) );
  OAI211_X1 U9187 ( .C1(n8248), .C2(n7558), .A(n7554), .B(n7553), .ZN(P2_U3474) );
  INV_X1 U9188 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n9693) );
  MUX2_X1 U9189 ( .A(n9693), .B(n7555), .S(n9775), .Z(n7557) );
  AOI22_X1 U9190 ( .A1(n7976), .A2(n9751), .B1(n9770), .B2(n7988), .ZN(n7556)
         );
  OAI211_X1 U9191 ( .C1(n7558), .C2(n8208), .A(n7557), .B(n7556), .ZN(P2_U3218) );
  NAND2_X1 U9192 ( .A1(n9607), .A2(n7559), .ZN(n7561) );
  AOI22_X1 U9193 ( .A1(n7562), .A2(n7561), .B1(n8747), .B2(n7560), .ZN(n7583)
         );
  AOI21_X1 U9194 ( .B1(n7568), .B2(n9614), .A(n7583), .ZN(n7564) );
  NOR2_X2 U9195 ( .A1(n7564), .A2(n7563), .ZN(n7825) );
  NAND2_X1 U9196 ( .A1(n7823), .A2(n8384), .ZN(n8464) );
  NAND2_X1 U9197 ( .A1(n7843), .A2(n8464), .ZN(n8641) );
  XNOR2_X1 U9198 ( .A(n7825), .B(n8641), .ZN(n9298) );
  INV_X1 U9199 ( .A(n9298), .ZN(n7582) );
  AND2_X1 U9200 ( .A1(n8692), .A2(n8693), .ZN(n7566) );
  AOI21_X2 U9201 ( .B1(n7567), .B2(n7566), .A(n7565), .ZN(n7591) );
  XNOR2_X1 U9202 ( .A(n8338), .B(n8519), .ZN(n8524) );
  NAND2_X1 U9203 ( .A1(n7591), .A2(n8524), .ZN(n7571) );
  INV_X1 U9204 ( .A(n7571), .ZN(n7569) );
  AND2_X1 U9205 ( .A1(n8338), .A2(n7568), .ZN(n8526) );
  OAI21_X1 U9206 ( .B1(n7569), .B2(n8526), .A(n8641), .ZN(n7572) );
  NOR2_X1 U9207 ( .A1(n8641), .A2(n8526), .ZN(n7570) );
  NAND2_X1 U9208 ( .A1(n7571), .A2(n7570), .ZN(n7842) );
  NAND3_X1 U9209 ( .A1(n7572), .A2(n7842), .A3(n9493), .ZN(n7574) );
  INV_X1 U9210 ( .A(n9061), .ZN(n8746) );
  AOI22_X1 U9211 ( .A1(n9489), .A2(n8519), .B1(n8746), .B2(n9490), .ZN(n7573)
         );
  NAND2_X1 U9212 ( .A1(n7574), .A2(n7573), .ZN(n9297) );
  INV_X1 U9213 ( .A(n7585), .ZN(n7576) );
  INV_X1 U9214 ( .A(n9079), .ZN(n7575) );
  OAI211_X1 U9215 ( .C1(n9295), .C2(n7576), .A(n7575), .B(n9496), .ZN(n9294)
         );
  INV_X1 U9216 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n9418) );
  INV_X1 U9217 ( .A(n7577), .ZN(n8457) );
  OAI22_X1 U9218 ( .A1(n9510), .A2(n9418), .B1(n8457), .B2(n9499), .ZN(n7578)
         );
  AOI21_X1 U9219 ( .B1(n7823), .B2(n9472), .A(n7578), .ZN(n7579) );
  OAI21_X1 U9220 ( .B1(n9294), .B2(n9085), .A(n7579), .ZN(n7580) );
  AOI21_X1 U9221 ( .B1(n9297), .B2(n9510), .A(n7580), .ZN(n7581) );
  OAI21_X1 U9222 ( .B1(n7582), .B2(n9071), .A(n7581), .ZN(P1_U3278) );
  INV_X1 U9223 ( .A(n8524), .ZN(n8640) );
  XNOR2_X1 U9224 ( .A(n7583), .B(n8640), .ZN(n9616) );
  AOI21_X1 U9225 ( .B1(n7584), .B2(n8338), .A(n9568), .ZN(n7586) );
  NAND2_X1 U9226 ( .A1(n7586), .A2(n7585), .ZN(n9611) );
  INV_X1 U9227 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n7588) );
  INV_X1 U9228 ( .A(n7587), .ZN(n8336) );
  OAI22_X1 U9229 ( .A1(n9510), .A2(n7588), .B1(n8336), .B2(n9499), .ZN(n7589)
         );
  AOI21_X1 U9230 ( .B1(n8338), .B2(n9472), .A(n7589), .ZN(n7590) );
  OAI21_X1 U9231 ( .B1(n9611), .B2(n9085), .A(n7590), .ZN(n7594) );
  OAI21_X1 U9232 ( .B1(n7591), .B2(n8524), .A(n7571), .ZN(n7592) );
  AOI222_X1 U9233 ( .A1(n9493), .A2(n7592), .B1(n9076), .B2(n9490), .C1(n8747), 
        .C2(n9489), .ZN(n9612) );
  NOR2_X1 U9234 ( .A1(n9612), .A2(n9485), .ZN(n7593) );
  AOI211_X1 U9235 ( .C1(n9482), .C2(n9616), .A(n7594), .B(n7593), .ZN(n7595)
         );
  INV_X1 U9236 ( .A(n7595), .ZN(P1_U3279) );
  INV_X1 U9237 ( .A(n7596), .ZN(n8445) );
  INV_X1 U9238 ( .A(n7597), .ZN(n7598) );
  INV_X1 U9239 ( .A(n8914), .ZN(n7603) );
  OAI22_X1 U9240 ( .A1(n7603), .A2(n8458), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n7602), .ZN(n7605) );
  OAI22_X1 U9241 ( .A1(n8867), .A2(n8427), .B1(n8876), .B2(n8426), .ZN(n7604)
         );
  AOI211_X1 U9242 ( .C1(n9109), .C2(n8460), .A(n7605), .B(n7604), .ZN(n7606)
         );
  OAI21_X1 U9243 ( .B1(n7607), .B2(n8462), .A(n7606), .ZN(P1_U3214) );
  MUX2_X1 U9244 ( .A(n8094), .B(n8086), .S(n7747), .Z(n7743) );
  MUX2_X1 U9245 ( .A(n7727), .B(n7728), .S(n7732), .Z(n7608) );
  AND2_X1 U9246 ( .A1(n8090), .A2(n7608), .ZN(n7736) );
  MUX2_X1 U9247 ( .A(n7610), .B(n7609), .S(n7732), .Z(n7698) );
  NAND3_X1 U9248 ( .A1(n7613), .A2(n7612), .A3(n7616), .ZN(n7614) );
  MUX2_X1 U9249 ( .A(n7614), .B(n7613), .S(n7732), .Z(n7621) );
  INV_X1 U9250 ( .A(n7618), .ZN(n7620) );
  NAND3_X1 U9251 ( .A1(n7621), .A2(n7620), .A3(n7619), .ZN(n7629) );
  NAND2_X1 U9252 ( .A1(n8004), .A2(n7622), .ZN(n7631) );
  NAND2_X1 U9253 ( .A1(n9745), .A2(n9769), .ZN(n7623) );
  NAND2_X1 U9254 ( .A1(n7631), .A2(n7623), .ZN(n7626) );
  NAND2_X1 U9255 ( .A1(n7638), .A2(n7624), .ZN(n7625) );
  MUX2_X1 U9256 ( .A(n7626), .B(n7625), .S(n7747), .Z(n7627) );
  INV_X1 U9257 ( .A(n7627), .ZN(n7628) );
  NAND2_X1 U9258 ( .A1(n7629), .A2(n7628), .ZN(n7630) );
  NAND2_X1 U9259 ( .A1(n7630), .A2(n7773), .ZN(n7642) );
  INV_X1 U9260 ( .A(n7631), .ZN(n7633) );
  OAI211_X1 U9261 ( .C1(n7642), .C2(n7633), .A(n7644), .B(n7632), .ZN(n7637)
         );
  INV_X1 U9262 ( .A(n7639), .ZN(n7634) );
  AOI21_X1 U9263 ( .B1(n7635), .B2(n7634), .A(n7643), .ZN(n7636) );
  NAND2_X1 U9264 ( .A1(n7637), .A2(n7636), .ZN(n7647) );
  INV_X1 U9265 ( .A(n7638), .ZN(n7641) );
  OAI211_X1 U9266 ( .C1(n7642), .C2(n7641), .A(n7640), .B(n7639), .ZN(n7645)
         );
  AOI21_X1 U9267 ( .B1(n7645), .B2(n7644), .A(n7643), .ZN(n7646) );
  MUX2_X1 U9268 ( .A(n7647), .B(n7646), .S(n7732), .Z(n7652) );
  NAND3_X1 U9269 ( .A1(n7649), .A2(n7732), .A3(n7648), .ZN(n7651) );
  AND2_X1 U9270 ( .A1(n7654), .A2(n7747), .ZN(n7650) );
  NAND2_X1 U9271 ( .A1(n7657), .A2(n7650), .ZN(n7662) );
  NAND2_X1 U9272 ( .A1(n7651), .A2(n7662), .ZN(n7656) );
  NAND3_X1 U9273 ( .A1(n7652), .A2(n7779), .A3(n7656), .ZN(n7667) );
  NAND2_X1 U9274 ( .A1(n7654), .A2(n7653), .ZN(n7655) );
  NAND2_X1 U9275 ( .A1(n7656), .A2(n7655), .ZN(n7658) );
  NAND3_X1 U9276 ( .A1(n7658), .A2(n7657), .A3(n7671), .ZN(n7659) );
  MUX2_X1 U9277 ( .A(n7660), .B(n7659), .S(n7732), .Z(n7661) );
  INV_X1 U9278 ( .A(n7661), .ZN(n7666) );
  INV_X1 U9279 ( .A(n7662), .ZN(n7664) );
  NAND2_X1 U9280 ( .A1(n7664), .A2(n7663), .ZN(n7665) );
  NAND4_X1 U9281 ( .A1(n7667), .A2(n7782), .A3(n7666), .A4(n7665), .ZN(n7678)
         );
  INV_X1 U9282 ( .A(n7668), .ZN(n7669) );
  NAND2_X1 U9283 ( .A1(n7672), .A2(n7669), .ZN(n7670) );
  AND2_X1 U9284 ( .A1(n7670), .A2(n7673), .ZN(n7676) );
  NAND2_X1 U9285 ( .A1(n7672), .A2(n7671), .ZN(n7674) );
  NAND2_X1 U9286 ( .A1(n7674), .A2(n7673), .ZN(n7675) );
  MUX2_X1 U9287 ( .A(n7676), .B(n7675), .S(n7747), .Z(n7677) );
  NAND2_X1 U9288 ( .A1(n7678), .A2(n7677), .ZN(n7679) );
  NAND2_X1 U9289 ( .A1(n7679), .A2(n7787), .ZN(n7684) );
  NAND2_X1 U9290 ( .A1(n9834), .A2(n5500), .ZN(n7680) );
  MUX2_X1 U9291 ( .A(n7681), .B(n7680), .S(n7747), .Z(n7683) );
  AOI21_X1 U9292 ( .B1(n7684), .B2(n7683), .A(n7682), .ZN(n7688) );
  MUX2_X1 U9293 ( .A(n7686), .B(n7685), .S(n7732), .Z(n7687) );
  OAI21_X1 U9294 ( .B1(n7688), .B2(n7687), .A(n7790), .ZN(n7693) );
  MUX2_X1 U9295 ( .A(n7690), .B(n7689), .S(n7747), .Z(n7691) );
  MUX2_X1 U9296 ( .A(n7695), .B(n7694), .S(n7732), .Z(n7696) );
  NAND2_X1 U9297 ( .A1(n7699), .A2(n7702), .ZN(n7700) );
  NAND2_X1 U9298 ( .A1(n7700), .A2(n7771), .ZN(n7705) );
  NAND3_X1 U9299 ( .A1(n7709), .A2(n7772), .A3(n7703), .ZN(n7704) );
  MUX2_X1 U9300 ( .A(n7705), .B(n7704), .S(n7732), .Z(n7712) );
  NAND3_X1 U9301 ( .A1(n7712), .A2(n7706), .A3(n7713), .ZN(n7707) );
  NAND3_X1 U9302 ( .A1(n7716), .A2(n7710), .A3(n7707), .ZN(n7708) );
  OAI211_X1 U9303 ( .C1(n7712), .C2(n7711), .A(n7710), .B(n7709), .ZN(n7715)
         );
  NAND3_X1 U9304 ( .A1(n7715), .A2(n7714), .A3(n7713), .ZN(n7717) );
  MUX2_X1 U9305 ( .A(n7719), .B(n7718), .S(n7747), .Z(n7720) );
  INV_X1 U9306 ( .A(n7720), .ZN(n7721) );
  MUX2_X1 U9307 ( .A(n7722), .B(n7732), .S(n7723), .Z(n7726) );
  OAI21_X1 U9308 ( .B1(n7723), .B2(n7770), .A(n7769), .ZN(n7724) );
  NAND2_X1 U9309 ( .A1(n7724), .A2(n7732), .ZN(n7725) );
  MUX2_X1 U9310 ( .A(n7730), .B(n7729), .S(n7747), .Z(n7731) );
  NOR2_X1 U9311 ( .A1(n8080), .A2(n7732), .ZN(n7734) );
  NOR2_X1 U9312 ( .A1(n8102), .A2(n7747), .ZN(n7733) );
  MUX2_X1 U9313 ( .A(n7734), .B(n7733), .S(n8257), .Z(n7735) );
  NAND2_X1 U9314 ( .A1(n7855), .A2(n7751), .ZN(n7739) );
  NAND2_X1 U9315 ( .A1(n7752), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n7738) );
  NAND2_X1 U9316 ( .A1(n7739), .A2(n7738), .ZN(n8073) );
  NAND2_X1 U9317 ( .A1(n8073), .A2(n7741), .ZN(n7802) );
  AND2_X1 U9318 ( .A1(n7802), .A2(n7740), .ZN(n7764) );
  OR2_X1 U9319 ( .A1(n8073), .A2(n7741), .ZN(n7803) );
  AND2_X1 U9320 ( .A1(n7803), .A2(n7762), .ZN(n7742) );
  AND2_X1 U9321 ( .A1(n7744), .A2(n7743), .ZN(n7745) );
  NAND2_X1 U9322 ( .A1(n7750), .A2(n7802), .ZN(n7748) );
  NAND2_X1 U9323 ( .A1(n8322), .A2(n7751), .ZN(n7754) );
  NAND2_X1 U9324 ( .A1(n7752), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n7753) );
  INV_X1 U9325 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n7758) );
  NAND2_X1 U9326 ( .A1(n5398), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n7756) );
  NAND2_X1 U9327 ( .A1(n5416), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n7755) );
  OAI211_X1 U9328 ( .C1(n7758), .C2(n7757), .A(n7756), .B(n7755), .ZN(n7759)
         );
  INV_X1 U9329 ( .A(n7759), .ZN(n7760) );
  NOR2_X1 U9330 ( .A1(n9279), .A2(n8069), .ZN(n7801) );
  INV_X1 U9331 ( .A(n9279), .ZN(n8072) );
  INV_X1 U9332 ( .A(n8069), .ZN(n7993) );
  OAI21_X1 U9333 ( .B1(n7993), .B2(n8073), .A(n8072), .ZN(n7763) );
  INV_X1 U9334 ( .A(n7808), .ZN(n7766) );
  NOR2_X1 U9335 ( .A1(n7767), .A2(n7766), .ZN(n7811) );
  INV_X1 U9336 ( .A(n8090), .ZN(n8092) );
  NAND2_X1 U9337 ( .A1(n7770), .A2(n8128), .ZN(n8136) );
  INV_X1 U9338 ( .A(n8179), .ZN(n8177) );
  NAND2_X1 U9339 ( .A1(n7772), .A2(n7771), .ZN(n8190) );
  NAND3_X1 U9340 ( .A1(n5704), .A2(n7774), .A3(n7773), .ZN(n7777) );
  INV_X1 U9341 ( .A(n7775), .ZN(n7776) );
  INV_X1 U9342 ( .A(n9750), .ZN(n9742) );
  NOR4_X1 U9343 ( .A1(n7777), .A2(n9759), .A3(n7776), .A4(n9742), .ZN(n7781)
         );
  NAND4_X1 U9344 ( .A1(n7781), .A2(n7780), .A3(n7779), .A4(n7778), .ZN(n7786)
         );
  INV_X1 U9345 ( .A(n7782), .ZN(n7785) );
  NOR4_X1 U9346 ( .A1(n7786), .A2(n7785), .A3(n7784), .A4(n7783), .ZN(n7789)
         );
  NAND4_X1 U9347 ( .A1(n7790), .A2(n7789), .A3(n7788), .A4(n7787), .ZN(n7791)
         );
  NOR4_X1 U9348 ( .A1(n8190), .A2(n7793), .A3(n7792), .A4(n7791), .ZN(n7794)
         );
  NAND4_X1 U9349 ( .A1(n7795), .A2(n8200), .A3(n8177), .A4(n7794), .ZN(n7796)
         );
  NOR4_X1 U9350 ( .A1(n8136), .A2(n8145), .A3(n7797), .A4(n7796), .ZN(n7798)
         );
  NAND4_X1 U9351 ( .A1(n8101), .A2(n8117), .A3(n8132), .A4(n7798), .ZN(n7799)
         );
  NOR4_X1 U9352 ( .A1(n7800), .A2(n8077), .A3(n8092), .A4(n7799), .ZN(n7805)
         );
  INV_X1 U9353 ( .A(n7801), .ZN(n7804) );
  NAND4_X1 U9354 ( .A1(n7805), .A2(n7804), .A3(n7803), .A4(n7802), .ZN(n7809)
         );
  NOR2_X1 U9355 ( .A1(n7811), .A2(n7810), .ZN(n7812) );
  XNOR2_X1 U9356 ( .A(n7813), .B(n8020), .ZN(n7820) );
  NAND3_X1 U9357 ( .A1(n7815), .A2(n7814), .A3(n8046), .ZN(n7816) );
  OAI211_X1 U9358 ( .C1(n7817), .C2(n7819), .A(n7816), .B(P2_B_REG_SCAN_IN), 
        .ZN(n7818) );
  OAI21_X1 U9359 ( .B1(n7820), .B2(n7819), .A(n7818), .ZN(P2_U3296) );
  OAI222_X1 U9360 ( .A1(n9195), .A2(n7822), .B1(P1_U3086), .B2(n5287), .C1(
        n7821), .C2(n9193), .ZN(P1_U3328) );
  NAND2_X1 U9361 ( .A1(n7823), .A2(n9076), .ZN(n7824) );
  NAND2_X1 U9362 ( .A1(n7825), .A2(n7824), .ZN(n7827) );
  NAND2_X1 U9363 ( .A1(n9295), .A2(n8384), .ZN(n7826) );
  NAND2_X1 U9364 ( .A1(n7829), .A2(n7828), .ZN(n7830) );
  NAND2_X1 U9365 ( .A1(n9068), .A2(n8383), .ZN(n7831) );
  NAND2_X1 U9366 ( .A1(n7832), .A2(n7831), .ZN(n9039) );
  NAND2_X1 U9367 ( .A1(n9017), .A2(n9026), .ZN(n7833) );
  NAND2_X1 U9368 ( .A1(n9140), .A2(n8745), .ZN(n7834) );
  NAND2_X1 U9369 ( .A1(n8988), .A2(n7834), .ZN(n7836) );
  INV_X1 U9370 ( .A(n9140), .ZN(n8991) );
  NAND2_X1 U9371 ( .A1(n8991), .A2(n9010), .ZN(n7835) );
  NAND2_X1 U9372 ( .A1(n8971), .A2(n8980), .ZN(n7837) );
  NOR2_X1 U9373 ( .A1(n8957), .A2(n8964), .ZN(n7839) );
  NAND2_X1 U9374 ( .A1(n8957), .A2(n8964), .ZN(n7838) );
  OAI21_X2 U9375 ( .B1(n8945), .B2(n7839), .A(n7838), .ZN(n8875) );
  OR2_X1 U9376 ( .A1(n9119), .A2(n8950), .ZN(n8599) );
  NAND2_X1 U9377 ( .A1(n9119), .A2(n8950), .ZN(n8860) );
  XNOR2_X1 U9378 ( .A(n8875), .B(n8647), .ZN(n9122) );
  AOI211_X1 U9379 ( .C1(n9119), .C2(n8951), .A(n9568), .B(n4492), .ZN(n9118)
         );
  INV_X1 U9380 ( .A(n8369), .ZN(n7840) );
  AOI22_X1 U9381 ( .A1(n7840), .A2(n9471), .B1(P1_REG2_REG_25__SCAN_IN), .B2(
        n9485), .ZN(n7841) );
  OAI21_X1 U9382 ( .B1(n8873), .B2(n9067), .A(n7841), .ZN(n7853) );
  NAND2_X1 U9383 ( .A1(n7842), .A2(n7843), .ZN(n9074) );
  NAND2_X1 U9384 ( .A1(n8528), .A2(n7843), .ZN(n8518) );
  NAND2_X1 U9385 ( .A1(n8518), .A2(n8465), .ZN(n8699) );
  OR2_X1 U9386 ( .A1(n7829), .A2(n8383), .ZN(n8540) );
  NAND2_X1 U9387 ( .A1(n7829), .A2(n8383), .ZN(n8533) );
  NAND2_X1 U9388 ( .A1(n8540), .A2(n8533), .ZN(n9057) );
  NAND2_X1 U9389 ( .A1(n9054), .A2(n8533), .ZN(n9044) );
  INV_X1 U9390 ( .A(n9034), .ZN(n9059) );
  OR2_X1 U9391 ( .A1(n9154), .A2(n9059), .ZN(n8541) );
  NAND2_X1 U9392 ( .A1(n9154), .A2(n9059), .ZN(n9027) );
  NAND2_X1 U9393 ( .A1(n9044), .A2(n9046), .ZN(n9045) );
  OR2_X1 U9394 ( .A1(n9148), .A2(n9009), .ZN(n8615) );
  NAND2_X1 U9395 ( .A1(n9148), .A2(n9009), .ZN(n8665) );
  NAND2_X1 U9396 ( .A1(n8615), .A2(n8665), .ZN(n9031) );
  INV_X1 U9397 ( .A(n9027), .ZN(n7844) );
  NOR2_X1 U9398 ( .A1(n9031), .A2(n7844), .ZN(n7845) );
  OR2_X1 U9399 ( .A1(n9145), .A2(n9026), .ZN(n8626) );
  AND2_X1 U9400 ( .A1(n8626), .A2(n8615), .ZN(n8537) );
  NAND2_X1 U9401 ( .A1(n9145), .A2(n9026), .ZN(n8996) );
  OR2_X1 U9402 ( .A1(n9140), .A2(n9010), .ZN(n8601) );
  NAND2_X1 U9403 ( .A1(n9140), .A2(n9010), .ZN(n8550) );
  INV_X1 U9404 ( .A(n8550), .ZN(n7846) );
  INV_X1 U9405 ( .A(n8744), .ZN(n9002) );
  OR2_X1 U9406 ( .A1(n9135), .A2(n9002), .ZN(n8554) );
  NAND2_X1 U9407 ( .A1(n9135), .A2(n9002), .ZN(n8556) );
  NAND2_X1 U9408 ( .A1(n8554), .A2(n8556), .ZN(n8977) );
  INV_X1 U9409 ( .A(n8556), .ZN(n7847) );
  NAND2_X1 U9410 ( .A1(n9130), .A2(n8980), .ZN(n8593) );
  NAND2_X1 U9411 ( .A1(n8558), .A2(n8593), .ZN(n8961) );
  NAND2_X1 U9412 ( .A1(n9125), .A2(n8964), .ZN(n8605) );
  NAND2_X1 U9413 ( .A1(n8596), .A2(n8605), .ZN(n8944) );
  NOR3_X1 U9414 ( .A1(n8946), .A2(n4565), .A3(n8944), .ZN(n7849) );
  INV_X1 U9415 ( .A(n8596), .ZN(n7848) );
  NAND2_X1 U9416 ( .A1(n7850), .A2(n8647), .ZN(n8861) );
  OAI21_X1 U9417 ( .B1(n8647), .B2(n7850), .A(n8861), .ZN(n7851) );
  AOI222_X1 U9418 ( .A1(n9493), .A2(n7851), .B1(n8921), .B2(n9490), .C1(n8742), 
        .C2(n9489), .ZN(n9121) );
  NOR2_X1 U9419 ( .A1(n9121), .A2(n9485), .ZN(n7852) );
  AOI211_X1 U9420 ( .C1(n9118), .C2(n9480), .A(n7853), .B(n7852), .ZN(n7854)
         );
  OAI21_X1 U9421 ( .B1(n9122), .B2(n9071), .A(n7854), .ZN(P1_U3268) );
  INV_X1 U9422 ( .A(n7855), .ZN(n8329) );
  INV_X1 U9423 ( .A(n5903), .ZN(n7856) );
  OAI222_X1 U9424 ( .A1(n7858), .A2(n7857), .B1(n9193), .B2(n8329), .C1(
        P1_U3086), .C2(n7856), .ZN(P1_U3325) );
  INV_X1 U9425 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n7860) );
  NAND2_X1 U9426 ( .A1(n7859), .A2(n9770), .ZN(n8070) );
  OAI21_X1 U9427 ( .B1(n9775), .B2(n7860), .A(n8070), .ZN(n7863) );
  NOR2_X1 U9428 ( .A1(n7861), .A2(n8208), .ZN(n7862) );
  AOI211_X1 U9429 ( .C1(n9751), .C2(n5683), .A(n7863), .B(n7862), .ZN(n7864)
         );
  OAI21_X1 U9430 ( .B1(n7865), .B2(n9777), .A(n7864), .ZN(P2_U3204) );
  XOR2_X1 U9431 ( .A(n7867), .B(n7866), .Z(n7874) );
  NAND2_X1 U9432 ( .A1(n7987), .A2(n7868), .ZN(n7870) );
  AOI22_X1 U9433 ( .A1(n7982), .A2(n7997), .B1(P2_REG3_REG_14__SCAN_IN), .B2(
        P2_U3151), .ZN(n7869) );
  OAI211_X1 U9434 ( .C1(n7912), .C2(n7984), .A(n7870), .B(n7869), .ZN(n7871)
         );
  AOI21_X1 U9435 ( .B1(n7872), .B2(n7973), .A(n7871), .ZN(n7873) );
  OAI21_X1 U9436 ( .B1(n7874), .B2(n7977), .A(n7873), .ZN(P2_U3155) );
  AOI21_X1 U9437 ( .B1(n8149), .B2(n7875), .A(n4388), .ZN(n7880) );
  AOI22_X1 U9438 ( .A1(n8161), .A2(n7982), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        n9917), .ZN(n7877) );
  NAND2_X1 U9439 ( .A1(n8141), .A2(n7987), .ZN(n7876) );
  OAI211_X1 U9440 ( .C1(n7903), .C2(n7984), .A(n7877), .B(n7876), .ZN(n7878)
         );
  AOI21_X1 U9441 ( .B1(n8280), .B2(n7973), .A(n7878), .ZN(n7879) );
  OAI21_X1 U9442 ( .B1(n7880), .B2(n7977), .A(n7879), .ZN(P2_U3156) );
  XOR2_X1 U9443 ( .A(n7881), .B(n7882), .Z(n7888) );
  INV_X1 U9444 ( .A(n7893), .ZN(n8181) );
  AOI22_X1 U9445 ( .A1(n8181), .A2(n7968), .B1(P2_REG3_REG_19__SCAN_IN), .B2(
        P2_U3151), .ZN(n7884) );
  NAND2_X1 U9446 ( .A1(n7987), .A2(n8184), .ZN(n7883) );
  OAI211_X1 U9447 ( .C1(n7885), .C2(n7971), .A(n7884), .B(n7883), .ZN(n7886)
         );
  AOI21_X1 U9448 ( .B1(n8304), .B2(n7973), .A(n7886), .ZN(n7887) );
  OAI21_X1 U9449 ( .B1(n7888), .B2(n7977), .A(n7887), .ZN(P2_U3159) );
  XOR2_X1 U9450 ( .A(n7890), .B(n7889), .Z(n7896) );
  AOI22_X1 U9451 ( .A1(n8161), .A2(n7968), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        n9917), .ZN(n7892) );
  NAND2_X1 U9452 ( .A1(n7987), .A2(n8164), .ZN(n7891) );
  OAI211_X1 U9453 ( .C1(n7893), .C2(n7971), .A(n7892), .B(n7891), .ZN(n7894)
         );
  AOI21_X1 U9454 ( .B1(n8292), .B2(n7973), .A(n7894), .ZN(n7895) );
  OAI21_X1 U9455 ( .B1(n7896), .B2(n7977), .A(n7895), .ZN(P2_U3163) );
  INV_X1 U9456 ( .A(n7897), .ZN(n7935) );
  INV_X1 U9457 ( .A(n7898), .ZN(n7900) );
  OAI21_X1 U9458 ( .B1(n7902), .B2(n7901), .A(n7954), .ZN(n7908) );
  OAI22_X1 U9459 ( .A1(n7903), .A2(n7971), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10050), .ZN(n7906) );
  NOR2_X1 U9460 ( .A1(n7904), .A2(n7984), .ZN(n7905) );
  AOI211_X1 U9461 ( .C1(n8115), .C2(n7987), .A(n7906), .B(n7905), .ZN(n7907)
         );
  OAI211_X1 U9462 ( .C1(n8108), .C2(n7991), .A(n7908), .B(n7907), .ZN(P2_U3165) );
  INV_X1 U9463 ( .A(n7909), .ZN(n7922) );
  AOI21_X1 U9464 ( .B1(n7911), .B2(n7910), .A(n7922), .ZN(n7919) );
  NOR2_X1 U9465 ( .A1(n7912), .A2(n7971), .ZN(n7914) );
  OAI22_X1 U9466 ( .A1(n7994), .A2(n7984), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10066), .ZN(n7913) );
  AOI211_X1 U9467 ( .C1(n7915), .C2(n7987), .A(n7914), .B(n7913), .ZN(n7918)
         );
  NAND2_X1 U9468 ( .A1(n7916), .A2(n7973), .ZN(n7917) );
  OAI211_X1 U9469 ( .C1(n7919), .C2(n7977), .A(n7918), .B(n7917), .ZN(P2_U3166) );
  INV_X1 U9470 ( .A(n7920), .ZN(n7921) );
  NOR3_X1 U9471 ( .A1(n7922), .A2(n7921), .A3(n7923), .ZN(n7926) );
  NAND2_X1 U9472 ( .A1(n7924), .A2(n7923), .ZN(n7965) );
  INV_X1 U9473 ( .A(n7965), .ZN(n7925) );
  OAI21_X1 U9474 ( .B1(n7926), .B2(n7925), .A(n7954), .ZN(n7930) );
  AOI22_X1 U9475 ( .A1(n8203), .A2(n7968), .B1(P2_REG3_REG_17__SCAN_IN), .B2(
        P2_U3151), .ZN(n7927) );
  OAI21_X1 U9476 ( .B1(n7985), .B2(n7971), .A(n7927), .ZN(n7928) );
  AOI21_X1 U9477 ( .B1(n8205), .B2(n7987), .A(n7928), .ZN(n7929) );
  OAI211_X1 U9478 ( .C1(n7931), .C2(n7991), .A(n7930), .B(n7929), .ZN(P2_U3168) );
  INV_X1 U9479 ( .A(n7932), .ZN(n7934) );
  NOR3_X1 U9480 ( .A1(n4388), .A2(n7934), .A3(n7933), .ZN(n7936) );
  OAI21_X1 U9481 ( .B1(n7936), .B2(n7935), .A(n7954), .ZN(n7942) );
  INV_X1 U9482 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n7937) );
  OAI22_X1 U9483 ( .A1(n7958), .A2(n7971), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7937), .ZN(n7940) );
  NOR2_X1 U9484 ( .A1(n7938), .A2(n7984), .ZN(n7939) );
  AOI211_X1 U9485 ( .C1(n8127), .C2(n7987), .A(n7940), .B(n7939), .ZN(n7941)
         );
  OAI211_X1 U9486 ( .C1(n8121), .C2(n7991), .A(n7942), .B(n7941), .ZN(P2_U3169) );
  XOR2_X1 U9487 ( .A(n7943), .B(n7944), .Z(n7950) );
  AOI22_X1 U9488 ( .A1(n8171), .A2(n7968), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3151), .ZN(n7946) );
  NAND2_X1 U9489 ( .A1(n7987), .A2(n8174), .ZN(n7945) );
  OAI211_X1 U9490 ( .C1(n7947), .C2(n7971), .A(n7946), .B(n7945), .ZN(n7948)
         );
  AOI21_X1 U9491 ( .B1(n8298), .B2(n7973), .A(n7948), .ZN(n7949) );
  OAI21_X1 U9492 ( .B1(n7950), .B2(n7977), .A(n7949), .ZN(P2_U3173) );
  XNOR2_X1 U9493 ( .A(n7952), .B(n8161), .ZN(n7953) );
  XNOR2_X1 U9494 ( .A(n7951), .B(n7953), .ZN(n7955) );
  NAND2_X1 U9495 ( .A1(n7955), .A2(n7954), .ZN(n7962) );
  INV_X1 U9496 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n7956) );
  OAI22_X1 U9497 ( .A1(n7957), .A2(n7971), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7956), .ZN(n7960) );
  NOR2_X1 U9498 ( .A1(n7958), .A2(n7984), .ZN(n7959) );
  AOI211_X1 U9499 ( .C1(n8152), .C2(n7987), .A(n7960), .B(n7959), .ZN(n7961)
         );
  OAI211_X1 U9500 ( .C1(n7963), .C2(n7991), .A(n7962), .B(n7961), .ZN(P2_U3175) );
  NAND2_X1 U9501 ( .A1(n7965), .A2(n7964), .ZN(n7966) );
  XOR2_X1 U9502 ( .A(n7967), .B(n7966), .Z(n7975) );
  AOI22_X1 U9503 ( .A1(n8193), .A2(n7968), .B1(P2_REG3_REG_18__SCAN_IN), .B2(
        n9917), .ZN(n7970) );
  NAND2_X1 U9504 ( .A1(n7987), .A2(n8196), .ZN(n7969) );
  OAI211_X1 U9505 ( .C1(n7994), .C2(n7971), .A(n7970), .B(n7969), .ZN(n7972)
         );
  AOI21_X1 U9506 ( .B1(n8310), .B2(n7973), .A(n7972), .ZN(n7974) );
  OAI21_X1 U9507 ( .B1(n7975), .B2(n7977), .A(n7974), .ZN(P2_U3178) );
  INV_X1 U9508 ( .A(n7976), .ZN(n7992) );
  AOI21_X1 U9509 ( .B1(n7979), .B2(n7978), .A(n7977), .ZN(n7981) );
  NAND2_X1 U9510 ( .A1(n7981), .A2(n7980), .ZN(n7990) );
  NAND2_X1 U9511 ( .A1(n7996), .A2(n7982), .ZN(n7983) );
  NAND2_X1 U9512 ( .A1(n9917), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n9697) );
  OAI211_X1 U9513 ( .C1(n7985), .C2(n7984), .A(n7983), .B(n9697), .ZN(n7986)
         );
  AOI21_X1 U9514 ( .B1(n7988), .B2(n7987), .A(n7986), .ZN(n7989) );
  OAI211_X1 U9515 ( .C1(n7992), .C2(n7991), .A(n7990), .B(n7989), .ZN(P2_U3181) );
  MUX2_X1 U9516 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n7993), .S(P2_U3893), .Z(
        P2_U3522) );
  MUX2_X1 U9517 ( .A(n8094), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8005), .Z(
        P2_U3519) );
  MUX2_X1 U9518 ( .A(n8102), .B(P2_DATAO_REG_27__SCAN_IN), .S(n8005), .Z(
        P2_U3518) );
  MUX2_X1 U9519 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n8111), .S(P2_U3893), .Z(
        P2_U3517) );
  MUX2_X1 U9520 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8123), .S(P2_U3893), .Z(
        P2_U3516) );
  MUX2_X1 U9521 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n8138), .S(P2_U3893), .Z(
        P2_U3515) );
  MUX2_X1 U9522 ( .A(n8149), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8005), .Z(
        P2_U3514) );
  MUX2_X1 U9523 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8161), .S(P2_U3893), .Z(
        P2_U3513) );
  MUX2_X1 U9524 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8171), .S(P2_U3893), .Z(
        P2_U3512) );
  MUX2_X1 U9525 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8181), .S(P2_U3893), .Z(
        P2_U3511) );
  MUX2_X1 U9526 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8193), .S(P2_U3893), .Z(
        P2_U3510) );
  MUX2_X1 U9527 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n8203), .S(P2_U3893), .Z(
        P2_U3509) );
  INV_X1 U9528 ( .A(n7994), .ZN(n8192) );
  MUX2_X1 U9529 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8192), .S(P2_U3893), .Z(
        P2_U3508) );
  MUX2_X1 U9530 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8202), .S(P2_U3893), .Z(
        P2_U3507) );
  MUX2_X1 U9531 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n7995), .S(P2_U3893), .Z(
        P2_U3506) );
  MUX2_X1 U9532 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n7996), .S(P2_U3893), .Z(
        P2_U3505) );
  MUX2_X1 U9533 ( .A(n7997), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8005), .Z(
        P2_U3504) );
  MUX2_X1 U9534 ( .A(n7998), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8005), .Z(
        P2_U3503) );
  MUX2_X1 U9535 ( .A(n7999), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8005), .Z(
        P2_U3502) );
  MUX2_X1 U9536 ( .A(n8000), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8005), .Z(
        P2_U3501) );
  MUX2_X1 U9537 ( .A(n8001), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8005), .Z(
        P2_U3500) );
  MUX2_X1 U9538 ( .A(n8002), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8005), .Z(
        P2_U3499) );
  MUX2_X1 U9539 ( .A(n5434), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8005), .Z(
        P2_U3497) );
  MUX2_X1 U9540 ( .A(n8003), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8005), .Z(
        P2_U3496) );
  MUX2_X1 U9541 ( .A(n9747), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8005), .Z(
        P2_U3495) );
  MUX2_X1 U9542 ( .A(n8004), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8005), .Z(
        P2_U3494) );
  MUX2_X1 U9543 ( .A(n9745), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8005), .Z(
        P2_U3493) );
  MUX2_X1 U9544 ( .A(n5373), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8005), .Z(
        P2_U3492) );
  MUX2_X1 U9545 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n8006), .S(P2_U3893), .Z(
        P2_U3491) );
  INV_X1 U9546 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8241) );
  AOI22_X1 U9547 ( .A1(P2_REG1_REG_18__SCAN_IN), .A2(n9206), .B1(n9204), .B2(
        n8241), .ZN(n9199) );
  AOI22_X1 U9548 ( .A1(P2_REG1_REG_16__SCAN_IN), .A2(n9701), .B1(n8040), .B2(
        n8016), .ZN(n9705) );
  NAND2_X1 U9549 ( .A1(P2_REG1_REG_14__SCAN_IN), .A2(n9665), .ZN(n8013) );
  AOI22_X1 U9550 ( .A1(P2_REG1_REG_14__SCAN_IN), .A2(n9665), .B1(n8044), .B2(
        n8007), .ZN(n9669) );
  NAND2_X1 U9551 ( .A1(P2_REG1_REG_12__SCAN_IN), .A2(n8008), .ZN(n8010) );
  NAND2_X1 U9552 ( .A1(n9647), .A2(n8011), .ZN(n8012) );
  NAND2_X1 U9553 ( .A1(P2_REG1_REG_13__SCAN_IN), .A2(n9650), .ZN(n9649) );
  NAND2_X1 U9554 ( .A1(n4759), .A2(n8014), .ZN(n8015) );
  NAND2_X1 U9555 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n9686), .ZN(n9685) );
  NAND2_X1 U9556 ( .A1(n8030), .A2(n8017), .ZN(n8018) );
  NAND2_X1 U9557 ( .A1(P2_REG1_REG_17__SCAN_IN), .A2(n9724), .ZN(n9723) );
  NAND2_X1 U9558 ( .A1(n8018), .A2(n9723), .ZN(n9198) );
  NAND2_X1 U9559 ( .A1(n9199), .A2(n9198), .ZN(n9197) );
  OAI21_X1 U9560 ( .B1(n9204), .B2(n8241), .A(n9197), .ZN(n8019) );
  XNOR2_X1 U9561 ( .A(n8064), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n8036) );
  XNOR2_X1 U9562 ( .A(n8019), .B(n8036), .ZN(n8067) );
  XNOR2_X1 U9563 ( .A(n8020), .B(P2_REG2_REG_19__SCAN_IN), .ZN(n8038) );
  NOR2_X1 U9564 ( .A1(n8050), .A2(n8023), .ZN(n8024) );
  XNOR2_X1 U9565 ( .A(n8023), .B(n8050), .ZN(n9658) );
  NOR2_X1 U9566 ( .A1(n9657), .A2(n9658), .ZN(n9656) );
  NAND2_X1 U9567 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n9665), .ZN(n8025) );
  OAI21_X1 U9568 ( .B1(n9665), .B2(P2_REG2_REG_14__SCAN_IN), .A(n8025), .ZN(
        n9676) );
  NAND2_X1 U9569 ( .A1(P2_REG2_REG_16__SCAN_IN), .A2(n9701), .ZN(n8027) );
  OAI21_X1 U9570 ( .B1(n9701), .B2(P2_REG2_REG_16__SCAN_IN), .A(n8027), .ZN(
        n9712) );
  NOR2_X1 U9571 ( .A1(n9713), .A2(n9712), .ZN(n9711) );
  INV_X1 U9572 ( .A(n8027), .ZN(n8028) );
  INV_X1 U9573 ( .A(n8031), .ZN(n8029) );
  NOR2_X1 U9574 ( .A1(n8039), .A2(n8029), .ZN(n8032) );
  INV_X1 U9575 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n9733) );
  INV_X1 U9576 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8195) );
  OR2_X1 U9577 ( .A1(n9204), .A2(n8195), .ZN(n8033) );
  OAI21_X1 U9578 ( .B1(n9206), .B2(P2_REG2_REG_18__SCAN_IN), .A(n8033), .ZN(
        n9212) );
  INV_X1 U9579 ( .A(n9211), .ZN(n8034) );
  NAND2_X1 U9580 ( .A1(n8034), .A2(n8033), .ZN(n8035) );
  INV_X1 U9581 ( .A(n8036), .ZN(n8037) );
  MUX2_X1 U9582 ( .A(n8038), .B(n8037), .S(n8057), .Z(n8063) );
  MUX2_X1 U9583 ( .A(P2_REG2_REG_17__SCAN_IN), .B(P2_REG1_REG_17__SCAN_IN), 
        .S(n8057), .Z(n8056) );
  XNOR2_X1 U9584 ( .A(n8056), .B(n8039), .ZN(n9727) );
  MUX2_X1 U9585 ( .A(P2_REG2_REG_16__SCAN_IN), .B(P2_REG1_REG_16__SCAN_IN), 
        .S(n8046), .Z(n8041) );
  OR2_X1 U9586 ( .A1(n8041), .A2(n9701), .ZN(n8055) );
  XNOR2_X1 U9587 ( .A(n8041), .B(n8040), .ZN(n9708) );
  MUX2_X1 U9588 ( .A(P2_REG2_REG_15__SCAN_IN), .B(P2_REG1_REG_15__SCAN_IN), 
        .S(n8046), .Z(n8043) );
  OR2_X1 U9589 ( .A1(n8043), .A2(n4759), .ZN(n8054) );
  XNOR2_X1 U9590 ( .A(n8043), .B(n8042), .ZN(n9689) );
  MUX2_X1 U9591 ( .A(P2_REG2_REG_14__SCAN_IN), .B(P2_REG1_REG_14__SCAN_IN), 
        .S(n8046), .Z(n8045) );
  OR2_X1 U9592 ( .A1(n8045), .A2(n9665), .ZN(n8053) );
  XNOR2_X1 U9593 ( .A(n8045), .B(n8044), .ZN(n9672) );
  MUX2_X1 U9594 ( .A(P2_REG2_REG_13__SCAN_IN), .B(P2_REG1_REG_13__SCAN_IN), 
        .S(n8046), .Z(n8051) );
  OR2_X1 U9595 ( .A1(n8051), .A2(n9647), .ZN(n8052) );
  AOI21_X1 U9596 ( .B1(n8049), .B2(n8048), .A(n8047), .ZN(n9652) );
  XNOR2_X1 U9597 ( .A(n8051), .B(n8050), .ZN(n9653) );
  NAND2_X1 U9598 ( .A1(n9652), .A2(n9653), .ZN(n9651) );
  NAND2_X1 U9599 ( .A1(n8052), .A2(n9651), .ZN(n9671) );
  NAND2_X1 U9600 ( .A1(n9708), .A2(n9707), .ZN(n9706) );
  MUX2_X1 U9601 ( .A(n8195), .B(n8241), .S(n8057), .Z(n8059) );
  NAND2_X1 U9602 ( .A1(n9203), .A2(n9206), .ZN(n9210) );
  INV_X1 U9603 ( .A(n8058), .ZN(n8061) );
  INV_X1 U9604 ( .A(n8059), .ZN(n8060) );
  NAND2_X1 U9605 ( .A1(n8061), .A2(n8060), .ZN(n9202) );
  NAND2_X1 U9606 ( .A1(n9210), .A2(n9202), .ZN(n8062) );
  OAI21_X1 U9607 ( .B1(n9777), .B2(n9280), .A(n8070), .ZN(n8074) );
  AOI21_X1 U9608 ( .B1(n9777), .B2(P2_REG2_REG_31__SCAN_IN), .A(n8074), .ZN(
        n8071) );
  OAI21_X1 U9609 ( .B1(n8072), .B2(n8076), .A(n8071), .ZN(P2_U3202) );
  INV_X1 U9610 ( .A(n8073), .ZN(n9281) );
  AOI21_X1 U9611 ( .B1(n9777), .B2(P2_REG2_REG_30__SCAN_IN), .A(n8074), .ZN(
        n8075) );
  OAI21_X1 U9612 ( .B1(n9281), .B2(n8076), .A(n8075), .ZN(P2_U3203) );
  XOR2_X1 U9613 ( .A(n8077), .B(n4419), .Z(n8251) );
  INV_X1 U9614 ( .A(n8251), .ZN(n8089) );
  INV_X1 U9615 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n8084) );
  INV_X1 U9616 ( .A(n8077), .ZN(n8078) );
  XNOR2_X1 U9617 ( .A(n8079), .B(n8078), .ZN(n8083) );
  OAI22_X1 U9618 ( .A1(n8081), .A2(n9760), .B1(n8080), .B2(n9762), .ZN(n8082)
         );
  AOI21_X1 U9619 ( .B1(n8083), .B2(n9765), .A(n8082), .ZN(n8249) );
  MUX2_X1 U9620 ( .A(n8084), .B(n8249), .S(n9775), .Z(n8088) );
  AOI22_X1 U9621 ( .A1(n8086), .A2(n9751), .B1(n9770), .B2(n8085), .ZN(n8087)
         );
  OAI211_X1 U9622 ( .C1(n8089), .C2(n8208), .A(n8088), .B(n8087), .ZN(P2_U3205) );
  XNOR2_X1 U9623 ( .A(n8091), .B(n8090), .ZN(n8258) );
  INV_X1 U9624 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n8095) );
  MUX2_X1 U9625 ( .A(n8095), .B(n8255), .S(n9775), .Z(n8098) );
  AOI22_X1 U9626 ( .A1(n8257), .A2(n9751), .B1(n9770), .B2(n8096), .ZN(n8097)
         );
  OAI211_X1 U9627 ( .C1(n8258), .C2(n8208), .A(n8098), .B(n8097), .ZN(P2_U3206) );
  XOR2_X1 U9628 ( .A(n8101), .B(n8099), .Z(n8264) );
  INV_X1 U9629 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n8104) );
  XOR2_X1 U9630 ( .A(n8101), .B(n8100), .Z(n8103) );
  AOI222_X1 U9631 ( .A1(n9765), .A2(n8103), .B1(n8123), .B2(n9744), .C1(n8102), 
        .C2(n9746), .ZN(n8259) );
  MUX2_X1 U9632 ( .A(n8104), .B(n8259), .S(n9775), .Z(n8107) );
  AOI22_X1 U9633 ( .A1(n8261), .A2(n9751), .B1(n9770), .B2(n8105), .ZN(n8106)
         );
  OAI211_X1 U9634 ( .C1(n8264), .C2(n8208), .A(n8107), .B(n8106), .ZN(P2_U3207) );
  NOR2_X1 U9635 ( .A1(n8108), .A2(n8120), .ZN(n8114) );
  OAI21_X1 U9636 ( .B1(n8110), .B2(n5636), .A(n8109), .ZN(n8112) );
  AOI222_X1 U9637 ( .A1(n9765), .A2(n8112), .B1(n8138), .B2(n9744), .C1(n8111), 
        .C2(n9746), .ZN(n8265) );
  INV_X1 U9638 ( .A(n8265), .ZN(n8113) );
  AOI211_X1 U9639 ( .C1(n9770), .C2(n8115), .A(n8114), .B(n8113), .ZN(n8119)
         );
  XOR2_X1 U9640 ( .A(n8117), .B(n8116), .Z(n8268) );
  AOI22_X1 U9641 ( .A1(n8268), .A2(n9753), .B1(P2_REG2_REG_25__SCAN_IN), .B2(
        n9777), .ZN(n8118) );
  OAI21_X1 U9642 ( .B1(n8119), .B2(n9777), .A(n8118), .ZN(P2_U3208) );
  NOR2_X1 U9643 ( .A1(n8121), .A2(n8120), .ZN(n8126) );
  XNOR2_X1 U9644 ( .A(n8122), .B(n8132), .ZN(n8124) );
  AOI222_X1 U9645 ( .A1(n9765), .A2(n8124), .B1(n8149), .B2(n9744), .C1(n8123), 
        .C2(n9746), .ZN(n8271) );
  INV_X1 U9646 ( .A(n8271), .ZN(n8125) );
  AOI211_X1 U9647 ( .C1(n9770), .C2(n8127), .A(n8126), .B(n8125), .ZN(n8134)
         );
  INV_X1 U9648 ( .A(n8128), .ZN(n8129) );
  NOR2_X1 U9649 ( .A1(n8130), .A2(n8129), .ZN(n8131) );
  XOR2_X1 U9650 ( .A(n8132), .B(n8131), .Z(n8275) );
  AOI22_X1 U9651 ( .A1(n8275), .A2(n9753), .B1(P2_REG2_REG_24__SCAN_IN), .B2(
        n9777), .ZN(n8133) );
  OAI21_X1 U9652 ( .B1(n8134), .B2(n9777), .A(n8133), .ZN(P2_U3209) );
  XOR2_X1 U9653 ( .A(n8136), .B(n8135), .Z(n8283) );
  INV_X1 U9654 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n8140) );
  XNOR2_X1 U9655 ( .A(n8137), .B(n8136), .ZN(n8139) );
  AOI222_X1 U9656 ( .A1(n9765), .A2(n8139), .B1(n8138), .B2(n9746), .C1(n8161), 
        .C2(n9744), .ZN(n8278) );
  MUX2_X1 U9657 ( .A(n8140), .B(n8278), .S(n9775), .Z(n8143) );
  AOI22_X1 U9658 ( .A1(n8280), .A2(n9751), .B1(n9770), .B2(n8141), .ZN(n8142)
         );
  OAI211_X1 U9659 ( .C1(n8283), .C2(n8208), .A(n8143), .B(n8142), .ZN(P2_U3210) );
  XNOR2_X1 U9660 ( .A(n8144), .B(n8145), .ZN(n8289) );
  INV_X1 U9661 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n8151) );
  OR3_X1 U9662 ( .A1(n8156), .A2(n8146), .A3(n8145), .ZN(n8147) );
  NAND2_X1 U9663 ( .A1(n8148), .A2(n8147), .ZN(n8150) );
  AOI222_X1 U9664 ( .A1(n9765), .A2(n8150), .B1(n8171), .B2(n9744), .C1(n8149), 
        .C2(n9746), .ZN(n8284) );
  MUX2_X1 U9665 ( .A(n8151), .B(n8284), .S(n9775), .Z(n8154) );
  AOI22_X1 U9666 ( .A1(n8286), .A2(n9751), .B1(n9770), .B2(n8152), .ZN(n8153)
         );
  OAI211_X1 U9667 ( .C1(n8289), .C2(n8208), .A(n8154), .B(n8153), .ZN(P2_U3211) );
  XNOR2_X1 U9668 ( .A(n8155), .B(n8158), .ZN(n8295) );
  INV_X1 U9669 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n8163) );
  INV_X1 U9670 ( .A(n8156), .ZN(n8160) );
  NAND3_X1 U9671 ( .A1(n8168), .A2(n8158), .A3(n8157), .ZN(n8159) );
  NAND2_X1 U9672 ( .A1(n8160), .A2(n8159), .ZN(n8162) );
  AOI222_X1 U9673 ( .A1(n9765), .A2(n8162), .B1(n8161), .B2(n9746), .C1(n8181), 
        .C2(n9744), .ZN(n8290) );
  MUX2_X1 U9674 ( .A(n8163), .B(n8290), .S(n9775), .Z(n8166) );
  AOI22_X1 U9675 ( .A1(n8292), .A2(n9751), .B1(n9770), .B2(n8164), .ZN(n8165)
         );
  OAI211_X1 U9676 ( .C1(n8295), .C2(n8208), .A(n8166), .B(n8165), .ZN(P2_U3212) );
  XNOR2_X1 U9677 ( .A(n8167), .B(n8169), .ZN(n8301) );
  INV_X1 U9678 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n8173) );
  OAI21_X1 U9679 ( .B1(n8170), .B2(n8169), .A(n8168), .ZN(n8172) );
  AOI222_X1 U9680 ( .A1(n9765), .A2(n8172), .B1(n8171), .B2(n9746), .C1(n8193), 
        .C2(n9744), .ZN(n8296) );
  MUX2_X1 U9681 ( .A(n8173), .B(n8296), .S(n9775), .Z(n8176) );
  AOI22_X1 U9682 ( .A1(n8298), .A2(n9751), .B1(n9770), .B2(n8174), .ZN(n8175)
         );
  OAI211_X1 U9683 ( .C1(n8301), .C2(n8208), .A(n8176), .B(n8175), .ZN(P2_U3213) );
  XNOR2_X1 U9684 ( .A(n8178), .B(n8177), .ZN(n8307) );
  INV_X1 U9685 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n8183) );
  XNOR2_X1 U9686 ( .A(n8180), .B(n8179), .ZN(n8182) );
  AOI222_X1 U9687 ( .A1(n9765), .A2(n8182), .B1(n8203), .B2(n9744), .C1(n8181), 
        .C2(n9746), .ZN(n8302) );
  MUX2_X1 U9688 ( .A(n8183), .B(n8302), .S(n9775), .Z(n8186) );
  AOI22_X1 U9689 ( .A1(n8304), .A2(n9751), .B1(n9770), .B2(n8184), .ZN(n8185)
         );
  OAI211_X1 U9690 ( .C1(n8307), .C2(n8208), .A(n8186), .B(n8185), .ZN(P2_U3214) );
  NAND2_X1 U9691 ( .A1(n8188), .A2(n8187), .ZN(n8189) );
  XOR2_X1 U9692 ( .A(n8190), .B(n8189), .Z(n8313) );
  XOR2_X1 U9693 ( .A(n8191), .B(n8190), .Z(n8194) );
  AOI222_X1 U9694 ( .A1(n9765), .A2(n8194), .B1(n8193), .B2(n9746), .C1(n8192), 
        .C2(n9744), .ZN(n8308) );
  MUX2_X1 U9695 ( .A(n8195), .B(n8308), .S(n9775), .Z(n8198) );
  AOI22_X1 U9696 ( .A1(n8310), .A2(n9751), .B1(n9770), .B2(n8196), .ZN(n8197)
         );
  OAI211_X1 U9697 ( .C1(n8313), .C2(n8208), .A(n8198), .B(n8197), .ZN(P2_U3215) );
  XNOR2_X1 U9698 ( .A(n8199), .B(n8200), .ZN(n8321) );
  XOR2_X1 U9699 ( .A(n8201), .B(n8200), .Z(n8204) );
  AOI222_X1 U9700 ( .A1(n9765), .A2(n8204), .B1(n8203), .B2(n9746), .C1(n8202), 
        .C2(n9744), .ZN(n8314) );
  MUX2_X1 U9701 ( .A(n9733), .B(n8314), .S(n9775), .Z(n8207) );
  AOI22_X1 U9702 ( .A1(n8317), .A2(n9751), .B1(n9770), .B2(n8205), .ZN(n8206)
         );
  OAI211_X1 U9703 ( .C1(n8321), .C2(n8208), .A(n8207), .B(n8206), .ZN(P2_U3216) );
  MUX2_X1 U9704 ( .A(n8209), .B(n8249), .S(n9854), .Z(n8211) );
  NAND2_X1 U9705 ( .A1(n8251), .A2(n8223), .ZN(n8210) );
  OAI211_X1 U9706 ( .C1(n4721), .C2(n8212), .A(n8211), .B(n8210), .ZN(P2_U3487) );
  MUX2_X1 U9707 ( .A(n8213), .B(n8255), .S(n9854), .Z(n8215) );
  NAND2_X1 U9708 ( .A1(n8257), .A2(n8245), .ZN(n8214) );
  OAI211_X1 U9709 ( .C1(n8258), .C2(n8248), .A(n8215), .B(n8214), .ZN(P2_U3486) );
  MUX2_X1 U9710 ( .A(n8216), .B(n8259), .S(n9854), .Z(n8218) );
  NAND2_X1 U9711 ( .A1(n8261), .A2(n8245), .ZN(n8217) );
  OAI211_X1 U9712 ( .C1(n8264), .C2(n8248), .A(n8218), .B(n8217), .ZN(P2_U3485) );
  MUX2_X1 U9713 ( .A(n8219), .B(n8265), .S(n9854), .Z(n8221) );
  AOI22_X1 U9714 ( .A1(n8268), .A2(n8223), .B1(n8245), .B2(n8267), .ZN(n8220)
         );
  NAND2_X1 U9715 ( .A1(n8221), .A2(n8220), .ZN(P2_U3484) );
  MUX2_X1 U9716 ( .A(n8222), .B(n8271), .S(n9854), .Z(n8225) );
  AOI22_X1 U9717 ( .A1(n8275), .A2(n8223), .B1(n8245), .B2(n8273), .ZN(n8224)
         );
  NAND2_X1 U9718 ( .A1(n8225), .A2(n8224), .ZN(P2_U3483) );
  MUX2_X1 U9719 ( .A(n8226), .B(n8278), .S(n9854), .Z(n8228) );
  NAND2_X1 U9720 ( .A1(n8280), .A2(n8245), .ZN(n8227) );
  OAI211_X1 U9721 ( .C1(n8283), .C2(n8248), .A(n8228), .B(n8227), .ZN(P2_U3482) );
  MUX2_X1 U9722 ( .A(n8229), .B(n8284), .S(n9854), .Z(n8231) );
  NAND2_X1 U9723 ( .A1(n8286), .A2(n8245), .ZN(n8230) );
  OAI211_X1 U9724 ( .C1(n8289), .C2(n8248), .A(n8231), .B(n8230), .ZN(P2_U3481) );
  INV_X1 U9725 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n8232) );
  MUX2_X1 U9726 ( .A(n8232), .B(n8290), .S(n9854), .Z(n8234) );
  NAND2_X1 U9727 ( .A1(n8292), .A2(n8245), .ZN(n8233) );
  OAI211_X1 U9728 ( .C1(n8248), .C2(n8295), .A(n8234), .B(n8233), .ZN(P2_U3480) );
  INV_X1 U9729 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n8235) );
  MUX2_X1 U9730 ( .A(n8235), .B(n8296), .S(n9854), .Z(n8237) );
  NAND2_X1 U9731 ( .A1(n8298), .A2(n8245), .ZN(n8236) );
  OAI211_X1 U9732 ( .C1(n8248), .C2(n8301), .A(n8237), .B(n8236), .ZN(P2_U3479) );
  INV_X1 U9733 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n8238) );
  MUX2_X1 U9734 ( .A(n8238), .B(n8302), .S(n9854), .Z(n8240) );
  NAND2_X1 U9735 ( .A1(n8304), .A2(n8245), .ZN(n8239) );
  OAI211_X1 U9736 ( .C1(n8248), .C2(n8307), .A(n8240), .B(n8239), .ZN(P2_U3478) );
  MUX2_X1 U9737 ( .A(n8241), .B(n8308), .S(n9854), .Z(n8243) );
  NAND2_X1 U9738 ( .A1(n8310), .A2(n8245), .ZN(n8242) );
  OAI211_X1 U9739 ( .C1(n8313), .C2(n8248), .A(n8243), .B(n8242), .ZN(P2_U3477) );
  INV_X1 U9740 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n8244) );
  MUX2_X1 U9741 ( .A(n8244), .B(n8314), .S(n9854), .Z(n8247) );
  NAND2_X1 U9742 ( .A1(n8317), .A2(n8245), .ZN(n8246) );
  OAI211_X1 U9743 ( .C1(n8321), .C2(n8248), .A(n8247), .B(n8246), .ZN(P2_U3476) );
  INV_X1 U9744 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n8250) );
  MUX2_X1 U9745 ( .A(n8250), .B(n8249), .S(n9836), .Z(n8253) );
  NAND2_X1 U9746 ( .A1(n8251), .A2(n8274), .ZN(n8252) );
  OAI211_X1 U9747 ( .C1(n4721), .C2(n8254), .A(n8253), .B(n8252), .ZN(P2_U3455) );
  INV_X1 U9748 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n8256) );
  INV_X1 U9749 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n8260) );
  MUX2_X1 U9750 ( .A(n8260), .B(n8259), .S(n9836), .Z(n8263) );
  NAND2_X1 U9751 ( .A1(n8261), .A2(n8316), .ZN(n8262) );
  OAI211_X1 U9752 ( .C1(n8264), .C2(n8320), .A(n8263), .B(n8262), .ZN(P2_U3453) );
  INV_X1 U9753 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n8266) );
  MUX2_X1 U9754 ( .A(n8266), .B(n8265), .S(n9836), .Z(n8270) );
  AOI22_X1 U9755 ( .A1(n8268), .A2(n8274), .B1(n8316), .B2(n8267), .ZN(n8269)
         );
  NAND2_X1 U9756 ( .A1(n8270), .A2(n8269), .ZN(P2_U3452) );
  INV_X1 U9757 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n8272) );
  MUX2_X1 U9758 ( .A(n8272), .B(n8271), .S(n9836), .Z(n8277) );
  AOI22_X1 U9759 ( .A1(n8275), .A2(n8274), .B1(n8316), .B2(n8273), .ZN(n8276)
         );
  NAND2_X1 U9760 ( .A1(n8277), .A2(n8276), .ZN(P2_U3451) );
  INV_X1 U9761 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n8279) );
  MUX2_X1 U9762 ( .A(n8279), .B(n8278), .S(n9836), .Z(n8282) );
  NAND2_X1 U9763 ( .A1(n8280), .A2(n8316), .ZN(n8281) );
  OAI211_X1 U9764 ( .C1(n8283), .C2(n8320), .A(n8282), .B(n8281), .ZN(P2_U3450) );
  INV_X1 U9765 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n8285) );
  MUX2_X1 U9766 ( .A(n8285), .B(n8284), .S(n9836), .Z(n8288) );
  NAND2_X1 U9767 ( .A1(n8286), .A2(n8316), .ZN(n8287) );
  OAI211_X1 U9768 ( .C1(n8289), .C2(n8320), .A(n8288), .B(n8287), .ZN(P2_U3449) );
  INV_X1 U9769 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n8291) );
  MUX2_X1 U9770 ( .A(n8291), .B(n8290), .S(n9836), .Z(n8294) );
  NAND2_X1 U9771 ( .A1(n8292), .A2(n8316), .ZN(n8293) );
  OAI211_X1 U9772 ( .C1(n8295), .C2(n8320), .A(n8294), .B(n8293), .ZN(P2_U3448) );
  INV_X1 U9773 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n8297) );
  MUX2_X1 U9774 ( .A(n8297), .B(n8296), .S(n9836), .Z(n8300) );
  NAND2_X1 U9775 ( .A1(n8298), .A2(n8316), .ZN(n8299) );
  OAI211_X1 U9776 ( .C1(n8301), .C2(n8320), .A(n8300), .B(n8299), .ZN(P2_U3447) );
  INV_X1 U9777 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n8303) );
  MUX2_X1 U9778 ( .A(n8303), .B(n8302), .S(n9836), .Z(n8306) );
  NAND2_X1 U9779 ( .A1(n8304), .A2(n8316), .ZN(n8305) );
  OAI211_X1 U9780 ( .C1(n8307), .C2(n8320), .A(n8306), .B(n8305), .ZN(P2_U3446) );
  INV_X1 U9781 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n8309) );
  MUX2_X1 U9782 ( .A(n8309), .B(n8308), .S(n9836), .Z(n8312) );
  NAND2_X1 U9783 ( .A1(n8310), .A2(n8316), .ZN(n8311) );
  OAI211_X1 U9784 ( .C1(n8313), .C2(n8320), .A(n8312), .B(n8311), .ZN(P2_U3444) );
  INV_X1 U9785 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n8315) );
  MUX2_X1 U9786 ( .A(n8315), .B(n8314), .S(n9836), .Z(n8319) );
  NAND2_X1 U9787 ( .A1(n8317), .A2(n8316), .ZN(n8318) );
  OAI211_X1 U9788 ( .C1(n8321), .C2(n8320), .A(n8319), .B(n8318), .ZN(P2_U3441) );
  INV_X1 U9789 ( .A(n8322), .ZN(n9191) );
  NOR4_X1 U9790 ( .A1(n8323), .A2(P2_IR_REG_30__SCAN_IN), .A3(n9917), .A4(
        n5330), .ZN(n8324) );
  AOI21_X1 U9791 ( .B1(n8326), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n8324), .ZN(
        n8325) );
  OAI21_X1 U9792 ( .B1(n9191), .B2(n8328), .A(n8325), .ZN(P2_U3264) );
  AOI22_X1 U9793 ( .A1(n5334), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n8326), .ZN(n8327) );
  OAI21_X1 U9794 ( .B1(n8329), .B2(n8328), .A(n8327), .ZN(P2_U3265) );
  MUX2_X1 U9795 ( .A(n8330), .B(P2_IR_REG_0__SCAN_IN), .S(P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  INV_X1 U9796 ( .A(n8332), .ZN(n8333) );
  AOI21_X1 U9797 ( .B1(n8331), .B2(n8334), .A(n8333), .ZN(n8340) );
  AOI22_X1 U9798 ( .A1(n8455), .A2(n8747), .B1(n8454), .B2(n9076), .ZN(n8335)
         );
  NAND2_X1 U9799 ( .A1(P1_U3086), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n9410) );
  OAI211_X1 U9800 ( .C1(n8458), .C2(n8336), .A(n8335), .B(n9410), .ZN(n8337)
         );
  AOI21_X1 U9801 ( .B1(n8338), .B2(n8460), .A(n8337), .ZN(n8339) );
  OAI21_X1 U9802 ( .B1(n8340), .B2(n8462), .A(n8339), .ZN(P1_U3215) );
  INV_X1 U9803 ( .A(n8400), .ZN(n8343) );
  NOR3_X1 U9804 ( .A1(n8423), .A2(n8418), .A3(n8341), .ZN(n8342) );
  OAI21_X1 U9805 ( .B1(n8343), .B2(n8342), .A(n8444), .ZN(n8347) );
  NOR2_X1 U9806 ( .A1(n8458), .A2(n8967), .ZN(n8345) );
  OAI22_X1 U9807 ( .A1(n8964), .A2(n8427), .B1(n9002), .B2(n8426), .ZN(n8344)
         );
  AOI211_X1 U9808 ( .C1(P1_REG3_REG_23__SCAN_IN), .C2(P1_U3086), .A(n8345), 
        .B(n8344), .ZN(n8346) );
  OAI211_X1 U9809 ( .C1(n8971), .C2(n8407), .A(n8347), .B(n8346), .ZN(P1_U3216) );
  INV_X1 U9810 ( .A(n8349), .ZN(n8350) );
  XOR2_X1 U9811 ( .A(n8348), .B(n8349), .Z(n8435) );
  NOR2_X1 U9812 ( .A1(n8435), .A2(n8434), .ZN(n8433) );
  AOI21_X1 U9813 ( .B1(n8350), .B2(n8348), .A(n8433), .ZN(n8354) );
  XNOR2_X1 U9814 ( .A(n8352), .B(n8351), .ZN(n8353) );
  XNOR2_X1 U9815 ( .A(n8354), .B(n8353), .ZN(n8355) );
  NAND2_X1 U9816 ( .A1(n8355), .A2(n8444), .ZN(n8358) );
  AND2_X1 U9817 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n8850) );
  OAI22_X1 U9818 ( .A1(n9059), .A2(n8426), .B1(n8427), .B2(n9026), .ZN(n8356)
         );
  AOI211_X1 U9819 ( .C1(n8446), .C2(n9023), .A(n8850), .B(n8356), .ZN(n8357)
         );
  OAI211_X1 U9820 ( .C1(n9025), .C2(n8407), .A(n8358), .B(n8357), .ZN(P1_U3219) );
  XOR2_X1 U9821 ( .A(n8359), .B(n8360), .Z(n8365) );
  OAI22_X1 U9822 ( .A1(n8458), .A2(n8992), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8361), .ZN(n8363) );
  OAI22_X1 U9823 ( .A1(n9026), .A2(n8426), .B1(n8427), .B2(n9002), .ZN(n8362)
         );
  AOI211_X1 U9824 ( .C1(n9140), .C2(n8460), .A(n8363), .B(n8362), .ZN(n8364)
         );
  OAI21_X1 U9825 ( .B1(n8365), .B2(n8462), .A(n8364), .ZN(P1_U3223) );
  AOI21_X1 U9826 ( .B1(n4384), .B2(n8367), .A(n8366), .ZN(n8373) );
  OAI22_X1 U9827 ( .A1(n8369), .A2(n8458), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8368), .ZN(n8371) );
  OAI22_X1 U9828 ( .A1(n8876), .A2(n8427), .B1(n8964), .B2(n8426), .ZN(n8370)
         );
  AOI211_X1 U9829 ( .C1(n9119), .C2(n8460), .A(n8371), .B(n8370), .ZN(n8372)
         );
  OAI21_X1 U9830 ( .B1(n8373), .B2(n8462), .A(n8372), .ZN(P1_U3225) );
  INV_X1 U9831 ( .A(n8375), .ZN(n8376) );
  XOR2_X1 U9832 ( .A(n8374), .B(n8375), .Z(n8453) );
  NOR2_X1 U9833 ( .A1(n8453), .A2(n8452), .ZN(n8451) );
  AOI21_X1 U9834 ( .B1(n8376), .B2(n8374), .A(n8451), .ZN(n8380) );
  XNOR2_X1 U9835 ( .A(n8378), .B(n8377), .ZN(n8379) );
  XNOR2_X1 U9836 ( .A(n8380), .B(n8379), .ZN(n8381) );
  NAND2_X1 U9837 ( .A1(n8381), .A2(n8444), .ZN(n8387) );
  NOR2_X1 U9838 ( .A1(n8382), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9430) );
  OAI22_X1 U9839 ( .A1(n8384), .A2(n8426), .B1(n8427), .B2(n8383), .ZN(n8385)
         );
  AOI211_X1 U9840 ( .C1(n8446), .C2(n9080), .A(n9430), .B(n8385), .ZN(n8386)
         );
  OAI211_X1 U9841 ( .C1(n9164), .C2(n8407), .A(n8387), .B(n8386), .ZN(P1_U3226) );
  INV_X1 U9842 ( .A(n8388), .ZN(n8390) );
  NOR2_X1 U9843 ( .A1(n8390), .A2(n8389), .ZN(n8391) );
  XNOR2_X1 U9844 ( .A(n8392), .B(n8391), .ZN(n8397) );
  INV_X1 U9845 ( .A(n9064), .ZN(n8394) );
  AOI22_X1 U9846 ( .A1(n8454), .A2(n9034), .B1(n8455), .B2(n8746), .ZN(n8393)
         );
  NAND2_X1 U9847 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9448) );
  OAI211_X1 U9848 ( .C1(n8458), .C2(n8394), .A(n8393), .B(n9448), .ZN(n8395)
         );
  AOI21_X1 U9849 ( .B1(n7829), .B2(n8460), .A(n8395), .ZN(n8396) );
  OAI21_X1 U9850 ( .B1(n8397), .B2(n8462), .A(n8396), .ZN(P1_U3228) );
  AND3_X1 U9851 ( .A1(n8400), .A2(n8399), .A3(n8398), .ZN(n8401) );
  OAI21_X1 U9852 ( .B1(n8402), .B2(n8401), .A(n8444), .ZN(n8406) );
  NOR2_X1 U9853 ( .A1(n8458), .A2(n8953), .ZN(n8404) );
  OAI22_X1 U9854 ( .A1(n8950), .A2(n8427), .B1(n8980), .B2(n8426), .ZN(n8403)
         );
  AOI211_X1 U9855 ( .C1(P1_REG3_REG_24__SCAN_IN), .C2(P1_U3086), .A(n8404), 
        .B(n8403), .ZN(n8405) );
  OAI211_X1 U9856 ( .C1(n8957), .C2(n8407), .A(n8406), .B(n8405), .ZN(P1_U3229) );
  XNOR2_X1 U9857 ( .A(n8409), .B(n8408), .ZN(n8410) );
  XNOR2_X1 U9858 ( .A(n8411), .B(n8410), .ZN(n8417) );
  INV_X1 U9859 ( .A(n9014), .ZN(n8413) );
  OAI22_X1 U9860 ( .A1(n8458), .A2(n8413), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8412), .ZN(n8415) );
  OAI22_X1 U9861 ( .A1(n9009), .A2(n8426), .B1(n8427), .B2(n9010), .ZN(n8414)
         );
  AOI211_X1 U9862 ( .C1(n9145), .C2(n8430), .A(n8415), .B(n8414), .ZN(n8416)
         );
  OAI21_X1 U9863 ( .B1(n8417), .B2(n8462), .A(n8416), .ZN(P1_U3233) );
  INV_X1 U9864 ( .A(n8418), .ZN(n8422) );
  OR2_X1 U9865 ( .A1(n8419), .A2(n8418), .ZN(n8420) );
  AOI22_X1 U9866 ( .A1(n8423), .A2(n8422), .B1(n8421), .B2(n8420), .ZN(n8432)
         );
  INV_X1 U9867 ( .A(n8982), .ZN(n8425) );
  OAI22_X1 U9868 ( .A1(n8458), .A2(n8425), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8424), .ZN(n8429) );
  OAI22_X1 U9869 ( .A1(n8980), .A2(n8427), .B1(n8426), .B2(n9010), .ZN(n8428)
         );
  AOI211_X1 U9870 ( .C1(n9135), .C2(n8430), .A(n8429), .B(n8428), .ZN(n8431)
         );
  OAI21_X1 U9871 ( .B1(n8432), .B2(n8462), .A(n8431), .ZN(P1_U3235) );
  AOI21_X1 U9872 ( .B1(n8435), .B2(n8434), .A(n8433), .ZN(n8440) );
  INV_X1 U9873 ( .A(n9041), .ZN(n8437) );
  AOI22_X1 U9874 ( .A1(n8455), .A2(n7828), .B1(n8454), .B2(n9047), .ZN(n8436)
         );
  NAND2_X1 U9875 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9464) );
  OAI211_X1 U9876 ( .C1(n8458), .C2(n8437), .A(n8436), .B(n9464), .ZN(n8438)
         );
  AOI21_X1 U9877 ( .B1(n9154), .B2(n8460), .A(n8438), .ZN(n8439) );
  OAI21_X1 U9878 ( .B1(n8440), .B2(n8462), .A(n8439), .ZN(P1_U3238) );
  OAI21_X1 U9879 ( .B1(n8366), .B2(n8442), .A(n8441), .ZN(n8443) );
  NAND3_X1 U9880 ( .A1(n8445), .A2(n8444), .A3(n8443), .ZN(n8450) );
  AOI22_X1 U9881 ( .A1(n8932), .A2(n8446), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3086), .ZN(n8449) );
  AOI22_X1 U9882 ( .A1(n8939), .A2(n8454), .B1(n8455), .B2(n8938), .ZN(n8448)
         );
  NAND2_X1 U9883 ( .A1(n9114), .A2(n8460), .ZN(n8447) );
  NAND4_X1 U9884 ( .A1(n8450), .A2(n8449), .A3(n8448), .A4(n8447), .ZN(
        P1_U3240) );
  AOI21_X1 U9885 ( .B1(n8453), .B2(n8452), .A(n8451), .ZN(n8463) );
  AOI22_X1 U9886 ( .A1(n8455), .A2(n8519), .B1(n8454), .B2(n8746), .ZN(n8456)
         );
  NAND2_X1 U9887 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9423) );
  OAI211_X1 U9888 ( .C1(n8458), .C2(n8457), .A(n8456), .B(n9423), .ZN(n8459)
         );
  AOI21_X1 U9889 ( .B1(n7823), .B2(n8460), .A(n8459), .ZN(n8461) );
  OAI21_X1 U9890 ( .B1(n8463), .B2(n8462), .A(n8461), .ZN(P1_U3241) );
  NAND2_X1 U9891 ( .A1(n8587), .A2(n8619), .ZN(n8717) );
  AOI22_X1 U9892 ( .A1(n8527), .A2(n8528), .B1(n8734), .B2(n9295), .ZN(n8532)
         );
  AOI21_X1 U9893 ( .B1(n8465), .B2(n9076), .A(n8514), .ZN(n8531) );
  INV_X1 U9894 ( .A(n8477), .ZN(n8467) );
  OAI21_X1 U9895 ( .B1(n7043), .B2(n8467), .A(n8466), .ZN(n8470) );
  NAND2_X1 U9896 ( .A1(n8466), .A2(n8468), .ZN(n8675) );
  AOI21_X1 U9897 ( .B1(n4367), .B2(n8672), .A(n8675), .ZN(n8469) );
  NAND2_X1 U9898 ( .A1(n8480), .A2(n8478), .ZN(n8472) );
  AND2_X1 U9899 ( .A1(n8678), .A2(n8471), .ZN(n8479) );
  NAND2_X1 U9900 ( .A1(n8472), .A2(n8479), .ZN(n8473) );
  NAND2_X1 U9901 ( .A1(n8473), .A2(n7163), .ZN(n8476) );
  NAND2_X1 U9902 ( .A1(n8476), .A2(n4906), .ZN(n8500) );
  NAND2_X1 U9903 ( .A1(n8478), .A2(n8477), .ZN(n8679) );
  OAI21_X1 U9904 ( .B1(n8480), .B2(n8679), .A(n8479), .ZN(n8498) );
  AND4_X1 U9905 ( .A1(n7163), .A2(n8482), .A3(n8481), .A4(n8514), .ZN(n8497)
         );
  NAND2_X1 U9906 ( .A1(n8483), .A2(n8734), .ZN(n8485) );
  OAI21_X1 U9907 ( .B1(n8485), .B2(n8752), .A(n8491), .ZN(n8489) );
  OR2_X1 U9908 ( .A1(n8483), .A2(n8734), .ZN(n8492) );
  OAI21_X1 U9909 ( .B1(n8492), .B2(n8490), .A(n9561), .ZN(n8488) );
  NAND2_X1 U9910 ( .A1(n8490), .A2(n8734), .ZN(n8484) );
  OAI21_X1 U9911 ( .B1(n8485), .B2(n9561), .A(n8484), .ZN(n8487) );
  AOI22_X1 U9912 ( .A1(n8489), .A2(n8488), .B1(n8487), .B2(n8486), .ZN(n8495)
         );
  OAI22_X1 U9913 ( .A1(n8492), .A2(n8491), .B1(n8734), .B2(n8490), .ZN(n8493)
         );
  NAND2_X1 U9914 ( .A1(n8493), .A2(n9567), .ZN(n8494) );
  NAND4_X1 U9915 ( .A1(n8495), .A2(n8506), .A3(n8501), .A4(n8494), .ZN(n8496)
         );
  AOI21_X1 U9916 ( .B1(n8498), .B2(n8497), .A(n8496), .ZN(n8499) );
  NAND2_X1 U9917 ( .A1(n8500), .A2(n8499), .ZN(n8507) );
  NAND2_X1 U9918 ( .A1(n8507), .A2(n8501), .ZN(n8502) );
  NAND2_X1 U9919 ( .A1(n8502), .A2(n8508), .ZN(n8504) );
  NAND2_X1 U9920 ( .A1(n8505), .A2(n8734), .ZN(n8517) );
  NAND2_X1 U9921 ( .A1(n8507), .A2(n8506), .ZN(n8510) );
  NAND2_X1 U9922 ( .A1(n8509), .A2(n8508), .ZN(n8686) );
  AOI21_X1 U9923 ( .B1(n8510), .B2(n8684), .A(n8686), .ZN(n8513) );
  NAND2_X1 U9924 ( .A1(n8512), .A2(n8511), .ZN(n8689) );
  OAI21_X1 U9925 ( .B1(n8513), .B2(n8689), .A(n8693), .ZN(n8515) );
  NAND2_X1 U9926 ( .A1(n8517), .A2(n8516), .ZN(n8523) );
  NAND2_X1 U9927 ( .A1(n8524), .A2(n8692), .ZN(n8522) );
  INV_X1 U9928 ( .A(n8518), .ZN(n8521) );
  AND2_X1 U9929 ( .A1(n9614), .A2(n8519), .ZN(n8695) );
  AOI21_X1 U9930 ( .B1(n8524), .B2(n7565), .A(n8695), .ZN(n8520) );
  OAI211_X1 U9931 ( .C1(n8523), .C2(n8522), .A(n8521), .B(n8520), .ZN(n8530)
         );
  NAND2_X1 U9932 ( .A1(n8523), .A2(n8692), .ZN(n8525) );
  OAI21_X1 U9933 ( .B1(n8701), .B2(n8696), .A(n8528), .ZN(n8529) );
  INV_X1 U9934 ( .A(n9057), .ZN(n9052) );
  AND2_X1 U9935 ( .A1(n9027), .A2(n8533), .ZN(n8705) );
  NAND2_X1 U9936 ( .A1(n8615), .A2(n8541), .ZN(n8703) );
  AOI21_X1 U9937 ( .B1(n8543), .B2(n8705), .A(n8703), .ZN(n8539) );
  NAND2_X1 U9938 ( .A1(n8996), .A2(n9025), .ZN(n8534) );
  NAND2_X1 U9939 ( .A1(n8534), .A2(n8514), .ZN(n8536) );
  AND2_X1 U9940 ( .A1(n9047), .A2(n8514), .ZN(n8535) );
  AOI22_X1 U9941 ( .A1(n8537), .A2(n8536), .B1(n8535), .B2(n8996), .ZN(n8538)
         );
  AND2_X1 U9942 ( .A1(n8541), .A2(n8540), .ZN(n8700) );
  NAND2_X1 U9943 ( .A1(n8665), .A2(n9027), .ZN(n8542) );
  AOI21_X1 U9944 ( .B1(n8543), .B2(n8700), .A(n8542), .ZN(n8544) );
  NAND2_X1 U9945 ( .A1(n8544), .A2(n8734), .ZN(n8545) );
  NAND2_X1 U9946 ( .A1(n8546), .A2(n8545), .ZN(n8549) );
  NAND2_X1 U9947 ( .A1(n8601), .A2(n8626), .ZN(n8611) );
  NAND2_X1 U9948 ( .A1(n8550), .A2(n8996), .ZN(n8602) );
  MUX2_X1 U9949 ( .A(n8611), .B(n8602), .S(n8734), .Z(n8547) );
  INV_X1 U9950 ( .A(n8547), .ZN(n8548) );
  NAND2_X1 U9951 ( .A1(n8549), .A2(n8548), .ZN(n8552) );
  MUX2_X1 U9952 ( .A(n8550), .B(n8601), .S(n8734), .Z(n8551) );
  NAND2_X1 U9953 ( .A1(n8552), .A2(n8551), .ZN(n8553) );
  INV_X1 U9954 ( .A(n8977), .ZN(n8974) );
  NAND2_X1 U9955 ( .A1(n8558), .A2(n8554), .ZN(n8594) );
  NAND2_X1 U9956 ( .A1(n8594), .A2(n8734), .ZN(n8555) );
  NAND2_X1 U9957 ( .A1(n8593), .A2(n8556), .ZN(n8600) );
  NAND2_X1 U9958 ( .A1(n8600), .A2(n8514), .ZN(n8557) );
  NOR2_X1 U9959 ( .A1(n8558), .A2(n8734), .ZN(n8559) );
  NOR2_X1 U9960 ( .A1(n8944), .A2(n8559), .ZN(n8560) );
  NAND2_X1 U9961 ( .A1(n8561), .A2(n8560), .ZN(n8563) );
  MUX2_X1 U9962 ( .A(n8605), .B(n8596), .S(n8734), .Z(n8562) );
  NAND2_X1 U9963 ( .A1(n8563), .A2(n8562), .ZN(n8568) );
  NAND2_X1 U9964 ( .A1(n8568), .A2(n8599), .ZN(n8565) );
  NAND2_X1 U9965 ( .A1(n9114), .A2(n8876), .ZN(n8862) );
  AND2_X1 U9966 ( .A1(n8862), .A2(n8860), .ZN(n8566) );
  INV_X1 U9967 ( .A(n8625), .ZN(n8564) );
  AOI21_X1 U9968 ( .B1(n8565), .B2(n8566), .A(n8564), .ZN(n8570) );
  INV_X1 U9969 ( .A(n8599), .ZN(n8567) );
  NAND2_X1 U9970 ( .A1(n9103), .A2(n8867), .ZN(n8864) );
  NAND2_X1 U9971 ( .A1(n9109), .A2(n8897), .ZN(n8863) );
  NAND2_X1 U9972 ( .A1(n8864), .A2(n8863), .ZN(n8610) );
  INV_X1 U9973 ( .A(n8624), .ZN(n8573) );
  OAI21_X1 U9974 ( .B1(n8610), .B2(n8706), .A(n8624), .ZN(n8571) );
  NAND2_X1 U9975 ( .A1(n8571), .A2(n8734), .ZN(n8572) );
  NAND2_X1 U9976 ( .A1(n8890), .A2(n8898), .ZN(n8618) );
  MUX2_X1 U9977 ( .A(n8618), .B(n8591), .S(n8734), .Z(n8574) );
  INV_X1 U9978 ( .A(n8574), .ZN(n8575) );
  NAND2_X1 U9979 ( .A1(n8856), .A2(n8514), .ZN(n8577) );
  OAI21_X1 U9980 ( .B1(n8582), .B2(n8856), .A(n8577), .ZN(n8586) );
  NAND2_X1 U9981 ( .A1(n8578), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n8581) );
  NAND2_X1 U9982 ( .A1(n5959), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n8580) );
  NAND2_X1 U9983 ( .A1(n5958), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n8579) );
  AND3_X1 U9984 ( .A1(n8581), .A2(n8580), .A3(n8579), .ZN(n8869) );
  AOI21_X1 U9985 ( .B1(n8587), .B2(n8869), .A(n8619), .ZN(n8585) );
  MUX2_X1 U9986 ( .A(n8514), .B(n8582), .S(n8856), .Z(n8583) );
  INV_X1 U9987 ( .A(n8869), .ZN(n8741) );
  NAND3_X1 U9988 ( .A1(n8583), .A2(n8741), .A3(n8587), .ZN(n8584) );
  OAI211_X1 U9989 ( .C1(n8586), .C2(n8585), .A(n8584), .B(n8717), .ZN(n8739)
         );
  OAI21_X1 U9990 ( .B1(n8717), .B2(n8514), .A(n8739), .ZN(n8729) );
  OR2_X1 U9991 ( .A1(n8587), .A2(n8619), .ZN(n8719) );
  NOR2_X1 U9992 ( .A1(n8719), .A2(n4453), .ZN(n8590) );
  NOR4_X1 U9993 ( .A1(n8590), .A2(n8589), .A3(n8732), .A4(n8588), .ZN(n8728)
         );
  NAND2_X1 U9994 ( .A1(n8591), .A2(n8624), .ZN(n8663) );
  INV_X1 U9995 ( .A(n8862), .ZN(n8592) );
  AND2_X1 U9996 ( .A1(n8706), .A2(n8592), .ZN(n8609) );
  NAND2_X1 U9997 ( .A1(n8594), .A2(n8593), .ZN(n8595) );
  NAND2_X1 U9998 ( .A1(n8596), .A2(n8595), .ZN(n8597) );
  NAND2_X1 U9999 ( .A1(n8597), .A2(n8605), .ZN(n8598) );
  NAND2_X1 U10000 ( .A1(n8599), .A2(n8598), .ZN(n8612) );
  INV_X1 U10001 ( .A(n8600), .ZN(n8604) );
  NAND2_X1 U10002 ( .A1(n8602), .A2(n8601), .ZN(n8603) );
  AND3_X1 U10003 ( .A1(n8605), .A2(n8604), .A3(n8603), .ZN(n8606) );
  OAI21_X1 U10004 ( .B1(n8612), .B2(n8606), .A(n8860), .ZN(n8607) );
  AND3_X1 U10005 ( .A1(n8706), .A2(n8625), .A3(n8607), .ZN(n8608) );
  OR3_X1 U10006 ( .A1(n8610), .A2(n8609), .A3(n8608), .ZN(n8664) );
  INV_X1 U10007 ( .A(n8611), .ZN(n8614) );
  INV_X1 U10008 ( .A(n8612), .ZN(n8613) );
  AND3_X1 U10009 ( .A1(n8625), .A2(n8614), .A3(n8613), .ZN(n8707) );
  AND2_X1 U10010 ( .A1(n9028), .A2(n8615), .ZN(n9006) );
  NOR2_X1 U10011 ( .A1(n8664), .A2(n4915), .ZN(n8617) );
  NAND2_X1 U10012 ( .A1(n8856), .A2(n8619), .ZN(n8616) );
  OAI21_X1 U10013 ( .B1(n8663), .B2(n8617), .A(n8616), .ZN(n8620) );
  NAND2_X1 U10014 ( .A1(n8856), .A2(n8869), .ZN(n8650) );
  NAND2_X1 U10015 ( .A1(n8650), .A2(n8618), .ZN(n8662) );
  OR2_X1 U10016 ( .A1(n8856), .A2(n8869), .ZN(n8716) );
  OAI22_X1 U10017 ( .A1(n8620), .A2(n8662), .B1(n8619), .B2(n8716), .ZN(n8621)
         );
  NAND2_X1 U10018 ( .A1(n8621), .A2(n8719), .ZN(n8623) );
  NAND3_X1 U10019 ( .A1(n8623), .A2(n8622), .A3(n8717), .ZN(n8653) );
  INV_X1 U10020 ( .A(n8944), .ZN(n8947) );
  AND2_X1 U10021 ( .A1(n8626), .A2(n8996), .ZN(n9007) );
  NOR2_X1 U10022 ( .A1(n7042), .A2(n8627), .ZN(n8630) );
  NOR2_X1 U10023 ( .A1(n9514), .A2(n8735), .ZN(n8629) );
  NOR2_X1 U10024 ( .A1(n7028), .A2(n9488), .ZN(n8628) );
  NAND4_X1 U10025 ( .A1(n8630), .A2(n8629), .A3(n7157), .A4(n8628), .ZN(n8633)
         );
  NOR4_X1 U10026 ( .A1(n8633), .A2(n8632), .A3(n8631), .A4(n9475), .ZN(n8636)
         );
  NAND4_X1 U10027 ( .A1(n8636), .A2(n8635), .A3(n4872), .A4(n4628), .ZN(n8637)
         );
  OR2_X1 U10028 ( .A1(n8638), .A2(n8637), .ZN(n8639) );
  NOR3_X1 U10029 ( .A1(n8641), .A2(n8640), .A3(n8639), .ZN(n8642) );
  NAND4_X1 U10030 ( .A1(n9046), .A2(n9052), .A3(n9075), .A4(n8642), .ZN(n8643)
         );
  NOR2_X1 U10031 ( .A1(n9031), .A2(n8643), .ZN(n8644) );
  NAND4_X1 U10032 ( .A1(n8974), .A2(n4433), .A3(n9007), .A4(n8644), .ZN(n8645)
         );
  NOR2_X1 U10033 ( .A1(n8645), .A2(n8961), .ZN(n8646) );
  NAND4_X1 U10034 ( .A1(n8937), .A2(n8947), .A3(n8647), .A4(n8646), .ZN(n8648)
         );
  NOR2_X1 U10035 ( .A1(n8878), .A2(n8648), .ZN(n8649) );
  AND2_X1 U10036 ( .A1(n8900), .A2(n8649), .ZN(n8651) );
  AND4_X1 U10037 ( .A1(n8882), .A2(n8716), .A3(n8651), .A4(n8650), .ZN(n8652)
         );
  NAND3_X1 U10038 ( .A1(n8652), .A2(n8719), .A3(n8717), .ZN(n8736) );
  NAND2_X1 U10039 ( .A1(n8653), .A2(n8736), .ZN(n8654) );
  INV_X1 U10040 ( .A(n8732), .ZN(n8721) );
  NAND4_X1 U10041 ( .A1(n8654), .A2(n8721), .A3(n8730), .A4(n4453), .ZN(n8727)
         );
  INV_X1 U10042 ( .A(n8655), .ZN(n8656) );
  NAND3_X1 U10043 ( .A1(n8657), .A2(n9302), .A3(n8656), .ZN(n8661) );
  NAND2_X1 U10044 ( .A1(n8721), .A2(n8658), .ZN(n8659) );
  OAI211_X1 U10045 ( .C1(n8661), .C2(n8660), .A(P1_B_REG_SCAN_IN), .B(n8659), 
        .ZN(n8726) );
  INV_X1 U10046 ( .A(n8662), .ZN(n8715) );
  INV_X1 U10047 ( .A(n8663), .ZN(n8713) );
  INV_X1 U10048 ( .A(n8664), .ZN(n8711) );
  INV_X1 U10049 ( .A(n8665), .ZN(n8709) );
  INV_X1 U10050 ( .A(n8667), .ZN(n8669) );
  AND3_X1 U10051 ( .A1(n8669), .A2(n8735), .A3(n8668), .ZN(n8671) );
  OAI21_X1 U10052 ( .B1(n8666), .B2(n8671), .A(n8670), .ZN(n8677) );
  INV_X1 U10053 ( .A(n8672), .ZN(n8674) );
  NOR2_X1 U10054 ( .A1(n8674), .A2(n8673), .ZN(n8676) );
  AOI21_X1 U10055 ( .B1(n8677), .B2(n8676), .A(n8675), .ZN(n8680) );
  OAI21_X1 U10056 ( .B1(n8680), .B2(n8679), .A(n8678), .ZN(n8682) );
  NAND3_X1 U10057 ( .A1(n8682), .A2(n7163), .A3(n8681), .ZN(n8685) );
  NAND3_X1 U10058 ( .A1(n8685), .A2(n8684), .A3(n8683), .ZN(n8688) );
  INV_X1 U10059 ( .A(n8686), .ZN(n8687) );
  NAND2_X1 U10060 ( .A1(n8688), .A2(n8687), .ZN(n8691) );
  INV_X1 U10061 ( .A(n8689), .ZN(n8690) );
  NAND2_X1 U10062 ( .A1(n8691), .A2(n8690), .ZN(n8694) );
  NAND3_X1 U10063 ( .A1(n8694), .A2(n8693), .A3(n8692), .ZN(n8698) );
  INV_X1 U10064 ( .A(n8695), .ZN(n8697) );
  AND3_X1 U10065 ( .A1(n8698), .A2(n8697), .A3(n8696), .ZN(n8702) );
  OAI211_X1 U10066 ( .C1(n8702), .C2(n8701), .A(n8700), .B(n8699), .ZN(n8704)
         );
  AOI21_X1 U10067 ( .B1(n8705), .B2(n8704), .A(n8703), .ZN(n8708) );
  OAI211_X1 U10068 ( .C1(n8709), .C2(n8708), .A(n8707), .B(n8706), .ZN(n8710)
         );
  NAND2_X1 U10069 ( .A1(n8711), .A2(n8710), .ZN(n8712) );
  NAND2_X1 U10070 ( .A1(n8713), .A2(n8712), .ZN(n8714) );
  NAND2_X1 U10071 ( .A1(n8715), .A2(n8714), .ZN(n8718) );
  NAND3_X1 U10072 ( .A1(n8718), .A2(n8717), .A3(n8716), .ZN(n8720) );
  NAND2_X1 U10073 ( .A1(n8720), .A2(n8719), .ZN(n8723) );
  NAND3_X1 U10074 ( .A1(n8723), .A2(n8722), .A3(n8721), .ZN(n8725) );
  OR4_X1 U10075 ( .A1(n8723), .A2(n8730), .A3(n8732), .A4(n4453), .ZN(n8724)
         );
  NAND2_X1 U10076 ( .A1(n8731), .A2(n8730), .ZN(n8733) );
  AOI211_X1 U10077 ( .C1(n8735), .C2(n8734), .A(n8733), .B(n8732), .ZN(n8737)
         );
  OAI211_X1 U10078 ( .C1(n8739), .C2(n8738), .A(n8737), .B(n8736), .ZN(n8740)
         );
  MUX2_X1 U10079 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n8741), .S(P1_U3973), .Z(
        P1_U3584) );
  INV_X1 U10080 ( .A(n8867), .ZN(n8920) );
  MUX2_X1 U10081 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n8920), .S(P1_U3973), .Z(
        P1_U3582) );
  MUX2_X1 U10082 ( .A(n8939), .B(P1_DATAO_REG_27__SCAN_IN), .S(n8755), .Z(
        P1_U3581) );
  MUX2_X1 U10083 ( .A(n8921), .B(P1_DATAO_REG_26__SCAN_IN), .S(n8755), .Z(
        P1_U3580) );
  MUX2_X1 U10084 ( .A(n8938), .B(P1_DATAO_REG_25__SCAN_IN), .S(n8755), .Z(
        P1_U3579) );
  MUX2_X1 U10085 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n8742), .S(P1_U3973), .Z(
        P1_U3578) );
  MUX2_X1 U10086 ( .A(n8743), .B(P1_DATAO_REG_23__SCAN_IN), .S(n8755), .Z(
        P1_U3577) );
  MUX2_X1 U10087 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n8744), .S(P1_U3973), .Z(
        P1_U3576) );
  MUX2_X1 U10088 ( .A(n8745), .B(P1_DATAO_REG_21__SCAN_IN), .S(n8755), .Z(
        P1_U3575) );
  MUX2_X1 U10089 ( .A(n9047), .B(P1_DATAO_REG_19__SCAN_IN), .S(n8755), .Z(
        P1_U3573) );
  MUX2_X1 U10090 ( .A(n9034), .B(P1_DATAO_REG_18__SCAN_IN), .S(n8755), .Z(
        P1_U3572) );
  MUX2_X1 U10091 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n7828), .S(P1_U3973), .Z(
        P1_U3571) );
  MUX2_X1 U10092 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n8746), .S(P1_U3973), .Z(
        P1_U3570) );
  MUX2_X1 U10093 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9076), .S(P1_U3973), .Z(
        P1_U3569) );
  MUX2_X1 U10094 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n8747), .S(P1_U3973), .Z(
        P1_U3567) );
  MUX2_X1 U10095 ( .A(n8748), .B(P1_DATAO_REG_12__SCAN_IN), .S(n8755), .Z(
        P1_U3566) );
  MUX2_X1 U10096 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n8749), .S(P1_U3973), .Z(
        P1_U3565) );
  MUX2_X1 U10097 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n7359), .S(P1_U3973), .Z(
        P1_U3564) );
  MUX2_X1 U10098 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n8751), .S(P1_U3973), .Z(
        P1_U3563) );
  MUX2_X1 U10099 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n8752), .S(P1_U3973), .Z(
        P1_U3562) );
  MUX2_X1 U10100 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n9468), .S(P1_U3973), .Z(
        P1_U3561) );
  MUX2_X1 U10101 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n8753), .S(P1_U3973), .Z(
        P1_U3560) );
  MUX2_X1 U10102 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n7068), .S(P1_U3973), .Z(
        P1_U3559) );
  MUX2_X1 U10103 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n9491), .S(P1_U3973), .Z(
        P1_U3557) );
  MUX2_X1 U10104 ( .A(n8754), .B(P1_DATAO_REG_2__SCAN_IN), .S(n8755), .Z(
        P1_U3556) );
  MUX2_X1 U10105 ( .A(n6898), .B(P1_DATAO_REG_1__SCAN_IN), .S(n8755), .Z(
        P1_U3555) );
  MUX2_X1 U10106 ( .A(n8756), .B(P1_DATAO_REG_0__SCAN_IN), .S(n8755), .Z(
        P1_U3554) );
  OAI211_X1 U10107 ( .C1(n8759), .C2(n8758), .A(n9446), .B(n8757), .ZN(n8767)
         );
  AOI22_X1 U10108 ( .A1(n9431), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n8766) );
  OAI211_X1 U10109 ( .C1(n8762), .C2(n8761), .A(n9454), .B(n8760), .ZN(n8765)
         );
  NAND2_X1 U10110 ( .A1(n9443), .A2(n8763), .ZN(n8764) );
  NAND4_X1 U10111 ( .A1(n8767), .A2(n8766), .A3(n8765), .A4(n8764), .ZN(
        P1_U3244) );
  INV_X1 U10112 ( .A(n8776), .ZN(n8817) );
  INV_X1 U10113 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n8770) );
  INV_X1 U10114 ( .A(n8768), .ZN(n8769) );
  OAI21_X1 U10115 ( .B1(n9466), .B2(n8770), .A(n8769), .ZN(n8771) );
  AOI21_X1 U10116 ( .B1(n8817), .B2(n9443), .A(n8771), .ZN(n8784) );
  MUX2_X1 U10117 ( .A(n6909), .B(P1_REG2_REG_3__SCAN_IN), .S(n8776), .Z(n8775)
         );
  NAND2_X1 U10118 ( .A1(n8777), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n8772) );
  NAND2_X1 U10119 ( .A1(n8773), .A2(n8772), .ZN(n8774) );
  NAND2_X1 U10120 ( .A1(n8774), .A2(n8775), .ZN(n8819) );
  OAI211_X1 U10121 ( .C1(n8775), .C2(n8774), .A(n9446), .B(n8819), .ZN(n8783)
         );
  INV_X1 U10122 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n9626) );
  MUX2_X1 U10123 ( .A(n9626), .B(P1_REG1_REG_3__SCAN_IN), .S(n8776), .Z(n8781)
         );
  NAND2_X1 U10124 ( .A1(n8777), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n8778) );
  NAND2_X1 U10125 ( .A1(n8779), .A2(n8778), .ZN(n8780) );
  NAND2_X1 U10126 ( .A1(n8780), .A2(n8781), .ZN(n8791) );
  OAI211_X1 U10127 ( .C1(n8781), .C2(n8780), .A(n9454), .B(n8791), .ZN(n8782)
         );
  NAND3_X1 U10128 ( .A1(n8784), .A2(n8783), .A3(n8782), .ZN(P1_U3246) );
  INV_X1 U10129 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n8785) );
  AOI22_X1 U10130 ( .A1(n9435), .A2(P1_REG1_REG_16__SCAN_IN), .B1(n8785), .B2(
        n8838), .ZN(n9434) );
  INV_X1 U10131 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n8786) );
  MUX2_X1 U10132 ( .A(n8786), .B(P1_REG1_REG_13__SCAN_IN), .S(n8833), .Z(n9388) );
  OR2_X1 U10133 ( .A1(n8832), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n8803) );
  OR2_X1 U10134 ( .A1(n8830), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n8788) );
  NAND2_X1 U10135 ( .A1(n8830), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n8787) );
  NAND2_X1 U10136 ( .A1(n8788), .A2(n8787), .ZN(n9224) );
  OR2_X1 U10137 ( .A1(n8829), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n8800) );
  NOR2_X1 U10138 ( .A1(n8829), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n8789) );
  AOI21_X1 U10139 ( .B1(n8829), .B2(P1_REG1_REG_9__SCAN_IN), .A(n8789), .ZN(
        n9269) );
  NAND2_X1 U10140 ( .A1(n8817), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n8790) );
  NAND2_X1 U10141 ( .A1(n8791), .A2(n8790), .ZN(n9308) );
  NAND2_X1 U10142 ( .A1(n9318), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n8792) );
  OAI21_X1 U10143 ( .B1(n9318), .B2(P1_REG1_REG_4__SCAN_IN), .A(n8792), .ZN(
        n9310) );
  INV_X1 U10144 ( .A(n9310), .ZN(n8793) );
  AND2_X1 U10145 ( .A1(n9318), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n8794) );
  NOR2_X1 U10146 ( .A1(n9309), .A2(n8794), .ZN(n9328) );
  INV_X1 U10147 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n8795) );
  MUX2_X1 U10148 ( .A(n8795), .B(P1_REG1_REG_5__SCAN_IN), .S(n8823), .Z(n9327)
         );
  NOR2_X1 U10149 ( .A1(n9328), .A2(n9327), .ZN(n9326) );
  AOI21_X1 U10150 ( .B1(n8823), .B2(P1_REG1_REG_5__SCAN_IN), .A(n9326), .ZN(
        n9342) );
  NAND2_X1 U10151 ( .A1(n8825), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n8796) );
  OAI21_X1 U10152 ( .B1(n8825), .B2(P1_REG1_REG_6__SCAN_IN), .A(n8796), .ZN(
        n9341) );
  NOR2_X1 U10153 ( .A1(n9342), .A2(n9341), .ZN(n9340) );
  AOI21_X1 U10154 ( .B1(n8825), .B2(P1_REG1_REG_6__SCAN_IN), .A(n9340), .ZN(
        n9238) );
  INV_X1 U10155 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n8797) );
  MUX2_X1 U10156 ( .A(n8797), .B(P1_REG1_REG_7__SCAN_IN), .S(n8826), .Z(n9239)
         );
  NOR2_X1 U10157 ( .A1(n9238), .A2(n9239), .ZN(n9237) );
  AOI21_X1 U10158 ( .B1(n8826), .B2(P1_REG1_REG_7__SCAN_IN), .A(n9237), .ZN(
        n9253) );
  OR2_X1 U10159 ( .A1(n8828), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n8799) );
  NAND2_X1 U10160 ( .A1(n8828), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n8798) );
  NAND2_X1 U10161 ( .A1(n8799), .A2(n8798), .ZN(n9254) );
  NOR2_X1 U10162 ( .A1(n9253), .A2(n9254), .ZN(n9252) );
  AOI21_X1 U10163 ( .B1(n8828), .B2(P1_REG1_REG_8__SCAN_IN), .A(n9252), .ZN(
        n9268) );
  NAND2_X1 U10164 ( .A1(n9269), .A2(n9268), .ZN(n9267) );
  NAND2_X1 U10165 ( .A1(n8800), .A2(n9267), .ZN(n9223) );
  NOR2_X1 U10166 ( .A1(n9224), .A2(n9223), .ZN(n9222) );
  AOI21_X1 U10167 ( .B1(n8830), .B2(P1_REG1_REG_10__SCAN_IN), .A(n9222), .ZN(
        n9357) );
  INV_X1 U10168 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n8801) );
  MUX2_X1 U10169 ( .A(n8801), .B(P1_REG1_REG_11__SCAN_IN), .S(n9351), .Z(n9358) );
  NOR2_X1 U10170 ( .A1(n9357), .A2(n9358), .ZN(n9356) );
  AOI21_X1 U10171 ( .B1(n9351), .B2(P1_REG1_REG_11__SCAN_IN), .A(n9356), .ZN(
        n9372) );
  INV_X1 U10172 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n8802) );
  MUX2_X1 U10173 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n8802), .S(n8832), .Z(n9373) );
  NAND2_X1 U10174 ( .A1(n9372), .A2(n9373), .ZN(n9371) );
  NAND2_X1 U10175 ( .A1(n8803), .A2(n9371), .ZN(n9387) );
  NOR2_X1 U10176 ( .A1(n9388), .A2(n9387), .ZN(n9386) );
  AOI21_X1 U10177 ( .B1(n8833), .B2(P1_REG1_REG_13__SCAN_IN), .A(n9386), .ZN(
        n9404) );
  INV_X1 U10178 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n8804) );
  OR2_X1 U10179 ( .A1(n9397), .A2(n8804), .ZN(n8806) );
  NAND2_X1 U10180 ( .A1(n9397), .A2(n8804), .ZN(n8805) );
  AND2_X1 U10181 ( .A1(n8806), .A2(n8805), .ZN(n9403) );
  NOR2_X1 U10182 ( .A1(n9404), .A2(n9403), .ZN(n9402) );
  AOI21_X1 U10183 ( .B1(P1_REG1_REG_14__SCAN_IN), .B2(n9397), .A(n9402), .ZN(
        n8807) );
  NOR2_X1 U10184 ( .A1(n8807), .A2(n8836), .ZN(n8808) );
  INV_X1 U10185 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n9415) );
  XNOR2_X1 U10186 ( .A(n8836), .B(n8807), .ZN(n9416) );
  NOR2_X1 U10187 ( .A1(n9415), .A2(n9416), .ZN(n9414) );
  NOR2_X1 U10188 ( .A1(n8808), .A2(n9414), .ZN(n9433) );
  NAND2_X1 U10189 ( .A1(n9434), .A2(n9433), .ZN(n9432) );
  OAI21_X1 U10190 ( .B1(n9435), .B2(P1_REG1_REG_16__SCAN_IN), .A(n9432), .ZN(
        n9442) );
  INV_X1 U10191 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n8810) );
  XNOR2_X1 U10192 ( .A(n9444), .B(n8810), .ZN(n9441) );
  AOI22_X1 U10193 ( .A1(n9442), .A2(n9441), .B1(n8810), .B2(n8809), .ZN(n9457)
         );
  INV_X1 U10194 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n8811) );
  AND2_X1 U10195 ( .A1(n8842), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n8812) );
  AOI21_X1 U10196 ( .B1(n8811), .B2(n9459), .A(n8812), .ZN(n9456) );
  NAND2_X1 U10197 ( .A1(n9457), .A2(n9456), .ZN(n9455) );
  INV_X1 U10198 ( .A(n8812), .ZN(n8813) );
  NAND2_X1 U10199 ( .A1(n9455), .A2(n8813), .ZN(n8814) );
  XOR2_X1 U10200 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n8814), .Z(n8846) );
  AOI22_X1 U10201 ( .A1(n8833), .A2(n7489), .B1(P1_REG2_REG_13__SCAN_IN), .B2(
        n9392), .ZN(n9384) );
  AOI22_X1 U10202 ( .A1(n8832), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n7405), .B2(
        n9377), .ZN(n9369) );
  NAND2_X1 U10203 ( .A1(n8830), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n8815) );
  OAI21_X1 U10204 ( .B1(n8830), .B2(P1_REG2_REG_10__SCAN_IN), .A(n8815), .ZN(
        n9220) );
  NOR2_X1 U10205 ( .A1(n8829), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n8816) );
  AOI21_X1 U10206 ( .B1(P1_REG2_REG_9__SCAN_IN), .B2(n8829), .A(n8816), .ZN(
        n9265) );
  NAND2_X1 U10207 ( .A1(n8817), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n8818) );
  NAND2_X1 U10208 ( .A1(n8819), .A2(n8818), .ZN(n9312) );
  NAND2_X1 U10209 ( .A1(n9318), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n8820) );
  OAI21_X1 U10210 ( .B1(n9318), .B2(P1_REG2_REG_4__SCAN_IN), .A(n8820), .ZN(
        n9314) );
  INV_X1 U10211 ( .A(n9314), .ZN(n8821) );
  INV_X1 U10212 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n8822) );
  AOI22_X1 U10213 ( .A1(n8823), .A2(n8822), .B1(P1_REG2_REG_5__SCAN_IN), .B2(
        n9332), .ZN(n9324) );
  NAND2_X1 U10214 ( .A1(n8825), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n8824) );
  OAI21_X1 U10215 ( .B1(n8825), .B2(P1_REG2_REG_6__SCAN_IN), .A(n8824), .ZN(
        n9338) );
  NOR2_X1 U10216 ( .A1(n4395), .A2(n9338), .ZN(n9337) );
  AOI21_X1 U10217 ( .B1(P1_REG2_REG_6__SCAN_IN), .B2(n8825), .A(n9337), .ZN(
        n9234) );
  AOI22_X1 U10218 ( .A1(n8826), .A2(n7210), .B1(P1_REG2_REG_7__SCAN_IN), .B2(
        n9243), .ZN(n9235) );
  NOR2_X1 U10219 ( .A1(n9234), .A2(n9235), .ZN(n9233) );
  NAND2_X1 U10220 ( .A1(n8828), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n8827) );
  OAI21_X1 U10221 ( .B1(n8828), .B2(P1_REG2_REG_8__SCAN_IN), .A(n8827), .ZN(
        n9250) );
  OAI21_X1 U10222 ( .B1(n8829), .B2(P1_REG2_REG_9__SCAN_IN), .A(n9263), .ZN(
        n9219) );
  NOR2_X1 U10223 ( .A1(n9220), .A2(n9219), .ZN(n9218) );
  NAND2_X1 U10224 ( .A1(n9351), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n8831) );
  OAI21_X1 U10225 ( .B1(n9351), .B2(P1_REG2_REG_11__SCAN_IN), .A(n8831), .ZN(
        n9354) );
  OAI21_X1 U10226 ( .B1(n8832), .B2(P1_REG2_REG_12__SCAN_IN), .A(n9367), .ZN(
        n9383) );
  NOR2_X1 U10227 ( .A1(n9384), .A2(n9383), .ZN(n9382) );
  NAND2_X1 U10228 ( .A1(n9397), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n8834) );
  OAI21_X1 U10229 ( .B1(n9397), .B2(P1_REG2_REG_14__SCAN_IN), .A(n8834), .ZN(
        n9400) );
  NOR2_X1 U10230 ( .A1(n8835), .A2(n8836), .ZN(n8837) );
  NOR2_X1 U10231 ( .A1(n9418), .A2(n9419), .ZN(n9417) );
  NOR2_X1 U10232 ( .A1(n8837), .A2(n9417), .ZN(n9428) );
  INV_X1 U10233 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n8839) );
  AOI22_X1 U10234 ( .A1(n9435), .A2(n8839), .B1(P1_REG2_REG_16__SCAN_IN), .B2(
        n8838), .ZN(n9427) );
  NOR2_X1 U10235 ( .A1(n9428), .A2(n9427), .ZN(n9426) );
  INV_X1 U10236 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n8840) );
  XNOR2_X1 U10237 ( .A(n9444), .B(n8840), .ZN(n9439) );
  OR2_X1 U10238 ( .A1(n9444), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n8841) );
  NAND2_X1 U10239 ( .A1(n8842), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n8843) );
  OAI21_X1 U10240 ( .B1(n8842), .B2(P1_REG2_REG_18__SCAN_IN), .A(n8843), .ZN(
        n9452) );
  NAND2_X1 U10241 ( .A1(n9462), .A2(n8843), .ZN(n8844) );
  XNOR2_X1 U10242 ( .A(n8844), .B(P1_REG2_REG_19__SCAN_IN), .ZN(n8848) );
  NAND2_X1 U10243 ( .A1(n8848), .A2(n9446), .ZN(n8845) );
  INV_X1 U10244 ( .A(n8846), .ZN(n8847) );
  OAI22_X1 U10245 ( .A1(n8848), .A2(n9451), .B1(n8847), .B2(n9413), .ZN(n8849)
         );
  NOR2_X1 U10246 ( .A1(n9093), .A2(n9485), .ZN(n8857) );
  NOR2_X1 U10247 ( .A1(n8851), .A2(n9067), .ZN(n8852) );
  AOI211_X1 U10248 ( .C1(n9485), .C2(P1_REG2_REG_31__SCAN_IN), .A(n8857), .B(
        n8852), .ZN(n8853) );
  OAI21_X1 U10249 ( .B1(n8854), .B2(n9085), .A(n8853), .ZN(P1_U3263) );
  INV_X1 U10250 ( .A(n8856), .ZN(n9095) );
  AOI21_X1 U10251 ( .B1(n8856), .B2(n8886), .A(n8855), .ZN(n9092) );
  NAND2_X1 U10252 ( .A1(n9092), .A2(n9037), .ZN(n8859) );
  AOI21_X1 U10253 ( .B1(n9485), .B2(P1_REG2_REG_30__SCAN_IN), .A(n8857), .ZN(
        n8858) );
  OAI211_X1 U10254 ( .C1(n9095), .C2(n9067), .A(n8859), .B(n8858), .ZN(
        P1_U3264) );
  NAND2_X1 U10255 ( .A1(n8861), .A2(n8860), .ZN(n8936) );
  NAND2_X1 U10256 ( .A1(n8936), .A2(n8937), .ZN(n8935) );
  NAND2_X1 U10257 ( .A1(n8935), .A2(n8862), .ZN(n8918) );
  INV_X1 U10258 ( .A(n8882), .ZN(n8865) );
  XNOR2_X1 U10259 ( .A(n8866), .B(n8865), .ZN(n8872) );
  NOR2_X1 U10260 ( .A1(n9119), .A2(n8938), .ZN(n8874) );
  NOR2_X1 U10261 ( .A1(n8934), .A2(n8876), .ZN(n8877) );
  OAI22_X2 U10262 ( .A1(n8929), .A2(n8877), .B1(n8921), .B2(n9114), .ZN(n8910)
         );
  NAND2_X1 U10263 ( .A1(n8916), .A2(n8897), .ZN(n8879) );
  INV_X1 U10264 ( .A(n8900), .ZN(n8880) );
  NAND2_X1 U10265 ( .A1(n9103), .A2(n8920), .ZN(n8881) );
  NAND2_X1 U10266 ( .A1(n8902), .A2(n8881), .ZN(n8883) );
  XNOR2_X1 U10267 ( .A(n8883), .B(n8882), .ZN(n9096) );
  NAND2_X1 U10268 ( .A1(n9096), .A2(n9482), .ZN(n8892) );
  OAI22_X1 U10269 ( .A1(n8885), .A2(n9499), .B1(n8884), .B2(n9510), .ZN(n8889)
         );
  NOR2_X1 U10270 ( .A1(n9098), .A2(n8887), .ZN(n8888) );
  AOI211_X1 U10271 ( .C1(n9472), .C2(n8890), .A(n8889), .B(n8888), .ZN(n8891)
         );
  OAI211_X1 U10272 ( .C1(n4399), .C2(n9485), .A(n8892), .B(n8891), .ZN(
        P1_U3356) );
  OAI21_X1 U10273 ( .B1(n8900), .B2(n8894), .A(n8893), .ZN(n8895) );
  INV_X1 U10274 ( .A(n8895), .ZN(n8896) );
  OAI222_X1 U10275 ( .A1(n9060), .A2(n8898), .B1(n9062), .B2(n8897), .C1(n9516), .C2(n8896), .ZN(n9101) );
  INV_X1 U10276 ( .A(n9101), .ZN(n8909) );
  NAND2_X1 U10277 ( .A1(n8899), .A2(n8900), .ZN(n8901) );
  NAND2_X1 U10278 ( .A1(n9102), .A2(n9482), .ZN(n8908) );
  AOI211_X1 U10279 ( .C1(n9103), .C2(n8911), .A(n9568), .B(n8903), .ZN(n9105)
         );
  AOI22_X1 U10280 ( .A1(n8904), .A2(n9471), .B1(P1_REG2_REG_28__SCAN_IN), .B2(
        n9485), .ZN(n8905) );
  OAI21_X1 U10281 ( .B1(n4482), .B2(n9067), .A(n8905), .ZN(n8906) );
  AOI21_X1 U10282 ( .B1(n9105), .B2(n9480), .A(n8906), .ZN(n8907) );
  OAI211_X1 U10283 ( .C1(n9485), .C2(n8909), .A(n8908), .B(n8907), .ZN(
        P1_U3265) );
  XNOR2_X1 U10284 ( .A(n8910), .B(n8919), .ZN(n9112) );
  INV_X1 U10285 ( .A(n8930), .ZN(n8913) );
  INV_X1 U10286 ( .A(n8911), .ZN(n8912) );
  AOI211_X1 U10287 ( .C1(n9109), .C2(n8913), .A(n9568), .B(n8912), .ZN(n9108)
         );
  AOI22_X1 U10288 ( .A1(n8914), .A2(n9471), .B1(P1_REG2_REG_27__SCAN_IN), .B2(
        n9485), .ZN(n8915) );
  OAI21_X1 U10289 ( .B1(n8916), .B2(n9067), .A(n8915), .ZN(n8927) );
  OAI21_X1 U10290 ( .B1(n8919), .B2(n8918), .A(n8917), .ZN(n8925) );
  NAND2_X1 U10291 ( .A1(n8921), .A2(n9489), .ZN(n8922) );
  AOI211_X1 U10292 ( .C1(n9480), .C2(n9108), .A(n8927), .B(n8926), .ZN(n8928)
         );
  OAI21_X1 U10293 ( .B1(n9112), .B2(n9071), .A(n8928), .ZN(P1_U3266) );
  XOR2_X1 U10294 ( .A(n8937), .B(n8929), .Z(n9117) );
  AOI211_X1 U10295 ( .C1(n9114), .C2(n8931), .A(n9568), .B(n8930), .ZN(n9113)
         );
  AOI22_X1 U10296 ( .A1(n8932), .A2(n9471), .B1(P1_REG2_REG_26__SCAN_IN), .B2(
        n9485), .ZN(n8933) );
  OAI21_X1 U10297 ( .B1(n8934), .B2(n9067), .A(n8933), .ZN(n8942) );
  OAI21_X1 U10298 ( .B1(n8937), .B2(n8936), .A(n8935), .ZN(n8940) );
  AOI222_X1 U10299 ( .A1(n9493), .A2(n8940), .B1(n8939), .B2(n9490), .C1(n8938), .C2(n9489), .ZN(n9116) );
  NOR2_X1 U10300 ( .A1(n9116), .A2(n9485), .ZN(n8941) );
  AOI211_X1 U10301 ( .C1(n9113), .C2(n9480), .A(n8942), .B(n8941), .ZN(n8943)
         );
  OAI21_X1 U10302 ( .B1(n9117), .B2(n9071), .A(n8943), .ZN(P1_U3267) );
  XNOR2_X1 U10303 ( .A(n8945), .B(n8944), .ZN(n9127) );
  NOR2_X1 U10304 ( .A1(n8946), .A2(n4565), .ZN(n8948) );
  XNOR2_X1 U10305 ( .A(n8948), .B(n8947), .ZN(n8949) );
  OAI222_X1 U10306 ( .A1(n9060), .A2(n8950), .B1(n9062), .B2(n8980), .C1(n8949), .C2(n9516), .ZN(n9123) );
  INV_X1 U10307 ( .A(n8965), .ZN(n8952) );
  AOI211_X1 U10308 ( .C1(n9125), .C2(n8952), .A(n9568), .B(n4488), .ZN(n9124)
         );
  NAND2_X1 U10309 ( .A1(n9124), .A2(n9480), .ZN(n8956) );
  INV_X1 U10310 ( .A(n8953), .ZN(n8954) );
  AOI22_X1 U10311 ( .A1(n8954), .A2(n9471), .B1(P1_REG2_REG_24__SCAN_IN), .B2(
        n9485), .ZN(n8955) );
  OAI211_X1 U10312 ( .C1(n8957), .C2(n9067), .A(n8956), .B(n8955), .ZN(n8958)
         );
  AOI21_X1 U10313 ( .B1(n9123), .B2(n9510), .A(n8958), .ZN(n8959) );
  OAI21_X1 U10314 ( .B1(n9127), .B2(n9071), .A(n8959), .ZN(P1_U3269) );
  XNOR2_X1 U10315 ( .A(n8960), .B(n8961), .ZN(n9132) );
  AOI21_X1 U10316 ( .B1(n8962), .B2(n8961), .A(n8946), .ZN(n8963) );
  OAI222_X1 U10317 ( .A1(n9062), .A2(n9002), .B1(n9060), .B2(n8964), .C1(n9516), .C2(n8963), .ZN(n9128) );
  INV_X1 U10318 ( .A(n8981), .ZN(n8966) );
  AOI211_X1 U10319 ( .C1(n9130), .C2(n8966), .A(n9568), .B(n8965), .ZN(n9129)
         );
  NAND2_X1 U10320 ( .A1(n9129), .A2(n9480), .ZN(n8970) );
  INV_X1 U10321 ( .A(n8967), .ZN(n8968) );
  AOI22_X1 U10322 ( .A1(n8968), .A2(n9471), .B1(n9485), .B2(
        P1_REG2_REG_23__SCAN_IN), .ZN(n8969) );
  OAI211_X1 U10323 ( .C1(n8971), .C2(n9067), .A(n8970), .B(n8969), .ZN(n8972)
         );
  AOI21_X1 U10324 ( .B1(n9128), .B2(n9510), .A(n8972), .ZN(n8973) );
  OAI21_X1 U10325 ( .B1(n9132), .B2(n9071), .A(n8973), .ZN(P1_U3270) );
  XNOR2_X1 U10326 ( .A(n8975), .B(n8974), .ZN(n9137) );
  AOI21_X1 U10327 ( .B1(n8978), .B2(n8977), .A(n8976), .ZN(n8979) );
  OAI222_X1 U10328 ( .A1(n9060), .A2(n8980), .B1(n9062), .B2(n9010), .C1(n9516), .C2(n8979), .ZN(n9133) );
  INV_X1 U10329 ( .A(n9135), .ZN(n8985) );
  AOI211_X1 U10330 ( .C1(n9135), .C2(n8989), .A(n9568), .B(n8981), .ZN(n9134)
         );
  NAND2_X1 U10331 ( .A1(n9134), .A2(n9480), .ZN(n8984) );
  AOI22_X1 U10332 ( .A1(n9485), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n8982), .B2(
        n9471), .ZN(n8983) );
  OAI211_X1 U10333 ( .C1(n8985), .C2(n9067), .A(n8984), .B(n8983), .ZN(n8986)
         );
  AOI21_X1 U10334 ( .B1(n9133), .B2(n9510), .A(n8986), .ZN(n8987) );
  OAI21_X1 U10335 ( .B1(n9137), .B2(n9071), .A(n8987), .ZN(P1_U3271) );
  XNOR2_X1 U10336 ( .A(n8988), .B(n4433), .ZN(n9142) );
  INV_X1 U10337 ( .A(n8989), .ZN(n8990) );
  AOI211_X1 U10338 ( .C1(n9140), .C2(n9011), .A(n9568), .B(n8990), .ZN(n9139)
         );
  NOR2_X1 U10339 ( .A1(n8991), .A2(n9067), .ZN(n8995) );
  OAI22_X1 U10340 ( .A1(n9510), .A2(n8993), .B1(n8992), .B2(n9499), .ZN(n8994)
         );
  AOI211_X1 U10341 ( .C1(n9139), .C2(n9480), .A(n8995), .B(n8994), .ZN(n9004)
         );
  INV_X1 U10342 ( .A(n8996), .ZN(n8997) );
  NOR2_X1 U10343 ( .A1(n4433), .A2(n8997), .ZN(n9000) );
  AOI21_X1 U10344 ( .B1(n9000), .B2(n8999), .A(n8998), .ZN(n9001) );
  OAI222_X1 U10345 ( .A1(n9060), .A2(n9002), .B1(n9062), .B2(n9026), .C1(n9516), .C2(n9001), .ZN(n9138) );
  NAND2_X1 U10346 ( .A1(n9138), .A2(n9510), .ZN(n9003) );
  OAI211_X1 U10347 ( .C1(n9142), .C2(n9071), .A(n9004), .B(n9003), .ZN(
        P1_U3272) );
  XOR2_X1 U10348 ( .A(n9007), .B(n9005), .Z(n9147) );
  XOR2_X1 U10349 ( .A(n9007), .B(n9006), .Z(n9008) );
  OAI222_X1 U10350 ( .A1(n9060), .A2(n9010), .B1(n9062), .B2(n9009), .C1(n9516), .C2(n9008), .ZN(n9143) );
  INV_X1 U10351 ( .A(n9021), .ZN(n9013) );
  INV_X1 U10352 ( .A(n9011), .ZN(n9012) );
  AOI211_X1 U10353 ( .C1(n9145), .C2(n9013), .A(n9568), .B(n9012), .ZN(n9144)
         );
  NAND2_X1 U10354 ( .A1(n9144), .A2(n9480), .ZN(n9016) );
  AOI22_X1 U10355 ( .A1(n9485), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9014), .B2(
        n9471), .ZN(n9015) );
  OAI211_X1 U10356 ( .C1(n9017), .C2(n9067), .A(n9016), .B(n9015), .ZN(n9018)
         );
  AOI21_X1 U10357 ( .B1(n9143), .B2(n9510), .A(n9018), .ZN(n9019) );
  OAI21_X1 U10358 ( .B1(n9147), .B2(n9071), .A(n9019), .ZN(P1_U3273) );
  XOR2_X1 U10359 ( .A(n9020), .B(n9031), .Z(n9152) );
  INV_X1 U10360 ( .A(n9040), .ZN(n9022) );
  AOI21_X1 U10361 ( .B1(n9148), .B2(n9022), .A(n9021), .ZN(n9149) );
  AOI22_X1 U10362 ( .A1(n9485), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9023), .B2(
        n9471), .ZN(n9024) );
  OAI21_X1 U10363 ( .B1(n9025), .B2(n9067), .A(n9024), .ZN(n9036) );
  NOR2_X1 U10364 ( .A1(n9026), .A2(n9060), .ZN(n9033) );
  NAND2_X1 U10365 ( .A1(n9045), .A2(n9027), .ZN(n9030) );
  INV_X1 U10366 ( .A(n9028), .ZN(n9029) );
  AOI211_X1 U10367 ( .C1(n9031), .C2(n9030), .A(n9516), .B(n9029), .ZN(n9032)
         );
  AOI211_X1 U10368 ( .C1(n9489), .C2(n9034), .A(n9033), .B(n9032), .ZN(n9151)
         );
  NOR2_X1 U10369 ( .A1(n9151), .A2(n9485), .ZN(n9035) );
  AOI211_X1 U10370 ( .C1(n9149), .C2(n9037), .A(n9036), .B(n9035), .ZN(n9038)
         );
  OAI21_X1 U10371 ( .B1(n9152), .B2(n9071), .A(n9038), .ZN(P1_U3274) );
  XNOR2_X1 U10372 ( .A(n9039), .B(n9046), .ZN(n9157) );
  AOI211_X1 U10373 ( .C1(n9154), .C2(n9063), .A(n9568), .B(n9040), .ZN(n9153)
         );
  INV_X1 U10374 ( .A(n9154), .ZN(n9043) );
  AOI22_X1 U10375 ( .A1(n9485), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9041), .B2(
        n9471), .ZN(n9042) );
  OAI21_X1 U10376 ( .B1(n9043), .B2(n9067), .A(n9042), .ZN(n9050) );
  OAI21_X1 U10377 ( .B1(n9046), .B2(n9044), .A(n9045), .ZN(n9048) );
  AOI222_X1 U10378 ( .A1(n9493), .A2(n9048), .B1(n9047), .B2(n9490), .C1(n7828), .C2(n9489), .ZN(n9156) );
  NOR2_X1 U10379 ( .A1(n9156), .A2(n9485), .ZN(n9049) );
  AOI211_X1 U10380 ( .C1(n9153), .C2(n9480), .A(n9050), .B(n9049), .ZN(n9051)
         );
  OAI21_X1 U10381 ( .B1(n9157), .B2(n9071), .A(n9051), .ZN(P1_U3275) );
  XNOR2_X1 U10382 ( .A(n9053), .B(n9052), .ZN(n9161) );
  INV_X1 U10383 ( .A(n9054), .ZN(n9055) );
  AOI21_X1 U10384 ( .B1(n9057), .B2(n9056), .A(n9055), .ZN(n9058) );
  OAI222_X1 U10385 ( .A1(n9062), .A2(n9061), .B1(n9060), .B2(n9059), .C1(n9516), .C2(n9058), .ZN(n9158) );
  AOI211_X1 U10386 ( .C1(n7829), .C2(n9078), .A(n9568), .B(n5182), .ZN(n9159)
         );
  NAND2_X1 U10387 ( .A1(n9159), .A2(n9480), .ZN(n9066) );
  AOI22_X1 U10388 ( .A1(n9485), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9064), .B2(
        n9471), .ZN(n9065) );
  OAI211_X1 U10389 ( .C1(n9068), .C2(n9067), .A(n9066), .B(n9065), .ZN(n9069)
         );
  AOI21_X1 U10390 ( .B1(n9158), .B2(n9510), .A(n9069), .ZN(n9070) );
  OAI21_X1 U10391 ( .B1(n9161), .B2(n9071), .A(n9070), .ZN(P1_U3276) );
  AOI21_X1 U10392 ( .B1(n9075), .B2(n9073), .A(n9072), .ZN(n9166) );
  XOR2_X1 U10393 ( .A(n9074), .B(n9075), .Z(n9077) );
  AOI222_X1 U10394 ( .A1(n9493), .A2(n9077), .B1(n7828), .B2(n9490), .C1(n9076), .C2(n9489), .ZN(n9163) );
  NOR2_X1 U10395 ( .A1(n9163), .A2(n9485), .ZN(n9087) );
  OAI211_X1 U10396 ( .C1(n9079), .C2(n9164), .A(n9496), .B(n9078), .ZN(n9162)
         );
  INV_X1 U10397 ( .A(n9080), .ZN(n9081) );
  OAI22_X1 U10398 ( .A1(n9510), .A2(n8839), .B1(n9081), .B2(n9499), .ZN(n9082)
         );
  AOI21_X1 U10399 ( .B1(n9083), .B2(n9472), .A(n9082), .ZN(n9084) );
  OAI21_X1 U10400 ( .B1(n9162), .B2(n9085), .A(n9084), .ZN(n9086) );
  AOI211_X1 U10401 ( .C1(n9166), .C2(n9482), .A(n9087), .B(n9086), .ZN(n9088)
         );
  INV_X1 U10402 ( .A(n9088), .ZN(P1_U3277) );
  INV_X2 U10403 ( .A(n9644), .ZN(n9630) );
  MUX2_X1 U10404 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n9091), .S(n9630), .Z(
        P1_U3553) );
  NAND2_X1 U10405 ( .A1(n9092), .A2(n9496), .ZN(n9094) );
  OAI211_X1 U10406 ( .C1(n9095), .C2(n9613), .A(n9094), .B(n9093), .ZN(n9168)
         );
  MUX2_X1 U10407 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n9168), .S(n9630), .Z(
        P1_U3552) );
  INV_X1 U10408 ( .A(n9565), .ZN(n9593) );
  NAND2_X1 U10409 ( .A1(n9096), .A2(n9617), .ZN(n9100) );
  OAI22_X1 U10410 ( .A1(n9098), .A2(n9568), .B1(n9097), .B2(n9613), .ZN(n9099)
         );
  MUX2_X1 U10411 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n9169), .S(n9630), .Z(
        P1_U3551) );
  NAND2_X1 U10412 ( .A1(n9102), .A2(n9617), .ZN(n9107) );
  NAND3_X1 U10413 ( .A1(n8909), .A2(n9107), .A3(n9106), .ZN(n9170) );
  MUX2_X1 U10414 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9170), .S(n9630), .Z(
        P1_U3550) );
  OAI211_X1 U10415 ( .C1(n9112), .C2(n9538), .A(n9111), .B(n9110), .ZN(n9171)
         );
  MUX2_X1 U10416 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9171), .S(n9630), .Z(
        P1_U3549) );
  AOI21_X1 U10417 ( .B1(n9591), .B2(n9114), .A(n9113), .ZN(n9115) );
  OAI211_X1 U10418 ( .C1(n9117), .C2(n9538), .A(n9116), .B(n9115), .ZN(n9172)
         );
  MUX2_X1 U10419 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9172), .S(n9630), .Z(
        P1_U3548) );
  AOI21_X1 U10420 ( .B1(n9591), .B2(n9119), .A(n9118), .ZN(n9120) );
  OAI211_X1 U10421 ( .C1(n9122), .C2(n9538), .A(n9121), .B(n9120), .ZN(n9173)
         );
  MUX2_X1 U10422 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9173), .S(n9630), .Z(
        P1_U3547) );
  AOI211_X1 U10423 ( .C1(n9591), .C2(n9125), .A(n9124), .B(n9123), .ZN(n9126)
         );
  OAI21_X1 U10424 ( .B1(n9127), .B2(n9538), .A(n9126), .ZN(n9174) );
  MUX2_X1 U10425 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9174), .S(n9630), .Z(
        P1_U3546) );
  AOI211_X1 U10426 ( .C1(n9591), .C2(n9130), .A(n9129), .B(n9128), .ZN(n9131)
         );
  OAI21_X1 U10427 ( .B1(n9132), .B2(n9538), .A(n9131), .ZN(n9175) );
  MUX2_X1 U10428 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9175), .S(n9630), .Z(
        P1_U3545) );
  AOI211_X1 U10429 ( .C1(n9591), .C2(n9135), .A(n9134), .B(n9133), .ZN(n9136)
         );
  OAI21_X1 U10430 ( .B1(n9137), .B2(n9538), .A(n9136), .ZN(n9176) );
  MUX2_X1 U10431 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9176), .S(n9630), .Z(
        P1_U3544) );
  AOI211_X1 U10432 ( .C1(n9591), .C2(n9140), .A(n9139), .B(n9138), .ZN(n9141)
         );
  OAI21_X1 U10433 ( .B1(n9142), .B2(n9538), .A(n9141), .ZN(n9177) );
  MUX2_X1 U10434 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9177), .S(n9630), .Z(
        P1_U3543) );
  AOI211_X1 U10435 ( .C1(n9591), .C2(n9145), .A(n9144), .B(n9143), .ZN(n9146)
         );
  OAI21_X1 U10436 ( .B1(n9147), .B2(n9538), .A(n9146), .ZN(n9178) );
  MUX2_X1 U10437 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9178), .S(n9630), .Z(
        P1_U3542) );
  AOI22_X1 U10438 ( .A1(n9149), .A2(n9496), .B1(n9591), .B2(n9148), .ZN(n9150)
         );
  OAI211_X1 U10439 ( .C1(n9152), .C2(n9538), .A(n9151), .B(n9150), .ZN(n9179)
         );
  MUX2_X1 U10440 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9179), .S(n9630), .Z(
        P1_U3541) );
  AOI21_X1 U10441 ( .B1(n9591), .B2(n9154), .A(n9153), .ZN(n9155) );
  OAI211_X1 U10442 ( .C1(n9157), .C2(n9538), .A(n9156), .B(n9155), .ZN(n9180)
         );
  MUX2_X1 U10443 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9180), .S(n9630), .Z(
        P1_U3540) );
  AOI211_X1 U10444 ( .C1(n9591), .C2(n7829), .A(n9159), .B(n9158), .ZN(n9160)
         );
  OAI21_X1 U10445 ( .B1(n9161), .B2(n9538), .A(n9160), .ZN(n9181) );
  MUX2_X1 U10446 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9181), .S(n9630), .Z(
        P1_U3539) );
  OAI211_X1 U10447 ( .C1(n9164), .C2(n9613), .A(n9163), .B(n9162), .ZN(n9165)
         );
  AOI21_X1 U10448 ( .B1(n9166), .B2(n9617), .A(n9165), .ZN(n9167) );
  INV_X1 U10449 ( .A(n9167), .ZN(n9182) );
  MUX2_X1 U10450 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9182), .S(n9630), .Z(
        P1_U3538) );
  MUX2_X1 U10451 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n9168), .S(n9546), .Z(
        P1_U3520) );
  MUX2_X1 U10452 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n9170), .S(n9546), .Z(
        P1_U3518) );
  MUX2_X1 U10453 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9171), .S(n9546), .Z(
        P1_U3517) );
  MUX2_X1 U10454 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9172), .S(n9546), .Z(
        P1_U3516) );
  MUX2_X1 U10455 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9173), .S(n9546), .Z(
        P1_U3515) );
  MUX2_X1 U10456 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9174), .S(n9546), .Z(
        P1_U3514) );
  MUX2_X1 U10457 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9175), .S(n9546), .Z(
        P1_U3513) );
  MUX2_X1 U10458 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9176), .S(n9546), .Z(
        P1_U3512) );
  MUX2_X1 U10459 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9177), .S(n9546), .Z(
        P1_U3511) );
  MUX2_X1 U10460 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9178), .S(n9546), .Z(
        P1_U3510) );
  MUX2_X1 U10461 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9179), .S(n9546), .Z(
        P1_U3509) );
  MUX2_X1 U10462 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9180), .S(n9546), .Z(
        P1_U3507) );
  MUX2_X1 U10463 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9181), .S(n9546), .Z(
        P1_U3504) );
  MUX2_X1 U10464 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n9182), .S(n9546), .Z(
        P1_U3501) );
  MUX2_X1 U10465 ( .A(n9183), .B(P1_D_REG_1__SCAN_IN), .S(n9512), .Z(P1_U3440)
         );
  MUX2_X1 U10466 ( .A(n9184), .B(P1_D_REG_0__SCAN_IN), .S(n9512), .Z(P1_U3439)
         );
  INV_X1 U10467 ( .A(n9185), .ZN(n9187) );
  NOR4_X1 U10468 ( .A1(n9187), .A2(P1_IR_REG_30__SCAN_IN), .A3(n5278), .A4(
        P1_U3086), .ZN(n9188) );
  AOI21_X1 U10469 ( .B1(n9189), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9188), .ZN(
        n9190) );
  OAI21_X1 U10470 ( .B1(n9191), .B2(n9193), .A(n9190), .ZN(P1_U3324) );
  OAI222_X1 U10471 ( .A1(n9195), .A2(n9194), .B1(n9193), .B2(n9192), .C1(n5282), .C2(P1_U3086), .ZN(P1_U3326) );
  MUX2_X1 U10472 ( .A(n9196), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  OAI21_X1 U10473 ( .B1(n9199), .B2(n9198), .A(n9197), .ZN(n9201) );
  AOI22_X1 U10474 ( .A1(n9201), .A2(n9730), .B1(n9200), .B2(
        P2_ADDR_REG_18__SCAN_IN), .ZN(n9217) );
  INV_X1 U10475 ( .A(n9202), .ZN(n9209) );
  NAND3_X1 U10476 ( .A1(n9203), .A2(n9202), .A3(P2_U3893), .ZN(n9205) );
  NAND3_X1 U10477 ( .A1(n9205), .A2(n9204), .A3(n9721), .ZN(n9208) );
  NAND2_X1 U10478 ( .A1(n4472), .A2(n9206), .ZN(n9207) );
  OAI211_X1 U10479 ( .C1(n9210), .C2(n9209), .A(n9208), .B(n9207), .ZN(n9216)
         );
  NAND2_X1 U10480 ( .A1(P2_REG3_REG_18__SCAN_IN), .A2(P2_U3151), .ZN(n9215) );
  AOI21_X1 U10481 ( .B1(n4397), .B2(n9212), .A(n9211), .ZN(n9213) );
  OR2_X1 U10482 ( .A1(n9213), .A2(n9736), .ZN(n9214) );
  NAND4_X1 U10483 ( .A1(n9217), .A2(n9216), .A3(n9215), .A4(n9214), .ZN(
        P2_U3200) );
  INV_X1 U10484 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n9232) );
  AOI21_X1 U10485 ( .B1(n9220), .B2(n9219), .A(n9218), .ZN(n9221) );
  NAND2_X1 U10486 ( .A1(n9446), .A2(n9221), .ZN(n9227) );
  AOI21_X1 U10487 ( .B1(n9224), .B2(n9223), .A(n9222), .ZN(n9225) );
  NAND2_X1 U10488 ( .A1(n9454), .A2(n9225), .ZN(n9226) );
  OAI211_X1 U10489 ( .C1(n9460), .C2(n9228), .A(n9227), .B(n9226), .ZN(n9229)
         );
  INV_X1 U10490 ( .A(n9229), .ZN(n9231) );
  OAI211_X1 U10491 ( .C1(n9466), .C2(n9232), .A(n9231), .B(n9230), .ZN(
        P1_U3253) );
  INV_X1 U10492 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n9247) );
  AOI21_X1 U10493 ( .B1(n9235), .B2(n9234), .A(n9233), .ZN(n9236) );
  NAND2_X1 U10494 ( .A1(n9446), .A2(n9236), .ZN(n9242) );
  AOI21_X1 U10495 ( .B1(n9239), .B2(n9238), .A(n9237), .ZN(n9240) );
  NAND2_X1 U10496 ( .A1(n9454), .A2(n9240), .ZN(n9241) );
  OAI211_X1 U10497 ( .C1(n9460), .C2(n9243), .A(n9242), .B(n9241), .ZN(n9244)
         );
  INV_X1 U10498 ( .A(n9244), .ZN(n9246) );
  OAI211_X1 U10499 ( .C1(n9466), .C2(n9247), .A(n9246), .B(n9245), .ZN(
        P1_U3250) );
  INV_X1 U10500 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n9262) );
  AOI21_X1 U10501 ( .B1(n9250), .B2(n9249), .A(n9248), .ZN(n9251) );
  NAND2_X1 U10502 ( .A1(n9446), .A2(n9251), .ZN(n9257) );
  AOI21_X1 U10503 ( .B1(n9254), .B2(n9253), .A(n9252), .ZN(n9255) );
  NAND2_X1 U10504 ( .A1(n9454), .A2(n9255), .ZN(n9256) );
  OAI211_X1 U10505 ( .C1(n9460), .C2(n9258), .A(n9257), .B(n9256), .ZN(n9259)
         );
  INV_X1 U10506 ( .A(n9259), .ZN(n9261) );
  OAI211_X1 U10507 ( .C1(n9466), .C2(n9262), .A(n9261), .B(n9260), .ZN(
        P1_U3251) );
  INV_X1 U10508 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n9277) );
  OAI21_X1 U10509 ( .B1(n9265), .B2(n9264), .A(n9263), .ZN(n9266) );
  NAND2_X1 U10510 ( .A1(n9446), .A2(n9266), .ZN(n9272) );
  OAI21_X1 U10511 ( .B1(n9269), .B2(n9268), .A(n9267), .ZN(n9270) );
  NAND2_X1 U10512 ( .A1(n9454), .A2(n9270), .ZN(n9271) );
  OAI211_X1 U10513 ( .C1(n9460), .C2(n9273), .A(n9272), .B(n9271), .ZN(n9274)
         );
  INV_X1 U10514 ( .A(n9274), .ZN(n9276) );
  OAI211_X1 U10515 ( .C1(n9466), .C2(n9277), .A(n9276), .B(n9275), .ZN(
        P1_U3252) );
  INV_X1 U10516 ( .A(n9280), .ZN(n9278) );
  AOI21_X1 U10517 ( .B1(n9279), .B2(n9835), .A(n9278), .ZN(n9288) );
  AOI22_X1 U10518 ( .A1(n9854), .A2(n9288), .B1(n7758), .B2(n9852), .ZN(
        P2_U3490) );
  OAI21_X1 U10519 ( .B1(n9281), .B2(n9807), .A(n9280), .ZN(n9290) );
  OAI22_X1 U10520 ( .A1(n9852), .A2(n9290), .B1(P2_REG1_REG_30__SCAN_IN), .B2(
        n9854), .ZN(n9282) );
  INV_X1 U10521 ( .A(n9282), .ZN(P2_U3489) );
  AND2_X1 U10522 ( .A1(n9283), .A2(n9831), .ZN(n9285) );
  AOI211_X1 U10523 ( .C1(n9835), .C2(n9286), .A(n9285), .B(n9284), .ZN(n9292)
         );
  INV_X1 U10524 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n9287) );
  AOI22_X1 U10525 ( .A1(n9854), .A2(n9292), .B1(n9287), .B2(n9852), .ZN(
        P2_U3472) );
  INV_X1 U10526 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n9289) );
  AOI22_X1 U10527 ( .A1(n9838), .A2(n9289), .B1(n9288), .B2(n9836), .ZN(
        P2_U3458) );
  OAI22_X1 U10528 ( .A1(n9836), .A2(P2_REG0_REG_30__SCAN_IN), .B1(n9290), .B2(
        n9838), .ZN(n9291) );
  INV_X1 U10529 ( .A(n9291), .ZN(P2_U3457) );
  INV_X1 U10530 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n9293) );
  AOI22_X1 U10531 ( .A1(n9838), .A2(n9293), .B1(n9292), .B2(n9836), .ZN(
        P2_U3429) );
  OAI21_X1 U10532 ( .B1(n9295), .B2(n9613), .A(n9294), .ZN(n9296) );
  AOI211_X1 U10533 ( .C1(n9298), .C2(n9617), .A(n9297), .B(n9296), .ZN(n9300)
         );
  AOI22_X1 U10534 ( .A1(n9630), .A2(n9300), .B1(n9415), .B2(n9644), .ZN(
        P1_U3537) );
  INV_X1 U10535 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n9299) );
  AOI22_X1 U10536 ( .A1(n9546), .A2(n9300), .B1(n9299), .B2(n9618), .ZN(
        P1_U3498) );
  INV_X1 U10537 ( .A(P2_WR_REG_SCAN_IN), .ZN(n9931) );
  XOR2_X1 U10538 ( .A(n9931), .B(P1_WR_REG_SCAN_IN), .Z(U123) );
  INV_X1 U10539 ( .A(P2_RD_REG_SCAN_IN), .ZN(n10053) );
  XOR2_X1 U10540 ( .A(P1_RD_REG_SCAN_IN), .B(n10053), .Z(U126) );
  OAI21_X1 U10541 ( .B1(P1_REG1_REG_0__SCAN_IN), .B2(n9302), .A(n9301), .ZN(
        n9303) );
  XOR2_X1 U10542 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9303), .Z(n9306) );
  AOI22_X1 U10543 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(n9431), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n9304) );
  OAI21_X1 U10544 ( .B1(n9306), .B2(n9305), .A(n9304), .ZN(P1_U3243) );
  AOI21_X1 U10545 ( .B1(P1_ADDR_REG_4__SCAN_IN), .B2(n9431), .A(n9307), .ZN(
        n9321) );
  INV_X1 U10546 ( .A(n9308), .ZN(n9311) );
  AOI211_X1 U10547 ( .C1(n9311), .C2(n9310), .A(n9309), .B(n9413), .ZN(n9317)
         );
  INV_X1 U10548 ( .A(n9312), .ZN(n9315) );
  AOI211_X1 U10549 ( .C1(n9315), .C2(n9314), .A(n9313), .B(n9451), .ZN(n9316)
         );
  AOI211_X1 U10550 ( .C1(n9443), .C2(n9318), .A(n9317), .B(n9316), .ZN(n9320)
         );
  NAND3_X1 U10551 ( .A1(n9321), .A2(n9320), .A3(n9319), .ZN(P1_U3247) );
  INV_X1 U10552 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n9336) );
  AOI21_X1 U10553 ( .B1(n9324), .B2(n9323), .A(n9322), .ZN(n9325) );
  NAND2_X1 U10554 ( .A1(n9446), .A2(n9325), .ZN(n9331) );
  AOI21_X1 U10555 ( .B1(n9328), .B2(n9327), .A(n9326), .ZN(n9329) );
  NAND2_X1 U10556 ( .A1(n9454), .A2(n9329), .ZN(n9330) );
  OAI211_X1 U10557 ( .C1(n9460), .C2(n9332), .A(n9331), .B(n9330), .ZN(n9333)
         );
  INV_X1 U10558 ( .A(n9333), .ZN(n9335) );
  OAI211_X1 U10559 ( .C1(n9466), .C2(n9336), .A(n9335), .B(n9334), .ZN(
        P1_U3248) );
  INV_X1 U10560 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n9350) );
  AOI21_X1 U10561 ( .B1(n9338), .B2(n4395), .A(n9337), .ZN(n9339) );
  NAND2_X1 U10562 ( .A1(n9446), .A2(n9339), .ZN(n9345) );
  AOI21_X1 U10563 ( .B1(n9342), .B2(n9341), .A(n9340), .ZN(n9343) );
  NAND2_X1 U10564 ( .A1(n9454), .A2(n9343), .ZN(n9344) );
  OAI211_X1 U10565 ( .C1(n9460), .C2(n9346), .A(n9345), .B(n9344), .ZN(n9347)
         );
  INV_X1 U10566 ( .A(n9347), .ZN(n9349) );
  OAI211_X1 U10567 ( .C1(n9466), .C2(n9350), .A(n9349), .B(n9348), .ZN(
        P1_U3249) );
  INV_X1 U10568 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n9366) );
  INV_X1 U10569 ( .A(n9351), .ZN(n9362) );
  AOI21_X1 U10570 ( .B1(n9354), .B2(n9353), .A(n9352), .ZN(n9355) );
  NAND2_X1 U10571 ( .A1(n9446), .A2(n9355), .ZN(n9361) );
  AOI21_X1 U10572 ( .B1(n9358), .B2(n9357), .A(n9356), .ZN(n9359) );
  NAND2_X1 U10573 ( .A1(n9454), .A2(n9359), .ZN(n9360) );
  OAI211_X1 U10574 ( .C1(n9460), .C2(n9362), .A(n9361), .B(n9360), .ZN(n9363)
         );
  INV_X1 U10575 ( .A(n9363), .ZN(n9365) );
  OAI211_X1 U10576 ( .C1(n9466), .C2(n9366), .A(n9365), .B(n9364), .ZN(
        P1_U3254) );
  INV_X1 U10577 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n9381) );
  OAI21_X1 U10578 ( .B1(n9369), .B2(n9368), .A(n9367), .ZN(n9370) );
  NAND2_X1 U10579 ( .A1(n9446), .A2(n9370), .ZN(n9376) );
  OAI21_X1 U10580 ( .B1(n9373), .B2(n9372), .A(n9371), .ZN(n9374) );
  NAND2_X1 U10581 ( .A1(n9454), .A2(n9374), .ZN(n9375) );
  OAI211_X1 U10582 ( .C1(n9460), .C2(n9377), .A(n9376), .B(n9375), .ZN(n9378)
         );
  INV_X1 U10583 ( .A(n9378), .ZN(n9380) );
  OAI211_X1 U10584 ( .C1(n9466), .C2(n9381), .A(n9380), .B(n9379), .ZN(
        P1_U3255) );
  INV_X1 U10585 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n9396) );
  AOI21_X1 U10586 ( .B1(n9384), .B2(n9383), .A(n9382), .ZN(n9385) );
  NAND2_X1 U10587 ( .A1(n9446), .A2(n9385), .ZN(n9391) );
  AOI21_X1 U10588 ( .B1(n9388), .B2(n9387), .A(n9386), .ZN(n9389) );
  NAND2_X1 U10589 ( .A1(n9454), .A2(n9389), .ZN(n9390) );
  OAI211_X1 U10590 ( .C1(n9460), .C2(n9392), .A(n9391), .B(n9390), .ZN(n9393)
         );
  INV_X1 U10591 ( .A(n9393), .ZN(n9395) );
  OAI211_X1 U10592 ( .C1(n9466), .C2(n9396), .A(n9395), .B(n9394), .ZN(
        P1_U3256) );
  INV_X1 U10593 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n9412) );
  INV_X1 U10594 ( .A(n9397), .ZN(n9408) );
  AOI21_X1 U10595 ( .B1(n9400), .B2(n9399), .A(n9398), .ZN(n9401) );
  NAND2_X1 U10596 ( .A1(n9446), .A2(n9401), .ZN(n9407) );
  AOI21_X1 U10597 ( .B1(n9404), .B2(n9403), .A(n9402), .ZN(n9405) );
  NAND2_X1 U10598 ( .A1(n9454), .A2(n9405), .ZN(n9406) );
  OAI211_X1 U10599 ( .C1(n9460), .C2(n9408), .A(n9407), .B(n9406), .ZN(n9409)
         );
  INV_X1 U10600 ( .A(n9409), .ZN(n9411) );
  OAI211_X1 U10601 ( .C1(n9466), .C2(n9412), .A(n9411), .B(n9410), .ZN(
        P1_U3257) );
  INV_X1 U10602 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n9425) );
  AOI211_X1 U10603 ( .C1(n9416), .C2(n9415), .A(n9414), .B(n9413), .ZN(n9421)
         );
  AOI211_X1 U10604 ( .C1(n9419), .C2(n9418), .A(n9417), .B(n9451), .ZN(n9420)
         );
  AOI211_X1 U10605 ( .C1(n9443), .C2(n9422), .A(n9421), .B(n9420), .ZN(n9424)
         );
  OAI211_X1 U10606 ( .C1(n9466), .C2(n9425), .A(n9424), .B(n9423), .ZN(
        P1_U3258) );
  AOI211_X1 U10607 ( .C1(n9428), .C2(n9427), .A(n9426), .B(n9451), .ZN(n9429)
         );
  AOI211_X1 U10608 ( .C1(n9431), .C2(P1_ADDR_REG_16__SCAN_IN), .A(n9430), .B(
        n9429), .ZN(n9438) );
  OAI21_X1 U10609 ( .B1(n9434), .B2(n9433), .A(n9432), .ZN(n9436) );
  AOI22_X1 U10610 ( .A1(n9436), .A2(n9454), .B1(n9435), .B2(n9443), .ZN(n9437)
         );
  NAND2_X1 U10611 ( .A1(n9438), .A2(n9437), .ZN(P1_U3259) );
  INV_X1 U10612 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n9450) );
  XNOR2_X1 U10613 ( .A(n9440), .B(n9439), .ZN(n9447) );
  XNOR2_X1 U10614 ( .A(n9442), .B(n9441), .ZN(n9445) );
  AOI222_X1 U10615 ( .A1(n9447), .A2(n9446), .B1(n9454), .B2(n9445), .C1(n9444), .C2(n9443), .ZN(n9449) );
  OAI211_X1 U10616 ( .C1(n9466), .C2(n9450), .A(n9449), .B(n9448), .ZN(
        P1_U3260) );
  INV_X1 U10617 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n10097) );
  AOI21_X1 U10618 ( .B1(n9453), .B2(n9452), .A(n9451), .ZN(n9463) );
  OAI211_X1 U10619 ( .C1(n9457), .C2(n9456), .A(n9455), .B(n9454), .ZN(n9458)
         );
  OAI21_X1 U10620 ( .B1(n9460), .B2(n9459), .A(n9458), .ZN(n9461) );
  AOI21_X1 U10621 ( .B1(n9463), .B2(n9462), .A(n9461), .ZN(n9465) );
  OAI211_X1 U10622 ( .C1(n9466), .C2(n10097), .A(n9465), .B(n9464), .ZN(
        P1_U3261) );
  XOR2_X1 U10623 ( .A(n9467), .B(n9475), .Z(n9469) );
  AOI222_X1 U10624 ( .A1(n9493), .A2(n9469), .B1(n7068), .B2(n9489), .C1(n9468), .C2(n9490), .ZN(n9555) );
  AOI222_X1 U10625 ( .A1(n9473), .A2(n9472), .B1(P1_REG2_REG_6__SCAN_IN), .B2(
        n9485), .C1(n9471), .C2(n9470), .ZN(n9484) );
  XNOR2_X1 U10626 ( .A(n9475), .B(n9474), .ZN(n9558) );
  INV_X1 U10627 ( .A(n9476), .ZN(n9479) );
  INV_X1 U10628 ( .A(n9477), .ZN(n9478) );
  OAI211_X1 U10629 ( .C1(n9554), .C2(n9479), .A(n9478), .B(n9496), .ZN(n9553)
         );
  INV_X1 U10630 ( .A(n9553), .ZN(n9481) );
  AOI22_X1 U10631 ( .A1(n9558), .A2(n9482), .B1(n9481), .B2(n9480), .ZN(n9483)
         );
  OAI211_X1 U10632 ( .C1(n9485), .C2(n9555), .A(n9484), .B(n9483), .ZN(
        P1_U3287) );
  INV_X1 U10633 ( .A(n9488), .ZN(n9487) );
  XNOR2_X1 U10634 ( .A(n9486), .B(n9487), .ZN(n9530) );
  XOR2_X1 U10635 ( .A(n8666), .B(n9488), .Z(n9492) );
  AOI222_X1 U10636 ( .A1(n9493), .A2(n9492), .B1(n9491), .B2(n9490), .C1(n6898), .C2(n9489), .ZN(n9529) );
  NAND2_X1 U10637 ( .A1(n9494), .A2(n9527), .ZN(n9495) );
  AND3_X1 U10638 ( .A1(n9497), .A2(n9496), .A3(n9495), .ZN(n9526) );
  INV_X1 U10639 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n9498) );
  OAI22_X1 U10640 ( .A1(n9501), .A2(n9500), .B1(n9499), .B2(n9498), .ZN(n9502)
         );
  AOI21_X1 U10641 ( .B1(n9526), .B2(n4453), .A(n9502), .ZN(n9504) );
  OAI211_X1 U10642 ( .C1(n9505), .C2(n9530), .A(n9529), .B(n9504), .ZN(n9508)
         );
  INV_X1 U10643 ( .A(n9530), .ZN(n9507) );
  AOI22_X1 U10644 ( .A1(n9508), .A2(n9510), .B1(n9507), .B2(n9506), .ZN(n9509)
         );
  OAI21_X1 U10645 ( .B1(n9511), .B2(n9510), .A(n9509), .ZN(P1_U3291) );
  AND2_X1 U10646 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n9512), .ZN(P1_U3294) );
  AND2_X1 U10647 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n9512), .ZN(P1_U3295) );
  AND2_X1 U10648 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n9512), .ZN(P1_U3296) );
  AND2_X1 U10649 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n9512), .ZN(P1_U3297) );
  AND2_X1 U10650 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n9512), .ZN(P1_U3298) );
  AND2_X1 U10651 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n9512), .ZN(P1_U3299) );
  AND2_X1 U10652 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n9512), .ZN(P1_U3300) );
  AND2_X1 U10653 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9512), .ZN(P1_U3301) );
  AND2_X1 U10654 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n9512), .ZN(P1_U3302) );
  AND2_X1 U10655 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n9512), .ZN(P1_U3303) );
  AND2_X1 U10656 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n9512), .ZN(P1_U3304) );
  AND2_X1 U10657 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n9512), .ZN(P1_U3305) );
  AND2_X1 U10658 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n9512), .ZN(P1_U3306) );
  AND2_X1 U10659 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n9512), .ZN(P1_U3307) );
  AND2_X1 U10660 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n9512), .ZN(P1_U3308) );
  AND2_X1 U10661 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n9512), .ZN(P1_U3309) );
  AND2_X1 U10662 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n9512), .ZN(P1_U3310) );
  AND2_X1 U10663 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n9512), .ZN(P1_U3311) );
  AND2_X1 U10664 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n9512), .ZN(P1_U3312) );
  AND2_X1 U10665 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n9512), .ZN(P1_U3313) );
  AND2_X1 U10666 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n9512), .ZN(P1_U3314) );
  AND2_X1 U10667 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n9512), .ZN(P1_U3315) );
  AND2_X1 U10668 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n9512), .ZN(P1_U3316) );
  AND2_X1 U10669 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n9512), .ZN(P1_U3317) );
  AND2_X1 U10670 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n9512), .ZN(P1_U3318) );
  AND2_X1 U10671 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n9512), .ZN(P1_U3319) );
  AND2_X1 U10672 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n9512), .ZN(P1_U3320) );
  AND2_X1 U10673 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n9512), .ZN(P1_U3321) );
  AND2_X1 U10674 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n9512), .ZN(P1_U3322) );
  AND2_X1 U10675 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n9512), .ZN(P1_U3323) );
  INV_X1 U10676 ( .A(n9513), .ZN(n9520) );
  INV_X1 U10677 ( .A(n9514), .ZN(n9515) );
  AOI21_X1 U10678 ( .B1(n9538), .B2(n9516), .A(n9515), .ZN(n9517) );
  AOI211_X1 U10679 ( .C1(n9520), .C2(n9519), .A(n9518), .B(n9517), .ZN(n9621)
         );
  AOI22_X1 U10680 ( .A1(n9546), .A2(n9621), .B1(n5905), .B2(n9618), .ZN(
        P1_U3453) );
  AOI211_X1 U10681 ( .C1(n9565), .C2(n9524), .A(n9523), .B(n9522), .ZN(n9623)
         );
  INV_X1 U10682 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n9525) );
  AOI22_X1 U10683 ( .A1(n9546), .A2(n9623), .B1(n9525), .B2(n9618), .ZN(
        P1_U3456) );
  AOI21_X1 U10684 ( .B1(n9591), .B2(n9527), .A(n9526), .ZN(n9528) );
  OAI211_X1 U10685 ( .C1(n9538), .C2(n9530), .A(n9529), .B(n9528), .ZN(n9531)
         );
  INV_X1 U10686 ( .A(n9531), .ZN(n9625) );
  INV_X1 U10687 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n9532) );
  AOI22_X1 U10688 ( .A1(n9546), .A2(n9625), .B1(n9532), .B2(n9618), .ZN(
        P1_U3459) );
  AOI21_X1 U10689 ( .B1(n9591), .B2(n9534), .A(n9533), .ZN(n9535) );
  OAI211_X1 U10690 ( .C1(n9538), .C2(n9537), .A(n9536), .B(n9535), .ZN(n9539)
         );
  INV_X1 U10691 ( .A(n9539), .ZN(n9627) );
  AOI22_X1 U10692 ( .A1(n9546), .A2(n9627), .B1(n5950), .B2(n9618), .ZN(
        P1_U3462) );
  OAI21_X1 U10693 ( .B1(n9541), .B2(n9613), .A(n9540), .ZN(n9543) );
  AOI211_X1 U10694 ( .C1(n9617), .C2(n9544), .A(n9543), .B(n9542), .ZN(n9629)
         );
  INV_X1 U10695 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n9545) );
  AOI22_X1 U10696 ( .A1(n9546), .A2(n9629), .B1(n9545), .B2(n9618), .ZN(
        P1_U3465) );
  OAI21_X1 U10697 ( .B1(n9548), .B2(n9613), .A(n9547), .ZN(n9550) );
  AOI211_X1 U10698 ( .C1(n9617), .C2(n9551), .A(n9550), .B(n9549), .ZN(n9631)
         );
  INV_X1 U10699 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n9552) );
  AOI22_X1 U10700 ( .A1(n9546), .A2(n9631), .B1(n9552), .B2(n9618), .ZN(
        P1_U3468) );
  OAI21_X1 U10701 ( .B1(n9554), .B2(n9613), .A(n9553), .ZN(n9557) );
  INV_X1 U10702 ( .A(n9555), .ZN(n9556) );
  AOI211_X1 U10703 ( .C1(n9617), .C2(n9558), .A(n9557), .B(n9556), .ZN(n9633)
         );
  INV_X1 U10704 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n9559) );
  AOI22_X1 U10705 ( .A1(n9546), .A2(n9633), .B1(n9559), .B2(n9618), .ZN(
        P1_U3471) );
  OAI21_X1 U10706 ( .B1(n9561), .B2(n9613), .A(n9560), .ZN(n9563) );
  AOI211_X1 U10707 ( .C1(n9565), .C2(n9564), .A(n9563), .B(n9562), .ZN(n9634)
         );
  INV_X1 U10708 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n9566) );
  AOI22_X1 U10709 ( .A1(n9546), .A2(n9634), .B1(n9566), .B2(n9618), .ZN(
        P1_U3474) );
  OAI22_X1 U10710 ( .A1(n9569), .A2(n9568), .B1(n9567), .B2(n9613), .ZN(n9570)
         );
  AOI21_X1 U10711 ( .B1(n9571), .B2(n9617), .A(n9570), .ZN(n9572) );
  AND2_X1 U10712 ( .A1(n9573), .A2(n9572), .ZN(n9636) );
  INV_X1 U10713 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n9574) );
  AOI22_X1 U10714 ( .A1(n9546), .A2(n9636), .B1(n9574), .B2(n9618), .ZN(
        P1_U3477) );
  OAI21_X1 U10715 ( .B1(n9576), .B2(n9613), .A(n9575), .ZN(n9577) );
  AOI21_X1 U10716 ( .B1(n9578), .B2(n9617), .A(n9577), .ZN(n9579) );
  AND2_X1 U10717 ( .A1(n9580), .A2(n9579), .ZN(n9638) );
  INV_X1 U10718 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n9581) );
  AOI22_X1 U10719 ( .A1(n9546), .A2(n9638), .B1(n9581), .B2(n9618), .ZN(
        P1_U3480) );
  OAI211_X1 U10720 ( .C1(n9584), .C2(n9613), .A(n9583), .B(n9582), .ZN(n9585)
         );
  AOI21_X1 U10721 ( .B1(n9617), .B2(n9586), .A(n9585), .ZN(n9640) );
  INV_X1 U10722 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n9587) );
  AOI22_X1 U10723 ( .A1(n9546), .A2(n9640), .B1(n9587), .B2(n9618), .ZN(
        P1_U3483) );
  INV_X1 U10724 ( .A(n9594), .ZN(n9596) );
  AOI211_X1 U10725 ( .C1(n9591), .C2(n9590), .A(n9589), .B(n9588), .ZN(n9592)
         );
  OAI21_X1 U10726 ( .B1(n9594), .B2(n9593), .A(n9592), .ZN(n9595) );
  AOI21_X1 U10727 ( .B1(n9597), .B2(n9596), .A(n9595), .ZN(n9641) );
  INV_X1 U10728 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n9598) );
  AOI22_X1 U10729 ( .A1(n9546), .A2(n9641), .B1(n9598), .B2(n9618), .ZN(
        P1_U3486) );
  OAI211_X1 U10730 ( .C1(n9601), .C2(n9613), .A(n9600), .B(n9599), .ZN(n9602)
         );
  AOI21_X1 U10731 ( .B1(n9617), .B2(n9603), .A(n9602), .ZN(n9642) );
  INV_X1 U10732 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n9604) );
  AOI22_X1 U10733 ( .A1(n9546), .A2(n9642), .B1(n9604), .B2(n9618), .ZN(
        P1_U3489) );
  OAI211_X1 U10734 ( .C1(n9607), .C2(n9613), .A(n9606), .B(n9605), .ZN(n9608)
         );
  AOI21_X1 U10735 ( .B1(n9617), .B2(n9609), .A(n9608), .ZN(n9643) );
  INV_X1 U10736 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n9610) );
  AOI22_X1 U10737 ( .A1(n9546), .A2(n9643), .B1(n9610), .B2(n9618), .ZN(
        P1_U3492) );
  OAI211_X1 U10738 ( .C1(n9614), .C2(n9613), .A(n9612), .B(n9611), .ZN(n9615)
         );
  AOI21_X1 U10739 ( .B1(n9617), .B2(n9616), .A(n9615), .ZN(n9645) );
  INV_X1 U10740 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n9619) );
  AOI22_X1 U10741 ( .A1(n9546), .A2(n9645), .B1(n9619), .B2(n9618), .ZN(
        P1_U3495) );
  AOI22_X1 U10742 ( .A1(n9630), .A2(n9621), .B1(n9620), .B2(n9644), .ZN(
        P1_U3522) );
  AOI22_X1 U10743 ( .A1(n9630), .A2(n9623), .B1(n9622), .B2(n9644), .ZN(
        P1_U3523) );
  AOI22_X1 U10744 ( .A1(n9630), .A2(n9625), .B1(n9624), .B2(n9644), .ZN(
        P1_U3524) );
  AOI22_X1 U10745 ( .A1(n9630), .A2(n9627), .B1(n9626), .B2(n9644), .ZN(
        P1_U3525) );
  INV_X1 U10746 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n9628) );
  AOI22_X1 U10747 ( .A1(n9630), .A2(n9629), .B1(n9628), .B2(n9644), .ZN(
        P1_U3526) );
  AOI22_X1 U10748 ( .A1(n9630), .A2(n9631), .B1(n8795), .B2(n9644), .ZN(
        P1_U3527) );
  INV_X1 U10749 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n9632) );
  AOI22_X1 U10750 ( .A1(n9630), .A2(n9633), .B1(n9632), .B2(n9644), .ZN(
        P1_U3528) );
  AOI22_X1 U10751 ( .A1(n9630), .A2(n9634), .B1(n8797), .B2(n9644), .ZN(
        P1_U3529) );
  INV_X1 U10752 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n9635) );
  AOI22_X1 U10753 ( .A1(n9630), .A2(n9636), .B1(n9635), .B2(n9644), .ZN(
        P1_U3530) );
  INV_X1 U10754 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n9637) );
  AOI22_X1 U10755 ( .A1(n9630), .A2(n9638), .B1(n9637), .B2(n9644), .ZN(
        P1_U3531) );
  INV_X1 U10756 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n9639) );
  AOI22_X1 U10757 ( .A1(n9630), .A2(n9640), .B1(n9639), .B2(n9644), .ZN(
        P1_U3532) );
  AOI22_X1 U10758 ( .A1(n9630), .A2(n9641), .B1(n8801), .B2(n9644), .ZN(
        P1_U3533) );
  AOI22_X1 U10759 ( .A1(n9630), .A2(n9642), .B1(n8802), .B2(n9644), .ZN(
        P1_U3534) );
  AOI22_X1 U10760 ( .A1(n9630), .A2(n9643), .B1(n8786), .B2(n9644), .ZN(
        P1_U3535) );
  AOI22_X1 U10761 ( .A1(n9630), .A2(n9645), .B1(n8804), .B2(n9644), .ZN(
        P1_U3536) );
  INV_X1 U10762 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n9646) );
  OAI22_X1 U10763 ( .A1(n9647), .A2(n9721), .B1(n9720), .B2(n9646), .ZN(n9648)
         );
  INV_X1 U10764 ( .A(n9648), .ZN(n9663) );
  OAI21_X1 U10765 ( .B1(P2_REG1_REG_13__SCAN_IN), .B2(n9650), .A(n9649), .ZN(
        n9655) );
  OAI21_X1 U10766 ( .B1(n9653), .B2(n9652), .A(n9651), .ZN(n9654) );
  AOI22_X1 U10767 ( .A1(n9655), .A2(n9730), .B1(n9729), .B2(n9654), .ZN(n9662)
         );
  NAND2_X1 U10768 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(n9917), .ZN(n9661) );
  AOI21_X1 U10769 ( .B1(n9658), .B2(n9657), .A(n9656), .ZN(n9659) );
  OR2_X1 U10770 ( .A1(n9659), .A2(n9736), .ZN(n9660) );
  NAND4_X1 U10771 ( .A1(n9663), .A2(n9662), .A3(n9661), .A4(n9660), .ZN(
        P2_U3195) );
  INV_X1 U10772 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n9664) );
  OAI22_X1 U10773 ( .A1(n9665), .A2(n9721), .B1(n9720), .B2(n9664), .ZN(n9666)
         );
  INV_X1 U10774 ( .A(n9666), .ZN(n9682) );
  OAI21_X1 U10775 ( .B1(n9669), .B2(n9668), .A(n9667), .ZN(n9674) );
  OAI21_X1 U10776 ( .B1(n9672), .B2(n9671), .A(n9670), .ZN(n9673) );
  AOI22_X1 U10777 ( .A1(n9674), .A2(n9730), .B1(n9729), .B2(n9673), .ZN(n9681)
         );
  NAND2_X1 U10778 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(n9917), .ZN(n9680) );
  AOI21_X1 U10779 ( .B1(n9677), .B2(n9676), .A(n9675), .ZN(n9678) );
  OR2_X1 U10780 ( .A1(n9678), .A2(n9736), .ZN(n9679) );
  NAND4_X1 U10781 ( .A1(n9682), .A2(n9681), .A3(n9680), .A4(n9679), .ZN(
        P2_U3196) );
  INV_X1 U10782 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n9683) );
  OAI22_X1 U10783 ( .A1(n4759), .A2(n9721), .B1(n9720), .B2(n9683), .ZN(n9684)
         );
  INV_X1 U10784 ( .A(n9684), .ZN(n9699) );
  OAI21_X1 U10785 ( .B1(P2_REG1_REG_15__SCAN_IN), .B2(n9686), .A(n9685), .ZN(
        n9691) );
  OAI21_X1 U10786 ( .B1(n9689), .B2(n9688), .A(n9687), .ZN(n9690) );
  AOI22_X1 U10787 ( .A1(n9691), .A2(n9730), .B1(n9729), .B2(n9690), .ZN(n9698)
         );
  AOI21_X1 U10788 ( .B1(n9694), .B2(n9693), .A(n9692), .ZN(n9695) );
  OR2_X1 U10789 ( .A1(n9736), .A2(n9695), .ZN(n9696) );
  NAND4_X1 U10790 ( .A1(n9699), .A2(n9698), .A3(n9697), .A4(n9696), .ZN(
        P2_U3197) );
  INV_X1 U10791 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n9700) );
  OAI22_X1 U10792 ( .A1(n9701), .A2(n9721), .B1(n9720), .B2(n9700), .ZN(n9702)
         );
  INV_X1 U10793 ( .A(n9702), .ZN(n9718) );
  OAI21_X1 U10794 ( .B1(n9705), .B2(n9704), .A(n9703), .ZN(n9710) );
  OAI21_X1 U10795 ( .B1(n9708), .B2(n9707), .A(n9706), .ZN(n9709) );
  AOI22_X1 U10796 ( .A1(n9710), .A2(n9730), .B1(n9729), .B2(n9709), .ZN(n9717)
         );
  NAND2_X1 U10797 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(P2_U3151), .ZN(n9716) );
  AOI21_X1 U10798 ( .B1(n9713), .B2(n9712), .A(n9711), .ZN(n9714) );
  OR2_X1 U10799 ( .A1(n9714), .A2(n9736), .ZN(n9715) );
  NAND4_X1 U10800 ( .A1(n9718), .A2(n9717), .A3(n9716), .A4(n9715), .ZN(
        P2_U3198) );
  INV_X1 U10801 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n9719) );
  OAI22_X1 U10802 ( .A1(n8030), .A2(n9721), .B1(n9720), .B2(n9719), .ZN(n9722)
         );
  INV_X1 U10803 ( .A(n9722), .ZN(n9740) );
  OAI21_X1 U10804 ( .B1(P2_REG1_REG_17__SCAN_IN), .B2(n9724), .A(n9723), .ZN(
        n9731) );
  OAI21_X1 U10805 ( .B1(n9727), .B2(n9726), .A(n9725), .ZN(n9728) );
  AOI22_X1 U10806 ( .A1(n9731), .A2(n9730), .B1(n9729), .B2(n9728), .ZN(n9739)
         );
  NAND2_X1 U10807 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(n9917), .ZN(n9738) );
  AOI21_X1 U10808 ( .B1(n9734), .B2(n9733), .A(n9732), .ZN(n9735) );
  OR2_X1 U10809 ( .A1(n9736), .A2(n9735), .ZN(n9737) );
  NAND4_X1 U10810 ( .A1(n9740), .A2(n9739), .A3(n9738), .A4(n9737), .ZN(
        P2_U3199) );
  NAND2_X1 U10811 ( .A1(n9757), .A2(n9741), .ZN(n9743) );
  XNOR2_X1 U10812 ( .A(n9743), .B(n9742), .ZN(n9748) );
  AOI222_X1 U10813 ( .A1(n9765), .A2(n9748), .B1(n9747), .B2(n9746), .C1(n9745), .C2(n9744), .ZN(n9792) );
  INV_X1 U10814 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n9755) );
  XNOR2_X1 U10815 ( .A(n9749), .B(n9750), .ZN(n9790) );
  AOI222_X1 U10816 ( .A1(n9790), .A2(n9753), .B1(n9752), .B2(n9770), .C1(n9789), .C2(n9751), .ZN(n9754) );
  OAI221_X1 U10817 ( .B1(n9777), .B2(n9792), .C1(n9775), .C2(n9755), .A(n9754), 
        .ZN(P2_U3230) );
  XNOR2_X1 U10818 ( .A(n9756), .B(n9759), .ZN(n9784) );
  OAI21_X1 U10819 ( .B1(n9759), .B2(n9758), .A(n9757), .ZN(n9766) );
  OAI22_X1 U10820 ( .A1(n9763), .A2(n9762), .B1(n9761), .B2(n9760), .ZN(n9764)
         );
  AOI21_X1 U10821 ( .B1(n9766), .B2(n9765), .A(n9764), .ZN(n9767) );
  OAI21_X1 U10822 ( .B1(n9784), .B2(n9768), .A(n9767), .ZN(n9785) );
  NOR2_X1 U10823 ( .A1(n9769), .A2(n9807), .ZN(n9786) );
  AOI22_X1 U10824 ( .A1(n9786), .A2(n9771), .B1(P2_REG3_REG_2__SCAN_IN), .B2(
        n9770), .ZN(n9772) );
  OAI21_X1 U10825 ( .B1(n9784), .B2(n9773), .A(n9772), .ZN(n9774) );
  NOR2_X1 U10826 ( .A1(n9785), .A2(n9774), .ZN(n9776) );
  AOI22_X1 U10827 ( .A1(n9777), .A2(n4460), .B1(n9776), .B2(n9775), .ZN(
        P2_U3231) );
  INV_X1 U10828 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n9783) );
  INV_X1 U10829 ( .A(n9778), .ZN(n9782) );
  OAI22_X1 U10830 ( .A1(n9780), .A2(n9796), .B1(n9779), .B2(n9807), .ZN(n9781)
         );
  NOR2_X1 U10831 ( .A1(n9782), .A2(n9781), .ZN(n9839) );
  AOI22_X1 U10832 ( .A1(n9838), .A2(n9783), .B1(n9839), .B2(n9836), .ZN(
        P2_U3393) );
  INV_X1 U10833 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n9788) );
  INV_X1 U10834 ( .A(n9819), .ZN(n9805) );
  INV_X1 U10835 ( .A(n9784), .ZN(n9787) );
  AOI211_X1 U10836 ( .C1(n9805), .C2(n9787), .A(n9786), .B(n9785), .ZN(n9840)
         );
  AOI22_X1 U10837 ( .A1(n9838), .A2(n9788), .B1(n9840), .B2(n9836), .ZN(
        P2_U3396) );
  INV_X1 U10838 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n9793) );
  AOI22_X1 U10839 ( .A1(n9790), .A2(n9831), .B1(n9835), .B2(n9789), .ZN(n9791)
         );
  AND2_X1 U10840 ( .A1(n9792), .A2(n9791), .ZN(n9841) );
  AOI22_X1 U10841 ( .A1(n9838), .A2(n9793), .B1(n9841), .B2(n9836), .ZN(
        P2_U3399) );
  INV_X1 U10842 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n9800) );
  INV_X1 U10843 ( .A(n9794), .ZN(n9799) );
  OAI22_X1 U10844 ( .A1(n9797), .A2(n9796), .B1(n9795), .B2(n9807), .ZN(n9798)
         );
  NOR2_X1 U10845 ( .A1(n9799), .A2(n9798), .ZN(n9842) );
  AOI22_X1 U10846 ( .A1(n9838), .A2(n9800), .B1(n9842), .B2(n9836), .ZN(
        P2_U3402) );
  INV_X1 U10847 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n9806) );
  NOR2_X1 U10848 ( .A1(n9801), .A2(n9807), .ZN(n9803) );
  AOI211_X1 U10849 ( .C1(n9805), .C2(n9804), .A(n9803), .B(n9802), .ZN(n9844)
         );
  AOI22_X1 U10850 ( .A1(n9838), .A2(n9806), .B1(n9844), .B2(n9836), .ZN(
        P2_U3405) );
  INV_X1 U10851 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n9812) );
  OAI22_X1 U10852 ( .A1(n9809), .A2(n9819), .B1(n9808), .B2(n9807), .ZN(n9810)
         );
  NOR2_X1 U10853 ( .A1(n9811), .A2(n9810), .ZN(n9846) );
  AOI22_X1 U10854 ( .A1(n9838), .A2(n9812), .B1(n9846), .B2(n9836), .ZN(
        P2_U3411) );
  INV_X1 U10855 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n9818) );
  AND2_X1 U10856 ( .A1(n9813), .A2(n9831), .ZN(n9816) );
  AND2_X1 U10857 ( .A1(n9814), .A2(n9835), .ZN(n9815) );
  NOR3_X1 U10858 ( .A1(n9817), .A2(n9816), .A3(n9815), .ZN(n9848) );
  AOI22_X1 U10859 ( .A1(n9838), .A2(n9818), .B1(n9848), .B2(n9836), .ZN(
        P2_U3414) );
  INV_X1 U10860 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n9824) );
  NOR2_X1 U10861 ( .A1(n9820), .A2(n9819), .ZN(n9822) );
  AOI211_X1 U10862 ( .C1(n9835), .C2(n9823), .A(n9822), .B(n9821), .ZN(n9849)
         );
  AOI22_X1 U10863 ( .A1(n9838), .A2(n9824), .B1(n9849), .B2(n9836), .ZN(
        P2_U3417) );
  INV_X1 U10864 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n9829) );
  AOI22_X1 U10865 ( .A1(n9826), .A2(n9831), .B1(n9835), .B2(n9825), .ZN(n9827)
         );
  AND2_X1 U10866 ( .A1(n9828), .A2(n9827), .ZN(n9851) );
  AOI22_X1 U10867 ( .A1(n9838), .A2(n9829), .B1(n9851), .B2(n9836), .ZN(
        P2_U3423) );
  INV_X1 U10868 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n9837) );
  AND3_X1 U10869 ( .A1(n7349), .A2(n9831), .A3(n9830), .ZN(n9833) );
  AOI211_X1 U10870 ( .C1(n9835), .C2(n9834), .A(n9833), .B(n9832), .ZN(n9853)
         );
  AOI22_X1 U10871 ( .A1(n9838), .A2(n9837), .B1(n9853), .B2(n9836), .ZN(
        P2_U3426) );
  AOI22_X1 U10872 ( .A1(n9854), .A2(n9839), .B1(n6413), .B2(n9852), .ZN(
        P2_U3460) );
  AOI22_X1 U10873 ( .A1(n9854), .A2(n9840), .B1(n6527), .B2(n9852), .ZN(
        P2_U3461) );
  AOI22_X1 U10874 ( .A1(n9854), .A2(n9841), .B1(n6561), .B2(n9852), .ZN(
        P2_U3462) );
  AOI22_X1 U10875 ( .A1(n9854), .A2(n9842), .B1(n6651), .B2(n9852), .ZN(
        P2_U3463) );
  INV_X1 U10876 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n9843) );
  AOI22_X1 U10877 ( .A1(n9854), .A2(n9844), .B1(n9843), .B2(n9852), .ZN(
        P2_U3464) );
  INV_X1 U10878 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n9845) );
  AOI22_X1 U10879 ( .A1(n9854), .A2(n9846), .B1(n9845), .B2(n9852), .ZN(
        P2_U3466) );
  AOI22_X1 U10880 ( .A1(n9854), .A2(n9848), .B1(n9847), .B2(n9852), .ZN(
        P2_U3467) );
  AOI22_X1 U10881 ( .A1(n9854), .A2(n9849), .B1(n7288), .B2(n9852), .ZN(
        P2_U3468) );
  INV_X1 U10882 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n9850) );
  AOI22_X1 U10883 ( .A1(n9854), .A2(n9851), .B1(n9850), .B2(n9852), .ZN(
        P2_U3470) );
  AOI22_X1 U10884 ( .A1(n9854), .A2(n9853), .B1(n7419), .B2(n9852), .ZN(
        P2_U3471) );
  NAND3_X1 U10885 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(P1_ADDR_REG_0__SCAN_IN), 
        .A3(P2_ADDR_REG_0__SCAN_IN), .ZN(n9857) );
  AND2_X1 U10886 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .ZN(n9855) );
  NOR2_X1 U10887 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(n9855), .ZN(n9856) );
  INV_X1 U10888 ( .A(n9856), .ZN(n9873) );
  NAND2_X1 U10889 ( .A1(n9858), .A2(n9857), .ZN(n9872) );
  OAI222_X1 U10890 ( .A1(n9858), .A2(n9857), .B1(n9858), .B2(n9873), .C1(n9856), .C2(n9872), .ZN(ADD_1068_U5) );
  XOR2_X1 U10891 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1068_U46) );
  NOR2_X1 U10892 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n9859) );
  AOI21_X1 U10893 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n9859), .ZN(n9880) );
  NOR2_X1 U10894 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n9860) );
  AOI21_X1 U10895 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n9860), .ZN(n9883) );
  NOR2_X1 U10896 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n9861) );
  AOI21_X1 U10897 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n9861), .ZN(n9886) );
  NOR2_X1 U10898 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n9862) );
  AOI21_X1 U10899 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n9862), .ZN(n9889) );
  NOR2_X1 U10900 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n9863) );
  AOI21_X1 U10901 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n9863), .ZN(n9892) );
  NOR2_X1 U10902 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n9864) );
  AOI21_X1 U10903 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n9864), .ZN(n9895) );
  NOR2_X1 U10904 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n9865) );
  AOI21_X1 U10905 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n9865), .ZN(n9898) );
  NOR2_X1 U10906 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n9866) );
  AOI21_X1 U10907 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n9866), .ZN(n9901) );
  NOR2_X1 U10908 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n9867) );
  AOI21_X1 U10909 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(P2_ADDR_REG_9__SCAN_IN), 
        .A(n9867), .ZN(n10109) );
  NOR2_X1 U10910 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n9868) );
  AOI21_X1 U10911 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(P2_ADDR_REG_8__SCAN_IN), 
        .A(n9868), .ZN(n10112) );
  NOR2_X1 U10912 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n9869) );
  AOI21_X1 U10913 ( .B1(P1_ADDR_REG_7__SCAN_IN), .B2(P2_ADDR_REG_7__SCAN_IN), 
        .A(n9869), .ZN(n10115) );
  NOR2_X1 U10914 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n9870) );
  AOI21_X1 U10915 ( .B1(P1_ADDR_REG_6__SCAN_IN), .B2(P2_ADDR_REG_6__SCAN_IN), 
        .A(n9870), .ZN(n10118) );
  NOR2_X1 U10916 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(P2_ADDR_REG_5__SCAN_IN), 
        .ZN(n9871) );
  AOI21_X1 U10917 ( .B1(P2_ADDR_REG_5__SCAN_IN), .B2(P1_ADDR_REG_5__SCAN_IN), 
        .A(n9871), .ZN(n10121) );
  NAND2_X1 U10918 ( .A1(n9873), .A2(n9872), .ZN(n10106) );
  NAND2_X1 U10919 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n9874) );
  OAI21_X1 U10920 ( .B1(P1_ADDR_REG_2__SCAN_IN), .B2(P2_ADDR_REG_2__SCAN_IN), 
        .A(n9874), .ZN(n10105) );
  NOR2_X1 U10921 ( .A1(n10106), .A2(n10105), .ZN(n10104) );
  AOI21_X1 U10922 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(P1_ADDR_REG_2__SCAN_IN), 
        .A(n10104), .ZN(n10124) );
  NAND2_X1 U10923 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n9875) );
  OAI21_X1 U10924 ( .B1(P1_ADDR_REG_3__SCAN_IN), .B2(P2_ADDR_REG_3__SCAN_IN), 
        .A(n9875), .ZN(n10123) );
  NOR2_X1 U10925 ( .A1(n10124), .A2(n10123), .ZN(n10122) );
  AOI21_X1 U10926 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(P1_ADDR_REG_3__SCAN_IN), 
        .A(n10122), .ZN(n10127) );
  NOR2_X1 U10927 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n9876) );
  AOI21_X1 U10928 ( .B1(P2_ADDR_REG_4__SCAN_IN), .B2(P1_ADDR_REG_4__SCAN_IN), 
        .A(n9876), .ZN(n10126) );
  NAND2_X1 U10929 ( .A1(n10127), .A2(n10126), .ZN(n10125) );
  OAI21_X1 U10930 ( .B1(P1_ADDR_REG_4__SCAN_IN), .B2(P2_ADDR_REG_4__SCAN_IN), 
        .A(n10125), .ZN(n10120) );
  NAND2_X1 U10931 ( .A1(n10121), .A2(n10120), .ZN(n10119) );
  OAI21_X1 U10932 ( .B1(P1_ADDR_REG_5__SCAN_IN), .B2(P2_ADDR_REG_5__SCAN_IN), 
        .A(n10119), .ZN(n10117) );
  NAND2_X1 U10933 ( .A1(n10118), .A2(n10117), .ZN(n10116) );
  OAI21_X1 U10934 ( .B1(P2_ADDR_REG_6__SCAN_IN), .B2(P1_ADDR_REG_6__SCAN_IN), 
        .A(n10116), .ZN(n10114) );
  NAND2_X1 U10935 ( .A1(n10115), .A2(n10114), .ZN(n10113) );
  OAI21_X1 U10936 ( .B1(P2_ADDR_REG_7__SCAN_IN), .B2(P1_ADDR_REG_7__SCAN_IN), 
        .A(n10113), .ZN(n10111) );
  NAND2_X1 U10937 ( .A1(n10112), .A2(n10111), .ZN(n10110) );
  OAI21_X1 U10938 ( .B1(P2_ADDR_REG_8__SCAN_IN), .B2(P1_ADDR_REG_8__SCAN_IN), 
        .A(n10110), .ZN(n10108) );
  NAND2_X1 U10939 ( .A1(n10109), .A2(n10108), .ZN(n10107) );
  OAI21_X1 U10940 ( .B1(P2_ADDR_REG_9__SCAN_IN), .B2(P1_ADDR_REG_9__SCAN_IN), 
        .A(n10107), .ZN(n9900) );
  NAND2_X1 U10941 ( .A1(n9901), .A2(n9900), .ZN(n9899) );
  OAI21_X1 U10942 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n9899), .ZN(n9897) );
  NAND2_X1 U10943 ( .A1(n9898), .A2(n9897), .ZN(n9896) );
  OAI21_X1 U10944 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n9896), .ZN(n9894) );
  NAND2_X1 U10945 ( .A1(n9895), .A2(n9894), .ZN(n9893) );
  OAI21_X1 U10946 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n9893), .ZN(n9891) );
  NAND2_X1 U10947 ( .A1(n9892), .A2(n9891), .ZN(n9890) );
  OAI21_X1 U10948 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n9890), .ZN(n9888) );
  NAND2_X1 U10949 ( .A1(n9889), .A2(n9888), .ZN(n9887) );
  OAI21_X1 U10950 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n9887), .ZN(n9885) );
  NAND2_X1 U10951 ( .A1(n9886), .A2(n9885), .ZN(n9884) );
  OAI21_X1 U10952 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n9884), .ZN(n9882) );
  NAND2_X1 U10953 ( .A1(n9883), .A2(n9882), .ZN(n9881) );
  OAI21_X1 U10954 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n9881), .ZN(n9879) );
  NAND2_X1 U10955 ( .A1(n9880), .A2(n9879), .ZN(n9878) );
  OAI21_X1 U10956 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n9878), .ZN(n10096) );
  NAND2_X1 U10957 ( .A1(n10097), .A2(n10096), .ZN(n10098) );
  OAI21_X1 U10958 ( .B1(n10096), .B2(n10097), .A(n10098), .ZN(n9877) );
  XNOR2_X1 U10959 ( .A(n9877), .B(P2_ADDR_REG_18__SCAN_IN), .ZN(ADD_1068_U55)
         );
  OAI21_X1 U10960 ( .B1(n9880), .B2(n9879), .A(n9878), .ZN(ADD_1068_U56) );
  OAI21_X1 U10961 ( .B1(n9883), .B2(n9882), .A(n9881), .ZN(ADD_1068_U57) );
  OAI21_X1 U10962 ( .B1(n9886), .B2(n9885), .A(n9884), .ZN(ADD_1068_U58) );
  OAI21_X1 U10963 ( .B1(n9889), .B2(n9888), .A(n9887), .ZN(ADD_1068_U59) );
  OAI21_X1 U10964 ( .B1(n9892), .B2(n9891), .A(n9890), .ZN(ADD_1068_U60) );
  OAI21_X1 U10965 ( .B1(n9895), .B2(n9894), .A(n9893), .ZN(ADD_1068_U61) );
  OAI21_X1 U10966 ( .B1(n9898), .B2(n9897), .A(n9896), .ZN(ADD_1068_U62) );
  OAI21_X1 U10967 ( .B1(n9901), .B2(n9900), .A(n9899), .ZN(ADD_1068_U63) );
  INV_X1 U10968 ( .A(SI_30_), .ZN(n10027) );
  AOI22_X1 U10969 ( .A1(n5544), .A2(keyinput_g50), .B1(keyinput_g2), .B2(
        n10027), .ZN(n9902) );
  OAI221_X1 U10970 ( .B1(n5544), .B2(keyinput_g50), .C1(n10027), .C2(
        keyinput_g2), .A(n9902), .ZN(n9912) );
  XNOR2_X1 U10971 ( .A(n9903), .B(keyinput_g30), .ZN(n9911) );
  INV_X1 U10972 ( .A(SI_20_), .ZN(n9904) );
  XNOR2_X1 U10973 ( .A(keyinput_g12), .B(n9904), .ZN(n9910) );
  XNOR2_X1 U10974 ( .A(SI_1_), .B(keyinput_g31), .ZN(n9908) );
  XNOR2_X1 U10975 ( .A(SI_14_), .B(keyinput_g18), .ZN(n9907) );
  XNOR2_X1 U10976 ( .A(SI_4_), .B(keyinput_g28), .ZN(n9906) );
  XNOR2_X1 U10977 ( .A(SI_29_), .B(keyinput_g3), .ZN(n9905) );
  NAND4_X1 U10978 ( .A1(n9908), .A2(n9907), .A3(n9906), .A4(n9905), .ZN(n9909)
         );
  NOR4_X1 U10979 ( .A1(n9912), .A2(n9911), .A3(n9910), .A4(n9909), .ZN(n9953)
         );
  INV_X1 U10980 ( .A(SI_12_), .ZN(n10049) );
  AOI22_X1 U10981 ( .A1(n10049), .A2(keyinput_g20), .B1(n10019), .B2(
        keyinput_g45), .ZN(n9913) );
  OAI221_X1 U10982 ( .B1(n10049), .B2(keyinput_g20), .C1(n10019), .C2(
        keyinput_g45), .A(n9913), .ZN(n9924) );
  AOI22_X1 U10983 ( .A1(SI_31_), .A2(keyinput_g1), .B1(P2_REG3_REG_20__SCAN_IN), .B2(keyinput_g55), .ZN(n9914) );
  OAI221_X1 U10984 ( .B1(SI_31_), .B2(keyinput_g1), .C1(
        P2_REG3_REG_20__SCAN_IN), .C2(keyinput_g55), .A(n9914), .ZN(n9923) );
  INV_X1 U10985 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n9916) );
  AOI22_X1 U10986 ( .A1(P2_U3151), .A2(keyinput_g34), .B1(n9916), .B2(
        keyinput_g38), .ZN(n9915) );
  OAI221_X1 U10987 ( .B1(n9917), .B2(keyinput_g34), .C1(n9916), .C2(
        keyinput_g38), .A(n9915), .ZN(n9922) );
  INV_X1 U10988 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n9919) );
  AOI22_X1 U10989 ( .A1(n9920), .A2(keyinput_g58), .B1(n9919), .B2(
        keyinput_g36), .ZN(n9918) );
  OAI221_X1 U10990 ( .B1(n9920), .B2(keyinput_g58), .C1(n9919), .C2(
        keyinput_g36), .A(n9918), .ZN(n9921) );
  NOR4_X1 U10991 ( .A1(n9924), .A2(n9923), .A3(n9922), .A4(n9921), .ZN(n9952)
         );
  AOI22_X1 U10992 ( .A1(n10058), .A2(keyinput_g49), .B1(keyinput_g15), .B2(
        n9926), .ZN(n9925) );
  OAI221_X1 U10993 ( .B1(n10058), .B2(keyinput_g49), .C1(n9926), .C2(
        keyinput_g15), .A(n9925), .ZN(n9936) );
  INV_X1 U10994 ( .A(SI_6_), .ZN(n10035) );
  AOI22_X1 U10995 ( .A1(n10035), .A2(keyinput_g26), .B1(n10042), .B2(
        keyinput_g35), .ZN(n9927) );
  OAI221_X1 U10996 ( .B1(n10035), .B2(keyinput_g26), .C1(n10042), .C2(
        keyinput_g35), .A(n9927), .ZN(n9935) );
  AOI22_X1 U10997 ( .A1(n9752), .A2(keyinput_g40), .B1(n9929), .B2(
        keyinput_g52), .ZN(n9928) );
  OAI221_X1 U10998 ( .B1(n9752), .B2(keyinput_g40), .C1(n9929), .C2(
        keyinput_g52), .A(n9928), .ZN(n9934) );
  AOI22_X1 U10999 ( .A1(n9932), .A2(keyinput_g21), .B1(keyinput_g0), .B2(n9931), .ZN(n9930) );
  OAI221_X1 U11000 ( .B1(n9932), .B2(keyinput_g21), .C1(n9931), .C2(
        keyinput_g0), .A(n9930), .ZN(n9933) );
  NOR4_X1 U11001 ( .A1(n9936), .A2(n9935), .A3(n9934), .A4(n9933), .ZN(n9951)
         );
  AOI22_X1 U11002 ( .A1(n10053), .A2(keyinput_g33), .B1(keyinput_g8), .B2(
        n9938), .ZN(n9937) );
  OAI221_X1 U11003 ( .B1(n10053), .B2(keyinput_g33), .C1(n9938), .C2(
        keyinput_g8), .A(n9937), .ZN(n9949) );
  AOI22_X1 U11004 ( .A1(n9940), .A2(keyinput_g43), .B1(n5336), .B2(
        keyinput_g53), .ZN(n9939) );
  OAI221_X1 U11005 ( .B1(n9940), .B2(keyinput_g43), .C1(n5336), .C2(
        keyinput_g53), .A(n9939), .ZN(n9948) );
  AOI22_X1 U11006 ( .A1(n10066), .A2(keyinput_g48), .B1(n9942), .B2(
        keyinput_g62), .ZN(n9941) );
  OAI221_X1 U11007 ( .B1(n10066), .B2(keyinput_g48), .C1(n9942), .C2(
        keyinput_g62), .A(n9941), .ZN(n9947) );
  AOI22_X1 U11008 ( .A1(n9945), .A2(keyinput_g6), .B1(keyinput_g7), .B2(n9944), 
        .ZN(n9943) );
  OAI221_X1 U11009 ( .B1(n9945), .B2(keyinput_g6), .C1(n9944), .C2(keyinput_g7), .A(n9943), .ZN(n9946) );
  NOR4_X1 U11010 ( .A1(n9949), .A2(n9948), .A3(n9947), .A4(n9946), .ZN(n9950)
         );
  AND4_X1 U11011 ( .A1(n9953), .A2(n9952), .A3(n9951), .A4(n9950), .ZN(n10095)
         );
  OAI22_X1 U11012 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(keyinput_g46), .B1(
        keyinput_g23), .B2(SI_9_), .ZN(n9954) );
  AOI221_X1 U11013 ( .B1(P2_REG3_REG_12__SCAN_IN), .B2(keyinput_g46), .C1(
        SI_9_), .C2(keyinput_g23), .A(n9954), .ZN(n9961) );
  OAI22_X1 U11014 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(keyinput_g37), .B1(SI_3_), .B2(keyinput_g29), .ZN(n9955) );
  AOI221_X1 U11015 ( .B1(P2_REG3_REG_14__SCAN_IN), .B2(keyinput_g37), .C1(
        keyinput_g29), .C2(SI_3_), .A(n9955), .ZN(n9960) );
  OAI22_X1 U11016 ( .A1(P2_REG3_REG_22__SCAN_IN), .A2(keyinput_g57), .B1(
        P2_REG3_REG_19__SCAN_IN), .B2(keyinput_g41), .ZN(n9956) );
  AOI221_X1 U11017 ( .B1(P2_REG3_REG_22__SCAN_IN), .B2(keyinput_g57), .C1(
        keyinput_g41), .C2(P2_REG3_REG_19__SCAN_IN), .A(n9956), .ZN(n9959) );
  OAI22_X1 U11018 ( .A1(SI_13_), .A2(keyinput_g19), .B1(SI_10_), .B2(
        keyinput_g22), .ZN(n9957) );
  AOI221_X1 U11019 ( .B1(SI_13_), .B2(keyinput_g19), .C1(keyinput_g22), .C2(
        SI_10_), .A(n9957), .ZN(n9958) );
  NAND4_X1 U11020 ( .A1(n9961), .A2(n9960), .A3(n9959), .A4(n9958), .ZN(n9988)
         );
  OAI22_X1 U11021 ( .A1(SI_21_), .A2(keyinput_g11), .B1(SI_15_), .B2(
        keyinput_g17), .ZN(n9962) );
  AOI221_X1 U11022 ( .B1(SI_21_), .B2(keyinput_g11), .C1(keyinput_g17), .C2(
        SI_15_), .A(n9962), .ZN(n9968) );
  OAI22_X1 U11023 ( .A1(SI_23_), .A2(keyinput_g9), .B1(SI_22_), .B2(
        keyinput_g10), .ZN(n9963) );
  AOI221_X1 U11024 ( .B1(SI_23_), .B2(keyinput_g9), .C1(keyinput_g10), .C2(
        SI_22_), .A(n9963), .ZN(n9967) );
  OAI22_X1 U11025 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(keyinput_g61), .B1(
        keyinput_g5), .B2(SI_27_), .ZN(n9964) );
  AOI221_X1 U11026 ( .B1(P2_REG3_REG_6__SCAN_IN), .B2(keyinput_g61), .C1(
        SI_27_), .C2(keyinput_g5), .A(n9964), .ZN(n9966) );
  XNOR2_X1 U11027 ( .A(P2_REG3_REG_28__SCAN_IN), .B(keyinput_g42), .ZN(n9965)
         );
  NAND4_X1 U11028 ( .A1(n9968), .A2(n9967), .A3(n9966), .A4(n9965), .ZN(n9987)
         );
  OAI22_X1 U11029 ( .A1(SI_19_), .A2(keyinput_g13), .B1(P2_REG3_REG_1__SCAN_IN), .B2(keyinput_g44), .ZN(n9969) );
  AOI221_X1 U11030 ( .B1(SI_19_), .B2(keyinput_g13), .C1(keyinput_g44), .C2(
        P2_REG3_REG_1__SCAN_IN), .A(n9969), .ZN(n9976) );
  OAI22_X1 U11031 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(keyinput_g56), .B1(
        keyinput_g4), .B2(SI_28_), .ZN(n9970) );
  AOI221_X1 U11032 ( .B1(P2_REG3_REG_13__SCAN_IN), .B2(keyinput_g56), .C1(
        SI_28_), .C2(keyinput_g4), .A(n9970), .ZN(n9975) );
  OAI22_X1 U11033 ( .A1(P2_REG3_REG_24__SCAN_IN), .A2(keyinput_g51), .B1(SI_0_), .B2(keyinput_g32), .ZN(n9971) );
  AOI221_X1 U11034 ( .B1(P2_REG3_REG_24__SCAN_IN), .B2(keyinput_g51), .C1(
        keyinput_g32), .C2(SI_0_), .A(n9971), .ZN(n9974) );
  OAI22_X1 U11035 ( .A1(P2_REG3_REG_18__SCAN_IN), .A2(keyinput_g60), .B1(SI_7_), .B2(keyinput_g25), .ZN(n9972) );
  AOI221_X1 U11036 ( .B1(P2_REG3_REG_18__SCAN_IN), .B2(keyinput_g60), .C1(
        keyinput_g25), .C2(SI_7_), .A(n9972), .ZN(n9973) );
  NAND4_X1 U11037 ( .A1(n9976), .A2(n9975), .A3(n9974), .A4(n9973), .ZN(n9986)
         );
  OAI22_X1 U11038 ( .A1(P2_REG3_REG_15__SCAN_IN), .A2(keyinput_g63), .B1(
        P2_REG3_REG_10__SCAN_IN), .B2(keyinput_g39), .ZN(n9977) );
  AOI221_X1 U11039 ( .B1(P2_REG3_REG_15__SCAN_IN), .B2(keyinput_g63), .C1(
        keyinput_g39), .C2(P2_REG3_REG_10__SCAN_IN), .A(n9977), .ZN(n9984) );
  OAI22_X1 U11040 ( .A1(SI_16_), .A2(keyinput_g16), .B1(P2_REG3_REG_0__SCAN_IN), .B2(keyinput_g54), .ZN(n9978) );
  AOI221_X1 U11041 ( .B1(SI_16_), .B2(keyinput_g16), .C1(keyinput_g54), .C2(
        P2_REG3_REG_0__SCAN_IN), .A(n9978), .ZN(n9983) );
  OAI22_X1 U11042 ( .A1(SI_18_), .A2(keyinput_g14), .B1(keyinput_g27), .B2(
        SI_5_), .ZN(n9979) );
  AOI221_X1 U11043 ( .B1(SI_18_), .B2(keyinput_g14), .C1(SI_5_), .C2(
        keyinput_g27), .A(n9979), .ZN(n9982) );
  OAI22_X1 U11044 ( .A1(P2_REG3_REG_25__SCAN_IN), .A2(keyinput_g47), .B1(
        keyinput_g59), .B2(P2_REG3_REG_2__SCAN_IN), .ZN(n9980) );
  AOI221_X1 U11045 ( .B1(P2_REG3_REG_25__SCAN_IN), .B2(keyinput_g47), .C1(
        P2_REG3_REG_2__SCAN_IN), .C2(keyinput_g59), .A(n9980), .ZN(n9981) );
  NAND4_X1 U11046 ( .A1(n9984), .A2(n9983), .A3(n9982), .A4(n9981), .ZN(n9985)
         );
  NOR4_X1 U11047 ( .A1(n9988), .A2(n9987), .A3(n9986), .A4(n9985), .ZN(n10094)
         );
  AOI22_X1 U11048 ( .A1(SI_20_), .A2(keyinput_f12), .B1(
        P2_REG3_REG_23__SCAN_IN), .B2(keyinput_f38), .ZN(n9989) );
  OAI221_X1 U11049 ( .B1(SI_20_), .B2(keyinput_f12), .C1(
        P2_REG3_REG_23__SCAN_IN), .C2(keyinput_f38), .A(n9989), .ZN(n9996) );
  AOI22_X1 U11050 ( .A1(keyinput_f0), .A2(P2_WR_REG_SCAN_IN), .B1(
        P2_STATE_REG_SCAN_IN), .B2(keyinput_f34), .ZN(n9990) );
  OAI221_X1 U11051 ( .B1(keyinput_f0), .B2(P2_WR_REG_SCAN_IN), .C1(
        P2_STATE_REG_SCAN_IN), .C2(keyinput_f34), .A(n9990), .ZN(n9995) );
  AOI22_X1 U11052 ( .A1(SI_3_), .A2(keyinput_f29), .B1(P2_REG3_REG_24__SCAN_IN), .B2(keyinput_f51), .ZN(n9991) );
  OAI221_X1 U11053 ( .B1(SI_3_), .B2(keyinput_f29), .C1(
        P2_REG3_REG_24__SCAN_IN), .C2(keyinput_f51), .A(n9991), .ZN(n9994) );
  AOI22_X1 U11054 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(keyinput_f40), .B1(
        P2_REG3_REG_18__SCAN_IN), .B2(keyinput_f60), .ZN(n9992) );
  OAI221_X1 U11055 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(keyinput_f40), .C1(
        P2_REG3_REG_18__SCAN_IN), .C2(keyinput_f60), .A(n9992), .ZN(n9993) );
  NOR4_X1 U11056 ( .A1(n9996), .A2(n9995), .A3(n9994), .A4(n9993), .ZN(n10087)
         );
  AOI22_X1 U11057 ( .A1(SI_24_), .A2(keyinput_f8), .B1(P2_REG3_REG_17__SCAN_IN), .B2(keyinput_f50), .ZN(n9997) );
  OAI221_X1 U11058 ( .B1(SI_24_), .B2(keyinput_f8), .C1(
        P2_REG3_REG_17__SCAN_IN), .C2(keyinput_f50), .A(n9997), .ZN(n10004) );
  AOI22_X1 U11059 ( .A1(SI_19_), .A2(keyinput_f13), .B1(SI_23_), .B2(
        keyinput_f9), .ZN(n9998) );
  OAI221_X1 U11060 ( .B1(SI_19_), .B2(keyinput_f13), .C1(SI_23_), .C2(
        keyinput_f9), .A(n9998), .ZN(n10003) );
  AOI22_X1 U11061 ( .A1(P2_REG3_REG_0__SCAN_IN), .A2(keyinput_f54), .B1(SI_26_), .B2(keyinput_f6), .ZN(n9999) );
  OAI221_X1 U11062 ( .B1(P2_REG3_REG_0__SCAN_IN), .B2(keyinput_f54), .C1(
        SI_26_), .C2(keyinput_f6), .A(n9999), .ZN(n10002) );
  AOI22_X1 U11063 ( .A1(SI_25_), .A2(keyinput_f7), .B1(P2_REG3_REG_11__SCAN_IN), .B2(keyinput_f58), .ZN(n10000) );
  OAI221_X1 U11064 ( .B1(SI_25_), .B2(keyinput_f7), .C1(
        P2_REG3_REG_11__SCAN_IN), .C2(keyinput_f58), .A(n10000), .ZN(n10001)
         );
  NOR4_X1 U11065 ( .A1(n10004), .A2(n10003), .A3(n10002), .A4(n10001), .ZN(
        n10086) );
  AOI22_X1 U11066 ( .A1(SI_11_), .A2(keyinput_f21), .B1(
        P2_REG3_REG_27__SCAN_IN), .B2(keyinput_f36), .ZN(n10005) );
  OAI221_X1 U11067 ( .B1(SI_11_), .B2(keyinput_f21), .C1(
        P2_REG3_REG_27__SCAN_IN), .C2(keyinput_f36), .A(n10005), .ZN(n10084)
         );
  AOI22_X1 U11068 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(keyinput_f52), .B1(
        P2_REG3_REG_28__SCAN_IN), .B2(keyinput_f42), .ZN(n10006) );
  OAI221_X1 U11069 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(keyinput_f52), .C1(
        P2_REG3_REG_28__SCAN_IN), .C2(keyinput_f42), .A(n10006), .ZN(n10083)
         );
  AOI22_X1 U11070 ( .A1(SI_4_), .A2(keyinput_f28), .B1(P2_REG3_REG_9__SCAN_IN), 
        .B2(keyinput_f53), .ZN(n10007) );
  OAI221_X1 U11071 ( .B1(SI_4_), .B2(keyinput_f28), .C1(P2_REG3_REG_9__SCAN_IN), .C2(keyinput_f53), .A(n10007), .ZN(n10014) );
  AOI22_X1 U11072 ( .A1(P2_REG3_REG_1__SCAN_IN), .A2(keyinput_f44), .B1(
        P2_REG3_REG_22__SCAN_IN), .B2(keyinput_f57), .ZN(n10008) );
  OAI221_X1 U11073 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(keyinput_f44), .C1(
        P2_REG3_REG_22__SCAN_IN), .C2(keyinput_f57), .A(n10008), .ZN(n10013)
         );
  AOI22_X1 U11074 ( .A1(SI_22_), .A2(keyinput_f10), .B1(
        P2_REG3_REG_19__SCAN_IN), .B2(keyinput_f41), .ZN(n10009) );
  OAI221_X1 U11075 ( .B1(SI_22_), .B2(keyinput_f10), .C1(
        P2_REG3_REG_19__SCAN_IN), .C2(keyinput_f41), .A(n10009), .ZN(n10012)
         );
  AOI22_X1 U11076 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(keyinput_f61), .B1(
        P2_REG3_REG_26__SCAN_IN), .B2(keyinput_f62), .ZN(n10010) );
  OAI221_X1 U11077 ( .B1(P2_REG3_REG_6__SCAN_IN), .B2(keyinput_f61), .C1(
        P2_REG3_REG_26__SCAN_IN), .C2(keyinput_f62), .A(n10010), .ZN(n10011)
         );
  NOR4_X1 U11078 ( .A1(n10014), .A2(n10013), .A3(n10012), .A4(n10011), .ZN(
        n10018) );
  AOI22_X1 U11079 ( .A1(SI_5_), .A2(keyinput_f27), .B1(P2_REG3_REG_12__SCAN_IN), .B2(keyinput_f46), .ZN(n10015) );
  OAI221_X1 U11080 ( .B1(SI_5_), .B2(keyinput_f27), .C1(
        P2_REG3_REG_12__SCAN_IN), .C2(keyinput_f46), .A(n10015), .ZN(n10016)
         );
  AOI21_X1 U11081 ( .B1(keyinput_f45), .B2(n10019), .A(n10016), .ZN(n10017) );
  OAI211_X1 U11082 ( .C1(keyinput_f45), .C2(n10019), .A(n10018), .B(n10017), 
        .ZN(n10082) );
  AOI22_X1 U11083 ( .A1(n5157), .A2(keyinput_f17), .B1(n10021), .B2(
        keyinput_f55), .ZN(n10020) );
  OAI221_X1 U11084 ( .B1(n5157), .B2(keyinput_f17), .C1(n10021), .C2(
        keyinput_f55), .A(n10020), .ZN(n10033) );
  AOI22_X1 U11085 ( .A1(n5337), .A2(keyinput_f56), .B1(keyinput_f25), .B2(
        n10023), .ZN(n10022) );
  OAI221_X1 U11086 ( .B1(n5337), .B2(keyinput_f56), .C1(n10023), .C2(
        keyinput_f25), .A(n10022), .ZN(n10032) );
  AOI22_X1 U11087 ( .A1(n10026), .A2(keyinput_f18), .B1(n10025), .B2(
        keyinput_f5), .ZN(n10024) );
  OAI221_X1 U11088 ( .B1(n10026), .B2(keyinput_f18), .C1(n10025), .C2(
        keyinput_f5), .A(n10024), .ZN(n10031) );
  XOR2_X1 U11089 ( .A(n10027), .B(keyinput_f2), .Z(n10029) );
  XNOR2_X1 U11090 ( .A(P2_REG3_REG_2__SCAN_IN), .B(keyinput_f59), .ZN(n10028)
         );
  NAND2_X1 U11091 ( .A1(n10029), .A2(n10028), .ZN(n10030) );
  NOR4_X1 U11092 ( .A1(n10033), .A2(n10032), .A3(n10031), .A4(n10030), .ZN(
        n10080) );
  AOI22_X1 U11093 ( .A1(n10036), .A2(keyinput_f39), .B1(keyinput_f26), .B2(
        n10035), .ZN(n10034) );
  OAI221_X1 U11094 ( .B1(n10036), .B2(keyinput_f39), .C1(n10035), .C2(
        keyinput_f26), .A(n10034), .ZN(n10047) );
  INV_X1 U11095 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n10038) );
  AOI22_X1 U11096 ( .A1(SI_2_), .A2(keyinput_f30), .B1(n10038), .B2(
        keyinput_f63), .ZN(n10037) );
  OAI221_X1 U11097 ( .B1(SI_2_), .B2(keyinput_f30), .C1(n10038), .C2(
        keyinput_f63), .A(n10037), .ZN(n10046) );
  AOI22_X1 U11098 ( .A1(n4734), .A2(keyinput_f19), .B1(keyinput_f22), .B2(
        n10040), .ZN(n10039) );
  OAI221_X1 U11099 ( .B1(n4734), .B2(keyinput_f19), .C1(n10040), .C2(
        keyinput_f22), .A(n10039), .ZN(n10045) );
  AOI22_X1 U11100 ( .A1(n10043), .A2(keyinput_f3), .B1(n10042), .B2(
        keyinput_f35), .ZN(n10041) );
  OAI221_X1 U11101 ( .B1(n10043), .B2(keyinput_f3), .C1(n10042), .C2(
        keyinput_f35), .A(n10041), .ZN(n10044) );
  NOR4_X1 U11102 ( .A1(n10047), .A2(n10046), .A3(n10045), .A4(n10044), .ZN(
        n10079) );
  AOI22_X1 U11103 ( .A1(n10050), .A2(keyinput_f47), .B1(keyinput_f20), .B2(
        n10049), .ZN(n10048) );
  OAI221_X1 U11104 ( .B1(n10050), .B2(keyinput_f47), .C1(n10049), .C2(
        keyinput_f20), .A(n10048), .ZN(n10063) );
  AOI22_X1 U11105 ( .A1(n10053), .A2(keyinput_f33), .B1(keyinput_f14), .B2(
        n10052), .ZN(n10051) );
  OAI221_X1 U11106 ( .B1(n10053), .B2(keyinput_f33), .C1(n10052), .C2(
        keyinput_f14), .A(n10051), .ZN(n10062) );
  AOI22_X1 U11107 ( .A1(n10056), .A2(keyinput_f1), .B1(n10055), .B2(
        keyinput_f11), .ZN(n10054) );
  OAI221_X1 U11108 ( .B1(n10056), .B2(keyinput_f1), .C1(n10055), .C2(
        keyinput_f11), .A(n10054), .ZN(n10061) );
  INV_X1 U11109 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n10059) );
  AOI22_X1 U11110 ( .A1(n10059), .A2(keyinput_f37), .B1(keyinput_f49), .B2(
        n10058), .ZN(n10057) );
  OAI221_X1 U11111 ( .B1(n10059), .B2(keyinput_f37), .C1(n10058), .C2(
        keyinput_f49), .A(n10057), .ZN(n10060) );
  NOR4_X1 U11112 ( .A1(n10063), .A2(n10062), .A3(n10061), .A4(n10060), .ZN(
        n10078) );
  AOI22_X1 U11113 ( .A1(n10066), .A2(keyinput_f48), .B1(keyinput_f23), .B2(
        n10065), .ZN(n10064) );
  OAI221_X1 U11114 ( .B1(n10066), .B2(keyinput_f48), .C1(n10065), .C2(
        keyinput_f23), .A(n10064), .ZN(n10076) );
  AOI22_X1 U11115 ( .A1(n10069), .A2(keyinput_f16), .B1(n10068), .B2(
        keyinput_f4), .ZN(n10067) );
  OAI221_X1 U11116 ( .B1(n10069), .B2(keyinput_f16), .C1(n10068), .C2(
        keyinput_f4), .A(n10067), .ZN(n10075) );
  XNOR2_X1 U11117 ( .A(SI_17_), .B(keyinput_f15), .ZN(n10073) );
  XNOR2_X1 U11118 ( .A(SI_1_), .B(keyinput_f31), .ZN(n10072) );
  XNOR2_X1 U11119 ( .A(P2_REG3_REG_8__SCAN_IN), .B(keyinput_f43), .ZN(n10071)
         );
  XNOR2_X1 U11120 ( .A(SI_0_), .B(keyinput_f32), .ZN(n10070) );
  NAND4_X1 U11121 ( .A1(n10073), .A2(n10072), .A3(n10071), .A4(n10070), .ZN(
        n10074) );
  NOR3_X1 U11122 ( .A1(n10076), .A2(n10075), .A3(n10074), .ZN(n10077) );
  NAND4_X1 U11123 ( .A1(n10080), .A2(n10079), .A3(n10078), .A4(n10077), .ZN(
        n10081) );
  NOR4_X1 U11124 ( .A1(n10084), .A2(n10083), .A3(n10082), .A4(n10081), .ZN(
        n10085) );
  NAND3_X1 U11125 ( .A1(n10087), .A2(n10086), .A3(n10085), .ZN(n10089) );
  AOI21_X1 U11126 ( .B1(keyinput_f24), .B2(n10089), .A(keyinput_g24), .ZN(
        n10091) );
  INV_X1 U11127 ( .A(keyinput_f24), .ZN(n10088) );
  AOI21_X1 U11128 ( .B1(n10089), .B2(n10088), .A(n10092), .ZN(n10090) );
  AOI22_X1 U11129 ( .A1(n10092), .A2(n10091), .B1(keyinput_g24), .B2(n10090), 
        .ZN(n10093) );
  AOI21_X1 U11130 ( .B1(n10095), .B2(n10094), .A(n10093), .ZN(n10103) );
  NOR2_X1 U11131 ( .A1(n10097), .A2(n10096), .ZN(n10099) );
  OAI21_X1 U11132 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(n10099), .A(n10098), 
        .ZN(n10101) );
  XNOR2_X1 U11133 ( .A(P1_ADDR_REG_19__SCAN_IN), .B(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n10100) );
  XNOR2_X1 U11134 ( .A(n10101), .B(n10100), .ZN(n10102) );
  XNOR2_X1 U11135 ( .A(n10103), .B(n10102), .ZN(ADD_1068_U4) );
  AOI21_X1 U11136 ( .B1(n10106), .B2(n10105), .A(n10104), .ZN(ADD_1068_U54) );
  OAI21_X1 U11137 ( .B1(n10109), .B2(n10108), .A(n10107), .ZN(ADD_1068_U47) );
  OAI21_X1 U11138 ( .B1(n10112), .B2(n10111), .A(n10110), .ZN(ADD_1068_U48) );
  OAI21_X1 U11139 ( .B1(n10115), .B2(n10114), .A(n10113), .ZN(ADD_1068_U49) );
  OAI21_X1 U11140 ( .B1(n10118), .B2(n10117), .A(n10116), .ZN(ADD_1068_U50) );
  OAI21_X1 U11141 ( .B1(n10121), .B2(n10120), .A(n10119), .ZN(ADD_1068_U51) );
  AOI21_X1 U11142 ( .B1(n10124), .B2(n10123), .A(n10122), .ZN(ADD_1068_U53) );
  OAI21_X1 U11143 ( .B1(n10127), .B2(n10126), .A(n10125), .ZN(ADD_1068_U52) );
  CLKBUF_X1 U4866 ( .A(n5858), .Z(n4355) );
  CLKBUF_X1 U4867 ( .A(n5801), .Z(n4357) );
endmodule

