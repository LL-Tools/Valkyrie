

module b14_C_2inp_gates_syn ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, U3352, U3351, U3350, U3349, 
        U3348, U3347, U3346, U3345, U3344, U3343, U3342, U3341, U3340, U3339, 
        U3338, U3337, U3336, U3335, U3334, U3333, U3332, U3331, U3330, U3329, 
        U3328, U3327, U3326, U3325, U3324, U3323, U3322, U3321, U3458, U3459, 
        U3320, U3319, U3318, U3317, U3316, U3315, U3314, U3313, U3312, U3311, 
        U3310, U3309, U3308, U3307, U3306, U3305, U3304, U3303, U3302, U3301, 
        U3300, U3299, U3298, U3297, U3296, U3295, U3294, U3293, U3292, U3291, 
        U3467, U3469, U3471, U3473, U3475, U3477, U3479, U3481, U3483, U3485, 
        U3487, U3489, U3491, U3493, U3495, U3497, U3499, U3501, U3503, U3505, 
        U3506, U3507, U3508, U3509, U3510, U3511, U3512, U3513, U3514, U3515, 
        U3516, U3517, U3518, U3519, U3520, U3521, U3522, U3523, U3524, U3525, 
        U3526, U3527, U3528, U3529, U3530, U3531, U3532, U3533, U3534, U3535, 
        U3536, U3537, U3538, U3539, U3540, U3541, U3542, U3543, U3544, U3545, 
        U3546, U3547, U3548, U3549, U3290, U3289, U3288, U3287, U3286, U3285, 
        U3284, U3283, U3282, U3281, U3280, U3279, U3278, U3277, U3276, U3275, 
        U3274, U3273, U3272, U3271, U3270, U3269, U3268, U3267, U3266, U3265, 
        U3264, U3263, U3262, U3354, U3261, U3260, U3259, U3258, U3257, U3256, 
        U3255, U3254, U3253, U3252, U3251, U3250, U3249, U3248, U3247, U3246, 
        U3245, U3244, U3243, U3242, U3241, U3240, U3550, U3551, U3552, U3553, 
        U3554, U3555, U3556, U3557, U3558, U3559, U3560, U3561, U3562, U3563, 
        U3564, U3565, U3566, U3567, U3568, U3569, U3570, U3571, U3572, U3573, 
        U3574, U3575, U3576, U3577, U3578, U3579, U3580, U3581, U3239, U3238, 
        U3237, U3236, U3235, U3234, U3233, U3232, U3231, U3230, U3229, U3228, 
        U3227, U3226, U3225, U3224, U3223, U3222, U3221, U3220, U3219, U3218, 
        U3217, U3216, U3215, U3214, U3213, U3212, U3211, U3210, U3149, U3148, 
        U4043, keyinput127, keyinput126, keyinput125, keyinput124, keyinput123, 
        keyinput122, keyinput121, keyinput120, keyinput119, keyinput118, 
        keyinput117, keyinput116, keyinput115, keyinput114, keyinput113, 
        keyinput112, keyinput111, keyinput110, keyinput109, keyinput108, 
        keyinput107, keyinput106, keyinput105, keyinput104, keyinput103, 
        keyinput102, keyinput101, keyinput100, keyinput99, keyinput98, 
        keyinput97, keyinput96, keyinput95, keyinput94, keyinput93, keyinput92, 
        keyinput91, keyinput90, keyinput89, keyinput88, keyinput87, keyinput86, 
        keyinput85, keyinput84, keyinput83, keyinput82, keyinput81, keyinput80, 
        keyinput79, keyinput78, keyinput77, keyinput76, keyinput75, keyinput74, 
        keyinput73, keyinput72, keyinput71, keyinput70, keyinput69, keyinput68, 
        keyinput67, keyinput66, keyinput65, keyinput64, keyinput63, keyinput62, 
        keyinput61, keyinput60, keyinput59, keyinput58, keyinput57, keyinput56, 
        keyinput55, keyinput54, keyinput53, keyinput52, keyinput51, keyinput50, 
        keyinput49, keyinput48, keyinput47, keyinput46, keyinput45, keyinput44, 
        keyinput43, keyinput42, keyinput41, keyinput40, keyinput39, keyinput38, 
        keyinput37, keyinput36, keyinput35, keyinput34, keyinput33, keyinput32, 
        keyinput31, keyinput30, keyinput29, keyinput28, keyinput27, keyinput26, 
        keyinput25, keyinput24, keyinput23, keyinput22, keyinput21, keyinput20, 
        keyinput19, keyinput18, keyinput17, keyinput16, keyinput15, keyinput14, 
        keyinput13, keyinput12, keyinput11, keyinput10, keyinput9, keyinput8, 
        keyinput7, keyinput6, keyinput5, keyinput4, keyinput3, keyinput2, 
        keyinput1, keyinput0 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN, keyinput127, keyinput126, keyinput125,
         keyinput124, keyinput123, keyinput122, keyinput121, keyinput120,
         keyinput119, keyinput118, keyinput117, keyinput116, keyinput115,
         keyinput114, keyinput113, keyinput112, keyinput111, keyinput110,
         keyinput109, keyinput108, keyinput107, keyinput106, keyinput105,
         keyinput104, keyinput103, keyinput102, keyinput101, keyinput100,
         keyinput99, keyinput98, keyinput97, keyinput96, keyinput95,
         keyinput94, keyinput93, keyinput92, keyinput91, keyinput90,
         keyinput89, keyinput88, keyinput87, keyinput86, keyinput85,
         keyinput84, keyinput83, keyinput82, keyinput81, keyinput80,
         keyinput79, keyinput78, keyinput77, keyinput76, keyinput75,
         keyinput74, keyinput73, keyinput72, keyinput71, keyinput70,
         keyinput69, keyinput68, keyinput67, keyinput66, keyinput65,
         keyinput64, keyinput63, keyinput62, keyinput61, keyinput60,
         keyinput59, keyinput58, keyinput57, keyinput56, keyinput55,
         keyinput54, keyinput53, keyinput52, keyinput51, keyinput50,
         keyinput49, keyinput48, keyinput47, keyinput46, keyinput45,
         keyinput44, keyinput43, keyinput42, keyinput41, keyinput40,
         keyinput39, keyinput38, keyinput37, keyinput36, keyinput35,
         keyinput34, keyinput33, keyinput32, keyinput31, keyinput30,
         keyinput29, keyinput28, keyinput27, keyinput26, keyinput25,
         keyinput24, keyinput23, keyinput22, keyinput21, keyinput20,
         keyinput19, keyinput18, keyinput17, keyinput16, keyinput15,
         keyinput14, keyinput13, keyinput12, keyinput11, keyinput10, keyinput9,
         keyinput8, keyinput7, keyinput6, keyinput5, keyinput4, keyinput3,
         keyinput2, keyinput1, keyinput0;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155,
         n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165,
         n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175,
         n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185,
         n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195,
         n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205,
         n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215,
         n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225,
         n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235,
         n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245,
         n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255,
         n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265,
         n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275,
         n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285,
         n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295,
         n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305,
         n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315,
         n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325,
         n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335,
         n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345,
         n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355,
         n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365,
         n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375,
         n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385,
         n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395,
         n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405,
         n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415,
         n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425,
         n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435,
         n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445,
         n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455,
         n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465,
         n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475,
         n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485,
         n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495,
         n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505,
         n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515,
         n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525,
         n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535,
         n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545,
         n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555,
         n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565,
         n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575,
         n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585,
         n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595,
         n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605,
         n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615,
         n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625,
         n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635,
         n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645,
         n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655,
         n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665,
         n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675,
         n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685,
         n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695,
         n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705,
         n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715,
         n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725,
         n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735,
         n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745,
         n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755,
         n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765,
         n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775,
         n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785,
         n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795,
         n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805,
         n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815,
         n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825,
         n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835,
         n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845,
         n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855,
         n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865,
         n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875,
         n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885,
         n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895,
         n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905,
         n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915,
         n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925,
         n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935,
         n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945,
         n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955,
         n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965,
         n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975,
         n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985,
         n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995,
         n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005,
         n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015,
         n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025,
         n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035,
         n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045,
         n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055,
         n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065,
         n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075,
         n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085,
         n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095,
         n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105,
         n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115,
         n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125,
         n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135,
         n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145,
         n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155,
         n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3165, n3166,
         n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176,
         n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186,
         n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196,
         n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206,
         n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216,
         n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226,
         n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236,
         n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246,
         n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256,
         n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266,
         n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276,
         n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286,
         n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296,
         n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306,
         n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316,
         n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326,
         n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336,
         n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346,
         n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356,
         n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366,
         n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376,
         n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386,
         n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396,
         n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406,
         n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416,
         n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426,
         n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436,
         n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446,
         n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456,
         n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466,
         n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476,
         n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486,
         n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496,
         n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506,
         n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516,
         n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526,
         n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536,
         n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546,
         n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556,
         n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566,
         n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576,
         n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586,
         n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596,
         n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606,
         n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616,
         n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626,
         n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636,
         n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646,
         n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656,
         n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666,
         n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676,
         n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686,
         n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696,
         n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706,
         n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716,
         n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726,
         n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736,
         n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746,
         n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756,
         n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766,
         n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776,
         n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786,
         n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796,
         n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806,
         n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816,
         n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826,
         n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836,
         n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846,
         n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856,
         n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866,
         n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876,
         n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886,
         n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896,
         n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906,
         n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916,
         n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926,
         n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936,
         n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946,
         n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956,
         n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966,
         n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976,
         n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986,
         n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996,
         n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006,
         n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016,
         n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026,
         n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036,
         n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046,
         n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056,
         n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066,
         n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076,
         n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086,
         n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096,
         n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106,
         n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116,
         n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126,
         n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136,
         n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146,
         n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156,
         n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166,
         n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176,
         n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186,
         n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196,
         n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206,
         n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216,
         n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226,
         n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236,
         n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246,
         n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256,
         n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266,
         n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276,
         n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286,
         n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296,
         n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306,
         n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316,
         n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326,
         n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336,
         n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346,
         n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356,
         n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366,
         n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376,
         n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386,
         n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396,
         n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406,
         n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416,
         n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426,
         n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436,
         n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446,
         n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456,
         n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466,
         n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476,
         n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486,
         n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496,
         n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506,
         n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516,
         n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526,
         n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536,
         n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546,
         n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556,
         n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566,
         n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576,
         n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586,
         n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596,
         n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606,
         n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616,
         n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626,
         n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636,
         n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646,
         n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656,
         n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666,
         n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676,
         n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686,
         n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696,
         n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706,
         n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716,
         n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726,
         n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736,
         n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746,
         n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756,
         n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766,
         n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776,
         n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786,
         n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796,
         n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806,
         n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816,
         n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826,
         n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836,
         n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846,
         n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856,
         n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866,
         n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876,
         n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886,
         n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896,
         n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906,
         n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916,
         n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926,
         n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936,
         n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946,
         n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956,
         n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966,
         n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976,
         n4977, n4978, n4979, n4980, n4981, n4982, n4983;

  INV_X1 U2389 ( .A(n2446), .ZN(n2757) );
  AND2_X1 U2390 ( .A1(n2356), .A2(n3083), .ZN(n2426) );
  AND2_X1 U2391 ( .A1(n2351), .A2(n2350), .ZN(n3081) );
  NOR4_X1 U2392 ( .A1(n3952), .A2(n4241), .A3(n3951), .A4(n3950), .ZN(n3974)
         );
  INV_X1 U2393 ( .A(n2844), .ZN(n2858) );
  OAI21_X1 U2394 ( .B1(n3909), .B2(n3190), .A(n2416), .ZN(n3167) );
  INV_X1 U2396 ( .A(n2355), .ZN(n3083) );
  AOI21_X2 U2397 ( .B1(n4143), .B2(n4667), .A(n3043), .ZN(n3069) );
  NOR2_X2 U2398 ( .A1(n2699), .A2(n4926), .ZN(n2718) );
  OAI21_X2 U2399 ( .B1(n4317), .B2(n3892), .A(n3895), .ZN(n4273) );
  NAND2_X1 U2400 ( .A1(n4582), .A2(n4952), .ZN(n4581) );
  NAND2_X1 U2401 ( .A1(n4538), .A2(n4094), .ZN(n4551) );
  OR2_X1 U2402 ( .A1(n3277), .A2(n2226), .ZN(n2225) );
  NAND2_X2 U2403 ( .A1(n3353), .A2(n4332), .ZN(n4357) );
  OR2_X1 U2404 ( .A1(n2804), .A2(n3789), .ZN(n2819) );
  AND2_X1 U2405 ( .A1(n3278), .A2(n4493), .ZN(n2226) );
  AND2_X1 U2406 ( .A1(n2755), .A2(REG3_REG_22__SCAN_IN), .ZN(n2779) );
  XNOR2_X1 U2407 ( .A(n4086), .B(n4106), .ZN(n4088) );
  NAND2_X1 U2408 ( .A1(n2968), .A2(n3977), .ZN(n2965) );
  OAI21_X1 U2409 ( .B1(n3206), .B2(n2231), .A(n2230), .ZN(n3234) );
  NAND3_X1 U2410 ( .A1(n2395), .A2(n2394), .A3(n2393), .ZN(n3462) );
  AND2_X2 U2411 ( .A1(n2899), .A2(n2963), .ZN(n2844) );
  NAND2_X1 U2412 ( .A1(n4489), .A2(n4049), .ZN(n2963) );
  NAND2_X1 U2413 ( .A1(n2382), .A2(n2381), .ZN(n2927) );
  CLKBUF_X3 U2414 ( .A(n2409), .Z(n2906) );
  NAND2_X1 U2415 ( .A1(n2355), .A2(n3081), .ZN(n2446) );
  AOI21_X1 U2416 ( .B1(n3139), .B2(REG2_REG_3__SCAN_IN), .A(n2234), .ZN(n3140)
         );
  XNOR2_X1 U2417 ( .A(n2236), .B(n2235), .ZN(n3139) );
  MUX2_X1 U2418 ( .A(IR_REG_31__SCAN_IN), .B(n2349), .S(IR_REG_29__SCAN_IN), 
        .Z(n2351) );
  AND3_X1 U2419 ( .A1(n2340), .A2(n2474), .A3(n2216), .ZN(n2348) );
  AND2_X1 U2420 ( .A1(n2311), .A2(n2163), .ZN(n2217) );
  AND3_X1 U2421 ( .A1(n2511), .A2(n2253), .A3(n2252), .ZN(n2688) );
  NOR2_X1 U2422 ( .A1(IR_REG_21__SCAN_IN), .A2(IR_REG_24__SCAN_IN), .ZN(n2342)
         );
  NOR2_X1 U2423 ( .A1(IR_REG_18__SCAN_IN), .A2(IR_REG_20__SCAN_IN), .ZN(n2341)
         );
  NOR2_X1 U2424 ( .A1(n3234), .A2(n2326), .ZN(n3276) );
  NOR2_X1 U2425 ( .A1(n4570), .A2(n2233), .ZN(n4099) );
  AND2_X1 U2426 ( .A1(n4104), .A2(REG2_REG_15__SCAN_IN), .ZN(n2233) );
  INV_X1 U2427 ( .A(n2200), .ZN(n2198) );
  NOR2_X1 U2428 ( .A1(n2330), .A2(n2172), .ZN(n2203) );
  INV_X1 U2429 ( .A(n2210), .ZN(n2208) );
  NOR2_X1 U2430 ( .A1(n2955), .A2(n2173), .ZN(n2213) );
  AOI21_X1 U2431 ( .B1(n3233), .B2(REG2_REG_5__SCAN_IN), .A(n3230), .ZN(n3281)
         );
  AOI21_X1 U2432 ( .B1(n3634), .B2(n2190), .A(n2189), .ZN(n3721) );
  NOR2_X1 U2433 ( .A1(n2193), .A2(n2149), .ZN(n2190) );
  OAI21_X1 U2434 ( .B1(n2191), .B2(n2149), .A(n2168), .ZN(n2189) );
  AND2_X1 U2435 ( .A1(n2912), .A2(n2389), .ZN(n3368) );
  AND2_X1 U2436 ( .A1(n3096), .A2(n4488), .ZN(n4374) );
  NAND2_X1 U2437 ( .A1(n2350), .A2(IR_REG_31__SCAN_IN), .ZN(n2346) );
  AND2_X1 U2438 ( .A1(n2155), .A2(n2217), .ZN(n2216) );
  INV_X1 U2439 ( .A(n3669), .ZN(n2292) );
  NOR2_X1 U2440 ( .A1(IR_REG_10__SCAN_IN), .A2(IR_REG_11__SCAN_IN), .ZN(n2611)
         );
  NAND2_X1 U2441 ( .A1(n2299), .A2(n2298), .ZN(n2297) );
  INV_X1 U2442 ( .A(n3572), .ZN(n2298) );
  INV_X1 U2443 ( .A(n3571), .ZN(n2299) );
  AND2_X1 U2444 ( .A1(n3571), .A2(n3572), .ZN(n2295) );
  INV_X1 U2445 ( .A(n3081), .ZN(n2356) );
  INV_X1 U2446 ( .A(n3192), .ZN(n2223) );
  NAND2_X1 U2447 ( .A1(n2147), .A2(n2219), .ZN(n2218) );
  NOR2_X1 U2448 ( .A1(n3134), .A2(n3133), .ZN(n3136) );
  AND2_X1 U2449 ( .A1(n3132), .A2(n4495), .ZN(n3133) );
  NAND2_X1 U2450 ( .A1(n2224), .A2(n2147), .ZN(n3132) );
  NAND2_X1 U2451 ( .A1(n4507), .A2(n4111), .ZN(n4113) );
  INV_X1 U2452 ( .A(n4068), .ZN(n2930) );
  NAND2_X1 U2453 ( .A1(n2930), .A2(n3167), .ZN(n3981) );
  NAND2_X1 U2454 ( .A1(n3984), .A2(n3981), .ZN(n2970) );
  INV_X1 U2455 ( .A(n3704), .ZN(n3015) );
  AND2_X1 U2456 ( .A1(n3422), .A2(n3318), .ZN(n2314) );
  AND2_X1 U2457 ( .A1(n4489), .A2(n4057), .ZN(n3096) );
  NOR2_X1 U2458 ( .A1(IR_REG_25__SCAN_IN), .A2(IR_REG_26__SCAN_IN), .ZN(n2311)
         );
  NAND2_X1 U2459 ( .A1(n2361), .A2(n2305), .ZN(n2304) );
  NOR2_X1 U2460 ( .A1(IR_REG_18__SCAN_IN), .A2(IR_REG_21__SCAN_IN), .ZN(n2305)
         );
  INV_X1 U2461 ( .A(IR_REG_11__SCAN_IN), .ZN(n2578) );
  NOR2_X1 U2462 ( .A1(n3668), .A2(n2295), .ZN(n2294) );
  INV_X1 U2463 ( .A(n2278), .ZN(n2277) );
  OAI21_X1 U2464 ( .B1(n2279), .B2(n2165), .A(n3847), .ZN(n2278) );
  NAND2_X1 U2465 ( .A1(n2831), .A2(n2830), .ZN(n2301) );
  NAND2_X1 U2466 ( .A1(n2380), .A2(n3116), .ZN(n2382) );
  AND2_X1 U2467 ( .A1(n2697), .A2(n2696), .ZN(n3807) );
  AOI21_X1 U2468 ( .B1(n3754), .B2(n2793), .A(n2320), .ZN(n3816) );
  NOR2_X1 U2469 ( .A1(n2321), .A2(n2800), .ZN(n2801) );
  XNOR2_X1 U2470 ( .A(n2438), .B(n2844), .ZN(n2460) );
  NOR2_X1 U2471 ( .A1(n3475), .A2(n2265), .ZN(n2264) );
  INV_X1 U2472 ( .A(n2267), .ZN(n2265) );
  NAND2_X1 U2473 ( .A1(n3826), .A2(n3827), .ZN(n3825) );
  INV_X1 U2474 ( .A(n4344), .ZN(n3852) );
  AND2_X1 U2475 ( .A1(n2487), .A2(REG3_REG_6__SCAN_IN), .ZN(n2507) );
  OR2_X1 U2476 ( .A1(n2847), .A2(n2837), .ZN(n3749) );
  BUF_X1 U2478 ( .A(n3904), .Z(n2849) );
  NAND2_X1 U2479 ( .A1(n2368), .A2(n3089), .ZN(n3070) );
  NAND2_X1 U2480 ( .A1(n2238), .A2(n2237), .ZN(n2236) );
  NAND2_X1 U2481 ( .A1(n3186), .A2(n3185), .ZN(n2238) );
  XNOR2_X1 U2482 ( .A(n3136), .B(n3135), .ZN(n3206) );
  OAI21_X1 U2483 ( .B1(n2225), .B2(REG1_REG_7__SCAN_IN), .A(n4492), .ZN(n3336)
         );
  NAND2_X1 U2484 ( .A1(n4527), .A2(n4116), .ZN(n4118) );
  NAND2_X1 U2485 ( .A1(n4539), .A2(REG2_REG_12__SCAN_IN), .ZN(n4538) );
  NAND2_X1 U2486 ( .A1(n4555), .A2(n4120), .ZN(n4121) );
  NAND2_X1 U2487 ( .A1(n4575), .A2(n4123), .ZN(n4124) );
  NAND2_X1 U2488 ( .A1(n4581), .A2(n4100), .ZN(n4589) );
  NOR2_X1 U2489 ( .A1(n2250), .A2(n4602), .ZN(n4601) );
  NOR2_X1 U2490 ( .A1(n2819), .A2(n3861), .ZN(n2836) );
  AOI21_X1 U2491 ( .B1(n2203), .B2(n2201), .A(n2174), .ZN(n2200) );
  INV_X1 U2492 ( .A(n2961), .ZN(n2201) );
  AND2_X1 U2493 ( .A1(n4261), .A2(n4246), .ZN(n2959) );
  AOI21_X1 U2494 ( .B1(n2213), .B2(n2211), .A(n2176), .ZN(n2210) );
  INV_X1 U2495 ( .A(n2956), .ZN(n2211) );
  INV_X1 U2496 ( .A(n2213), .ZN(n2212) );
  AND2_X1 U2497 ( .A1(n4029), .A2(n4237), .ZN(n4276) );
  NAND2_X1 U2498 ( .A1(n2953), .A2(n4351), .ZN(n2954) );
  AND2_X1 U2499 ( .A1(n3582), .A2(n2169), .ZN(n2194) );
  AOI21_X1 U2500 ( .B1(n2188), .B2(n2186), .A(n2178), .ZN(n2185) );
  INV_X1 U2501 ( .A(n2188), .ZN(n2187) );
  OR2_X1 U2502 ( .A1(n2328), .A2(n2942), .ZN(n3408) );
  NAND2_X1 U2503 ( .A1(n3248), .A2(n2932), .ZN(n2184) );
  OR2_X1 U2504 ( .A1(n3383), .A2(n3258), .ZN(n2933) );
  OR2_X1 U2505 ( .A1(n4655), .A2(n4489), .ZN(n3008) );
  NAND2_X1 U2506 ( .A1(n3045), .A2(n3912), .ZN(n4365) );
  OR2_X1 U2507 ( .A1(n3016), .A2(n3975), .ZN(n3058) );
  AND2_X1 U2508 ( .A1(n3448), .A2(n3528), .ZN(n3520) );
  AND2_X1 U2509 ( .A1(n3368), .A2(n4049), .ZN(n4437) );
  INV_X1 U2510 ( .A(n3088), .ZN(n2867) );
  NAND2_X1 U2511 ( .A1(n2866), .A2(n3088), .ZN(n3087) );
  AND2_X1 U2512 ( .A1(n2161), .A2(n2340), .ZN(n2365) );
  NAND2_X1 U2513 ( .A1(n2361), .A2(n2303), .ZN(n2302) );
  INV_X1 U2514 ( .A(IR_REG_18__SCAN_IN), .ZN(n2303) );
  AND2_X1 U2515 ( .A1(n2477), .A2(n2476), .ZN(n3233) );
  INV_X1 U2516 ( .A(n4067), .ZN(n3296) );
  INV_X1 U2517 ( .A(n4280), .ZN(n4404) );
  NAND2_X1 U2518 ( .A1(n2322), .A2(n2918), .ZN(n2919) );
  AND2_X1 U2519 ( .A1(n2819), .A2(n2805), .ZN(n4213) );
  INV_X1 U2520 ( .A(n3885), .ZN(n3866) );
  NAND2_X1 U2521 ( .A1(n4556), .A2(n4557), .ZN(n4555) );
  NOR2_X1 U2522 ( .A1(n4586), .A2(n4126), .ZN(n4595) );
  OAI21_X1 U2523 ( .B1(n4601), .B2(n2248), .A(n2247), .ZN(n2246) );
  AOI21_X1 U2524 ( .B1(n4604), .B2(ADDR_REG_18__SCAN_IN), .A(n4603), .ZN(n2247) );
  NAND2_X1 U2525 ( .A1(n2249), .A2(n4549), .ZN(n2248) );
  NAND2_X1 U2526 ( .A1(n2250), .A2(n4602), .ZN(n2249) );
  INV_X1 U2527 ( .A(n4148), .ZN(n4285) );
  NAND2_X1 U2528 ( .A1(n4357), .A2(n3355), .ZN(n4360) );
  INV_X1 U2529 ( .A(n4331), .ZN(n4621) );
  NAND2_X1 U2530 ( .A1(n2310), .A2(n4365), .ZN(n4152) );
  NAND2_X1 U2531 ( .A1(n3059), .A2(n4149), .ZN(n2310) );
  INV_X1 U2532 ( .A(IR_REG_29__SCAN_IN), .ZN(n2344) );
  INV_X1 U2533 ( .A(n4103), .ZN(n4632) );
  NOR2_X1 U2534 ( .A1(n2288), .A2(n2292), .ZN(n2287) );
  INV_X1 U2535 ( .A(n2297), .ZN(n2288) );
  INV_X1 U2536 ( .A(n2291), .ZN(n2290) );
  OAI21_X1 U2537 ( .B1(n2294), .B2(n2292), .A(n3700), .ZN(n2291) );
  CLKBUF_X1 U2538 ( .A(n2968), .Z(n3980) );
  OR2_X1 U2539 ( .A1(n3848), .A2(n2280), .ZN(n2279) );
  INV_X1 U2540 ( .A(n2283), .ZN(n2280) );
  AND2_X1 U2541 ( .A1(n3871), .A2(n2274), .ZN(n2271) );
  NOR2_X1 U2542 ( .A1(n2279), .A2(n2275), .ZN(n2274) );
  INV_X1 U2543 ( .A(n3797), .ZN(n2275) );
  INV_X1 U2544 ( .A(IR_REG_4__SCAN_IN), .ZN(n4904) );
  AND2_X1 U2545 ( .A1(n2836), .A2(REG3_REG_27__SCAN_IN), .ZN(n2847) );
  AOI21_X1 U2546 ( .B1(n3962), .B2(n2948), .A(n2177), .ZN(n2188) );
  INV_X1 U2547 ( .A(n2948), .ZN(n2186) );
  INV_X1 U2548 ( .A(n3087), .ZN(n2880) );
  NOR2_X1 U2549 ( .A1(n3058), .A2(n3044), .ZN(n3045) );
  NOR2_X1 U2550 ( .A1(n4246), .A2(n2313), .ZN(n2312) );
  INV_X1 U2551 ( .A(n4265), .ZN(n2313) );
  OR2_X1 U2552 ( .A1(n3723), .A2(n4430), .ZN(n3722) );
  NOR2_X1 U2553 ( .A1(n2318), .A2(n3677), .ZN(n2317) );
  INV_X1 U2554 ( .A(n2319), .ZN(n2318) );
  NOR2_X1 U2555 ( .A1(n3619), .A2(n3547), .ZN(n2319) );
  NOR2_X1 U2556 ( .A1(n3457), .A2(n3167), .ZN(n3166) );
  INV_X1 U2557 ( .A(IR_REG_28__SCAN_IN), .ZN(n2903) );
  NAND2_X1 U2558 ( .A1(n2157), .A2(IR_REG_31__SCAN_IN), .ZN(n2884) );
  INV_X1 U2559 ( .A(IR_REG_23__SCAN_IN), .ZN(n2883) );
  INV_X1 U2560 ( .A(IR_REG_20__SCAN_IN), .ZN(n4912) );
  INV_X1 U2561 ( .A(IR_REG_8__SCAN_IN), .ZN(n2253) );
  OR2_X1 U2562 ( .A1(n2613), .A2(n2612), .ZN(n2628) );
  INV_X1 U2563 ( .A(IR_REG_6__SCAN_IN), .ZN(n2511) );
  NOR2_X1 U2564 ( .A1(IR_REG_4__SCAN_IN), .A2(IR_REG_3__SCAN_IN), .ZN(n2306)
         );
  INV_X1 U2565 ( .A(IR_REG_1__SCAN_IN), .ZN(n2307) );
  INV_X1 U2566 ( .A(IR_REG_2__SCAN_IN), .ZN(n2308) );
  AND2_X1 U2567 ( .A1(n2766), .A2(n3837), .ZN(n3755) );
  XNOR2_X1 U2568 ( .A(n2388), .B(n2844), .ZN(n2405) );
  OR2_X1 U2569 ( .A1(n2572), .A2(n4923), .ZN(n2593) );
  INV_X1 U2570 ( .A(REG3_REG_12__SCAN_IN), .ZN(n2592) );
  INV_X1 U2571 ( .A(n2600), .ZN(n2861) );
  NAND2_X1 U2572 ( .A1(n3329), .A2(n3330), .ZN(n2267) );
  NAND2_X1 U2573 ( .A1(n2270), .A2(n2269), .ZN(n2268) );
  INV_X1 U2574 ( .A(n3330), .ZN(n2269) );
  INV_X1 U2575 ( .A(n3329), .ZN(n2270) );
  AND2_X1 U2576 ( .A1(n2606), .A2(REG3_REG_13__SCAN_IN), .ZN(n2622) );
  INV_X1 U2577 ( .A(n2295), .ZN(n2293) );
  NOR2_X1 U2578 ( .A1(n2167), .A2(n2263), .ZN(n2262) );
  INV_X1 U2579 ( .A(n3829), .ZN(n2263) );
  NAND2_X1 U2580 ( .A1(n2256), .A2(n2255), .ZN(n2257) );
  NAND2_X1 U2581 ( .A1(n2424), .A2(n2423), .ZN(n2425) );
  NAND2_X1 U2582 ( .A1(n2285), .A2(n2284), .ZN(n2283) );
  INV_X1 U2583 ( .A(n3807), .ZN(n2284) );
  INV_X1 U2584 ( .A(n3808), .ZN(n2285) );
  INV_X1 U2585 ( .A(n2679), .ZN(n2281) );
  AND2_X1 U2586 ( .A1(n3871), .A2(n3797), .ZN(n2272) );
  OR2_X1 U2587 ( .A1(n2683), .A2(n2682), .ZN(n2699) );
  NAND2_X1 U2588 ( .A1(n2622), .A2(REG3_REG_14__SCAN_IN), .ZN(n2644) );
  INV_X1 U2589 ( .A(REG3_REG_15__SCAN_IN), .ZN(n2643) );
  OR2_X1 U2590 ( .A1(n2644), .A2(n2643), .ZN(n2683) );
  NAND4_X1 U2591 ( .A1(n2221), .A2(n2160), .A3(n2220), .A4(n2218), .ZN(n3119)
         );
  NOR2_X1 U2592 ( .A1(n3119), .A2(n3120), .ZN(n3134) );
  NOR2_X1 U2593 ( .A1(n3206), .A2(n2447), .ZN(n3205) );
  AND2_X1 U2594 ( .A1(n2236), .A2(n4495), .ZN(n2234) );
  XNOR2_X1 U2595 ( .A(n3276), .B(n3232), .ZN(n3235) );
  NOR2_X1 U2596 ( .A1(n3235), .A2(n3321), .ZN(n3277) );
  NOR2_X1 U2597 ( .A1(n3284), .A2(n2242), .ZN(n2241) );
  NOR2_X1 U2598 ( .A1(n3284), .A2(n3232), .ZN(n2240) );
  AND2_X1 U2599 ( .A1(n2244), .A2(n2243), .ZN(n4086) );
  NAND2_X1 U2600 ( .A1(n4492), .A2(REG2_REG_7__SCAN_IN), .ZN(n2243) );
  OAI22_X1 U2601 ( .A1(n4108), .A2(n4934), .B1(n4107), .B2(n4106), .ZN(n4508)
         );
  NAND2_X1 U2602 ( .A1(n4508), .A2(n4509), .ZN(n4507) );
  XNOR2_X1 U2603 ( .A(n4113), .B(n4644), .ZN(n4519) );
  NAND2_X1 U2604 ( .A1(n4519), .A2(REG1_REG_10__SCAN_IN), .ZN(n4518) );
  XNOR2_X1 U2605 ( .A(n4093), .B(n4641), .ZN(n4539) );
  AOI21_X1 U2606 ( .B1(n4551), .B2(n4095), .A(n2245), .ZN(n4096) );
  AND2_X1 U2607 ( .A1(n4548), .A2(REG2_REG_13__SCAN_IN), .ZN(n2245) );
  XNOR2_X1 U2608 ( .A(n4099), .B(n4125), .ZN(n4582) );
  INV_X1 U2609 ( .A(n4594), .ZN(n2229) );
  NAND2_X1 U2610 ( .A1(n4590), .A2(n2251), .ZN(n2250) );
  OR2_X1 U2611 ( .A1(n4633), .A2(REG2_REG_17__SCAN_IN), .ZN(n2251) );
  OAI21_X1 U2612 ( .B1(n4204), .B2(n4036), .A(n3001), .ZN(n3002) );
  NAND2_X1 U2613 ( .A1(n2197), .A2(n2196), .ZN(n3027) );
  AOI21_X1 U2614 ( .B1(n2146), .B2(n2202), .A(n2170), .ZN(n2196) );
  NAND2_X1 U2615 ( .A1(n2207), .A2(n2206), .ZN(n4256) );
  AOI21_X1 U2616 ( .B1(n2166), .B2(n2212), .A(n2152), .ZN(n2206) );
  NAND2_X1 U2617 ( .A1(n4315), .A2(n2956), .ZN(n2214) );
  OR2_X1 U2618 ( .A1(n3038), .A2(IR_REG_28__SCAN_IN), .ZN(n2378) );
  NAND2_X1 U2619 ( .A1(n3738), .A2(n4430), .ZN(n2951) );
  OR2_X1 U2620 ( .A1(n3654), .A2(n3933), .ZN(n3655) );
  AOI21_X1 U2621 ( .B1(n2194), .B2(n2192), .A(n2175), .ZN(n2191) );
  INV_X1 U2622 ( .A(n2949), .ZN(n2192) );
  INV_X1 U2623 ( .A(n2194), .ZN(n2193) );
  OR2_X1 U2624 ( .A1(n3512), .A2(n3962), .ZN(n3510) );
  AND2_X1 U2625 ( .A1(n3602), .A2(n2982), .ZN(n3962) );
  CLKBUF_X1 U2626 ( .A(n3509), .Z(n3600) );
  OR2_X1 U2627 ( .A1(n3404), .A2(n4006), .ZN(n2980) );
  NOR2_X1 U2628 ( .A1(n2537), .A2(n2536), .ZN(n2551) );
  OR2_X1 U2629 ( .A1(n3418), .A2(n2976), .ZN(n2977) );
  OR2_X1 U2630 ( .A1(n4066), .A2(n3360), .ZN(n2939) );
  INV_X1 U2631 ( .A(n3309), .ZN(n3422) );
  AND2_X1 U2632 ( .A1(n3993), .A2(n3995), .ZN(n3968) );
  INV_X1 U2633 ( .A(n4145), .ZN(n4281) );
  OR2_X1 U2634 ( .A1(n3381), .A2(n2972), .ZN(n2973) );
  AND2_X1 U2635 ( .A1(REG3_REG_3__SCAN_IN), .A2(REG3_REG_4__SCAN_IN), .ZN(
        n2466) );
  NAND2_X1 U2636 ( .A1(n2183), .A2(n2970), .ZN(n3178) );
  INV_X1 U2637 ( .A(n2970), .ZN(n3967) );
  NOR2_X1 U2638 ( .A1(n4365), .A2(n4366), .ZN(n4364) );
  AND2_X1 U2639 ( .A1(n3923), .A2(n4138), .ZN(n3040) );
  AND2_X1 U2640 ( .A1(n4264), .A2(n2154), .ZN(n4209) );
  NAND2_X1 U2641 ( .A1(n4264), .A2(n2153), .ZN(n4226) );
  NAND2_X1 U2642 ( .A1(n4264), .A2(n2312), .ZN(n4248) );
  NAND2_X1 U2643 ( .A1(n4264), .A2(n4265), .ZN(n4267) );
  NOR2_X1 U2644 ( .A1(n4328), .A2(n4298), .ZN(n4306) );
  OR2_X1 U2645 ( .A1(n4350), .A2(n3771), .ZN(n4328) );
  NOR2_X1 U2646 ( .A1(n3722), .A2(n4420), .ZN(n4352) );
  AND2_X1 U2647 ( .A1(n3520), .A2(n2315), .ZN(n3658) );
  NOR2_X1 U2648 ( .A1(n2316), .A2(n3015), .ZN(n2315) );
  INV_X1 U2649 ( .A(n2317), .ZN(n2316) );
  NAND2_X1 U2650 ( .A1(n3520), .A2(n2317), .ZN(n3648) );
  NAND2_X1 U2651 ( .A1(n3520), .A2(n2319), .ZN(n3646) );
  NAND2_X1 U2652 ( .A1(n3520), .A2(n3519), .ZN(n3593) );
  INV_X1 U2653 ( .A(n3490), .ZN(n3528) );
  AND2_X1 U2654 ( .A1(n3319), .A2(n2179), .ZN(n3448) );
  NAND2_X1 U2655 ( .A1(n3319), .A2(n2314), .ZN(n3551) );
  NAND2_X1 U2656 ( .A1(n3319), .A2(n2150), .ZN(n3552) );
  AND2_X1 U2657 ( .A1(n3319), .A2(n3318), .ZN(n3423) );
  OR2_X1 U2658 ( .A1(n3256), .A2(n3382), .ZN(n3390) );
  NOR2_X1 U2659 ( .A1(n3390), .A2(n3435), .ZN(n3319) );
  INV_X1 U2660 ( .A(n4378), .ZN(n4431) );
  INV_X1 U2661 ( .A(n4374), .ZN(n4434) );
  INV_X1 U2662 ( .A(n4437), .ZN(n4654) );
  NAND2_X1 U2663 ( .A1(n2375), .A2(IR_REG_31__SCAN_IN), .ZN(n3038) );
  XNOR2_X1 U2664 ( .A(n2386), .B(n2385), .ZN(n2912) );
  NAND2_X1 U2665 ( .A1(n2158), .A2(IR_REG_31__SCAN_IN), .ZN(n2386) );
  NAND2_X1 U2666 ( .A1(n2156), .A2(IR_REG_31__SCAN_IN), .ZN(n2387) );
  AND2_X1 U2667 ( .A1(n2665), .A2(n2653), .ZN(n4104) );
  AND2_X1 U2668 ( .A1(n2580), .A2(n2597), .ZN(n4115) );
  AND2_X1 U2669 ( .A1(n2545), .A2(n2613), .ZN(n4110) );
  INV_X1 U2670 ( .A(IR_REG_7__SCAN_IN), .ZN(n2252) );
  CLKBUF_X1 U2671 ( .A(n2474), .Z(n2475) );
  INV_X1 U2672 ( .A(IR_REG_3__SCAN_IN), .ZN(n2433) );
  NOR2_X1 U2673 ( .A1(n3262), .A2(n2260), .ZN(n2259) );
  INV_X1 U2674 ( .A(n2486), .ZN(n2260) );
  NAND2_X1 U2675 ( .A1(n2296), .A2(n2294), .ZN(n2289) );
  NAND2_X1 U2676 ( .A1(n2301), .A2(n2151), .ZN(n2923) );
  CLKBUF_X1 U2677 ( .A(n2927), .Z(n3461) );
  INV_X1 U2678 ( .A(n3741), .ZN(n4420) );
  INV_X1 U2679 ( .A(n4298), .ZN(n4308) );
  NOR2_X1 U2680 ( .A1(n2905), .A2(n3114), .ZN(n3798) );
  NAND2_X1 U2681 ( .A1(n2276), .A2(n2283), .ZN(n3851) );
  NAND2_X1 U2682 ( .A1(n2282), .A2(n2165), .ZN(n2276) );
  INV_X1 U2683 ( .A(n3880), .ZN(n3862) );
  AND2_X1 U2684 ( .A1(n2901), .A2(n3106), .ZN(n3885) );
  INV_X1 U2685 ( .A(n3798), .ZN(n3877) );
  INV_X1 U2686 ( .A(n3869), .ZN(n3874) );
  NAND2_X1 U2687 ( .A1(n2855), .A2(n2854), .ZN(n4174) );
  NAND2_X1 U2688 ( .A1(n2811), .A2(n2810), .ZN(n4385) );
  NAND2_X1 U2689 ( .A1(n2771), .A2(n2770), .ZN(n4261) );
  OR2_X1 U2690 ( .A1(n2737), .A2(n2736), .ZN(n4280) );
  OR2_X1 U2691 ( .A1(n2721), .A2(n2720), .ZN(n4344) );
  NAND4_X1 U2692 ( .A1(n2526), .A2(n2525), .A3(n2524), .A4(n2523), .ZN(n3496)
         );
  OR2_X1 U2693 ( .A1(n2510), .A2(n2509), .ZN(n4065) );
  OR2_X1 U2694 ( .A1(n2449), .A2(n2448), .ZN(n4067) );
  AND3_X1 U2695 ( .A1(n2429), .A2(n2428), .A3(n2427), .ZN(n2431) );
  AND2_X1 U2696 ( .A1(n2412), .A2(n2411), .ZN(n2413) );
  AND2_X1 U2697 ( .A1(n3113), .A2(n3112), .ZN(n4503) );
  NAND2_X1 U2698 ( .A1(n4076), .A2(n3115), .ZN(n3186) );
  INV_X1 U2699 ( .A(REG2_REG_2__SCAN_IN), .ZN(n2239) );
  INV_X1 U2700 ( .A(n2224), .ZN(n3191) );
  NAND2_X1 U2701 ( .A1(n2232), .A2(REG1_REG_4__SCAN_IN), .ZN(n2231) );
  NAND2_X1 U2702 ( .A1(n2327), .A2(n2232), .ZN(n2230) );
  INV_X1 U2703 ( .A(n3138), .ZN(n2232) );
  INV_X1 U2704 ( .A(n2225), .ZN(n3337) );
  AOI21_X1 U2705 ( .B1(n3283), .B2(REG2_REG_6__SCAN_IN), .A(n2181), .ZN(n3285)
         );
  NAND2_X1 U2706 ( .A1(n4565), .A2(n4122), .ZN(n4576) );
  NAND2_X1 U2707 ( .A1(n4576), .A2(n4577), .ZN(n4575) );
  XNOR2_X1 U2708 ( .A(n4124), .B(n4125), .ZN(n4585) );
  OR2_X1 U2709 ( .A1(n2820), .A2(n2836), .ZN(n4198) );
  OR2_X1 U2710 ( .A1(n4315), .A2(n2212), .ZN(n2209) );
  NAND2_X1 U2711 ( .A1(n2195), .A2(n2194), .ZN(n3581) );
  NAND2_X1 U2712 ( .A1(n2950), .A2(n2949), .ZN(n2195) );
  INV_X1 U2713 ( .A(n4360), .ZN(n4277) );
  OR2_X1 U2714 ( .A1(n4355), .A2(n4654), .ZN(n4331) );
  OR2_X1 U2715 ( .A1(n3346), .A2(n3008), .ZN(n4332) );
  INV_X1 U2716 ( .A(REG1_REG_0__SCAN_IN), .ZN(n4676) );
  AND2_X1 U2717 ( .A1(n4167), .A2(n3055), .ZN(n3056) );
  INV_X1 U2718 ( .A(n4630), .ZN(n3092) );
  XNOR2_X1 U2719 ( .A(n2254), .B(IR_REG_24__SCAN_IN), .ZN(n3089) );
  NAND2_X1 U2720 ( .A1(n2882), .A2(IR_REG_31__SCAN_IN), .ZN(n2254) );
  NAND2_X1 U2721 ( .A1(n3087), .A2(n3107), .ZN(n4628) );
  AND2_X1 U2722 ( .A1(n2364), .A2(n2375), .ZN(n3088) );
  NAND2_X1 U2723 ( .A1(n3095), .A2(STATE_REG_SCAN_IN), .ZN(n4630) );
  INV_X1 U2724 ( .A(n2912), .ZN(n4057) );
  AND2_X1 U2725 ( .A1(n2371), .A2(n2158), .ZN(n4489) );
  OR2_X1 U2726 ( .A1(n2360), .A2(n2302), .ZN(n2369) );
  XNOR2_X1 U2727 ( .A(n2387), .B(IR_REG_19__SCAN_IN), .ZN(n4490) );
  INV_X1 U2728 ( .A(n4117), .ZN(n4641) );
  INV_X1 U2729 ( .A(n4115), .ZN(n4643) );
  XNOR2_X1 U2730 ( .A(n2415), .B(IR_REG_2__SCAN_IN), .ZN(n4496) );
  OAI21_X1 U2731 ( .B1(IR_REG_0__SCAN_IN), .B2(IR_REG_1__SCAN_IN), .A(
        IR_REG_31__SCAN_IN), .ZN(n2415) );
  NOR2_X1 U2732 ( .A1(n4595), .A2(n4594), .ZN(n4596) );
  INV_X1 U2733 ( .A(n2246), .ZN(n4609) );
  AOI211_X1 U2734 ( .C1(n4621), .C2(n4170), .A(n4169), .B(n4168), .ZN(n4171)
         );
  INV_X1 U2735 ( .A(n3067), .ZN(n3068) );
  OR2_X1 U2736 ( .A1(n4173), .A2(n4428), .ZN(n3018) );
  OAI21_X1 U2737 ( .B1(n4152), .B2(n4485), .A(n3046), .ZN(n3047) );
  NAND2_X1 U2738 ( .A1(n4673), .A2(REG0_REG_29__SCAN_IN), .ZN(n3046) );
  OR2_X1 U2739 ( .A1(n4173), .A2(n4485), .ZN(n3024) );
  NAND2_X1 U2740 ( .A1(n2675), .A2(n2272), .ZN(n2282) );
  AND2_X1 U2741 ( .A1(n2204), .A2(n2205), .ZN(n4207) );
  NOR2_X1 U2742 ( .A1(n2962), .A2(n2198), .ZN(n2146) );
  NAND2_X1 U2743 ( .A1(n4496), .A2(REG1_REG_2__SCAN_IN), .ZN(n2147) );
  INV_X1 U2744 ( .A(IR_REG_25__SCAN_IN), .ZN(n2366) );
  OR2_X1 U2745 ( .A1(n2304), .A2(IR_REG_22__SCAN_IN), .ZN(n2148) );
  AND2_X1 U2746 ( .A1(n4061), .A2(n3881), .ZN(n2149) );
  AND2_X1 U2747 ( .A1(n2214), .A2(n2215), .ZN(n4291) );
  AND2_X1 U2748 ( .A1(n2314), .A2(n3553), .ZN(n2150) );
  NOR2_X1 U2749 ( .A1(n3747), .A2(n2300), .ZN(n2151) );
  AND2_X1 U2750 ( .A1(n4300), .A2(n4286), .ZN(n2152) );
  AND2_X1 U2751 ( .A1(n2312), .A2(n4231), .ZN(n2153) );
  AND2_X1 U2752 ( .A1(n2153), .A2(n4216), .ZN(n2154) );
  INV_X1 U2753 ( .A(n2455), .ZN(n2695) );
  NAND2_X1 U2754 ( .A1(n2340), .A2(n2474), .ZN(n2360) );
  AND2_X2 U2755 ( .A1(n3070), .A2(n2963), .ZN(n2600) );
  AND4_X1 U2756 ( .A1(n2343), .A2(n2342), .A3(n2341), .A4(n2385), .ZN(n2155)
         );
  NAND2_X1 U2757 ( .A1(n3825), .A2(n2262), .ZN(n3754) );
  AOI21_X1 U2758 ( .B1(n4126), .B2(n2229), .A(n4128), .ZN(n2228) );
  OR2_X1 U2759 ( .A1(n2360), .A2(IR_REG_18__SCAN_IN), .ZN(n2156) );
  OR2_X1 U2760 ( .A1(n2360), .A2(n2148), .ZN(n2157) );
  NAND2_X1 U2761 ( .A1(n3825), .A2(n3829), .ZN(n3774) );
  NAND2_X1 U2762 ( .A1(n2199), .A2(n2200), .ZN(n4184) );
  OR2_X1 U2763 ( .A1(n2360), .A2(n2304), .ZN(n2158) );
  NOR2_X1 U2764 ( .A1(n4064), .A2(n3495), .ZN(n2159) );
  INV_X1 U2765 ( .A(IR_REG_22__SCAN_IN), .ZN(n2385) );
  OR2_X1 U2766 ( .A1(n2147), .A2(n2235), .ZN(n2160) );
  AND2_X1 U2767 ( .A1(n2474), .A2(n2155), .ZN(n2161) );
  NAND2_X1 U2768 ( .A1(n4064), .A2(n3495), .ZN(n2162) );
  AND2_X1 U2769 ( .A1(n4941), .A2(n2903), .ZN(n2163) );
  AND2_X1 U2770 ( .A1(n2227), .A2(n2228), .ZN(n2164) );
  INV_X1 U2771 ( .A(n2419), .ZN(n2900) );
  NOR2_X1 U2772 ( .A1(n2698), .A2(n2281), .ZN(n2165) );
  AND2_X1 U2773 ( .A1(n4306), .A2(n4286), .ZN(n4264) );
  NAND2_X1 U2774 ( .A1(n2289), .A2(n3669), .ZN(n3699) );
  NAND2_X1 U2775 ( .A1(n2282), .A2(n2679), .ZN(n3806) );
  NAND2_X1 U2776 ( .A1(n2209), .A2(n2210), .ZN(n4275) );
  NAND2_X1 U2777 ( .A1(n2296), .A2(n2293), .ZN(n3667) );
  NOR2_X1 U2778 ( .A1(n2957), .A2(n2208), .ZN(n2166) );
  AND2_X1 U2779 ( .A1(n3776), .A2(n3775), .ZN(n2167) );
  OR2_X1 U2780 ( .A1(n4061), .A2(n3881), .ZN(n2168) );
  OR2_X1 U2781 ( .A1(n3623), .A2(n2984), .ZN(n2169) );
  AND2_X1 U2782 ( .A1(n4379), .A2(n4196), .ZN(n2170) );
  OR2_X1 U2783 ( .A1(n2596), .A2(n2595), .ZN(n3513) );
  INV_X1 U2784 ( .A(n3513), .ZN(n3675) );
  AND2_X1 U2785 ( .A1(n2334), .A2(n2325), .ZN(n2171) );
  NOR2_X1 U2786 ( .A1(n4385), .A2(n4373), .ZN(n2172) );
  NOR2_X1 U2787 ( .A1(n4280), .A2(n4298), .ZN(n2173) );
  AND2_X1 U2788 ( .A1(n4385), .A2(n4373), .ZN(n2174) );
  NOR2_X1 U2789 ( .A1(n3674), .A2(n3015), .ZN(n2175) );
  NOR2_X1 U2790 ( .A1(n4404), .A2(n4308), .ZN(n2176) );
  NOR2_X1 U2791 ( .A1(n3675), .A2(n3575), .ZN(n2177) );
  AND2_X1 U2792 ( .A1(n3675), .A2(n3575), .ZN(n2178) );
  INV_X1 U2793 ( .A(n3858), .ZN(n2300) );
  AND2_X1 U2794 ( .A1(n2150), .A2(n2979), .ZN(n2179) );
  INV_X1 U2795 ( .A(n2330), .ZN(n2205) );
  OAI21_X1 U2796 ( .B1(n3312), .B2(n2940), .A(n2939), .ZN(n3406) );
  NAND2_X1 U2797 ( .A1(n2266), .A2(n2264), .ZN(n3473) );
  NOR3_X1 U2798 ( .A1(n2900), .A2(n4630), .A3(n2899), .ZN(n2180) );
  NAND2_X1 U2799 ( .A1(n3510), .A2(n2948), .ZN(n3592) );
  NAND2_X1 U2800 ( .A1(n2261), .A2(n2486), .ZN(n3260) );
  NAND2_X1 U2801 ( .A1(n2266), .A2(n2267), .ZN(n3472) );
  AND2_X1 U2802 ( .A1(n2195), .A2(n2169), .ZN(n3580) );
  NAND2_X1 U2803 ( .A1(n2184), .A2(n2933), .ZN(n3378) );
  INV_X1 U2804 ( .A(n3089), .ZN(n2864) );
  INV_X1 U2805 ( .A(n2955), .ZN(n2215) );
  AND2_X1 U2806 ( .A1(n3282), .A2(n4493), .ZN(n2181) );
  INV_X1 U2807 ( .A(n4549), .ZN(n4600) );
  AND2_X1 U2808 ( .A1(n4503), .A2(n4055), .ZN(n4549) );
  INV_X1 U2809 ( .A(n4216), .ZN(n4373) );
  NOR2_X1 U2810 ( .A1(n3205), .A2(n2327), .ZN(n2182) );
  AND2_X1 U2811 ( .A1(n2450), .A2(n2435), .ZN(n4495) );
  INV_X1 U2812 ( .A(n4495), .ZN(n2235) );
  INV_X1 U2813 ( .A(REG2_REG_6__SCAN_IN), .ZN(n2242) );
  INV_X1 U2814 ( .A(n3176), .ZN(n2183) );
  NAND2_X1 U2815 ( .A1(n3460), .A2(n2929), .ZN(n3176) );
  NAND2_X1 U2816 ( .A1(n2965), .A2(n3458), .ZN(n3460) );
  NAND3_X1 U2817 ( .A1(n2184), .A2(n2933), .A3(n3379), .ZN(n3377) );
  OAI21_X1 U2818 ( .B1(n3512), .B2(n2187), .A(n2185), .ZN(n3634) );
  OAI21_X1 U2819 ( .B1(n2950), .B2(n2193), .A(n2191), .ZN(n3657) );
  OR2_X1 U2820 ( .A1(n4224), .A2(n2202), .ZN(n2199) );
  NAND2_X1 U2821 ( .A1(n4224), .A2(n2146), .ZN(n2197) );
  NAND2_X1 U2822 ( .A1(n4224), .A2(n2961), .ZN(n2204) );
  INV_X1 U2823 ( .A(n2203), .ZN(n2202) );
  NAND2_X1 U2824 ( .A1(n4315), .A2(n2166), .ZN(n2207) );
  NAND4_X1 U2825 ( .A1(n2340), .A2(n2474), .A3(n2155), .A4(n2311), .ZN(n2375)
         );
  NAND2_X1 U2826 ( .A1(n4543), .A2(n4119), .ZN(n4556) );
  NAND2_X1 U2827 ( .A1(n4544), .A2(REG1_REG_12__SCAN_IN), .ZN(n4543) );
  NAND2_X1 U2828 ( .A1(n2223), .A2(n2222), .ZN(n2224) );
  NOR2_X1 U2829 ( .A1(n2222), .A2(n4495), .ZN(n2219) );
  NAND3_X1 U2830 ( .A1(n2223), .A2(n2222), .A3(n4495), .ZN(n2220) );
  NAND3_X1 U2831 ( .A1(n3192), .A2(n2147), .A3(n2235), .ZN(n2221) );
  INV_X1 U2832 ( .A(n3193), .ZN(n2222) );
  NAND3_X1 U2833 ( .A1(n2227), .A2(n4607), .A3(n2228), .ZN(n4605) );
  NAND2_X1 U2834 ( .A1(n4586), .A2(n2229), .ZN(n2227) );
  NAND2_X1 U2835 ( .A1(n4496), .A2(REG2_REG_2__SCAN_IN), .ZN(n2237) );
  XNOR2_X1 U2836 ( .A(n4496), .B(n2239), .ZN(n3185) );
  AOI22_X1 U2837 ( .A1(n3283), .A2(n2241), .B1(n3282), .B2(n2240), .ZN(n2244)
         );
  INV_X1 U2838 ( .A(n2244), .ZN(n3338) );
  NAND2_X1 U2839 ( .A1(n3103), .A2(n3104), .ZN(n2258) );
  NAND4_X1 U2840 ( .A1(n2258), .A2(n2257), .A3(n2408), .A4(n2425), .ZN(n3126)
         );
  INV_X1 U2841 ( .A(n2423), .ZN(n2255) );
  INV_X1 U2842 ( .A(n2424), .ZN(n2256) );
  NAND2_X1 U2843 ( .A1(n2257), .A2(n2425), .ZN(n3128) );
  NAND2_X1 U2844 ( .A1(n2258), .A2(n2408), .ZN(n3125) );
  NAND2_X1 U2845 ( .A1(n2261), .A2(n2259), .ZN(n2504) );
  NAND2_X1 U2846 ( .A1(n3222), .A2(n3223), .ZN(n2261) );
  NAND2_X1 U2847 ( .A1(n3328), .A2(n2268), .ZN(n2266) );
  NAND2_X1 U2848 ( .A1(n2675), .A2(n2271), .ZN(n2273) );
  NAND2_X1 U2849 ( .A1(n2273), .A2(n2277), .ZN(n3767) );
  NAND2_X1 U2850 ( .A1(n3570), .A2(n2297), .ZN(n2296) );
  NAND2_X1 U2851 ( .A1(n2286), .A2(n2290), .ZN(n2636) );
  NAND2_X1 U2852 ( .A1(n3570), .A2(n2287), .ZN(n2286) );
  NAND2_X1 U2853 ( .A1(n2301), .A2(n3858), .ZN(n3748) );
  INV_X1 U2854 ( .A(n2923), .ZN(n2921) );
  NAND3_X1 U2855 ( .A1(n2309), .A2(n2307), .A3(n2308), .ZN(n2432) );
  NAND4_X1 U2856 ( .A1(n2306), .A2(n2309), .A3(n2308), .A4(n2307), .ZN(n2472)
         );
  INV_X2 U2857 ( .A(IR_REG_0__SCAN_IN), .ZN(n2309) );
  NAND2_X1 U2858 ( .A1(n2365), .A2(n2366), .ZN(n2362) );
  NAND2_X1 U2859 ( .A1(n3070), .A2(n3092), .ZN(n3346) );
  NAND2_X1 U2860 ( .A1(n4352), .A2(n4351), .ZN(n4350) );
  NAND2_X1 U2861 ( .A1(n3658), .A2(n3662), .ZN(n3723) );
  NAND2_X1 U2862 ( .A1(n4209), .A2(n4196), .ZN(n3016) );
  AND2_X4 U2863 ( .A1(n3070), .A2(n3354), .ZN(n2419) );
  AND2_X1 U2864 ( .A1(n3462), .A2(n2966), .ZN(n3458) );
  OAI21_X1 U2865 ( .B1(n4152), .B2(n4428), .A(n3066), .ZN(n3067) );
  AND2_X1 U2866 ( .A1(n3909), .A2(DATAI_20_), .ZN(n4298) );
  NAND2_X1 U2867 ( .A1(n3909), .A2(DATAI_2_), .ZN(n2416) );
  INV_X2 U2868 ( .A(n4680), .ZN(n4682) );
  OR2_X1 U2869 ( .A1(n3021), .A2(n3352), .ZN(n4680) );
  INV_X2 U2870 ( .A(n4673), .ZN(n4675) );
  NOR2_X1 U2871 ( .A1(n2792), .A2(n3756), .ZN(n2320) );
  NOR2_X1 U2872 ( .A1(n2799), .A2(n3756), .ZN(n2321) );
  OR3_X1 U2873 ( .A1(n2893), .A2(n3869), .A3(n2325), .ZN(n2322) );
  AND2_X1 U2874 ( .A1(n4432), .A2(n4420), .ZN(n2323) );
  AND2_X1 U2875 ( .A1(n3116), .A2(REG1_REG_1__SCAN_IN), .ZN(n2324) );
  NAND2_X1 U2876 ( .A1(n2892), .A2(n2891), .ZN(n2325) );
  AND2_X1 U2877 ( .A1(n3233), .A2(REG1_REG_5__SCAN_IN), .ZN(n2326) );
  INV_X1 U2878 ( .A(n3623), .ZN(n4062) );
  AND2_X1 U2879 ( .A1(n2609), .A2(n2608), .ZN(n3623) );
  INV_X1 U2880 ( .A(IR_REG_30__SCAN_IN), .ZN(n2345) );
  NAND2_X1 U2881 ( .A1(n2802), .A2(n2801), .ZN(n3815) );
  AND2_X1 U2882 ( .A1(n3137), .A2(n4494), .ZN(n2327) );
  INV_X1 U2883 ( .A(n2984), .ZN(n3677) );
  NOR2_X1 U2884 ( .A1(n3496), .A2(n3558), .ZN(n2328) );
  INV_X1 U2885 ( .A(IR_REG_27__SCAN_IN), .ZN(n4941) );
  OR2_X1 U2886 ( .A1(n3780), .A2(n4265), .ZN(n2329) );
  AND2_X1 U2887 ( .A1(n4245), .A2(n4231), .ZN(n2330) );
  INV_X1 U2888 ( .A(n3881), .ZN(n3662) );
  OR2_X1 U2889 ( .A1(n4159), .A2(n4485), .ZN(n2331) );
  OR2_X1 U2890 ( .A1(n4159), .A2(n4428), .ZN(n2332) );
  OR2_X1 U2891 ( .A1(n4146), .A2(n4166), .ZN(n2333) );
  NOR2_X1 U2892 ( .A1(n2922), .A2(n3869), .ZN(n2334) );
  XNOR2_X1 U2893 ( .A(n2405), .B(n2406), .ZN(n3103) );
  NAND2_X1 U2894 ( .A1(n3987), .A2(n3990), .ZN(n3379) );
  INV_X1 U2895 ( .A(n4421), .ZN(n2953) );
  OR2_X1 U2896 ( .A1(n2664), .A2(n2663), .ZN(n3738) );
  INV_X1 U2897 ( .A(IR_REG_17__SCAN_IN), .ZN(n2338) );
  AND2_X1 U2898 ( .A1(n3852), .A2(n4329), .ZN(n2955) );
  INV_X1 U2899 ( .A(n3379), .ZN(n2934) );
  NOR2_X1 U2900 ( .A1(IR_REG_19__SCAN_IN), .A2(IR_REG_20__SCAN_IN), .ZN(n2361)
         );
  NAND2_X1 U2901 ( .A1(n3909), .A2(DATAI_1_), .ZN(n2381) );
  OR2_X1 U2902 ( .A1(n2734), .A2(n3832), .ZN(n2747) );
  NAND2_X1 U2903 ( .A1(n2779), .A2(n2778), .ZN(n2804) );
  NOR2_X1 U2904 ( .A1(n2747), .A2(n3779), .ZN(n2755) );
  INV_X1 U2905 ( .A(n4494), .ZN(n3135) );
  OAI22_X1 U2906 ( .A1(n3444), .A2(n2947), .B1(n3545), .B2(n3528), .ZN(n3512)
         );
  INV_X1 U2907 ( .A(n4061), .ZN(n4435) );
  INV_X1 U2908 ( .A(IR_REG_24__SCAN_IN), .ZN(n4940) );
  NOR2_X1 U2909 ( .A1(n2628), .A2(IR_REG_13__SCAN_IN), .ZN(n2649) );
  INV_X1 U2910 ( .A(n3303), .ZN(n2518) );
  XNOR2_X1 U2911 ( .A(n2460), .B(n2458), .ZN(n3241) );
  INV_X1 U2912 ( .A(n4212), .ZN(n4379) );
  AND2_X1 U2913 ( .A1(n2466), .A2(REG3_REG_5__SCAN_IN), .ZN(n2487) );
  NOR2_X1 U2914 ( .A1(n2593), .A2(n2592), .ZN(n2606) );
  INV_X1 U2915 ( .A(n3360), .ZN(n3318) );
  INV_X1 U2916 ( .A(n3738), .ZN(n4424) );
  OR2_X1 U2917 ( .A1(n4162), .A2(n2906), .ZN(n2855) );
  AND2_X1 U2918 ( .A1(n2686), .A2(n2685), .ZN(n4346) );
  NOR2_X1 U2919 ( .A1(n4070), .A2(n2324), .ZN(n3193) );
  INV_X1 U2920 ( .A(REG3_REG_11__SCAN_IN), .ZN(n4923) );
  INV_X1 U2921 ( .A(REG3_REG_18__SCAN_IN), .ZN(n4926) );
  INV_X1 U2922 ( .A(n4323), .ZN(n4429) );
  INV_X1 U2923 ( .A(n3002), .ZN(n3003) );
  INV_X1 U2924 ( .A(n4375), .ZN(n4245) );
  INV_X1 U2925 ( .A(n4490), .ZN(n4133) );
  INV_X1 U2926 ( .A(n3761), .ZN(n4246) );
  INV_X1 U2927 ( .A(n3575), .ZN(n3619) );
  OR2_X1 U2928 ( .A1(n2544), .A2(IR_REG_9__SCAN_IN), .ZN(n2613) );
  NAND2_X1 U2929 ( .A1(n2507), .A2(REG3_REG_7__SCAN_IN), .ZN(n2537) );
  NAND2_X1 U2930 ( .A1(n2718), .A2(REG3_REG_19__SCAN_IN), .ZN(n2734) );
  NOR2_X1 U2931 ( .A1(n2905), .A2(n4488), .ZN(n3799) );
  OR2_X1 U2932 ( .A1(n3819), .A2(n2906), .ZN(n2785) );
  INV_X1 U2933 ( .A(n4346), .ZN(n4432) );
  AND2_X1 U2934 ( .A1(n4357), .A2(n4429), .ZN(n4148) );
  INV_X1 U2935 ( .A(n4332), .ZN(n4619) );
  NAND2_X1 U2936 ( .A1(n2869), .A2(n2868), .ZN(n3352) );
  NAND2_X1 U2937 ( .A1(n4304), .A2(n4655), .ZN(n4667) );
  INV_X1 U2938 ( .A(n3352), .ZN(n3020) );
  INV_X1 U2939 ( .A(n3346), .ZN(n3107) );
  OR2_X1 U2940 ( .A1(n2512), .A2(n2347), .ZN(n2527) );
  AND2_X1 U2941 ( .A1(n3113), .A2(n3098), .ZN(n4604) );
  INV_X1 U2942 ( .A(n3799), .ZN(n3876) );
  OR2_X1 U2943 ( .A1(n2914), .A2(n2888), .ZN(n3869) );
  OAI21_X1 U2944 ( .B1(n3749), .B2(n2906), .A(n2841), .ZN(n4161) );
  NAND2_X1 U2945 ( .A1(n2785), .A2(n2784), .ZN(n4375) );
  OR2_X1 U2946 ( .A1(n2647), .A2(n2646), .ZN(n4061) );
  OR2_X1 U2947 ( .A1(n3070), .A2(n4630), .ZN(n4975) );
  INV_X1 U2948 ( .A(n4606), .ZN(n4069) );
  INV_X1 U2949 ( .A(n4638), .ZN(n4569) );
  NAND2_X1 U2950 ( .A1(n4503), .A2(n3114), .ZN(n4610) );
  INV_X1 U2951 ( .A(n4357), .ZN(n4612) );
  INV_X1 U2952 ( .A(n4357), .ZN(n4627) );
  NAND2_X1 U2953 ( .A1(n4682), .A2(n4437), .ZN(n4428) );
  NAND2_X1 U2954 ( .A1(n4675), .A2(n4437), .ZN(n4485) );
  OR2_X1 U2955 ( .A1(n3021), .A2(n3020), .ZN(n4673) );
  INV_X1 U2956 ( .A(n4628), .ZN(n4629) );
  INV_X1 U2957 ( .A(n4548), .ZN(n4640) );
  INV_X2 U2958 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  NOR2_X1 U2959 ( .A1(IR_REG_14__SCAN_IN), .A2(IR_REG_12__SCAN_IN), .ZN(n2337)
         );
  NOR2_X1 U2960 ( .A1(IR_REG_9__SCAN_IN), .A2(IR_REG_13__SCAN_IN), .ZN(n2336)
         );
  NOR2_X1 U2961 ( .A1(IR_REG_16__SCAN_IN), .A2(IR_REG_15__SCAN_IN), .ZN(n2335)
         );
  NAND4_X1 U2962 ( .A1(n2611), .A2(n2337), .A3(n2336), .A4(n2335), .ZN(n2687)
         );
  NAND2_X1 U2963 ( .A1(n2338), .A2(n2688), .ZN(n2339) );
  NOR2_X2 U2964 ( .A1(n2687), .A2(n2339), .ZN(n2340) );
  NOR2_X2 U2965 ( .A1(n2472), .A2(IR_REG_5__SCAN_IN), .ZN(n2474) );
  NOR2_X1 U2966 ( .A1(IR_REG_19__SCAN_IN), .A2(IR_REG_23__SCAN_IN), .ZN(n2343)
         );
  NAND2_X1 U2967 ( .A1(n2348), .A2(n2344), .ZN(n2350) );
  XNOR2_X2 U2968 ( .A(n2346), .B(n2345), .ZN(n2355) );
  INV_X1 U2969 ( .A(IR_REG_31__SCAN_IN), .ZN(n2347) );
  OR2_X1 U2970 ( .A1(n2348), .A2(n2347), .ZN(n2349) );
  INV_X1 U2971 ( .A(REG1_REG_1__SCAN_IN), .ZN(n2353) );
  NAND2_X2 U2972 ( .A1(n3083), .A2(n3081), .ZN(n2409) );
  INV_X1 U2973 ( .A(REG3_REG_1__SCAN_IN), .ZN(n2352) );
  OAI22_X1 U2974 ( .A1(n2446), .A2(n2353), .B1(n2409), .B2(n2352), .ZN(n2354)
         );
  INV_X1 U2975 ( .A(n2354), .ZN(n2359) );
  AND2_X2 U2976 ( .A1(n2356), .A2(n2355), .ZN(n2489) );
  NAND2_X1 U2977 ( .A1(n2489), .A2(REG0_REG_1__SCAN_IN), .ZN(n2358) );
  NAND2_X1 U2978 ( .A1(n2426), .A2(REG2_REG_1__SCAN_IN), .ZN(n2357) );
  NAND3_X2 U2979 ( .A1(n2359), .A2(n2358), .A3(n2357), .ZN(n2928) );
  NAND2_X1 U2980 ( .A1(n2884), .A2(n2883), .ZN(n2882) );
  NAND2_X1 U2981 ( .A1(n2362), .A2(IR_REG_31__SCAN_IN), .ZN(n2363) );
  MUX2_X1 U2982 ( .A(IR_REG_31__SCAN_IN), .B(n2363), .S(IR_REG_26__SCAN_IN), 
        .Z(n2364) );
  OR2_X1 U2983 ( .A1(n2365), .A2(n2347), .ZN(n2367) );
  XNOR2_X1 U2984 ( .A(n2367), .B(n2366), .ZN(n3074) );
  NOR2_X1 U2985 ( .A1(n2867), .A2(n3074), .ZN(n2368) );
  NAND2_X1 U2986 ( .A1(n2369), .A2(IR_REG_31__SCAN_IN), .ZN(n2370) );
  MUX2_X1 U2987 ( .A(IR_REG_31__SCAN_IN), .B(n2370), .S(IR_REG_21__SCAN_IN), 
        .Z(n2371) );
  INV_X1 U2988 ( .A(IR_REG_19__SCAN_IN), .ZN(n2372) );
  NAND2_X1 U2989 ( .A1(n2387), .A2(n2372), .ZN(n2373) );
  NAND2_X1 U2990 ( .A1(n2373), .A2(IR_REG_31__SCAN_IN), .ZN(n2374) );
  XNOR2_X2 U2991 ( .A(n2374), .B(n4912), .ZN(n4049) );
  INV_X1 U2992 ( .A(n2963), .ZN(n3354) );
  NAND2_X1 U2993 ( .A1(n2928), .A2(n2419), .ZN(n2384) );
  NAND2_X1 U2994 ( .A1(n3038), .A2(IR_REG_27__SCAN_IN), .ZN(n2377) );
  NAND2_X1 U2995 ( .A1(n4941), .A2(IR_REG_28__SCAN_IN), .ZN(n2376) );
  NAND3_X4 U2996 ( .A1(n2378), .A2(n2377), .A3(n2376), .ZN(n3909) );
  INV_X1 U2997 ( .A(n3909), .ZN(n2380) );
  NAND2_X1 U2998 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n2379)
         );
  XNOR2_X1 U2999 ( .A(IR_REG_1__SCAN_IN), .B(n2379), .ZN(n3116) );
  NAND2_X1 U3000 ( .A1(n2600), .A2(n2927), .ZN(n2383) );
  NAND2_X1 U3001 ( .A1(n2384), .A2(n2383), .ZN(n2388) );
  NAND2_X1 U3002 ( .A1(n4057), .A2(n4133), .ZN(n2899) );
  INV_X1 U3003 ( .A(n4489), .ZN(n2389) );
  AND2_X4 U3004 ( .A1(n2600), .A2(n4654), .ZN(n2455) );
  NAND2_X1 U3005 ( .A1(n2928), .A2(n2455), .ZN(n2391) );
  NAND2_X1 U3006 ( .A1(n2419), .A2(n3461), .ZN(n2390) );
  NAND2_X1 U3007 ( .A1(n2391), .A2(n2390), .ZN(n2406) );
  INV_X1 U3008 ( .A(REG3_REG_0__SCAN_IN), .ZN(n4906) );
  OAI22_X1 U3009 ( .A1(n2446), .A2(n4676), .B1(n2409), .B2(n4906), .ZN(n2392)
         );
  INV_X1 U3010 ( .A(n2392), .ZN(n2395) );
  NAND2_X1 U3011 ( .A1(n2489), .A2(REG0_REG_0__SCAN_IN), .ZN(n2394) );
  NAND2_X1 U3012 ( .A1(n2426), .A2(REG2_REG_0__SCAN_IN), .ZN(n2393) );
  NAND2_X1 U3013 ( .A1(n3462), .A2(n2419), .ZN(n2397) );
  MUX2_X1 U3014 ( .A(IR_REG_0__SCAN_IN), .B(DATAI_0_), .S(n3909), .Z(n2966) );
  NAND2_X1 U3015 ( .A1(n2600), .A2(n2966), .ZN(n2396) );
  AND2_X1 U3016 ( .A1(n2397), .A2(n2396), .ZN(n2402) );
  OR2_X1 U3017 ( .A1(n3070), .A2(n4676), .ZN(n2398) );
  NAND2_X1 U3018 ( .A1(n2402), .A2(n2398), .ZN(n3149) );
  NAND2_X1 U3019 ( .A1(n3462), .A2(n2455), .ZN(n2401) );
  INV_X1 U3020 ( .A(n3070), .ZN(n2399) );
  AOI22_X1 U3021 ( .A1(n2419), .A2(n2966), .B1(n2399), .B2(IR_REG_0__SCAN_IN), 
        .ZN(n2400) );
  NAND2_X1 U3022 ( .A1(n2401), .A2(n2400), .ZN(n3150) );
  NAND2_X1 U3023 ( .A1(n3149), .A2(n3150), .ZN(n2404) );
  NAND2_X1 U3024 ( .A1(n2402), .A2(n2844), .ZN(n2403) );
  NAND2_X1 U3025 ( .A1(n2404), .A2(n2403), .ZN(n3104) );
  INV_X1 U3026 ( .A(n2405), .ZN(n2407) );
  NAND2_X1 U3027 ( .A1(n2407), .A2(n2406), .ZN(n2408) );
  INV_X1 U3028 ( .A(REG3_REG_2__SCAN_IN), .ZN(n3187) );
  INV_X1 U3029 ( .A(REG1_REG_2__SCAN_IN), .ZN(n3117) );
  OAI22_X1 U3030 ( .A1(n2409), .A2(n3187), .B1(n2446), .B2(n3117), .ZN(n2410)
         );
  INV_X1 U3031 ( .A(n2410), .ZN(n2414) );
  NAND2_X1 U3032 ( .A1(n2426), .A2(REG2_REG_2__SCAN_IN), .ZN(n2412) );
  NAND2_X1 U3033 ( .A1(n2489), .A2(REG0_REG_2__SCAN_IN), .ZN(n2411) );
  NAND2_X2 U3034 ( .A1(n2414), .A2(n2413), .ZN(n4068) );
  NAND2_X1 U3035 ( .A1(n4068), .A2(n2455), .ZN(n2418) );
  NAND2_X1 U3036 ( .A1(n2419), .A2(n3167), .ZN(n2417) );
  AND2_X1 U3037 ( .A1(n2418), .A2(n2417), .ZN(n2424) );
  NAND2_X1 U3038 ( .A1(n4068), .A2(n2419), .ZN(n2421) );
  NAND2_X1 U3039 ( .A1(n2600), .A2(n3167), .ZN(n2420) );
  NAND2_X1 U3040 ( .A1(n2421), .A2(n2420), .ZN(n2422) );
  XNOR2_X1 U3041 ( .A(n2422), .B(n2844), .ZN(n2423) );
  NAND2_X1 U3042 ( .A1(n3126), .A2(n2425), .ZN(n3240) );
  NAND2_X1 U3043 ( .A1(n2757), .A2(REG1_REG_3__SCAN_IN), .ZN(n2429) );
  NAND2_X1 U3044 ( .A1(n3904), .A2(REG2_REG_3__SCAN_IN), .ZN(n2428) );
  NAND2_X1 U3045 ( .A1(n2489), .A2(REG0_REG_3__SCAN_IN), .ZN(n2427) );
  INV_X2 U3046 ( .A(n2906), .ZN(n2806) );
  INV_X1 U3047 ( .A(REG3_REG_3__SCAN_IN), .ZN(n3242) );
  NAND2_X1 U3048 ( .A1(n2806), .A2(n3242), .ZN(n2430) );
  NAND2_X2 U3049 ( .A1(n2431), .A2(n2430), .ZN(n3383) );
  NAND2_X1 U3050 ( .A1(n3383), .A2(n2419), .ZN(n2437) );
  NAND2_X1 U3051 ( .A1(n2432), .A2(IR_REG_31__SCAN_IN), .ZN(n2434) );
  NAND2_X1 U3052 ( .A1(n2434), .A2(n2433), .ZN(n2450) );
  OR2_X1 U3053 ( .A1(n2434), .A2(n2433), .ZN(n2435) );
  MUX2_X1 U3054 ( .A(n4495), .B(DATAI_3_), .S(n3909), .Z(n3258) );
  NAND2_X1 U3055 ( .A1(n2600), .A2(n3258), .ZN(n2436) );
  NAND2_X1 U3056 ( .A1(n2437), .A2(n2436), .ZN(n2438) );
  NAND2_X1 U3057 ( .A1(n3383), .A2(n2455), .ZN(n2440) );
  NAND2_X1 U3058 ( .A1(n2419), .A2(n3258), .ZN(n2439) );
  NAND2_X1 U3059 ( .A1(n2440), .A2(n2439), .ZN(n2458) );
  NAND2_X1 U3060 ( .A1(n3240), .A2(n3241), .ZN(n3215) );
  NAND2_X1 U3061 ( .A1(n3904), .A2(REG2_REG_4__SCAN_IN), .ZN(n2442) );
  NAND2_X1 U3062 ( .A1(n2489), .A2(REG0_REG_4__SCAN_IN), .ZN(n2441) );
  NAND2_X1 U3063 ( .A1(n2442), .A2(n2441), .ZN(n2449) );
  INV_X1 U3064 ( .A(n2466), .ZN(n2445) );
  INV_X1 U3065 ( .A(REG3_REG_4__SCAN_IN), .ZN(n2443) );
  NAND2_X1 U3066 ( .A1(n3242), .A2(n2443), .ZN(n2444) );
  NAND2_X1 U3067 ( .A1(n2445), .A2(n2444), .ZN(n3393) );
  INV_X1 U3068 ( .A(REG1_REG_4__SCAN_IN), .ZN(n2447) );
  OAI22_X1 U3069 ( .A1(n2409), .A2(n3393), .B1(n3908), .B2(n2447), .ZN(n2448)
         );
  NAND2_X1 U3070 ( .A1(n4067), .A2(n2419), .ZN(n2453) );
  NAND2_X1 U3071 ( .A1(n2450), .A2(IR_REG_31__SCAN_IN), .ZN(n2451) );
  XNOR2_X1 U3072 ( .A(n2451), .B(IR_REG_4__SCAN_IN), .ZN(n4494) );
  MUX2_X1 U3073 ( .A(n4494), .B(DATAI_4_), .S(n3909), .Z(n3382) );
  NAND2_X1 U3074 ( .A1(n2600), .A2(n3382), .ZN(n2452) );
  NAND2_X1 U3075 ( .A1(n2453), .A2(n2452), .ZN(n2454) );
  XNOR2_X1 U3076 ( .A(n2454), .B(n2844), .ZN(n2462) );
  NAND2_X1 U3077 ( .A1(n4067), .A2(n2455), .ZN(n2457) );
  NAND2_X1 U3078 ( .A1(n2419), .A2(n3382), .ZN(n2456) );
  NAND2_X1 U3079 ( .A1(n2457), .A2(n2456), .ZN(n2463) );
  XNOR2_X1 U3080 ( .A(n2462), .B(n2463), .ZN(n3218) );
  INV_X1 U3081 ( .A(n2458), .ZN(n2459) );
  NAND2_X1 U3082 ( .A1(n2460), .A2(n2459), .ZN(n3216) );
  AND2_X1 U3083 ( .A1(n3218), .A2(n3216), .ZN(n2461) );
  NAND2_X1 U3084 ( .A1(n3215), .A2(n2461), .ZN(n3217) );
  INV_X1 U3085 ( .A(n2462), .ZN(n2464) );
  NAND2_X1 U3086 ( .A1(n2464), .A2(n2463), .ZN(n2465) );
  NAND2_X1 U3087 ( .A1(n3217), .A2(n2465), .ZN(n3222) );
  NAND2_X1 U3088 ( .A1(n2757), .A2(REG1_REG_5__SCAN_IN), .ZN(n2471) );
  NOR2_X1 U3089 ( .A1(n2466), .A2(REG3_REG_5__SCAN_IN), .ZN(n2467) );
  NOR2_X1 U3090 ( .A1(n2487), .A2(n2467), .ZN(n3432) );
  NAND2_X1 U3091 ( .A1(n2806), .A2(n3432), .ZN(n2470) );
  NAND2_X1 U3092 ( .A1(n2489), .A2(REG0_REG_5__SCAN_IN), .ZN(n2469) );
  NAND2_X1 U3093 ( .A1(n2849), .A2(REG2_REG_5__SCAN_IN), .ZN(n2468) );
  NAND4_X1 U3094 ( .A1(n2471), .A2(n2470), .A3(n2469), .A4(n2468), .ZN(n3384)
         );
  NAND2_X1 U3095 ( .A1(n3384), .A2(n2419), .ZN(n2479) );
  NAND2_X1 U3096 ( .A1(n2472), .A2(IR_REG_31__SCAN_IN), .ZN(n2473) );
  MUX2_X1 U3097 ( .A(IR_REG_31__SCAN_IN), .B(n2473), .S(IR_REG_5__SCAN_IN), 
        .Z(n2477) );
  INV_X1 U3098 ( .A(n2475), .ZN(n2476) );
  MUX2_X1 U3099 ( .A(n3233), .B(DATAI_5_), .S(n3909), .Z(n3435) );
  NAND2_X1 U3100 ( .A1(n2600), .A2(n3435), .ZN(n2478) );
  NAND2_X1 U3101 ( .A1(n2479), .A2(n2478), .ZN(n2480) );
  XNOR2_X1 U3102 ( .A(n2480), .B(n2844), .ZN(n2483) );
  NAND2_X1 U3103 ( .A1(n3384), .A2(n2455), .ZN(n2482) );
  NAND2_X1 U3104 ( .A1(n2419), .A2(n3435), .ZN(n2481) );
  NAND2_X1 U3105 ( .A1(n2482), .A2(n2481), .ZN(n2484) );
  XNOR2_X1 U3106 ( .A(n2483), .B(n2484), .ZN(n3223) );
  INV_X1 U3107 ( .A(n2483), .ZN(n2485) );
  NAND2_X1 U3108 ( .A1(n2485), .A2(n2484), .ZN(n2486) );
  NOR2_X1 U3109 ( .A1(n2487), .A2(REG3_REG_6__SCAN_IN), .ZN(n2488) );
  NOR2_X1 U3110 ( .A1(n2507), .A2(n2488), .ZN(n3357) );
  NAND2_X1 U3111 ( .A1(n2806), .A2(n3357), .ZN(n2493) );
  NAND2_X1 U3112 ( .A1(n2757), .A2(REG1_REG_6__SCAN_IN), .ZN(n2492) );
  NAND2_X1 U3113 ( .A1(n2849), .A2(REG2_REG_6__SCAN_IN), .ZN(n2491) );
  NAND2_X1 U3114 ( .A1(n2489), .A2(REG0_REG_6__SCAN_IN), .ZN(n2490) );
  NAND4_X1 U3115 ( .A1(n2493), .A2(n2492), .A3(n2491), .A4(n2490), .ZN(n4066)
         );
  NAND2_X1 U3116 ( .A1(n4066), .A2(n2419), .ZN(n2496) );
  OR2_X1 U3117 ( .A1(n2475), .A2(n2347), .ZN(n2494) );
  XNOR2_X1 U3118 ( .A(n2494), .B(IR_REG_6__SCAN_IN), .ZN(n4493) );
  MUX2_X1 U3119 ( .A(n4493), .B(DATAI_6_), .S(n3909), .Z(n3360) );
  NAND2_X1 U3120 ( .A1(n2600), .A2(n3360), .ZN(n2495) );
  NAND2_X1 U3121 ( .A1(n2496), .A2(n2495), .ZN(n2497) );
  XNOR2_X1 U3122 ( .A(n2497), .B(n2858), .ZN(n2500) );
  NAND2_X1 U3123 ( .A1(n4066), .A2(n2455), .ZN(n2499) );
  NAND2_X1 U3124 ( .A1(n2419), .A2(n3360), .ZN(n2498) );
  NAND2_X1 U3125 ( .A1(n2499), .A2(n2498), .ZN(n2501) );
  AND2_X1 U3126 ( .A1(n2500), .A2(n2501), .ZN(n3262) );
  INV_X1 U3127 ( .A(n2500), .ZN(n2503) );
  INV_X1 U3128 ( .A(n2501), .ZN(n2502) );
  NAND2_X1 U3129 ( .A1(n2503), .A2(n2502), .ZN(n3261) );
  NAND2_X1 U3130 ( .A1(n2504), .A2(n3261), .ZN(n3302) );
  INV_X1 U3131 ( .A(n3302), .ZN(n2519) );
  NAND2_X1 U3132 ( .A1(n3904), .A2(REG2_REG_7__SCAN_IN), .ZN(n2506) );
  NAND2_X1 U3133 ( .A1(n2489), .A2(REG0_REG_7__SCAN_IN), .ZN(n2505) );
  NAND2_X1 U3134 ( .A1(n2506), .A2(n2505), .ZN(n2510) );
  OAI21_X1 U3135 ( .B1(n2507), .B2(REG3_REG_7__SCAN_IN), .A(n2537), .ZN(n3424)
         );
  INV_X1 U3136 ( .A(REG1_REG_7__SCAN_IN), .ZN(n2508) );
  OAI22_X1 U3137 ( .A1(n2906), .A2(n3424), .B1(n3908), .B2(n2508), .ZN(n2509)
         );
  NAND2_X1 U3138 ( .A1(n4065), .A2(n2419), .ZN(n2514) );
  AND2_X1 U3139 ( .A1(n2475), .A2(n2511), .ZN(n2512) );
  XNOR2_X1 U3140 ( .A(n2527), .B(IR_REG_7__SCAN_IN), .ZN(n4492) );
  MUX2_X1 U3141 ( .A(n4492), .B(DATAI_7_), .S(n3909), .Z(n3309) );
  NAND2_X1 U3142 ( .A1(n2600), .A2(n3309), .ZN(n2513) );
  NAND2_X1 U3143 ( .A1(n2514), .A2(n2513), .ZN(n2515) );
  XNOR2_X1 U3144 ( .A(n2515), .B(n2858), .ZN(n2521) );
  NAND2_X1 U3145 ( .A1(n4065), .A2(n2455), .ZN(n2517) );
  NAND2_X1 U3146 ( .A1(n2419), .A2(n3309), .ZN(n2516) );
  NAND2_X1 U3147 ( .A1(n2517), .A2(n2516), .ZN(n2520) );
  XNOR2_X1 U31480 ( .A(n2521), .B(n2520), .ZN(n3303) );
  NAND2_X1 U31490 ( .A1(n2519), .A2(n2518), .ZN(n3304) );
  NAND2_X1 U3150 ( .A1(n2521), .A2(n2520), .ZN(n2522) );
  NAND2_X1 U3151 ( .A1(n3304), .A2(n2522), .ZN(n3328) );
  NAND2_X1 U3152 ( .A1(n2757), .A2(REG1_REG_8__SCAN_IN), .ZN(n2526) );
  XNOR2_X1 U3153 ( .A(n2537), .B(REG3_REG_8__SCAN_IN), .ZN(n4611) );
  NAND2_X1 U3154 ( .A1(n2806), .A2(n4611), .ZN(n2525) );
  NAND2_X1 U3155 ( .A1(n2489), .A2(REG0_REG_8__SCAN_IN), .ZN(n2524) );
  NAND2_X1 U3156 ( .A1(n3904), .A2(REG2_REG_8__SCAN_IN), .ZN(n2523) );
  NAND2_X1 U3157 ( .A1(n3496), .A2(n2455), .ZN(n2531) );
  NAND2_X1 U3158 ( .A1(n2527), .A2(n2252), .ZN(n2528) );
  NAND2_X1 U3159 ( .A1(n2528), .A2(IR_REG_31__SCAN_IN), .ZN(n2529) );
  XNOR2_X1 U3160 ( .A(n2529), .B(IR_REG_8__SCAN_IN), .ZN(n4491) );
  MUX2_X1 U3161 ( .A(n4491), .B(DATAI_8_), .S(n3909), .Z(n3558) );
  NAND2_X1 U3162 ( .A1(n2419), .A2(n3558), .ZN(n2530) );
  NAND2_X1 U3163 ( .A1(n2531), .A2(n2530), .ZN(n3330) );
  NAND2_X1 U3164 ( .A1(n3496), .A2(n2419), .ZN(n2533) );
  NAND2_X1 U3165 ( .A1(n2600), .A2(n3558), .ZN(n2532) );
  NAND2_X1 U3166 ( .A1(n2533), .A2(n2532), .ZN(n2534) );
  XNOR2_X1 U3167 ( .A(n2534), .B(n2858), .ZN(n3329) );
  INV_X1 U3168 ( .A(n2537), .ZN(n2535) );
  AOI21_X1 U3169 ( .B1(n2535), .B2(REG3_REG_8__SCAN_IN), .A(
        REG3_REG_9__SCAN_IN), .ZN(n2538) );
  NAND2_X1 U3170 ( .A1(REG3_REG_8__SCAN_IN), .A2(REG3_REG_9__SCAN_IN), .ZN(
        n2536) );
  OR2_X1 U3171 ( .A1(n2538), .A2(n2551), .ZN(n3413) );
  INV_X1 U3172 ( .A(n3413), .ZN(n3478) );
  NAND2_X1 U3173 ( .A1(n2806), .A2(n3478), .ZN(n2542) );
  NAND2_X1 U3174 ( .A1(n2757), .A2(REG1_REG_9__SCAN_IN), .ZN(n2541) );
  NAND2_X1 U3175 ( .A1(n3905), .A2(REG0_REG_9__SCAN_IN), .ZN(n2540) );
  NAND2_X1 U3176 ( .A1(n2849), .A2(REG2_REG_9__SCAN_IN), .ZN(n2539) );
  NAND4_X1 U3177 ( .A1(n2542), .A2(n2541), .A3(n2540), .A4(n2539), .ZN(n4064)
         );
  NAND2_X1 U3178 ( .A1(n4064), .A2(n2419), .ZN(n2547) );
  NAND2_X1 U3179 ( .A1(n2475), .A2(n2688), .ZN(n2544) );
  NAND2_X1 U3180 ( .A1(n2544), .A2(IR_REG_31__SCAN_IN), .ZN(n2543) );
  MUX2_X1 U3181 ( .A(IR_REG_31__SCAN_IN), .B(n2543), .S(IR_REG_9__SCAN_IN), 
        .Z(n2545) );
  MUX2_X1 U3182 ( .A(n4110), .B(DATAI_9_), .S(n3909), .Z(n3495) );
  NAND2_X1 U3183 ( .A1(n2600), .A2(n3495), .ZN(n2546) );
  NAND2_X1 U3184 ( .A1(n2547), .A2(n2546), .ZN(n2548) );
  XNOR2_X1 U3185 ( .A(n2548), .B(n2858), .ZN(n2563) );
  NAND2_X1 U3186 ( .A1(n4064), .A2(n2455), .ZN(n2550) );
  NAND2_X1 U3187 ( .A1(n2419), .A2(n3495), .ZN(n2549) );
  NAND2_X1 U3188 ( .A1(n2550), .A2(n2549), .ZN(n2564) );
  XNOR2_X1 U3189 ( .A(n2563), .B(n2564), .ZN(n3475) );
  NAND2_X1 U3190 ( .A1(n2757), .A2(REG1_REG_10__SCAN_IN), .ZN(n2556) );
  NAND2_X1 U3191 ( .A1(n2551), .A2(REG3_REG_10__SCAN_IN), .ZN(n2572) );
  OR2_X1 U3192 ( .A1(n2551), .A2(REG3_REG_10__SCAN_IN), .ZN(n2552) );
  AND2_X1 U3193 ( .A1(n2572), .A2(n2552), .ZN(n3482) );
  NAND2_X1 U3194 ( .A1(n2806), .A2(n3482), .ZN(n2555) );
  NAND2_X1 U3195 ( .A1(n3905), .A2(REG0_REG_10__SCAN_IN), .ZN(n2554) );
  NAND2_X1 U3196 ( .A1(n2849), .A2(REG2_REG_10__SCAN_IN), .ZN(n2553) );
  NAND4_X1 U3197 ( .A1(n2556), .A2(n2555), .A3(n2554), .A4(n2553), .ZN(n4063)
         );
  NAND2_X1 U3198 ( .A1(n4063), .A2(n2419), .ZN(n2559) );
  NAND2_X1 U3199 ( .A1(n2613), .A2(IR_REG_31__SCAN_IN), .ZN(n2557) );
  XNOR2_X1 U3200 ( .A(n2557), .B(IR_REG_10__SCAN_IN), .ZN(n4112) );
  MUX2_X1 U3201 ( .A(n4112), .B(DATAI_10_), .S(n3909), .Z(n3490) );
  NAND2_X1 U3202 ( .A1(n2600), .A2(n3490), .ZN(n2558) );
  NAND2_X1 U3203 ( .A1(n2559), .A2(n2558), .ZN(n2560) );
  XNOR2_X1 U3204 ( .A(n2560), .B(n2844), .ZN(n2568) );
  NAND2_X1 U3205 ( .A1(n4063), .A2(n2455), .ZN(n2562) );
  NAND2_X1 U3206 ( .A1(n2419), .A2(n3490), .ZN(n2561) );
  NAND2_X1 U3207 ( .A1(n2562), .A2(n2561), .ZN(n2569) );
  XNOR2_X1 U3208 ( .A(n2568), .B(n2569), .ZN(n3485) );
  INV_X1 U3209 ( .A(n2563), .ZN(n2566) );
  INV_X1 U32100 ( .A(n2564), .ZN(n2565) );
  NAND2_X1 U32110 ( .A1(n2566), .A2(n2565), .ZN(n3483) );
  AND2_X1 U32120 ( .A1(n3485), .A2(n3483), .ZN(n2567) );
  NAND2_X1 U32130 ( .A1(n3473), .A2(n2567), .ZN(n3484) );
  INV_X1 U32140 ( .A(n2568), .ZN(n2570) );
  NAND2_X1 U32150 ( .A1(n2570), .A2(n2569), .ZN(n2571) );
  NAND2_X1 U32160 ( .A1(n3484), .A2(n2571), .ZN(n3540) );
  NAND2_X1 U32170 ( .A1(n2757), .A2(REG1_REG_11__SCAN_IN), .ZN(n2577) );
  NAND2_X1 U32180 ( .A1(n2572), .A2(n4923), .ZN(n2573) );
  AND2_X1 U32190 ( .A1(n2593), .A2(n2573), .ZN(n3521) );
  NAND2_X1 U32200 ( .A1(n2806), .A2(n3521), .ZN(n2576) );
  NAND2_X1 U32210 ( .A1(n3905), .A2(REG0_REG_11__SCAN_IN), .ZN(n2575) );
  NAND2_X1 U32220 ( .A1(n2849), .A2(REG2_REG_11__SCAN_IN), .ZN(n2574) );
  NAND4_X1 U32230 ( .A1(n2577), .A2(n2576), .A3(n2575), .A4(n2574), .ZN(n3620)
         );
  NAND2_X1 U32240 ( .A1(n3620), .A2(n2419), .ZN(n2582) );
  OAI21_X1 U32250 ( .B1(n2613), .B2(IR_REG_10__SCAN_IN), .A(IR_REG_31__SCAN_IN), .ZN(n2579) );
  OR2_X1 U32260 ( .A1(n2579), .A2(n2578), .ZN(n2580) );
  NAND2_X1 U32270 ( .A1(n2579), .A2(n2578), .ZN(n2597) );
  INV_X1 U32280 ( .A(DATAI_11_), .ZN(n4642) );
  MUX2_X1 U32290 ( .A(n4643), .B(n4642), .S(n3909), .Z(n3519) );
  INV_X1 U32300 ( .A(n3519), .ZN(n3547) );
  NAND2_X1 U32310 ( .A1(n2600), .A2(n3547), .ZN(n2581) );
  NAND2_X1 U32320 ( .A1(n2582), .A2(n2581), .ZN(n2583) );
  XNOR2_X1 U32330 ( .A(n2583), .B(n2844), .ZN(n2585) );
  NOR2_X1 U32340 ( .A1(n2900), .A2(n3519), .ZN(n2584) );
  AOI21_X1 U32350 ( .B1(n3620), .B2(n2455), .A(n2584), .ZN(n2586) );
  NAND2_X1 U32360 ( .A1(n2585), .A2(n2586), .ZN(n3541) );
  NAND2_X1 U32370 ( .A1(n3540), .A2(n3541), .ZN(n2589) );
  INV_X1 U32380 ( .A(n2585), .ZN(n2588) );
  INV_X1 U32390 ( .A(n2586), .ZN(n2587) );
  NAND2_X1 U32400 ( .A1(n2588), .A2(n2587), .ZN(n3542) );
  NAND2_X1 U32410 ( .A1(n2589), .A2(n3542), .ZN(n3570) );
  NAND2_X1 U32420 ( .A1(n2849), .A2(REG2_REG_12__SCAN_IN), .ZN(n2591) );
  NAND2_X1 U32430 ( .A1(n3905), .A2(REG0_REG_12__SCAN_IN), .ZN(n2590) );
  NAND2_X1 U32440 ( .A1(n2591), .A2(n2590), .ZN(n2596) );
  AND2_X1 U32450 ( .A1(n2593), .A2(n2592), .ZN(n2594) );
  OR2_X1 U32460 ( .A1(n2594), .A2(n2606), .ZN(n3595) );
  INV_X1 U32470 ( .A(REG1_REG_12__SCAN_IN), .ZN(n4935) );
  OAI22_X1 U32480 ( .A1(n2906), .A2(n3595), .B1(n3908), .B2(n4935), .ZN(n2595)
         );
  NAND2_X1 U32490 ( .A1(n3513), .A2(n2419), .ZN(n2602) );
  NAND2_X1 U32500 ( .A1(n2597), .A2(IR_REG_31__SCAN_IN), .ZN(n2598) );
  XNOR2_X1 U32510 ( .A(n2598), .B(IR_REG_12__SCAN_IN), .ZN(n4117) );
  INV_X1 U32520 ( .A(DATAI_12_), .ZN(n2599) );
  MUX2_X1 U32530 ( .A(n4641), .B(n2599), .S(n3909), .Z(n3575) );
  NAND2_X1 U32540 ( .A1(n2600), .A2(n3619), .ZN(n2601) );
  NAND2_X1 U32550 ( .A1(n2602), .A2(n2601), .ZN(n2603) );
  XNOR2_X1 U32560 ( .A(n2603), .B(n2858), .ZN(n3571) );
  NAND2_X1 U32570 ( .A1(n3513), .A2(n2455), .ZN(n2605) );
  NAND2_X1 U32580 ( .A1(n2419), .A2(n3619), .ZN(n2604) );
  NAND2_X1 U32590 ( .A1(n2605), .A2(n2604), .ZN(n3572) );
  AOI22_X1 U32600 ( .A1(n2757), .A2(REG1_REG_13__SCAN_IN), .B1(n3905), .B2(
        REG0_REG_13__SCAN_IN), .ZN(n2609) );
  NOR2_X1 U32610 ( .A1(n2606), .A2(REG3_REG_13__SCAN_IN), .ZN(n2607) );
  OR2_X1 U32620 ( .A1(n2622), .A2(n2607), .ZN(n3680) );
  INV_X1 U32630 ( .A(n3680), .ZN(n3649) );
  AOI22_X1 U32640 ( .A1(n2806), .A2(n3649), .B1(n2849), .B2(
        REG2_REG_13__SCAN_IN), .ZN(n2608) );
  INV_X1 U32650 ( .A(IR_REG_12__SCAN_IN), .ZN(n2610) );
  NAND2_X1 U32660 ( .A1(n2611), .A2(n2610), .ZN(n2612) );
  NAND2_X1 U32670 ( .A1(n2628), .A2(IR_REG_31__SCAN_IN), .ZN(n2614) );
  XNOR2_X1 U32680 ( .A(n2614), .B(IR_REG_13__SCAN_IN), .ZN(n4548) );
  INV_X1 U32690 ( .A(DATAI_13_), .ZN(n4697) );
  MUX2_X1 U32700 ( .A(n4640), .B(n4697), .S(n3909), .Z(n2984) );
  OAI22_X1 U32710 ( .A1(n3623), .A2(n2900), .B1(n2861), .B2(n2984), .ZN(n2615)
         );
  XNOR2_X1 U32720 ( .A(n2615), .B(n2858), .ZN(n2618) );
  OR2_X1 U32730 ( .A1(n3623), .A2(n2695), .ZN(n2617) );
  NAND2_X1 U32740 ( .A1(n2419), .A2(n3677), .ZN(n2616) );
  NAND2_X1 U32750 ( .A1(n2617), .A2(n2616), .ZN(n2619) );
  AND2_X1 U32760 ( .A1(n2618), .A2(n2619), .ZN(n3668) );
  INV_X1 U32770 ( .A(n2618), .ZN(n2621) );
  INV_X1 U32780 ( .A(n2619), .ZN(n2620) );
  NAND2_X1 U32790 ( .A1(n2621), .A2(n2620), .ZN(n3669) );
  NAND2_X1 U32800 ( .A1(n2757), .A2(REG1_REG_14__SCAN_IN), .ZN(n2627) );
  OR2_X1 U32810 ( .A1(n2622), .A2(REG3_REG_14__SCAN_IN), .ZN(n2623) );
  AND2_X1 U32820 ( .A1(n2644), .A2(n2623), .ZN(n3706) );
  NAND2_X1 U32830 ( .A1(n2806), .A2(n3706), .ZN(n2626) );
  NAND2_X1 U32840 ( .A1(n3905), .A2(REG0_REG_14__SCAN_IN), .ZN(n2625) );
  NAND2_X1 U32850 ( .A1(n2849), .A2(REG2_REG_14__SCAN_IN), .ZN(n2624) );
  NAND4_X1 U32860 ( .A1(n2627), .A2(n2626), .A3(n2625), .A4(n2624), .ZN(n3674)
         );
  NAND2_X1 U32870 ( .A1(n3674), .A2(n2419), .ZN(n2632) );
  OR2_X1 U32880 ( .A1(n2649), .A2(n2347), .ZN(n2629) );
  XNOR2_X1 U32890 ( .A(n2629), .B(IR_REG_14__SCAN_IN), .ZN(n4638) );
  INV_X1 U32900 ( .A(DATAI_14_), .ZN(n2630) );
  MUX2_X1 U32910 ( .A(n4569), .B(n2630), .S(n3909), .Z(n3704) );
  NAND2_X1 U32920 ( .A1(n2600), .A2(n3015), .ZN(n2631) );
  NAND2_X1 U32930 ( .A1(n2632), .A2(n2631), .ZN(n2633) );
  XNOR2_X1 U32940 ( .A(n2633), .B(n2844), .ZN(n3700) );
  NAND2_X1 U32950 ( .A1(n3674), .A2(n2455), .ZN(n2635) );
  NAND2_X1 U32960 ( .A1(n2419), .A2(n3015), .ZN(n2634) );
  NAND2_X1 U32970 ( .A1(n2635), .A2(n2634), .ZN(n3701) );
  NAND2_X1 U32980 ( .A1(n2636), .A2(n3701), .ZN(n2640) );
  INV_X1 U32990 ( .A(n3699), .ZN(n2638) );
  INV_X1 U33000 ( .A(n3700), .ZN(n2637) );
  NAND2_X1 U33010 ( .A1(n2638), .A2(n2637), .ZN(n2639) );
  NAND2_X1 U33020 ( .A1(n2640), .A2(n2639), .ZN(n2674) );
  INV_X1 U33030 ( .A(n2674), .ZN(n2657) );
  NAND2_X1 U33040 ( .A1(n3904), .A2(REG2_REG_15__SCAN_IN), .ZN(n2642) );
  NAND2_X1 U33050 ( .A1(n3905), .A2(REG0_REG_15__SCAN_IN), .ZN(n2641) );
  NAND2_X1 U33060 ( .A1(n2642), .A2(n2641), .ZN(n2647) );
  NAND2_X1 U33070 ( .A1(n2644), .A2(n2643), .ZN(n2645) );
  NAND2_X1 U33080 ( .A1(n2683), .A2(n2645), .ZN(n3884) );
  INV_X1 U33090 ( .A(REG1_REG_15__SCAN_IN), .ZN(n3716) );
  OAI22_X1 U33100 ( .A1(n2906), .A2(n3884), .B1(n3908), .B2(n3716), .ZN(n2646)
         );
  NAND2_X1 U33110 ( .A1(n4061), .A2(n2419), .ZN(n2655) );
  INV_X1 U33120 ( .A(IR_REG_14__SCAN_IN), .ZN(n2648) );
  NAND2_X1 U33130 ( .A1(n2649), .A2(n2648), .ZN(n2650) );
  NAND2_X1 U33140 ( .A1(n2650), .A2(IR_REG_31__SCAN_IN), .ZN(n2652) );
  INV_X1 U33150 ( .A(IR_REG_15__SCAN_IN), .ZN(n2651) );
  NAND2_X1 U33160 ( .A1(n2652), .A2(n2651), .ZN(n2665) );
  OR2_X1 U33170 ( .A1(n2652), .A2(n2651), .ZN(n2653) );
  MUX2_X1 U33180 ( .A(n4104), .B(DATAI_15_), .S(n3909), .Z(n3881) );
  NAND2_X1 U33190 ( .A1(n2600), .A2(n3881), .ZN(n2654) );
  NAND2_X1 U33200 ( .A1(n2655), .A2(n2654), .ZN(n2656) );
  XNOR2_X1 U33210 ( .A(n2656), .B(n2844), .ZN(n2672) );
  NAND2_X1 U33220 ( .A1(n2657), .A2(n2672), .ZN(n3794) );
  NAND2_X1 U33230 ( .A1(n4061), .A2(n2455), .ZN(n2659) );
  NAND2_X1 U33240 ( .A1(n2419), .A2(n3881), .ZN(n2658) );
  NAND2_X1 U33250 ( .A1(n2659), .A2(n2658), .ZN(n3872) );
  NAND2_X1 U33260 ( .A1(n3794), .A2(n3872), .ZN(n2675) );
  NAND2_X1 U33270 ( .A1(n2849), .A2(REG2_REG_16__SCAN_IN), .ZN(n2661) );
  NAND2_X1 U33280 ( .A1(n3905), .A2(REG0_REG_16__SCAN_IN), .ZN(n2660) );
  NAND2_X1 U33290 ( .A1(n2661), .A2(n2660), .ZN(n2664) );
  INV_X1 U33300 ( .A(REG3_REG_16__SCAN_IN), .ZN(n2681) );
  XNOR2_X1 U33310 ( .A(n2683), .B(n2681), .ZN(n3724) );
  INV_X1 U33320 ( .A(REG1_REG_16__SCAN_IN), .ZN(n2662) );
  OAI22_X1 U33330 ( .A1(n2906), .A2(n3724), .B1(n3908), .B2(n2662), .ZN(n2663)
         );
  NAND2_X1 U33340 ( .A1(n3738), .A2(n2419), .ZN(n2668) );
  NAND2_X1 U33350 ( .A1(n2665), .A2(IR_REG_31__SCAN_IN), .ZN(n2666) );
  XNOR2_X1 U33360 ( .A(n2666), .B(IR_REG_16__SCAN_IN), .ZN(n4125) );
  MUX2_X1 U33370 ( .A(n4125), .B(DATAI_16_), .S(n3909), .Z(n4430) );
  NAND2_X1 U33380 ( .A1(n2600), .A2(n4430), .ZN(n2667) );
  NAND2_X1 U33390 ( .A1(n2668), .A2(n2667), .ZN(n2669) );
  XNOR2_X1 U33400 ( .A(n2669), .B(n2844), .ZN(n2678) );
  NAND2_X1 U33410 ( .A1(n3738), .A2(n2455), .ZN(n2671) );
  NAND2_X1 U33420 ( .A1(n2419), .A2(n4430), .ZN(n2670) );
  NAND2_X1 U33430 ( .A1(n2671), .A2(n2670), .ZN(n2676) );
  XNOR2_X1 U33440 ( .A(n2678), .B(n2676), .ZN(n3797) );
  INV_X1 U33450 ( .A(n2672), .ZN(n2673) );
  NAND2_X1 U33460 ( .A1(n2674), .A2(n2673), .ZN(n3871) );
  INV_X1 U33470 ( .A(n2676), .ZN(n2677) );
  NAND2_X1 U33480 ( .A1(n2678), .A2(n2677), .ZN(n2679) );
  AOI22_X1 U33490 ( .A1(n2757), .A2(REG1_REG_17__SCAN_IN), .B1(n3905), .B2(
        REG0_REG_17__SCAN_IN), .ZN(n2686) );
  INV_X1 U33500 ( .A(REG3_REG_17__SCAN_IN), .ZN(n2680) );
  OAI21_X1 U33510 ( .B1(n2683), .B2(n2681), .A(n2680), .ZN(n2684) );
  NAND2_X1 U33520 ( .A1(REG3_REG_16__SCAN_IN), .A2(REG3_REG_17__SCAN_IN), .ZN(
        n2682) );
  AND2_X1 U3353 ( .A1(n2684), .A2(n2699), .ZN(n3811) );
  AOI22_X1 U33540 ( .A1(n2806), .A2(n3811), .B1(n2849), .B2(
        REG2_REG_17__SCAN_IN), .ZN(n2685) );
  INV_X1 U3355 ( .A(n2687), .ZN(n2689) );
  AND2_X1 U3356 ( .A1(n2689), .A2(n2688), .ZN(n2690) );
  NAND2_X1 U3357 ( .A1(n2475), .A2(n2690), .ZN(n2691) );
  NAND2_X1 U3358 ( .A1(n2691), .A2(IR_REG_31__SCAN_IN), .ZN(n2692) );
  XNOR2_X1 U3359 ( .A(n2692), .B(IR_REG_17__SCAN_IN), .ZN(n4633) );
  INV_X1 U3360 ( .A(n4633), .ZN(n4599) );
  INV_X1 U3361 ( .A(DATAI_17_), .ZN(n2693) );
  MUX2_X1 U3362 ( .A(n4599), .B(n2693), .S(n3909), .Z(n3741) );
  OAI22_X1 U3363 ( .A1(n4346), .A2(n2900), .B1(n3741), .B2(n2861), .ZN(n2694)
         );
  XNOR2_X1 U3364 ( .A(n2694), .B(n2844), .ZN(n3808) );
  OR2_X1 U3365 ( .A1(n4346), .A2(n2695), .ZN(n2697) );
  NAND2_X1 U3366 ( .A1(n2419), .A2(n4420), .ZN(n2696) );
  AND2_X1 U3367 ( .A1(n3808), .A2(n3807), .ZN(n2698) );
  NAND2_X1 U3368 ( .A1(n2757), .A2(REG1_REG_18__SCAN_IN), .ZN(n2704) );
  AND2_X1 U3369 ( .A1(n2699), .A2(n4926), .ZN(n2700) );
  NOR2_X1 U3370 ( .A1(n2718), .A2(n2700), .ZN(n4353) );
  NAND2_X1 U3371 ( .A1(n2806), .A2(n4353), .ZN(n2703) );
  NAND2_X1 U3372 ( .A1(n3905), .A2(REG0_REG_18__SCAN_IN), .ZN(n2702) );
  NAND2_X1 U3373 ( .A1(n3904), .A2(REG2_REG_18__SCAN_IN), .ZN(n2701) );
  NAND4_X1 U3374 ( .A1(n2704), .A2(n2703), .A3(n2702), .A4(n2701), .ZN(n4421)
         );
  NAND2_X1 U3375 ( .A1(n4421), .A2(n2419), .ZN(n2708) );
  NAND2_X1 U3376 ( .A1(n2360), .A2(IR_REG_31__SCAN_IN), .ZN(n2705) );
  XNOR2_X1 U3377 ( .A(n2705), .B(IR_REG_18__SCAN_IN), .ZN(n4103) );
  INV_X1 U3378 ( .A(DATAI_18_), .ZN(n2706) );
  MUX2_X1 U3379 ( .A(n4632), .B(n2706), .S(n3909), .Z(n4351) );
  INV_X1 U3380 ( .A(n4351), .ZN(n4343) );
  NAND2_X1 U3381 ( .A1(n2600), .A2(n4343), .ZN(n2707) );
  NAND2_X1 U3382 ( .A1(n2708), .A2(n2707), .ZN(n2709) );
  XNOR2_X1 U3383 ( .A(n2709), .B(n2858), .ZN(n2712) );
  NAND2_X1 U3384 ( .A1(n4421), .A2(n2455), .ZN(n2711) );
  NAND2_X1 U3385 ( .A1(n2419), .A2(n4343), .ZN(n2710) );
  NAND2_X1 U3386 ( .A1(n2711), .A2(n2710), .ZN(n2713) );
  AND2_X1 U3387 ( .A1(n2712), .A2(n2713), .ZN(n3848) );
  INV_X1 U3388 ( .A(n2712), .ZN(n2715) );
  INV_X1 U3389 ( .A(n2713), .ZN(n2714) );
  NAND2_X1 U3390 ( .A1(n2715), .A2(n2714), .ZN(n3847) );
  NAND2_X1 U3391 ( .A1(n2849), .A2(REG2_REG_19__SCAN_IN), .ZN(n2717) );
  NAND2_X1 U3392 ( .A1(n3905), .A2(REG0_REG_19__SCAN_IN), .ZN(n2716) );
  NAND2_X1 U3393 ( .A1(n2717), .A2(n2716), .ZN(n2721) );
  OR2_X1 U3394 ( .A1(n2718), .A2(REG3_REG_19__SCAN_IN), .ZN(n2719) );
  NAND2_X1 U3395 ( .A1(n2734), .A2(n2719), .ZN(n4333) );
  INV_X1 U3396 ( .A(REG1_REG_19__SCAN_IN), .ZN(n4415) );
  OAI22_X1 U3397 ( .A1(n2906), .A2(n4333), .B1(n3908), .B2(n4415), .ZN(n2720)
         );
  NAND2_X1 U3398 ( .A1(n4344), .A2(n2419), .ZN(n2723) );
  MUX2_X1 U3399 ( .A(n4490), .B(DATAI_19_), .S(n3909), .Z(n3771) );
  NAND2_X1 U3400 ( .A1(n2600), .A2(n3771), .ZN(n2722) );
  NAND2_X1 U3401 ( .A1(n2723), .A2(n2722), .ZN(n2724) );
  XNOR2_X1 U3402 ( .A(n2724), .B(n2844), .ZN(n2729) );
  NAND2_X1 U3403 ( .A1(n4344), .A2(n2455), .ZN(n2726) );
  NAND2_X1 U3404 ( .A1(n2419), .A2(n3771), .ZN(n2725) );
  NAND2_X1 U3405 ( .A1(n2726), .A2(n2725), .ZN(n2727) );
  XNOR2_X1 U3406 ( .A(n2729), .B(n2727), .ZN(n3768) );
  NAND2_X1 U3407 ( .A1(n3767), .A2(n3768), .ZN(n2731) );
  INV_X1 U3408 ( .A(n2727), .ZN(n2728) );
  NAND2_X1 U3409 ( .A1(n2729), .A2(n2728), .ZN(n2730) );
  NAND2_X1 U3410 ( .A1(n2731), .A2(n2730), .ZN(n3826) );
  NAND2_X1 U3411 ( .A1(n3904), .A2(REG2_REG_20__SCAN_IN), .ZN(n2733) );
  NAND2_X1 U3412 ( .A1(n3905), .A2(REG0_REG_20__SCAN_IN), .ZN(n2732) );
  NAND2_X1 U3413 ( .A1(n2733), .A2(n2732), .ZN(n2737) );
  INV_X1 U3414 ( .A(REG3_REG_20__SCAN_IN), .ZN(n3832) );
  NAND2_X1 U3415 ( .A1(n2734), .A2(n3832), .ZN(n2735) );
  NAND2_X1 U3416 ( .A1(n2747), .A2(n2735), .ZN(n3831) );
  INV_X1 U3417 ( .A(REG1_REG_20__SCAN_IN), .ZN(n4411) );
  OAI22_X1 U3418 ( .A1(n2906), .A2(n3831), .B1(n3908), .B2(n4411), .ZN(n2736)
         );
  NAND2_X1 U3419 ( .A1(n4280), .A2(n2419), .ZN(n2739) );
  OR2_X1 U3420 ( .A1(n4308), .A2(n2861), .ZN(n2738) );
  NAND2_X1 U3421 ( .A1(n2739), .A2(n2738), .ZN(n2740) );
  XNOR2_X1 U3422 ( .A(n2740), .B(n2858), .ZN(n2743) );
  NAND2_X1 U3423 ( .A1(n4280), .A2(n2455), .ZN(n2742) );
  OR2_X1 U3424 ( .A1(n4308), .A2(n2900), .ZN(n2741) );
  NAND2_X1 U3425 ( .A1(n2742), .A2(n2741), .ZN(n2744) );
  NAND2_X1 U3426 ( .A1(n2743), .A2(n2744), .ZN(n3827) );
  INV_X1 U3427 ( .A(n2743), .ZN(n2746) );
  INV_X1 U3428 ( .A(n2744), .ZN(n2745) );
  NAND2_X1 U3429 ( .A1(n2746), .A2(n2745), .ZN(n3829) );
  INV_X1 U3430 ( .A(REG3_REG_21__SCAN_IN), .ZN(n3779) );
  AND2_X1 U3431 ( .A1(n2747), .A2(n3779), .ZN(n2748) );
  OR2_X1 U3432 ( .A1(n2748), .A2(n2755), .ZN(n3778) );
  AOI22_X1 U3433 ( .A1(n3904), .A2(REG2_REG_21__SCAN_IN), .B1(n3905), .B2(
        REG0_REG_21__SCAN_IN), .ZN(n2750) );
  NAND2_X1 U3434 ( .A1(n2757), .A2(REG1_REG_21__SCAN_IN), .ZN(n2749) );
  OAI211_X1 U3435 ( .C1(n3778), .C2(n2906), .A(n2750), .B(n2749), .ZN(n3160)
         );
  NAND2_X1 U3436 ( .A1(n3160), .A2(n2419), .ZN(n2752) );
  NAND2_X1 U3437 ( .A1(n3909), .A2(DATAI_21_), .ZN(n4286) );
  OR2_X1 U3438 ( .A1(n2861), .A2(n4286), .ZN(n2751) );
  NAND2_X1 U3439 ( .A1(n2752), .A2(n2751), .ZN(n2753) );
  XNOR2_X1 U3440 ( .A(n2753), .B(n2844), .ZN(n3776) );
  NOR2_X1 U3441 ( .A1(n2900), .A2(n4286), .ZN(n2754) );
  AOI21_X1 U3442 ( .B1(n3160), .B2(n2455), .A(n2754), .ZN(n3775) );
  NOR2_X1 U3443 ( .A1(n2755), .A2(REG3_REG_22__SCAN_IN), .ZN(n2756) );
  OR2_X1 U3444 ( .A1(n2779), .A2(n2756), .ZN(n3842) );
  AOI22_X1 U3445 ( .A1(n2757), .A2(REG1_REG_22__SCAN_IN), .B1(n3905), .B2(
        REG0_REG_22__SCAN_IN), .ZN(n2759) );
  NAND2_X1 U3446 ( .A1(n3904), .A2(REG2_REG_22__SCAN_IN), .ZN(n2758) );
  OAI211_X1 U3447 ( .C1(n3842), .C2(n2906), .A(n2759), .B(n2758), .ZN(n4401)
         );
  NAND2_X1 U3448 ( .A1(n4401), .A2(n2419), .ZN(n2761) );
  NAND2_X1 U3449 ( .A1(n3909), .A2(DATAI_22_), .ZN(n4265) );
  OR2_X1 U3450 ( .A1(n2861), .A2(n4265), .ZN(n2760) );
  NAND2_X1 U3451 ( .A1(n2761), .A2(n2760), .ZN(n2762) );
  XNOR2_X1 U3452 ( .A(n2762), .B(n2844), .ZN(n2791) );
  NOR2_X1 U3453 ( .A1(n2900), .A2(n4265), .ZN(n2763) );
  AOI21_X1 U3454 ( .B1(n4401), .B2(n2455), .A(n2763), .ZN(n2790) );
  XNOR2_X1 U3455 ( .A(n2791), .B(n2790), .ZN(n3841) );
  INV_X1 U3456 ( .A(n3841), .ZN(n2766) );
  INV_X1 U3457 ( .A(n3776), .ZN(n2765) );
  INV_X1 U34580 ( .A(n3775), .ZN(n2764) );
  NAND2_X1 U34590 ( .A1(n2765), .A2(n2764), .ZN(n3837) );
  INV_X1 U3460 ( .A(REG3_REG_23__SCAN_IN), .ZN(n3760) );
  XNOR2_X1 U3461 ( .A(n2779), .B(n3760), .ZN(n4249) );
  NAND2_X1 U3462 ( .A1(n4249), .A2(n2806), .ZN(n2771) );
  INV_X1 U3463 ( .A(REG1_REG_23__SCAN_IN), .ZN(n4394) );
  NAND2_X1 U3464 ( .A1(n3905), .A2(REG0_REG_23__SCAN_IN), .ZN(n2768) );
  NAND2_X1 U3465 ( .A1(n3904), .A2(REG2_REG_23__SCAN_IN), .ZN(n2767) );
  OAI211_X1 U3466 ( .C1(n3908), .C2(n4394), .A(n2768), .B(n2767), .ZN(n2769)
         );
  INV_X1 U34670 ( .A(n2769), .ZN(n2770) );
  NAND2_X1 U3468 ( .A1(n4261), .A2(n2419), .ZN(n2773) );
  NAND2_X1 U34690 ( .A1(n3909), .A2(DATAI_23_), .ZN(n3761) );
  OR2_X1 U3470 ( .A1(n2861), .A2(n3761), .ZN(n2772) );
  NAND2_X1 U34710 ( .A1(n2773), .A2(n2772), .ZN(n2774) );
  XNOR2_X1 U3472 ( .A(n2774), .B(n2858), .ZN(n2789) );
  NOR2_X1 U34730 ( .A1(n2900), .A2(n3761), .ZN(n2775) );
  AOI21_X1 U3474 ( .B1(n4261), .B2(n2455), .A(n2775), .ZN(n2788) );
  INV_X1 U34750 ( .A(n2788), .ZN(n2776) );
  NAND2_X1 U3476 ( .A1(n2789), .A2(n2776), .ZN(n2798) );
  NAND2_X1 U34770 ( .A1(n2779), .A2(REG3_REG_23__SCAN_IN), .ZN(n2777) );
  INV_X1 U3478 ( .A(REG3_REG_24__SCAN_IN), .ZN(n3820) );
  NAND2_X1 U34790 ( .A1(n2777), .A2(n3820), .ZN(n2780) );
  AND2_X1 U3480 ( .A1(REG3_REG_23__SCAN_IN), .A2(REG3_REG_24__SCAN_IN), .ZN(
        n2778) );
  NAND2_X1 U34810 ( .A1(n2780), .A2(n2804), .ZN(n3819) );
  INV_X1 U3482 ( .A(REG1_REG_24__SCAN_IN), .ZN(n4949) );
  NAND2_X1 U34830 ( .A1(n3904), .A2(REG2_REG_24__SCAN_IN), .ZN(n2782) );
  NAND2_X1 U3484 ( .A1(n3905), .A2(REG0_REG_24__SCAN_IN), .ZN(n2781) );
  OAI211_X1 U34850 ( .C1(n4949), .C2(n3908), .A(n2782), .B(n2781), .ZN(n2783)
         );
  INV_X1 U3486 ( .A(n2783), .ZN(n2784) );
  NAND2_X1 U34870 ( .A1(n3909), .A2(DATAI_24_), .ZN(n4231) );
  NOR2_X1 U3488 ( .A1(n2900), .A2(n4231), .ZN(n2786) );
  AOI21_X1 U34890 ( .B1(n4375), .B2(n2455), .A(n2786), .ZN(n2800) );
  AND2_X1 U3490 ( .A1(n2798), .A2(n2800), .ZN(n2787) );
  AND2_X1 U34910 ( .A1(n3755), .A2(n2787), .ZN(n2793) );
  INV_X1 U3492 ( .A(n2787), .ZN(n2792) );
  XNOR2_X1 U34930 ( .A(n2789), .B(n2788), .ZN(n3758) );
  NAND2_X1 U3494 ( .A1(n2791), .A2(n2790), .ZN(n3759) );
  AND2_X1 U34950 ( .A1(n3758), .A2(n3759), .ZN(n3756) );
  NAND2_X1 U3496 ( .A1(n4375), .A2(n2419), .ZN(n2795) );
  OR2_X1 U34970 ( .A1(n2861), .A2(n4231), .ZN(n2794) );
  NAND2_X1 U3498 ( .A1(n2795), .A2(n2794), .ZN(n2796) );
  XNOR2_X1 U34990 ( .A(n2796), .B(n2858), .ZN(n3818) );
  NAND2_X1 U3500 ( .A1(n3816), .A2(n3818), .ZN(n2803) );
  AND2_X1 U35010 ( .A1(n3755), .A2(n2798), .ZN(n2797) );
  NAND2_X1 U3502 ( .A1(n3754), .A2(n2797), .ZN(n2802) );
  INV_X1 U35030 ( .A(n2798), .ZN(n2799) );
  NAND2_X1 U3504 ( .A1(n2803), .A2(n3815), .ZN(n3787) );
  INV_X1 U35050 ( .A(REG3_REG_25__SCAN_IN), .ZN(n3789) );
  NAND2_X1 U35060 ( .A1(n2804), .A2(n3789), .ZN(n2805) );
  NAND2_X1 U35070 ( .A1(n4213), .A2(n2806), .ZN(n2811) );
  INV_X1 U35080 ( .A(REG1_REG_25__SCAN_IN), .ZN(n4382) );
  NAND2_X1 U35090 ( .A1(n3905), .A2(REG0_REG_25__SCAN_IN), .ZN(n2808) );
  NAND2_X1 U35100 ( .A1(n2849), .A2(REG2_REG_25__SCAN_IN), .ZN(n2807) );
  OAI211_X1 U35110 ( .C1(n3908), .C2(n4382), .A(n2808), .B(n2807), .ZN(n2809)
         );
  INV_X1 U35120 ( .A(n2809), .ZN(n2810) );
  NAND2_X1 U35130 ( .A1(n4385), .A2(n2419), .ZN(n2813) );
  NAND2_X1 U35140 ( .A1(n3909), .A2(DATAI_25_), .ZN(n4216) );
  OR2_X1 U35150 ( .A1(n2861), .A2(n4216), .ZN(n2812) );
  NAND2_X1 U35160 ( .A1(n2813), .A2(n2812), .ZN(n2814) );
  XNOR2_X1 U35170 ( .A(n2814), .B(n2844), .ZN(n2817) );
  NOR2_X1 U35180 ( .A1(n2900), .A2(n4216), .ZN(n2815) );
  AOI21_X1 U35190 ( .B1(n4385), .B2(n2455), .A(n2815), .ZN(n2816) );
  NAND2_X1 U35200 ( .A1(n2817), .A2(n2816), .ZN(n3785) );
  NAND2_X1 U35210 ( .A1(n3787), .A2(n3785), .ZN(n2818) );
  OR2_X1 U35220 ( .A1(n2817), .A2(n2816), .ZN(n3786) );
  NAND2_X1 U35230 ( .A1(n2818), .A2(n3786), .ZN(n3857) );
  INV_X1 U35240 ( .A(n3857), .ZN(n2831) );
  INV_X1 U35250 ( .A(REG3_REG_26__SCAN_IN), .ZN(n3861) );
  AND2_X1 U35260 ( .A1(n2819), .A2(n3861), .ZN(n2820) );
  INV_X1 U35270 ( .A(REG1_REG_26__SCAN_IN), .ZN(n4798) );
  NAND2_X1 U35280 ( .A1(n3905), .A2(REG0_REG_26__SCAN_IN), .ZN(n2822) );
  NAND2_X1 U35290 ( .A1(n3904), .A2(REG2_REG_26__SCAN_IN), .ZN(n2821) );
  OAI211_X1 U35300 ( .C1(n3908), .C2(n4798), .A(n2822), .B(n2821), .ZN(n2823)
         );
  INV_X1 U35310 ( .A(n2823), .ZN(n2824) );
  OAI21_X1 U35320 ( .B1(n4198), .B2(n2906), .A(n2824), .ZN(n4212) );
  NAND2_X1 U35330 ( .A1(n4212), .A2(n2419), .ZN(n2826) );
  NAND2_X1 U35340 ( .A1(n3909), .A2(DATAI_26_), .ZN(n4196) );
  OR2_X1 U35350 ( .A1(n2861), .A2(n4196), .ZN(n2825) );
  NAND2_X1 U35360 ( .A1(n2826), .A2(n2825), .ZN(n2827) );
  XNOR2_X1 U35370 ( .A(n2827), .B(n2858), .ZN(n2832) );
  NAND2_X1 U35380 ( .A1(n4212), .A2(n2455), .ZN(n2829) );
  OR2_X1 U35390 ( .A1(n2900), .A2(n4196), .ZN(n2828) );
  NAND2_X1 U35400 ( .A1(n2829), .A2(n2828), .ZN(n2833) );
  AND2_X1 U35410 ( .A1(n2832), .A2(n2833), .ZN(n3859) );
  INV_X1 U35420 ( .A(n3859), .ZN(n2830) );
  INV_X1 U35430 ( .A(n2832), .ZN(n2835) );
  INV_X1 U35440 ( .A(n2833), .ZN(n2834) );
  NAND2_X1 U35450 ( .A1(n2835), .A2(n2834), .ZN(n3858) );
  NOR2_X1 U35460 ( .A1(n2836), .A2(REG3_REG_27__SCAN_IN), .ZN(n2837) );
  INV_X1 U35470 ( .A(REG1_REG_27__SCAN_IN), .ZN(n3012) );
  NAND2_X1 U35480 ( .A1(n3905), .A2(REG0_REG_27__SCAN_IN), .ZN(n2839) );
  NAND2_X1 U35490 ( .A1(n2849), .A2(REG2_REG_27__SCAN_IN), .ZN(n2838) );
  OAI211_X1 U35500 ( .C1(n3908), .C2(n3012), .A(n2839), .B(n2838), .ZN(n2840)
         );
  INV_X1 U35510 ( .A(n2840), .ZN(n2841) );
  NAND2_X1 U35520 ( .A1(n4161), .A2(n2419), .ZN(n2843) );
  AND2_X1 U35530 ( .A1(n3909), .A2(DATAI_27_), .ZN(n3975) );
  INV_X1 U35540 ( .A(n3975), .ZN(n4178) );
  OR2_X1 U35550 ( .A1(n4178), .A2(n2861), .ZN(n2842) );
  NAND2_X1 U35560 ( .A1(n2843), .A2(n2842), .ZN(n2845) );
  XNOR2_X1 U35570 ( .A(n2845), .B(n2844), .ZN(n2889) );
  NOR2_X1 U35580 ( .A1(n2900), .A2(n4178), .ZN(n2846) );
  AOI21_X1 U35590 ( .B1(n4161), .B2(n2455), .A(n2846), .ZN(n2890) );
  XNOR2_X1 U35600 ( .A(n2889), .B(n2890), .ZN(n3747) );
  NAND2_X1 U35610 ( .A1(n2847), .A2(REG3_REG_28__SCAN_IN), .ZN(n4151) );
  OR2_X1 U35620 ( .A1(n2847), .A2(REG3_REG_28__SCAN_IN), .ZN(n2848) );
  NAND2_X1 U35630 ( .A1(n4151), .A2(n2848), .ZN(n4162) );
  INV_X1 U35640 ( .A(REG1_REG_28__SCAN_IN), .ZN(n2852) );
  NAND2_X1 U35650 ( .A1(n2489), .A2(REG0_REG_28__SCAN_IN), .ZN(n2851) );
  NAND2_X1 U35660 ( .A1(n2849), .A2(REG2_REG_28__SCAN_IN), .ZN(n2850) );
  OAI211_X1 U35670 ( .C1(n3908), .C2(n2852), .A(n2851), .B(n2850), .ZN(n2853)
         );
  INV_X1 U35680 ( .A(n2853), .ZN(n2854) );
  NAND2_X1 U35690 ( .A1(n4174), .A2(n2455), .ZN(n2857) );
  NAND2_X1 U35700 ( .A1(n3909), .A2(DATAI_28_), .ZN(n4166) );
  OR2_X1 U35710 ( .A1(n2900), .A2(n4166), .ZN(n2856) );
  NAND2_X1 U35720 ( .A1(n2857), .A2(n2856), .ZN(n2859) );
  XNOR2_X1 U35730 ( .A(n2859), .B(n2858), .ZN(n2863) );
  NAND2_X1 U35740 ( .A1(n4174), .A2(n2419), .ZN(n2860) );
  OAI21_X1 U35750 ( .B1(n2861), .B2(n4166), .A(n2860), .ZN(n2862) );
  XNOR2_X1 U35760 ( .A(n2863), .B(n2862), .ZN(n2922) );
  INV_X1 U35770 ( .A(n2922), .ZN(n2893) );
  NAND2_X1 U35780 ( .A1(n2864), .A2(n3074), .ZN(n2865) );
  MUX2_X1 U35790 ( .A(n2864), .B(n2865), .S(B_REG_SCAN_IN), .Z(n2866) );
  NAND2_X1 U35800 ( .A1(n2867), .A2(n3074), .ZN(n3347) );
  OAI21_X1 U35810 ( .B1(n3087), .B2(D_REG_1__SCAN_IN), .A(n3347), .ZN(n3011)
         );
  INV_X1 U3582 ( .A(n3011), .ZN(n2881) );
  INV_X1 U3583 ( .A(D_REG_0__SCAN_IN), .ZN(n3091) );
  NAND2_X1 U3584 ( .A1(n2880), .A2(n3091), .ZN(n2869) );
  NAND2_X1 U3585 ( .A1(n2864), .A2(n2867), .ZN(n2868) );
  NOR4_X1 U3586 ( .A1(D_REG_2__SCAN_IN), .A2(D_REG_5__SCAN_IN), .A3(
        D_REG_7__SCAN_IN), .A4(D_REG_16__SCAN_IN), .ZN(n2871) );
  NOR4_X1 U3587 ( .A1(D_REG_20__SCAN_IN), .A2(D_REG_28__SCAN_IN), .A3(
        D_REG_27__SCAN_IN), .A4(D_REG_9__SCAN_IN), .ZN(n2870) );
  INV_X1 U3588 ( .A(D_REG_17__SCAN_IN), .ZN(n4749) );
  INV_X1 U3589 ( .A(D_REG_21__SCAN_IN), .ZN(n4753) );
  NAND4_X1 U3590 ( .A1(n2871), .A2(n2870), .A3(n4749), .A4(n4753), .ZN(n4927)
         );
  NOR4_X1 U3591 ( .A1(D_REG_24__SCAN_IN), .A2(D_REG_22__SCAN_IN), .A3(
        D_REG_11__SCAN_IN), .A4(D_REG_4__SCAN_IN), .ZN(n2875) );
  NOR4_X1 U3592 ( .A1(D_REG_3__SCAN_IN), .A2(D_REG_6__SCAN_IN), .A3(
        D_REG_10__SCAN_IN), .A4(D_REG_18__SCAN_IN), .ZN(n2874) );
  NOR4_X1 U3593 ( .A1(D_REG_14__SCAN_IN), .A2(D_REG_15__SCAN_IN), .A3(
        D_REG_23__SCAN_IN), .A4(D_REG_25__SCAN_IN), .ZN(n2873) );
  NOR4_X1 U3594 ( .A1(D_REG_8__SCAN_IN), .A2(D_REG_12__SCAN_IN), .A3(
        D_REG_13__SCAN_IN), .A4(D_REG_19__SCAN_IN), .ZN(n2872) );
  NAND4_X1 U3595 ( .A1(n2875), .A2(n2874), .A3(n2873), .A4(n2872), .ZN(n2876)
         );
  NOR2_X1 U3596 ( .A1(n4927), .A2(n2876), .ZN(n2878) );
  NOR4_X1 U3597 ( .A1(D_REG_26__SCAN_IN), .A2(D_REG_29__SCAN_IN), .A3(
        D_REG_30__SCAN_IN), .A4(D_REG_31__SCAN_IN), .ZN(n2877) );
  NAND2_X1 U3598 ( .A1(n2878), .A2(n2877), .ZN(n2879) );
  NAND2_X1 U3599 ( .A1(n2880), .A2(n2879), .ZN(n3349) );
  NAND3_X1 U3600 ( .A1(n2881), .A2(n3020), .A3(n3349), .ZN(n2914) );
  OR2_X1 U3601 ( .A1(n2884), .A2(n2883), .ZN(n2885) );
  NAND2_X1 U3602 ( .A1(n2882), .A2(n2885), .ZN(n3095) );
  INV_X1 U3603 ( .A(n3096), .ZN(n2887) );
  NAND2_X1 U3604 ( .A1(n4049), .A2(n4133), .ZN(n2896) );
  NAND2_X1 U3605 ( .A1(n3368), .A2(n2896), .ZN(n2886) );
  NAND2_X1 U3606 ( .A1(n2887), .A2(n2886), .ZN(n2894) );
  OR2_X1 U3607 ( .A1(n3346), .A2(n2894), .ZN(n2888) );
  NOR2_X1 U3608 ( .A1(n2893), .A2(n3869), .ZN(n2920) );
  INV_X1 U3609 ( .A(n2889), .ZN(n2892) );
  INV_X1 U3610 ( .A(n2890), .ZN(n2891) );
  INV_X1 U3611 ( .A(n4049), .ZN(n3078) );
  NAND2_X1 U3612 ( .A1(n3368), .A2(n3078), .ZN(n4323) );
  NAND2_X1 U3613 ( .A1(n2894), .A2(n4323), .ZN(n2895) );
  NAND2_X1 U3614 ( .A1(n2914), .A2(n2895), .ZN(n2897) );
  NAND2_X1 U3615 ( .A1(n3096), .A2(n2896), .ZN(n3348) );
  NAND2_X1 U3616 ( .A1(n2897), .A2(n3348), .ZN(n3105) );
  NAND2_X1 U3617 ( .A1(n3070), .A2(n3095), .ZN(n2898) );
  OAI21_X1 U3618 ( .B1(n3105), .B2(n2898), .A(STATE_REG_SCAN_IN), .ZN(n2901)
         );
  NAND2_X1 U3619 ( .A1(n2914), .A2(n2180), .ZN(n3106) );
  INV_X1 U3620 ( .A(n2914), .ZN(n2902) );
  NAND2_X1 U3621 ( .A1(n2902), .A2(n2180), .ZN(n2905) );
  OAI21_X1 U3622 ( .B1(n2375), .B2(IR_REG_27__SCAN_IN), .A(IR_REG_31__SCAN_IN), 
        .ZN(n2904) );
  XNOR2_X1 U3623 ( .A(n2904), .B(n2903), .ZN(n3114) );
  INV_X1 U3624 ( .A(n3114), .ZN(n4488) );
  OR2_X1 U3625 ( .A1(n4151), .A2(n2906), .ZN(n2911) );
  INV_X1 U3626 ( .A(REG1_REG_29__SCAN_IN), .ZN(n3065) );
  NAND2_X1 U3627 ( .A1(n3904), .A2(REG2_REG_29__SCAN_IN), .ZN(n2908) );
  NAND2_X1 U3628 ( .A1(n3905), .A2(REG0_REG_29__SCAN_IN), .ZN(n2907) );
  OAI211_X1 U3629 ( .C1(n3908), .C2(n3065), .A(n2908), .B(n2907), .ZN(n2909)
         );
  INV_X1 U3630 ( .A(n2909), .ZN(n2910) );
  NAND2_X1 U3631 ( .A1(n2911), .A2(n2910), .ZN(n4160) );
  AOI22_X1 U3632 ( .A1(n4161), .A2(n3798), .B1(n3799), .B2(n4160), .ZN(n2916)
         );
  NAND2_X1 U3633 ( .A1(n3107), .A2(n4429), .ZN(n2913) );
  AND2_X1 U3634 ( .A1(n4049), .A2(n4490), .ZN(n3371) );
  NAND2_X1 U3635 ( .A1(n3371), .A2(n2912), .ZN(n4655) );
  OAI21_X2 U3636 ( .B1(n2914), .B2(n2913), .A(n4332), .ZN(n3880) );
  INV_X1 U3637 ( .A(n4166), .ZN(n3044) );
  AOI22_X1 U3638 ( .A1(n3880), .A2(n3044), .B1(REG3_REG_28__SCAN_IN), .B2(
        U3149), .ZN(n2915) );
  OAI211_X1 U3639 ( .C1(n3885), .C2(n4162), .A(n2916), .B(n2915), .ZN(n2917)
         );
  INV_X1 U3640 ( .A(n2917), .ZN(n2918) );
  AOI21_X1 U3641 ( .B1(n2921), .B2(n2920), .A(n2919), .ZN(n2925) );
  NAND2_X1 U3642 ( .A1(n2923), .A2(n2171), .ZN(n2924) );
  NAND2_X1 U3643 ( .A1(n2925), .A2(n2924), .ZN(U3217) );
  XNOR2_X1 U3644 ( .A(n4161), .B(n3975), .ZN(n3945) );
  INV_X1 U3645 ( .A(n2928), .ZN(n2926) );
  NAND2_X1 U3646 ( .A1(n2926), .A2(n2927), .ZN(n2968) );
  INV_X1 U3647 ( .A(n2927), .ZN(n3013) );
  NAND2_X1 U3648 ( .A1(n3013), .A2(n2928), .ZN(n3977) );
  NAND2_X1 U3649 ( .A1(n2928), .A2(n3461), .ZN(n2929) );
  INV_X1 U3650 ( .A(n3167), .ZN(n3173) );
  NAND2_X1 U3651 ( .A1(n4068), .A2(n3173), .ZN(n3984) );
  NAND2_X1 U3652 ( .A1(n2930), .A2(n3173), .ZN(n2931) );
  NAND2_X1 U3653 ( .A1(n3178), .A2(n2931), .ZN(n3248) );
  NAND2_X1 U3654 ( .A1(n3383), .A2(n3258), .ZN(n2932) );
  NAND2_X1 U3655 ( .A1(n3296), .A2(n3382), .ZN(n3987) );
  INV_X1 U3656 ( .A(n3382), .ZN(n3391) );
  NAND2_X1 U3657 ( .A1(n4067), .A2(n3391), .ZN(n3990) );
  NAND2_X1 U3658 ( .A1(n4067), .A2(n3382), .ZN(n2935) );
  NAND2_X1 U3659 ( .A1(n3377), .A2(n2935), .ZN(n3291) );
  OR2_X1 U3660 ( .A1(n3384), .A2(n3435), .ZN(n2936) );
  NAND2_X1 U3661 ( .A1(n3291), .A2(n2936), .ZN(n2938) );
  NAND2_X1 U3662 ( .A1(n3384), .A2(n3435), .ZN(n2937) );
  NAND2_X1 U3663 ( .A1(n2938), .A2(n2937), .ZN(n3312) );
  AND2_X1 U3664 ( .A1(n4066), .A2(n3360), .ZN(n2940) );
  INV_X1 U3665 ( .A(n4065), .ZN(n3313) );
  NAND2_X1 U3666 ( .A1(n3313), .A2(n3309), .ZN(n3993) );
  NAND2_X1 U3667 ( .A1(n4065), .A2(n3422), .ZN(n3995) );
  OR2_X1 U3668 ( .A1(n3968), .A2(n2328), .ZN(n3407) );
  OR2_X1 U3669 ( .A1(n3407), .A2(n2159), .ZN(n2945) );
  NAND2_X1 U3670 ( .A1(n4065), .A2(n3309), .ZN(n3555) );
  NAND2_X1 U3671 ( .A1(n3496), .A2(n3558), .ZN(n2941) );
  AND2_X1 U3672 ( .A1(n3555), .A2(n2941), .ZN(n2942) );
  AND2_X1 U3673 ( .A1(n2162), .A2(n3408), .ZN(n2943) );
  OR2_X1 U3674 ( .A1(n2159), .A2(n2943), .ZN(n2944) );
  OAI21_X1 U3675 ( .B1(n3406), .B2(n2945), .A(n2944), .ZN(n2946) );
  INV_X1 U3676 ( .A(n2946), .ZN(n3444) );
  NOR2_X1 U3677 ( .A1(n4063), .A2(n3490), .ZN(n2947) );
  INV_X1 U3678 ( .A(n4063), .ZN(n3545) );
  OR2_X1 U3679 ( .A1(n3620), .A2(n3519), .ZN(n3602) );
  NAND2_X1 U3680 ( .A1(n3620), .A2(n3519), .ZN(n2982) );
  OR2_X1 U3681 ( .A1(n3620), .A2(n3547), .ZN(n2948) );
  INV_X1 U3682 ( .A(n3634), .ZN(n2950) );
  NAND2_X1 U3683 ( .A1(n3623), .A2(n2984), .ZN(n2949) );
  OR2_X1 U3684 ( .A1(n3674), .A2(n3704), .ZN(n3886) );
  NAND2_X1 U3685 ( .A1(n3674), .A2(n3704), .ZN(n3887) );
  NAND2_X1 U3686 ( .A1(n3886), .A2(n3887), .ZN(n3582) );
  NAND2_X1 U3687 ( .A1(n4424), .A2(n4430), .ZN(n4027) );
  INV_X1 U3688 ( .A(n4430), .ZN(n3801) );
  NAND2_X1 U3689 ( .A1(n3738), .A2(n3801), .ZN(n4023) );
  NAND2_X1 U3690 ( .A1(n4027), .A2(n4023), .ZN(n3720) );
  NAND2_X1 U3691 ( .A1(n3721), .A2(n3720), .ZN(n3719) );
  NAND2_X1 U3692 ( .A1(n3719), .A2(n2951), .ZN(n3735) );
  NAND2_X1 U3693 ( .A1(n4346), .A2(n3741), .ZN(n2952) );
  AOI21_X1 U3694 ( .B1(n3735), .B2(n2952), .A(n2323), .ZN(n4339) );
  OR2_X1 U3695 ( .A1(n4421), .A2(n4351), .ZN(n4318) );
  NAND2_X1 U3696 ( .A1(n4421), .A2(n4351), .ZN(n4319) );
  NAND2_X1 U3697 ( .A1(n4318), .A2(n4319), .ZN(n4342) );
  NAND2_X1 U3698 ( .A1(n4339), .A2(n4342), .ZN(n4338) );
  NAND2_X1 U3699 ( .A1(n4338), .A2(n2954), .ZN(n4315) );
  NAND2_X1 U3700 ( .A1(n4344), .A2(n3771), .ZN(n2956) );
  INV_X1 U3701 ( .A(n3771), .ZN(n4329) );
  INV_X1 U3702 ( .A(n3160), .ZN(n4300) );
  NOR2_X1 U3703 ( .A1(n4300), .A2(n4286), .ZN(n2957) );
  INV_X1 U3704 ( .A(n4286), .ZN(n4400) );
  INV_X1 U3705 ( .A(n4256), .ZN(n4254) );
  OR2_X1 U3706 ( .A1(n4401), .A2(n4265), .ZN(n4239) );
  NAND2_X1 U3707 ( .A1(n4401), .A2(n4265), .ZN(n2997) );
  NAND2_X1 U3708 ( .A1(n4239), .A2(n2997), .ZN(n4259) );
  NAND2_X1 U3709 ( .A1(n4254), .A2(n4259), .ZN(n2958) );
  INV_X1 U3710 ( .A(n4401), .ZN(n3780) );
  NAND2_X1 U3711 ( .A1(n2958), .A2(n2329), .ZN(n4236) );
  INV_X1 U3712 ( .A(n4261), .ZN(n4388) );
  NAND2_X1 U3713 ( .A1(n4388), .A2(n3761), .ZN(n2960) );
  AOI21_X1 U3714 ( .B1(n4236), .B2(n2960), .A(n2959), .ZN(n4224) );
  INV_X1 U3715 ( .A(n4231), .ZN(n4384) );
  NAND2_X1 U3716 ( .A1(n4375), .A2(n4384), .ZN(n2961) );
  NOR2_X1 U3717 ( .A1(n4379), .A2(n4196), .ZN(n2962) );
  XOR2_X1 U3718 ( .A(n3945), .B(n3027), .Z(n4172) );
  XNOR2_X1 U3719 ( .A(n2963), .B(n4057), .ZN(n2964) );
  NAND2_X1 U3720 ( .A1(n2964), .A2(n4133), .ZN(n4304) );
  INV_X1 U3721 ( .A(n4174), .ZN(n4146) );
  NAND2_X1 U3722 ( .A1(n3096), .A2(n3114), .ZN(n4378) );
  INV_X1 U3723 ( .A(n3462), .ZN(n2967) );
  NAND2_X1 U3724 ( .A1(n2967), .A2(n2966), .ZN(n3976) );
  OR2_X1 U3725 ( .A1(n2965), .A2(n3976), .ZN(n2969) );
  NAND2_X1 U3726 ( .A1(n2969), .A2(n3980), .ZN(n3170) );
  NAND2_X1 U3727 ( .A1(n3170), .A2(n3967), .ZN(n3169) );
  NAND2_X1 U3728 ( .A1(n3169), .A2(n3981), .ZN(n3250) );
  INV_X1 U3729 ( .A(n3258), .ZN(n3014) );
  OR2_X1 U3730 ( .A1(n3383), .A2(n3014), .ZN(n3986) );
  NAND2_X1 U3731 ( .A1(n3383), .A2(n3014), .ZN(n3983) );
  NAND2_X1 U3732 ( .A1(n3986), .A2(n3983), .ZN(n3956) );
  INV_X1 U3733 ( .A(n3956), .ZN(n3249) );
  NAND2_X1 U3734 ( .A1(n3250), .A2(n3249), .ZN(n2971) );
  NAND2_X1 U3735 ( .A1(n2971), .A2(n3986), .ZN(n3381) );
  INV_X1 U3736 ( .A(n3987), .ZN(n2972) );
  NAND2_X1 U3737 ( .A1(n2973), .A2(n3990), .ZN(n3293) );
  INV_X1 U3738 ( .A(n3435), .ZN(n2974) );
  AND2_X1 U3739 ( .A1(n3384), .A2(n2974), .ZN(n3292) );
  OR2_X1 U3740 ( .A1(n3384), .A2(n2974), .ZN(n4005) );
  OAI21_X1 U3741 ( .B1(n3293), .B2(n3292), .A(n4005), .ZN(n3314) );
  NAND2_X1 U3742 ( .A1(n4066), .A2(n3318), .ZN(n4004) );
  NAND2_X1 U3743 ( .A1(n3314), .A2(n4004), .ZN(n2975) );
  OR2_X1 U3744 ( .A1(n4066), .A2(n3318), .ZN(n3992) );
  NAND2_X1 U3745 ( .A1(n2975), .A2(n3992), .ZN(n3418) );
  INV_X1 U3746 ( .A(n3993), .ZN(n2976) );
  NAND2_X1 U3747 ( .A1(n2977), .A2(n3995), .ZN(n3557) );
  INV_X1 U3748 ( .A(n3558), .ZN(n3553) );
  OR2_X1 U3749 ( .A1(n3496), .A2(n3553), .ZN(n3997) );
  NAND2_X1 U3750 ( .A1(n3557), .A2(n3997), .ZN(n2978) );
  NAND2_X1 U3751 ( .A1(n3496), .A2(n3553), .ZN(n3996) );
  NAND2_X1 U3752 ( .A1(n2978), .A2(n3996), .ZN(n3404) );
  INV_X1 U3753 ( .A(n3495), .ZN(n2979) );
  AND2_X1 U3754 ( .A1(n4064), .A2(n2979), .ZN(n4006) );
  OR2_X1 U3755 ( .A1(n4064), .A2(n2979), .ZN(n3998) );
  NAND2_X1 U3756 ( .A1(n2980), .A2(n3998), .ZN(n3446) );
  NAND2_X1 U3757 ( .A1(n4063), .A2(n3528), .ZN(n4012) );
  NAND2_X1 U3758 ( .A1(n3446), .A2(n4012), .ZN(n2981) );
  OR2_X1 U3759 ( .A1(n4063), .A2(n3528), .ZN(n4009) );
  NAND2_X1 U3760 ( .A1(n2981), .A2(n4009), .ZN(n3509) );
  NAND2_X1 U3761 ( .A1(n3513), .A2(n3575), .ZN(n3639) );
  NAND2_X1 U3762 ( .A1(n4062), .A2(n2984), .ZN(n3635) );
  NAND2_X1 U3763 ( .A1(n3639), .A2(n3635), .ZN(n2983) );
  INV_X1 U3764 ( .A(n2982), .ZN(n3601) );
  NOR2_X1 U3765 ( .A1(n2983), .A2(n3601), .ZN(n4013) );
  NAND2_X1 U3766 ( .A1(n3509), .A2(n4013), .ZN(n2987) );
  NAND2_X1 U3767 ( .A1(n3675), .A2(n3619), .ZN(n3638) );
  NAND2_X1 U3768 ( .A1(n3638), .A2(n3602), .ZN(n2986) );
  INV_X1 U3769 ( .A(n2983), .ZN(n2985) );
  NOR2_X1 U3770 ( .A1(n4062), .A2(n2984), .ZN(n3637) );
  AOI21_X1 U3771 ( .B1(n2986), .B2(n2985), .A(n3637), .ZN(n4022) );
  NAND2_X1 U3772 ( .A1(n2987), .A2(n4022), .ZN(n3890) );
  INV_X1 U3773 ( .A(n3582), .ZN(n3935) );
  NAND2_X1 U3774 ( .A1(n3890), .A2(n3935), .ZN(n2988) );
  NAND2_X1 U3775 ( .A1(n2988), .A2(n3886), .ZN(n3654) );
  NAND2_X1 U3776 ( .A1(n4435), .A2(n3881), .ZN(n3889) );
  NAND2_X1 U3777 ( .A1(n4061), .A2(n3662), .ZN(n3888) );
  NAND2_X1 U3778 ( .A1(n3889), .A2(n3888), .ZN(n3933) );
  NAND2_X1 U3779 ( .A1(n3655), .A2(n3888), .ZN(n3728) );
  INV_X1 U3780 ( .A(n3720), .ZN(n3936) );
  NAND2_X1 U3781 ( .A1(n3728), .A2(n3936), .ZN(n3727) );
  NAND2_X1 U3782 ( .A1(n3727), .A2(n4023), .ZN(n3733) );
  AND2_X1 U3783 ( .A1(n4432), .A2(n3741), .ZN(n3891) );
  NOR2_X1 U3784 ( .A1(n3733), .A2(n3891), .ZN(n2989) );
  INV_X1 U3785 ( .A(n2989), .ZN(n4317) );
  NAND2_X1 U3786 ( .A1(n4344), .A2(n4329), .ZN(n3940) );
  AND2_X1 U3787 ( .A1(n4319), .A2(n3940), .ZN(n4293) );
  NAND2_X1 U3788 ( .A1(n4280), .A2(n4308), .ZN(n2990) );
  NAND2_X1 U3789 ( .A1(n4293), .A2(n2990), .ZN(n3892) );
  OR2_X1 U3790 ( .A1(n4432), .A2(n3741), .ZN(n4316) );
  NAND2_X1 U3791 ( .A1(n4318), .A2(n4316), .ZN(n2991) );
  NAND2_X1 U3792 ( .A1(n4293), .A2(n2991), .ZN(n2992) );
  NAND2_X1 U3793 ( .A1(n3852), .A2(n3771), .ZN(n3941) );
  NAND2_X1 U3794 ( .A1(n2992), .A2(n3941), .ZN(n2994) );
  NAND2_X1 U3795 ( .A1(n2994), .A2(n4298), .ZN(n2993) );
  NAND2_X1 U3796 ( .A1(n2993), .A2(n4280), .ZN(n2996) );
  INV_X1 U3797 ( .A(n2994), .ZN(n4294) );
  NAND2_X1 U3798 ( .A1(n4294), .A2(n4308), .ZN(n2995) );
  NAND2_X1 U3799 ( .A1(n2996), .A2(n2995), .ZN(n3895) );
  OR2_X1 U3800 ( .A1(n3160), .A2(n4286), .ZN(n4237) );
  NAND2_X1 U3801 ( .A1(n4239), .A2(n4237), .ZN(n4032) );
  NAND2_X1 U3802 ( .A1(n4261), .A2(n3761), .ZN(n3931) );
  AND2_X1 U3803 ( .A1(n3931), .A2(n2997), .ZN(n4038) );
  AND2_X1 U3804 ( .A1(n3160), .A2(n4286), .ZN(n3953) );
  NAND2_X1 U3805 ( .A1(n4239), .A2(n3953), .ZN(n2998) );
  AND2_X1 U3806 ( .A1(n4038), .A2(n2998), .ZN(n3897) );
  OAI21_X1 U3807 ( .B1(n4273), .B2(n4032), .A(n3897), .ZN(n2999) );
  OR2_X1 U3808 ( .A1(n4261), .A2(n3761), .ZN(n3932) );
  NAND2_X1 U3809 ( .A1(n2999), .A2(n3932), .ZN(n4222) );
  NOR2_X1 U3810 ( .A1(n4375), .A2(n4231), .ZN(n3939) );
  OR2_X2 U3811 ( .A1(n4222), .A2(n3939), .ZN(n4204) );
  OR2_X1 U3812 ( .A1(n4212), .A2(n4196), .ZN(n3000) );
  OR2_X1 U3813 ( .A1(n4385), .A2(n4216), .ZN(n4185) );
  NAND2_X1 U3814 ( .A1(n3000), .A2(n4185), .ZN(n4036) );
  NAND2_X1 U3815 ( .A1(n4385), .A2(n4216), .ZN(n3937) );
  NAND2_X1 U3816 ( .A1(n4375), .A2(n4231), .ZN(n4203) );
  AND2_X1 U3817 ( .A1(n3937), .A2(n4203), .ZN(n4187) );
  NAND2_X1 U3818 ( .A1(n4212), .A2(n4196), .ZN(n3915) );
  OAI21_X1 U3819 ( .B1(n4036), .B2(n4187), .A(n3915), .ZN(n4041) );
  INV_X1 U3820 ( .A(n4041), .ZN(n3001) );
  NAND2_X1 U3821 ( .A1(n3003), .A2(n3945), .ZN(n3032) );
  OAI21_X1 U3822 ( .B1(n3945), .B2(n3003), .A(n3032), .ZN(n3005) );
  NAND2_X1 U3823 ( .A1(n4057), .A2(n4490), .ZN(n3004) );
  NAND2_X1 U3824 ( .A1(n4489), .A2(n3078), .ZN(n3922) );
  NAND2_X2 U3825 ( .A1(n3004), .A2(n3922), .ZN(n4348) );
  NAND2_X1 U3826 ( .A1(n3005), .A2(n4348), .ZN(n4183) );
  AOI22_X1 U3827 ( .A1(n4212), .A2(n4374), .B1(n3975), .B2(n4429), .ZN(n3006)
         );
  OAI211_X1 U3828 ( .C1(n4146), .C2(n4378), .A(n4183), .B(n3006), .ZN(n3007)
         );
  AOI21_X1 U3829 ( .B1(n4172), .B2(n4667), .A(n3007), .ZN(n3022) );
  NAND2_X1 U3830 ( .A1(n3008), .A2(n3348), .ZN(n3009) );
  NOR2_X1 U3831 ( .A1(n3346), .A2(n3009), .ZN(n3010) );
  NAND3_X1 U3832 ( .A1(n3011), .A2(n3010), .A3(n3349), .ZN(n3021) );
  MUX2_X1 U3833 ( .A(n3012), .B(n3022), .S(n4682), .Z(n3019) );
  INV_X1 U3834 ( .A(n2966), .ZN(n3369) );
  NAND2_X1 U3835 ( .A1(n3013), .A2(n3369), .ZN(n3457) );
  NAND2_X1 U3836 ( .A1(n3166), .A2(n3014), .ZN(n3256) );
  NAND2_X1 U3837 ( .A1(n3016), .A2(n3975), .ZN(n3017) );
  NAND2_X1 U3838 ( .A1(n3058), .A2(n3017), .ZN(n4173) );
  NAND2_X1 U3839 ( .A1(n3019), .A2(n3018), .ZN(U3545) );
  INV_X1 U3840 ( .A(REG0_REG_27__SCAN_IN), .ZN(n3023) );
  MUX2_X1 U3841 ( .A(n3023), .B(n3022), .S(n4675), .Z(n3025) );
  NAND2_X1 U3842 ( .A1(n3025), .A2(n3024), .ZN(U3513) );
  NOR2_X1 U3843 ( .A1(n4161), .A2(n3975), .ZN(n3026) );
  INV_X1 U3844 ( .A(n4161), .ZN(n4195) );
  OAI22_X1 U3845 ( .A1(n3027), .A2(n3026), .B1(n4195), .B2(n4178), .ZN(n3049)
         );
  NOR2_X1 U3846 ( .A1(n4174), .A2(n4166), .ZN(n3903) );
  INV_X1 U3847 ( .A(n3903), .ZN(n3028) );
  NAND2_X1 U3848 ( .A1(n4174), .A2(n4166), .ZN(n3914) );
  NAND2_X1 U3849 ( .A1(n3028), .A2(n3914), .ZN(n3952) );
  NAND2_X1 U3850 ( .A1(n3049), .A2(n3952), .ZN(n3029) );
  NAND2_X1 U3851 ( .A1(n3029), .A2(n2333), .ZN(n3030) );
  NAND2_X1 U3852 ( .A1(n3909), .A2(DATAI_29_), .ZN(n3912) );
  XOR2_X1 U3853 ( .A(n3912), .B(n4160), .Z(n3946) );
  XNOR2_X1 U3854 ( .A(n3030), .B(n3946), .ZN(n4143) );
  NOR2_X1 U3855 ( .A1(n4161), .A2(n4178), .ZN(n3902) );
  INV_X1 U3856 ( .A(n3902), .ZN(n3031) );
  NAND2_X1 U3857 ( .A1(n3032), .A2(n3031), .ZN(n3051) );
  AOI21_X1 U3858 ( .B1(n3051), .B2(n3914), .A(n3903), .ZN(n3034) );
  INV_X1 U3859 ( .A(n3946), .ZN(n3033) );
  XNOR2_X1 U3860 ( .A(n3034), .B(n3033), .ZN(n3041) );
  INV_X1 U3861 ( .A(REG1_REG_30__SCAN_IN), .ZN(n3037) );
  NAND2_X1 U3862 ( .A1(n3904), .A2(REG2_REG_30__SCAN_IN), .ZN(n3036) );
  NAND2_X1 U3863 ( .A1(n3905), .A2(REG0_REG_30__SCAN_IN), .ZN(n3035) );
  OAI211_X1 U3864 ( .C1(n3908), .C2(n3037), .A(n3036), .B(n3035), .ZN(n3923)
         );
  XNOR2_X1 U3865 ( .A(n3038), .B(IR_REG_27__SCAN_IN), .ZN(n4501) );
  AND2_X1 U3866 ( .A1(n4501), .A2(B_REG_SCAN_IN), .ZN(n3039) );
  NOR2_X1 U3867 ( .A1(n4378), .A2(n3039), .ZN(n4138) );
  AOI21_X2 U3868 ( .B1(n3041), .B2(n4348), .A(n3040), .ZN(n4150) );
  NAND2_X1 U3869 ( .A1(n4174), .A2(n4374), .ZN(n3042) );
  OAI211_X1 U3870 ( .C1(n3912), .C2(n4323), .A(n4150), .B(n3042), .ZN(n3043)
         );
  INV_X1 U3871 ( .A(n3045), .ZN(n3059) );
  INV_X1 U3872 ( .A(n3912), .ZN(n4149) );
  INV_X1 U3873 ( .A(n3047), .ZN(n3048) );
  OAI21_X1 U3874 ( .B1(n3069), .B2(n4673), .A(n3048), .ZN(U3515) );
  XNOR2_X1 U3875 ( .A(n3049), .B(n3952), .ZN(n4158) );
  INV_X1 U3876 ( .A(n4667), .ZN(n4441) );
  INV_X1 U3877 ( .A(n3952), .ZN(n3050) );
  XNOR2_X1 U3878 ( .A(n3051), .B(n3050), .ZN(n3052) );
  NAND2_X1 U3879 ( .A1(n3052), .A2(n4348), .ZN(n4167) );
  INV_X1 U3880 ( .A(n4160), .ZN(n3053) );
  OAI22_X1 U3881 ( .A1(n3053), .A2(n4378), .B1(n4323), .B2(n4166), .ZN(n3054)
         );
  AOI21_X1 U3882 ( .B1(n4374), .B2(n4161), .A(n3054), .ZN(n3055) );
  OAI21_X1 U3883 ( .B1(n4158), .B2(n4441), .A(n3056), .ZN(n3062) );
  MUX2_X1 U3884 ( .A(REG1_REG_28__SCAN_IN), .B(n3062), .S(n4682), .Z(n3057) );
  INV_X1 U3885 ( .A(n3057), .ZN(n3061) );
  INV_X1 U3886 ( .A(n3058), .ZN(n3060) );
  OAI21_X1 U3887 ( .B1(n3060), .B2(n4166), .A(n3059), .ZN(n4159) );
  NAND2_X1 U3888 ( .A1(n3061), .A2(n2332), .ZN(U3546) );
  MUX2_X1 U3889 ( .A(REG0_REG_28__SCAN_IN), .B(n3062), .S(n4675), .Z(n3063) );
  INV_X1 U3890 ( .A(n3063), .ZN(n3064) );
  NAND2_X1 U3891 ( .A1(n3064), .A2(n2331), .ZN(U3514) );
  OR2_X1 U3892 ( .A1(n4682), .A2(n3065), .ZN(n3066) );
  OAI21_X1 U3893 ( .B1(n3069), .B2(n4680), .A(n3068), .ZN(U3547) );
  INV_X2 U3894 ( .A(n4975), .ZN(U4043) );
  INV_X1 U3895 ( .A(n3233), .ZN(n3145) );
  INV_X1 U3896 ( .A(DATAI_5_), .ZN(n3071) );
  MUX2_X1 U3897 ( .A(n3145), .B(n3071), .S(U3149), .Z(n3072) );
  INV_X1 U3898 ( .A(n3072), .ZN(U3347) );
  NAND2_X1 U3899 ( .A1(U3149), .A2(DATAI_25_), .ZN(n3073) );
  OAI21_X1 U3900 ( .B1(n3074), .B2(U3149), .A(n3073), .ZN(U3327) );
  INV_X1 U3901 ( .A(DATAI_26_), .ZN(n4903) );
  NAND2_X1 U3902 ( .A1(n3088), .A2(STATE_REG_SCAN_IN), .ZN(n3075) );
  OAI21_X1 U3903 ( .B1(STATE_REG_SCAN_IN), .B2(n4903), .A(n3075), .ZN(U3326)
         );
  INV_X1 U3904 ( .A(DATAI_27_), .ZN(n3077) );
  NAND2_X1 U3905 ( .A1(n4501), .A2(STATE_REG_SCAN_IN), .ZN(n3076) );
  OAI21_X1 U3906 ( .B1(STATE_REG_SCAN_IN), .B2(n3077), .A(n3076), .ZN(U3325)
         );
  INV_X1 U3907 ( .A(DATAI_20_), .ZN(n4901) );
  NAND2_X1 U3908 ( .A1(n3078), .A2(STATE_REG_SCAN_IN), .ZN(n3079) );
  OAI21_X1 U3909 ( .B1(STATE_REG_SCAN_IN), .B2(n4901), .A(n3079), .ZN(U3332)
         );
  INV_X1 U3910 ( .A(DATAI_22_), .ZN(n4689) );
  NAND2_X1 U3911 ( .A1(n4057), .A2(STATE_REG_SCAN_IN), .ZN(n3080) );
  OAI21_X1 U3912 ( .B1(STATE_REG_SCAN_IN), .B2(n4689), .A(n3080), .ZN(U3330)
         );
  INV_X1 U3913 ( .A(DATAI_29_), .ZN(n4686) );
  NAND2_X1 U3914 ( .A1(n3081), .A2(STATE_REG_SCAN_IN), .ZN(n3082) );
  OAI21_X1 U3915 ( .B1(STATE_REG_SCAN_IN), .B2(n4686), .A(n3082), .ZN(U3323)
         );
  INV_X1 U3916 ( .A(DATAI_30_), .ZN(n4684) );
  NAND2_X1 U3917 ( .A1(n3083), .A2(STATE_REG_SCAN_IN), .ZN(n3084) );
  OAI21_X1 U3918 ( .B1(STATE_REG_SCAN_IN), .B2(n4684), .A(n3084), .ZN(U3322)
         );
  INV_X1 U3919 ( .A(DATAI_24_), .ZN(n3085) );
  MUX2_X1 U3920 ( .A(n3085), .B(n2864), .S(STATE_REG_SCAN_IN), .Z(n3086) );
  INV_X1 U3921 ( .A(n3086), .ZN(U3328) );
  NOR3_X1 U3922 ( .A1(n3089), .A2(n3088), .A3(n4630), .ZN(n3090) );
  AOI21_X1 U3923 ( .B1(n4628), .B2(n3091), .A(n3090), .ZN(U3458) );
  INV_X1 U3924 ( .A(D_REG_1__SCAN_IN), .ZN(n4733) );
  INV_X1 U3925 ( .A(n3347), .ZN(n3093) );
  AOI22_X1 U3926 ( .A1(n4628), .A2(n4733), .B1(n3093), .B2(n3092), .ZN(U3459)
         );
  INV_X1 U3927 ( .A(n3095), .ZN(n3094) );
  NAND2_X1 U3928 ( .A1(n3094), .A2(STATE_REG_SCAN_IN), .ZN(n4059) );
  NAND2_X1 U3929 ( .A1(n3346), .A2(n4059), .ZN(n3113) );
  NAND2_X1 U3930 ( .A1(n3096), .A2(n3095), .ZN(n3097) );
  AND2_X1 U3931 ( .A1(n3097), .A2(n3909), .ZN(n3112) );
  INV_X1 U3932 ( .A(n3112), .ZN(n3098) );
  NOR2_X1 U3933 ( .A1(n4604), .A2(U4043), .ZN(U3148) );
  INV_X1 U3934 ( .A(DATAO_REG_11__SCAN_IN), .ZN(n4918) );
  NAND2_X1 U3935 ( .A1(n3620), .A2(U4043), .ZN(n3099) );
  OAI21_X1 U3936 ( .B1(U4043), .B2(n4918), .A(n3099), .ZN(U3561) );
  INV_X1 U3937 ( .A(DATAO_REG_0__SCAN_IN), .ZN(n4840) );
  NAND2_X1 U3938 ( .A1(n3462), .A2(U4043), .ZN(n3100) );
  OAI21_X1 U3939 ( .B1(U4043), .B2(n4840), .A(n3100), .ZN(U3550) );
  INV_X1 U3940 ( .A(DATAO_REG_12__SCAN_IN), .ZN(n4845) );
  NAND2_X1 U3941 ( .A1(n3513), .A2(U4043), .ZN(n3101) );
  OAI21_X1 U3942 ( .B1(U4043), .B2(n4845), .A(n3101), .ZN(U3562) );
  INV_X1 U3943 ( .A(DATAO_REG_16__SCAN_IN), .ZN(n4928) );
  NAND2_X1 U3944 ( .A1(n3738), .A2(U4043), .ZN(n3102) );
  OAI21_X1 U3945 ( .B1(U4043), .B2(n4928), .A(n3102), .ZN(U3566) );
  XNOR2_X1 U3946 ( .A(n3104), .B(n3103), .ZN(n3111) );
  INV_X1 U3947 ( .A(n3105), .ZN(n3108) );
  NAND3_X1 U3948 ( .A1(n3108), .A2(n3107), .A3(n3106), .ZN(n3151) );
  AOI22_X1 U3949 ( .A1(n3151), .A2(REG3_REG_1__SCAN_IN), .B1(n3799), .B2(n4068), .ZN(n3110) );
  AOI22_X1 U3950 ( .A1(n3798), .A2(n3462), .B1(n3461), .B2(n3880), .ZN(n3109)
         );
  OAI211_X1 U3951 ( .C1(n3111), .C2(n3869), .A(n3110), .B(n3109), .ZN(U3219)
         );
  INV_X1 U3952 ( .A(n4501), .ZN(n3197) );
  NOR2_X1 U3953 ( .A1(n3197), .A2(n3114), .ZN(n4055) );
  INV_X1 U3954 ( .A(REG2_REG_1__SCAN_IN), .ZN(n4075) );
  AND2_X1 U3955 ( .A1(IR_REG_0__SCAN_IN), .A2(REG2_REG_0__SCAN_IN), .ZN(n4078)
         );
  NAND2_X1 U3956 ( .A1(n3116), .A2(REG2_REG_1__SCAN_IN), .ZN(n3115) );
  OAI211_X1 U3957 ( .C1(n3116), .C2(REG2_REG_1__SCAN_IN), .A(n4078), .B(n3115), 
        .ZN(n4076) );
  INV_X1 U3958 ( .A(REG2_REG_3__SCAN_IN), .ZN(n3398) );
  XNOR2_X1 U3959 ( .A(n3139), .B(n3398), .ZN(n3122) );
  INV_X1 U3960 ( .A(REG1_REG_3__SCAN_IN), .ZN(n3120) );
  XNOR2_X1 U3961 ( .A(n3116), .B(REG1_REG_1__SCAN_IN), .ZN(n4071) );
  NOR3_X1 U3962 ( .A1(n4071), .A2(n2309), .A3(n4676), .ZN(n4070) );
  MUX2_X1 U3963 ( .A(n3117), .B(REG1_REG_2__SCAN_IN), .S(n4496), .Z(n3192) );
  INV_X1 U3964 ( .A(n4503), .ZN(n3118) );
  NOR2_X2 U3965 ( .A1(n3118), .A2(n4501), .ZN(n4606) );
  AOI211_X1 U3966 ( .C1(n3120), .C2(n3119), .A(n3134), .B(n4069), .ZN(n3121)
         );
  AOI21_X1 U3967 ( .B1(n4549), .B2(n3122), .A(n3121), .ZN(n3124) );
  AOI22_X1 U3968 ( .A1(n4604), .A2(ADDR_REG_3__SCAN_IN), .B1(
        REG3_REG_3__SCAN_IN), .B2(U3149), .ZN(n3123) );
  OAI211_X1 U3969 ( .C1(n2235), .C2(n4610), .A(n3124), .B(n3123), .ZN(U3243)
         );
  INV_X1 U3970 ( .A(n3126), .ZN(n3127) );
  AOI21_X1 U3971 ( .B1(n3125), .B2(n3128), .A(n3127), .ZN(n3131) );
  AOI22_X1 U3972 ( .A1(n3798), .A2(n2928), .B1(n3167), .B2(n3880), .ZN(n3130)
         );
  AOI22_X1 U3973 ( .A1(n3151), .A2(REG3_REG_2__SCAN_IN), .B1(n3799), .B2(n3383), .ZN(n3129) );
  OAI211_X1 U3974 ( .C1(n3131), .C2(n3869), .A(n3130), .B(n3129), .ZN(U3234)
         );
  INV_X1 U3975 ( .A(n3136), .ZN(n3137) );
  XNOR2_X1 U3976 ( .A(n3233), .B(REG1_REG_5__SCAN_IN), .ZN(n3138) );
  AOI211_X1 U3977 ( .C1(n2182), .C2(n3138), .A(n4069), .B(n3234), .ZN(n3148)
         );
  XNOR2_X1 U3978 ( .A(n3140), .B(n4494), .ZN(n3203) );
  INV_X1 U3979 ( .A(n3140), .ZN(n3141) );
  AOI22_X1 U3980 ( .A1(n3203), .A2(REG2_REG_4__SCAN_IN), .B1(n4494), .B2(n3141), .ZN(n3143) );
  INV_X1 U3981 ( .A(REG2_REG_5__SCAN_IN), .ZN(n4801) );
  MUX2_X1 U3982 ( .A(n4801), .B(REG2_REG_5__SCAN_IN), .S(n3233), .Z(n3142) );
  NOR2_X1 U3983 ( .A1(n3143), .A2(n3142), .ZN(n3230) );
  AOI211_X1 U3984 ( .C1(n3143), .C2(n3142), .A(n3230), .B(n4600), .ZN(n3147)
         );
  AND2_X1 U3985 ( .A1(U3149), .A2(REG3_REG_5__SCAN_IN), .ZN(n3225) );
  AOI21_X1 U3986 ( .B1(n4604), .B2(ADDR_REG_5__SCAN_IN), .A(n3225), .ZN(n3144)
         );
  OAI21_X1 U3987 ( .B1(n4610), .B2(n3145), .A(n3144), .ZN(n3146) );
  OR3_X1 U3988 ( .A1(n3148), .A2(n3147), .A3(n3146), .ZN(U3245) );
  XOR2_X1 U3989 ( .A(n3150), .B(n3149), .Z(n3201) );
  AOI22_X1 U3990 ( .A1(n3201), .A2(n3874), .B1(n3880), .B2(n2966), .ZN(n3153)
         );
  NAND2_X1 U3991 ( .A1(n3151), .A2(REG3_REG_0__SCAN_IN), .ZN(n3152) );
  OAI211_X1 U3992 ( .C1(n3876), .C2(n2926), .A(n3153), .B(n3152), .ZN(U3229)
         );
  INV_X1 U3993 ( .A(DATAO_REG_18__SCAN_IN), .ZN(n4920) );
  NAND2_X1 U3994 ( .A1(n4421), .A2(U4043), .ZN(n3154) );
  OAI21_X1 U3995 ( .B1(U4043), .B2(n4920), .A(n3154), .ZN(U3568) );
  INV_X1 U3996 ( .A(DATAO_REG_23__SCAN_IN), .ZN(n4854) );
  NAND2_X1 U3997 ( .A1(n4261), .A2(U4043), .ZN(n3155) );
  OAI21_X1 U3998 ( .B1(U4043), .B2(n4854), .A(n3155), .ZN(U3573) );
  INV_X1 U3999 ( .A(DATAO_REG_17__SCAN_IN), .ZN(n4852) );
  NAND2_X1 U4000 ( .A1(n4432), .A2(U4043), .ZN(n3156) );
  OAI21_X1 U4001 ( .B1(U4043), .B2(n4852), .A(n3156), .ZN(U3567) );
  INV_X1 U4002 ( .A(DATAO_REG_8__SCAN_IN), .ZN(n4842) );
  NAND2_X1 U4003 ( .A1(n3496), .A2(U4043), .ZN(n3157) );
  OAI21_X1 U4004 ( .B1(U4043), .B2(n4842), .A(n3157), .ZN(U3558) );
  INV_X1 U4005 ( .A(DATAO_REG_30__SCAN_IN), .ZN(n4922) );
  NAND2_X1 U4006 ( .A1(n3923), .A2(U4043), .ZN(n3158) );
  OAI21_X1 U4007 ( .B1(U4043), .B2(n4922), .A(n3158), .ZN(U3580) );
  INV_X1 U4008 ( .A(DATAO_REG_3__SCAN_IN), .ZN(n4843) );
  NAND2_X1 U4009 ( .A1(n3383), .A2(U4043), .ZN(n3159) );
  OAI21_X1 U4010 ( .B1(U4043), .B2(n4843), .A(n3159), .ZN(U3553) );
  INV_X1 U4011 ( .A(DATAO_REG_21__SCAN_IN), .ZN(n4856) );
  NAND2_X1 U4012 ( .A1(n3160), .A2(U4043), .ZN(n3161) );
  OAI21_X1 U4013 ( .B1(U4043), .B2(n4856), .A(n3161), .ZN(U3571) );
  INV_X1 U4014 ( .A(DATAO_REG_14__SCAN_IN), .ZN(n4844) );
  NAND2_X1 U4015 ( .A1(n3674), .A2(U4043), .ZN(n3162) );
  OAI21_X1 U4016 ( .B1(U4043), .B2(n4844), .A(n3162), .ZN(U3564) );
  INV_X1 U4017 ( .A(DATAO_REG_19__SCAN_IN), .ZN(n4850) );
  NAND2_X1 U4018 ( .A1(n4344), .A2(U4043), .ZN(n3163) );
  OAI21_X1 U4019 ( .B1(U4043), .B2(n4850), .A(n3163), .ZN(U3569) );
  INV_X1 U4020 ( .A(DATAO_REG_20__SCAN_IN), .ZN(n4857) );
  NAND2_X1 U4021 ( .A1(n4280), .A2(U4043), .ZN(n3165) );
  OAI21_X1 U4022 ( .B1(U4043), .B2(n4857), .A(n3165), .ZN(U3570) );
  INV_X1 U4023 ( .A(n3166), .ZN(n3257) );
  NAND2_X1 U4024 ( .A1(n3457), .A2(n3167), .ZN(n3168) );
  NAND2_X1 U4025 ( .A1(n3257), .A2(n3168), .ZN(n3273) );
  OAI21_X1 U4026 ( .B1(n3967), .B2(n3170), .A(n3169), .ZN(n3175) );
  NAND2_X1 U4027 ( .A1(n3383), .A2(n4431), .ZN(n3172) );
  NAND2_X1 U4028 ( .A1(n2928), .A2(n4374), .ZN(n3171) );
  OAI211_X1 U4029 ( .C1(n4323), .C2(n3173), .A(n3172), .B(n3171), .ZN(n3174)
         );
  AOI21_X1 U4030 ( .B1(n3175), .B2(n4348), .A(n3174), .ZN(n3181) );
  NAND2_X1 U4031 ( .A1(n3176), .A2(n3967), .ZN(n3177) );
  NAND2_X1 U4032 ( .A1(n3178), .A2(n3177), .ZN(n4623) );
  INV_X1 U4033 ( .A(n4304), .ZN(n3179) );
  NAND2_X1 U4034 ( .A1(n4623), .A2(n3179), .ZN(n3180) );
  AND2_X1 U4035 ( .A1(n3181), .A2(n3180), .ZN(n4626) );
  INV_X1 U4036 ( .A(n4655), .ZN(n4664) );
  NAND2_X1 U4037 ( .A1(n4623), .A2(n4664), .ZN(n3182) );
  NAND2_X1 U4038 ( .A1(n4626), .A2(n3182), .ZN(n3272) );
  MUX2_X1 U4039 ( .A(REG1_REG_2__SCAN_IN), .B(n3272), .S(n4682), .Z(n3183) );
  INV_X1 U4040 ( .A(n3183), .ZN(n3184) );
  OAI21_X1 U4041 ( .B1(n4428), .B2(n3273), .A(n3184), .ZN(U3520) );
  XOR2_X1 U4042 ( .A(n3186), .B(n3185), .Z(n3196) );
  INV_X1 U40430 ( .A(n4496), .ZN(n3190) );
  NOR2_X1 U4044 ( .A1(n3187), .A2(STATE_REG_SCAN_IN), .ZN(n3188) );
  AOI21_X1 U4045 ( .B1(n4604), .B2(ADDR_REG_2__SCAN_IN), .A(n3188), .ZN(n3189)
         );
  OAI21_X1 U4046 ( .B1(n4610), .B2(n3190), .A(n3189), .ZN(n3195) );
  AOI211_X1 U4047 ( .C1(n3193), .C2(n3192), .A(n3191), .B(n4069), .ZN(n3194)
         );
  AOI211_X1 U4048 ( .C1(n4549), .C2(n3196), .A(n3195), .B(n3194), .ZN(n3202)
         );
  NAND2_X1 U4049 ( .A1(n4488), .A2(n3197), .ZN(n3200) );
  INV_X1 U4050 ( .A(REG2_REG_0__SCAN_IN), .ZN(n3376) );
  NAND2_X1 U4051 ( .A1(n4501), .A2(n3376), .ZN(n3198) );
  NAND2_X1 U4052 ( .A1(n4488), .A2(n3198), .ZN(n4502) );
  AOI22_X1 U4053 ( .A1(n4055), .A2(n4078), .B1(n4502), .B2(n2309), .ZN(n3199)
         );
  OAI211_X1 U4054 ( .C1(n3201), .C2(n3200), .A(U4043), .B(n3199), .ZN(n3210)
         );
  NAND2_X1 U4055 ( .A1(n3202), .A2(n3210), .ZN(U3242) );
  XOR2_X1 U4056 ( .A(REG2_REG_4__SCAN_IN), .B(n3203), .Z(n3209) );
  AND2_X1 U4057 ( .A1(U3149), .A2(REG3_REG_4__SCAN_IN), .ZN(n3214) );
  AOI21_X1 U4058 ( .B1(n4604), .B2(ADDR_REG_4__SCAN_IN), .A(n3214), .ZN(n3204)
         );
  OAI21_X1 U4059 ( .B1(n4610), .B2(n3135), .A(n3204), .ZN(n3208) );
  AOI211_X1 U4060 ( .C1(n2447), .C2(n3206), .A(n4069), .B(n3205), .ZN(n3207)
         );
  AOI211_X1 U4061 ( .C1(n4549), .C2(n3209), .A(n3208), .B(n3207), .ZN(n3211)
         );
  NAND2_X1 U4062 ( .A1(n3211), .A2(n3210), .ZN(U3244) );
  INV_X1 U4063 ( .A(n3384), .ZN(n4981) );
  INV_X1 U4064 ( .A(n3383), .ZN(n3212) );
  OAI22_X1 U4065 ( .A1(n4981), .A2(n3876), .B1(n3877), .B2(n3212), .ZN(n3213)
         );
  AOI211_X1 U4066 ( .C1(n3382), .C2(n3880), .A(n3214), .B(n3213), .ZN(n3221)
         );
  AND2_X1 U4067 ( .A1(n3215), .A2(n3216), .ZN(n3219) );
  OAI211_X1 U4068 ( .C1(n3219), .C2(n3218), .A(n3874), .B(n3217), .ZN(n3220)
         );
  OAI211_X1 U4069 ( .C1(n3885), .C2(n3393), .A(n3221), .B(n3220), .ZN(U3227)
         );
  XNOR2_X1 U4070 ( .A(n3222), .B(n3223), .ZN(n3228) );
  INV_X1 U4071 ( .A(n4066), .ZN(n3306) );
  OAI22_X1 U4072 ( .A1(n3296), .A2(n3877), .B1(n3876), .B2(n3306), .ZN(n3224)
         );
  AOI211_X1 U4073 ( .C1(n3435), .C2(n3880), .A(n3225), .B(n3224), .ZN(n3227)
         );
  NAND2_X1 U4074 ( .A1(n3866), .A2(n3432), .ZN(n3226) );
  OAI211_X1 U4075 ( .C1(n3228), .C2(n3869), .A(n3227), .B(n3226), .ZN(U3224)
         );
  INV_X1 U4076 ( .A(DATAO_REG_28__SCAN_IN), .ZN(n4855) );
  NAND2_X1 U4077 ( .A1(n4174), .A2(U4043), .ZN(n3229) );
  OAI21_X1 U4078 ( .B1(U4043), .B2(n4855), .A(n3229), .ZN(U3578) );
  XNOR2_X1 U4079 ( .A(n3281), .B(n4493), .ZN(n3283) );
  XOR2_X1 U4080 ( .A(REG2_REG_6__SCAN_IN), .B(n3283), .Z(n3238) );
  INV_X1 U4081 ( .A(n4493), .ZN(n3232) );
  NAND2_X1 U4082 ( .A1(U3149), .A2(REG3_REG_6__SCAN_IN), .ZN(n3265) );
  NAND2_X1 U4083 ( .A1(n4604), .A2(ADDR_REG_6__SCAN_IN), .ZN(n3231) );
  OAI211_X1 U4084 ( .C1(n4610), .C2(n3232), .A(n3265), .B(n3231), .ZN(n3237)
         );
  INV_X1 U4085 ( .A(REG1_REG_6__SCAN_IN), .ZN(n3321) );
  AOI211_X1 U4086 ( .C1(n3235), .C2(n3321), .A(n4069), .B(n3277), .ZN(n3236)
         );
  AOI211_X1 U4087 ( .C1(n4549), .C2(n3238), .A(n3237), .B(n3236), .ZN(n3239)
         );
  INV_X1 U4088 ( .A(n3239), .ZN(U3246) );
  OAI21_X1 U4089 ( .B1(n3241), .B2(n3240), .A(n3215), .ZN(n3246) );
  MUX2_X1 U4090 ( .A(STATE_REG_SCAN_IN), .B(n3885), .S(n3242), .Z(n3244) );
  AOI22_X1 U4091 ( .A1(n3798), .A2(n4068), .B1(n3258), .B2(n3880), .ZN(n3243)
         );
  OAI211_X1 U4092 ( .C1(n3296), .C2(n3876), .A(n3244), .B(n3243), .ZN(n3245)
         );
  AOI21_X1 U4093 ( .B1(n3246), .B2(n3874), .A(n3245), .ZN(n3247) );
  INV_X1 U4094 ( .A(n3247), .ZN(U3215) );
  XNOR2_X1 U4095 ( .A(n3248), .B(n3249), .ZN(n3403) );
  INV_X1 U4096 ( .A(n3403), .ZN(n3255) );
  XNOR2_X1 U4097 ( .A(n3250), .B(n3249), .ZN(n3253) );
  AOI22_X1 U4098 ( .A1(n4068), .A2(n4374), .B1(n4429), .B2(n3258), .ZN(n3251)
         );
  OAI21_X1 U4099 ( .B1(n3296), .B2(n4378), .A(n3251), .ZN(n3252) );
  AOI21_X1 U4100 ( .B1(n3253), .B2(n4348), .A(n3252), .ZN(n3254) );
  OAI21_X1 U4101 ( .B1(n3403), .B2(n4304), .A(n3254), .ZN(n3397) );
  AOI21_X1 U4102 ( .B1(n4664), .B2(n3255), .A(n3397), .ZN(n3271) );
  INV_X1 U4103 ( .A(n4428), .ZN(n3502) );
  INV_X1 U4104 ( .A(n3256), .ZN(n3392) );
  AOI21_X1 U4105 ( .B1(n3258), .B2(n3257), .A(n3392), .ZN(n3400) );
  AOI22_X1 U4106 ( .A1(n3502), .A2(n3400), .B1(REG1_REG_3__SCAN_IN), .B2(n4680), .ZN(n3259) );
  OAI21_X1 U4107 ( .B1(n3271), .B2(n4680), .A(n3259), .ZN(U3521) );
  INV_X1 U4108 ( .A(n3261), .ZN(n3263) );
  NOR2_X1 U4109 ( .A1(n3263), .A2(n3262), .ZN(n3264) );
  XNOR2_X1 U4110 ( .A(n3260), .B(n3264), .ZN(n3269) );
  AOI22_X1 U4111 ( .A1(n3798), .A2(n3384), .B1(n3799), .B2(n4065), .ZN(n3266)
         );
  OAI211_X1 U4112 ( .C1(n3862), .C2(n3318), .A(n3266), .B(n3265), .ZN(n3267)
         );
  AOI21_X1 U4113 ( .B1(n3357), .B2(n3866), .A(n3267), .ZN(n3268) );
  OAI21_X1 U4114 ( .B1(n3269), .B2(n3869), .A(n3268), .ZN(U3236) );
  INV_X1 U4115 ( .A(n4485), .ZN(n3506) );
  AOI22_X1 U4116 ( .A1(n3506), .A2(n3400), .B1(REG0_REG_3__SCAN_IN), .B2(n4673), .ZN(n3270) );
  OAI21_X1 U4117 ( .B1(n3271), .B2(n4673), .A(n3270), .ZN(U3473) );
  INV_X1 U4118 ( .A(n3272), .ZN(n3275) );
  INV_X1 U4119 ( .A(n3273), .ZN(n4620) );
  AOI22_X1 U4120 ( .A1(n3506), .A2(n4620), .B1(REG0_REG_2__SCAN_IN), .B2(n4673), .ZN(n3274) );
  OAI21_X1 U4121 ( .B1(n3275), .B2(n4673), .A(n3274), .ZN(U3471) );
  INV_X1 U4122 ( .A(n3276), .ZN(n3278) );
  MUX2_X1 U4123 ( .A(n2508), .B(REG1_REG_7__SCAN_IN), .S(n4492), .Z(n3280) );
  OAI21_X1 U4124 ( .B1(n3337), .B2(n3280), .A(n4606), .ZN(n3279) );
  AOI21_X1 U4125 ( .B1(n3337), .B2(n3280), .A(n3279), .ZN(n3290) );
  INV_X1 U4126 ( .A(n3281), .ZN(n3282) );
  INV_X1 U4127 ( .A(REG2_REG_7__SCAN_IN), .ZN(n3425) );
  MUX2_X1 U4128 ( .A(n3425), .B(REG2_REG_7__SCAN_IN), .S(n4492), .Z(n3284) );
  AOI211_X1 U4129 ( .C1(n3285), .C2(n3284), .A(n4600), .B(n3338), .ZN(n3289)
         );
  INV_X1 U4130 ( .A(n4492), .ZN(n3287) );
  AND2_X1 U4131 ( .A1(U3149), .A2(REG3_REG_7__SCAN_IN), .ZN(n3308) );
  AOI21_X1 U4132 ( .B1(n4604), .B2(ADDR_REG_7__SCAN_IN), .A(n3308), .ZN(n3286)
         );
  OAI21_X1 U4133 ( .B1(n4610), .B2(n3287), .A(n3286), .ZN(n3288) );
  OR3_X1 U4134 ( .A1(n3290), .A2(n3289), .A3(n3288), .ZN(U3247) );
  INV_X1 U4135 ( .A(n3292), .ZN(n3989) );
  NAND2_X1 U4136 ( .A1(n3989), .A2(n4005), .ZN(n3964) );
  XOR2_X1 U4137 ( .A(n3291), .B(n3964), .Z(n3442) );
  XNOR2_X1 U4138 ( .A(n3293), .B(n3964), .ZN(n3294) );
  NAND2_X1 U4139 ( .A1(n3294), .A2(n4348), .ZN(n3439) );
  AOI22_X1 U4140 ( .A1(n4066), .A2(n4431), .B1(n4429), .B2(n3435), .ZN(n3295)
         );
  OAI211_X1 U4141 ( .C1(n3296), .C2(n4434), .A(n3439), .B(n3295), .ZN(n3297)
         );
  AOI21_X1 U4142 ( .B1(n3442), .B2(n4667), .A(n3297), .ZN(n3301) );
  AND2_X1 U4143 ( .A1(n3390), .A2(n3435), .ZN(n3298) );
  NOR2_X1 U4144 ( .A1(n3319), .A2(n3298), .ZN(n3431) );
  AOI22_X1 U4145 ( .A1(n3431), .A2(n3502), .B1(REG1_REG_5__SCAN_IN), .B2(n4680), .ZN(n3299) );
  OAI21_X1 U4146 ( .B1(n3301), .B2(n4680), .A(n3299), .ZN(U3523) );
  AOI22_X1 U4147 ( .A1(n3431), .A2(n3506), .B1(REG0_REG_5__SCAN_IN), .B2(n4673), .ZN(n3300) );
  OAI21_X1 U4148 ( .B1(n3301), .B2(n4673), .A(n3300), .ZN(U3477) );
  AOI21_X1 U4149 ( .B1(n3302), .B2(n3303), .A(n3869), .ZN(n3305) );
  NAND2_X1 U4150 ( .A1(n3305), .A2(n3304), .ZN(n3311) );
  INV_X1 U4151 ( .A(n3496), .ZN(n3476) );
  OAI22_X1 U4152 ( .A1(n3476), .A2(n3876), .B1(n3877), .B2(n3306), .ZN(n3307)
         );
  AOI211_X1 U4153 ( .C1(n3309), .C2(n3880), .A(n3308), .B(n3307), .ZN(n3310)
         );
  OAI211_X1 U4154 ( .C1(n3885), .C2(n3424), .A(n3311), .B(n3310), .ZN(U3210)
         );
  NAND2_X1 U4155 ( .A1(n3992), .A2(n4004), .ZN(n3954) );
  XNOR2_X1 U4156 ( .A(n3312), .B(n3954), .ZN(n3367) );
  OAI22_X1 U4157 ( .A1(n3313), .A2(n4378), .B1(n4323), .B2(n3318), .ZN(n3316)
         );
  XNOR2_X1 U4158 ( .A(n3314), .B(n3954), .ZN(n3356) );
  INV_X1 U4159 ( .A(n4348), .ZN(n4326) );
  NOR2_X1 U4160 ( .A1(n3356), .A2(n4326), .ZN(n3315) );
  AOI211_X1 U4161 ( .C1(n4374), .C2(n3384), .A(n3316), .B(n3315), .ZN(n3317)
         );
  OAI21_X1 U4162 ( .B1(n4441), .B2(n3367), .A(n3317), .ZN(n3326) );
  NOR2_X1 U4163 ( .A1(n3319), .A2(n3318), .ZN(n3320) );
  OR2_X1 U4164 ( .A1(n3423), .A2(n3320), .ZN(n3363) );
  OAI22_X1 U4165 ( .A1(n3363), .A2(n4428), .B1(n4682), .B2(n3321), .ZN(n3322)
         );
  AOI21_X1 U4166 ( .B1(n3326), .B2(n4682), .A(n3322), .ZN(n3323) );
  INV_X1 U4167 ( .A(n3323), .ZN(U3524) );
  INV_X1 U4168 ( .A(REG0_REG_6__SCAN_IN), .ZN(n3324) );
  OAI22_X1 U4169 ( .A1(n3363), .A2(n4485), .B1(n4675), .B2(n3324), .ZN(n3325)
         );
  AOI21_X1 U4170 ( .B1(n3326), .B2(n4675), .A(n3325), .ZN(n3327) );
  INV_X1 U4171 ( .A(n3327), .ZN(U3479) );
  XOR2_X1 U4172 ( .A(n3330), .B(n3329), .Z(n3331) );
  XNOR2_X1 U4173 ( .A(n3328), .B(n3331), .ZN(n3335) );
  AOI22_X1 U4174 ( .A1(n3798), .A2(n4065), .B1(n3799), .B2(n4064), .ZN(n3332)
         );
  NAND2_X1 U4175 ( .A1(REG3_REG_8__SCAN_IN), .A2(U3149), .ZN(n3341) );
  OAI211_X1 U4176 ( .C1(n3862), .C2(n3553), .A(n3332), .B(n3341), .ZN(n3333)
         );
  AOI21_X1 U4177 ( .B1(n4611), .B2(n3866), .A(n3333), .ZN(n3334) );
  OAI21_X1 U4178 ( .B1(n3335), .B2(n3869), .A(n3334), .ZN(U3218) );
  OAI21_X1 U4179 ( .B1(n3337), .B2(n2508), .A(n3336), .ZN(n4105) );
  XNOR2_X1 U4180 ( .A(n4105), .B(n4491), .ZN(n4108) );
  XOR2_X1 U4181 ( .A(REG1_REG_8__SCAN_IN), .B(n4108), .Z(n3345) );
  INV_X1 U4182 ( .A(n4491), .ZN(n4106) );
  XNOR2_X1 U4183 ( .A(REG2_REG_8__SCAN_IN), .B(n4088), .ZN(n3339) );
  NAND2_X1 U4184 ( .A1(n4549), .A2(n3339), .ZN(n3340) );
  NAND2_X1 U4185 ( .A1(n3341), .A2(n3340), .ZN(n3342) );
  AOI21_X1 U4186 ( .B1(n4604), .B2(ADDR_REG_8__SCAN_IN), .A(n3342), .ZN(n3344)
         );
  INV_X1 U4187 ( .A(n4610), .ZN(n4074) );
  NAND2_X1 U4188 ( .A1(n4074), .A2(n4491), .ZN(n3343) );
  OAI211_X1 U4189 ( .C1(n3345), .C2(n4069), .A(n3344), .B(n3343), .ZN(U3248)
         );
  OAI21_X1 U4190 ( .B1(n3346), .B2(n4733), .A(n4628), .ZN(n3351) );
  AND2_X1 U4191 ( .A1(n3348), .A2(n3347), .ZN(n3350) );
  NAND4_X1 U4192 ( .A1(n3352), .A2(n3351), .A3(n3350), .A4(n3349), .ZN(n3353)
         );
  NAND2_X1 U4193 ( .A1(n3354), .A2(n4490), .ZN(n3373) );
  NAND2_X1 U4194 ( .A1(n4304), .A2(n3373), .ZN(n3355) );
  INV_X1 U4195 ( .A(n3356), .ZN(n3365) );
  NAND2_X1 U4196 ( .A1(n4357), .A2(n4348), .ZN(n3591) );
  INV_X1 U4197 ( .A(n3591), .ZN(n3453) );
  NAND2_X1 U4198 ( .A1(n4357), .A2(n4133), .ZN(n4355) );
  INV_X1 U4199 ( .A(n3357), .ZN(n3358) );
  OAI22_X1 U4200 ( .A1(n4357), .A2(n2242), .B1(n3358), .B2(n4332), .ZN(n3359)
         );
  AOI21_X1 U4201 ( .B1(n3360), .B2(n4148), .A(n3359), .ZN(n3362) );
  NAND2_X1 U4202 ( .A1(n4357), .A2(n4374), .ZN(n4145) );
  AND2_X1 U4203 ( .A1(n4357), .A2(n4431), .ZN(n4279) );
  AOI22_X1 U4204 ( .A1(n4281), .A2(n3384), .B1(n4279), .B2(n4065), .ZN(n3361)
         );
  OAI211_X1 U4205 ( .C1(n3363), .C2(n4331), .A(n3362), .B(n3361), .ZN(n3364)
         );
  AOI21_X1 U4206 ( .B1(n3365), .B2(n3453), .A(n3364), .ZN(n3366) );
  OAI21_X1 U4207 ( .B1(n4360), .B2(n3367), .A(n3366), .ZN(U3284) );
  NAND2_X1 U4208 ( .A1(n2966), .A2(n3368), .ZN(n4647) );
  NAND2_X1 U4209 ( .A1(n3462), .A2(n3369), .ZN(n3978) );
  NAND2_X1 U4210 ( .A1(n3976), .A2(n3978), .ZN(n4651) );
  NAND2_X1 U4211 ( .A1(n4304), .A2(n4326), .ZN(n3370) );
  AOI22_X1 U4212 ( .A1(n4651), .A2(n3370), .B1(n4431), .B2(n2928), .ZN(n4648)
         );
  OAI21_X1 U4213 ( .B1(n3371), .B2(n4647), .A(n4648), .ZN(n3372) );
  AOI22_X1 U4214 ( .A1(n3372), .A2(n4357), .B1(REG3_REG_0__SCAN_IN), .B2(n4619), .ZN(n3375) );
  NOR2_X1 U4215 ( .A1(n4612), .A2(n3373), .ZN(n4622) );
  NAND2_X1 U4216 ( .A1(n4622), .A2(n4651), .ZN(n3374) );
  OAI211_X1 U4217 ( .C1(n4357), .C2(n3376), .A(n3375), .B(n3374), .ZN(U3290)
         );
  NAND2_X1 U4218 ( .A1(n3378), .A2(n2934), .ZN(n3380) );
  NAND2_X1 U4219 ( .A1(n3377), .A2(n3380), .ZN(n4660) );
  INV_X1 U4220 ( .A(n4622), .ZN(n3468) );
  XNOR2_X1 U4221 ( .A(n3381), .B(n2934), .ZN(n3388) );
  AOI22_X1 U4222 ( .A1(n3383), .A2(n4374), .B1(n3382), .B2(n4429), .ZN(n3386)
         );
  NAND2_X1 U4223 ( .A1(n3384), .A2(n4431), .ZN(n3385) );
  OAI211_X1 U4224 ( .C1(n4660), .C2(n4304), .A(n3386), .B(n3385), .ZN(n3387)
         );
  AOI21_X1 U4225 ( .B1(n3388), .B2(n4348), .A(n3387), .ZN(n3389) );
  INV_X1 U4226 ( .A(n3389), .ZN(n4662) );
  OAI211_X1 U4227 ( .C1(n3392), .C2(n3391), .A(n4437), .B(n3390), .ZN(n4661)
         );
  OAI22_X1 U4228 ( .A1(n4661), .A2(n4490), .B1(n4332), .B2(n3393), .ZN(n3394)
         );
  OAI21_X1 U4229 ( .B1(n4662), .B2(n3394), .A(n4357), .ZN(n3396) );
  NAND2_X1 U4230 ( .A1(n4612), .A2(REG2_REG_4__SCAN_IN), .ZN(n3395) );
  OAI211_X1 U4231 ( .C1(n4660), .C2(n3468), .A(n3396), .B(n3395), .ZN(U3286)
         );
  NAND2_X1 U4232 ( .A1(n3397), .A2(n4357), .ZN(n3402) );
  OAI22_X1 U4233 ( .A1(n4357), .A2(n3398), .B1(REG3_REG_3__SCAN_IN), .B2(n4332), .ZN(n3399) );
  AOI21_X1 U4234 ( .B1(n4621), .B2(n3400), .A(n3399), .ZN(n3401) );
  OAI211_X1 U4235 ( .C1(n3403), .C2(n3468), .A(n3402), .B(n3401), .ZN(U3287)
         );
  INV_X1 U4236 ( .A(n4006), .ZN(n4001) );
  NAND2_X1 U4237 ( .A1(n4001), .A2(n3998), .ZN(n3955) );
  XNOR2_X1 U4238 ( .A(n3404), .B(n3955), .ZN(n3405) );
  NAND2_X1 U4239 ( .A1(n3405), .A2(n4348), .ZN(n3498) );
  OR2_X1 U4240 ( .A1(n3406), .A2(n3407), .ZN(n3409) );
  NAND2_X1 U4241 ( .A1(n3409), .A2(n3408), .ZN(n3411) );
  INV_X1 U4242 ( .A(n3955), .ZN(n3410) );
  XNOR2_X1 U4243 ( .A(n3411), .B(n3410), .ZN(n3494) );
  NAND2_X1 U4244 ( .A1(n3494), .A2(n4277), .ZN(n3417) );
  AOI21_X1 U4245 ( .B1(n3495), .B2(n3552), .A(n3448), .ZN(n3507) );
  AOI22_X1 U4246 ( .A1(n4148), .A2(n3495), .B1(n4279), .B2(n4063), .ZN(n3412)
         );
  OAI21_X1 U4247 ( .B1(n3476), .B2(n4145), .A(n3412), .ZN(n3415) );
  INV_X1 U4248 ( .A(REG2_REG_9__SCAN_IN), .ZN(n4950) );
  OAI22_X1 U4249 ( .A1(n3413), .A2(n4332), .B1(n4950), .B2(n4357), .ZN(n3414)
         );
  AOI211_X1 U4250 ( .C1(n3507), .C2(n4621), .A(n3415), .B(n3414), .ZN(n3416)
         );
  OAI211_X1 U4251 ( .C1(n4627), .C2(n3498), .A(n3417), .B(n3416), .ZN(U3281)
         );
  OAI22_X1 U4252 ( .A1(n3476), .A2(n4378), .B1(n3422), .B2(n4323), .ZN(n3421)
         );
  XOR2_X1 U4253 ( .A(n3418), .B(n3968), .Z(n3419) );
  NOR2_X1 U4254 ( .A1(n3419), .A2(n4326), .ZN(n3420) );
  AOI211_X1 U4255 ( .C1(n4374), .C2(n4066), .A(n3421), .B(n3420), .ZN(n4672)
         );
  OAI211_X1 U4256 ( .C1(n3423), .C2(n3422), .A(n4437), .B(n3551), .ZN(n4671)
         );
  INV_X1 U4257 ( .A(n4671), .ZN(n3428) );
  INV_X1 U4258 ( .A(n4355), .ZN(n3427) );
  OAI22_X1 U4259 ( .A1(n4357), .A2(n3425), .B1(n3424), .B2(n4332), .ZN(n3426)
         );
  AOI21_X1 U4260 ( .B1(n3428), .B2(n3427), .A(n3426), .ZN(n3430) );
  OR2_X1 U4261 ( .A1(n3406), .A2(n3968), .ZN(n4669) );
  NAND2_X1 U4262 ( .A1(n3406), .A2(n3968), .ZN(n4668) );
  NAND3_X1 U4263 ( .A1(n4669), .A2(n4668), .A3(n4277), .ZN(n3429) );
  OAI211_X1 U4264 ( .C1(n4672), .C2(n4612), .A(n3430), .B(n3429), .ZN(U3283)
         );
  NAND2_X1 U4265 ( .A1(n3431), .A2(n4621), .ZN(n3438) );
  INV_X1 U4266 ( .A(n3432), .ZN(n3433) );
  OAI22_X1 U4267 ( .A1(n4357), .A2(n4801), .B1(n3433), .B2(n4332), .ZN(n3434)
         );
  AOI21_X1 U4268 ( .B1(n3435), .B2(n4148), .A(n3434), .ZN(n3437) );
  AOI22_X1 U4269 ( .A1(n4281), .A2(n4067), .B1(n4279), .B2(n4066), .ZN(n3436)
         );
  NAND3_X1 U4270 ( .A1(n3438), .A2(n3437), .A3(n3436), .ZN(n3441) );
  NOR2_X1 U4271 ( .A1(n3439), .A2(n4627), .ZN(n3440) );
  AOI211_X1 U4272 ( .C1(n3442), .C2(n4277), .A(n3441), .B(n3440), .ZN(n3443)
         );
  INV_X1 U4273 ( .A(n3443), .ZN(U3285) );
  NAND2_X1 U4274 ( .A1(n4009), .A2(n4012), .ZN(n3958) );
  XNOR2_X1 U4275 ( .A(n3444), .B(n3958), .ZN(n3531) );
  INV_X1 U4276 ( .A(n3531), .ZN(n3455) );
  INV_X1 U4277 ( .A(n3958), .ZN(n3445) );
  XNOR2_X1 U4278 ( .A(n3446), .B(n3445), .ZN(n3530) );
  INV_X1 U4279 ( .A(n3520), .ZN(n3447) );
  OAI21_X1 U4280 ( .B1(n3448), .B2(n3528), .A(n3447), .ZN(n3539) );
  NOR2_X1 U4281 ( .A1(n3539), .A2(n4331), .ZN(n3452) );
  AOI22_X1 U4282 ( .A1(n4281), .A2(n4064), .B1(n4279), .B2(n3620), .ZN(n3450)
         );
  AOI22_X1 U4283 ( .A1(n4612), .A2(REG2_REG_10__SCAN_IN), .B1(n3482), .B2(
        n4619), .ZN(n3449) );
  OAI211_X1 U4284 ( .C1(n3528), .C2(n4285), .A(n3450), .B(n3449), .ZN(n3451)
         );
  AOI211_X1 U4285 ( .C1(n3530), .C2(n3453), .A(n3452), .B(n3451), .ZN(n3454)
         );
  OAI21_X1 U4286 ( .B1(n3455), .B2(n4360), .A(n3454), .ZN(U3280) );
  NAND2_X1 U4287 ( .A1(n3461), .A2(n2966), .ZN(n3456) );
  NAND2_X1 U4288 ( .A1(n3457), .A2(n3456), .ZN(n4653) );
  XNOR2_X1 U4289 ( .A(n2965), .B(n3976), .ZN(n3466) );
  OR2_X1 U4290 ( .A1(n2965), .A2(n3458), .ZN(n3459) );
  NAND2_X1 U4291 ( .A1(n3460), .A2(n3459), .ZN(n4656) );
  AOI22_X1 U4292 ( .A1(n4068), .A2(n4431), .B1(n4429), .B2(n3461), .ZN(n3464)
         );
  NAND2_X1 U4293 ( .A1(n3462), .A2(n4374), .ZN(n3463) );
  OAI211_X1 U4294 ( .C1(n4656), .C2(n4304), .A(n3464), .B(n3463), .ZN(n3465)
         );
  AOI21_X1 U4295 ( .B1(n4348), .B2(n3466), .A(n3465), .ZN(n3467) );
  INV_X1 U4296 ( .A(n3467), .ZN(n4658) );
  OAI22_X1 U4297 ( .A1(n4357), .A2(n4075), .B1(n2352), .B2(n4332), .ZN(n3470)
         );
  NOR2_X1 U4298 ( .A1(n3468), .A2(n4656), .ZN(n3469) );
  AOI211_X1 U4299 ( .C1(n4658), .C2(n4357), .A(n3470), .B(n3469), .ZN(n3471)
         );
  OAI21_X1 U4300 ( .B1(n4331), .B2(n4653), .A(n3471), .ZN(U3289) );
  INV_X1 U4301 ( .A(n3473), .ZN(n3474) );
  AOI21_X1 U4302 ( .B1(n3475), .B2(n3472), .A(n3474), .ZN(n3481) );
  INV_X1 U4303 ( .A(REG3_REG_9__SCAN_IN), .ZN(n4911) );
  NOR2_X1 U4304 ( .A1(STATE_REG_SCAN_IN), .A2(n4911), .ZN(n4516) );
  OAI22_X1 U4305 ( .A1(n3476), .A2(n3877), .B1(n3876), .B2(n3545), .ZN(n3477)
         );
  AOI211_X1 U4306 ( .C1(n3495), .C2(n3880), .A(n4516), .B(n3477), .ZN(n3480)
         );
  NAND2_X1 U4307 ( .A1(n3866), .A2(n3478), .ZN(n3479) );
  OAI211_X1 U4308 ( .C1(n3481), .C2(n3869), .A(n3480), .B(n3479), .ZN(U3228)
         );
  INV_X1 U4309 ( .A(n3482), .ZN(n3493) );
  AND2_X1 U4310 ( .A1(n3473), .A2(n3483), .ZN(n3486) );
  OAI211_X1 U4311 ( .C1(n3486), .C2(n3485), .A(n3874), .B(n3484), .ZN(n3492)
         );
  INV_X1 U4312 ( .A(REG3_REG_10__SCAN_IN), .ZN(n3487) );
  NOR2_X1 U4313 ( .A1(STATE_REG_SCAN_IN), .A2(n3487), .ZN(n4525) );
  INV_X1 U4314 ( .A(n4064), .ZN(n3560) );
  INV_X1 U4315 ( .A(n3620), .ZN(n3488) );
  OAI22_X1 U4316 ( .A1(n3560), .A2(n3877), .B1(n3876), .B2(n3488), .ZN(n3489)
         );
  AOI211_X1 U4317 ( .C1(n3490), .C2(n3880), .A(n4525), .B(n3489), .ZN(n3491)
         );
  OAI211_X1 U4318 ( .C1(n3885), .C2(n3493), .A(n3492), .B(n3491), .ZN(U3214)
         );
  NAND2_X1 U4319 ( .A1(n3494), .A2(n4667), .ZN(n3500) );
  AOI22_X1 U4320 ( .A1(n4063), .A2(n4431), .B1(n4429), .B2(n3495), .ZN(n3499)
         );
  NAND2_X1 U4321 ( .A1(n3496), .A2(n4374), .ZN(n3497) );
  NAND4_X1 U4322 ( .A1(n3500), .A2(n3499), .A3(n3498), .A4(n3497), .ZN(n3504)
         );
  MUX2_X1 U4323 ( .A(REG1_REG_9__SCAN_IN), .B(n3504), .S(n4682), .Z(n3501) );
  AOI21_X1 U4324 ( .B1(n3502), .B2(n3507), .A(n3501), .ZN(n3503) );
  INV_X1 U4325 ( .A(n3503), .ZN(U3527) );
  MUX2_X1 U4326 ( .A(REG0_REG_9__SCAN_IN), .B(n3504), .S(n4675), .Z(n3505) );
  AOI21_X1 U4327 ( .B1(n3507), .B2(n3506), .A(n3505), .ZN(n3508) );
  INV_X1 U4328 ( .A(n3508), .ZN(U3485) );
  XNOR2_X1 U4329 ( .A(n3600), .B(n3962), .ZN(n3517) );
  INV_X1 U4330 ( .A(n3510), .ZN(n3511) );
  AOI21_X1 U4331 ( .B1(n3962), .B2(n3512), .A(n3511), .ZN(n3518) );
  AOI22_X1 U4332 ( .A1(n4063), .A2(n4374), .B1(n3547), .B2(n4429), .ZN(n3515)
         );
  NAND2_X1 U4333 ( .A1(n3513), .A2(n4431), .ZN(n3514) );
  OAI211_X1 U4334 ( .C1(n3518), .C2(n4304), .A(n3515), .B(n3514), .ZN(n3516)
         );
  AOI21_X1 U4335 ( .B1(n3517), .B2(n4348), .A(n3516), .ZN(n3609) );
  INV_X1 U4336 ( .A(n3518), .ZN(n3611) );
  OAI21_X1 U4337 ( .B1(n3520), .B2(n3519), .A(n3593), .ZN(n3617) );
  NOR2_X1 U4338 ( .A1(n3617), .A2(n4331), .ZN(n3524) );
  INV_X1 U4339 ( .A(REG2_REG_11__SCAN_IN), .ZN(n3522) );
  INV_X1 U4340 ( .A(n3521), .ZN(n3550) );
  OAI22_X1 U4341 ( .A1(n4357), .A2(n3522), .B1(n3550), .B2(n4332), .ZN(n3523)
         );
  AOI211_X1 U4342 ( .C1(n3611), .C2(n4622), .A(n3524), .B(n3523), .ZN(n3525)
         );
  OAI21_X1 U4343 ( .B1(n3609), .B2(n4627), .A(n3525), .ZN(U3279) );
  NAND2_X1 U4344 ( .A1(n4064), .A2(n4374), .ZN(n3527) );
  NAND2_X1 U4345 ( .A1(n3620), .A2(n4431), .ZN(n3526) );
  OAI211_X1 U4346 ( .C1(n4323), .C2(n3528), .A(n3527), .B(n3526), .ZN(n3529)
         );
  AOI21_X1 U4347 ( .B1(n3530), .B2(n4348), .A(n3529), .ZN(n3533) );
  NAND2_X1 U4348 ( .A1(n3531), .A2(n4667), .ZN(n3532) );
  NAND2_X1 U4349 ( .A1(n3533), .A2(n3532), .ZN(n3536) );
  MUX2_X1 U4350 ( .A(REG0_REG_10__SCAN_IN), .B(n3536), .S(n4675), .Z(n3534) );
  INV_X1 U4351 ( .A(n3534), .ZN(n3535) );
  OAI21_X1 U4352 ( .B1(n3539), .B2(n4485), .A(n3535), .ZN(U3487) );
  MUX2_X1 U4353 ( .A(REG1_REG_10__SCAN_IN), .B(n3536), .S(n4682), .Z(n3537) );
  INV_X1 U4354 ( .A(n3537), .ZN(n3538) );
  OAI21_X1 U4355 ( .B1(n4428), .B2(n3539), .A(n3538), .ZN(U3528) );
  NAND2_X1 U4356 ( .A1(n3542), .A2(n3541), .ZN(n3543) );
  XNOR2_X1 U4357 ( .A(n3540), .B(n3543), .ZN(n3544) );
  NAND2_X1 U4358 ( .A1(n3544), .A2(n3874), .ZN(n3549) );
  NOR2_X1 U4359 ( .A1(STATE_REG_SCAN_IN), .A2(n4923), .ZN(n4536) );
  OAI22_X1 U4360 ( .A1(n3675), .A2(n3876), .B1(n3877), .B2(n3545), .ZN(n3546)
         );
  AOI211_X1 U4361 ( .C1(n3547), .C2(n3880), .A(n4536), .B(n3546), .ZN(n3548)
         );
  OAI211_X1 U4362 ( .C1(n3885), .C2(n3550), .A(n3549), .B(n3548), .ZN(U3233)
         );
  INV_X1 U4363 ( .A(n3551), .ZN(n3554) );
  OAI21_X1 U4364 ( .B1(n3554), .B2(n3553), .A(n3552), .ZN(n4613) );
  INV_X1 U4365 ( .A(REG0_REG_8__SCAN_IN), .ZN(n3566) );
  NAND2_X1 U4366 ( .A1(n4669), .A2(n3555), .ZN(n3556) );
  NAND2_X1 U4367 ( .A1(n3997), .A2(n3996), .ZN(n3963) );
  XNOR2_X1 U4368 ( .A(n3556), .B(n3963), .ZN(n3561) );
  INV_X1 U4369 ( .A(n3561), .ZN(n4615) );
  XNOR2_X1 U4370 ( .A(n3557), .B(n3963), .ZN(n3564) );
  AOI22_X1 U4371 ( .A1(n4065), .A2(n4374), .B1(n4429), .B2(n3558), .ZN(n3559)
         );
  OAI21_X1 U4372 ( .B1(n3560), .B2(n4378), .A(n3559), .ZN(n3563) );
  NOR2_X1 U4373 ( .A1(n3561), .A2(n4304), .ZN(n3562) );
  AOI211_X1 U4374 ( .C1(n4348), .C2(n3564), .A(n3563), .B(n3562), .ZN(n4618)
         );
  INV_X1 U4375 ( .A(n4618), .ZN(n3565) );
  AOI21_X1 U4376 ( .B1(n4664), .B2(n4615), .A(n3565), .ZN(n3568) );
  MUX2_X1 U4377 ( .A(n3566), .B(n3568), .S(n4675), .Z(n3567) );
  OAI21_X1 U4378 ( .B1(n4613), .B2(n4485), .A(n3567), .ZN(U3483) );
  INV_X1 U4379 ( .A(REG1_REG_8__SCAN_IN), .ZN(n4934) );
  MUX2_X1 U4380 ( .A(n4934), .B(n3568), .S(n4682), .Z(n3569) );
  OAI21_X1 U4381 ( .B1(n4613), .B2(n4428), .A(n3569), .ZN(U3526) );
  XOR2_X1 U4382 ( .A(n3572), .B(n3571), .Z(n3573) );
  XNOR2_X1 U4383 ( .A(n3570), .B(n3573), .ZN(n3579) );
  INV_X1 U4384 ( .A(n3595), .ZN(n3577) );
  AOI22_X1 U4385 ( .A1(n3798), .A2(n3620), .B1(n3799), .B2(n4062), .ZN(n3574)
         );
  NAND2_X1 U4386 ( .A1(REG3_REG_12__SCAN_IN), .A2(U3149), .ZN(n4540) );
  OAI211_X1 U4387 ( .C1(n3862), .C2(n3575), .A(n3574), .B(n4540), .ZN(n3576)
         );
  AOI21_X1 U4388 ( .B1(n3577), .B2(n3866), .A(n3576), .ZN(n3578) );
  OAI21_X1 U4389 ( .B1(n3579), .B2(n3869), .A(n3578), .ZN(U3221) );
  XNOR2_X1 U4390 ( .A(n3890), .B(n3582), .ZN(n3683) );
  OAI21_X1 U4391 ( .B1(n3580), .B2(n3582), .A(n3581), .ZN(n3685) );
  NAND2_X1 U4392 ( .A1(n3685), .A2(n4277), .ZN(n3590) );
  INV_X1 U4393 ( .A(n3648), .ZN(n3584) );
  INV_X1 U4394 ( .A(n3658), .ZN(n3583) );
  OAI21_X1 U4395 ( .B1(n3584), .B2(n3704), .A(n3583), .ZN(n3690) );
  INV_X1 U4396 ( .A(n3690), .ZN(n3588) );
  AOI22_X1 U4397 ( .A1(n4281), .A2(n4062), .B1(n4279), .B2(n4061), .ZN(n3586)
         );
  AOI22_X1 U4398 ( .A1(n4612), .A2(REG2_REG_14__SCAN_IN), .B1(n3706), .B2(
        n4619), .ZN(n3585) );
  OAI211_X1 U4399 ( .C1(n3704), .C2(n4285), .A(n3586), .B(n3585), .ZN(n3587)
         );
  AOI21_X1 U4400 ( .B1(n3588), .B2(n4621), .A(n3587), .ZN(n3589) );
  OAI211_X1 U4401 ( .C1(n3683), .C2(n3591), .A(n3590), .B(n3589), .ZN(U3276)
         );
  NAND2_X1 U4402 ( .A1(n3638), .A2(n3639), .ZN(n3959) );
  XNOR2_X1 U4403 ( .A(n3592), .B(n3959), .ZN(n3618) );
  NAND2_X1 U4404 ( .A1(n3593), .A2(n3619), .ZN(n3594) );
  NAND2_X1 U4405 ( .A1(n3646), .A2(n3594), .ZN(n3633) );
  INV_X1 U4406 ( .A(REG2_REG_12__SCAN_IN), .ZN(n3596) );
  OAI22_X1 U4407 ( .A1(n4357), .A2(n3596), .B1(n3595), .B2(n4332), .ZN(n3597)
         );
  AOI21_X1 U4408 ( .B1(n3619), .B2(n4148), .A(n3597), .ZN(n3599) );
  AOI22_X1 U4409 ( .A1(n4281), .A2(n3620), .B1(n4279), .B2(n4062), .ZN(n3598)
         );
  OAI211_X1 U4410 ( .C1(n3633), .C2(n4331), .A(n3599), .B(n3598), .ZN(n3607)
         );
  INV_X1 U4411 ( .A(n3600), .ZN(n3603) );
  AOI21_X1 U4412 ( .B1(n3603), .B2(n3602), .A(n3601), .ZN(n3641) );
  INV_X1 U4413 ( .A(n3959), .ZN(n3604) );
  XNOR2_X1 U4414 ( .A(n3641), .B(n3604), .ZN(n3605) );
  NAND2_X1 U4415 ( .A1(n3605), .A2(n4348), .ZN(n3625) );
  NOR2_X1 U4416 ( .A1(n3625), .A2(n4627), .ZN(n3606) );
  AOI211_X1 U4417 ( .C1(n4277), .C2(n3618), .A(n3607), .B(n3606), .ZN(n3608)
         );
  INV_X1 U4418 ( .A(n3608), .ZN(U3278) );
  INV_X1 U4419 ( .A(REG0_REG_11__SCAN_IN), .ZN(n3612) );
  INV_X1 U4420 ( .A(n3609), .ZN(n3610) );
  AOI21_X1 U4421 ( .B1(n4664), .B2(n3611), .A(n3610), .ZN(n3614) );
  MUX2_X1 U4422 ( .A(n3612), .B(n3614), .S(n4675), .Z(n3613) );
  OAI21_X1 U4423 ( .B1(n3617), .B2(n4485), .A(n3613), .ZN(U3489) );
  INV_X1 U4424 ( .A(REG1_REG_11__SCAN_IN), .ZN(n3615) );
  MUX2_X1 U4425 ( .A(n3615), .B(n3614), .S(n4682), .Z(n3616) );
  OAI21_X1 U4426 ( .B1(n4428), .B2(n3617), .A(n3616), .ZN(U3529) );
  NAND2_X1 U4427 ( .A1(n3618), .A2(n4667), .ZN(n3627) );
  NAND2_X1 U4428 ( .A1(n3619), .A2(n4429), .ZN(n3622) );
  NAND2_X1 U4429 ( .A1(n3620), .A2(n4374), .ZN(n3621) );
  OAI211_X1 U4430 ( .C1(n3623), .C2(n4378), .A(n3622), .B(n3621), .ZN(n3624)
         );
  INV_X1 U4431 ( .A(n3624), .ZN(n3626) );
  NAND3_X1 U4432 ( .A1(n3627), .A2(n3626), .A3(n3625), .ZN(n3630) );
  MUX2_X1 U4433 ( .A(n3630), .B(REG0_REG_12__SCAN_IN), .S(n4673), .Z(n3628) );
  INV_X1 U4434 ( .A(n3628), .ZN(n3629) );
  OAI21_X1 U4435 ( .B1(n3633), .B2(n4485), .A(n3629), .ZN(U3491) );
  MUX2_X1 U4436 ( .A(REG1_REG_12__SCAN_IN), .B(n3630), .S(n4682), .Z(n3631) );
  INV_X1 U4437 ( .A(n3631), .ZN(n3632) );
  OAI21_X1 U4438 ( .B1(n4428), .B2(n3633), .A(n3632), .ZN(U3530) );
  INV_X1 U4439 ( .A(n3635), .ZN(n3636) );
  OR2_X1 U4440 ( .A1(n3637), .A2(n3636), .ZN(n3960) );
  XNOR2_X1 U4441 ( .A(n3634), .B(n3960), .ZN(n3692) );
  INV_X1 U4442 ( .A(n3692), .ZN(n3653) );
  INV_X1 U4443 ( .A(n3638), .ZN(n3640) );
  OAI21_X1 U4444 ( .B1(n3641), .B2(n3640), .A(n3639), .ZN(n3642) );
  XNOR2_X1 U4445 ( .A(n3642), .B(n3960), .ZN(n3643) );
  NAND2_X1 U4446 ( .A1(n3643), .A2(n4348), .ZN(n3645) );
  AOI22_X1 U4447 ( .A1(n3674), .A2(n4431), .B1(n4429), .B2(n3677), .ZN(n3644)
         );
  OAI211_X1 U4448 ( .C1(n3675), .C2(n4434), .A(n3645), .B(n3644), .ZN(n3691)
         );
  NAND2_X1 U4449 ( .A1(n3646), .A2(n3677), .ZN(n3647) );
  NAND2_X1 U4450 ( .A1(n3648), .A2(n3647), .ZN(n3698) );
  AOI22_X1 U4451 ( .A1(n4612), .A2(REG2_REG_13__SCAN_IN), .B1(n3649), .B2(
        n4619), .ZN(n3650) );
  OAI21_X1 U4452 ( .B1(n3698), .B2(n4331), .A(n3650), .ZN(n3651) );
  AOI21_X1 U4453 ( .B1(n3691), .B2(n4357), .A(n3651), .ZN(n3652) );
  OAI21_X1 U4454 ( .B1(n3653), .B2(n4360), .A(n3652), .ZN(U3277) );
  AOI21_X1 U4455 ( .B1(n3654), .B2(n3933), .A(n4326), .ZN(n3656) );
  NAND2_X1 U4456 ( .A1(n3656), .A2(n3655), .ZN(n3710) );
  XNOR2_X1 U4457 ( .A(n3657), .B(n3933), .ZN(n3712) );
  NAND2_X1 U4458 ( .A1(n3712), .A2(n4277), .ZN(n3666) );
  OAI21_X1 U4459 ( .B1(n3658), .B2(n3662), .A(n3723), .ZN(n3718) );
  INV_X1 U4460 ( .A(n3718), .ZN(n3664) );
  AOI22_X1 U4461 ( .A1(n4281), .A2(n3674), .B1(n4279), .B2(n3738), .ZN(n3661)
         );
  INV_X1 U4462 ( .A(n3884), .ZN(n3659) );
  AOI22_X1 U4463 ( .A1(n4612), .A2(REG2_REG_15__SCAN_IN), .B1(n3659), .B2(
        n4619), .ZN(n3660) );
  OAI211_X1 U4464 ( .C1(n3662), .C2(n4285), .A(n3661), .B(n3660), .ZN(n3663)
         );
  AOI21_X1 U4465 ( .B1(n3664), .B2(n4621), .A(n3663), .ZN(n3665) );
  OAI211_X1 U4466 ( .C1(n4612), .C2(n3710), .A(n3666), .B(n3665), .ZN(U3275)
         );
  INV_X1 U4467 ( .A(n3668), .ZN(n3670) );
  NAND2_X1 U4468 ( .A1(n3670), .A2(n3669), .ZN(n3671) );
  XNOR2_X1 U4469 ( .A(n3667), .B(n3671), .ZN(n3672) );
  NAND2_X1 U4470 ( .A1(n3672), .A2(n3874), .ZN(n3679) );
  INV_X1 U4471 ( .A(REG3_REG_13__SCAN_IN), .ZN(n3673) );
  NOR2_X1 U4472 ( .A1(STATE_REG_SCAN_IN), .A2(n3673), .ZN(n4553) );
  INV_X1 U4473 ( .A(n3674), .ZN(n3878) );
  OAI22_X1 U4474 ( .A1(n3675), .A2(n3877), .B1(n3876), .B2(n3878), .ZN(n3676)
         );
  AOI211_X1 U4475 ( .C1(n3677), .C2(n3880), .A(n4553), .B(n3676), .ZN(n3678)
         );
  OAI211_X1 U4476 ( .C1(n3885), .C2(n3680), .A(n3679), .B(n3678), .ZN(U3231)
         );
  INV_X1 U4477 ( .A(REG0_REG_14__SCAN_IN), .ZN(n4769) );
  OAI22_X1 U4478 ( .A1(n4435), .A2(n4378), .B1(n3704), .B2(n4323), .ZN(n3681)
         );
  AOI21_X1 U4479 ( .B1(n4374), .B2(n4062), .A(n3681), .ZN(n3682) );
  OAI21_X1 U4480 ( .B1(n3683), .B2(n4326), .A(n3682), .ZN(n3684) );
  AOI21_X1 U4481 ( .B1(n3685), .B2(n4667), .A(n3684), .ZN(n3687) );
  MUX2_X1 U4482 ( .A(n4769), .B(n3687), .S(n4675), .Z(n3686) );
  OAI21_X1 U4483 ( .B1(n3690), .B2(n4485), .A(n3686), .ZN(U3495) );
  INV_X1 U4484 ( .A(REG1_REG_14__SCAN_IN), .ZN(n3688) );
  MUX2_X1 U4485 ( .A(n3688), .B(n3687), .S(n4682), .Z(n3689) );
  OAI21_X1 U4486 ( .B1(n4428), .B2(n3690), .A(n3689), .ZN(U3532) );
  INV_X1 U4487 ( .A(REG1_REG_13__SCAN_IN), .ZN(n3693) );
  AOI21_X1 U4488 ( .B1(n4667), .B2(n3692), .A(n3691), .ZN(n3695) );
  MUX2_X1 U4489 ( .A(n3693), .B(n3695), .S(n4682), .Z(n3694) );
  OAI21_X1 U4490 ( .B1(n4428), .B2(n3698), .A(n3694), .ZN(U3531) );
  INV_X1 U4491 ( .A(REG0_REG_13__SCAN_IN), .ZN(n3696) );
  MUX2_X1 U4492 ( .A(n3696), .B(n3695), .S(n4675), .Z(n3697) );
  OAI21_X1 U4493 ( .B1(n3698), .B2(n4485), .A(n3697), .ZN(U3493) );
  XOR2_X1 U4494 ( .A(n3701), .B(n3700), .Z(n3702) );
  XNOR2_X1 U4495 ( .A(n3699), .B(n3702), .ZN(n3708) );
  AOI22_X1 U4496 ( .A1(n3799), .A2(n4061), .B1(n3798), .B2(n4062), .ZN(n3703)
         );
  NAND2_X1 U4497 ( .A1(REG3_REG_14__SCAN_IN), .A2(U3149), .ZN(n4560) );
  OAI211_X1 U4498 ( .C1(n3862), .C2(n3704), .A(n3703), .B(n4560), .ZN(n3705)
         );
  AOI21_X1 U4499 ( .B1(n3706), .B2(n3866), .A(n3705), .ZN(n3707) );
  OAI21_X1 U4500 ( .B1(n3708), .B2(n3869), .A(n3707), .ZN(U3212) );
  INV_X1 U4501 ( .A(REG0_REG_15__SCAN_IN), .ZN(n3713) );
  AOI22_X1 U4502 ( .A1(n3738), .A2(n4431), .B1(n4429), .B2(n3881), .ZN(n3709)
         );
  OAI211_X1 U4503 ( .C1(n3878), .C2(n4434), .A(n3710), .B(n3709), .ZN(n3711)
         );
  AOI21_X1 U4504 ( .B1(n3712), .B2(n4667), .A(n3711), .ZN(n3715) );
  MUX2_X1 U4505 ( .A(n3713), .B(n3715), .S(n4675), .Z(n3714) );
  OAI21_X1 U4506 ( .B1(n3718), .B2(n4485), .A(n3714), .ZN(U3497) );
  MUX2_X1 U4507 ( .A(n3716), .B(n3715), .S(n4682), .Z(n3717) );
  OAI21_X1 U4508 ( .B1(n4428), .B2(n3718), .A(n3717), .ZN(U3533) );
  OAI21_X1 U4509 ( .B1(n3721), .B2(n3720), .A(n3719), .ZN(n4442) );
  INV_X1 U4510 ( .A(n3722), .ZN(n3737) );
  AOI21_X1 U4511 ( .B1(n4430), .B2(n3723), .A(n3737), .ZN(n4438) );
  AOI22_X1 U4512 ( .A1(n4281), .A2(n4061), .B1(n4279), .B2(n4432), .ZN(n3726)
         );
  INV_X1 U4513 ( .A(n3724), .ZN(n3803) );
  AOI22_X1 U4514 ( .A1(n4612), .A2(REG2_REG_16__SCAN_IN), .B1(n3803), .B2(
        n4619), .ZN(n3725) );
  OAI211_X1 U4515 ( .C1(n3801), .C2(n4285), .A(n3726), .B(n3725), .ZN(n3730)
         );
  OAI211_X1 U4516 ( .C1(n3728), .C2(n3936), .A(n3727), .B(n4348), .ZN(n4439)
         );
  NOR2_X1 U4517 ( .A1(n4439), .A2(n4627), .ZN(n3729) );
  AOI211_X1 U4518 ( .C1(n4438), .C2(n4621), .A(n3730), .B(n3729), .ZN(n3731)
         );
  OAI21_X1 U4519 ( .B1(n4442), .B2(n4360), .A(n3731), .ZN(U3274) );
  INV_X1 U4520 ( .A(n3891), .ZN(n3732) );
  NAND2_X1 U4521 ( .A1(n3732), .A2(n4316), .ZN(n3961) );
  XNOR2_X1 U4522 ( .A(n3733), .B(n3961), .ZN(n3734) );
  NAND2_X1 U4523 ( .A1(n3734), .A2(n4348), .ZN(n4423) );
  XOR2_X1 U4524 ( .A(n3961), .B(n3735), .Z(n4426) );
  NAND2_X1 U4525 ( .A1(n4426), .A2(n4277), .ZN(n3745) );
  INV_X1 U4526 ( .A(n4352), .ZN(n3736) );
  OAI21_X1 U4527 ( .B1(n3737), .B2(n3741), .A(n3736), .ZN(n4486) );
  INV_X1 U4528 ( .A(n4486), .ZN(n3743) );
  AOI22_X1 U4529 ( .A1(n4281), .A2(n3738), .B1(n4279), .B2(n4421), .ZN(n3740)
         );
  AOI22_X1 U4530 ( .A1(n4612), .A2(REG2_REG_17__SCAN_IN), .B1(n3811), .B2(
        n4619), .ZN(n3739) );
  OAI211_X1 U4531 ( .C1(n3741), .C2(n4285), .A(n3740), .B(n3739), .ZN(n3742)
         );
  AOI21_X1 U4532 ( .B1(n3743), .B2(n4621), .A(n3742), .ZN(n3744) );
  OAI211_X1 U4533 ( .C1(n4627), .C2(n4423), .A(n3745), .B(n3744), .ZN(U3273)
         );
  NAND3_X1 U4534 ( .A1(n2345), .A2(IR_REG_31__SCAN_IN), .A3(STATE_REG_SCAN_IN), 
        .ZN(n3746) );
  INV_X1 U4535 ( .A(DATAI_31_), .ZN(n4902) );
  OAI22_X1 U4536 ( .A1(n2350), .A2(n3746), .B1(STATE_REG_SCAN_IN), .B2(n4902), 
        .ZN(U3321) );
  XNOR2_X1 U4537 ( .A(n3748), .B(n3747), .ZN(n3753) );
  INV_X1 U4538 ( .A(n3749), .ZN(n4175) );
  INV_X1 U4539 ( .A(REG3_REG_27__SCAN_IN), .ZN(n4908) );
  OAI22_X1 U4540 ( .A1(n3862), .A2(n4178), .B1(STATE_REG_SCAN_IN), .B2(n4908), 
        .ZN(n3751) );
  OAI22_X1 U4541 ( .A1(n4146), .A2(n3876), .B1(n3877), .B2(n4379), .ZN(n3750)
         );
  AOI211_X1 U4542 ( .C1(n4175), .C2(n3866), .A(n3751), .B(n3750), .ZN(n3752)
         );
  OAI21_X1 U4543 ( .B1(n3753), .B2(n3869), .A(n3752), .ZN(U3211) );
  NAND2_X1 U4544 ( .A1(n3754), .A2(n3755), .ZN(n3838) );
  NAND2_X1 U4545 ( .A1(n3838), .A2(n3756), .ZN(n3757) );
  NAND2_X1 U4546 ( .A1(n3757), .A2(n3874), .ZN(n3766) );
  AOI21_X1 U4547 ( .B1(n3838), .B2(n3759), .A(n3758), .ZN(n3765) );
  OAI22_X1 U4548 ( .A1(n3862), .A2(n3761), .B1(STATE_REG_SCAN_IN), .B2(n3760), 
        .ZN(n3763) );
  OAI22_X1 U4549 ( .A1(n3780), .A2(n3877), .B1(n3876), .B2(n4245), .ZN(n3762)
         );
  AOI211_X1 U4550 ( .C1(n4249), .C2(n3866), .A(n3763), .B(n3762), .ZN(n3764)
         );
  OAI21_X1 U4551 ( .B1(n3766), .B2(n3765), .A(n3764), .ZN(U3213) );
  XNOR2_X1 U4552 ( .A(n3767), .B(n3768), .ZN(n3769) );
  NAND2_X1 U4553 ( .A1(n3769), .A2(n3874), .ZN(n3773) );
  AND2_X1 U4554 ( .A1(U3149), .A2(REG3_REG_19__SCAN_IN), .ZN(n4131) );
  OAI22_X1 U4555 ( .A1(n2953), .A2(n3877), .B1(n3876), .B2(n4404), .ZN(n3770)
         );
  AOI211_X1 U4556 ( .C1(n3771), .C2(n3880), .A(n4131), .B(n3770), .ZN(n3772)
         );
  OAI211_X1 U4557 ( .C1(n3885), .C2(n4333), .A(n3773), .B(n3772), .ZN(U3216)
         );
  XNOR2_X1 U4558 ( .A(n3776), .B(n3775), .ZN(n3777) );
  XNOR2_X1 U4559 ( .A(n3774), .B(n3777), .ZN(n3784) );
  INV_X1 U4560 ( .A(n3778), .ZN(n4282) );
  OAI22_X1 U4561 ( .A1(n3862), .A2(n4286), .B1(STATE_REG_SCAN_IN), .B2(n3779), 
        .ZN(n3782) );
  OAI22_X1 U4562 ( .A1(n4404), .A2(n3877), .B1(n3876), .B2(n3780), .ZN(n3781)
         );
  AOI211_X1 U4563 ( .C1(n4282), .C2(n3866), .A(n3782), .B(n3781), .ZN(n3783)
         );
  OAI21_X1 U4564 ( .B1(n3784), .B2(n3869), .A(n3783), .ZN(U3220) );
  NAND2_X1 U4565 ( .A1(n3786), .A2(n3785), .ZN(n3788) );
  XOR2_X1 U4566 ( .A(n3788), .B(n3787), .Z(n3793) );
  OAI22_X1 U4567 ( .A1(n3862), .A2(n4216), .B1(STATE_REG_SCAN_IN), .B2(n3789), 
        .ZN(n3791) );
  OAI22_X1 U4568 ( .A1(n4245), .A2(n3877), .B1(n3876), .B2(n4379), .ZN(n3790)
         );
  AOI211_X1 U4569 ( .C1(n4213), .C2(n3866), .A(n3791), .B(n3790), .ZN(n3792)
         );
  OAI21_X1 U4570 ( .B1(n3793), .B2(n3869), .A(n3792), .ZN(U3222) );
  INV_X1 U4571 ( .A(n3871), .ZN(n3795) );
  OAI21_X1 U4572 ( .B1(n3795), .B2(n3872), .A(n3794), .ZN(n3796) );
  XOR2_X1 U4573 ( .A(n3797), .B(n3796), .Z(n3805) );
  AOI22_X1 U4574 ( .A1(n3799), .A2(n4432), .B1(n3798), .B2(n4061), .ZN(n3800)
         );
  NAND2_X1 U4575 ( .A1(REG3_REG_16__SCAN_IN), .A2(U3149), .ZN(n4580) );
  OAI211_X1 U4576 ( .C1(n3862), .C2(n3801), .A(n3800), .B(n4580), .ZN(n3802)
         );
  AOI21_X1 U4577 ( .B1(n3803), .B2(n3866), .A(n3802), .ZN(n3804) );
  OAI21_X1 U4578 ( .B1(n3805), .B2(n3869), .A(n3804), .ZN(U3223) );
  XNOR2_X1 U4579 ( .A(n3808), .B(n3807), .ZN(n3809) );
  XNOR2_X1 U4580 ( .A(n3806), .B(n3809), .ZN(n3814) );
  NOR2_X1 U4581 ( .A1(STATE_REG_SCAN_IN), .A2(n2680), .ZN(n4593) );
  OAI22_X1 U4582 ( .A1(n4424), .A2(n3877), .B1(n3876), .B2(n2953), .ZN(n3810)
         );
  AOI211_X1 U4583 ( .C1(n4420), .C2(n3880), .A(n4593), .B(n3810), .ZN(n3813)
         );
  NAND2_X1 U4584 ( .A1(n3866), .A2(n3811), .ZN(n3812) );
  OAI211_X1 U4585 ( .C1(n3814), .C2(n3869), .A(n3813), .B(n3812), .ZN(U3225)
         );
  NAND2_X1 U4586 ( .A1(n3815), .A2(n3816), .ZN(n3817) );
  XOR2_X1 U4587 ( .A(n3818), .B(n3817), .Z(n3824) );
  INV_X1 U4588 ( .A(n3819), .ZN(n4228) );
  OAI22_X1 U4589 ( .A1(n3862), .A2(n4231), .B1(STATE_REG_SCAN_IN), .B2(n3820), 
        .ZN(n3822) );
  INV_X1 U4590 ( .A(n4385), .ZN(n3863) );
  OAI22_X1 U4591 ( .A1(n4388), .A2(n3877), .B1(n3876), .B2(n3863), .ZN(n3821)
         );
  AOI211_X1 U4592 ( .C1(n4228), .C2(n3866), .A(n3822), .B(n3821), .ZN(n3823)
         );
  OAI21_X1 U4593 ( .B1(n3824), .B2(n3869), .A(n3823), .ZN(U3226) );
  INV_X1 U4594 ( .A(n3825), .ZN(n3830) );
  AOI21_X1 U4595 ( .B1(n3829), .B2(n3827), .A(n3826), .ZN(n3828) );
  AOI21_X1 U4596 ( .B1(n3830), .B2(n3829), .A(n3828), .ZN(n3836) );
  INV_X1 U4597 ( .A(n3831), .ZN(n4310) );
  OAI22_X1 U4598 ( .A1(n3862), .A2(n4308), .B1(STATE_REG_SCAN_IN), .B2(n3832), 
        .ZN(n3834) );
  OAI22_X1 U4599 ( .A1(n3852), .A2(n3877), .B1(n3876), .B2(n4300), .ZN(n3833)
         );
  AOI211_X1 U4600 ( .C1(n4310), .C2(n3866), .A(n3834), .B(n3833), .ZN(n3835)
         );
  OAI21_X1 U4601 ( .B1(n3836), .B2(n3869), .A(n3835), .ZN(U3230) );
  NAND2_X1 U4602 ( .A1(n3754), .A2(n3837), .ZN(n3840) );
  INV_X1 U4603 ( .A(n3838), .ZN(n3839) );
  AOI21_X1 U4604 ( .B1(n3841), .B2(n3840), .A(n3839), .ZN(n3846) );
  INV_X1 U4605 ( .A(n3842), .ZN(n4268) );
  INV_X1 U4606 ( .A(REG3_REG_22__SCAN_IN), .ZN(n4877) );
  OAI22_X1 U4607 ( .A1(n3862), .A2(n4265), .B1(STATE_REG_SCAN_IN), .B2(n4877), 
        .ZN(n3844) );
  OAI22_X1 U4608 ( .A1(n4388), .A2(n3876), .B1(n3877), .B2(n4300), .ZN(n3843)
         );
  AOI211_X1 U4609 ( .C1(n4268), .C2(n3866), .A(n3844), .B(n3843), .ZN(n3845)
         );
  OAI21_X1 U4610 ( .B1(n3846), .B2(n3869), .A(n3845), .ZN(U3232) );
  INV_X1 U4611 ( .A(n3847), .ZN(n3849) );
  NOR2_X1 U4612 ( .A1(n3849), .A2(n3848), .ZN(n3850) );
  XNOR2_X1 U4613 ( .A(n3851), .B(n3850), .ZN(n3856) );
  NOR2_X1 U4614 ( .A1(STATE_REG_SCAN_IN), .A2(n4926), .ZN(n4603) );
  OAI22_X1 U4615 ( .A1(n3852), .A2(n3876), .B1(n3877), .B2(n4346), .ZN(n3853)
         );
  AOI211_X1 U4616 ( .C1(n4343), .C2(n3880), .A(n4603), .B(n3853), .ZN(n3855)
         );
  NAND2_X1 U4617 ( .A1(n3866), .A2(n4353), .ZN(n3854) );
  OAI211_X1 U4618 ( .C1(n3856), .C2(n3869), .A(n3855), .B(n3854), .ZN(U3235)
         );
  NOR2_X1 U4619 ( .A1(n2300), .A2(n3859), .ZN(n3860) );
  XNOR2_X1 U4620 ( .A(n3857), .B(n3860), .ZN(n3870) );
  INV_X1 U4621 ( .A(n4198), .ZN(n3867) );
  OAI22_X1 U4622 ( .A1(n3862), .A2(n4196), .B1(STATE_REG_SCAN_IN), .B2(n3861), 
        .ZN(n3865) );
  OAI22_X1 U4623 ( .A1(n4195), .A2(n3876), .B1(n3877), .B2(n3863), .ZN(n3864)
         );
  AOI211_X1 U4624 ( .C1(n3867), .C2(n3866), .A(n3865), .B(n3864), .ZN(n3868)
         );
  OAI21_X1 U4625 ( .B1(n3870), .B2(n3869), .A(n3868), .ZN(U3237) );
  NAND2_X1 U4626 ( .A1(n3794), .A2(n3871), .ZN(n3873) );
  XNOR2_X1 U4627 ( .A(n3873), .B(n3872), .ZN(n3875) );
  NAND2_X1 U4628 ( .A1(n3875), .A2(n3874), .ZN(n3883) );
  AND2_X1 U4629 ( .A1(U3149), .A2(REG3_REG_15__SCAN_IN), .ZN(n4574) );
  OAI22_X1 U4630 ( .A1(n3878), .A2(n3877), .B1(n3876), .B2(n4424), .ZN(n3879)
         );
  AOI211_X1 U4631 ( .C1(n3881), .C2(n3880), .A(n4574), .B(n3879), .ZN(n3882)
         );
  OAI211_X1 U4632 ( .C1(n3885), .C2(n3884), .A(n3883), .B(n3882), .ZN(U3238)
         );
  NAND2_X1 U4633 ( .A1(n3889), .A2(n3886), .ZN(n4018) );
  NAND2_X1 U4634 ( .A1(n3888), .A2(n3887), .ZN(n4000) );
  NAND2_X1 U4635 ( .A1(n4000), .A2(n3889), .ZN(n4019) );
  OAI21_X1 U4636 ( .B1(n3890), .B2(n4018), .A(n4019), .ZN(n3894) );
  INV_X1 U4637 ( .A(n4023), .ZN(n3893) );
  OR2_X1 U4638 ( .A1(n3892), .A2(n3891), .ZN(n4026) );
  AOI211_X1 U4639 ( .C1(n3894), .C2(n4027), .A(n3893), .B(n4026), .ZN(n3896)
         );
  INV_X1 U4640 ( .A(n3895), .ZN(n4030) );
  NOR3_X1 U4641 ( .A1(n3896), .A2(n4030), .A3(n4032), .ZN(n3901) );
  INV_X1 U4642 ( .A(n3897), .ZN(n3900) );
  INV_X1 U4643 ( .A(n3932), .ZN(n3898) );
  OR2_X1 U4644 ( .A1(n3939), .A2(n3898), .ZN(n4035) );
  INV_X1 U4645 ( .A(n4035), .ZN(n3899) );
  OAI21_X1 U4646 ( .B1(n3901), .B2(n3900), .A(n3899), .ZN(n3911) );
  OR2_X1 U4647 ( .A1(n3903), .A2(n3902), .ZN(n3917) );
  INV_X1 U4648 ( .A(REG1_REG_31__SCAN_IN), .ZN(n4361) );
  NAND2_X1 U4649 ( .A1(n3904), .A2(REG2_REG_31__SCAN_IN), .ZN(n3907) );
  NAND2_X1 U4650 ( .A1(n3905), .A2(REG0_REG_31__SCAN_IN), .ZN(n3906) );
  OAI211_X1 U4651 ( .C1(n3908), .C2(n4361), .A(n3907), .B(n3906), .ZN(n4139)
         );
  AND2_X1 U4652 ( .A1(n3909), .A2(DATAI_31_), .ZN(n3925) );
  INV_X1 U4653 ( .A(n3925), .ZN(n4140) );
  AND2_X1 U4654 ( .A1(n4139), .A2(n4140), .ZN(n4045) );
  AND2_X1 U4655 ( .A1(n3909), .A2(DATAI_30_), .ZN(n4366) );
  INV_X1 U4656 ( .A(n4366), .ZN(n3921) );
  NOR2_X1 U4657 ( .A1(n3923), .A2(n3921), .ZN(n3910) );
  NOR2_X1 U4658 ( .A1(n4045), .A2(n3910), .ZN(n3944) );
  OAI21_X1 U4659 ( .B1(n4160), .B2(n3912), .A(n3944), .ZN(n3916) );
  AOI211_X1 U4660 ( .C1(n4187), .C2(n3911), .A(n3917), .B(n3916), .ZN(n3920)
         );
  INV_X1 U4661 ( .A(n4036), .ZN(n3919) );
  NAND2_X1 U4662 ( .A1(n4160), .A2(n3912), .ZN(n3913) );
  AND2_X1 U4663 ( .A1(n3914), .A2(n3913), .ZN(n4039) );
  NAND3_X1 U4664 ( .A1(n3945), .A2(n4039), .A3(n3915), .ZN(n3918) );
  AOI21_X1 U4665 ( .B1(n4039), .B2(n3917), .A(n3916), .ZN(n4044) );
  AOI22_X1 U4666 ( .A1(n3920), .A2(n3919), .B1(n3918), .B2(n4044), .ZN(n3930)
         );
  NOR2_X1 U4667 ( .A1(n4139), .A2(n3921), .ZN(n3929) );
  INV_X1 U4668 ( .A(n3922), .ZN(n3928) );
  INV_X1 U4669 ( .A(n3923), .ZN(n3924) );
  NOR2_X1 U4670 ( .A1(n3924), .A2(n4366), .ZN(n3943) );
  INV_X1 U4671 ( .A(n4139), .ZN(n3926) );
  OAI21_X1 U4672 ( .B1(n3943), .B2(n3926), .A(n3925), .ZN(n3927) );
  OAI211_X1 U4673 ( .C1(n3930), .C2(n3929), .A(n3928), .B(n3927), .ZN(n4053)
         );
  NAND2_X1 U4674 ( .A1(n3932), .A2(n3931), .ZN(n4241) );
  INV_X1 U4675 ( .A(n4259), .ZN(n4257) );
  INV_X1 U4676 ( .A(n3933), .ZN(n3934) );
  NAND4_X1 U4677 ( .A1(n4257), .A2(n3936), .A3(n3935), .A4(n3934), .ZN(n3951)
         );
  NAND2_X1 U4678 ( .A1(n4185), .A2(n3937), .ZN(n4208) );
  INV_X1 U4679 ( .A(n4208), .ZN(n3949) );
  INV_X1 U4680 ( .A(n4203), .ZN(n3938) );
  OR2_X1 U4681 ( .A1(n3939), .A2(n3938), .ZN(n4225) );
  INV_X1 U4682 ( .A(n4225), .ZN(n4221) );
  XNOR2_X1 U4683 ( .A(n4280), .B(n4308), .ZN(n4292) );
  INV_X1 U4684 ( .A(n4292), .ZN(n4296) );
  NAND2_X1 U4685 ( .A1(n3941), .A2(n3940), .ZN(n4322) );
  NOR2_X1 U4686 ( .A1(n4139), .A2(n4140), .ZN(n3942) );
  NOR2_X1 U4687 ( .A1(n3943), .A2(n3942), .ZN(n4046) );
  NAND4_X1 U4688 ( .A1(n3946), .A2(n3945), .A3(n3944), .A4(n4046), .ZN(n3947)
         );
  NOR4_X1 U4689 ( .A1(n4651), .A2(n4322), .A3(n4489), .A4(n3947), .ZN(n3948)
         );
  NAND4_X1 U4690 ( .A1(n3949), .A2(n4221), .A3(n4296), .A4(n3948), .ZN(n3950)
         );
  XNOR2_X1 U4691 ( .A(n4379), .B(n4196), .ZN(n4188) );
  INV_X1 U4692 ( .A(n3953), .ZN(n4029) );
  INV_X1 U4693 ( .A(n4276), .ZN(n3957) );
  NOR4_X1 U4694 ( .A1(n3957), .A2(n3956), .A3(n3955), .A4(n3954), .ZN(n3972)
         );
  NOR4_X1 U4695 ( .A1(n3961), .A2(n3960), .A3(n3959), .A4(n3958), .ZN(n3971)
         );
  INV_X1 U4696 ( .A(n3962), .ZN(n3965) );
  NOR4_X1 U4697 ( .A1(n3965), .A2(n3964), .A3(n4342), .A4(n3963), .ZN(n3970)
         );
  INV_X1 U4698 ( .A(n2965), .ZN(n3966) );
  AND4_X1 U4699 ( .A1(n3968), .A2(n2934), .A3(n3967), .A4(n3966), .ZN(n3969)
         );
  AND4_X1 U4700 ( .A1(n3972), .A2(n3971), .A3(n3970), .A4(n3969), .ZN(n3973)
         );
  NAND3_X1 U4701 ( .A1(n3974), .A2(n4188), .A3(n3973), .ZN(n4051) );
  NOR2_X1 U4702 ( .A1(n4195), .A2(n3975), .ZN(n4043) );
  INV_X1 U4703 ( .A(n3976), .ZN(n3979) );
  OAI211_X1 U4704 ( .C1(n3979), .C2(n4489), .A(n3978), .B(n3977), .ZN(n3982)
         );
  NAND3_X1 U4705 ( .A1(n3982), .A2(n3981), .A3(n3980), .ZN(n3985) );
  NAND3_X1 U4706 ( .A1(n3985), .A2(n3984), .A3(n3983), .ZN(n3988) );
  NAND3_X1 U4707 ( .A1(n3988), .A2(n3987), .A3(n3986), .ZN(n3991) );
  NAND4_X1 U4708 ( .A1(n3991), .A2(n3990), .A3(n3989), .A4(n4004), .ZN(n3994)
         );
  AND3_X1 U4709 ( .A1(n3994), .A2(n3993), .A3(n3992), .ZN(n3999) );
  NAND2_X1 U4710 ( .A1(n3996), .A2(n3995), .ZN(n4007) );
  OAI211_X1 U4711 ( .C1(n3999), .C2(n4007), .A(n3998), .B(n3997), .ZN(n4003)
         );
  INV_X1 U4712 ( .A(n4000), .ZN(n4002) );
  NAND3_X1 U4713 ( .A1(n4003), .A2(n4002), .A3(n4001), .ZN(n4017) );
  INV_X1 U4714 ( .A(n4004), .ZN(n4008) );
  NOR4_X1 U4715 ( .A1(n4008), .A2(n4007), .A3(n4006), .A4(n4005), .ZN(n4011)
         );
  INV_X1 U4716 ( .A(n4009), .ZN(n4010) );
  OAI21_X1 U4717 ( .B1(n4011), .B2(n4010), .A(n4019), .ZN(n4016) );
  INV_X1 U4718 ( .A(n4012), .ZN(n4015) );
  INV_X1 U4719 ( .A(n4013), .ZN(n4014) );
  AOI211_X1 U4720 ( .C1(n4017), .C2(n4016), .A(n4015), .B(n4014), .ZN(n4025)
         );
  INV_X1 U4721 ( .A(n4018), .ZN(n4021) );
  INV_X1 U4722 ( .A(n4019), .ZN(n4020) );
  AOI21_X1 U4723 ( .B1(n4022), .B2(n4021), .A(n4020), .ZN(n4024) );
  OAI21_X1 U4724 ( .B1(n4025), .B2(n4024), .A(n4023), .ZN(n4028) );
  AOI21_X1 U4725 ( .B1(n4028), .B2(n4027), .A(n4026), .ZN(n4031) );
  OAI21_X1 U4726 ( .B1(n4031), .B2(n4030), .A(n4029), .ZN(n4034) );
  INV_X1 U4727 ( .A(n4032), .ZN(n4033) );
  NAND2_X1 U4728 ( .A1(n4034), .A2(n4033), .ZN(n4037) );
  AOI211_X1 U4729 ( .C1(n4038), .C2(n4037), .A(n4036), .B(n4035), .ZN(n4042)
         );
  INV_X1 U4730 ( .A(n4039), .ZN(n4040) );
  NOR4_X1 U4731 ( .A1(n4043), .A2(n4042), .A3(n4041), .A4(n4040), .ZN(n4048)
         );
  INV_X1 U4732 ( .A(n4044), .ZN(n4047) );
  OAI22_X1 U4733 ( .A1(n4048), .A2(n4047), .B1(n4046), .B2(n4045), .ZN(n4050)
         );
  MUX2_X1 U4734 ( .A(n4051), .B(n4050), .S(n4049), .Z(n4052) );
  NAND2_X1 U4735 ( .A1(n4053), .A2(n4052), .ZN(n4054) );
  XNOR2_X1 U4736 ( .A(n4054), .B(n4490), .ZN(n4060) );
  NAND2_X1 U4737 ( .A1(n2180), .A2(n4055), .ZN(n4056) );
  OAI211_X1 U4738 ( .C1(n4057), .C2(n4059), .A(n4056), .B(B_REG_SCAN_IN), .ZN(
        n4058) );
  OAI21_X1 U4739 ( .B1(n4060), .B2(n4059), .A(n4058), .ZN(U3239) );
  MUX2_X1 U4740 ( .A(n4139), .B(DATAO_REG_31__SCAN_IN), .S(n4975), .Z(U3581)
         );
  MUX2_X1 U4741 ( .A(n4160), .B(DATAO_REG_29__SCAN_IN), .S(n4975), .Z(U3579)
         );
  MUX2_X1 U4742 ( .A(n4161), .B(DATAO_REG_27__SCAN_IN), .S(n4975), .Z(U3577)
         );
  MUX2_X1 U4743 ( .A(n4212), .B(DATAO_REG_26__SCAN_IN), .S(n4975), .Z(U3576)
         );
  MUX2_X1 U4744 ( .A(n4385), .B(DATAO_REG_25__SCAN_IN), .S(n4975), .Z(U3575)
         );
  MUX2_X1 U4745 ( .A(n4375), .B(DATAO_REG_24__SCAN_IN), .S(n4975), .Z(U3574)
         );
  MUX2_X1 U4746 ( .A(n4401), .B(DATAO_REG_22__SCAN_IN), .S(n4975), .Z(U3572)
         );
  MUX2_X1 U4747 ( .A(n4061), .B(DATAO_REG_15__SCAN_IN), .S(n4975), .Z(U3565)
         );
  MUX2_X1 U4748 ( .A(DATAO_REG_13__SCAN_IN), .B(n4062), .S(U4043), .Z(U3563)
         );
  MUX2_X1 U4749 ( .A(n4063), .B(DATAO_REG_10__SCAN_IN), .S(n4975), .Z(U3560)
         );
  MUX2_X1 U4750 ( .A(n4064), .B(DATAO_REG_9__SCAN_IN), .S(n4975), .Z(U3559) );
  MUX2_X1 U4751 ( .A(n4065), .B(DATAO_REG_7__SCAN_IN), .S(n4975), .Z(U3557) );
  MUX2_X1 U4752 ( .A(n4066), .B(DATAO_REG_6__SCAN_IN), .S(n4975), .Z(U3556) );
  MUX2_X1 U4753 ( .A(n4067), .B(DATAO_REG_4__SCAN_IN), .S(n4975), .Z(U3554) );
  MUX2_X1 U4754 ( .A(n4068), .B(DATAO_REG_2__SCAN_IN), .S(n4975), .Z(U3552) );
  MUX2_X1 U4755 ( .A(n2928), .B(DATAO_REG_1__SCAN_IN), .S(n4975), .Z(U3551) );
  NAND2_X1 U4756 ( .A1(IR_REG_0__SCAN_IN), .A2(REG1_REG_0__SCAN_IN), .ZN(n4072) );
  AOI211_X1 U4757 ( .C1(n4072), .C2(n4071), .A(n4070), .B(n4069), .ZN(n4073)
         );
  INV_X1 U4758 ( .A(n4073), .ZN(n4082) );
  AOI22_X1 U4759 ( .A1(n4604), .A2(ADDR_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(U3149), .ZN(n4081) );
  NAND2_X1 U4760 ( .A1(n4074), .A2(n3116), .ZN(n4080) );
  MUX2_X1 U4761 ( .A(REG2_REG_1__SCAN_IN), .B(n4075), .S(n3116), .Z(n4077) );
  OAI211_X1 U4762 ( .C1(n4078), .C2(n4077), .A(n4549), .B(n4076), .ZN(n4079)
         );
  NAND4_X1 U4763 ( .A1(n4082), .A2(n4081), .A3(n4080), .A4(n4079), .ZN(U3241)
         );
  INV_X1 U4764 ( .A(REG2_REG_19__SCAN_IN), .ZN(n4083) );
  MUX2_X1 U4765 ( .A(REG2_REG_19__SCAN_IN), .B(n4083), .S(n4490), .Z(n4102) );
  INV_X1 U4766 ( .A(REG2_REG_18__SCAN_IN), .ZN(n4084) );
  AOI22_X1 U4767 ( .A1(REG2_REG_18__SCAN_IN), .A2(n4632), .B1(n4103), .B2(
        n4084), .ZN(n4602) );
  NOR2_X1 U4768 ( .A1(n4633), .A2(REG2_REG_17__SCAN_IN), .ZN(n4085) );
  AOI21_X1 U4769 ( .B1(REG2_REG_17__SCAN_IN), .B2(n4633), .A(n4085), .ZN(n4591) );
  NAND2_X1 U4770 ( .A1(REG2_REG_11__SCAN_IN), .A2(n4115), .ZN(n4092) );
  AOI22_X1 U4771 ( .A1(REG2_REG_11__SCAN_IN), .A2(n4115), .B1(n4643), .B2(
        n3522), .ZN(n4532) );
  NAND2_X1 U4772 ( .A1(n4110), .A2(REG2_REG_9__SCAN_IN), .ZN(n4089) );
  INV_X1 U4773 ( .A(n4110), .ZN(n4646) );
  AOI22_X1 U4774 ( .A1(n4110), .A2(REG2_REG_9__SCAN_IN), .B1(n4950), .B2(n4646), .ZN(n4512) );
  INV_X1 U4775 ( .A(REG2_REG_8__SCAN_IN), .ZN(n4087) );
  OAI22_X1 U4776 ( .A1(n4088), .A2(n4087), .B1(n4086), .B2(n4106), .ZN(n4511)
         );
  NAND2_X1 U4777 ( .A1(n4512), .A2(n4511), .ZN(n4510) );
  NAND2_X1 U4778 ( .A1(n4089), .A2(n4510), .ZN(n4090) );
  NAND2_X1 U4779 ( .A1(n4112), .A2(n4090), .ZN(n4091) );
  INV_X1 U4780 ( .A(n4112), .ZN(n4644) );
  XNOR2_X1 U4781 ( .A(n4090), .B(n4644), .ZN(n4521) );
  NAND2_X1 U4782 ( .A1(REG2_REG_10__SCAN_IN), .A2(n4521), .ZN(n4520) );
  NAND2_X1 U4783 ( .A1(n4091), .A2(n4520), .ZN(n4531) );
  NAND2_X1 U4784 ( .A1(n4532), .A2(n4531), .ZN(n4530) );
  NAND2_X1 U4785 ( .A1(n4092), .A2(n4530), .ZN(n4093) );
  NAND2_X1 U4786 ( .A1(n4117), .A2(n4093), .ZN(n4094) );
  INV_X1 U4787 ( .A(REG2_REG_13__SCAN_IN), .ZN(n4547) );
  NAND2_X1 U4788 ( .A1(n4547), .A2(n4640), .ZN(n4095) );
  NOR2_X1 U4789 ( .A1(n4096), .A2(n4569), .ZN(n4097) );
  INV_X1 U4790 ( .A(REG2_REG_14__SCAN_IN), .ZN(n4810) );
  XOR2_X1 U4791 ( .A(n4096), .B(n4638), .Z(n4562) );
  NOR2_X1 U4792 ( .A1(n4810), .A2(n4562), .ZN(n4561) );
  NOR2_X1 U4793 ( .A1(n4097), .A2(n4561), .ZN(n4572) );
  NAND2_X1 U4794 ( .A1(REG2_REG_15__SCAN_IN), .A2(n4104), .ZN(n4098) );
  OAI21_X1 U4795 ( .B1(REG2_REG_15__SCAN_IN), .B2(n4104), .A(n4098), .ZN(n4571) );
  NOR2_X1 U4796 ( .A1(n4572), .A2(n4571), .ZN(n4570) );
  INV_X1 U4797 ( .A(n4125), .ZN(n4636) );
  NAND2_X1 U4798 ( .A1(n4099), .A2(n4636), .ZN(n4100) );
  INV_X1 U4799 ( .A(REG2_REG_16__SCAN_IN), .ZN(n4952) );
  NAND2_X1 U4800 ( .A1(n4591), .A2(n4589), .ZN(n4590) );
  AOI21_X1 U4801 ( .B1(n4103), .B2(REG2_REG_18__SCAN_IN), .A(n4601), .ZN(n4101) );
  XOR2_X1 U4802 ( .A(n4102), .B(n4101), .Z(n4137) );
  INV_X1 U4803 ( .A(REG1_REG_18__SCAN_IN), .ZN(n4791) );
  AOI22_X1 U4804 ( .A1(REG1_REG_18__SCAN_IN), .A2(n4103), .B1(n4632), .B2(
        n4791), .ZN(n4607) );
  NOR2_X1 U4805 ( .A1(n4633), .A2(REG1_REG_17__SCAN_IN), .ZN(n4128) );
  NAND2_X1 U4806 ( .A1(REG1_REG_15__SCAN_IN), .A2(n4104), .ZN(n4123) );
  INV_X1 U4807 ( .A(n4104), .ZN(n4637) );
  AOI22_X1 U4808 ( .A1(REG1_REG_15__SCAN_IN), .A2(n4104), .B1(n4637), .B2(
        n3716), .ZN(n4577) );
  NAND2_X1 U4809 ( .A1(n4110), .A2(REG1_REG_9__SCAN_IN), .ZN(n4111) );
  INV_X1 U4810 ( .A(n4105), .ZN(n4107) );
  INV_X1 U4811 ( .A(REG1_REG_9__SCAN_IN), .ZN(n4109) );
  AOI22_X1 U4812 ( .A1(n4110), .A2(REG1_REG_9__SCAN_IN), .B1(n4109), .B2(n4646), .ZN(n4509) );
  NAND2_X1 U4813 ( .A1(n4112), .A2(n4113), .ZN(n4114) );
  NAND2_X1 U4814 ( .A1(n4114), .A2(n4518), .ZN(n4528) );
  AOI22_X1 U4815 ( .A1(REG1_REG_11__SCAN_IN), .A2(n4115), .B1(n4643), .B2(
        n3615), .ZN(n4529) );
  NAND2_X1 U4816 ( .A1(n4528), .A2(n4529), .ZN(n4527) );
  NAND2_X1 U4817 ( .A1(REG1_REG_11__SCAN_IN), .A2(n4115), .ZN(n4116) );
  NAND2_X1 U4818 ( .A1(n4117), .A2(n4118), .ZN(n4119) );
  XNOR2_X1 U4819 ( .A(n4118), .B(n4641), .ZN(n4544) );
  AOI22_X1 U4820 ( .A1(REG1_REG_13__SCAN_IN), .A2(n4548), .B1(n4640), .B2(
        n3693), .ZN(n4557) );
  NAND2_X1 U4821 ( .A1(REG1_REG_13__SCAN_IN), .A2(n4548), .ZN(n4120) );
  NAND2_X1 U4822 ( .A1(n4638), .A2(n4121), .ZN(n4122) );
  XNOR2_X1 U4823 ( .A(n4121), .B(n4569), .ZN(n4566) );
  NAND2_X1 U4824 ( .A1(REG1_REG_14__SCAN_IN), .A2(n4566), .ZN(n4565) );
  NOR2_X1 U4825 ( .A1(REG1_REG_16__SCAN_IN), .A2(n4585), .ZN(n4586) );
  NOR2_X1 U4826 ( .A1(n4125), .A2(n4124), .ZN(n4126) );
  INV_X1 U4827 ( .A(REG1_REG_17__SCAN_IN), .ZN(n4127) );
  AOI22_X1 U4828 ( .A1(n4633), .A2(n4127), .B1(REG1_REG_17__SCAN_IN), .B2(
        n4599), .ZN(n4594) );
  OAI21_X1 U4829 ( .B1(n4791), .B2(n4632), .A(n4605), .ZN(n4130) );
  MUX2_X1 U4830 ( .A(n4415), .B(REG1_REG_19__SCAN_IN), .S(n4490), .Z(n4129) );
  XNOR2_X1 U4831 ( .A(n4130), .B(n4129), .ZN(n4135) );
  AOI21_X1 U4832 ( .B1(n4604), .B2(ADDR_REG_19__SCAN_IN), .A(n4131), .ZN(n4132) );
  OAI21_X1 U4833 ( .B1(n4610), .B2(n4133), .A(n4132), .ZN(n4134) );
  AOI21_X1 U4834 ( .B1(n4135), .B2(n4606), .A(n4134), .ZN(n4136) );
  OAI21_X1 U4835 ( .B1(n4137), .B2(n4600), .A(n4136), .ZN(U3259) );
  XNOR2_X1 U4836 ( .A(n4364), .B(n4140), .ZN(n4446) );
  NAND2_X1 U4837 ( .A1(n4139), .A2(n4138), .ZN(n4368) );
  OAI21_X1 U4838 ( .B1(n4140), .B2(n4323), .A(n4368), .ZN(n4443) );
  NAND2_X1 U4839 ( .A1(n4357), .A2(n4443), .ZN(n4142) );
  NAND2_X1 U4840 ( .A1(n4612), .A2(REG2_REG_31__SCAN_IN), .ZN(n4141) );
  OAI211_X1 U4841 ( .C1(n4446), .C2(n4331), .A(n4142), .B(n4141), .ZN(U3260)
         );
  INV_X1 U4842 ( .A(n4143), .ZN(n4157) );
  INV_X1 U4843 ( .A(REG2_REG_29__SCAN_IN), .ZN(n4144) );
  OAI22_X1 U4844 ( .A1(n4146), .A2(n4145), .B1(n4144), .B2(n4357), .ZN(n4147)
         );
  AOI21_X1 U4845 ( .B1(n4149), .B2(n4148), .A(n4147), .ZN(n4156) );
  INV_X1 U4846 ( .A(n4150), .ZN(n4154) );
  OAI22_X1 U4847 ( .A1(n4152), .A2(n4331), .B1(n4151), .B2(n4332), .ZN(n4153)
         );
  OAI21_X1 U4848 ( .B1(n4154), .B2(n4153), .A(n4357), .ZN(n4155) );
  OAI211_X1 U4849 ( .C1(n4157), .C2(n4360), .A(n4156), .B(n4155), .ZN(U3354)
         );
  INV_X1 U4850 ( .A(n4159), .ZN(n4170) );
  AOI22_X1 U4851 ( .A1(n4161), .A2(n4281), .B1(n4160), .B2(n4279), .ZN(n4165)
         );
  INV_X1 U4852 ( .A(n4162), .ZN(n4163) );
  AOI22_X1 U4853 ( .A1(n4163), .A2(n4619), .B1(REG2_REG_28__SCAN_IN), .B2(
        n4627), .ZN(n4164) );
  OAI211_X1 U4854 ( .C1(n4166), .C2(n4285), .A(n4165), .B(n4164), .ZN(n4169)
         );
  NOR2_X1 U4855 ( .A1(n4167), .A2(n4627), .ZN(n4168) );
  OAI21_X1 U4856 ( .B1(n4158), .B2(n4360), .A(n4171), .ZN(U3262) );
  NAND2_X1 U4857 ( .A1(n4172), .A2(n4277), .ZN(n4182) );
  INV_X1 U4858 ( .A(n4173), .ZN(n4180) );
  AOI22_X1 U4859 ( .A1(n4174), .A2(n4279), .B1(n4281), .B2(n4212), .ZN(n4177)
         );
  AOI22_X1 U4860 ( .A1(n4175), .A2(n4619), .B1(REG2_REG_27__SCAN_IN), .B2(
        n4627), .ZN(n4176) );
  OAI211_X1 U4861 ( .C1(n4178), .C2(n4285), .A(n4177), .B(n4176), .ZN(n4179)
         );
  AOI21_X1 U4862 ( .B1(n4180), .B2(n4621), .A(n4179), .ZN(n4181) );
  OAI211_X1 U4863 ( .C1(n4627), .C2(n4183), .A(n4182), .B(n4181), .ZN(U3263)
         );
  XNOR2_X1 U4864 ( .A(n4184), .B(n4188), .ZN(n4371) );
  INV_X1 U4865 ( .A(n4371), .ZN(n4202) );
  INV_X1 U4866 ( .A(n4185), .ZN(n4186) );
  AOI21_X1 U4867 ( .B1(n4204), .B2(n4187), .A(n4186), .ZN(n4190) );
  INV_X1 U4868 ( .A(n4188), .ZN(n4189) );
  XNOR2_X1 U4869 ( .A(n4190), .B(n4189), .ZN(n4191) );
  NAND2_X1 U4870 ( .A1(n4191), .A2(n4348), .ZN(n4194) );
  INV_X1 U4871 ( .A(n4196), .ZN(n4192) );
  AOI22_X1 U4872 ( .A1(n4385), .A2(n4374), .B1(n4192), .B2(n4429), .ZN(n4193)
         );
  OAI211_X1 U4873 ( .C1(n4195), .C2(n4378), .A(n4194), .B(n4193), .ZN(n4370)
         );
  OAI21_X1 U4874 ( .B1(n4209), .B2(n4196), .A(n3016), .ZN(n4453) );
  NOR2_X1 U4875 ( .A1(n4453), .A2(n4331), .ZN(n4200) );
  INV_X1 U4876 ( .A(REG2_REG_26__SCAN_IN), .ZN(n4197) );
  OAI22_X1 U4877 ( .A1(n4198), .A2(n4332), .B1(n4357), .B2(n4197), .ZN(n4199)
         );
  AOI211_X1 U4878 ( .C1(n4370), .C2(n4357), .A(n4200), .B(n4199), .ZN(n4201)
         );
  OAI21_X1 U4879 ( .B1(n4202), .B2(n4360), .A(n4201), .ZN(U3264) );
  NAND2_X1 U4880 ( .A1(n4204), .A2(n4203), .ZN(n4205) );
  XNOR2_X1 U4881 ( .A(n4205), .B(n4208), .ZN(n4206) );
  NAND2_X1 U4882 ( .A1(n4206), .A2(n4348), .ZN(n4377) );
  XOR2_X1 U4883 ( .A(n4208), .B(n4207), .Z(n4381) );
  NAND2_X1 U4884 ( .A1(n4381), .A2(n4277), .ZN(n4220) );
  INV_X1 U4885 ( .A(n4226), .ZN(n4211) );
  INV_X1 U4886 ( .A(n4209), .ZN(n4210) );
  OAI21_X1 U4887 ( .B1(n4211), .B2(n4216), .A(n4210), .ZN(n4457) );
  INV_X1 U4888 ( .A(n4457), .ZN(n4218) );
  AOI22_X1 U4889 ( .A1(n4212), .A2(n4279), .B1(n4281), .B2(n4375), .ZN(n4215)
         );
  AOI22_X1 U4890 ( .A1(n4612), .A2(REG2_REG_25__SCAN_IN), .B1(n4213), .B2(
        n4619), .ZN(n4214) );
  OAI211_X1 U4891 ( .C1(n4216), .C2(n4285), .A(n4215), .B(n4214), .ZN(n4217)
         );
  AOI21_X1 U4892 ( .B1(n4218), .B2(n4621), .A(n4217), .ZN(n4219) );
  OAI211_X1 U4893 ( .C1(n4627), .C2(n4377), .A(n4220), .B(n4219), .ZN(U3265)
         );
  XNOR2_X1 U4894 ( .A(n4222), .B(n4221), .ZN(n4223) );
  NAND2_X1 U4895 ( .A1(n4223), .A2(n4348), .ZN(n4387) );
  XNOR2_X1 U4896 ( .A(n4224), .B(n4225), .ZN(n4390) );
  NAND2_X1 U4897 ( .A1(n4390), .A2(n4277), .ZN(n4235) );
  INV_X1 U4898 ( .A(n4248), .ZN(n4227) );
  OAI21_X1 U4899 ( .B1(n4227), .B2(n4231), .A(n4226), .ZN(n4461) );
  INV_X1 U4900 ( .A(n4461), .ZN(n4233) );
  AOI22_X1 U4901 ( .A1(n4281), .A2(n4261), .B1(n4279), .B2(n4385), .ZN(n4230)
         );
  AOI22_X1 U4902 ( .A1(n4612), .A2(REG2_REG_24__SCAN_IN), .B1(n4228), .B2(
        n4619), .ZN(n4229) );
  OAI211_X1 U4903 ( .C1(n4231), .C2(n4285), .A(n4230), .B(n4229), .ZN(n4232)
         );
  AOI21_X1 U4904 ( .B1(n4233), .B2(n4621), .A(n4232), .ZN(n4234) );
  OAI211_X1 U4905 ( .C1(n4627), .C2(n4387), .A(n4235), .B(n4234), .ZN(U3266)
         );
  XOR2_X1 U4906 ( .A(n4241), .B(n4236), .Z(n4393) );
  INV_X1 U4907 ( .A(n4393), .ZN(n4253) );
  INV_X1 U4908 ( .A(n4237), .ZN(n4238) );
  AOI21_X1 U4909 ( .B1(n4273), .B2(n4276), .A(n4238), .ZN(n4258) );
  OAI21_X1 U4910 ( .B1(n4258), .B2(n4259), .A(n4239), .ZN(n4240) );
  XOR2_X1 U4911 ( .A(n4241), .B(n4240), .Z(n4242) );
  NAND2_X1 U4912 ( .A1(n4242), .A2(n4348), .ZN(n4244) );
  AOI22_X1 U4913 ( .A1(n4401), .A2(n4374), .B1(n4429), .B2(n4246), .ZN(n4243)
         );
  OAI211_X1 U4914 ( .C1(n4245), .C2(n4378), .A(n4244), .B(n4243), .ZN(n4392)
         );
  NAND2_X1 U4915 ( .A1(n4267), .A2(n4246), .ZN(n4247) );
  NAND2_X1 U4916 ( .A1(n4248), .A2(n4247), .ZN(n4465) );
  AOI22_X1 U4917 ( .A1(n4612), .A2(REG2_REG_23__SCAN_IN), .B1(n4249), .B2(
        n4619), .ZN(n4250) );
  OAI21_X1 U4918 ( .B1(n4465), .B2(n4331), .A(n4250), .ZN(n4251) );
  AOI21_X1 U4919 ( .B1(n4392), .B2(n4357), .A(n4251), .ZN(n4252) );
  OAI21_X1 U4920 ( .B1(n4253), .B2(n4360), .A(n4252), .ZN(U3267) );
  AND2_X1 U4921 ( .A1(n4254), .A2(n4259), .ZN(n4255) );
  AOI21_X1 U4922 ( .B1(n4257), .B2(n4256), .A(n4255), .ZN(n4397) );
  INV_X1 U4923 ( .A(n4397), .ZN(n4272) );
  XOR2_X1 U4924 ( .A(n4259), .B(n4258), .Z(n4263) );
  OAI22_X1 U4925 ( .A1(n4300), .A2(n4434), .B1(n4265), .B2(n4323), .ZN(n4260)
         );
  AOI21_X1 U4926 ( .B1(n4431), .B2(n4261), .A(n4260), .ZN(n4262) );
  OAI21_X1 U4927 ( .B1(n4263), .B2(n4326), .A(n4262), .ZN(n4396) );
  OR2_X1 U4928 ( .A1(n4264), .A2(n4265), .ZN(n4266) );
  NAND2_X1 U4929 ( .A1(n4267), .A2(n4266), .ZN(n4468) );
  AOI22_X1 U4930 ( .A1(n4612), .A2(REG2_REG_22__SCAN_IN), .B1(n4268), .B2(
        n4619), .ZN(n4269) );
  OAI21_X1 U4931 ( .B1(n4468), .B2(n4331), .A(n4269), .ZN(n4270) );
  AOI21_X1 U4932 ( .B1(n4396), .B2(n4357), .A(n4270), .ZN(n4271) );
  OAI21_X1 U4933 ( .B1(n4272), .B2(n4360), .A(n4271), .ZN(U3268) );
  XNOR2_X1 U4934 ( .A(n4273), .B(n4276), .ZN(n4274) );
  NAND2_X1 U4935 ( .A1(n4274), .A2(n4348), .ZN(n4403) );
  XNOR2_X1 U4936 ( .A(n4275), .B(n4276), .ZN(n4406) );
  NAND2_X1 U4937 ( .A1(n4406), .A2(n4277), .ZN(n4290) );
  INV_X1 U4938 ( .A(n4264), .ZN(n4278) );
  OAI21_X1 U4939 ( .B1(n4306), .B2(n4286), .A(n4278), .ZN(n4472) );
  INV_X1 U4940 ( .A(n4472), .ZN(n4288) );
  AOI22_X1 U4941 ( .A1(n4281), .A2(n4280), .B1(n4279), .B2(n4401), .ZN(n4284)
         );
  AOI22_X1 U4942 ( .A1(n4612), .A2(REG2_REG_21__SCAN_IN), .B1(n4282), .B2(
        n4619), .ZN(n4283) );
  OAI211_X1 U4943 ( .C1(n4286), .C2(n4285), .A(n4284), .B(n4283), .ZN(n4287)
         );
  AOI21_X1 U4944 ( .B1(n4288), .B2(n4621), .A(n4287), .ZN(n4289) );
  OAI211_X1 U4945 ( .C1(n4627), .C2(n4403), .A(n4290), .B(n4289), .ZN(U3269)
         );
  XNOR2_X1 U4946 ( .A(n4291), .B(n4292), .ZN(n4305) );
  INV_X1 U4947 ( .A(n4293), .ZN(n4295) );
  OAI21_X1 U4948 ( .B1(n4317), .B2(n4295), .A(n4294), .ZN(n4297) );
  XNOR2_X1 U4949 ( .A(n4297), .B(n4296), .ZN(n4302) );
  AOI22_X1 U4950 ( .A1(n4344), .A2(n4374), .B1(n4298), .B2(n4429), .ZN(n4299)
         );
  OAI21_X1 U4951 ( .B1(n4300), .B2(n4378), .A(n4299), .ZN(n4301) );
  AOI21_X1 U4952 ( .B1(n4302), .B2(n4348), .A(n4301), .ZN(n4303) );
  OAI21_X1 U4953 ( .B1(n4305), .B2(n4304), .A(n4303), .ZN(n4409) );
  INV_X1 U4954 ( .A(n4409), .ZN(n4314) );
  INV_X1 U4955 ( .A(n4305), .ZN(n4410) );
  INV_X1 U4956 ( .A(n4328), .ZN(n4309) );
  INV_X1 U4957 ( .A(n4306), .ZN(n4307) );
  OAI21_X1 U4958 ( .B1(n4309), .B2(n4308), .A(n4307), .ZN(n4476) );
  AOI22_X1 U4959 ( .A1(n4612), .A2(REG2_REG_20__SCAN_IN), .B1(n4310), .B2(
        n4619), .ZN(n4311) );
  OAI21_X1 U4960 ( .B1(n4476), .B2(n4331), .A(n4311), .ZN(n4312) );
  AOI21_X1 U4961 ( .B1(n4410), .B2(n4622), .A(n4312), .ZN(n4313) );
  OAI21_X1 U4962 ( .B1(n4314), .B2(n4627), .A(n4313), .ZN(U3270) );
  XNOR2_X1 U4963 ( .A(n4315), .B(n4322), .ZN(n4414) );
  INV_X1 U4964 ( .A(n4414), .ZN(n4337) );
  NAND2_X1 U4965 ( .A1(n4317), .A2(n4316), .ZN(n4341) );
  INV_X1 U4966 ( .A(n4318), .ZN(n4320) );
  OAI21_X1 U4967 ( .B1(n4341), .B2(n4320), .A(n4319), .ZN(n4321) );
  XOR2_X1 U4968 ( .A(n4322), .B(n4321), .Z(n4327) );
  OAI22_X1 U4969 ( .A1(n4404), .A2(n4378), .B1(n4323), .B2(n4329), .ZN(n4324)
         );
  AOI21_X1 U4970 ( .B1(n4374), .B2(n4421), .A(n4324), .ZN(n4325) );
  OAI21_X1 U4971 ( .B1(n4327), .B2(n4326), .A(n4325), .ZN(n4413) );
  INV_X1 U4972 ( .A(n4350), .ZN(n4330) );
  OAI21_X1 U4973 ( .B1(n4330), .B2(n4329), .A(n4328), .ZN(n4480) );
  NOR2_X1 U4974 ( .A1(n4480), .A2(n4331), .ZN(n4335) );
  OAI22_X1 U4975 ( .A1(n4357), .A2(n4083), .B1(n4333), .B2(n4332), .ZN(n4334)
         );
  AOI211_X1 U4976 ( .C1(n4413), .C2(n4357), .A(n4335), .B(n4334), .ZN(n4336)
         );
  OAI21_X1 U4977 ( .B1(n4337), .B2(n4360), .A(n4336), .ZN(U3271) );
  OAI21_X1 U4978 ( .B1(n4339), .B2(n4342), .A(n4338), .ZN(n4340) );
  INV_X1 U4979 ( .A(n4340), .ZN(n4419) );
  XOR2_X1 U4980 ( .A(n4342), .B(n4341), .Z(n4349) );
  AOI22_X1 U4981 ( .A1(n4344), .A2(n4431), .B1(n4343), .B2(n4429), .ZN(n4345)
         );
  OAI21_X1 U4982 ( .B1(n4346), .B2(n4434), .A(n4345), .ZN(n4347) );
  AOI21_X1 U4983 ( .B1(n4349), .B2(n4348), .A(n4347), .ZN(n4418) );
  INV_X1 U4984 ( .A(n4418), .ZN(n4358) );
  OAI211_X1 U4985 ( .C1(n4352), .C2(n4351), .A(n4437), .B(n4350), .ZN(n4417)
         );
  AOI22_X1 U4986 ( .A1(n4612), .A2(REG2_REG_18__SCAN_IN), .B1(n4353), .B2(
        n4619), .ZN(n4354) );
  OAI21_X1 U4987 ( .B1(n4417), .B2(n4355), .A(n4354), .ZN(n4356) );
  AOI21_X1 U4988 ( .B1(n4358), .B2(n4357), .A(n4356), .ZN(n4359) );
  OAI21_X1 U4989 ( .B1(n4419), .B2(n4360), .A(n4359), .ZN(U3272) );
  NOR2_X1 U4990 ( .A1(n4682), .A2(n4361), .ZN(n4362) );
  AOI21_X1 U4991 ( .B1(n4682), .B2(n4443), .A(n4362), .ZN(n4363) );
  OAI21_X1 U4992 ( .B1(n4446), .B2(n4428), .A(n4363), .ZN(U3549) );
  AOI21_X1 U4993 ( .B1(n4366), .B2(n4365), .A(n4364), .ZN(n4497) );
  INV_X1 U4994 ( .A(n4497), .ZN(n4449) );
  NAND2_X1 U4995 ( .A1(n4429), .A2(n4366), .ZN(n4367) );
  AND2_X1 U4996 ( .A1(n4368), .A2(n4367), .ZN(n4499) );
  MUX2_X1 U4997 ( .A(n4499), .B(n3037), .S(n4680), .Z(n4369) );
  OAI21_X1 U4998 ( .B1(n4449), .B2(n4428), .A(n4369), .ZN(U3548) );
  AOI21_X1 U4999 ( .B1(n4371), .B2(n4667), .A(n4370), .ZN(n4450) );
  MUX2_X1 U5000 ( .A(n4798), .B(n4450), .S(n4682), .Z(n4372) );
  OAI21_X1 U5001 ( .B1(n4428), .B2(n4453), .A(n4372), .ZN(U3544) );
  AOI22_X1 U5002 ( .A1(n4375), .A2(n4374), .B1(n4373), .B2(n4429), .ZN(n4376)
         );
  OAI211_X1 U5003 ( .C1(n4379), .C2(n4378), .A(n4377), .B(n4376), .ZN(n4380)
         );
  AOI21_X1 U5004 ( .B1(n4381), .B2(n4667), .A(n4380), .ZN(n4454) );
  MUX2_X1 U5005 ( .A(n4382), .B(n4454), .S(n4682), .Z(n4383) );
  OAI21_X1 U5006 ( .B1(n4428), .B2(n4457), .A(n4383), .ZN(U3543) );
  AOI22_X1 U5007 ( .A1(n4385), .A2(n4431), .B1(n4429), .B2(n4384), .ZN(n4386)
         );
  OAI211_X1 U5008 ( .C1(n4388), .C2(n4434), .A(n4387), .B(n4386), .ZN(n4389)
         );
  AOI21_X1 U5009 ( .B1(n4390), .B2(n4667), .A(n4389), .ZN(n4458) );
  MUX2_X1 U5010 ( .A(n4949), .B(n4458), .S(n4682), .Z(n4391) );
  OAI21_X1 U5011 ( .B1(n4428), .B2(n4461), .A(n4391), .ZN(U3542) );
  AOI21_X1 U5012 ( .B1(n4393), .B2(n4667), .A(n4392), .ZN(n4462) );
  MUX2_X1 U5013 ( .A(n4394), .B(n4462), .S(n4682), .Z(n4395) );
  OAI21_X1 U5014 ( .B1(n4428), .B2(n4465), .A(n4395), .ZN(U3541) );
  INV_X1 U5015 ( .A(REG1_REG_22__SCAN_IN), .ZN(n4398) );
  AOI21_X1 U5016 ( .B1(n4397), .B2(n4667), .A(n4396), .ZN(n4466) );
  MUX2_X1 U5017 ( .A(n4398), .B(n4466), .S(n4682), .Z(n4399) );
  OAI21_X1 U5018 ( .B1(n4428), .B2(n4468), .A(n4399), .ZN(U3540) );
  INV_X1 U5019 ( .A(REG1_REG_21__SCAN_IN), .ZN(n4407) );
  AOI22_X1 U5020 ( .A1(n4401), .A2(n4431), .B1(n4429), .B2(n4400), .ZN(n4402)
         );
  OAI211_X1 U5021 ( .C1(n4404), .C2(n4434), .A(n4403), .B(n4402), .ZN(n4405)
         );
  AOI21_X1 U5022 ( .B1(n4406), .B2(n4667), .A(n4405), .ZN(n4469) );
  MUX2_X1 U5023 ( .A(n4407), .B(n4469), .S(n4682), .Z(n4408) );
  OAI21_X1 U5024 ( .B1(n4428), .B2(n4472), .A(n4408), .ZN(U3539) );
  AOI21_X1 U5025 ( .B1(n4664), .B2(n4410), .A(n4409), .ZN(n4473) );
  MUX2_X1 U5026 ( .A(n4411), .B(n4473), .S(n4682), .Z(n4412) );
  OAI21_X1 U5027 ( .B1(n4428), .B2(n4476), .A(n4412), .ZN(U3538) );
  AOI21_X1 U5028 ( .B1(n4414), .B2(n4667), .A(n4413), .ZN(n4477) );
  MUX2_X1 U5029 ( .A(n4415), .B(n4477), .S(n4682), .Z(n4416) );
  OAI21_X1 U5030 ( .B1(n4428), .B2(n4480), .A(n4416), .ZN(U3537) );
  OAI211_X1 U5031 ( .C1(n4419), .C2(n4441), .A(n4418), .B(n4417), .ZN(n4481)
         );
  MUX2_X1 U5032 ( .A(REG1_REG_18__SCAN_IN), .B(n4481), .S(n4682), .Z(U3536) );
  AOI22_X1 U5033 ( .A1(n4421), .A2(n4431), .B1(n4429), .B2(n4420), .ZN(n4422)
         );
  OAI211_X1 U5034 ( .C1(n4424), .C2(n4434), .A(n4423), .B(n4422), .ZN(n4425)
         );
  AOI21_X1 U5035 ( .B1(n4426), .B2(n4667), .A(n4425), .ZN(n4482) );
  MUX2_X1 U5036 ( .A(n4127), .B(n4482), .S(n4682), .Z(n4427) );
  OAI21_X1 U5037 ( .B1(n4428), .B2(n4486), .A(n4427), .ZN(U3535) );
  AOI22_X1 U5038 ( .A1(n4432), .A2(n4431), .B1(n4430), .B2(n4429), .ZN(n4433)
         );
  OAI21_X1 U5039 ( .B1(n4435), .B2(n4434), .A(n4433), .ZN(n4436) );
  AOI21_X1 U5040 ( .B1(n4438), .B2(n4437), .A(n4436), .ZN(n4440) );
  OAI211_X1 U5041 ( .C1(n4442), .C2(n4441), .A(n4440), .B(n4439), .ZN(n4487)
         );
  MUX2_X1 U5042 ( .A(REG1_REG_16__SCAN_IN), .B(n4487), .S(n4682), .Z(U3534) );
  NAND2_X1 U5043 ( .A1(n4675), .A2(n4443), .ZN(n4445) );
  NAND2_X1 U5044 ( .A1(n4673), .A2(REG0_REG_31__SCAN_IN), .ZN(n4444) );
  OAI211_X1 U5045 ( .C1(n4446), .C2(n4485), .A(n4445), .B(n4444), .ZN(U3517)
         );
  INV_X1 U5046 ( .A(REG0_REG_30__SCAN_IN), .ZN(n4447) );
  MUX2_X1 U5047 ( .A(n4499), .B(n4447), .S(n4673), .Z(n4448) );
  OAI21_X1 U5048 ( .B1(n4449), .B2(n4485), .A(n4448), .ZN(U3516) );
  INV_X1 U5049 ( .A(REG0_REG_26__SCAN_IN), .ZN(n4451) );
  MUX2_X1 U5050 ( .A(n4451), .B(n4450), .S(n4675), .Z(n4452) );
  OAI21_X1 U5051 ( .B1(n4453), .B2(n4485), .A(n4452), .ZN(U3512) );
  INV_X1 U5052 ( .A(REG0_REG_25__SCAN_IN), .ZN(n4455) );
  MUX2_X1 U5053 ( .A(n4455), .B(n4454), .S(n4675), .Z(n4456) );
  OAI21_X1 U5054 ( .B1(n4457), .B2(n4485), .A(n4456), .ZN(U3511) );
  INV_X1 U5055 ( .A(REG0_REG_24__SCAN_IN), .ZN(n4459) );
  MUX2_X1 U5056 ( .A(n4459), .B(n4458), .S(n4675), .Z(n4460) );
  OAI21_X1 U5057 ( .B1(n4461), .B2(n4485), .A(n4460), .ZN(U3510) );
  INV_X1 U5058 ( .A(REG0_REG_23__SCAN_IN), .ZN(n4463) );
  MUX2_X1 U5059 ( .A(n4463), .B(n4462), .S(n4675), .Z(n4464) );
  OAI21_X1 U5060 ( .B1(n4465), .B2(n4485), .A(n4464), .ZN(U3509) );
  INV_X1 U5061 ( .A(REG0_REG_22__SCAN_IN), .ZN(n4932) );
  MUX2_X1 U5062 ( .A(n4932), .B(n4466), .S(n4675), .Z(n4467) );
  OAI21_X1 U5063 ( .B1(n4468), .B2(n4485), .A(n4467), .ZN(U3508) );
  INV_X1 U5064 ( .A(REG0_REG_21__SCAN_IN), .ZN(n4470) );
  MUX2_X1 U5065 ( .A(n4470), .B(n4469), .S(n4675), .Z(n4471) );
  OAI21_X1 U5066 ( .B1(n4472), .B2(n4485), .A(n4471), .ZN(U3507) );
  INV_X1 U5067 ( .A(REG0_REG_20__SCAN_IN), .ZN(n4474) );
  MUX2_X1 U5068 ( .A(n4474), .B(n4473), .S(n4675), .Z(n4475) );
  OAI21_X1 U5069 ( .B1(n4476), .B2(n4485), .A(n4475), .ZN(U3506) );
  INV_X1 U5070 ( .A(REG0_REG_19__SCAN_IN), .ZN(n4478) );
  MUX2_X1 U5071 ( .A(n4478), .B(n4477), .S(n4675), .Z(n4479) );
  OAI21_X1 U5072 ( .B1(n4480), .B2(n4485), .A(n4479), .ZN(U3505) );
  MUX2_X1 U5073 ( .A(REG0_REG_18__SCAN_IN), .B(n4481), .S(n4675), .Z(U3503) );
  INV_X1 U5074 ( .A(REG0_REG_17__SCAN_IN), .ZN(n4483) );
  MUX2_X1 U5075 ( .A(n4483), .B(n4482), .S(n4675), .Z(n4484) );
  OAI21_X1 U5076 ( .B1(n4486), .B2(n4485), .A(n4484), .ZN(U3501) );
  MUX2_X1 U5077 ( .A(REG0_REG_16__SCAN_IN), .B(n4487), .S(n4675), .Z(U3499) );
  MUX2_X1 U5078 ( .A(DATAI_28_), .B(n4488), .S(STATE_REG_SCAN_IN), .Z(U3324)
         );
  MUX2_X1 U5079 ( .A(n4489), .B(DATAI_21_), .S(U3149), .Z(U3331) );
  MUX2_X1 U5080 ( .A(n4490), .B(DATAI_19_), .S(U3149), .Z(U3333) );
  MUX2_X1 U5081 ( .A(n4491), .B(DATAI_8_), .S(U3149), .Z(U3344) );
  MUX2_X1 U5082 ( .A(n4492), .B(DATAI_7_), .S(U3149), .Z(U3345) );
  MUX2_X1 U5083 ( .A(n4493), .B(DATAI_6_), .S(U3149), .Z(U3346) );
  MUX2_X1 U5084 ( .A(DATAI_4_), .B(n4494), .S(STATE_REG_SCAN_IN), .Z(U3348) );
  MUX2_X1 U5085 ( .A(n4495), .B(DATAI_3_), .S(U3149), .Z(U3349) );
  MUX2_X1 U5086 ( .A(n4496), .B(DATAI_2_), .S(U3149), .Z(U3350) );
  MUX2_X1 U5087 ( .A(n3116), .B(DATAI_1_), .S(U3149), .Z(U3351) );
  AOI22_X1 U5088 ( .A1(n4497), .A2(n4621), .B1(REG2_REG_30__SCAN_IN), .B2(
        n4627), .ZN(n4498) );
  OAI21_X1 U5089 ( .B1(n4627), .B2(n4499), .A(n4498), .ZN(U3261) );
  INV_X1 U5090 ( .A(n4502), .ZN(n4500) );
  OAI211_X1 U5091 ( .C1(REG1_REG_0__SCAN_IN), .C2(n4501), .A(n4503), .B(n4500), 
        .ZN(n4506) );
  AOI22_X1 U5092 ( .A1(n4503), .A2(n4502), .B1(n4606), .B2(n4676), .ZN(n4505)
         );
  AOI22_X1 U5093 ( .A1(ADDR_REG_0__SCAN_IN), .A2(n4604), .B1(
        REG3_REG_0__SCAN_IN), .B2(U3149), .ZN(n4504) );
  OAI221_X1 U5094 ( .B1(IR_REG_0__SCAN_IN), .B2(n4506), .C1(n2309), .C2(n4505), 
        .A(n4504), .ZN(U3240) );
  OAI211_X1 U5095 ( .C1(n4509), .C2(n4508), .A(n4606), .B(n4507), .ZN(n4514)
         );
  OAI211_X1 U5096 ( .C1(n4512), .C2(n4511), .A(n4549), .B(n4510), .ZN(n4513)
         );
  OAI211_X1 U5097 ( .C1(n4610), .C2(n4646), .A(n4514), .B(n4513), .ZN(n4515)
         );
  AOI211_X1 U5098 ( .C1(n4604), .C2(ADDR_REG_9__SCAN_IN), .A(n4516), .B(n4515), 
        .ZN(n4517) );
  INV_X1 U5099 ( .A(n4517), .ZN(U3249) );
  OAI211_X1 U5100 ( .C1(REG1_REG_10__SCAN_IN), .C2(n4519), .A(n4606), .B(n4518), .ZN(n4523) );
  OAI211_X1 U5101 ( .C1(REG2_REG_10__SCAN_IN), .C2(n4521), .A(n4549), .B(n4520), .ZN(n4522) );
  OAI211_X1 U5102 ( .C1(n4610), .C2(n4644), .A(n4523), .B(n4522), .ZN(n4524)
         );
  AOI211_X1 U5103 ( .C1(n4604), .C2(ADDR_REG_10__SCAN_IN), .A(n4525), .B(n4524), .ZN(n4526) );
  INV_X1 U5104 ( .A(n4526), .ZN(U3250) );
  OAI211_X1 U5105 ( .C1(n4529), .C2(n4528), .A(n4606), .B(n4527), .ZN(n4534)
         );
  OAI211_X1 U5106 ( .C1(n4532), .C2(n4531), .A(n4549), .B(n4530), .ZN(n4533)
         );
  OAI211_X1 U5107 ( .C1(n4610), .C2(n4643), .A(n4534), .B(n4533), .ZN(n4535)
         );
  AOI211_X1 U5108 ( .C1(n4604), .C2(ADDR_REG_11__SCAN_IN), .A(n4536), .B(n4535), .ZN(n4537) );
  INV_X1 U5109 ( .A(n4537), .ZN(U3251) );
  OAI211_X1 U5110 ( .C1(REG2_REG_12__SCAN_IN), .C2(n4539), .A(n4549), .B(n4538), .ZN(n4541) );
  NAND2_X1 U5111 ( .A1(n4541), .A2(n4540), .ZN(n4542) );
  AOI21_X1 U5112 ( .B1(n4604), .B2(ADDR_REG_12__SCAN_IN), .A(n4542), .ZN(n4546) );
  OAI211_X1 U5113 ( .C1(REG1_REG_12__SCAN_IN), .C2(n4544), .A(n4606), .B(n4543), .ZN(n4545) );
  OAI211_X1 U5114 ( .C1(n4610), .C2(n4641), .A(n4546), .B(n4545), .ZN(U3252)
         );
  AOI22_X1 U5115 ( .A1(REG2_REG_13__SCAN_IN), .A2(n4548), .B1(n4640), .B2(
        n4547), .ZN(n4552) );
  OAI21_X1 U5116 ( .B1(n4552), .B2(n4551), .A(n4549), .ZN(n4550) );
  AOI21_X1 U5117 ( .B1(n4552), .B2(n4551), .A(n4550), .ZN(n4554) );
  AOI211_X1 U5118 ( .C1(n4604), .C2(ADDR_REG_13__SCAN_IN), .A(n4554), .B(n4553), .ZN(n4559) );
  OAI211_X1 U5119 ( .C1(n4557), .C2(n4556), .A(n4606), .B(n4555), .ZN(n4558)
         );
  OAI211_X1 U5120 ( .C1(n4610), .C2(n4640), .A(n4559), .B(n4558), .ZN(U3253)
         );
  INV_X1 U5121 ( .A(n4560), .ZN(n4564) );
  AOI211_X1 U5122 ( .C1(n4810), .C2(n4562), .A(n4561), .B(n4600), .ZN(n4563)
         );
  AOI211_X1 U5123 ( .C1(n4604), .C2(ADDR_REG_14__SCAN_IN), .A(n4564), .B(n4563), .ZN(n4568) );
  OAI211_X1 U5124 ( .C1(REG1_REG_14__SCAN_IN), .C2(n4566), .A(n4606), .B(n4565), .ZN(n4567) );
  OAI211_X1 U5125 ( .C1(n4610), .C2(n4569), .A(n4568), .B(n4567), .ZN(U3254)
         );
  AOI211_X1 U5126 ( .C1(n4572), .C2(n4571), .A(n4570), .B(n4600), .ZN(n4573)
         );
  AOI211_X1 U5127 ( .C1(n4604), .C2(ADDR_REG_15__SCAN_IN), .A(n4574), .B(n4573), .ZN(n4579) );
  OAI211_X1 U5128 ( .C1(n4577), .C2(n4576), .A(n4606), .B(n4575), .ZN(n4578)
         );
  OAI211_X1 U5129 ( .C1(n4610), .C2(n4637), .A(n4579), .B(n4578), .ZN(U3255)
         );
  INV_X1 U5130 ( .A(n4580), .ZN(n4584) );
  AOI221_X1 U5131 ( .B1(n4582), .B2(n4581), .C1(n4952), .C2(n4581), .A(n4600), 
        .ZN(n4583) );
  AOI211_X1 U5132 ( .C1(n4604), .C2(ADDR_REG_16__SCAN_IN), .A(n4584), .B(n4583), .ZN(n4588) );
  OAI221_X1 U5133 ( .B1(n4586), .B2(REG1_REG_16__SCAN_IN), .C1(n4586), .C2(
        n4585), .A(n4606), .ZN(n4587) );
  OAI211_X1 U5134 ( .C1(n4610), .C2(n4636), .A(n4588), .B(n4587), .ZN(U3256)
         );
  AOI221_X1 U5135 ( .B1(n4591), .B2(n4590), .C1(n4589), .C2(n4590), .A(n4600), 
        .ZN(n4592) );
  AOI211_X1 U5136 ( .C1(n4604), .C2(ADDR_REG_17__SCAN_IN), .A(n4593), .B(n4592), .ZN(n4598) );
  OAI221_X1 U5137 ( .B1(n4596), .B2(n4595), .C1(n4596), .C2(n4594), .A(n4606), 
        .ZN(n4597) );
  OAI211_X1 U5138 ( .C1(n4610), .C2(n4599), .A(n4598), .B(n4597), .ZN(U3257)
         );
  OAI211_X1 U5139 ( .C1(n4607), .C2(n2164), .A(n4606), .B(n4605), .ZN(n4608)
         );
  OAI211_X1 U5140 ( .C1(n4610), .C2(n4632), .A(n4609), .B(n4608), .ZN(U3258)
         );
  AOI22_X1 U5141 ( .A1(n4612), .A2(REG2_REG_8__SCAN_IN), .B1(n4611), .B2(n4619), .ZN(n4617) );
  INV_X1 U5142 ( .A(n4613), .ZN(n4614) );
  AOI22_X1 U5143 ( .A1(n4615), .A2(n4622), .B1(n4621), .B2(n4614), .ZN(n4616)
         );
  OAI211_X1 U5144 ( .C1(n4627), .C2(n4618), .A(n4617), .B(n4616), .ZN(U3282)
         );
  AOI22_X1 U5145 ( .A1(REG3_REG_2__SCAN_IN), .A2(n4619), .B1(
        REG2_REG_2__SCAN_IN), .B2(n4627), .ZN(n4625) );
  AOI22_X1 U5146 ( .A1(n4623), .A2(n4622), .B1(n4621), .B2(n4620), .ZN(n4624)
         );
  OAI211_X1 U5147 ( .C1(n4627), .C2(n4626), .A(n4625), .B(n4624), .ZN(U3288)
         );
  AND2_X1 U5148 ( .A1(D_REG_31__SCAN_IN), .A2(n4628), .ZN(U3291) );
  AND2_X1 U5149 ( .A1(D_REG_30__SCAN_IN), .A2(n4628), .ZN(U3292) );
  AND2_X1 U5150 ( .A1(D_REG_29__SCAN_IN), .A2(n4628), .ZN(U3293) );
  INV_X1 U5151 ( .A(D_REG_28__SCAN_IN), .ZN(n4758) );
  NOR2_X1 U5152 ( .A1(n4629), .A2(n4758), .ZN(U3294) );
  INV_X1 U5153 ( .A(D_REG_27__SCAN_IN), .ZN(n4757) );
  NOR2_X1 U5154 ( .A1(n4629), .A2(n4757), .ZN(U3295) );
  AND2_X1 U5155 ( .A1(D_REG_26__SCAN_IN), .A2(n4628), .ZN(U3296) );
  AND2_X1 U5156 ( .A1(D_REG_25__SCAN_IN), .A2(n4628), .ZN(U3297) );
  INV_X1 U5157 ( .A(D_REG_24__SCAN_IN), .ZN(n4755) );
  NOR2_X1 U5158 ( .A1(n4629), .A2(n4755), .ZN(U3298) );
  AND2_X1 U5159 ( .A1(D_REG_23__SCAN_IN), .A2(n4628), .ZN(U3299) );
  INV_X1 U5160 ( .A(D_REG_22__SCAN_IN), .ZN(n4948) );
  NOR2_X1 U5161 ( .A1(n4629), .A2(n4948), .ZN(U3300) );
  NOR2_X1 U5162 ( .A1(n4629), .A2(n4753), .ZN(U3301) );
  INV_X1 U5163 ( .A(D_REG_20__SCAN_IN), .ZN(n4752) );
  NOR2_X1 U5164 ( .A1(n4629), .A2(n4752), .ZN(U3302) );
  AND2_X1 U5165 ( .A1(D_REG_19__SCAN_IN), .A2(n4628), .ZN(U3303) );
  INV_X1 U5166 ( .A(D_REG_18__SCAN_IN), .ZN(n4750) );
  NOR2_X1 U5167 ( .A1(n4629), .A2(n4750), .ZN(U3304) );
  NOR2_X1 U5168 ( .A1(n4629), .A2(n4749), .ZN(U3305) );
  INV_X1 U5169 ( .A(D_REG_16__SCAN_IN), .ZN(n4742) );
  NOR2_X1 U5170 ( .A1(n4629), .A2(n4742), .ZN(U3306) );
  AND2_X1 U5171 ( .A1(D_REG_15__SCAN_IN), .A2(n4628), .ZN(U3307) );
  AND2_X1 U5172 ( .A1(D_REG_14__SCAN_IN), .A2(n4628), .ZN(U3308) );
  AND2_X1 U5173 ( .A1(D_REG_13__SCAN_IN), .A2(n4628), .ZN(U3309) );
  AND2_X1 U5174 ( .A1(D_REG_12__SCAN_IN), .A2(n4628), .ZN(U3310) );
  AND2_X1 U5175 ( .A1(D_REG_11__SCAN_IN), .A2(n4628), .ZN(U3311) );
  INV_X1 U5176 ( .A(D_REG_10__SCAN_IN), .ZN(n4743) );
  NOR2_X1 U5177 ( .A1(n4629), .A2(n4743), .ZN(U3312) );
  INV_X1 U5178 ( .A(D_REG_9__SCAN_IN), .ZN(n4876) );
  NOR2_X1 U5179 ( .A1(n4629), .A2(n4876), .ZN(U3313) );
  AND2_X1 U5180 ( .A1(D_REG_8__SCAN_IN), .A2(n4628), .ZN(U3314) );
  INV_X1 U5181 ( .A(D_REG_7__SCAN_IN), .ZN(n4740) );
  NOR2_X1 U5182 ( .A1(n4629), .A2(n4740), .ZN(U3315) );
  INV_X1 U5183 ( .A(D_REG_6__SCAN_IN), .ZN(n4739) );
  NOR2_X1 U5184 ( .A1(n4629), .A2(n4739), .ZN(U3316) );
  INV_X1 U5185 ( .A(D_REG_5__SCAN_IN), .ZN(n4736) );
  NOR2_X1 U5186 ( .A1(n4629), .A2(n4736), .ZN(U3317) );
  AND2_X1 U5187 ( .A1(D_REG_4__SCAN_IN), .A2(n4628), .ZN(U3318) );
  INV_X1 U5188 ( .A(D_REG_3__SCAN_IN), .ZN(n4737) );
  NOR2_X1 U5189 ( .A1(n4629), .A2(n4737), .ZN(U3319) );
  INV_X1 U5190 ( .A(D_REG_2__SCAN_IN), .ZN(n4734) );
  NOR2_X1 U5191 ( .A1(n4629), .A2(n4734), .ZN(U3320) );
  OAI21_X1 U5192 ( .B1(STATE_REG_SCAN_IN), .B2(DATAI_23_), .A(n4630), .ZN(
        n4631) );
  INV_X1 U5193 ( .A(n4631), .ZN(U3329) );
  AOI22_X1 U5194 ( .A1(STATE_REG_SCAN_IN), .A2(n4632), .B1(n2706), .B2(U3149), 
        .ZN(U3334) );
  OAI22_X1 U5195 ( .A1(U3149), .A2(n4633), .B1(DATAI_17_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4634) );
  INV_X1 U5196 ( .A(n4634), .ZN(U3335) );
  INV_X1 U5197 ( .A(DATAI_16_), .ZN(n4635) );
  AOI22_X1 U5198 ( .A1(STATE_REG_SCAN_IN), .A2(n4636), .B1(n4635), .B2(U3149), 
        .ZN(U3336) );
  INV_X1 U5199 ( .A(DATAI_15_), .ZN(n4698) );
  AOI22_X1 U5200 ( .A1(STATE_REG_SCAN_IN), .A2(n4637), .B1(n4698), .B2(U3149), 
        .ZN(U3337) );
  OAI22_X1 U5201 ( .A1(U3149), .A2(n4638), .B1(DATAI_14_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4639) );
  INV_X1 U5202 ( .A(n4639), .ZN(U3338) );
  AOI22_X1 U5203 ( .A1(STATE_REG_SCAN_IN), .A2(n4640), .B1(n4697), .B2(U3149), 
        .ZN(U3339) );
  AOI22_X1 U5204 ( .A1(STATE_REG_SCAN_IN), .A2(n4641), .B1(n2599), .B2(U3149), 
        .ZN(U3340) );
  AOI22_X1 U5205 ( .A1(STATE_REG_SCAN_IN), .A2(n4643), .B1(n4642), .B2(U3149), 
        .ZN(U3341) );
  INV_X1 U5206 ( .A(DATAI_10_), .ZN(n4900) );
  AOI22_X1 U5207 ( .A1(STATE_REG_SCAN_IN), .A2(n4644), .B1(n4900), .B2(U3149), 
        .ZN(U3342) );
  INV_X1 U5208 ( .A(DATAI_9_), .ZN(n4645) );
  AOI22_X1 U5209 ( .A1(STATE_REG_SCAN_IN), .A2(n4646), .B1(n4645), .B2(U3149), 
        .ZN(U3343) );
  INV_X1 U5210 ( .A(DATAI_0_), .ZN(n4704) );
  AOI22_X1 U5211 ( .A1(STATE_REG_SCAN_IN), .A2(n2309), .B1(n4704), .B2(U3149), 
        .ZN(U3352) );
  INV_X1 U5212 ( .A(n4647), .ZN(n4650) );
  INV_X1 U5213 ( .A(n4648), .ZN(n4649) );
  AOI211_X1 U5214 ( .C1(n4664), .C2(n4651), .A(n4650), .B(n4649), .ZN(n4677)
         );
  INV_X1 U5215 ( .A(REG0_REG_0__SCAN_IN), .ZN(n4652) );
  AOI22_X1 U5216 ( .A1(n4675), .A2(n4677), .B1(n4652), .B2(n4673), .ZN(U3467)
         );
  OAI22_X1 U5217 ( .A1(n4656), .A2(n4655), .B1(n4654), .B2(n4653), .ZN(n4657)
         );
  NOR2_X1 U5218 ( .A1(n4658), .A2(n4657), .ZN(n4678) );
  INV_X1 U5219 ( .A(REG0_REG_1__SCAN_IN), .ZN(n4659) );
  AOI22_X1 U5220 ( .A1(n4675), .A2(n4678), .B1(n4659), .B2(n4673), .ZN(U3469)
         );
  INV_X1 U5221 ( .A(n4660), .ZN(n4665) );
  INV_X1 U5222 ( .A(n4661), .ZN(n4663) );
  AOI211_X1 U5223 ( .C1(n4665), .C2(n4664), .A(n4663), .B(n4662), .ZN(n4679)
         );
  INV_X1 U5224 ( .A(REG0_REG_4__SCAN_IN), .ZN(n4666) );
  AOI22_X1 U5225 ( .A1(n4675), .A2(n4679), .B1(n4666), .B2(n4673), .ZN(U3475)
         );
  NAND3_X1 U5226 ( .A1(n4669), .A2(n4668), .A3(n4667), .ZN(n4670) );
  AND3_X1 U5227 ( .A1(n4672), .A2(n4671), .A3(n4670), .ZN(n4681) );
  INV_X1 U5228 ( .A(REG0_REG_7__SCAN_IN), .ZN(n4674) );
  AOI22_X1 U5229 ( .A1(n4675), .A2(n4681), .B1(n4674), .B2(n4673), .ZN(U3481)
         );
  AOI22_X1 U5230 ( .A1(n4682), .A2(n4677), .B1(n4676), .B2(n4680), .ZN(U3518)
         );
  AOI22_X1 U5231 ( .A1(n4682), .A2(n4678), .B1(n2353), .B2(n4680), .ZN(U3519)
         );
  AOI22_X1 U5232 ( .A1(n4682), .A2(n4679), .B1(n2447), .B2(n4680), .ZN(U3522)
         );
  AOI22_X1 U5233 ( .A1(n4682), .A2(n4681), .B1(n2508), .B2(n4680), .ZN(U3525)
         );
  AOI22_X1 U5234 ( .A1(n4902), .A2(keyinput32), .B1(n4684), .B2(keyinput61), 
        .ZN(n4683) );
  OAI221_X1 U5235 ( .B1(n4902), .B2(keyinput32), .C1(n4684), .C2(keyinput61), 
        .A(n4683), .ZN(n4695) );
  AOI22_X1 U5236 ( .A1(n4903), .A2(keyinput45), .B1(n4686), .B2(keyinput2), 
        .ZN(n4685) );
  OAI221_X1 U5237 ( .B1(n4903), .B2(keyinput45), .C1(n4686), .C2(keyinput2), 
        .A(n4685), .ZN(n4694) );
  INV_X1 U5238 ( .A(DATAI_21_), .ZN(n4688) );
  AOI22_X1 U5239 ( .A1(n4689), .A2(keyinput7), .B1(keyinput115), .B2(n4688), 
        .ZN(n4687) );
  OAI221_X1 U5240 ( .B1(n4689), .B2(keyinput7), .C1(n4688), .C2(keyinput115), 
        .A(n4687), .ZN(n4693) );
  INV_X1 U5241 ( .A(DATAI_19_), .ZN(n4691) );
  AOI22_X1 U5242 ( .A1(n4691), .A2(keyinput123), .B1(n4901), .B2(keyinput97), 
        .ZN(n4690) );
  OAI221_X1 U5243 ( .B1(n4691), .B2(keyinput123), .C1(n4901), .C2(keyinput97), 
        .A(n4690), .ZN(n4692) );
  NOR4_X1 U5244 ( .A1(n4695), .A2(n4694), .A3(n4693), .A4(n4692), .ZN(n4731)
         );
  AOI22_X1 U5245 ( .A1(n4698), .A2(keyinput50), .B1(keyinput96), .B2(n4697), 
        .ZN(n4696) );
  OAI221_X1 U5246 ( .B1(n4698), .B2(keyinput50), .C1(n4697), .C2(keyinput96), 
        .A(n4696), .ZN(n4708) );
  AOI22_X1 U5247 ( .A1(n2599), .A2(keyinput15), .B1(keyinput64), .B2(n4900), 
        .ZN(n4699) );
  OAI221_X1 U5248 ( .B1(n2599), .B2(keyinput15), .C1(n4900), .C2(keyinput64), 
        .A(n4699), .ZN(n4707) );
  INV_X1 U5249 ( .A(DATAI_6_), .ZN(n4702) );
  INV_X1 U5250 ( .A(DATAI_2_), .ZN(n4701) );
  AOI22_X1 U5251 ( .A1(n4702), .A2(keyinput21), .B1(keyinput35), .B2(n4701), 
        .ZN(n4700) );
  OAI221_X1 U5252 ( .B1(n4702), .B2(keyinput21), .C1(n4701), .C2(keyinput35), 
        .A(n4700), .ZN(n4706) );
  AOI22_X1 U5253 ( .A1(n4704), .A2(keyinput33), .B1(n4908), .B2(keyinput114), 
        .ZN(n4703) );
  OAI221_X1 U5254 ( .B1(n4704), .B2(keyinput33), .C1(n4908), .C2(keyinput114), 
        .A(n4703), .ZN(n4705) );
  NOR4_X1 U5255 ( .A1(n4708), .A2(n4707), .A3(n4706), .A4(n4705), .ZN(n4730)
         );
  INV_X1 U5256 ( .A(REG3_REG_28__SCAN_IN), .ZN(n4910) );
  INV_X1 U5257 ( .A(REG3_REG_19__SCAN_IN), .ZN(n4907) );
  AOI22_X1 U5258 ( .A1(n4910), .A2(keyinput48), .B1(keyinput63), .B2(n4907), 
        .ZN(n4709) );
  OAI221_X1 U5259 ( .B1(n4910), .B2(keyinput48), .C1(n4907), .C2(keyinput63), 
        .A(n4709), .ZN(n4717) );
  XNOR2_X1 U5260 ( .A(REG3_REG_0__SCAN_IN), .B(keyinput54), .ZN(n4713) );
  XNOR2_X1 U5261 ( .A(REG3_REG_1__SCAN_IN), .B(keyinput78), .ZN(n4712) );
  XNOR2_X1 U5262 ( .A(IR_REG_1__SCAN_IN), .B(keyinput87), .ZN(n4711) );
  XNOR2_X1 U5263 ( .A(REG3_REG_13__SCAN_IN), .B(keyinput25), .ZN(n4710) );
  NAND4_X1 U5264 ( .A1(n4713), .A2(n4712), .A3(n4711), .A4(n4710), .ZN(n4716)
         );
  XNOR2_X1 U5265 ( .A(keyinput55), .B(n2680), .ZN(n4715) );
  XNOR2_X1 U5266 ( .A(keyinput86), .B(n4911), .ZN(n4714) );
  NOR4_X1 U5267 ( .A1(n4717), .A2(n4716), .A3(n4715), .A4(n4714), .ZN(n4729)
         );
  XNOR2_X1 U5268 ( .A(IR_REG_5__SCAN_IN), .B(keyinput52), .ZN(n4721) );
  XNOR2_X1 U5269 ( .A(IR_REG_4__SCAN_IN), .B(keyinput1), .ZN(n4720) );
  XNOR2_X1 U5270 ( .A(IR_REG_20__SCAN_IN), .B(keyinput65), .ZN(n4719) );
  XNOR2_X1 U5271 ( .A(IR_REG_8__SCAN_IN), .B(keyinput101), .ZN(n4718) );
  NAND4_X1 U5272 ( .A1(n4721), .A2(n4720), .A3(n4719), .A4(n4718), .ZN(n4727)
         );
  XNOR2_X1 U5273 ( .A(IR_REG_24__SCAN_IN), .B(keyinput77), .ZN(n4725) );
  XNOR2_X1 U5274 ( .A(IR_REG_22__SCAN_IN), .B(keyinput108), .ZN(n4724) );
  XNOR2_X1 U5275 ( .A(IR_REG_28__SCAN_IN), .B(keyinput56), .ZN(n4723) );
  XNOR2_X1 U5276 ( .A(IR_REG_27__SCAN_IN), .B(keyinput120), .ZN(n4722) );
  NAND4_X1 U5277 ( .A1(n4725), .A2(n4724), .A3(n4723), .A4(n4722), .ZN(n4726)
         );
  NOR2_X1 U5278 ( .A1(n4727), .A2(n4726), .ZN(n4728) );
  NAND4_X1 U5279 ( .A1(n4731), .A2(n4730), .A3(n4729), .A4(n4728), .ZN(n4899)
         );
  AOI22_X1 U5280 ( .A1(n4734), .A2(keyinput109), .B1(n4733), .B2(keyinput60), 
        .ZN(n4732) );
  OAI221_X1 U5281 ( .B1(n4734), .B2(keyinput109), .C1(n4733), .C2(keyinput60), 
        .A(n4732), .ZN(n4747) );
  AOI22_X1 U5282 ( .A1(n4737), .A2(keyinput29), .B1(n4736), .B2(keyinput107), 
        .ZN(n4735) );
  OAI221_X1 U5283 ( .B1(n4737), .B2(keyinput29), .C1(n4736), .C2(keyinput107), 
        .A(n4735), .ZN(n4746) );
  AOI22_X1 U5284 ( .A1(n4740), .A2(keyinput105), .B1(keyinput75), .B2(n4739), 
        .ZN(n4738) );
  OAI221_X1 U5285 ( .B1(n4740), .B2(keyinput105), .C1(n4739), .C2(keyinput75), 
        .A(n4738), .ZN(n4745) );
  AOI22_X1 U5286 ( .A1(n4743), .A2(keyinput93), .B1(n4742), .B2(keyinput47), 
        .ZN(n4741) );
  OAI221_X1 U5287 ( .B1(n4743), .B2(keyinput93), .C1(n4742), .C2(keyinput47), 
        .A(n4741), .ZN(n4744) );
  NOR4_X1 U5288 ( .A1(n4747), .A2(n4746), .A3(n4745), .A4(n4744), .ZN(n4787)
         );
  AOI22_X1 U5289 ( .A1(n4750), .A2(keyinput94), .B1(n4749), .B2(keyinput90), 
        .ZN(n4748) );
  OAI221_X1 U5290 ( .B1(n4750), .B2(keyinput94), .C1(n4749), .C2(keyinput90), 
        .A(n4748), .ZN(n4762) );
  AOI22_X1 U5291 ( .A1(n4753), .A2(keyinput88), .B1(keyinput23), .B2(n4752), 
        .ZN(n4751) );
  OAI221_X1 U5292 ( .B1(n4753), .B2(keyinput88), .C1(n4752), .C2(keyinput23), 
        .A(n4751), .ZN(n4761) );
  AOI22_X1 U5293 ( .A1(n4755), .A2(keyinput39), .B1(keyinput5), .B2(n4948), 
        .ZN(n4754) );
  OAI221_X1 U5294 ( .B1(n4755), .B2(keyinput39), .C1(n4948), .C2(keyinput5), 
        .A(n4754), .ZN(n4760) );
  AOI22_X1 U5295 ( .A1(n4758), .A2(keyinput84), .B1(keyinput73), .B2(n4757), 
        .ZN(n4756) );
  OAI221_X1 U5296 ( .B1(n4758), .B2(keyinput84), .C1(n4757), .C2(keyinput73), 
        .A(n4756), .ZN(n4759) );
  NOR4_X1 U5297 ( .A1(n4762), .A2(n4761), .A3(n4760), .A4(n4759), .ZN(n4786)
         );
  INV_X1 U5298 ( .A(REG0_REG_2__SCAN_IN), .ZN(n4765) );
  INV_X1 U5299 ( .A(REG0_REG_5__SCAN_IN), .ZN(n4764) );
  AOI22_X1 U5300 ( .A1(n4765), .A2(keyinput116), .B1(n4764), .B2(keyinput89), 
        .ZN(n4763) );
  OAI221_X1 U5301 ( .B1(n4765), .B2(keyinput116), .C1(n4764), .C2(keyinput89), 
        .A(n4763), .ZN(n4774) );
  INV_X1 U5302 ( .A(REG0_REG_10__SCAN_IN), .ZN(n4767) );
  AOI22_X1 U5303 ( .A1(n4767), .A2(keyinput0), .B1(n3612), .B2(keyinput103), 
        .ZN(n4766) );
  OAI221_X1 U5304 ( .B1(n4767), .B2(keyinput0), .C1(n3612), .C2(keyinput103), 
        .A(n4766), .ZN(n4773) );
  AOI22_X1 U5305 ( .A1(n3713), .A2(keyinput49), .B1(keyinput71), .B2(n4769), 
        .ZN(n4768) );
  OAI221_X1 U5306 ( .B1(n3713), .B2(keyinput49), .C1(n4769), .C2(keyinput71), 
        .A(n4768), .ZN(n4772) );
  INV_X1 U5307 ( .A(REG0_REG_18__SCAN_IN), .ZN(n4933) );
  AOI22_X1 U5308 ( .A1(n4483), .A2(keyinput95), .B1(keyinput125), .B2(n4933), 
        .ZN(n4770) );
  OAI221_X1 U5309 ( .B1(n4483), .B2(keyinput95), .C1(n4933), .C2(keyinput125), 
        .A(n4770), .ZN(n4771) );
  NOR4_X1 U5310 ( .A1(n4774), .A2(n4773), .A3(n4772), .A4(n4771), .ZN(n4785)
         );
  AOI22_X1 U5311 ( .A1(n4470), .A2(keyinput124), .B1(n4932), .B2(keyinput69), 
        .ZN(n4775) );
  OAI221_X1 U5312 ( .B1(n4470), .B2(keyinput124), .C1(n4932), .C2(keyinput69), 
        .A(n4775), .ZN(n4783) );
  INV_X1 U5313 ( .A(REG0_REG_28__SCAN_IN), .ZN(n4777) );
  AOI22_X1 U5314 ( .A1(n4455), .A2(keyinput9), .B1(n4777), .B2(keyinput76), 
        .ZN(n4776) );
  OAI221_X1 U5315 ( .B1(n4455), .B2(keyinput9), .C1(n4777), .C2(keyinput76), 
        .A(n4776), .ZN(n4782) );
  AOI22_X1 U5316 ( .A1(n2353), .A2(keyinput79), .B1(n3117), .B2(keyinput34), 
        .ZN(n4778) );
  OAI221_X1 U5317 ( .B1(n2353), .B2(keyinput79), .C1(n3117), .C2(keyinput34), 
        .A(n4778), .ZN(n4781) );
  AOI22_X1 U5318 ( .A1(n2447), .A2(keyinput67), .B1(keyinput117), .B2(n2508), 
        .ZN(n4779) );
  OAI221_X1 U5319 ( .B1(n2447), .B2(keyinput67), .C1(n2508), .C2(keyinput117), 
        .A(n4779), .ZN(n4780) );
  NOR4_X1 U5320 ( .A1(n4783), .A2(n4782), .A3(n4781), .A4(n4780), .ZN(n4784)
         );
  NAND4_X1 U5321 ( .A1(n4787), .A2(n4786), .A3(n4785), .A4(n4784), .ZN(n4898)
         );
  AOI22_X1 U5322 ( .A1(n3615), .A2(keyinput42), .B1(keyinput62), .B2(n4934), 
        .ZN(n4788) );
  OAI221_X1 U5323 ( .B1(n3615), .B2(keyinput42), .C1(n4934), .C2(keyinput62), 
        .A(n4788), .ZN(n4796) );
  AOI22_X1 U5324 ( .A1(n3693), .A2(keyinput16), .B1(keyinput104), .B2(n4935), 
        .ZN(n4789) );
  OAI221_X1 U5325 ( .B1(n3693), .B2(keyinput16), .C1(n4935), .C2(keyinput104), 
        .A(n4789), .ZN(n4795) );
  AOI22_X1 U5326 ( .A1(n4791), .A2(keyinput72), .B1(n3716), .B2(keyinput57), 
        .ZN(n4790) );
  OAI221_X1 U5327 ( .B1(n4791), .B2(keyinput72), .C1(n3716), .C2(keyinput57), 
        .A(n4790), .ZN(n4794) );
  AOI22_X1 U5328 ( .A1(n4415), .A2(keyinput91), .B1(n4407), .B2(keyinput66), 
        .ZN(n4792) );
  OAI221_X1 U5329 ( .B1(n4415), .B2(keyinput91), .C1(n4407), .C2(keyinput66), 
        .A(n4792), .ZN(n4793) );
  NOR4_X1 U5330 ( .A1(n4796), .A2(n4795), .A3(n4794), .A4(n4793), .ZN(n4837)
         );
  AOI22_X1 U5331 ( .A1(n4798), .A2(keyinput126), .B1(n3065), .B2(keyinput98), 
        .ZN(n4797) );
  OAI221_X1 U5332 ( .B1(n4798), .B2(keyinput126), .C1(n3065), .C2(keyinput98), 
        .A(n4797), .ZN(n4807) );
  AOI22_X1 U5333 ( .A1(n3037), .A2(keyinput13), .B1(keyinput80), .B2(n4361), 
        .ZN(n4799) );
  OAI221_X1 U5334 ( .B1(n3037), .B2(keyinput13), .C1(n4361), .C2(keyinput80), 
        .A(n4799), .ZN(n4806) );
  AOI22_X1 U5335 ( .A1(n4949), .A2(keyinput44), .B1(n4382), .B2(keyinput3), 
        .ZN(n4800) );
  OAI221_X1 U5336 ( .B1(n4949), .B2(keyinput44), .C1(n4382), .C2(keyinput3), 
        .A(n4800), .ZN(n4805) );
  XOR2_X1 U5337 ( .A(n4801), .B(keyinput74), .Z(n4803) );
  XNOR2_X1 U5338 ( .A(REG2_REG_2__SCAN_IN), .B(keyinput68), .ZN(n4802) );
  NAND2_X1 U5339 ( .A1(n4803), .A2(n4802), .ZN(n4804) );
  NOR4_X1 U5340 ( .A1(n4807), .A2(n4806), .A3(n4805), .A4(n4804), .ZN(n4836)
         );
  AOI22_X1 U5341 ( .A1(n4087), .A2(keyinput121), .B1(n4950), .B2(keyinput118), 
        .ZN(n4808) );
  OAI221_X1 U5342 ( .B1(n4087), .B2(keyinput121), .C1(n4950), .C2(keyinput118), 
        .A(n4808), .ZN(n4820) );
  INV_X1 U5343 ( .A(REG2_REG_15__SCAN_IN), .ZN(n4811) );
  AOI22_X1 U5344 ( .A1(n4811), .A2(keyinput113), .B1(keyinput83), .B2(n4810), 
        .ZN(n4809) );
  OAI221_X1 U5345 ( .B1(n4811), .B2(keyinput113), .C1(n4810), .C2(keyinput83), 
        .A(n4809), .ZN(n4819) );
  INV_X1 U5346 ( .A(REG2_REG_20__SCAN_IN), .ZN(n4813) );
  AOI22_X1 U5347 ( .A1(n4813), .A2(keyinput81), .B1(keyinput24), .B2(n4952), 
        .ZN(n4812) );
  OAI221_X1 U5348 ( .B1(n4813), .B2(keyinput81), .C1(n4952), .C2(keyinput24), 
        .A(n4812), .ZN(n4818) );
  INV_X1 U5349 ( .A(REG2_REG_23__SCAN_IN), .ZN(n4816) );
  INV_X1 U5350 ( .A(REG2_REG_22__SCAN_IN), .ZN(n4815) );
  AOI22_X1 U5351 ( .A1(n4816), .A2(keyinput17), .B1(keyinput40), .B2(n4815), 
        .ZN(n4814) );
  OAI221_X1 U5352 ( .B1(n4816), .B2(keyinput17), .C1(n4815), .C2(keyinput40), 
        .A(n4814), .ZN(n4817) );
  NOR4_X1 U5353 ( .A1(n4820), .A2(n4819), .A3(n4818), .A4(n4817), .ZN(n4835)
         );
  INV_X1 U5354 ( .A(REG2_REG_25__SCAN_IN), .ZN(n4953) );
  AOI22_X1 U5355 ( .A1(n4953), .A2(keyinput59), .B1(n4197), .B2(keyinput28), 
        .ZN(n4821) );
  OAI221_X1 U5356 ( .B1(n4953), .B2(keyinput59), .C1(n4197), .C2(keyinput28), 
        .A(n4821), .ZN(n4833) );
  INV_X1 U5357 ( .A(ADDR_REG_17__SCAN_IN), .ZN(n4823) );
  INV_X1 U5358 ( .A(ADDR_REG_18__SCAN_IN), .ZN(n4951) );
  AOI22_X1 U5359 ( .A1(n4823), .A2(keyinput92), .B1(n4951), .B2(keyinput4), 
        .ZN(n4822) );
  OAI221_X1 U5360 ( .B1(n4823), .B2(keyinput92), .C1(n4951), .C2(keyinput4), 
        .A(n4822), .ZN(n4832) );
  INV_X1 U5361 ( .A(ADDR_REG_15__SCAN_IN), .ZN(n4826) );
  INV_X1 U5362 ( .A(ADDR_REG_13__SCAN_IN), .ZN(n4825) );
  AOI22_X1 U5363 ( .A1(n4826), .A2(keyinput43), .B1(keyinput10), .B2(n4825), 
        .ZN(n4824) );
  OAI221_X1 U5364 ( .B1(n4826), .B2(keyinput43), .C1(n4825), .C2(keyinput10), 
        .A(n4824), .ZN(n4831) );
  INV_X1 U5365 ( .A(ADDR_REG_10__SCAN_IN), .ZN(n4829) );
  INV_X1 U5366 ( .A(ADDR_REG_12__SCAN_IN), .ZN(n4828) );
  AOI22_X1 U5367 ( .A1(n4829), .A2(keyinput82), .B1(n4828), .B2(keyinput102), 
        .ZN(n4827) );
  OAI221_X1 U5368 ( .B1(n4829), .B2(keyinput82), .C1(n4828), .C2(keyinput102), 
        .A(n4827), .ZN(n4830) );
  NOR4_X1 U5369 ( .A1(n4833), .A2(n4832), .A3(n4831), .A4(n4830), .ZN(n4834)
         );
  NAND4_X1 U5370 ( .A1(n4837), .A2(n4836), .A3(n4835), .A4(n4834), .ZN(n4897)
         );
  INV_X1 U5371 ( .A(keyinput19), .ZN(n4839) );
  OAI22_X1 U5372 ( .A1(keyinput37), .A2(n4840), .B1(n4839), .B2(
        DATAO_REG_1__SCAN_IN), .ZN(n4838) );
  AOI221_X1 U5373 ( .B1(n4840), .B2(keyinput37), .C1(n4839), .C2(
        DATAO_REG_1__SCAN_IN), .A(n4838), .ZN(n4895) );
  OAI22_X1 U5374 ( .A1(keyinput14), .A2(n4918), .B1(n4842), .B2(keyinput36), 
        .ZN(n4841) );
  AOI221_X1 U5375 ( .B1(n4918), .B2(keyinput14), .C1(n4842), .C2(keyinput36), 
        .A(n4841), .ZN(n4894) );
  INV_X1 U5376 ( .A(DATAO_REG_5__SCAN_IN), .ZN(n4977) );
  XNOR2_X1 U5377 ( .A(keyinput70), .B(n4977), .ZN(n4849) );
  XNOR2_X1 U5378 ( .A(keyinput122), .B(n4843), .ZN(n4848) );
  XNOR2_X1 U5379 ( .A(keyinput111), .B(n4844), .ZN(n4847) );
  XNOR2_X1 U5380 ( .A(keyinput27), .B(n4845), .ZN(n4846) );
  NOR4_X1 U5381 ( .A1(n4849), .A2(n4848), .A3(n4847), .A4(n4846), .ZN(n4893)
         );
  XNOR2_X1 U5382 ( .A(keyinput20), .B(n4920), .ZN(n4891) );
  XNOR2_X1 U5383 ( .A(keyinput112), .B(n4850), .ZN(n4890) );
  OAI22_X1 U5384 ( .A1(keyinput119), .A2(n4928), .B1(n4852), .B2(keyinput22), 
        .ZN(n4851) );
  AOI221_X1 U5385 ( .B1(n4928), .B2(keyinput119), .C1(n4852), .C2(keyinput22), 
        .A(n4851), .ZN(n4861) );
  OAI22_X1 U5386 ( .A1(keyinput26), .A2(n4855), .B1(n4854), .B2(keyinput41), 
        .ZN(n4853) );
  AOI221_X1 U5387 ( .B1(n4855), .B2(keyinput26), .C1(n4854), .C2(keyinput41), 
        .A(n4853), .ZN(n4860) );
  XOR2_X1 U5388 ( .A(keyinput53), .B(n4856), .Z(n4859) );
  XOR2_X1 U5389 ( .A(keyinput8), .B(n4857), .Z(n4858) );
  NAND4_X1 U5390 ( .A1(n4861), .A2(n4860), .A3(n4859), .A4(n4858), .ZN(n4889)
         );
  INV_X1 U5391 ( .A(ADDR_REG_5__SCAN_IN), .ZN(n4863) );
  INV_X1 U5392 ( .A(ADDR_REG_6__SCAN_IN), .ZN(n4954) );
  OAI22_X1 U5393 ( .A1(keyinput106), .A2(n4863), .B1(n4954), .B2(keyinput46), 
        .ZN(n4862) );
  AOI221_X1 U5394 ( .B1(n4863), .B2(keyinput106), .C1(n4954), .C2(keyinput46), 
        .A(n4862), .ZN(n4887) );
  XOR2_X1 U5395 ( .A(keyinput100), .B(ADDR_REG_3__SCAN_IN), .Z(n4872) );
  XOR2_X1 U5396 ( .A(ADDR_REG_4__SCAN_IN), .B(keyinput12), .Z(n4871) );
  INV_X1 U5397 ( .A(ADDR_REG_9__SCAN_IN), .ZN(n4865) );
  INV_X1 U5398 ( .A(ADDR_REG_8__SCAN_IN), .ZN(n4955) );
  AOI22_X1 U5399 ( .A1(n4865), .A2(keyinput51), .B1(keyinput30), .B2(n4955), 
        .ZN(n4864) );
  OAI221_X1 U5400 ( .B1(n4865), .B2(keyinput51), .C1(n4955), .C2(keyinput30), 
        .A(n4864), .ZN(n4870) );
  INV_X1 U5401 ( .A(ADDR_REG_2__SCAN_IN), .ZN(n4868) );
  INV_X1 U5402 ( .A(keyinput31), .ZN(n4867) );
  AOI22_X1 U5403 ( .A1(n4868), .A2(keyinput11), .B1(ADDR_REG_0__SCAN_IN), .B2(
        n4867), .ZN(n4866) );
  OAI221_X1 U5404 ( .B1(n4868), .B2(keyinput11), .C1(n4867), .C2(
        ADDR_REG_0__SCAN_IN), .A(n4866), .ZN(n4869) );
  NOR4_X1 U5405 ( .A1(n4872), .A2(n4871), .A3(n4870), .A4(n4869), .ZN(n4886)
         );
  INV_X1 U5406 ( .A(DATAO_REG_29__SCAN_IN), .ZN(n4874) );
  OAI22_X1 U5407 ( .A1(keyinput85), .A2(n4922), .B1(n4874), .B2(keyinput58), 
        .ZN(n4873) );
  AOI221_X1 U5408 ( .B1(n4922), .B2(keyinput85), .C1(n4874), .C2(keyinput58), 
        .A(n4873), .ZN(n4885) );
  AOI22_X1 U5409 ( .A1(n4877), .A2(keyinput110), .B1(n4876), .B2(keyinput6), 
        .ZN(n4875) );
  OAI221_X1 U5410 ( .B1(n4877), .B2(keyinput110), .C1(n4876), .C2(keyinput6), 
        .A(n4875), .ZN(n4883) );
  AOI22_X1 U5411 ( .A1(n4923), .A2(keyinput38), .B1(n4926), .B2(keyinput99), 
        .ZN(n4878) );
  OAI221_X1 U5412 ( .B1(n4923), .B2(keyinput38), .C1(n4926), .C2(keyinput99), 
        .A(n4878), .ZN(n4882) );
  XNOR2_X1 U5413 ( .A(n2345), .B(keyinput18), .ZN(n4881) );
  INV_X1 U5414 ( .A(ADDR_REG_11__SCAN_IN), .ZN(n4879) );
  XNOR2_X1 U5415 ( .A(n4879), .B(keyinput127), .ZN(n4880) );
  NOR4_X1 U5416 ( .A1(n4883), .A2(n4882), .A3(n4881), .A4(n4880), .ZN(n4884)
         );
  NAND4_X1 U5417 ( .A1(n4887), .A2(n4886), .A3(n4885), .A4(n4884), .ZN(n4888)
         );
  NOR4_X1 U5418 ( .A1(n4891), .A2(n4890), .A3(n4889), .A4(n4888), .ZN(n4892)
         );
  NAND4_X1 U5419 ( .A1(n4895), .A2(n4894), .A3(n4893), .A4(n4892), .ZN(n4896)
         );
  NOR4_X1 U5420 ( .A1(n4899), .A2(n4898), .A3(n4897), .A4(n4896), .ZN(n4983)
         );
  NOR4_X1 U5421 ( .A1(DATAI_15_), .A2(DATAI_13_), .A3(DATAI_12_), .A4(n4900), 
        .ZN(n4974) );
  NOR4_X1 U5422 ( .A1(DATAI_22_), .A2(DATAI_21_), .A3(DATAI_19_), .A4(n4901), 
        .ZN(n4973) );
  NAND4_X1 U5423 ( .A1(DATAI_29_), .A2(DATAI_30_), .A3(n4903), .A4(n4902), 
        .ZN(n4917) );
  INV_X1 U5424 ( .A(IR_REG_5__SCAN_IN), .ZN(n4905) );
  NOR4_X1 U5425 ( .A1(n4905), .A2(n4904), .A3(n2253), .A4(IR_REG_1__SCAN_IN), 
        .ZN(n4915) );
  NOR4_X1 U5426 ( .A1(n4907), .A2(n4906), .A3(REG3_REG_17__SCAN_IN), .A4(
        REG3_REG_13__SCAN_IN), .ZN(n4914) );
  OR4_X1 U5427 ( .A1(DATAI_2_), .A2(DATAI_6_), .A3(DATAI_0_), .A4(n4908), .ZN(
        n4909) );
  NOR4_X1 U5428 ( .A1(n4912), .A2(n4911), .A3(n4910), .A4(n4909), .ZN(n4913)
         );
  NAND4_X1 U5429 ( .A1(n4915), .A2(REG3_REG_1__SCAN_IN), .A3(n4914), .A4(n4913), .ZN(n4916) );
  NOR4_X1 U5430 ( .A1(IR_REG_30__SCAN_IN), .A2(ADDR_REG_11__SCAN_IN), .A3(
        n4917), .A4(n4916), .ZN(n4972) );
  NAND4_X1 U5431 ( .A1(DATAO_REG_5__SCAN_IN), .A2(DATAO_REG_1__SCAN_IN), .A3(
        DATAO_REG_3__SCAN_IN), .A4(n4918), .ZN(n4970) );
  INV_X1 U5432 ( .A(ADDR_REG_0__SCAN_IN), .ZN(n4919) );
  NAND4_X1 U5433 ( .A1(ADDR_REG_3__SCAN_IN), .A2(ADDR_REG_2__SCAN_IN), .A3(
        DATAO_REG_0__SCAN_IN), .A4(n4919), .ZN(n4969) );
  NAND4_X1 U5434 ( .A1(DATAO_REG_17__SCAN_IN), .A2(DATAO_REG_19__SCAN_IN), 
        .A3(DATAO_REG_20__SCAN_IN), .A4(n4920), .ZN(n4921) );
  NOR3_X1 U5435 ( .A1(DATAO_REG_8__SCAN_IN), .A2(DATAO_REG_14__SCAN_IN), .A3(
        n4921), .ZN(n4930) );
  NOR4_X1 U5436 ( .A1(DATAO_REG_23__SCAN_IN), .A2(DATAO_REG_29__SCAN_IN), .A3(
        n4923), .A4(n4922), .ZN(n4924) );
  NAND3_X1 U5437 ( .A1(DATAO_REG_21__SCAN_IN), .A2(DATAO_REG_28__SCAN_IN), 
        .A3(n4924), .ZN(n4925) );
  NOR4_X1 U5438 ( .A1(REG3_REG_22__SCAN_IN), .A2(n4927), .A3(n4926), .A4(n4925), .ZN(n4929) );
  NAND4_X1 U5439 ( .A1(DATAO_REG_12__SCAN_IN), .A2(n4930), .A3(n4929), .A4(
        n4928), .ZN(n4968) );
  NOR4_X1 U5440 ( .A1(REG0_REG_10__SCAN_IN), .A2(REG0_REG_11__SCAN_IN), .A3(
        REG0_REG_5__SCAN_IN), .A4(n3713), .ZN(n4931) );
  NAND3_X1 U5441 ( .A1(D_REG_18__SCAN_IN), .A2(D_REG_24__SCAN_IN), .A3(n4931), 
        .ZN(n4947) );
  NAND4_X1 U5442 ( .A1(REG0_REG_28__SCAN_IN), .A2(REG1_REG_1__SCAN_IN), .A3(
        n4932), .A4(n4455), .ZN(n4939) );
  NAND4_X1 U5443 ( .A1(REG0_REG_17__SCAN_IN), .A2(REG0_REG_21__SCAN_IN), .A3(
        REG0_REG_14__SCAN_IN), .A4(n4933), .ZN(n4938) );
  NAND4_X1 U5444 ( .A1(REG1_REG_18__SCAN_IN), .A2(n3693), .A3(n4935), .A4(
        n4934), .ZN(n4937) );
  NAND4_X1 U5445 ( .A1(REG1_REG_4__SCAN_IN), .A2(REG1_REG_2__SCAN_IN), .A3(
        n3615), .A4(n2508), .ZN(n4936) );
  NOR4_X1 U5446 ( .A1(n4939), .A2(n4938), .A3(n4937), .A4(n4936), .ZN(n4945)
         );
  NAND4_X1 U5447 ( .A1(n4941), .A2(n4940), .A3(IR_REG_22__SCAN_IN), .A4(
        IR_REG_28__SCAN_IN), .ZN(n4943) );
  NAND4_X1 U5448 ( .A1(D_REG_1__SCAN_IN), .A2(D_REG_10__SCAN_IN), .A3(
        D_REG_3__SCAN_IN), .A4(D_REG_6__SCAN_IN), .ZN(n4942) );
  NOR2_X1 U5449 ( .A1(n4943), .A2(n4942), .ZN(n4944) );
  NAND2_X1 U5450 ( .A1(n4945), .A2(n4944), .ZN(n4946) );
  NOR4_X1 U5451 ( .A1(REG0_REG_2__SCAN_IN), .A2(n4948), .A3(n4947), .A4(n4946), 
        .ZN(n4966) );
  NOR4_X1 U5452 ( .A1(REG1_REG_29__SCAN_IN), .A2(REG1_REG_26__SCAN_IN), .A3(
        REG1_REG_25__SCAN_IN), .A4(REG1_REG_30__SCAN_IN), .ZN(n4965) );
  NOR4_X1 U5453 ( .A1(REG1_REG_15__SCAN_IN), .A2(n4415), .A3(n4407), .A4(n4949), .ZN(n4964) );
  NAND4_X1 U5454 ( .A1(REG2_REG_15__SCAN_IN), .A2(REG2_REG_20__SCAN_IN), .A3(
        REG2_REG_14__SCAN_IN), .A4(n4950), .ZN(n4962) );
  NAND4_X1 U5455 ( .A1(REG2_REG_5__SCAN_IN), .A2(REG2_REG_2__SCAN_IN), .A3(
        REG1_REG_31__SCAN_IN), .A4(n4087), .ZN(n4961) );
  NOR4_X1 U5456 ( .A1(ADDR_REG_17__SCAN_IN), .A2(ADDR_REG_15__SCAN_IN), .A3(
        n4951), .A4(n4197), .ZN(n4959) );
  NOR4_X1 U5457 ( .A1(REG2_REG_22__SCAN_IN), .A2(REG2_REG_23__SCAN_IN), .A3(
        n4953), .A4(n4952), .ZN(n4958) );
  NOR4_X1 U5458 ( .A1(ADDR_REG_4__SCAN_IN), .A2(ADDR_REG_9__SCAN_IN), .A3(
        ADDR_REG_5__SCAN_IN), .A4(n4954), .ZN(n4957) );
  NOR4_X1 U5459 ( .A1(ADDR_REG_13__SCAN_IN), .A2(ADDR_REG_12__SCAN_IN), .A3(
        ADDR_REG_10__SCAN_IN), .A4(n4955), .ZN(n4956) );
  NAND4_X1 U5460 ( .A1(n4959), .A2(n4958), .A3(n4957), .A4(n4956), .ZN(n4960)
         );
  NOR3_X1 U5461 ( .A1(n4962), .A2(n4961), .A3(n4960), .ZN(n4963) );
  NAND4_X1 U5462 ( .A1(n4966), .A2(n4965), .A3(n4964), .A4(n4963), .ZN(n4967)
         );
  NOR4_X1 U5463 ( .A1(n4970), .A2(n4969), .A3(n4968), .A4(n4967), .ZN(n4971)
         );
  NAND4_X1 U5464 ( .A1(n4974), .A2(n4973), .A3(n4972), .A4(n4971), .ZN(n4980)
         );
  NAND3_X1 U5465 ( .A1(n4981), .A2(U4043), .A3(n4980), .ZN(n4979) );
  INV_X1 U5466 ( .A(n4980), .ZN(n4976) );
  OAI21_X1 U5467 ( .B1(n4977), .B2(n4976), .A(n4975), .ZN(n4978) );
  OAI211_X1 U5468 ( .C1(n4981), .C2(n4980), .A(n4979), .B(n4978), .ZN(n4982)
         );
  XNOR2_X1 U5469 ( .A(n4983), .B(n4982), .ZN(U3555) );
  CLKBUF_X3 U2388 ( .A(n2426), .Z(n3904) );
  CLKBUF_X1 U2395 ( .A(n2489), .Z(n3905) );
  CLKBUF_X1 U2477 ( .A(n2446), .Z(n3908) );
endmodule

