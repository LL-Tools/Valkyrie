

module b14_C_gen_AntiSAT_k_256_6 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, keyinput_f0, keyinput_f1, 
        keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, 
        keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, 
        keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, 
        keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, 
        keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, 
        keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, 
        keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, 
        keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, 
        keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, 
        keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, 
        keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, 
        keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, 
        keyinput_f62, keyinput_f63, keyinput_f64, keyinput_f65, keyinput_f66, 
        keyinput_f67, keyinput_f68, keyinput_f69, keyinput_f70, keyinput_f71, 
        keyinput_f72, keyinput_f73, keyinput_f74, keyinput_f75, keyinput_f76, 
        keyinput_f77, keyinput_f78, keyinput_f79, keyinput_f80, keyinput_f81, 
        keyinput_f82, keyinput_f83, keyinput_f84, keyinput_f85, keyinput_f86, 
        keyinput_f87, keyinput_f88, keyinput_f89, keyinput_f90, keyinput_f91, 
        keyinput_f92, keyinput_f93, keyinput_f94, keyinput_f95, keyinput_f96, 
        keyinput_f97, keyinput_f98, keyinput_f99, keyinput_f100, keyinput_f101, 
        keyinput_f102, keyinput_f103, keyinput_f104, keyinput_f105, 
        keyinput_f106, keyinput_f107, keyinput_f108, keyinput_f109, 
        keyinput_f110, keyinput_f111, keyinput_f112, keyinput_f113, 
        keyinput_f114, keyinput_f115, keyinput_f116, keyinput_f117, 
        keyinput_f118, keyinput_f119, keyinput_f120, keyinput_f121, 
        keyinput_f122, keyinput_f123, keyinput_f124, keyinput_f125, 
        keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1, keyinput_g2, 
        keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7, 
        keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12, 
        keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17, 
        keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22, 
        keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27, 
        keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32, 
        keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37, 
        keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42, 
        keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47, 
        keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52, 
        keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57, 
        keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62, 
        keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66, keyinput_g67, 
        keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71, keyinput_g72, 
        keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76, keyinput_g77, 
        keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81, keyinput_g82, 
        keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86, keyinput_g87, 
        keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91, keyinput_g92, 
        keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96, keyinput_g97, 
        keyinput_g98, keyinput_g99, keyinput_g100, keyinput_g101, 
        keyinput_g102, keyinput_g103, keyinput_g104, keyinput_g105, 
        keyinput_g106, keyinput_g107, keyinput_g108, keyinput_g109, 
        keyinput_g110, keyinput_g111, keyinput_g112, keyinput_g113, 
        keyinput_g114, keyinput_g115, keyinput_g116, keyinput_g117, 
        keyinput_g118, keyinput_g119, keyinput_g120, keyinput_g121, 
        keyinput_g122, keyinput_g123, keyinput_g124, keyinput_g125, 
        keyinput_g126, keyinput_g127, U3352, U3351, U3350, U3349, U3348, U3347, 
        U3346, U3345, U3344, U3343, U3342, U3341, U3340, U3339, U3338, U3337, 
        U3336, U3335, U3334, U3333, U3332, U3331, U3330, U3329, U3328, U3327, 
        U3326, U3325, U3324, U3323, U3322, U3321, U3458, U3459, U3320, U3319, 
        U3318, U3317, U3316, U3315, U3314, U3313, U3312, U3311, U3310, U3309, 
        U3308, U3307, U3306, U3305, U3304, U3303, U3302, U3301, U3300, U3299, 
        U3298, U3297, U3296, U3295, U3294, U3293, U3292, U3291, U3467, U3469, 
        U3471, U3473, U3475, U3477, U3479, U3481, U3483, U3485, U3487, U3489, 
        U3491, U3493, U3495, U3497, U3499, U3501, U3503, U3505, U3506, U3507, 
        U3508, U3509, U3510, U3511, U3512, U3513, U3514, U3515, U3516, U3517, 
        U3518, U3519, U3520, U3521, U3522, U3523, U3524, U3525, U3526, U3527, 
        U3528, U3529, U3530, U3531, U3532, U3533, U3534, U3535, U3536, U3537, 
        U3538, U3539, U3540, U3541, U3542, U3543, U3544, U3545, U3546, U3547, 
        U3548, U3549, U3290, U3289, U3288, U3287, U3286, U3285, U3284, U3283, 
        U3282, U3281, U3280, U3279, U3278, U3277, U3276, U3275, U3274, U3273, 
        U3272, U3271, U3270, U3269, U3268, U3267, U3266, U3265, U3264, U3263, 
        U3262, U3354, U3261, U3260, U3259, U3258, U3257, U3256, U3255, U3254, 
        U3253, U3252, U3251, U3250, U3249, U3248, U3247, U3246, U3245, U3244, 
        U3243, U3242, U3241, U3240, U3550, U3551, U3552, U3553, U3554, U3555, 
        U3556, U3557, U3558, U3559, U3560, U3561, U3562, U3563, U3564, U3565, 
        U3566, U3567, U3568, U3569, U3570, U3571, U3572, U3573, U3574, U3575, 
        U3576, U3577, U3578, U3579, U3580, U3581, U3239, U3238, U3237, U3236, 
        U3235, U3234, U3233, U3232, U3231, U3230, U3229, U3228, U3227, U3226, 
        U3225, U3224, U3223, U3222, U3221, U3220, U3219, U3218, U3217, U3216, 
        U3215, U3214, U3213, U3212, U3211, U3210, U3149, U3148, U4043 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN, keyinput_f0, keyinput_f1, keyinput_f2,
         keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, keyinput_f7,
         keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, keyinput_f12,
         keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, keyinput_f17,
         keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, keyinput_f22,
         keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, keyinput_f27,
         keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, keyinput_f32,
         keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, keyinput_f37,
         keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, keyinput_f42,
         keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, keyinput_f47,
         keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, keyinput_f52,
         keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, keyinput_f57,
         keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, keyinput_f62,
         keyinput_f63, keyinput_f64, keyinput_f65, keyinput_f66, keyinput_f67,
         keyinput_f68, keyinput_f69, keyinput_f70, keyinput_f71, keyinput_f72,
         keyinput_f73, keyinput_f74, keyinput_f75, keyinput_f76, keyinput_f77,
         keyinput_f78, keyinput_f79, keyinput_f80, keyinput_f81, keyinput_f82,
         keyinput_f83, keyinput_f84, keyinput_f85, keyinput_f86, keyinput_f87,
         keyinput_f88, keyinput_f89, keyinput_f90, keyinput_f91, keyinput_f92,
         keyinput_f93, keyinput_f94, keyinput_f95, keyinput_f96, keyinput_f97,
         keyinput_f98, keyinput_f99, keyinput_f100, keyinput_f101,
         keyinput_f102, keyinput_f103, keyinput_f104, keyinput_f105,
         keyinput_f106, keyinput_f107, keyinput_f108, keyinput_f109,
         keyinput_f110, keyinput_f111, keyinput_f112, keyinput_f113,
         keyinput_f114, keyinput_f115, keyinput_f116, keyinput_f117,
         keyinput_f118, keyinput_f119, keyinput_f120, keyinput_f121,
         keyinput_f122, keyinput_f123, keyinput_f124, keyinput_f125,
         keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1, keyinput_g2,
         keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7,
         keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12,
         keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17,
         keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22,
         keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27,
         keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32,
         keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37,
         keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42,
         keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47,
         keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52,
         keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57,
         keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62,
         keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66, keyinput_g67,
         keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71, keyinput_g72,
         keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76, keyinput_g77,
         keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81, keyinput_g82,
         keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86, keyinput_g87,
         keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91, keyinput_g92,
         keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96, keyinput_g97,
         keyinput_g98, keyinput_g99, keyinput_g100, keyinput_g101,
         keyinput_g102, keyinput_g103, keyinput_g104, keyinput_g105,
         keyinput_g106, keyinput_g107, keyinput_g108, keyinput_g109,
         keyinput_g110, keyinput_g111, keyinput_g112, keyinput_g113,
         keyinput_g114, keyinput_g115, keyinput_g116, keyinput_g117,
         keyinput_g118, keyinput_g119, keyinput_g120, keyinput_g121,
         keyinput_g122, keyinput_g123, keyinput_g124, keyinput_g125,
         keyinput_g126, keyinput_g127;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227,
         n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237,
         n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247,
         n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257,
         n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267,
         n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277,
         n2278, n2279, n2280, n2281, n2282, n2284, n2285, n2286, n2287, n2288,
         n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298,
         n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308,
         n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318,
         n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328,
         n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338,
         n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348,
         n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358,
         n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368,
         n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378,
         n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388,
         n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398,
         n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408,
         n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418,
         n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428,
         n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438,
         n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448,
         n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458,
         n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468,
         n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478,
         n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488,
         n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498,
         n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508,
         n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518,
         n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528,
         n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538,
         n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548,
         n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558,
         n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568,
         n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578,
         n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588,
         n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598,
         n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608,
         n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618,
         n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628,
         n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638,
         n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648,
         n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658,
         n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668,
         n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678,
         n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688,
         n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698,
         n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708,
         n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718,
         n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728,
         n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738,
         n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748,
         n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758,
         n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768,
         n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778,
         n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788,
         n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798,
         n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808,
         n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818,
         n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828,
         n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838,
         n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848,
         n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858,
         n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868,
         n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878,
         n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888,
         n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898,
         n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908,
         n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918,
         n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928,
         n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938,
         n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948,
         n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958,
         n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968,
         n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978,
         n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988,
         n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998,
         n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008,
         n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018,
         n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028,
         n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038,
         n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048,
         n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058,
         n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068,
         n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078,
         n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088,
         n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098,
         n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108,
         n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118,
         n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128,
         n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138,
         n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148,
         n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158,
         n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168,
         n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178,
         n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188,
         n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198,
         n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208,
         n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218,
         n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228,
         n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238,
         n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248,
         n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258,
         n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268,
         n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278,
         n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288,
         n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298,
         n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308,
         n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318,
         n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328,
         n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338,
         n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348,
         n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358,
         n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368,
         n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378,
         n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388,
         n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398,
         n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408,
         n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418,
         n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428,
         n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438,
         n3439, n3440, n3441, n3442, n3443, n3445, n3446, n3447, n3448, n3449,
         n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459,
         n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469,
         n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479,
         n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489,
         n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499,
         n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509,
         n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519,
         n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529,
         n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539,
         n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549,
         n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559,
         n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569,
         n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579,
         n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589,
         n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599,
         n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609,
         n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619,
         n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629,
         n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639,
         n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649,
         n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659,
         n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669,
         n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679,
         n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689,
         n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699,
         n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709,
         n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719,
         n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729,
         n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739,
         n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749,
         n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759,
         n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769,
         n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779,
         n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789,
         n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799,
         n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809,
         n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819,
         n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829,
         n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839,
         n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849,
         n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859,
         n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869,
         n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879,
         n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889,
         n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899,
         n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909,
         n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919,
         n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929,
         n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939,
         n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949,
         n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959,
         n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969,
         n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979,
         n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989,
         n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999,
         n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009,
         n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019,
         n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029,
         n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039,
         n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049,
         n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059,
         n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069,
         n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079,
         n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089,
         n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099,
         n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109,
         n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119,
         n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129,
         n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139,
         n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149,
         n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159,
         n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169,
         n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179,
         n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189,
         n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199,
         n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209,
         n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219,
         n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229,
         n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239,
         n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249,
         n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259,
         n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269,
         n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279,
         n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289,
         n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299,
         n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309,
         n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319,
         n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329,
         n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339,
         n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349,
         n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359,
         n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369,
         n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379,
         n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389,
         n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399,
         n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409,
         n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419,
         n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429,
         n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439,
         n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449,
         n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459,
         n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469,
         n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479,
         n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489,
         n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499,
         n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509,
         n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519,
         n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529,
         n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539,
         n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549,
         n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559,
         n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569,
         n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579,
         n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589,
         n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599,
         n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609,
         n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619,
         n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629,
         n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639,
         n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649,
         n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659,
         n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669,
         n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679,
         n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689,
         n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699,
         n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709,
         n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719,
         n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729,
         n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739,
         n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749,
         n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759,
         n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769,
         n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779,
         n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789,
         n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799,
         n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809,
         n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819,
         n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829,
         n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839,
         n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849,
         n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859,
         n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869,
         n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879,
         n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889,
         n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899,
         n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909,
         n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919,
         n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929,
         n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939,
         n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949,
         n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959,
         n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969,
         n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979,
         n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989,
         n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999,
         n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009,
         n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018;

  CLKBUF_X2 U2460 ( .A(n2499), .Z(n2659) );
  BUF_X1 U2461 ( .A(n2485), .Z(n2218) );
  INV_X1 U2462 ( .A(n3438), .ZN(n2352) );
  NAND2_X1 U2464 ( .A1(n3774), .A2(n3703), .ZN(n2915) );
  AND2_X2 U2467 ( .A1(n2420), .A2(n2620), .ZN(n2669) );
  NOR2_X4 U2468 ( .A1(n2531), .A2(n2438), .ZN(n2620) );
  NAND2_X1 U2469 ( .A1(n2877), .A2(n4231), .ZN(n3621) );
  OAI21_X1 U2470 ( .B1(n2965), .B2(n2352), .A(n2351), .ZN(n2350) );
  NAND2_X1 U2471 ( .A1(n2483), .A2(n2895), .ZN(n2744) );
  NAND4_X1 U2472 ( .A1(n2497), .A2(n2496), .A3(n2495), .A4(n2494), .ZN(n3794)
         );
  AND2_X1 U2473 ( .A1(n4373), .A2(n2452), .ZN(n2485) );
  MUX2_X1 U2474 ( .A(REG0_REG_28__SCAN_IN), .B(n4248), .S(n4631), .Z(n2813) );
  MUX2_X1 U2475 ( .A(REG1_REG_28__SCAN_IN), .B(n4248), .S(n4646), .Z(n4249) );
  NOR2_X1 U2476 ( .A1(n2309), .A2(n2311), .ZN(n2307) );
  AND2_X1 U2477 ( .A1(n3952), .A2(n4622), .ZN(n2309) );
  OAI21_X1 U2478 ( .B1(n3132), .B2(n3131), .A(n3130), .ZN(n2354) );
  OAI21_X1 U2479 ( .B1(n3062), .B2(n2273), .A(n2239), .ZN(n2274) );
  NAND2_X1 U2480 ( .A1(n2401), .A2(n2542), .ZN(n3062) );
  NAND2_X1 U2481 ( .A1(n2396), .A2(n2221), .ZN(n2401) );
  NAND2_X1 U2482 ( .A1(n2333), .A2(n2332), .ZN(n3036) );
  NAND2_X1 U2483 ( .A1(n4631), .A2(n4629), .ZN(n4371) );
  NAND2_X1 U2484 ( .A1(n3705), .A2(n3708), .ZN(n3660) );
  NAND4_X1 U2485 ( .A1(n2507), .A2(n2506), .A3(n2505), .A4(n2504), .ZN(n3793)
         );
  NAND4_X1 U2486 ( .A1(n2475), .A2(n2474), .A3(n2473), .A4(n2472), .ZN(n2885)
         );
  AND2_X2 U2487 ( .A1(n3438), .A2(n4606), .ZN(n3282) );
  NAND2_X1 U2488 ( .A1(n2789), .A2(IR_REG_31__SCAN_IN), .ZN(n2790) );
  XNOR2_X1 U2489 ( .A(n2449), .B(IR_REG_29__SCAN_IN), .ZN(n2838) );
  XNOR2_X1 U2490 ( .A(n2740), .B(n2739), .ZN(n3774) );
  AND4_X1 U2491 ( .A1(n2420), .A2(n2620), .A3(n4801), .A4(n2670), .ZN(n2313)
         );
  AND2_X1 U2492 ( .A1(n2422), .A2(n2421), .ZN(n2420) );
  AND2_X1 U2493 ( .A1(n2236), .A2(n2423), .ZN(n2422) );
  AND2_X1 U2494 ( .A1(n2388), .A2(n2394), .ZN(n2477) );
  AND2_X1 U2495 ( .A1(n2439), .A2(n2424), .ZN(n2423) );
  INV_X1 U2496 ( .A(IR_REG_31__SCAN_IN), .ZN(n2459) );
  INV_X1 U2497 ( .A(IR_REG_19__SCAN_IN), .ZN(n2683) );
  INV_X1 U2498 ( .A(IR_REG_3__SCAN_IN), .ZN(n2519) );
  NOR2_X1 U2499 ( .A1(IR_REG_4__SCAN_IN), .A2(IR_REG_1__SCAN_IN), .ZN(n2393)
         );
  NOR2_X1 U2500 ( .A1(IR_REG_9__SCAN_IN), .A2(IR_REG_5__SCAN_IN), .ZN(n2437)
         );
  INV_X1 U2501 ( .A(IR_REG_16__SCAN_IN), .ZN(n4896) );
  NOR2_X1 U2502 ( .A1(IR_REG_10__SCAN_IN), .A2(IR_REG_6__SCAN_IN), .ZN(n2436)
         );
  NOR2_X1 U2503 ( .A1(IR_REG_7__SCAN_IN), .A2(IR_REG_8__SCAN_IN), .ZN(n2575)
         );
  NOR2_X1 U2504 ( .A1(IR_REG_11__SCAN_IN), .A2(IR_REG_12__SCAN_IN), .ZN(n2435)
         );
  INV_X4 U2505 ( .A(n2290), .ZN(n2502) );
  NAND2_X1 U2506 ( .A1(n2260), .A2(n2258), .ZN(n4187) );
  AOI21_X1 U2507 ( .B1(n2262), .B2(n2264), .A(n2259), .ZN(n2258) );
  INV_X1 U2508 ( .A(n3223), .ZN(n2259) );
  NAND2_X1 U2509 ( .A1(n3969), .A2(n3447), .ZN(n2828) );
  NAND2_X1 U2510 ( .A1(n2375), .A2(n2373), .ZN(n2372) );
  INV_X1 U2511 ( .A(n2378), .ZN(n2373) );
  OR2_X1 U2512 ( .A1(n3716), .A2(n2273), .ZN(n2272) );
  NAND2_X1 U2513 ( .A1(n2317), .A2(n2315), .ZN(n3083) );
  INV_X1 U2514 ( .A(n2316), .ZN(n2315) );
  OAI21_X1 U2515 ( .B1(n2319), .B2(n3711), .A(n3724), .ZN(n2316) );
  NAND2_X1 U2516 ( .A1(n3040), .A2(n3792), .ZN(n3714) );
  OR2_X1 U2517 ( .A1(n3794), .A2(n2984), .ZN(n3705) );
  NOR2_X1 U2518 ( .A1(n2430), .A2(IR_REG_22__SCAN_IN), .ZN(n2429) );
  NAND2_X1 U2519 ( .A1(n2431), .A2(n2441), .ZN(n2430) );
  INV_X1 U2520 ( .A(n2440), .ZN(n2431) );
  OAI21_X1 U2521 ( .B1(n3278), .B2(n2382), .A(n2380), .ZN(n3319) );
  AOI21_X1 U2522 ( .B1(n3305), .B2(n2383), .A(n2381), .ZN(n2380) );
  INV_X1 U2523 ( .A(n3305), .ZN(n2382) );
  NAND2_X1 U2524 ( .A1(n3381), .A2(n2885), .ZN(n2351) );
  NAND2_X1 U2525 ( .A1(n2338), .A2(n2337), .ZN(n2336) );
  INV_X1 U2526 ( .A(n2340), .ZN(n2338) );
  INV_X1 U2527 ( .A(n2345), .ZN(n2337) );
  XNOR2_X1 U2528 ( .A(n3907), .B(n2279), .ZN(n4445) );
  NAND2_X1 U2529 ( .A1(n4454), .A2(n4455), .ZN(n4453) );
  XNOR2_X1 U2530 ( .A(n3910), .B(n2281), .ZN(n4466) );
  NAND2_X1 U2531 ( .A1(n4475), .A2(n4476), .ZN(n4474) );
  XNOR2_X1 U2532 ( .A(n3913), .B(n2280), .ZN(n4487) );
  OAI22_X1 U2533 ( .A1(n4498), .A2(n4495), .B1(n3915), .B2(
        REG2_REG_13__SCAN_IN), .ZN(n3916) );
  NOR2_X1 U2534 ( .A1(n2407), .A2(n2405), .ZN(n2404) );
  NAND2_X1 U2535 ( .A1(n2268), .A2(n2267), .ZN(n4076) );
  OR2_X1 U2536 ( .A1(n2270), .A2(n3651), .ZN(n2267) );
  NAND2_X1 U2537 ( .A1(n4094), .A2(n2269), .ZN(n2268) );
  NAND2_X1 U2538 ( .A1(n2270), .A2(n3651), .ZN(n2269) );
  NAND2_X1 U2539 ( .A1(n4187), .A2(n2637), .ZN(n2426) );
  AND2_X1 U2540 ( .A1(n3662), .A2(n2636), .ZN(n2637) );
  NOR2_X1 U2541 ( .A1(n2533), .A2(n2400), .ZN(n2399) );
  INV_X1 U2542 ( .A(n2523), .ZN(n2400) );
  NAND2_X1 U2543 ( .A1(n2924), .A2(n3659), .ZN(n2524) );
  AND2_X1 U2544 ( .A1(n4050), .A2(n2232), .ZN(n3969) );
  AND2_X1 U2545 ( .A1(n3476), .A2(n2366), .ZN(n2365) );
  NAND2_X1 U2546 ( .A1(n2371), .A2(n2368), .ZN(n2366) );
  INV_X1 U2547 ( .A(n2368), .ZN(n2367) );
  NAND2_X1 U2548 ( .A1(n4478), .A2(n4479), .ZN(n4477) );
  NOR2_X1 U2549 ( .A1(n3962), .A2(n3629), .ZN(n2304) );
  AND2_X1 U2550 ( .A1(n3503), .A2(n2358), .ZN(n2357) );
  NAND2_X1 U2551 ( .A1(n2359), .A2(n3596), .ZN(n2358) );
  INV_X1 U2552 ( .A(n3597), .ZN(n2359) );
  AOI21_X1 U2553 ( .B1(n3484), .B2(n3485), .A(n2247), .ZN(n2349) );
  NAND2_X1 U2554 ( .A1(n3011), .A2(n2849), .ZN(n2943) );
  AND2_X1 U2555 ( .A1(n4019), .A2(n3679), .ZN(n3998) );
  NAND2_X1 U2556 ( .A1(n2759), .A2(n3738), .ZN(n4221) );
  NAND2_X1 U2557 ( .A1(n3722), .A2(n3093), .ZN(n2299) );
  OR2_X1 U2558 ( .A1(n3796), .A2(n2961), .ZN(n3700) );
  AND2_X1 U2559 ( .A1(n2304), .A2(n2817), .ZN(n2303) );
  AND2_X1 U2560 ( .A1(n3179), .A2(n3254), .ZN(n2325) );
  INV_X1 U2561 ( .A(n2429), .ZN(n2427) );
  INV_X1 U2562 ( .A(IR_REG_21__SCAN_IN), .ZN(n2441) );
  NAND4_X1 U2563 ( .A1(n2575), .A2(n2437), .A3(n2436), .A4(n2435), .ZN(n2438)
         );
  OR2_X1 U2564 ( .A1(n2598), .A2(IR_REG_10__SCAN_IN), .ZN(n2599) );
  INV_X1 U2565 ( .A(IR_REG_4__SCAN_IN), .ZN(n4800) );
  INV_X1 U2566 ( .A(IR_REG_0__SCAN_IN), .ZN(n2388) );
  INV_X1 U2567 ( .A(n2375), .ZN(n2374) );
  OAI21_X1 U2568 ( .B1(n2369), .B2(n3541), .A(n2249), .ZN(n2368) );
  INV_X1 U2569 ( .A(n3605), .ZN(n2369) );
  AND2_X1 U2570 ( .A1(n2882), .A2(n2915), .ZN(n3431) );
  NAND2_X1 U2571 ( .A1(n2346), .A2(n4394), .ZN(n2345) );
  INV_X1 U2572 ( .A(n3342), .ZN(n2346) );
  NAND2_X1 U2573 ( .A1(n4394), .A2(n2348), .ZN(n2347) );
  AOI21_X1 U2574 ( .B1(n2349), .B2(n2342), .A(n2341), .ZN(n2340) );
  INV_X1 U2575 ( .A(n4392), .ZN(n2341) );
  INV_X1 U2576 ( .A(n3485), .ZN(n2342) );
  INV_X1 U2577 ( .A(n2349), .ZN(n2343) );
  NAND2_X1 U2578 ( .A1(n2464), .A2(n2463), .ZN(n2499) );
  NAND2_X1 U2579 ( .A1(n2462), .A2(n2442), .ZN(n2463) );
  NOR2_X1 U2580 ( .A1(n2865), .A2(n2864), .ZN(n2869) );
  OR2_X1 U2581 ( .A1(n2716), .A2(n2715), .ZN(n2722) );
  OR2_X1 U2582 ( .A1(n2702), .A2(n4977), .ZN(n2716) );
  INV_X1 U2583 ( .A(n2493), .ZN(n2471) );
  NAND2_X1 U2584 ( .A1(n2451), .A2(n2838), .ZN(n2290) );
  NAND2_X1 U2585 ( .A1(n4417), .A2(n3902), .ZN(n3904) );
  OR2_X1 U2586 ( .A1(n4424), .A2(n4425), .ZN(n2391) );
  OAI21_X1 U2587 ( .B1(n4641), .B2(n4435), .A(n2389), .ZN(n3871) );
  NAND2_X1 U2588 ( .A1(n2390), .A2(n4432), .ZN(n2389) );
  NAND2_X1 U2589 ( .A1(n4435), .A2(n4641), .ZN(n2390) );
  NAND2_X1 U2590 ( .A1(n4438), .A2(n3906), .ZN(n3907) );
  NAND2_X1 U2591 ( .A1(n4453), .A2(n3873), .ZN(n3874) );
  NAND2_X1 U2592 ( .A1(n4456), .A2(n3909), .ZN(n3910) );
  NAND2_X1 U2593 ( .A1(n4474), .A2(n2252), .ZN(n3876) );
  NAND2_X1 U2594 ( .A1(n4521), .A2(n3882), .ZN(n3884) );
  INV_X1 U2595 ( .A(n3636), .ZN(n2405) );
  AND2_X1 U2596 ( .A1(n3966), .A2(n3459), .ZN(n2409) );
  NOR2_X1 U2597 ( .A1(n2408), .A2(n2237), .ZN(n2407) );
  NOR3_X1 U2598 ( .A1(n2726), .A2(n2721), .A3(n2220), .ZN(n2408) );
  OR2_X1 U2599 ( .A1(n3964), .A2(n3988), .ZN(n2721) );
  AOI22_X1 U2600 ( .A1(n4017), .A2(n2708), .B1(n4044), .B2(n4027), .ZN(n3995)
         );
  INV_X1 U2601 ( .A(n4004), .ZN(n4044) );
  OR2_X1 U2602 ( .A1(n4101), .A2(n3518), .ZN(n2415) );
  NOR2_X1 U2603 ( .A1(n2414), .A2(n2412), .ZN(n2411) );
  INV_X1 U2604 ( .A(n2415), .ZN(n2412) );
  NAND2_X1 U2605 ( .A1(n4133), .A2(n2673), .ZN(n2674) );
  INV_X1 U2606 ( .A(n4155), .ZN(n2673) );
  AND2_X1 U2607 ( .A1(n4169), .A2(n2639), .ZN(n2425) );
  INV_X1 U2608 ( .A(n2263), .ZN(n2262) );
  OAI21_X1 U2609 ( .B1(n3656), .B2(n2264), .A(n2265), .ZN(n2263) );
  NAND2_X1 U2610 ( .A1(n2274), .A2(n2416), .ZN(n3206) );
  AOI21_X1 U2611 ( .B1(n2417), .B2(n2565), .A(n2222), .ZN(n2416) );
  NAND2_X1 U2612 ( .A1(n3062), .A2(n3716), .ZN(n2271) );
  NAND2_X1 U2613 ( .A1(n2257), .A2(n2256), .ZN(n3040) );
  OR2_X1 U2614 ( .A1(n2659), .A2(n4379), .ZN(n2257) );
  NAND2_X1 U2615 ( .A1(n2659), .A2(n4846), .ZN(n2256) );
  NAND2_X1 U2616 ( .A1(n3711), .A2(n3714), .ZN(n3659) );
  NAND2_X1 U2617 ( .A1(n2747), .A2(n3710), .ZN(n2925) );
  NAND2_X1 U2618 ( .A1(n2974), .A2(n2501), .ZN(n2899) );
  AND2_X1 U2619 ( .A1(n2850), .A2(n2798), .ZN(n2937) );
  AND2_X1 U2620 ( .A1(n4066), .A2(n4048), .ZN(n4050) );
  NAND2_X1 U2621 ( .A1(n2659), .A2(DATAI_23_), .ZN(n4048) );
  AND2_X1 U2622 ( .A1(n4084), .A2(n4068), .ZN(n4066) );
  NOR2_X1 U2623 ( .A1(n4109), .A2(n3518), .ZN(n4084) );
  INV_X1 U2624 ( .A(n3084), .ZN(n3081) );
  AND2_X1 U2625 ( .A1(n2937), .A2(n3774), .ZN(n4629) );
  NAND2_X1 U2626 ( .A1(n2794), .A2(n2795), .ZN(n3398) );
  NAND2_X1 U2627 ( .A1(n3011), .A2(n4588), .ZN(n3397) );
  INV_X1 U2628 ( .A(IR_REG_28__SCAN_IN), .ZN(n4801) );
  NAND2_X1 U2629 ( .A1(n2429), .A2(n2445), .ZN(n2428) );
  AND2_X1 U2630 ( .A1(n4919), .A2(n2442), .ZN(n2443) );
  NOR2_X1 U2631 ( .A1(n2427), .A2(n2322), .ZN(n2323) );
  NAND2_X1 U2632 ( .A1(n2457), .A2(n2670), .ZN(n2322) );
  NAND2_X1 U2633 ( .A1(n2459), .A2(n2458), .ZN(n2785) );
  NAND2_X1 U2634 ( .A1(n3324), .A2(n3323), .ZN(n3487) );
  INV_X1 U2635 ( .A(n3317), .ZN(n3318) );
  NAND2_X1 U2636 ( .A1(n3004), .A2(n3003), .ZN(n2332) );
  AND2_X1 U2637 ( .A1(n2363), .A2(n3454), .ZN(n2362) );
  INV_X1 U2638 ( .A(n3616), .ZN(n4396) );
  NAND4_X1 U2639 ( .A1(n2518), .A2(n2517), .A3(n2516), .A4(n2515), .ZN(n3792)
         );
  NAND2_X1 U2640 ( .A1(n4418), .A2(n4419), .ZN(n4417) );
  NOR2_X1 U2641 ( .A1(n4414), .A2(n4413), .ZN(n4412) );
  XNOR2_X1 U2642 ( .A(n3904), .B(n4598), .ZN(n4429) );
  NAND2_X1 U2643 ( .A1(n4439), .A2(n4440), .ZN(n4438) );
  NAND2_X1 U2644 ( .A1(n4457), .A2(n4458), .ZN(n4456) );
  XNOR2_X1 U2645 ( .A(n3876), .B(n2280), .ZN(n4492) );
  NAND2_X1 U2646 ( .A1(n4486), .A2(n3914), .ZN(n4498) );
  NAND2_X1 U2647 ( .A1(n4503), .A2(n4504), .ZN(n4502) );
  XNOR2_X1 U2648 ( .A(n3916), .B(n4592), .ZN(n4508) );
  NOR2_X1 U2649 ( .A1(n4508), .A2(n4509), .ZN(n4507) );
  NOR2_X1 U2650 ( .A1(n4531), .A2(REG1_REG_16__SCAN_IN), .ZN(n4532) );
  XNOR2_X1 U2651 ( .A(n3884), .B(n3883), .ZN(n4531) );
  AND2_X1 U2652 ( .A1(n4537), .A2(n2288), .ZN(n2287) );
  OR2_X1 U2653 ( .A1(n3922), .A2(REG2_REG_17__SCAN_IN), .ZN(n2288) );
  AND2_X1 U2654 ( .A1(n2287), .A2(n2286), .ZN(n3935) );
  AND2_X1 U2655 ( .A1(n4408), .A2(n3809), .ZN(n4542) );
  NAND2_X1 U2656 ( .A1(n4241), .A2(n2829), .ZN(n3954) );
  NAND2_X1 U2657 ( .A1(n2307), .A2(n2312), .ZN(n2308) );
  OR2_X1 U2658 ( .A1(n3954), .A2(n4371), .ZN(n2833) );
  OR2_X1 U2659 ( .A1(n2992), .A2(n2320), .ZN(n2319) );
  INV_X1 U2660 ( .A(n3714), .ZN(n2320) );
  INV_X1 U2661 ( .A(n2319), .ZN(n2318) );
  INV_X1 U2662 ( .A(IR_REG_9__SCAN_IN), .ZN(n4933) );
  INV_X1 U2663 ( .A(IR_REG_6__SCAN_IN), .ZN(n2574) );
  NOR2_X1 U2664 ( .A1(n3388), .A2(n2379), .ZN(n2378) );
  INV_X1 U2665 ( .A(n3587), .ZN(n2379) );
  NAND2_X1 U2666 ( .A1(n4078), .A2(n3755), .ZN(n2770) );
  NAND2_X1 U2667 ( .A1(n2291), .A2(n3754), .ZN(n4078) );
  OAI21_X1 U2668 ( .B1(n4152), .B2(n2292), .A(n3676), .ZN(n2291) );
  NAND2_X1 U2669 ( .A1(n4098), .A2(n2293), .ZN(n2292) );
  INV_X1 U2670 ( .A(n2553), .ZN(n2273) );
  NOR2_X1 U2671 ( .A1(n2418), .A2(n2579), .ZN(n2417) );
  INV_X1 U2672 ( .A(n2566), .ZN(n2418) );
  AND2_X1 U2673 ( .A1(n3710), .A2(n3707), .ZN(n2898) );
  NOR2_X1 U2674 ( .A1(n3998), .A2(n3762), .ZN(n3979) );
  AOI21_X1 U2675 ( .B1(n2303), .B2(n2771), .A(n2244), .ZN(n2301) );
  OR2_X1 U2676 ( .A1(n3685), .A2(n3687), .ZN(n2302) );
  AND2_X1 U2677 ( .A1(n2305), .A2(n3685), .ZN(n2818) );
  NOR2_X1 U2678 ( .A1(n4003), .A2(n3568), .ZN(n2328) );
  NAND2_X1 U2679 ( .A1(n2277), .A2(IR_REG_31__SCAN_IN), .ZN(n2461) );
  NAND2_X1 U2680 ( .A1(n2365), .A2(n2367), .ZN(n2363) );
  INV_X1 U2681 ( .A(n4086), .ZN(n3518) );
  NAND2_X1 U2682 ( .A1(n2696), .A2(REG3_REG_23__SCAN_IN), .ZN(n2702) );
  NAND2_X1 U2683 ( .A1(n2356), .A2(n2355), .ZN(n3584) );
  AOI21_X1 U2684 ( .B1(n2357), .B2(n2360), .A(n2227), .ZN(n2355) );
  NAND2_X1 U2685 ( .A1(n3298), .A2(n3277), .ZN(n2383) );
  NOR2_X1 U2686 ( .A1(n3390), .A2(n2376), .ZN(n2375) );
  INV_X1 U2687 ( .A(n3387), .ZN(n2376) );
  NAND2_X1 U2688 ( .A1(n3583), .A2(n2378), .ZN(n2377) );
  NOR2_X1 U2689 ( .A1(n2950), .A2(n2433), .ZN(n2951) );
  NAND2_X1 U2690 ( .A1(n2951), .A2(n2952), .ZN(n2333) );
  NAND2_X1 U2691 ( .A1(n3595), .A2(n3597), .ZN(n3594) );
  OR2_X1 U2692 ( .A1(n3487), .A2(n3484), .ZN(n2344) );
  NAND2_X1 U2693 ( .A1(n2339), .A2(n2349), .ZN(n4391) );
  NAND2_X1 U2694 ( .A1(n3487), .A2(n3485), .ZN(n2339) );
  AND2_X1 U2695 ( .A1(n2736), .A2(n2735), .ZN(n3479) );
  OR2_X1 U2696 ( .A1(n3469), .A2(n2493), .ZN(n2736) );
  OR2_X1 U2697 ( .A1(n2723), .A2(n2727), .ZN(n3478) );
  NAND2_X1 U2698 ( .A1(n2502), .A2(REG1_REG_1__SCAN_IN), .ZN(n2473) );
  OR2_X1 U2699 ( .A1(n2493), .A2(n2880), .ZN(n2486) );
  OR2_X1 U2700 ( .A1(n2492), .A2(n2484), .ZN(n2489) );
  XNOR2_X1 U2701 ( .A(n3857), .B(n3843), .ZN(n3856) );
  NAND2_X1 U2702 ( .A1(n4449), .A2(n3872), .ZN(n4454) );
  NAND2_X1 U2703 ( .A1(n4470), .A2(n3875), .ZN(n4475) );
  NAND2_X1 U2704 ( .A1(n4477), .A2(n3912), .ZN(n3913) );
  NAND2_X1 U2705 ( .A1(n4502), .A2(n3878), .ZN(n3880) );
  NOR2_X1 U2706 ( .A1(n4516), .A2(n2282), .ZN(n3920) );
  AND2_X1 U2707 ( .A1(n3919), .A2(REG2_REG_15__SCAN_IN), .ZN(n2282) );
  NAND2_X1 U2708 ( .A1(n2499), .A2(n2845), .ZN(n3797) );
  NOR2_X1 U2709 ( .A1(n2722), .A2(n4957), .ZN(n2727) );
  INV_X1 U2710 ( .A(n2305), .ZN(n3961) );
  NAND2_X1 U2711 ( .A1(n2306), .A2(n3766), .ZN(n3963) );
  INV_X1 U2712 ( .A(n4010), .ZN(n4003) );
  NAND2_X1 U2713 ( .A1(n2266), .A2(n2410), .ZN(n4037) );
  AOI21_X1 U2714 ( .B1(n2411), .B2(n2694), .A(n2223), .ZN(n2410) );
  NAND2_X1 U2715 ( .A1(n4076), .A2(n2411), .ZN(n2266) );
  NOR2_X1 U2716 ( .A1(n2687), .A2(n3516), .ZN(n2688) );
  AND2_X1 U2717 ( .A1(n3653), .A2(n4038), .ZN(n4075) );
  INV_X1 U2718 ( .A(REG3_REG_20__SCAN_IN), .ZN(n4777) );
  OR2_X1 U2719 ( .A1(n2677), .A2(n4777), .ZN(n2687) );
  NAND2_X1 U2720 ( .A1(n2675), .A2(REG3_REG_19__SCAN_IN), .ZN(n2677) );
  AOI21_X1 U2721 ( .B1(n4150), .B2(n2661), .A(n2434), .ZN(n4144) );
  AND2_X1 U2722 ( .A1(n2663), .A2(REG3_REG_18__SCAN_IN), .ZN(n2675) );
  NAND2_X1 U2723 ( .A1(n4179), .A2(n2650), .ZN(n4150) );
  OR2_X1 U2724 ( .A1(n4159), .A2(n4386), .ZN(n2650) );
  NOR2_X1 U2725 ( .A1(n2622), .A2(n4744), .ZN(n2630) );
  INV_X1 U2726 ( .A(REG3_REG_14__SCAN_IN), .ZN(n4744) );
  NAND2_X1 U2727 ( .A1(n2248), .A2(n2601), .ZN(n2264) );
  INV_X1 U2728 ( .A(REG3_REG_12__SCAN_IN), .ZN(n4955) );
  OR2_X1 U2729 ( .A1(n2603), .A2(n4955), .ZN(n2614) );
  OAI21_X1 U2730 ( .B1(n3094), .B2(n2298), .A(n2294), .ZN(n3177) );
  AOI21_X1 U2731 ( .B1(n2297), .B2(n2296), .A(n2295), .ZN(n2294) );
  INV_X1 U2732 ( .A(n3722), .ZN(n2296) );
  AND2_X1 U2733 ( .A1(n2580), .A2(REG3_REG_10__SCAN_IN), .ZN(n2592) );
  INV_X1 U2734 ( .A(REG3_REG_9__SCAN_IN), .ZN(n2567) );
  OR2_X1 U2735 ( .A1(n2554), .A2(n4958), .ZN(n2568) );
  NAND2_X1 U2736 ( .A1(n2749), .A2(n3717), .ZN(n3057) );
  INV_X1 U2737 ( .A(REG3_REG_6__SCAN_IN), .ZN(n3073) );
  NAND2_X1 U2738 ( .A1(n2321), .A2(n3714), .ZN(n2996) );
  OR2_X1 U2739 ( .A1(n2925), .A2(n2748), .ZN(n2321) );
  AND2_X1 U2740 ( .A1(REG3_REG_3__SCAN_IN), .A2(REG3_REG_4__SCAN_IN), .ZN(
        n2526) );
  NAND2_X1 U2741 ( .A1(n2746), .A2(n3705), .ZN(n2900) );
  NAND2_X1 U2742 ( .A1(n2289), .A2(n2745), .ZN(n2746) );
  INV_X1 U2743 ( .A(n4158), .ZN(n4219) );
  INV_X1 U2744 ( .A(n2898), .ZN(n3661) );
  OAI21_X1 U2745 ( .B1(n3700), .B2(n2743), .A(n2744), .ZN(n2289) );
  OAI21_X1 U2746 ( .B1(n2499), .B2(n2482), .A(n2481), .ZN(n2965) );
  NAND2_X1 U2747 ( .A1(n2499), .A2(n2480), .ZN(n2481) );
  NAND2_X1 U2748 ( .A1(n2742), .A2(n3941), .ZN(n4227) );
  INV_X1 U2749 ( .A(n4216), .ZN(n4194) );
  OR2_X1 U2750 ( .A1(n2853), .A2(n2851), .ZN(n2908) );
  INV_X1 U2751 ( .A(n3691), .ZN(n2827) );
  OR2_X1 U2752 ( .A1(n2828), .A2(n2827), .ZN(n4241) );
  NOR2_X1 U2753 ( .A1(n4241), .A2(n4245), .ZN(n4240) );
  INV_X1 U2754 ( .A(n3689), .ZN(n4245) );
  NAND2_X1 U2755 ( .A1(n2499), .A2(DATAI_28_), .ZN(n3447) );
  NAND2_X1 U2756 ( .A1(n2659), .A2(DATAI_25_), .ZN(n4010) );
  NAND2_X1 U2757 ( .A1(n4050), .A2(n2328), .ZN(n4009) );
  NAND2_X1 U2758 ( .A1(n4050), .A2(n4027), .ZN(n4029) );
  NAND2_X1 U2759 ( .A1(n2659), .A2(DATAI_21_), .ZN(n4086) );
  OR2_X1 U2760 ( .A1(n2225), .A2(n4107), .ZN(n4109) );
  INV_X1 U2761 ( .A(n3506), .ZN(n4126) );
  NOR3_X1 U2762 ( .A1(n4201), .A2(n3558), .A3(n4176), .ZN(n4160) );
  NOR2_X1 U2763 ( .A1(n4201), .A2(n4176), .ZN(n4178) );
  OR2_X1 U2764 ( .A1(n4228), .A2(n3620), .ZN(n4201) );
  AND2_X1 U2765 ( .A1(n3205), .A2(n2250), .ZN(n4230) );
  INV_X1 U2766 ( .A(n3269), .ZN(n3254) );
  NAND2_X1 U2767 ( .A1(n3205), .A2(n3254), .ZN(n3204) );
  NOR2_X1 U2768 ( .A1(n3113), .A2(n3197), .ZN(n3205) );
  AND2_X1 U2769 ( .A1(n3128), .A2(n3081), .ZN(n2327) );
  OR2_X1 U2770 ( .A1(n3112), .A2(n3156), .ZN(n3113) );
  NAND2_X1 U2771 ( .A1(n2255), .A2(n2226), .ZN(n3080) );
  NAND2_X1 U2772 ( .A1(n2930), .A2(n3040), .ZN(n2994) );
  INV_X1 U2773 ( .A(n3019), .ZN(n2904) );
  AND2_X1 U2774 ( .A1(n2976), .A2(n2904), .ZN(n2930) );
  NAND2_X1 U2775 ( .A1(n4227), .A2(n4624), .ZN(n4622) );
  INV_X1 U2776 ( .A(n2428), .ZN(n2314) );
  NOR2_X1 U2777 ( .A1(n2427), .A2(IR_REG_18__SCAN_IN), .ZN(n2324) );
  INV_X1 U2778 ( .A(IR_REG_23__SCAN_IN), .ZN(n2797) );
  XNOR2_X1 U2779 ( .A(n2796), .B(n2797), .ZN(n3010) );
  XNOR2_X1 U2780 ( .A(n2737), .B(n4721), .ZN(n2850) );
  XNOR2_X1 U2781 ( .A(n2741), .B(n2441), .ZN(n2798) );
  NAND2_X1 U2782 ( .A1(n2682), .A2(IR_REG_31__SCAN_IN), .ZN(n2684) );
  NOR2_X1 U2783 ( .A1(n2477), .A2(n2459), .ZN(n2387) );
  NAND2_X1 U2784 ( .A1(n2479), .A2(n2478), .ZN(n3804) );
  NAND2_X1 U2785 ( .A1(n2364), .A2(n2368), .ZN(n3477) );
  NAND2_X1 U2786 ( .A1(n3594), .A2(n3596), .ZN(n3504) );
  NAND2_X1 U2787 ( .A1(n3583), .A2(n3587), .ZN(n3515) );
  NAND2_X1 U2788 ( .A1(n2335), .A2(n2334), .ZN(n3345) );
  AOI22_X1 U2789 ( .A1(n2340), .A2(n2343), .B1(n2345), .B2(n2347), .ZN(n2334)
         );
  OAI21_X1 U2790 ( .B1(n2499), .B2(n2395), .A(n2490), .ZN(n2862) );
  NAND2_X1 U2791 ( .A1(n2499), .A2(DATAI_0_), .ZN(n2490) );
  NAND2_X1 U2792 ( .A1(n2377), .A2(n3387), .ZN(n3389) );
  INV_X1 U2793 ( .A(n2984), .ZN(n2977) );
  OR2_X1 U2794 ( .A1(n2892), .A2(n2891), .ZN(n4384) );
  NAND2_X1 U2795 ( .A1(n2873), .A2(n2872), .ZN(n3616) );
  OR3_X1 U2796 ( .A1(n2707), .A2(n2706), .A3(n2705), .ZN(n4004) );
  OR2_X1 U2797 ( .A1(n2492), .A2(n4612), .ZN(n2495) );
  NAND2_X1 U2798 ( .A1(n2502), .A2(REG1_REG_2__SCAN_IN), .ZN(n2497) );
  CLKBUF_X1 U2799 ( .A(n2861), .Z(n3796) );
  NAND2_X1 U2800 ( .A1(n3803), .A2(n3810), .ZN(n3826) );
  NAND2_X1 U2801 ( .A1(n3855), .A2(REG1_REG_4__SCAN_IN), .ZN(n3867) );
  OAI22_X1 U2802 ( .A1(n3901), .A2(n3900), .B1(n3899), .B2(n3898), .ZN(n4418)
         );
  AND2_X1 U2803 ( .A1(n3867), .A2(n2386), .ZN(n4414) );
  NAND2_X1 U2804 ( .A1(n3868), .A2(n4379), .ZN(n2386) );
  INV_X1 U2805 ( .A(n2391), .ZN(n4423) );
  NAND2_X1 U2806 ( .A1(n4428), .A2(n3905), .ZN(n4439) );
  AND2_X1 U2807 ( .A1(n2391), .A2(n2245), .ZN(n4435) );
  XNOR2_X1 U2808 ( .A(n3871), .B(n2279), .ZN(n4450) );
  NAND2_X1 U2809 ( .A1(n4444), .A2(n3908), .ZN(n4457) );
  XNOR2_X1 U2810 ( .A(n3874), .B(n2281), .ZN(n4471) );
  NAND2_X1 U2811 ( .A1(n4465), .A2(n3911), .ZN(n4478) );
  NAND2_X1 U2812 ( .A1(n4491), .A2(n3877), .ZN(n4503) );
  XNOR2_X1 U2813 ( .A(n3880), .B(n4592), .ZN(n4513) );
  NOR2_X1 U2814 ( .A1(n3917), .A2(n4507), .ZN(n4518) );
  NOR2_X1 U2815 ( .A1(n4518), .A2(n4517), .ZN(n4516) );
  XNOR2_X1 U2816 ( .A(n3920), .B(n3883), .ZN(n4528) );
  NAND2_X1 U2817 ( .A1(n4528), .A2(n4526), .ZN(n4527) );
  NOR2_X1 U2818 ( .A1(n4532), .A2(n3885), .ZN(n4544) );
  INV_X1 U2819 ( .A(n3923), .ZN(n2286) );
  AOI21_X1 U2820 ( .B1(REG2_REG_18__SCAN_IN), .B2(n4378), .A(n3935), .ZN(n3938) );
  XNOR2_X1 U2821 ( .A(n2402), .B(n2278), .ZN(n3952) );
  OAI21_X1 U2822 ( .B1(n3977), .B2(n2243), .A(n2403), .ZN(n2402) );
  NOR2_X1 U2823 ( .A1(n2404), .A2(n2409), .ZN(n2403) );
  INV_X1 U2824 ( .A(n2406), .ZN(n3960) );
  NAND2_X1 U2825 ( .A1(n2413), .A2(n2415), .ZN(n4057) );
  OR2_X1 U2826 ( .A1(n4076), .A2(n2694), .ZN(n2413) );
  NAND2_X1 U2827 ( .A1(n2426), .A2(n2639), .ZN(n4181) );
  NAND2_X1 U2828 ( .A1(n2261), .A2(n2601), .ZN(n3170) );
  NAND2_X1 U2829 ( .A1(n3176), .A2(n3656), .ZN(n2261) );
  NAND2_X1 U2830 ( .A1(n2419), .A2(n2566), .ZN(n3098) );
  OR2_X1 U2831 ( .A1(n3116), .A2(n2565), .ZN(n2419) );
  NAND2_X1 U2832 ( .A1(n2396), .A2(n2397), .ZN(n3082) );
  INV_X1 U2833 ( .A(n4204), .ZN(n4569) );
  NAND2_X1 U2834 ( .A1(n2524), .A2(n2523), .ZN(n2993) );
  OR2_X1 U2835 ( .A1(n3397), .A2(n2876), .ZN(n4231) );
  INV_X1 U2836 ( .A(n4231), .ZN(n4565) );
  OR2_X1 U2837 ( .A1(n4050), .A2(n4049), .ZN(n4336) );
  OR2_X1 U2838 ( .A1(n2826), .A2(n2848), .ZN(n4630) );
  NAND2_X1 U2839 ( .A1(n2835), .A2(IR_REG_31__SCAN_IN), .ZN(n2392) );
  NOR2_X1 U2840 ( .A1(n2682), .A2(n2428), .ZN(n2774) );
  NAND2_X1 U2841 ( .A1(n2792), .A2(IR_REG_31__SCAN_IN), .ZN(n2793) );
  AOI21_X1 U2842 ( .B1(n2787), .B2(IR_REG_25__SCAN_IN), .A(n2786), .ZN(n3401)
         );
  AND2_X1 U2843 ( .A1(n2669), .A2(n2323), .ZN(n2784) );
  AND2_X1 U2844 ( .A1(n3010), .A2(STATE_REG_SCAN_IN), .ZN(n4588) );
  INV_X1 U2845 ( .A(n2850), .ZN(n4375) );
  INV_X1 U2846 ( .A(DATAI_16_), .ZN(n4989) );
  INV_X1 U2847 ( .A(n3891), .ZN(n4595) );
  INV_X2 U2848 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  OAI21_X1 U2849 ( .B1(n3545), .B2(n2367), .A(n2365), .ZN(n3467) );
  OAI21_X1 U2850 ( .B1(n2287), .B2(n2286), .A(n4496), .ZN(n2285) );
  AOI21_X1 U2851 ( .B1(n3929), .B2(n4542), .A(n3928), .ZN(n2284) );
  NAND2_X1 U2852 ( .A1(n2276), .A2(n2275), .ZN(U3515) );
  AND2_X1 U2853 ( .A1(n2833), .A2(n2253), .ZN(n2275) );
  NAND2_X1 U2854 ( .A1(n2308), .A2(n4631), .ZN(n2276) );
  OR2_X1 U2855 ( .A1(n4251), .A2(n4371), .ZN(n2814) );
  INV_X1 U2856 ( .A(n3534), .ZN(n3296) );
  NOR2_X1 U2857 ( .A1(n2385), .A2(n2384), .ZN(n3299) );
  AND2_X1 U2858 ( .A1(n3964), .A2(n3988), .ZN(n2220) );
  INV_X1 U2859 ( .A(n4081), .ZN(n3316) );
  NOR2_X1 U2860 ( .A1(n2398), .A2(n2543), .ZN(n2221) );
  NOR2_X1 U2861 ( .A1(n3208), .A2(n3196), .ZN(n2222) );
  AND2_X1 U2862 ( .A1(n4081), .A2(n2695), .ZN(n2223) );
  AND2_X1 U2863 ( .A1(n2669), .A2(n2324), .ZN(n2224) );
  INV_X1 U2864 ( .A(n4122), .ZN(n2270) );
  OR3_X1 U2865 ( .A1(n4201), .A2(n2331), .A3(n3506), .ZN(n2225) );
  AND2_X1 U2866 ( .A1(n3051), .A2(n3040), .ZN(n2226) );
  AND2_X1 U2867 ( .A1(n3371), .A2(n3370), .ZN(n2227) );
  AND2_X1 U2868 ( .A1(n2325), .A2(n3296), .ZN(n2228) );
  AND2_X1 U2869 ( .A1(n3205), .A2(n2325), .ZN(n2229) );
  AND2_X1 U2870 ( .A1(n2328), .A2(n3988), .ZN(n2230) );
  OR2_X1 U2871 ( .A1(n4646), .A2(REG1_REG_29__SCAN_IN), .ZN(n2231) );
  AND2_X1 U2872 ( .A1(n2230), .A2(n3971), .ZN(n2232) );
  INV_X1 U2873 ( .A(n4386), .ZN(n4176) );
  OAI211_X1 U2875 ( .C1(n2779), .C2(n2720), .A(n2719), .B(n2718), .ZN(n4002)
         );
  NAND2_X1 U2876 ( .A1(n2344), .A2(n3342), .ZN(n3618) );
  NAND2_X1 U2877 ( .A1(n2451), .A2(n2452), .ZN(n2492) );
  AND2_X1 U2878 ( .A1(n2377), .A2(n2375), .ZN(n2233) );
  INV_X1 U2879 ( .A(IR_REG_18__SCAN_IN), .ZN(n2670) );
  NAND2_X2 U2880 ( .A1(n4373), .A2(n2838), .ZN(n2493) );
  AOI22_X1 U2881 ( .A1(n3995), .A2(n2714), .B1(n4003), .B2(n4024), .ZN(n3977)
         );
  XNOR2_X1 U2882 ( .A(n2392), .B(IR_REG_30__SCAN_IN), .ZN(n4373) );
  OAI21_X1 U2883 ( .B1(n4037), .B2(n3637), .A(n3638), .ZN(n4017) );
  OR2_X1 U2884 ( .A1(n2726), .A2(n2220), .ZN(n2234) );
  INV_X1 U2885 ( .A(IR_REG_2__SCAN_IN), .ZN(n2498) );
  OR2_X1 U2886 ( .A1(n3045), .A2(n3044), .ZN(n2235) );
  AND2_X1 U2887 ( .A1(n2646), .A2(n4896), .ZN(n2236) );
  NOR2_X1 U2888 ( .A1(n3611), .A2(n3971), .ZN(n2237) );
  AND2_X1 U2889 ( .A1(n2413), .A2(n2411), .ZN(n2238) );
  INV_X1 U2890 ( .A(IR_REG_25__SCAN_IN), .ZN(n2458) );
  AND2_X1 U2891 ( .A1(n2417), .A2(n2272), .ZN(n2239) );
  AND2_X1 U2892 ( .A1(n3411), .A2(n2372), .ZN(n2240) );
  OR2_X1 U2893 ( .A1(n2682), .A2(n2430), .ZN(n2241) );
  OR2_X1 U2894 ( .A1(n2682), .A2(n2440), .ZN(n2242) );
  OR2_X1 U2895 ( .A1(n3040), .A2(n3792), .ZN(n3711) );
  INV_X1 U2896 ( .A(IR_REG_22__SCAN_IN), .ZN(n4721) );
  INV_X1 U2897 ( .A(n2298), .ZN(n2297) );
  NAND2_X1 U2898 ( .A1(n2299), .A2(n3736), .ZN(n2298) );
  OR2_X1 U2899 ( .A1(n2234), .A2(n2405), .ZN(n2243) );
  NAND2_X1 U2900 ( .A1(n2302), .A2(n3686), .ZN(n2244) );
  NOR2_X1 U2901 ( .A1(IR_REG_24__SCAN_IN), .A2(IR_REG_23__SCAN_IN), .ZN(n2457)
         );
  OR2_X1 U2902 ( .A1(n3870), .A2(n4598), .ZN(n2245) );
  INV_X1 U2903 ( .A(n2398), .ZN(n2397) );
  NOR2_X1 U2904 ( .A1(n3047), .A2(n3791), .ZN(n2398) );
  OAI21_X1 U2905 ( .B1(n2285), .B2(n3935), .A(n2284), .ZN(U3258) );
  AND2_X1 U2906 ( .A1(n3745), .A2(n3747), .ZN(n4180) );
  INV_X1 U2907 ( .A(n3321), .ZN(n2381) );
  INV_X1 U2908 ( .A(n3669), .ZN(n2278) );
  AND2_X1 U2909 ( .A1(n4103), .A2(n4126), .ZN(n2246) );
  AOI21_X1 U2910 ( .B1(n3153), .B2(n3152), .A(n3151), .ZN(n3190) );
  XNOR2_X1 U2911 ( .A(n3332), .B(n3331), .ZN(n2247) );
  AOI21_X1 U2912 ( .B1(n4116), .B2(n2686), .A(n2246), .ZN(n4094) );
  INV_X1 U2913 ( .A(n4058), .ZN(n2414) );
  INV_X1 U2914 ( .A(n4432), .ZN(n4597) );
  OR2_X1 U2915 ( .A1(n3784), .A2(n3534), .ZN(n2248) );
  INV_X1 U2916 ( .A(n4096), .ZN(n2293) );
  NAND2_X1 U2917 ( .A1(n2426), .A2(n2425), .ZN(n4179) );
  NAND2_X1 U2918 ( .A1(n2620), .A2(n2439), .ZN(n2628) );
  NAND2_X1 U2919 ( .A1(n4050), .A2(n2230), .ZN(n2329) );
  INV_X1 U2920 ( .A(n3277), .ZN(n2384) );
  NAND2_X1 U2921 ( .A1(n3437), .A2(n3436), .ZN(n2249) );
  INV_X1 U2922 ( .A(n2311), .ZN(n2310) );
  OAI21_X1 U2923 ( .B1(n3479), .B2(n4158), .A(n2825), .ZN(n2311) );
  INV_X2 U2924 ( .A(IR_REG_0__SCAN_IN), .ZN(n2395) );
  INV_X1 U2925 ( .A(n2371), .ZN(n2370) );
  NAND2_X1 U2926 ( .A1(n2249), .A2(n3542), .ZN(n2371) );
  INV_X1 U2927 ( .A(n3128), .ZN(n3133) );
  INV_X1 U2928 ( .A(n3179), .ZN(n3286) );
  AND2_X1 U2929 ( .A1(n2228), .A2(n3229), .ZN(n2250) );
  NAND2_X1 U2930 ( .A1(n2620), .A2(n2423), .ZN(n2251) );
  INV_X1 U2931 ( .A(IR_REG_26__SCAN_IN), .ZN(n4919) );
  INV_X1 U2932 ( .A(n3484), .ZN(n2348) );
  XNOR2_X1 U2933 ( .A(n2793), .B(IR_REG_26__SCAN_IN), .ZN(n2795) );
  INV_X1 U2934 ( .A(n3596), .ZN(n2360) );
  NAND2_X1 U2935 ( .A1(n2271), .A2(n2553), .ZN(n3116) );
  NAND2_X1 U2936 ( .A1(n2659), .A2(DATAI_24_), .ZN(n4027) );
  NAND2_X1 U2937 ( .A1(n2659), .A2(DATAI_22_), .ZN(n4068) );
  INV_X1 U2938 ( .A(n3733), .ZN(n2295) );
  NAND2_X1 U2939 ( .A1(n2620), .A2(n2422), .ZN(n2657) );
  INV_X1 U2940 ( .A(n3651), .ZN(n4107) );
  NAND2_X1 U2941 ( .A1(n2659), .A2(DATAI_20_), .ZN(n3651) );
  INV_X1 U2942 ( .A(n2330), .ZN(n4132) );
  NOR2_X1 U2943 ( .A1(n4201), .A2(n2331), .ZN(n2330) );
  OR2_X1 U2944 ( .A1(n4595), .A2(n4644), .ZN(n2252) );
  NAND2_X1 U2945 ( .A1(n3205), .A2(n2228), .ZN(n2326) );
  CLKBUF_X1 U2946 ( .A(n2885), .Z(n2887) );
  INV_X1 U2947 ( .A(n3883), .ZN(n4590) );
  INV_X2 U2948 ( .A(n4643), .ZN(n4646) );
  OR2_X1 U2949 ( .A1(n4631), .A2(n2832), .ZN(n2253) );
  AND2_X1 U2950 ( .A1(n4408), .A2(n3811), .ZN(n4496) );
  AND2_X1 U2951 ( .A1(n2930), .A2(n2226), .ZN(n2254) );
  INV_X1 U2952 ( .A(n3988), .ZN(n3428) );
  NAND2_X1 U2953 ( .A1(n2499), .A2(DATAI_26_), .ZN(n3988) );
  AND2_X1 U2954 ( .A1(n2930), .A2(n3081), .ZN(n2255) );
  INV_X1 U2955 ( .A(IR_REG_15__SCAN_IN), .ZN(n2646) );
  INV_X1 U2956 ( .A(n4485), .ZN(n2280) );
  INV_X1 U2957 ( .A(n4443), .ZN(n2279) );
  INV_X1 U2958 ( .A(n4464), .ZN(n2281) );
  INV_X1 U2959 ( .A(IR_REG_29__SCAN_IN), .ZN(n2446) );
  INV_X1 U2960 ( .A(IR_REG_20__SCAN_IN), .ZN(n2739) );
  INV_X1 U2961 ( .A(IR_REG_14__SCAN_IN), .ZN(n2424) );
  INV_X1 U2962 ( .A(IR_REG_1__SCAN_IN), .ZN(n2394) );
  INV_X1 U2963 ( .A(IR_REG_17__SCAN_IN), .ZN(n2421) );
  OAI21_X1 U2964 ( .B1(n3176), .B2(n2264), .A(n2262), .ZN(n3228) );
  NAND2_X1 U2965 ( .A1(n3176), .A2(n2262), .ZN(n2260) );
  OR2_X1 U2966 ( .A1(n3296), .A2(n3180), .ZN(n2265) );
  NAND3_X1 U2967 ( .A1(n2669), .A2(n2323), .A3(n2458), .ZN(n2792) );
  NAND4_X1 U2968 ( .A1(n2669), .A2(n2323), .A3(n2458), .A4(n4919), .ZN(n2277)
         );
  INV_X1 U2969 ( .A(n2461), .ZN(n2824) );
  XNOR2_X1 U2970 ( .A(n2289), .B(n3660), .ZN(n2988) );
  OAI21_X1 U2971 ( .B1(n3094), .B2(n3093), .A(n3722), .ZN(n3207) );
  OR2_X1 U2972 ( .A1(n3979), .A2(n2771), .ZN(n2306) );
  NAND2_X1 U2973 ( .A1(n2300), .A2(n2301), .ZN(n2819) );
  NAND2_X1 U2974 ( .A1(n3979), .A2(n2303), .ZN(n2300) );
  NAND2_X1 U2975 ( .A1(n2306), .A2(n2304), .ZN(n2305) );
  NAND2_X1 U2976 ( .A1(n2820), .A2(n4223), .ZN(n2312) );
  NAND2_X1 U2977 ( .A1(n2312), .A2(n2310), .ZN(n3956) );
  OAI21_X1 U2978 ( .B1(n2308), .B2(n4643), .A(n2231), .ZN(n2831) );
  NAND2_X1 U2979 ( .A1(n2314), .A2(n2313), .ZN(n2448) );
  NAND3_X1 U2980 ( .A1(n2420), .A2(n2620), .A3(n2670), .ZN(n2682) );
  NAND2_X1 U2981 ( .A1(n2925), .A2(n2318), .ZN(n2317) );
  NAND2_X1 U2982 ( .A1(n2763), .A2(n3747), .ZN(n4152) );
  NAND4_X1 U2983 ( .A1(n2489), .A2(n2488), .A3(n2487), .A4(n2486), .ZN(n2861)
         );
  MUX2_X1 U2984 ( .A(n4380), .B(DATAI_3_), .S(n2499), .Z(n3019) );
  INV_X1 U2985 ( .A(n2326), .ZN(n3230) );
  NAND3_X1 U2986 ( .A1(n2226), .A2(n2930), .A3(n2327), .ZN(n3112) );
  INV_X1 U2987 ( .A(n2329), .ZN(n3987) );
  NAND3_X1 U2988 ( .A1(n4162), .A2(n4133), .A3(n4386), .ZN(n2331) );
  OAI21_X1 U2989 ( .B1(n2951), .B2(n2952), .A(n2333), .ZN(n2953) );
  NAND2_X1 U2990 ( .A1(n3487), .A2(n2336), .ZN(n2335) );
  INV_X1 U2991 ( .A(n2965), .ZN(n2895) );
  XNOR2_X1 U2992 ( .A(n2350), .B(n3431), .ZN(n2946) );
  INV_X4 U2993 ( .A(n2943), .ZN(n3381) );
  NAND2_X1 U2994 ( .A1(n2354), .A2(n2353), .ZN(n3153) );
  NAND2_X1 U2995 ( .A1(n3132), .A2(n3131), .ZN(n2353) );
  NAND2_X1 U2996 ( .A1(n3069), .A2(n3068), .ZN(n3132) );
  NAND2_X1 U2997 ( .A1(n3595), .A2(n2357), .ZN(n2356) );
  NAND2_X1 U2998 ( .A1(n2361), .A2(n2362), .ZN(n3465) );
  NAND2_X1 U2999 ( .A1(n3545), .A2(n2365), .ZN(n2361) );
  NAND2_X1 U3000 ( .A1(n3545), .A2(n2370), .ZN(n2364) );
  AOI21_X1 U3001 ( .B1(n3545), .B2(n3542), .A(n3541), .ZN(n3607) );
  OAI21_X2 U3002 ( .B1(n3583), .B2(n2374), .A(n2240), .ZN(n3496) );
  INV_X1 U3003 ( .A(n3278), .ZN(n2385) );
  OAI21_X2 U3004 ( .B1(n2385), .B2(n2383), .A(n3305), .ZN(n3320) );
  XNOR2_X2 U3005 ( .A(n2387), .B(IR_REG_2__SCAN_IN), .ZN(n3836) );
  NAND3_X1 U3006 ( .A1(n2395), .A2(n2498), .A3(n2394), .ZN(n2508) );
  NAND4_X1 U3007 ( .A1(n2393), .A2(n2519), .A3(n2498), .A4(n2395), .ZN(n2531)
         );
  NAND2_X1 U3008 ( .A1(n2524), .A2(n2399), .ZN(n2396) );
  OAI21_X1 U3009 ( .B1(n3977), .B2(n2234), .A(n2407), .ZN(n2816) );
  AOI21_X1 U3010 ( .B1(n3977), .B2(n2721), .A(n2220), .ZN(n2406) );
  OR2_X1 U3011 ( .A1(n2224), .A2(n2459), .ZN(n2796) );
  AND2_X1 U3012 ( .A1(n2861), .A2(n3381), .ZN(n2865) );
  XNOR2_X1 U3013 ( .A(n3004), .B(n2945), .ZN(n2952) );
  NAND2_X1 U3014 ( .A1(n3322), .A2(n2381), .ZN(n3323) );
  NAND3_X2 U3015 ( .A1(n2795), .A2(n3401), .A3(n4374), .ZN(n3011) );
  INV_X1 U3016 ( .A(n2866), .ZN(n2870) );
  NAND2_X1 U3017 ( .A1(n2448), .A2(IR_REG_31__SCAN_IN), .ZN(n2449) );
  NAND2_X1 U3018 ( .A1(n2885), .A2(n2965), .ZN(n3701) );
  AOI22_X1 U3019 ( .A1(n3036), .A2(n3035), .B1(n3034), .B2(n3033), .ZN(n3576)
         );
  NAND2_X2 U3020 ( .A1(n2914), .A2(n4231), .ZN(n4207) );
  NAND2_X1 U3021 ( .A1(n3399), .A2(n3398), .ZN(n4575) );
  INV_X2 U3022 ( .A(n4575), .ZN(n4587) );
  NOR3_X1 U3023 ( .A1(n3448), .A2(n2882), .A3(n3400), .ZN(n2432) );
  INV_X1 U3024 ( .A(n3804), .ZN(n2482) );
  AND2_X1 U3025 ( .A1(n2949), .A2(n2948), .ZN(n2433) );
  AND2_X1 U3026 ( .A1(n3558), .A2(n4389), .ZN(n2434) );
  INV_X1 U3027 ( .A(n3401), .ZN(n2788) );
  AOI22_X1 U3028 ( .A1(n3282), .A2(n3794), .B1(n2977), .B2(n3381), .ZN(n3003)
         );
  AND2_X1 U3029 ( .A1(n4186), .A2(n2638), .ZN(n2636) );
  INV_X1 U3030 ( .A(n3267), .ZN(n3264) );
  INV_X1 U3031 ( .A(IR_REG_13__SCAN_IN), .ZN(n2439) );
  INV_X1 U3032 ( .A(n3320), .ZN(n3322) );
  INV_X1 U3033 ( .A(REG3_REG_24__SCAN_IN), .ZN(n4977) );
  AOI22_X1 U3034 ( .A1(n3381), .A2(n2862), .B1(IR_REG_0__SCAN_IN), .B2(n2858), 
        .ZN(n2859) );
  INV_X1 U3035 ( .A(REG3_REG_21__SCAN_IN), .ZN(n3516) );
  INV_X1 U3036 ( .A(REG3_REG_13__SCAN_IN), .ZN(n2613) );
  INV_X1 U3037 ( .A(n3259), .ZN(n3260) );
  INV_X1 U3038 ( .A(n3003), .ZN(n2945) );
  AND2_X1 U3039 ( .A1(n2688), .A2(REG3_REG_22__SCAN_IN), .ZN(n2696) );
  OR2_X1 U3040 ( .A1(n2614), .A2(n2613), .ZN(n2622) );
  INV_X1 U3041 ( .A(REG3_REG_8__SCAN_IN), .ZN(n4958) );
  AND2_X1 U3042 ( .A1(n2861), .A2(n2862), .ZN(n2960) );
  INV_X1 U3043 ( .A(REG3_REG_27__SCAN_IN), .ZN(n4957) );
  AOI21_X1 U3044 ( .B1(n3341), .B2(n3340), .A(n3343), .ZN(n4394) );
  INV_X1 U3045 ( .A(n4062), .ZN(n4022) );
  NOR2_X1 U3046 ( .A1(n2651), .A2(n4954), .ZN(n2663) );
  OR2_X1 U3047 ( .A1(n2892), .A2(n2874), .ZN(n3610) );
  INV_X1 U3048 ( .A(n2884), .ZN(n2868) );
  INV_X1 U3049 ( .A(REG3_REG_16__SCAN_IN), .ZN(n4383) );
  OR2_X1 U3050 ( .A1(n3978), .A2(n3650), .ZN(n3999) );
  OR2_X1 U3051 ( .A1(n4382), .A2(n2853), .ZN(n4158) );
  OAI21_X1 U3052 ( .B1(n3206), .B2(n2590), .A(n2589), .ZN(n3176) );
  INV_X1 U3053 ( .A(n4244), .ZN(n4215) );
  INV_X1 U3054 ( .A(n3308), .ZN(n3229) );
  INV_X1 U3055 ( .A(n4223), .ZN(n4199) );
  INV_X1 U3056 ( .A(n4618), .ZN(n4624) );
  NAND2_X1 U3057 ( .A1(n2792), .A2(n2785), .ZN(n2786) );
  OR2_X1 U3058 ( .A1(n2640), .A2(n4383), .ZN(n2651) );
  INV_X1 U3059 ( .A(n4384), .ZN(n3622) );
  INV_X1 U3060 ( .A(n3610), .ZN(n4390) );
  AND2_X1 U3061 ( .A1(n2722), .A2(n2717), .ZN(n3990) );
  AND2_X1 U3062 ( .A1(n3799), .A2(n3798), .ZN(n4408) );
  AND2_X1 U3063 ( .A1(n2937), .A2(n4376), .ZN(n4244) );
  NAND2_X1 U3064 ( .A1(n2773), .A2(n2772), .ZN(n4223) );
  INV_X1 U3065 ( .A(n3662), .ZN(n4222) );
  INV_X1 U3066 ( .A(n4377), .ZN(n3941) );
  AND2_X1 U3067 ( .A1(n4207), .A2(n2916), .ZN(n3951) );
  OAI22_X1 U3068 ( .A1(n3398), .A2(D_REG_0__SCAN_IN), .B1(n2795), .B2(n4374), 
        .ZN(n2910) );
  NAND2_X1 U3069 ( .A1(n2659), .A2(DATAI_27_), .ZN(n3971) );
  INV_X1 U3070 ( .A(n3620), .ZN(n4202) );
  INV_X1 U3071 ( .A(n4588), .ZN(n3400) );
  AND2_X1 U3072 ( .A1(n3798), .A2(n3797), .ZN(n4541) );
  AND2_X1 U3073 ( .A1(n3015), .A2(n3014), .ZN(n4401) );
  INV_X1 U3074 ( .A(n3479), .ZN(n3966) );
  NAND2_X1 U3075 ( .A1(n2713), .A2(n2712), .ZN(n4024) );
  NAND2_X1 U3076 ( .A1(n4408), .A2(n4382), .ZN(n4548) );
  NAND2_X1 U3077 ( .A1(n4207), .A2(n2917), .ZN(n4204) );
  INV_X1 U3078 ( .A(n3951), .ZN(n4211) );
  OR2_X1 U3079 ( .A1(n3954), .A2(n4309), .ZN(n2830) );
  NAND2_X1 U3080 ( .A1(n4646), .A2(n4629), .ZN(n4309) );
  OR2_X1 U3081 ( .A1(n2826), .A2(n2910), .ZN(n4643) );
  OR2_X1 U3082 ( .A1(n4230), .A2(n3231), .ZN(n3250) );
  INV_X2 U3083 ( .A(n4630), .ZN(n4631) );
  XNOR2_X1 U3084 ( .A(n2775), .B(n4801), .ZN(n4382) );
  AND2_X1 U3085 ( .A1(n2738), .A2(n2685), .ZN(n4377) );
  INV_X1 U3086 ( .A(n3879), .ZN(n4592) );
  INV_X1 U3087 ( .A(n3795), .ZN(U4043) );
  NAND2_X1 U3088 ( .A1(n2739), .A2(n2683), .ZN(n2440) );
  INV_X1 U3089 ( .A(IR_REG_27__SCAN_IN), .ZN(n2442) );
  AND2_X1 U3090 ( .A1(n2443), .A2(n2458), .ZN(n2444) );
  AND2_X1 U3091 ( .A1(n2457), .A2(n2444), .ZN(n2445) );
  INV_X1 U3092 ( .A(n2448), .ZN(n2447) );
  NAND2_X1 U3093 ( .A1(n2447), .A2(n2446), .ZN(n2835) );
  NAND2_X1 U3094 ( .A1(n2526), .A2(REG3_REG_5__SCAN_IN), .ZN(n2534) );
  NOR2_X1 U3095 ( .A1(n2534), .A2(n3073), .ZN(n2545) );
  NAND2_X1 U3096 ( .A1(n2545), .A2(REG3_REG_7__SCAN_IN), .ZN(n2554) );
  NOR2_X1 U3097 ( .A1(n2568), .A2(n2567), .ZN(n2580) );
  NAND2_X1 U3098 ( .A1(n2592), .A2(REG3_REG_11__SCAN_IN), .ZN(n2603) );
  NAND2_X1 U3099 ( .A1(n2630), .A2(REG3_REG_15__SCAN_IN), .ZN(n2640) );
  NOR2_X1 U3100 ( .A1(n2688), .A2(REG3_REG_22__SCAN_IN), .ZN(n2450) );
  OR2_X1 U3101 ( .A1(n2696), .A2(n2450), .ZN(n4069) );
  OR2_X1 U3102 ( .A1(n2493), .A2(n4069), .ZN(n2456) );
  INV_X1 U3103 ( .A(n4373), .ZN(n2451) );
  NAND2_X1 U3104 ( .A1(n2502), .A2(REG1_REG_22__SCAN_IN), .ZN(n2455) );
  INV_X1 U3105 ( .A(n2838), .ZN(n2452) );
  NAND2_X1 U3106 ( .A1(n2219), .A2(REG2_REG_22__SCAN_IN), .ZN(n2454) );
  INV_X1 U3107 ( .A(REG0_REG_22__SCAN_IN), .ZN(n4338) );
  OR2_X1 U3108 ( .A1(n3632), .A2(n4338), .ZN(n2453) );
  NAND4_X1 U3109 ( .A1(n2456), .A2(n2455), .A3(n2454), .A4(n2453), .ZN(n4081)
         );
  NAND2_X1 U3110 ( .A1(n2824), .A2(IR_REG_28__SCAN_IN), .ZN(n2460) );
  NAND2_X1 U3111 ( .A1(n2460), .A2(IR_REG_27__SCAN_IN), .ZN(n2464) );
  NAND2_X1 U3112 ( .A1(n2461), .A2(n4801), .ZN(n2462) );
  NAND2_X1 U3113 ( .A1(n2502), .A2(REG1_REG_20__SCAN_IN), .ZN(n2469) );
  NAND2_X1 U3114 ( .A1(n2218), .A2(REG2_REG_20__SCAN_IN), .ZN(n2468) );
  INV_X1 U3115 ( .A(REG0_REG_20__SCAN_IN), .ZN(n4346) );
  OR2_X1 U3116 ( .A1(n2492), .A2(n4346), .ZN(n2467) );
  NAND2_X1 U3117 ( .A1(n2677), .A2(n4777), .ZN(n2465) );
  NAND2_X1 U3118 ( .A1(n2687), .A2(n2465), .ZN(n4110) );
  OR2_X1 U3119 ( .A1(n2493), .A2(n4110), .ZN(n2466) );
  NAND4_X1 U3120 ( .A1(n2469), .A2(n2468), .A3(n2467), .A4(n2466), .ZN(n4122)
         );
  INV_X1 U3121 ( .A(REG0_REG_1__SCAN_IN), .ZN(n2470) );
  OR2_X1 U3122 ( .A1(n2492), .A2(n2470), .ZN(n2475) );
  NAND2_X1 U3123 ( .A1(n2471), .A2(REG3_REG_1__SCAN_IN), .ZN(n2474) );
  NAND2_X1 U3124 ( .A1(n2485), .A2(REG2_REG_1__SCAN_IN), .ZN(n2472) );
  INV_X1 U3125 ( .A(n2885), .ZN(n2483) );
  NAND2_X1 U3126 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n2476)
         );
  MUX2_X1 U3127 ( .A(IR_REG_31__SCAN_IN), .B(n2476), .S(IR_REG_1__SCAN_IN), 
        .Z(n2479) );
  INV_X1 U3128 ( .A(n2477), .ZN(n2478) );
  INV_X1 U3129 ( .A(DATAI_1_), .ZN(n2480) );
  NAND2_X1 U3130 ( .A1(n2744), .A2(n3701), .ZN(n2743) );
  INV_X1 U3131 ( .A(REG0_REG_0__SCAN_IN), .ZN(n2484) );
  NAND2_X1 U3132 ( .A1(n2502), .A2(REG1_REG_0__SCAN_IN), .ZN(n2488) );
  NAND2_X1 U3133 ( .A1(n2219), .A2(REG2_REG_0__SCAN_IN), .ZN(n2487) );
  INV_X1 U3134 ( .A(REG3_REG_0__SCAN_IN), .ZN(n2880) );
  NAND2_X1 U3135 ( .A1(n2743), .A2(n2960), .ZN(n2959) );
  NAND2_X1 U3136 ( .A1(n2887), .A2(n2895), .ZN(n2491) );
  AND2_X1 U3137 ( .A1(n2959), .A2(n2491), .ZN(n2975) );
  NAND2_X1 U3138 ( .A1(n2218), .A2(REG2_REG_2__SCAN_IN), .ZN(n2496) );
  INV_X1 U3139 ( .A(REG0_REG_2__SCAN_IN), .ZN(n4612) );
  INV_X1 U3140 ( .A(REG3_REG_2__SCAN_IN), .ZN(n2981) );
  OR2_X1 U3141 ( .A1(n2493), .A2(n2981), .ZN(n2494) );
  INV_X1 U3142 ( .A(DATAI_2_), .ZN(n2500) );
  MUX2_X1 U3143 ( .A(n3836), .B(n2500), .S(n2499), .Z(n2984) );
  NAND2_X1 U3144 ( .A1(n3794), .A2(n2984), .ZN(n3708) );
  NAND2_X1 U3145 ( .A1(n2975), .A2(n3660), .ZN(n2974) );
  OR2_X1 U3146 ( .A1(n3794), .A2(n2977), .ZN(n2501) );
  NAND2_X1 U3147 ( .A1(n2502), .A2(REG1_REG_3__SCAN_IN), .ZN(n2507) );
  NAND2_X1 U31480 ( .A1(n2219), .A2(REG2_REG_3__SCAN_IN), .ZN(n2506) );
  OR2_X1 U31490 ( .A1(n2493), .A2(REG3_REG_3__SCAN_IN), .ZN(n2505) );
  INV_X1 U3150 ( .A(REG0_REG_3__SCAN_IN), .ZN(n2503) );
  OR2_X1 U3151 ( .A1(n2492), .A2(n2503), .ZN(n2504) );
  NAND2_X1 U3152 ( .A1(n2508), .A2(IR_REG_31__SCAN_IN), .ZN(n2520) );
  XNOR2_X1 U3153 ( .A(n2520), .B(IR_REG_3__SCAN_IN), .ZN(n4380) );
  NOR2_X1 U3154 ( .A1(n3793), .A2(n3019), .ZN(n2510) );
  NAND2_X1 U3155 ( .A1(n3793), .A2(n3019), .ZN(n2509) );
  OAI21_X1 U3156 ( .B1(n2899), .B2(n2510), .A(n2509), .ZN(n2924) );
  NAND2_X1 U3157 ( .A1(n2502), .A2(REG1_REG_4__SCAN_IN), .ZN(n2518) );
  NAND2_X1 U3158 ( .A1(n2218), .A2(REG2_REG_4__SCAN_IN), .ZN(n2517) );
  INV_X1 U3159 ( .A(REG0_REG_4__SCAN_IN), .ZN(n2511) );
  OR2_X1 U3160 ( .A1(n2492), .A2(n2511), .ZN(n2516) );
  INV_X1 U3161 ( .A(n2526), .ZN(n2514) );
  INV_X1 U3162 ( .A(REG3_REG_3__SCAN_IN), .ZN(n3016) );
  INV_X1 U3163 ( .A(REG3_REG_4__SCAN_IN), .ZN(n2512) );
  NAND2_X1 U3164 ( .A1(n3016), .A2(n2512), .ZN(n2513) );
  NAND2_X1 U3165 ( .A1(n2514), .A2(n2513), .ZN(n3578) );
  OR2_X1 U3166 ( .A1(n2493), .A2(n3578), .ZN(n2515) );
  NAND2_X1 U3167 ( .A1(n2520), .A2(n2519), .ZN(n2521) );
  NAND2_X1 U3168 ( .A1(n2521), .A2(IR_REG_31__SCAN_IN), .ZN(n2522) );
  XNOR2_X1 U3169 ( .A(n2522), .B(n4800), .ZN(n3898) );
  INV_X1 U3170 ( .A(DATAI_4_), .ZN(n4846) );
  INV_X1 U3171 ( .A(n3040), .ZN(n3577) );
  NAND2_X1 U3172 ( .A1(n3792), .A2(n3577), .ZN(n2523) );
  NAND2_X1 U3173 ( .A1(n2502), .A2(REG1_REG_5__SCAN_IN), .ZN(n2530) );
  NAND2_X1 U3174 ( .A1(n2218), .A2(REG2_REG_5__SCAN_IN), .ZN(n2529) );
  INV_X1 U3175 ( .A(REG0_REG_5__SCAN_IN), .ZN(n2525) );
  OR2_X1 U3176 ( .A1(n2492), .A2(n2525), .ZN(n2528) );
  OAI21_X1 U3177 ( .B1(n2526), .B2(REG3_REG_5__SCAN_IN), .A(n2534), .ZN(n3055)
         );
  OR2_X1 U3178 ( .A1(n2493), .A2(n3055), .ZN(n2527) );
  NAND4_X1 U3179 ( .A1(n2530), .A2(n2529), .A3(n2528), .A4(n2527), .ZN(n3791)
         );
  NAND2_X1 U3180 ( .A1(n2531), .A2(IR_REG_31__SCAN_IN), .ZN(n2532) );
  XNOR2_X1 U3181 ( .A(n2532), .B(IR_REG_5__SCAN_IN), .ZN(n3896) );
  MUX2_X1 U3182 ( .A(n3896), .B(DATAI_5_), .S(n2659), .Z(n3047) );
  AND2_X1 U3183 ( .A1(n3791), .A2(n3047), .ZN(n2533) );
  NAND2_X1 U3184 ( .A1(n2502), .A2(REG1_REG_6__SCAN_IN), .ZN(n2540) );
  NAND2_X1 U3185 ( .A1(n2218), .A2(REG2_REG_6__SCAN_IN), .ZN(n2539) );
  AND2_X1 U3186 ( .A1(n2534), .A2(n3073), .ZN(n2535) );
  NOR2_X1 U3187 ( .A1(n2545), .A2(n2535), .ZN(n4566) );
  INV_X1 U3188 ( .A(n4566), .ZN(n3076) );
  OR2_X1 U3189 ( .A1(n2493), .A2(n3076), .ZN(n2538) );
  INV_X1 U3190 ( .A(REG0_REG_6__SCAN_IN), .ZN(n2536) );
  OR2_X1 U3191 ( .A1(n3632), .A2(n2536), .ZN(n2537) );
  NAND4_X1 U3192 ( .A1(n2540), .A2(n2539), .A3(n2538), .A4(n2537), .ZN(n3790)
         );
  NOR2_X1 U3193 ( .A1(n2531), .A2(IR_REG_5__SCAN_IN), .ZN(n2577) );
  OR2_X1 U3194 ( .A1(n2577), .A2(n2459), .ZN(n2541) );
  XNOR2_X1 U3195 ( .A(n2541), .B(IR_REG_6__SCAN_IN), .ZN(n3903) );
  MUX2_X1 U3196 ( .A(n3903), .B(DATAI_6_), .S(n2659), .Z(n3084) );
  NOR2_X1 U3197 ( .A1(n3790), .A2(n3084), .ZN(n2543) );
  NAND2_X1 U3198 ( .A1(n3790), .A2(n3084), .ZN(n2542) );
  NAND2_X1 U3199 ( .A1(n2502), .A2(REG1_REG_7__SCAN_IN), .ZN(n2550) );
  NAND2_X1 U3200 ( .A1(n2219), .A2(REG2_REG_7__SCAN_IN), .ZN(n2549) );
  INV_X1 U3201 ( .A(REG0_REG_7__SCAN_IN), .ZN(n2544) );
  OR2_X1 U3202 ( .A1(n2492), .A2(n2544), .ZN(n2548) );
  OR2_X1 U3203 ( .A1(n2545), .A2(REG3_REG_7__SCAN_IN), .ZN(n2546) );
  NAND2_X1 U3204 ( .A1(n2554), .A2(n2546), .ZN(n3136) );
  OR2_X1 U3205 ( .A1(n2493), .A2(n3136), .ZN(n2547) );
  NAND4_X1 U3206 ( .A1(n2550), .A2(n2549), .A3(n2548), .A4(n2547), .ZN(n3789)
         );
  NAND2_X1 U3207 ( .A1(n2577), .A2(n2574), .ZN(n2551) );
  NAND2_X1 U3208 ( .A1(n2551), .A2(IR_REG_31__SCAN_IN), .ZN(n2562) );
  XNOR2_X1 U3209 ( .A(n2562), .B(IR_REG_7__SCAN_IN), .ZN(n4432) );
  INV_X1 U32100 ( .A(DATAI_7_), .ZN(n2552) );
  MUX2_X1 U32110 ( .A(n4597), .B(n2552), .S(n2659), .Z(n3128) );
  NAND2_X1 U32120 ( .A1(n3789), .A2(n3128), .ZN(n3727) );
  OR2_X1 U32130 ( .A1(n3789), .A2(n3128), .ZN(n2750) );
  NAND2_X1 U32140 ( .A1(n3727), .A2(n2750), .ZN(n3716) );
  NAND2_X1 U32150 ( .A1(n3789), .A2(n3133), .ZN(n2553) );
  NAND2_X1 U32160 ( .A1(n2502), .A2(REG1_REG_8__SCAN_IN), .ZN(n2560) );
  NAND2_X1 U32170 ( .A1(n2219), .A2(REG2_REG_8__SCAN_IN), .ZN(n2559) );
  NAND2_X1 U32180 ( .A1(n2554), .A2(n4958), .ZN(n2555) );
  AND2_X1 U32190 ( .A1(n2568), .A2(n2555), .ZN(n4557) );
  INV_X1 U32200 ( .A(n4557), .ZN(n3159) );
  OR2_X1 U32210 ( .A1(n2493), .A2(n3159), .ZN(n2558) );
  INV_X1 U32220 ( .A(REG0_REG_8__SCAN_IN), .ZN(n2556) );
  OR2_X1 U32230 ( .A1(n3632), .A2(n2556), .ZN(n2557) );
  NAND4_X1 U32240 ( .A1(n2560), .A2(n2559), .A3(n2558), .A4(n2557), .ZN(n3788)
         );
  INV_X1 U32250 ( .A(IR_REG_7__SCAN_IN), .ZN(n2561) );
  NAND2_X1 U32260 ( .A1(n2562), .A2(n2561), .ZN(n2563) );
  NAND2_X1 U32270 ( .A1(n2563), .A2(IR_REG_31__SCAN_IN), .ZN(n2564) );
  XNOR2_X1 U32280 ( .A(n2564), .B(IR_REG_8__SCAN_IN), .ZN(n4443) );
  MUX2_X1 U32290 ( .A(n4443), .B(DATAI_8_), .S(n2659), .Z(n3156) );
  AND2_X1 U32300 ( .A1(n3788), .A2(n3156), .ZN(n2565) );
  OR2_X1 U32310 ( .A1(n3788), .A2(n3156), .ZN(n2566) );
  NAND2_X1 U32320 ( .A1(n2502), .A2(REG1_REG_9__SCAN_IN), .ZN(n2573) );
  NAND2_X1 U32330 ( .A1(n2219), .A2(REG2_REG_9__SCAN_IN), .ZN(n2572) );
  INV_X1 U32340 ( .A(REG0_REG_9__SCAN_IN), .ZN(n3106) );
  OR2_X1 U32350 ( .A1(n3632), .A2(n3106), .ZN(n2571) );
  AND2_X1 U32360 ( .A1(n2568), .A2(n2567), .ZN(n2569) );
  OR2_X1 U32370 ( .A1(n2569), .A2(n2580), .ZN(n3200) );
  OR2_X1 U32380 ( .A1(n2493), .A2(n3200), .ZN(n2570) );
  NAND4_X1 U32390 ( .A1(n2573), .A2(n2572), .A3(n2571), .A4(n2570), .ZN(n3787)
         );
  AND2_X1 U32400 ( .A1(n2575), .A2(n2574), .ZN(n2576) );
  AND2_X1 U32410 ( .A1(n2577), .A2(n2576), .ZN(n2587) );
  OR2_X1 U32420 ( .A1(n2587), .A2(n2459), .ZN(n2578) );
  XNOR2_X1 U32430 ( .A(n2578), .B(IR_REG_9__SCAN_IN), .ZN(n3893) );
  MUX2_X1 U32440 ( .A(n3893), .B(DATAI_9_), .S(n2659), .Z(n3197) );
  NOR2_X1 U32450 ( .A1(n3787), .A2(n3197), .ZN(n2579) );
  INV_X1 U32460 ( .A(n3787), .ZN(n3208) );
  INV_X1 U32470 ( .A(n3197), .ZN(n3196) );
  NAND2_X1 U32480 ( .A1(n2502), .A2(REG1_REG_10__SCAN_IN), .ZN(n2586) );
  NAND2_X1 U32490 ( .A1(n2218), .A2(REG2_REG_10__SCAN_IN), .ZN(n2585) );
  NOR2_X1 U32500 ( .A1(n2580), .A2(REG3_REG_10__SCAN_IN), .ZN(n2581) );
  OR2_X1 U32510 ( .A1(n2592), .A2(n2581), .ZN(n4549) );
  OR2_X1 U32520 ( .A1(n2493), .A2(n4549), .ZN(n2584) );
  INV_X1 U32530 ( .A(REG0_REG_10__SCAN_IN), .ZN(n2582) );
  OR2_X1 U32540 ( .A1(n3632), .A2(n2582), .ZN(n2583) );
  NAND4_X1 U32550 ( .A1(n2586), .A2(n2585), .A3(n2584), .A4(n2583), .ZN(n3786)
         );
  NAND2_X1 U32560 ( .A1(n2587), .A2(n4933), .ZN(n2598) );
  NAND2_X1 U32570 ( .A1(n2598), .A2(IR_REG_31__SCAN_IN), .ZN(n2588) );
  XNOR2_X1 U32580 ( .A(n2588), .B(IR_REG_10__SCAN_IN), .ZN(n4464) );
  MUX2_X1 U32590 ( .A(n4464), .B(DATAI_10_), .S(n2659), .Z(n3269) );
  AND2_X1 U32600 ( .A1(n3786), .A2(n3269), .ZN(n2590) );
  OR2_X1 U32610 ( .A1(n3786), .A2(n3269), .ZN(n2589) );
  NAND2_X1 U32620 ( .A1(n2502), .A2(REG1_REG_11__SCAN_IN), .ZN(n2597) );
  NAND2_X1 U32630 ( .A1(n2219), .A2(REG2_REG_11__SCAN_IN), .ZN(n2596) );
  INV_X1 U32640 ( .A(REG0_REG_11__SCAN_IN), .ZN(n2591) );
  OR2_X1 U32650 ( .A1(n3632), .A2(n2591), .ZN(n2595) );
  OR2_X1 U32660 ( .A1(n2592), .A2(REG3_REG_11__SCAN_IN), .ZN(n2593) );
  NAND2_X1 U32670 ( .A1(n2603), .A2(n2593), .ZN(n3289) );
  OR2_X1 U32680 ( .A1(n2493), .A2(n3289), .ZN(n2594) );
  NAND4_X1 U32690 ( .A1(n2597), .A2(n2596), .A3(n2595), .A4(n2594), .ZN(n3785)
         );
  NAND2_X1 U32700 ( .A1(n2599), .A2(IR_REG_31__SCAN_IN), .ZN(n2610) );
  XNOR2_X1 U32710 ( .A(n2610), .B(IR_REG_11__SCAN_IN), .ZN(n3891) );
  INV_X1 U32720 ( .A(DATAI_11_), .ZN(n2600) );
  MUX2_X1 U32730 ( .A(n4595), .B(n2600), .S(n2659), .Z(n3179) );
  OR2_X1 U32740 ( .A1(n3785), .A2(n3179), .ZN(n3163) );
  NAND2_X1 U32750 ( .A1(n3785), .A2(n3179), .ZN(n3165) );
  NAND2_X1 U32760 ( .A1(n3163), .A2(n3165), .ZN(n3656) );
  OR2_X1 U32770 ( .A1(n3785), .A2(n3286), .ZN(n2601) );
  NAND2_X1 U32780 ( .A1(n2502), .A2(REG1_REG_12__SCAN_IN), .ZN(n2608) );
  NAND2_X1 U32790 ( .A1(n2219), .A2(REG2_REG_12__SCAN_IN), .ZN(n2607) );
  INV_X1 U32800 ( .A(REG0_REG_12__SCAN_IN), .ZN(n2602) );
  OR2_X1 U32810 ( .A1(n3632), .A2(n2602), .ZN(n2606) );
  NAND2_X1 U32820 ( .A1(n2603), .A2(n4955), .ZN(n2604) );
  NAND2_X1 U32830 ( .A1(n2614), .A2(n2604), .ZN(n3537) );
  OR2_X1 U32840 ( .A1(n2493), .A2(n3537), .ZN(n2605) );
  NAND4_X1 U32850 ( .A1(n2608), .A2(n2607), .A3(n2606), .A4(n2605), .ZN(n3784)
         );
  INV_X1 U32860 ( .A(IR_REG_11__SCAN_IN), .ZN(n2609) );
  NAND2_X1 U32870 ( .A1(n2610), .A2(n2609), .ZN(n2611) );
  NAND2_X1 U32880 ( .A1(n2611), .A2(IR_REG_31__SCAN_IN), .ZN(n2612) );
  XNOR2_X1 U32890 ( .A(n2612), .B(IR_REG_12__SCAN_IN), .ZN(n4485) );
  MUX2_X1 U32900 ( .A(n4485), .B(DATAI_12_), .S(n2659), .Z(n3534) );
  INV_X1 U32910 ( .A(n3784), .ZN(n3180) );
  NAND2_X1 U32920 ( .A1(n2502), .A2(REG1_REG_13__SCAN_IN), .ZN(n2619) );
  NAND2_X1 U32930 ( .A1(n2218), .A2(REG2_REG_13__SCAN_IN), .ZN(n2618) );
  INV_X1 U32940 ( .A(REG0_REG_13__SCAN_IN), .ZN(n3248) );
  OR2_X1 U32950 ( .A1(n2492), .A2(n3248), .ZN(n2617) );
  NAND2_X1 U32960 ( .A1(n2614), .A2(n2613), .ZN(n2615) );
  NAND2_X1 U32970 ( .A1(n2622), .A2(n2615), .ZN(n3311) );
  OR2_X1 U32980 ( .A1(n2493), .A2(n3311), .ZN(n2616) );
  NAND4_X1 U32990 ( .A1(n2619), .A2(n2618), .A3(n2617), .A4(n2616), .ZN(n4218)
         );
  OR2_X1 U33000 ( .A1(n2620), .A2(n2459), .ZN(n2621) );
  XNOR2_X1 U33010 ( .A(n2621), .B(IR_REG_13__SCAN_IN), .ZN(n3915) );
  MUX2_X1 U33020 ( .A(n3915), .B(DATAI_13_), .S(n2659), .Z(n3308) );
  OR2_X1 U33030 ( .A1(n4218), .A2(n3308), .ZN(n3223) );
  NAND2_X1 U33040 ( .A1(n2502), .A2(REG1_REG_14__SCAN_IN), .ZN(n2627) );
  NAND2_X1 U33050 ( .A1(n2218), .A2(REG2_REG_14__SCAN_IN), .ZN(n2626) );
  INV_X1 U33060 ( .A(REG0_REG_14__SCAN_IN), .ZN(n4369) );
  OR2_X1 U33070 ( .A1(n3632), .A2(n4369), .ZN(n2625) );
  AND2_X1 U33080 ( .A1(n2622), .A2(n4744), .ZN(n2623) );
  OR2_X1 U33090 ( .A1(n2623), .A2(n2630), .ZN(n4232) );
  OR2_X1 U33100 ( .A1(n2493), .A2(n4232), .ZN(n2624) );
  NAND4_X1 U33110 ( .A1(n2627), .A2(n2626), .A3(n2625), .A4(n2624), .ZN(n4196)
         );
  NAND2_X1 U33120 ( .A1(n2628), .A2(IR_REG_31__SCAN_IN), .ZN(n2629) );
  XNOR2_X1 U33130 ( .A(n2629), .B(IR_REG_14__SCAN_IN), .ZN(n3879) );
  INV_X1 U33140 ( .A(DATAI_14_), .ZN(n4980) );
  MUX2_X1 U33150 ( .A(n4592), .B(n4980), .S(n2659), .Z(n4229) );
  OR2_X1 U33160 ( .A1(n4196), .A2(n4229), .ZN(n4190) );
  NAND2_X1 U33170 ( .A1(n4196), .A2(n4229), .ZN(n3671) );
  NAND2_X1 U33180 ( .A1(n4190), .A2(n3671), .ZN(n3662) );
  NAND2_X1 U33190 ( .A1(n4218), .A2(n3308), .ZN(n4186) );
  NAND2_X1 U33200 ( .A1(n2502), .A2(REG1_REG_15__SCAN_IN), .ZN(n2635) );
  NAND2_X1 U33210 ( .A1(n2218), .A2(REG2_REG_15__SCAN_IN), .ZN(n2634) );
  INV_X1 U33220 ( .A(REG0_REG_15__SCAN_IN), .ZN(n4365) );
  OR2_X1 U33230 ( .A1(n3632), .A2(n4365), .ZN(n2633) );
  OR2_X1 U33240 ( .A1(n2630), .A2(REG3_REG_15__SCAN_IN), .ZN(n2631) );
  NAND2_X1 U33250 ( .A1(n2640), .A2(n2631), .ZN(n4205) );
  OR2_X1 U33260 ( .A1(n2493), .A2(n4205), .ZN(n2632) );
  NAND4_X1 U33270 ( .A1(n2635), .A2(n2634), .A3(n2633), .A4(n2632), .ZN(n4171)
         );
  NAND2_X1 U33280 ( .A1(n2251), .A2(IR_REG_31__SCAN_IN), .ZN(n2647) );
  XNOR2_X1 U33290 ( .A(n2647), .B(IR_REG_15__SCAN_IN), .ZN(n3919) );
  MUX2_X1 U33300 ( .A(n3919), .B(DATAI_15_), .S(n2659), .Z(n3620) );
  NAND2_X1 U33310 ( .A1(n4171), .A2(n3620), .ZN(n2638) );
  INV_X1 U33320 ( .A(n4229), .ZN(n3488) );
  NOR2_X1 U33330 ( .A1(n4196), .A2(n3488), .ZN(n4188) );
  INV_X1 U33340 ( .A(n4171), .ZN(n4385) );
  AOI22_X1 U33350 ( .A1(n4188), .A2(n2638), .B1(n4385), .B2(n4202), .ZN(n2639)
         );
  NAND2_X1 U33360 ( .A1(n2502), .A2(REG1_REG_16__SCAN_IN), .ZN(n2645) );
  NAND2_X1 U33370 ( .A1(n2219), .A2(REG2_REG_16__SCAN_IN), .ZN(n2644) );
  NAND2_X1 U33380 ( .A1(n2640), .A2(n4383), .ZN(n2641) );
  NAND2_X1 U33390 ( .A1(n2651), .A2(n2641), .ZN(n4400) );
  OR2_X1 U33400 ( .A1(n2493), .A2(n4400), .ZN(n2643) );
  INV_X1 U33410 ( .A(REG0_REG_16__SCAN_IN), .ZN(n4360) );
  OR2_X1 U33420 ( .A1(n3632), .A2(n4360), .ZN(n2642) );
  NAND4_X1 U33430 ( .A1(n2645), .A2(n2644), .A3(n2643), .A4(n2642), .ZN(n4195)
         );
  NAND2_X1 U33440 ( .A1(n2647), .A2(n2646), .ZN(n2648) );
  NAND2_X1 U33450 ( .A1(n2648), .A2(IR_REG_31__SCAN_IN), .ZN(n2649) );
  XNOR2_X1 U33460 ( .A(n2649), .B(IR_REG_16__SCAN_IN), .ZN(n3883) );
  MUX2_X1 U33470 ( .A(n4590), .B(n4989), .S(n2659), .Z(n4386) );
  OR2_X1 U33480 ( .A1(n4195), .A2(n4386), .ZN(n3745) );
  NAND2_X1 U33490 ( .A1(n4195), .A2(n4386), .ZN(n3747) );
  INV_X1 U33500 ( .A(n4195), .ZN(n4159) );
  NAND2_X1 U33510 ( .A1(n2502), .A2(REG1_REG_17__SCAN_IN), .ZN(n2656) );
  NAND2_X1 U33520 ( .A1(n2218), .A2(REG2_REG_17__SCAN_IN), .ZN(n2655) );
  AND2_X1 U3353 ( .A1(n2651), .A2(n4954), .ZN(n2652) );
  OR2_X1 U33540 ( .A1(n2652), .A2(n2663), .ZN(n4163) );
  OR2_X1 U3355 ( .A1(n2493), .A2(n4163), .ZN(n2654) );
  INV_X1 U3356 ( .A(REG0_REG_17__SCAN_IN), .ZN(n4355) );
  OR2_X1 U3357 ( .A1(n3632), .A2(n4355), .ZN(n2653) );
  NAND4_X1 U3358 ( .A1(n2656), .A2(n2655), .A3(n2654), .A4(n2653), .ZN(n4389)
         );
  INV_X1 U3359 ( .A(n4389), .ZN(n4138) );
  NAND2_X1 U3360 ( .A1(n2657), .A2(IR_REG_31__SCAN_IN), .ZN(n2658) );
  XNOR2_X1 U3361 ( .A(n2658), .B(IR_REG_17__SCAN_IN), .ZN(n3922) );
  INV_X1 U3362 ( .A(n3922), .ZN(n4589) );
  INV_X1 U3363 ( .A(DATAI_17_), .ZN(n2660) );
  MUX2_X1 U3364 ( .A(n4589), .B(n2660), .S(n2659), .Z(n4162) );
  NAND2_X1 U3365 ( .A1(n4138), .A2(n4162), .ZN(n2661) );
  INV_X1 U3366 ( .A(n4162), .ZN(n3558) );
  NAND2_X1 U3367 ( .A1(n2502), .A2(REG1_REG_18__SCAN_IN), .ZN(n2668) );
  NAND2_X1 U3368 ( .A1(n2219), .A2(REG2_REG_18__SCAN_IN), .ZN(n2667) );
  INV_X1 U3369 ( .A(REG0_REG_18__SCAN_IN), .ZN(n2662) );
  OR2_X1 U3370 ( .A1(n3632), .A2(n2662), .ZN(n2666) );
  NOR2_X1 U3371 ( .A1(n2663), .A2(REG3_REG_18__SCAN_IN), .ZN(n2664) );
  OR2_X1 U3372 ( .A1(n2675), .A2(n2664), .ZN(n4141) );
  OR2_X1 U3373 ( .A1(n2493), .A2(n4141), .ZN(n2665) );
  NAND4_X1 U3374 ( .A1(n2668), .A2(n2667), .A3(n2666), .A4(n2665), .ZN(n4155)
         );
  OR2_X1 U3375 ( .A1(n2669), .A2(n2459), .ZN(n2671) );
  XNOR2_X1 U3376 ( .A(n2671), .B(n2670), .ZN(n3927) );
  INV_X1 U3377 ( .A(DATAI_18_), .ZN(n2672) );
  MUX2_X1 U3378 ( .A(n3927), .B(n2672), .S(n2659), .Z(n4133) );
  OR2_X1 U3379 ( .A1(n4155), .A2(n4133), .ZN(n2764) );
  NAND2_X1 U3380 ( .A1(n4155), .A2(n4133), .ZN(n4117) );
  NAND2_X1 U3381 ( .A1(n2764), .A2(n4117), .ZN(n4143) );
  NAND2_X1 U3382 ( .A1(n4144), .A2(n4143), .ZN(n4142) );
  INV_X1 U3383 ( .A(n4133), .ZN(n4135) );
  NAND2_X1 U3384 ( .A1(n4142), .A2(n2674), .ZN(n4116) );
  NAND2_X1 U3385 ( .A1(n2502), .A2(REG1_REG_19__SCAN_IN), .ZN(n2681) );
  NAND2_X1 U3386 ( .A1(n2219), .A2(REG2_REG_19__SCAN_IN), .ZN(n2680) );
  INV_X1 U3387 ( .A(REG0_REG_19__SCAN_IN), .ZN(n4350) );
  OR2_X1 U3388 ( .A1(n2492), .A2(n4350), .ZN(n2679) );
  OR2_X1 U3389 ( .A1(n2675), .A2(REG3_REG_19__SCAN_IN), .ZN(n2676) );
  NAND2_X1 U3390 ( .A1(n2677), .A2(n2676), .ZN(n4127) );
  OR2_X1 U3391 ( .A1(n2493), .A2(n4127), .ZN(n2678) );
  NAND4_X1 U3392 ( .A1(n2681), .A2(n2680), .A3(n2679), .A4(n2678), .ZN(n4136)
         );
  NAND2_X1 U3393 ( .A1(n2684), .A2(n2683), .ZN(n2738) );
  OR2_X1 U3394 ( .A1(n2684), .A2(n2683), .ZN(n2685) );
  MUX2_X1 U3395 ( .A(n4377), .B(DATAI_19_), .S(n2659), .Z(n3506) );
  NAND2_X1 U3396 ( .A1(n4136), .A2(n3506), .ZN(n2686) );
  INV_X1 U3397 ( .A(n4136), .ZN(n4103) );
  NAND2_X1 U3398 ( .A1(n2502), .A2(REG1_REG_21__SCAN_IN), .ZN(n2693) );
  NAND2_X1 U3399 ( .A1(n2219), .A2(REG2_REG_21__SCAN_IN), .ZN(n2692) );
  INV_X1 U3400 ( .A(REG0_REG_21__SCAN_IN), .ZN(n4342) );
  OR2_X1 U3401 ( .A1(n2492), .A2(n4342), .ZN(n2691) );
  AND2_X1 U3402 ( .A1(n2687), .A2(n3516), .ZN(n2689) );
  OR2_X1 U3403 ( .A1(n2689), .A2(n2688), .ZN(n4088) );
  OR2_X1 U3404 ( .A1(n2493), .A2(n4088), .ZN(n2690) );
  NAND4_X1 U3405 ( .A1(n2693), .A2(n2692), .A3(n2691), .A4(n2690), .ZN(n4101)
         );
  INV_X1 U3406 ( .A(n4101), .ZN(n4065) );
  NOR2_X1 U3407 ( .A1(n4065), .A2(n4086), .ZN(n2694) );
  INV_X1 U3408 ( .A(n4068), .ZN(n2695) );
  NAND2_X1 U3409 ( .A1(n3316), .A2(n2695), .ZN(n4041) );
  NAND2_X1 U3410 ( .A1(n4081), .A2(n4068), .ZN(n2768) );
  NAND2_X1 U3411 ( .A1(n4041), .A2(n2768), .ZN(n4058) );
  OR2_X1 U3412 ( .A1(n2696), .A2(REG3_REG_23__SCAN_IN), .ZN(n2697) );
  NAND2_X1 U3413 ( .A1(n2702), .A2(n2697), .ZN(n4051) );
  OR2_X1 U3414 ( .A1(n4051), .A2(n2493), .ZN(n2701) );
  NAND2_X1 U3415 ( .A1(n2502), .A2(REG1_REG_23__SCAN_IN), .ZN(n2700) );
  NAND2_X1 U3416 ( .A1(n2218), .A2(REG2_REG_23__SCAN_IN), .ZN(n2699) );
  INV_X1 U3417 ( .A(REG0_REG_23__SCAN_IN), .ZN(n4334) );
  OR2_X1 U3418 ( .A1(n3632), .A2(n4334), .ZN(n2698) );
  NAND4_X1 U3419 ( .A1(n2701), .A2(n2700), .A3(n2699), .A4(n2698), .ZN(n4062)
         );
  INV_X1 U3420 ( .A(n4048), .ZN(n3498) );
  AND2_X1 U3421 ( .A1(n4062), .A2(n3498), .ZN(n3637) );
  NAND2_X1 U3422 ( .A1(n4022), .A2(n4048), .ZN(n3638) );
  NAND2_X1 U3423 ( .A1(n2702), .A2(n4977), .ZN(n2703) );
  NAND2_X1 U3424 ( .A1(n2716), .A2(n2703), .ZN(n4030) );
  NOR2_X1 U3425 ( .A1(n4030), .A2(n2493), .ZN(n2707) );
  AND2_X1 U3426 ( .A1(n2218), .A2(REG2_REG_24__SCAN_IN), .ZN(n2706) );
  INV_X1 U3427 ( .A(REG0_REG_24__SCAN_IN), .ZN(n4330) );
  NAND2_X1 U3428 ( .A1(n2502), .A2(REG1_REG_24__SCAN_IN), .ZN(n2704) );
  OAI21_X1 U3429 ( .B1(n4330), .B2(n2492), .A(n2704), .ZN(n2705) );
  INV_X1 U3430 ( .A(n4027), .ZN(n3568) );
  NAND2_X1 U3431 ( .A1(n4004), .A2(n3568), .ZN(n2708) );
  XNOR2_X1 U3432 ( .A(n2716), .B(REG3_REG_25__SCAN_IN), .ZN(n4012) );
  NAND2_X1 U3433 ( .A1(n4012), .A2(n2471), .ZN(n2713) );
  INV_X1 U3434 ( .A(REG0_REG_25__SCAN_IN), .ZN(n4326) );
  NAND2_X1 U3435 ( .A1(n2502), .A2(REG1_REG_25__SCAN_IN), .ZN(n2710) );
  NAND2_X1 U3436 ( .A1(n2219), .A2(REG2_REG_25__SCAN_IN), .ZN(n2709) );
  OAI211_X1 U3437 ( .C1(n3632), .C2(n4326), .A(n2710), .B(n2709), .ZN(n2711)
         );
  INV_X1 U3438 ( .A(n2711), .ZN(n2712) );
  INV_X1 U3439 ( .A(n4024), .ZN(n3609) );
  NAND2_X1 U3440 ( .A1(n3609), .A2(n4010), .ZN(n2714) );
  INV_X1 U3441 ( .A(n2218), .ZN(n2779) );
  INV_X1 U3442 ( .A(REG2_REG_26__SCAN_IN), .ZN(n2720) );
  NAND2_X1 U3443 ( .A1(REG3_REG_25__SCAN_IN), .A2(REG3_REG_26__SCAN_IN), .ZN(
        n2715) );
  INV_X1 U3444 ( .A(REG3_REG_25__SCAN_IN), .ZN(n3546) );
  INV_X1 U3445 ( .A(REG3_REG_26__SCAN_IN), .ZN(n3608) );
  OAI21_X1 U3446 ( .B1(n2716), .B2(n3546), .A(n3608), .ZN(n2717) );
  NAND2_X1 U3447 ( .A1(n3990), .A2(n2471), .ZN(n2719) );
  INV_X1 U3448 ( .A(n3632), .ZN(n2776) );
  AOI22_X1 U3449 ( .A1(n2776), .A2(REG0_REG_26__SCAN_IN), .B1(n2502), .B2(
        REG1_REG_26__SCAN_IN), .ZN(n2718) );
  INV_X1 U3450 ( .A(n4002), .ZN(n3964) );
  AND2_X1 U3451 ( .A1(n2722), .A2(n4957), .ZN(n2723) );
  AOI22_X1 U3452 ( .A1(n2776), .A2(REG0_REG_27__SCAN_IN), .B1(n2502), .B2(
        REG1_REG_27__SCAN_IN), .ZN(n2725) );
  NAND2_X1 U3453 ( .A1(n2219), .A2(REG2_REG_27__SCAN_IN), .ZN(n2724) );
  OAI211_X1 U3454 ( .C1(n3478), .C2(n2493), .A(n2725), .B(n2724), .ZN(n3983)
         );
  INV_X1 U3455 ( .A(n3971), .ZN(n3439) );
  NOR2_X1 U3456 ( .A1(n3983), .A2(n3439), .ZN(n2726) );
  INV_X1 U3457 ( .A(n3983), .ZN(n3611) );
  NAND2_X1 U34580 ( .A1(n2727), .A2(REG3_REG_28__SCAN_IN), .ZN(n3953) );
  INV_X1 U34590 ( .A(n2727), .ZN(n2729) );
  INV_X1 U3460 ( .A(REG3_REG_28__SCAN_IN), .ZN(n2728) );
  NAND2_X1 U3461 ( .A1(n2729), .A2(n2728), .ZN(n2730) );
  NAND2_X1 U3462 ( .A1(n3953), .A2(n2730), .ZN(n3469) );
  INV_X1 U3463 ( .A(REG0_REG_28__SCAN_IN), .ZN(n2733) );
  NAND2_X1 U3464 ( .A1(n2218), .A2(REG2_REG_28__SCAN_IN), .ZN(n2732) );
  NAND2_X1 U3465 ( .A1(n2502), .A2(REG1_REG_28__SCAN_IN), .ZN(n2731) );
  OAI211_X1 U3466 ( .C1(n3632), .C2(n2733), .A(n2732), .B(n2731), .ZN(n2734)
         );
  INV_X1 U34670 ( .A(n2734), .ZN(n2735) );
  NAND2_X1 U3468 ( .A1(n3966), .A2(n3447), .ZN(n2817) );
  INV_X1 U34690 ( .A(n3447), .ZN(n3459) );
  NAND2_X1 U3470 ( .A1(n3479), .A2(n3459), .ZN(n3686) );
  NAND2_X1 U34710 ( .A1(n2817), .A2(n3686), .ZN(n3636) );
  XNOR2_X1 U3472 ( .A(n2816), .B(n3636), .ZN(n3475) );
  NAND2_X1 U34730 ( .A1(n2241), .A2(IR_REG_31__SCAN_IN), .ZN(n2737) );
  NAND2_X1 U3474 ( .A1(n2738), .A2(IR_REG_31__SCAN_IN), .ZN(n2740) );
  NAND2_X1 U34750 ( .A1(n2242), .A2(IR_REG_31__SCAN_IN), .ZN(n2741) );
  INV_X2 U3476 ( .A(n2798), .ZN(n3703) );
  XNOR2_X1 U34770 ( .A(n4375), .B(n2915), .ZN(n2742) );
  AND2_X1 U3478 ( .A1(n3774), .A2(n4377), .ZN(n2939) );
  AND2_X1 U34790 ( .A1(n2939), .A2(n2850), .ZN(n4618) );
  INV_X1 U3480 ( .A(n4622), .ZN(n4294) );
  INV_X1 U34810 ( .A(n2862), .ZN(n2961) );
  INV_X1 U3482 ( .A(n3660), .ZN(n2745) );
  OR2_X1 U34830 ( .A1(n3793), .A2(n2904), .ZN(n3710) );
  NAND2_X1 U3484 ( .A1(n3793), .A2(n2904), .ZN(n3707) );
  NAND2_X1 U34850 ( .A1(n2900), .A2(n2898), .ZN(n2747) );
  INV_X1 U3486 ( .A(n3711), .ZN(n2748) );
  INV_X1 U34870 ( .A(n3047), .ZN(n3051) );
  AND2_X1 U3488 ( .A1(n3791), .A2(n3051), .ZN(n2992) );
  OR2_X1 U34890 ( .A1(n3791), .A2(n3051), .ZN(n3724) );
  NAND2_X1 U3490 ( .A1(n3790), .A2(n3081), .ZN(n3725) );
  NAND2_X1 U34910 ( .A1(n3083), .A2(n3725), .ZN(n2749) );
  OR2_X1 U3492 ( .A1(n3790), .A2(n3081), .ZN(n3717) );
  INV_X1 U34930 ( .A(n2750), .ZN(n2751) );
  OAI21_X1 U3494 ( .B1(n3057), .B2(n2751), .A(n3727), .ZN(n3117) );
  INV_X1 U34950 ( .A(n3156), .ZN(n3114) );
  OR2_X1 U3496 ( .A1(n3788), .A2(n3114), .ZN(n3721) );
  NAND2_X1 U34970 ( .A1(n3117), .A2(n3721), .ZN(n2752) );
  NAND2_X1 U3498 ( .A1(n3788), .A2(n3114), .ZN(n3726) );
  NAND2_X1 U34990 ( .A1(n2752), .A2(n3726), .ZN(n3094) );
  AND2_X1 U3500 ( .A1(n3787), .A2(n3196), .ZN(n3093) );
  OR2_X1 U35010 ( .A1(n3787), .A2(n3196), .ZN(n3722) );
  NAND2_X1 U3502 ( .A1(n3786), .A2(n3254), .ZN(n3736) );
  OR2_X1 U35030 ( .A1(n3786), .A2(n3254), .ZN(n3733) );
  NAND2_X1 U3504 ( .A1(n3784), .A2(n3296), .ZN(n3219) );
  NAND2_X1 U35050 ( .A1(n4218), .A2(n3229), .ZN(n2753) );
  NAND2_X1 U35060 ( .A1(n3219), .A2(n2753), .ZN(n2755) );
  INV_X1 U35070 ( .A(n3165), .ZN(n2754) );
  NOR2_X1 U35080 ( .A1(n2755), .A2(n2754), .ZN(n3737) );
  NAND2_X1 U35090 ( .A1(n3177), .A2(n3737), .ZN(n2759) );
  INV_X1 U35100 ( .A(n2755), .ZN(n2758) );
  OR2_X1 U35110 ( .A1(n3784), .A2(n3296), .ZN(n3221) );
  NAND2_X1 U35120 ( .A1(n3163), .A2(n3221), .ZN(n2757) );
  NOR2_X1 U35130 ( .A1(n4218), .A2(n3229), .ZN(n2756) );
  AOI21_X1 U35140 ( .B1(n2758), .B2(n2757), .A(n2756), .ZN(n3738) );
  NAND2_X1 U35150 ( .A1(n4221), .A2(n4222), .ZN(n4220) );
  OR2_X1 U35160 ( .A1(n4171), .A2(n4202), .ZN(n3673) );
  NAND2_X1 U35170 ( .A1(n4171), .A2(n4202), .ZN(n3672) );
  NAND2_X1 U35180 ( .A1(n3673), .A2(n3672), .ZN(n4191) );
  INV_X1 U35190 ( .A(n4190), .ZN(n2760) );
  NOR2_X1 U35200 ( .A1(n4191), .A2(n2760), .ZN(n2761) );
  NAND2_X1 U35210 ( .A1(n4220), .A2(n2761), .ZN(n2762) );
  NAND2_X1 U35220 ( .A1(n2762), .A2(n3672), .ZN(n4170) );
  NAND2_X1 U35230 ( .A1(n4170), .A2(n4180), .ZN(n2763) );
  AND2_X1 U35240 ( .A1(n4389), .A2(n4162), .ZN(n4096) );
  NAND2_X1 U35250 ( .A1(n4136), .A2(n4126), .ZN(n3640) );
  NAND2_X1 U35260 ( .A1(n4117), .A2(n3640), .ZN(n3749) );
  INV_X1 U35270 ( .A(n3749), .ZN(n4098) );
  INV_X1 U35280 ( .A(n2764), .ZN(n4118) );
  NAND2_X1 U35290 ( .A1(n4098), .A2(n4118), .ZN(n2765) );
  OR2_X1 U35300 ( .A1(n4136), .A2(n4126), .ZN(n3641) );
  NAND2_X1 U35310 ( .A1(n2765), .A2(n3641), .ZN(n4097) );
  OR2_X1 U35320 ( .A1(n4389), .A2(n4162), .ZN(n4095) );
  OAI22_X1 U35330 ( .A1(n3749), .A2(n4095), .B1(n3651), .B2(n4122), .ZN(n2766)
         );
  NOR2_X1 U35340 ( .A1(n4097), .A2(n2766), .ZN(n3676) );
  NAND2_X1 U35350 ( .A1(n4122), .A2(n3651), .ZN(n3754) );
  NAND2_X1 U35360 ( .A1(n4065), .A2(n3518), .ZN(n4038) );
  AND2_X1 U35370 ( .A1(n4041), .A2(n4038), .ZN(n3755) );
  AND2_X1 U35380 ( .A1(n4101), .A2(n4086), .ZN(n3756) );
  NAND2_X1 U35390 ( .A1(n4041), .A2(n3756), .ZN(n2769) );
  NAND2_X1 U35400 ( .A1(n4062), .A2(n4048), .ZN(n2767) );
  AND2_X1 U35410 ( .A1(n2768), .A2(n2767), .ZN(n3760) );
  AND2_X1 U35420 ( .A1(n2769), .A2(n3760), .ZN(n3681) );
  NAND2_X1 U35430 ( .A1(n2770), .A2(n3681), .ZN(n4019) );
  NAND2_X1 U35440 ( .A1(n4044), .A2(n3568), .ZN(n3642) );
  NAND2_X1 U35450 ( .A1(n4022), .A2(n3498), .ZN(n4018) );
  AND2_X1 U35460 ( .A1(n3642), .A2(n4018), .ZN(n3679) );
  NAND2_X1 U35470 ( .A1(n4024), .A2(n4010), .ZN(n3649) );
  NAND2_X1 U35480 ( .A1(n4004), .A2(n4027), .ZN(n3996) );
  NAND2_X1 U35490 ( .A1(n3649), .A2(n3996), .ZN(n3762) );
  NOR2_X1 U35500 ( .A1(n4002), .A2(n3988), .ZN(n3628) );
  NOR2_X1 U35510 ( .A1(n4024), .A2(n4010), .ZN(n3978) );
  NOR2_X1 U35520 ( .A1(n3628), .A2(n3978), .ZN(n3761) );
  INV_X1 U35530 ( .A(n3761), .ZN(n2771) );
  NAND2_X1 U35540 ( .A1(n4002), .A2(n3988), .ZN(n3766) );
  OR2_X1 U35550 ( .A1(n3983), .A2(n3971), .ZN(n3685) );
  NAND2_X1 U35560 ( .A1(n3983), .A2(n3971), .ZN(n3765) );
  NAND2_X1 U35570 ( .A1(n3685), .A2(n3765), .ZN(n3962) );
  XNOR2_X1 U35580 ( .A(n2818), .B(n3636), .ZN(n2783) );
  NAND2_X1 U35590 ( .A1(n4375), .A2(n4377), .ZN(n2773) );
  INV_X1 U35600 ( .A(n3774), .ZN(n4376) );
  NAND2_X1 U35610 ( .A1(n4376), .A2(n3703), .ZN(n2772) );
  OR2_X1 U35620 ( .A1(n2774), .A2(n2459), .ZN(n2775) );
  NAND2_X1 U35630 ( .A1(n4375), .A2(n3703), .ZN(n2853) );
  NAND2_X1 U35640 ( .A1(n3983), .A2(n4219), .ZN(n2781) );
  INV_X1 U35650 ( .A(REG2_REG_29__SCAN_IN), .ZN(n3959) );
  OR2_X1 U35660 ( .A1(n3953), .A2(n2493), .ZN(n2778) );
  AOI22_X1 U35670 ( .A1(n2776), .A2(REG0_REG_29__SCAN_IN), .B1(n2502), .B2(
        REG1_REG_29__SCAN_IN), .ZN(n2777) );
  OAI211_X1 U35680 ( .C1(n2779), .C2(n3959), .A(n2778), .B(n2777), .ZN(n3783)
         );
  INV_X1 U35690 ( .A(n2853), .ZN(n2844) );
  NAND2_X1 U35700 ( .A1(n4382), .A2(n2844), .ZN(n4216) );
  NAND2_X1 U35710 ( .A1(n3783), .A2(n4194), .ZN(n2780) );
  OAI211_X1 U35720 ( .C1(n3447), .C2(n4215), .A(n2781), .B(n2780), .ZN(n2782)
         );
  AOI21_X1 U35730 ( .B1(n2783), .B2(n4223), .A(n2782), .ZN(n3470) );
  OAI21_X1 U35740 ( .B1(n3475), .B2(n4294), .A(n3470), .ZN(n4248) );
  NOR2_X1 U35750 ( .A1(n2784), .A2(n2459), .ZN(n2787) );
  NAND2_X1 U35760 ( .A1(n2788), .A2(B_REG_SCAN_IN), .ZN(n2791) );
  NAND2_X1 U35770 ( .A1(n2796), .A2(n2797), .ZN(n2789) );
  XNOR2_X2 U35780 ( .A(n2790), .B(IR_REG_24__SCAN_IN), .ZN(n4374) );
  MUX2_X1 U35790 ( .A(n2791), .B(B_REG_SCAN_IN), .S(n4374), .Z(n2794) );
  INV_X1 U35800 ( .A(n3398), .ZN(n2808) );
  INV_X1 U35810 ( .A(D_REG_1__SCAN_IN), .ZN(n3403) );
  NAND2_X1 U3582 ( .A1(n2808), .A2(n3403), .ZN(n2911) );
  INV_X1 U3583 ( .A(n2795), .ZN(n3405) );
  NAND2_X1 U3584 ( .A1(n2788), .A2(n3405), .ZN(n2846) );
  NAND2_X1 U3585 ( .A1(n2911), .A2(n2846), .ZN(n2812) );
  NAND2_X1 U3586 ( .A1(n4618), .A2(n2798), .ZN(n2876) );
  AND2_X1 U3587 ( .A1(n3774), .A2(n3941), .ZN(n2851) );
  NAND2_X1 U3588 ( .A1(n2876), .A2(n2908), .ZN(n2799) );
  NOR2_X1 U3589 ( .A1(n3397), .A2(n2799), .ZN(n2811) );
  NOR4_X1 U3590 ( .A1(D_REG_8__SCAN_IN), .A2(D_REG_29__SCAN_IN), .A3(
        D_REG_25__SCAN_IN), .A4(D_REG_4__SCAN_IN), .ZN(n2803) );
  NOR4_X1 U3591 ( .A1(D_REG_11__SCAN_IN), .A2(D_REG_19__SCAN_IN), .A3(
        D_REG_14__SCAN_IN), .A4(D_REG_6__SCAN_IN), .ZN(n2802) );
  NOR4_X1 U3592 ( .A1(D_REG_3__SCAN_IN), .A2(D_REG_21__SCAN_IN), .A3(
        D_REG_23__SCAN_IN), .A4(D_REG_12__SCAN_IN), .ZN(n2801) );
  NOR4_X1 U3593 ( .A1(D_REG_27__SCAN_IN), .A2(D_REG_28__SCAN_IN), .A3(
        D_REG_10__SCAN_IN), .A4(D_REG_9__SCAN_IN), .ZN(n2800) );
  NAND4_X1 U3594 ( .A1(n2803), .A2(n2802), .A3(n2801), .A4(n2800), .ZN(n2810)
         );
  NOR2_X1 U3595 ( .A1(D_REG_26__SCAN_IN), .A2(D_REG_24__SCAN_IN), .ZN(n2807)
         );
  NOR4_X1 U3596 ( .A1(D_REG_7__SCAN_IN), .A2(D_REG_30__SCAN_IN), .A3(
        D_REG_5__SCAN_IN), .A4(D_REG_2__SCAN_IN), .ZN(n2806) );
  NOR4_X1 U3597 ( .A1(D_REG_15__SCAN_IN), .A2(D_REG_18__SCAN_IN), .A3(
        D_REG_17__SCAN_IN), .A4(D_REG_20__SCAN_IN), .ZN(n2805) );
  NOR4_X1 U3598 ( .A1(D_REG_22__SCAN_IN), .A2(D_REG_16__SCAN_IN), .A3(
        D_REG_31__SCAN_IN), .A4(D_REG_13__SCAN_IN), .ZN(n2804) );
  NAND4_X1 U3599 ( .A1(n2807), .A2(n2806), .A3(n2805), .A4(n2804), .ZN(n2809)
         );
  OAI21_X1 U3600 ( .B1(n2810), .B2(n2809), .A(n2808), .ZN(n2847) );
  NAND3_X1 U3601 ( .A1(n2812), .A2(n2811), .A3(n2847), .ZN(n2826) );
  INV_X1 U3602 ( .A(n2910), .ZN(n2848) );
  INV_X1 U3603 ( .A(n2813), .ZN(n2815) );
  NAND2_X1 U3604 ( .A1(n2965), .A2(n2961), .ZN(n2978) );
  NOR2_X1 U3605 ( .A1(n2978), .A2(n2977), .ZN(n2976) );
  NAND2_X1 U3606 ( .A1(n4230), .A2(n4229), .ZN(n4228) );
  OAI21_X1 U3607 ( .B1(n3969), .B2(n3447), .A(n2828), .ZN(n4251) );
  NAND2_X1 U3608 ( .A1(n2815), .A2(n2814), .ZN(U3514) );
  NAND2_X1 U3609 ( .A1(n2659), .A2(DATAI_29_), .ZN(n3691) );
  XNOR2_X1 U3610 ( .A(n3783), .B(n3691), .ZN(n3669) );
  INV_X1 U3611 ( .A(n2817), .ZN(n3687) );
  XNOR2_X1 U3612 ( .A(n2819), .B(n2278), .ZN(n2820) );
  INV_X1 U3613 ( .A(REG0_REG_30__SCAN_IN), .ZN(n2823) );
  NAND2_X1 U3614 ( .A1(n2218), .A2(REG2_REG_30__SCAN_IN), .ZN(n2822) );
  NAND2_X1 U3615 ( .A1(n2502), .A2(REG1_REG_30__SCAN_IN), .ZN(n2821) );
  OAI211_X1 U3616 ( .C1(n3632), .C2(n2823), .A(n2822), .B(n2821), .ZN(n3782)
         );
  XNOR2_X1 U3617 ( .A(n2824), .B(n2442), .ZN(n4406) );
  AOI21_X1 U3618 ( .B1(B_REG_SCAN_IN), .B2(n4406), .A(n4216), .ZN(n3946) );
  AOI22_X1 U3619 ( .A1(n3782), .A2(n3946), .B1(n4244), .B2(n2827), .ZN(n2825)
         );
  NAND2_X1 U3620 ( .A1(n2828), .A2(n2827), .ZN(n2829) );
  NAND2_X1 U3621 ( .A1(n2831), .A2(n2830), .ZN(U3547) );
  INV_X1 U3622 ( .A(REG0_REG_29__SCAN_IN), .ZN(n2832) );
  OR2_X2 U3623 ( .A1(n3011), .A2(n3400), .ZN(n3795) );
  INV_X1 U3624 ( .A(DATAI_21_), .ZN(n4917) );
  NAND2_X1 U3625 ( .A1(n3703), .A2(STATE_REG_SCAN_IN), .ZN(n2834) );
  OAI21_X1 U3626 ( .B1(STATE_REG_SCAN_IN), .B2(n4917), .A(n2834), .ZN(U3331)
         );
  INV_X1 U3627 ( .A(IR_REG_30__SCAN_IN), .ZN(n2836) );
  NAND3_X1 U3628 ( .A1(n2836), .A2(IR_REG_31__SCAN_IN), .A3(STATE_REG_SCAN_IN), 
        .ZN(n2837) );
  INV_X1 U3629 ( .A(DATAI_31_), .ZN(n4969) );
  OAI22_X1 U3630 ( .A1(n2835), .A2(n2837), .B1(STATE_REG_SCAN_IN), .B2(n4969), 
        .ZN(U3321) );
  INV_X1 U3631 ( .A(DATAI_29_), .ZN(n4921) );
  NAND2_X1 U3632 ( .A1(n2838), .A2(STATE_REG_SCAN_IN), .ZN(n2839) );
  OAI21_X1 U3633 ( .B1(STATE_REG_SCAN_IN), .B2(n4921), .A(n2839), .ZN(U3323)
         );
  INV_X1 U3634 ( .A(DATAI_25_), .ZN(n2841) );
  NAND2_X1 U3635 ( .A1(n3401), .A2(STATE_REG_SCAN_IN), .ZN(n2840) );
  OAI21_X1 U3636 ( .B1(STATE_REG_SCAN_IN), .B2(n2841), .A(n2840), .ZN(U3327)
         );
  INV_X1 U3637 ( .A(DATAI_27_), .ZN(n4767) );
  NAND2_X1 U3638 ( .A1(n4406), .A2(STATE_REG_SCAN_IN), .ZN(n2842) );
  OAI21_X1 U3639 ( .B1(STATE_REG_SCAN_IN), .B2(n4767), .A(n2842), .ZN(U3325)
         );
  INV_X1 U3640 ( .A(n3010), .ZN(n2843) );
  NAND2_X1 U3641 ( .A1(n2843), .A2(STATE_REG_SCAN_IN), .ZN(n3780) );
  NAND2_X1 U3642 ( .A1(n3397), .A2(n3780), .ZN(n3798) );
  NAND2_X1 U3643 ( .A1(n3010), .A2(n2844), .ZN(n2845) );
  NOR2_X1 U3644 ( .A1(n4541), .A2(U4043), .ZN(U3148) );
  AND2_X1 U3645 ( .A1(n2847), .A2(n2846), .ZN(n2913) );
  NAND3_X1 U3646 ( .A1(n2913), .A2(n2848), .A3(n2911), .ZN(n2892) );
  INV_X1 U3647 ( .A(n2915), .ZN(n2849) );
  OR2_X1 U3648 ( .A1(n2850), .A2(n4377), .ZN(n2882) );
  NAND2_X1 U3649 ( .A1(n2892), .A2(n2432), .ZN(n3014) );
  INV_X1 U3650 ( .A(n3014), .ZN(n2857) );
  INV_X1 U3651 ( .A(n2851), .ZN(n2852) );
  NAND2_X1 U3652 ( .A1(n2937), .A2(n2852), .ZN(n2854) );
  NAND2_X1 U3653 ( .A1(n2854), .A2(n2853), .ZN(n2871) );
  NAND2_X1 U3654 ( .A1(n4215), .A2(n2871), .ZN(n2855) );
  NAND2_X1 U3655 ( .A1(n2892), .A2(n2855), .ZN(n2856) );
  NAND2_X1 U3656 ( .A1(n2856), .A2(n2908), .ZN(n3013) );
  NOR3_X1 U3657 ( .A1(n2857), .A2(n3013), .A3(n3397), .ZN(n2958) );
  AND2_X4 U3658 ( .A1(n3011), .A2(n2915), .ZN(n3438) );
  INV_X1 U3659 ( .A(n4629), .ZN(n4606) );
  NAND2_X1 U3660 ( .A1(n3282), .A2(n2861), .ZN(n2860) );
  INV_X1 U3661 ( .A(n3011), .ZN(n2858) );
  NAND2_X1 U3662 ( .A1(n2860), .A2(n2859), .ZN(n2866) );
  INV_X1 U3663 ( .A(REG1_REG_0__SCAN_IN), .ZN(n2863) );
  NAND2_X1 U3664 ( .A1(n2862), .A2(n3438), .ZN(n2881) );
  OAI21_X1 U3665 ( .B1(n2863), .B2(n3011), .A(n2881), .ZN(n2864) );
  INV_X1 U3666 ( .A(n2869), .ZN(n2867) );
  NAND2_X1 U3667 ( .A1(n2867), .A2(n2866), .ZN(n2884) );
  AOI21_X1 U3668 ( .B1(n2870), .B2(n2869), .A(n2868), .ZN(n3818) );
  INV_X1 U3669 ( .A(n2892), .ZN(n2873) );
  NOR2_X1 U3670 ( .A1(n3397), .A2(n2871), .ZN(n2872) );
  NAND2_X1 U3671 ( .A1(n3818), .A2(n4396), .ZN(n2879) );
  NAND2_X1 U3672 ( .A1(n2432), .A2(n4382), .ZN(n2874) );
  OR2_X1 U3673 ( .A1(n3397), .A2(n4215), .ZN(n2875) );
  OR2_X1 U3674 ( .A1(n2892), .A2(n2875), .ZN(n2877) );
  AOI22_X1 U3675 ( .A1(n4390), .A2(n2887), .B1(n3621), .B2(n2862), .ZN(n2878)
         );
  OAI211_X1 U3676 ( .C1(n2958), .C2(n2880), .A(n2879), .B(n2878), .ZN(U3229)
         );
  INV_X1 U3677 ( .A(REG3_REG_1__SCAN_IN), .ZN(n2962) );
  NAND2_X1 U3678 ( .A1(n2881), .A2(n3431), .ZN(n2883) );
  AND2_X1 U3679 ( .A1(n2884), .A2(n2883), .ZN(n2889) );
  INV_X2 U3680 ( .A(n3431), .ZN(n3332) );
  NOR2_X1 U3681 ( .A1(n2965), .A2(n2943), .ZN(n2886) );
  AOI21_X1 U3682 ( .B1(n2887), .B2(n3282), .A(n2886), .ZN(n2947) );
  XNOR2_X1 U3683 ( .A(n2946), .B(n2947), .ZN(n2888) );
  NOR2_X1 U3684 ( .A1(n2889), .A2(n2888), .ZN(n2950) );
  AOI211_X1 U3685 ( .C1(n2889), .C2(n2888), .A(n3616), .B(n2950), .ZN(n2890)
         );
  INV_X1 U3686 ( .A(n2890), .ZN(n2897) );
  INV_X1 U3687 ( .A(n3796), .ZN(n2893) );
  INV_X1 U3688 ( .A(n4382), .ZN(n3814) );
  NAND2_X1 U3689 ( .A1(n2432), .A2(n3814), .ZN(n2891) );
  INV_X1 U3690 ( .A(n3794), .ZN(n3009) );
  OAI22_X1 U3691 ( .A1(n2893), .A2(n4384), .B1(n3009), .B2(n3610), .ZN(n2894)
         );
  AOI21_X1 U3692 ( .B1(n2895), .B2(n3621), .A(n2894), .ZN(n2896) );
  OAI211_X1 U3693 ( .C1(n2958), .C2(n2962), .A(n2897), .B(n2896), .ZN(U3219)
         );
  XNOR2_X1 U3694 ( .A(n2899), .B(n3661), .ZN(n2921) );
  XNOR2_X1 U3695 ( .A(n2900), .B(n3661), .ZN(n2903) );
  INV_X1 U3696 ( .A(n3792), .ZN(n3008) );
  OAI22_X1 U3697 ( .A1(n3008), .A2(n4216), .B1(n4215), .B2(n2904), .ZN(n2901)
         );
  AOI21_X1 U3698 ( .B1(n4219), .B2(n3794), .A(n2901), .ZN(n2902) );
  OAI21_X1 U3699 ( .B1(n2903), .B2(n4199), .A(n2902), .ZN(n2907) );
  AOI21_X1 U3700 ( .B1(n4622), .B2(n2921), .A(n2907), .ZN(n3028) );
  NOR2_X1 U3701 ( .A1(n2976), .A2(n2904), .ZN(n2905) );
  NOR2_X1 U3702 ( .A1(n2905), .A2(n2930), .ZN(n3026) );
  INV_X1 U3703 ( .A(n4371), .ZN(n3024) );
  AOI22_X1 U3704 ( .A1(n3026), .A2(n3024), .B1(REG0_REG_3__SCAN_IN), .B2(n4630), .ZN(n2906) );
  OAI21_X1 U3705 ( .B1(n3028), .B2(n4630), .A(n2906), .ZN(U3473) );
  INV_X1 U3706 ( .A(n2907), .ZN(n2923) );
  INV_X1 U3707 ( .A(n2908), .ZN(n2909) );
  NOR2_X1 U3708 ( .A1(n3397), .A2(n2909), .ZN(n2912) );
  NAND4_X1 U3709 ( .A1(n2913), .A2(n2912), .A3(n2911), .A4(n2910), .ZN(n2914)
         );
  INV_X2 U3710 ( .A(n4207), .ZN(n4564) );
  OR2_X1 U3711 ( .A1(n2915), .A2(n3941), .ZN(n2933) );
  NAND2_X1 U3712 ( .A1(n4227), .A2(n2933), .ZN(n2916) );
  INV_X1 U3713 ( .A(n3026), .ZN(n2919) );
  AND2_X1 U3714 ( .A1(n4629), .A2(n3941), .ZN(n2917) );
  AOI22_X1 U3715 ( .A1(n4564), .A2(REG2_REG_3__SCAN_IN), .B1(n4565), .B2(n3016), .ZN(n2918) );
  OAI21_X1 U3716 ( .B1(n2919), .B2(n4204), .A(n2918), .ZN(n2920) );
  AOI21_X1 U3717 ( .B1(n2921), .B2(n3951), .A(n2920), .ZN(n2922) );
  OAI21_X1 U3718 ( .B1(n2923), .B2(n4564), .A(n2922), .ZN(U3287) );
  XNOR2_X1 U3719 ( .A(n2924), .B(n3659), .ZN(n2932) );
  XOR2_X1 U3720 ( .A(n3659), .B(n2925), .Z(n2928) );
  INV_X1 U3721 ( .A(n3793), .ZN(n2954) );
  AOI22_X1 U3722 ( .A1(n3791), .A2(n4194), .B1(n3577), .B2(n4244), .ZN(n2926)
         );
  OAI21_X1 U3723 ( .B1(n2954), .B2(n4158), .A(n2926), .ZN(n2927) );
  AOI21_X1 U3724 ( .B1(n2928), .B2(n4223), .A(n2927), .ZN(n2929) );
  OAI21_X1 U3725 ( .B1(n4227), .B2(n2932), .A(n2929), .ZN(n4616) );
  OAI211_X1 U3726 ( .C1(n2930), .C2(n3040), .A(n4629), .B(n2994), .ZN(n4615)
         );
  OAI22_X1 U3727 ( .A1(n4615), .A2(n4377), .B1(n4231), .B2(n3578), .ZN(n2931)
         );
  OAI21_X1 U3728 ( .B1(n4616), .B2(n2931), .A(n4207), .ZN(n2936) );
  INV_X1 U3729 ( .A(n2932), .ZN(n4619) );
  INV_X1 U3730 ( .A(n2933), .ZN(n2934) );
  NAND2_X1 U3731 ( .A1(n4207), .A2(n2934), .ZN(n4237) );
  INV_X1 U3732 ( .A(n4237), .ZN(n4570) );
  AOI22_X1 U3733 ( .A1(n4619), .A2(n4570), .B1(REG2_REG_4__SCAN_IN), .B2(n4564), .ZN(n2935) );
  NAND2_X1 U3734 ( .A1(n2936), .A2(n2935), .ZN(U3286) );
  NAND2_X1 U3735 ( .A1(n3796), .A2(n2961), .ZN(n3702) );
  NAND2_X1 U3736 ( .A1(n3700), .A2(n3702), .ZN(n3652) );
  INV_X1 U3737 ( .A(n3652), .ZN(n4603) );
  NAND2_X1 U3738 ( .A1(n2862), .A2(n2937), .ZN(n4601) );
  NAND2_X1 U3739 ( .A1(n4227), .A2(n4199), .ZN(n2938) );
  AOI22_X1 U3740 ( .A1(n3652), .A2(n2938), .B1(n4194), .B2(n2887), .ZN(n4602)
         );
  OAI21_X1 U3741 ( .B1(n2939), .B2(n4601), .A(n4602), .ZN(n2940) );
  NAND2_X1 U3742 ( .A1(n2940), .A2(n4207), .ZN(n2942) );
  AOI22_X1 U3743 ( .A1(n4564), .A2(REG2_REG_0__SCAN_IN), .B1(
        REG3_REG_0__SCAN_IN), .B2(n4565), .ZN(n2941) );
  OAI211_X1 U3744 ( .C1(n4603), .C2(n4237), .A(n2942), .B(n2941), .ZN(U3290)
         );
  AOI22_X1 U3745 ( .A1(n3794), .A2(n3381), .B1(n2977), .B2(n3438), .ZN(n2944)
         );
  XNOR2_X1 U3746 ( .A(n2944), .B(n3332), .ZN(n3004) );
  INV_X1 U3747 ( .A(n2946), .ZN(n2949) );
  INV_X1 U3748 ( .A(n2947), .ZN(n2948) );
  NAND2_X1 U3749 ( .A1(n2953), .A2(n4396), .ZN(n2957) );
  OAI22_X1 U3750 ( .A1(n2954), .A2(n3610), .B1(n2483), .B2(n4384), .ZN(n2955)
         );
  AOI21_X1 U3751 ( .B1(n2977), .B2(n3621), .A(n2955), .ZN(n2956) );
  OAI211_X1 U3752 ( .C1(n2958), .C2(n2981), .A(n2957), .B(n2956), .ZN(U3234)
         );
  OAI21_X1 U3753 ( .B1(n2743), .B2(n2960), .A(n2959), .ZN(n4607) );
  INV_X1 U3754 ( .A(n4607), .ZN(n2972) );
  OAI21_X1 U3755 ( .B1(n2961), .B2(n2965), .A(n2978), .ZN(n4605) );
  OAI22_X1 U3756 ( .A1(n4204), .A2(n4605), .B1(n2962), .B2(n4231), .ZN(n2971)
         );
  NAND2_X1 U3757 ( .A1(n3796), .A2(n4219), .ZN(n2964) );
  NAND2_X1 U3758 ( .A1(n3794), .A2(n4194), .ZN(n2963) );
  OAI211_X1 U3759 ( .C1(n4215), .C2(n2965), .A(n2964), .B(n2963), .ZN(n2966)
         );
  INV_X1 U3760 ( .A(n2966), .ZN(n2969) );
  XNOR2_X1 U3761 ( .A(n2743), .B(n3700), .ZN(n2967) );
  NAND2_X1 U3762 ( .A1(n2967), .A2(n4223), .ZN(n2968) );
  OAI211_X1 U3763 ( .C1(n4607), .C2(n4227), .A(n2969), .B(n2968), .ZN(n4609)
         );
  MUX2_X1 U3764 ( .A(n4609), .B(REG2_REG_1__SCAN_IN), .S(n4564), .Z(n2970) );
  AOI211_X1 U3765 ( .C1(n2972), .C2(n4570), .A(n2971), .B(n2970), .ZN(n2973)
         );
  INV_X1 U3766 ( .A(n2973), .ZN(U3289) );
  OAI21_X1 U3767 ( .B1(n2975), .B2(n3660), .A(n2974), .ZN(n4611) );
  INV_X1 U3768 ( .A(n2976), .ZN(n2980) );
  NAND2_X1 U3769 ( .A1(n2978), .A2(n2977), .ZN(n2979) );
  NAND2_X1 U3770 ( .A1(n2980), .A2(n2979), .ZN(n4635) );
  OAI22_X1 U3771 ( .A1(n4635), .A2(n4204), .B1(n2981), .B2(n4231), .ZN(n2990)
         );
  INV_X1 U3772 ( .A(n4227), .ZN(n3213) );
  NAND2_X1 U3773 ( .A1(n4611), .A2(n3213), .ZN(n2987) );
  NAND2_X1 U3774 ( .A1(n2887), .A2(n4219), .ZN(n2983) );
  NAND2_X1 U3775 ( .A1(n3793), .A2(n4194), .ZN(n2982) );
  OAI211_X1 U3776 ( .C1(n4215), .C2(n2984), .A(n2983), .B(n2982), .ZN(n2985)
         );
  INV_X1 U3777 ( .A(n2985), .ZN(n2986) );
  OAI211_X1 U3778 ( .C1(n4199), .C2(n2988), .A(n2987), .B(n2986), .ZN(n4610)
         );
  MUX2_X1 U3779 ( .A(n4610), .B(REG2_REG_2__SCAN_IN), .S(n4564), .Z(n2989) );
  AOI211_X1 U3780 ( .C1(n4570), .C2(n4611), .A(n2990), .B(n2989), .ZN(n2991)
         );
  INV_X1 U3781 ( .A(n2991), .ZN(U3288) );
  INV_X1 U3782 ( .A(n2992), .ZN(n3713) );
  NAND2_X1 U3783 ( .A1(n3713), .A2(n3724), .ZN(n3657) );
  XOR2_X1 U3784 ( .A(n3657), .B(n2993), .Z(n3023) );
  INV_X1 U3785 ( .A(n3023), .ZN(n3002) );
  AOI21_X1 U3786 ( .B1(n3047), .B2(n2994), .A(n2254), .ZN(n3029) );
  INV_X1 U3787 ( .A(REG2_REG_5__SCAN_IN), .ZN(n3895) );
  OAI22_X1 U3788 ( .A1(n4207), .A2(n3895), .B1(n3055), .B2(n4231), .ZN(n2995)
         );
  AOI21_X1 U3789 ( .B1(n3029), .B2(n4569), .A(n2995), .ZN(n3001) );
  XOR2_X1 U3790 ( .A(n3657), .B(n2996), .Z(n2999) );
  INV_X1 U3791 ( .A(n3790), .ZN(n3071) );
  OAI22_X1 U3792 ( .A1(n3071), .A2(n4216), .B1(n4215), .B2(n3051), .ZN(n2997)
         );
  AOI21_X1 U3793 ( .B1(n4219), .B2(n3792), .A(n2997), .ZN(n2998) );
  OAI21_X1 U3794 ( .B1(n2999), .B2(n4199), .A(n2998), .ZN(n3022) );
  NAND2_X1 U3795 ( .A1(n3022), .A2(n4207), .ZN(n3000) );
  OAI211_X1 U3796 ( .C1(n3002), .C2(n4211), .A(n3001), .B(n3000), .ZN(U3285)
         );
  NAND2_X1 U3797 ( .A1(n3793), .A2(n3381), .ZN(n3006) );
  NAND2_X1 U3798 ( .A1(n3019), .A2(n3438), .ZN(n3005) );
  NAND2_X1 U3799 ( .A1(n3006), .A2(n3005), .ZN(n3007) );
  XNOR2_X1 U3800 ( .A(n3007), .B(n3332), .ZN(n3032) );
  AOI22_X1 U3801 ( .A1(n3793), .A2(n3282), .B1(n3381), .B2(n3019), .ZN(n3033)
         );
  XNOR2_X1 U3802 ( .A(n3032), .B(n3033), .ZN(n3035) );
  XOR2_X1 U3803 ( .A(n3036), .B(n3035), .Z(n3021) );
  OAI22_X1 U3804 ( .A1(n3009), .A2(n4384), .B1(n3008), .B2(n3610), .ZN(n3018)
         );
  NAND2_X1 U3805 ( .A1(n3011), .A2(n3010), .ZN(n3012) );
  OAI21_X1 U3806 ( .B1(n3013), .B2(n3012), .A(STATE_REG_SCAN_IN), .ZN(n3015)
         );
  INV_X1 U3807 ( .A(n4401), .ZN(n3614) );
  MUX2_X1 U3808 ( .A(U3149), .B(n3614), .S(n3016), .Z(n3017) );
  AOI211_X1 U3809 ( .C1(n3019), .C2(n3621), .A(n3018), .B(n3017), .ZN(n3020)
         );
  OAI21_X1 U3810 ( .B1(n3021), .B2(n3616), .A(n3020), .ZN(U3215) );
  AOI21_X1 U3811 ( .B1(n3023), .B2(n4622), .A(n3022), .ZN(n3031) );
  AOI22_X1 U3812 ( .A1(n3029), .A2(n3024), .B1(REG0_REG_5__SCAN_IN), .B2(n4630), .ZN(n3025) );
  OAI21_X1 U3813 ( .B1(n3031), .B2(n4630), .A(n3025), .ZN(U3477) );
  INV_X1 U3814 ( .A(n4309), .ZN(n4299) );
  AOI22_X1 U3815 ( .A1(n3026), .A2(n4299), .B1(REG1_REG_3__SCAN_IN), .B2(n4643), .ZN(n3027) );
  OAI21_X1 U3816 ( .B1(n3028), .B2(n4643), .A(n3027), .ZN(U3521) );
  AOI22_X1 U3817 ( .A1(n3029), .A2(n4299), .B1(REG1_REG_5__SCAN_IN), .B2(n4643), .ZN(n3030) );
  OAI21_X1 U3818 ( .B1(n3031), .B2(n4643), .A(n3030), .ZN(U3523) );
  INV_X1 U3819 ( .A(n3032), .ZN(n3034) );
  NAND2_X1 U3820 ( .A1(n3792), .A2(n3381), .ZN(n3038) );
  NAND2_X1 U3821 ( .A1(n3577), .A2(n3438), .ZN(n3037) );
  NAND2_X1 U3822 ( .A1(n3038), .A2(n3037), .ZN(n3039) );
  XNOR2_X1 U3823 ( .A(n3039), .B(n3332), .ZN(n3043) );
  NOR2_X1 U3825 ( .A1(n3040), .A2(n3448), .ZN(n3041) );
  AOI21_X1 U3826 ( .B1(n3792), .B2(n3042), .A(n3041), .ZN(n3044) );
  XNOR2_X1 U3827 ( .A(n3043), .B(n3044), .ZN(n3575) );
  NAND2_X1 U3828 ( .A1(n3576), .A2(n3575), .ZN(n3574) );
  INV_X1 U3829 ( .A(n3043), .ZN(n3045) );
  NAND2_X1 U3830 ( .A1(n3574), .A2(n2235), .ZN(n3050) );
  NOR2_X1 U3831 ( .A1(n3051), .A2(n3448), .ZN(n3046) );
  AOI21_X1 U3832 ( .B1(n3791), .B2(n3042), .A(n3046), .ZN(n3066) );
  AOI22_X1 U3833 ( .A1(n3791), .A2(n3381), .B1(n3438), .B2(n3047), .ZN(n3048)
         );
  XNOR2_X1 U3834 ( .A(n3048), .B(n3332), .ZN(n3067) );
  XOR2_X1 U3835 ( .A(n3066), .B(n3067), .Z(n3049) );
  NAND2_X1 U3836 ( .A1(n3050), .A2(n3049), .ZN(n3069) );
  OAI211_X1 U3837 ( .C1(n3050), .C2(n3049), .A(n3069), .B(n4396), .ZN(n3054)
         );
  INV_X1 U3838 ( .A(REG3_REG_5__SCAN_IN), .ZN(n4780) );
  NOR2_X1 U3839 ( .A1(STATE_REG_SCAN_IN), .A2(n4780), .ZN(n4415) );
  INV_X1 U3840 ( .A(n3621), .ZN(n4387) );
  OAI22_X1 U3841 ( .A1(n4387), .A2(n3051), .B1(n3071), .B2(n3610), .ZN(n3052)
         );
  AOI211_X1 U3842 ( .C1(n3622), .C2(n3792), .A(n4415), .B(n3052), .ZN(n3053)
         );
  OAI211_X1 U3843 ( .C1(n4401), .C2(n3055), .A(n3054), .B(n3053), .ZN(U3224)
         );
  AOI21_X1 U3844 ( .B1(n3080), .B2(n3133), .A(n4606), .ZN(n3056) );
  AND2_X1 U3845 ( .A1(n3056), .A2(n3112), .ZN(n4621) );
  XNOR2_X1 U3846 ( .A(n3057), .B(n3716), .ZN(n3061) );
  NOR2_X1 U3847 ( .A1(n3128), .A2(n4215), .ZN(n3058) );
  AOI21_X1 U3848 ( .B1(n3788), .B2(n4194), .A(n3058), .ZN(n3060) );
  NAND2_X1 U3849 ( .A1(n3790), .A2(n4219), .ZN(n3059) );
  OAI211_X1 U3850 ( .C1(n3061), .C2(n4199), .A(n3060), .B(n3059), .ZN(n4620)
         );
  AOI21_X1 U3851 ( .B1(n4621), .B2(n3941), .A(n4620), .ZN(n3065) );
  XOR2_X1 U3852 ( .A(n3062), .B(n3716), .Z(n4623) );
  INV_X1 U3853 ( .A(REG2_REG_7__SCAN_IN), .ZN(n3894) );
  OAI22_X1 U3854 ( .A1(n4207), .A2(n3894), .B1(n3136), .B2(n4231), .ZN(n3063)
         );
  AOI21_X1 U3855 ( .B1(n4623), .B2(n3951), .A(n3063), .ZN(n3064) );
  OAI21_X1 U3856 ( .B1(n3065), .B2(n4564), .A(n3064), .ZN(U3283) );
  OR2_X1 U3857 ( .A1(n3067), .A2(n3066), .ZN(n3068) );
  AOI22_X1 U3858 ( .A1(n3790), .A2(n3381), .B1(n3438), .B2(n3084), .ZN(n3070)
         );
  XOR2_X1 U3859 ( .A(n3332), .B(n3070), .Z(n3130) );
  INV_X1 U3860 ( .A(n3282), .ZN(n3445) );
  OAI22_X1 U3861 ( .A1(n3071), .A2(n3445), .B1(n3448), .B2(n3081), .ZN(n3131)
         );
  XNOR2_X1 U3862 ( .A(n3130), .B(n3131), .ZN(n3072) );
  XNOR2_X1 U3863 ( .A(n3132), .B(n3072), .ZN(n3078) );
  NOR2_X1 U3864 ( .A1(STATE_REG_SCAN_IN), .A2(n3073), .ZN(n4426) );
  AOI21_X1 U3865 ( .B1(n4390), .B2(n3789), .A(n4426), .ZN(n3075) );
  AOI22_X1 U3866 ( .A1(n3622), .A2(n3791), .B1(n3621), .B2(n3084), .ZN(n3074)
         );
  OAI211_X1 U3867 ( .C1(n4401), .C2(n3076), .A(n3075), .B(n3074), .ZN(n3077)
         );
  AOI21_X1 U3868 ( .B1(n3078), .B2(n4396), .A(n3077), .ZN(n3079) );
  INV_X1 U3869 ( .A(n3079), .ZN(U3236) );
  OAI21_X1 U3870 ( .B1(n2254), .B2(n3081), .A(n3080), .ZN(n4567) );
  NAND2_X1 U3871 ( .A1(n3717), .A2(n3725), .ZN(n3654) );
  XNOR2_X1 U3872 ( .A(n3082), .B(n3654), .ZN(n4571) );
  XNOR2_X1 U3873 ( .A(n3083), .B(n3654), .ZN(n3087) );
  AOI22_X1 U3874 ( .A1(n3791), .A2(n4219), .B1(n3084), .B2(n4244), .ZN(n3086)
         );
  NAND2_X1 U3875 ( .A1(n3789), .A2(n4194), .ZN(n3085) );
  OAI211_X1 U3876 ( .C1(n3087), .C2(n4199), .A(n3086), .B(n3085), .ZN(n3088)
         );
  AOI21_X1 U3877 ( .B1(n3213), .B2(n4571), .A(n3088), .ZN(n4574) );
  INV_X1 U3878 ( .A(n4574), .ZN(n3089) );
  AOI21_X1 U3879 ( .B1(n4618), .B2(n4571), .A(n3089), .ZN(n3091) );
  MUX2_X1 U3880 ( .A(n2536), .B(n3091), .S(n4631), .Z(n3090) );
  OAI21_X1 U3881 ( .B1(n4567), .B2(n4371), .A(n3090), .ZN(U3479) );
  INV_X1 U3882 ( .A(REG1_REG_6__SCAN_IN), .ZN(n4425) );
  MUX2_X1 U3883 ( .A(n4425), .B(n3091), .S(n4646), .Z(n3092) );
  OAI21_X1 U3884 ( .B1(n4567), .B2(n4309), .A(n3092), .ZN(U3524) );
  INV_X1 U3885 ( .A(n3093), .ZN(n3734) );
  NAND2_X1 U3886 ( .A1(n3734), .A2(n3722), .ZN(n3658) );
  XOR2_X1 U3887 ( .A(n3658), .B(n3094), .Z(n3097) );
  AOI22_X1 U3888 ( .A1(n3786), .A2(n4194), .B1(n4244), .B2(n3197), .ZN(n3096)
         );
  NAND2_X1 U3889 ( .A1(n3788), .A2(n4219), .ZN(n3095) );
  OAI211_X1 U3890 ( .C1(n3097), .C2(n4199), .A(n3096), .B(n3095), .ZN(n3104)
         );
  INV_X1 U3891 ( .A(n3104), .ZN(n3103) );
  XNOR2_X1 U3892 ( .A(n3098), .B(n3658), .ZN(n3105) );
  INV_X1 U3893 ( .A(REG2_REG_9__SCAN_IN), .ZN(n3892) );
  OAI22_X1 U3894 ( .A1(n3200), .A2(n4231), .B1(n3892), .B2(n4207), .ZN(n3101)
         );
  AND2_X1 U3895 ( .A1(n3113), .A2(n3197), .ZN(n3099) );
  OR2_X1 U3896 ( .A1(n3099), .A2(n3205), .ZN(n3111) );
  NOR2_X1 U3897 ( .A1(n3111), .A2(n4204), .ZN(n3100) );
  AOI211_X1 U3898 ( .C1(n3105), .C2(n3951), .A(n3101), .B(n3100), .ZN(n3102)
         );
  OAI21_X1 U3899 ( .B1(n3103), .B2(n4564), .A(n3102), .ZN(U3281) );
  AOI21_X1 U3900 ( .B1(n4622), .B2(n3105), .A(n3104), .ZN(n3108) );
  MUX2_X1 U3901 ( .A(n3106), .B(n3108), .S(n4631), .Z(n3107) );
  OAI21_X1 U3902 ( .B1(n3111), .B2(n4371), .A(n3107), .ZN(U3485) );
  INV_X1 U3903 ( .A(REG1_REG_9__SCAN_IN), .ZN(n3109) );
  MUX2_X1 U3904 ( .A(n3109), .B(n3108), .S(n4646), .Z(n3110) );
  OAI21_X1 U3905 ( .B1(n4309), .B2(n3111), .A(n3110), .ZN(U3527) );
  INV_X1 U3906 ( .A(n3112), .ZN(n3115) );
  OAI21_X1 U3907 ( .B1(n3115), .B2(n3114), .A(n3113), .ZN(n4558) );
  NAND2_X1 U3908 ( .A1(n3721), .A2(n3726), .ZN(n3655) );
  XOR2_X1 U3909 ( .A(n3116), .B(n3655), .Z(n4560) );
  XNOR2_X1 U3910 ( .A(n3117), .B(n3655), .ZN(n3118) );
  NAND2_X1 U3911 ( .A1(n3118), .A2(n4223), .ZN(n3120) );
  AOI22_X1 U3912 ( .A1(n3789), .A2(n4219), .B1(n3156), .B2(n4244), .ZN(n3119)
         );
  OAI211_X1 U3913 ( .C1(n3208), .C2(n4216), .A(n3120), .B(n3119), .ZN(n3121)
         );
  AOI21_X1 U3914 ( .B1(n4560), .B2(n3213), .A(n3121), .ZN(n4563) );
  INV_X1 U3915 ( .A(n4563), .ZN(n3122) );
  AOI21_X1 U3916 ( .B1(n4618), .B2(n4560), .A(n3122), .ZN(n3124) );
  MUX2_X1 U3917 ( .A(n2556), .B(n3124), .S(n4631), .Z(n3123) );
  OAI21_X1 U3918 ( .B1(n4558), .B2(n4371), .A(n3123), .ZN(U3483) );
  INV_X1 U3919 ( .A(REG1_REG_8__SCAN_IN), .ZN(n3125) );
  MUX2_X1 U3920 ( .A(n3125), .B(n3124), .S(n4646), .Z(n3126) );
  OAI21_X1 U3921 ( .B1(n4558), .B2(n4309), .A(n3126), .ZN(U3526) );
  AOI22_X1 U3922 ( .A1(n3789), .A2(n3381), .B1(n3438), .B2(n3133), .ZN(n3127)
         );
  XNOR2_X1 U3923 ( .A(n3127), .B(n3332), .ZN(n3150) );
  NOR2_X1 U3924 ( .A1(n3128), .A2(n3448), .ZN(n3129) );
  AOI21_X1 U3925 ( .B1(n3789), .B2(n3282), .A(n3129), .ZN(n3149) );
  XOR2_X1 U3926 ( .A(n3150), .B(n3149), .Z(n3152) );
  XOR2_X1 U3927 ( .A(n3152), .B(n3153), .Z(n3138) );
  INV_X1 U3928 ( .A(REG3_REG_7__SCAN_IN), .ZN(n4789) );
  NOR2_X1 U3929 ( .A1(STATE_REG_SCAN_IN), .A2(n4789), .ZN(n4436) );
  AOI21_X1 U3930 ( .B1(n4390), .B2(n3788), .A(n4436), .ZN(n3135) );
  AOI22_X1 U3931 ( .A1(n3622), .A2(n3790), .B1(n3621), .B2(n3133), .ZN(n3134)
         );
  OAI211_X1 U3932 ( .C1(n4401), .C2(n3136), .A(n3135), .B(n3134), .ZN(n3137)
         );
  AOI21_X1 U3933 ( .B1(n3138), .B2(n4396), .A(n3137), .ZN(n3139) );
  INV_X1 U3934 ( .A(n3139), .ZN(U3210) );
  NAND2_X1 U3935 ( .A1(n3788), .A2(n3381), .ZN(n3141) );
  NAND2_X1 U3936 ( .A1(n3156), .A2(n3438), .ZN(n3140) );
  NAND2_X1 U3937 ( .A1(n3141), .A2(n3140), .ZN(n3142) );
  XNOR2_X1 U3938 ( .A(n3142), .B(n3332), .ZN(n3145) );
  NAND2_X1 U3939 ( .A1(n3788), .A2(n3042), .ZN(n3144) );
  NAND2_X1 U3940 ( .A1(n3156), .A2(n3381), .ZN(n3143) );
  NAND2_X1 U3941 ( .A1(n3144), .A2(n3143), .ZN(n3146) );
  NAND2_X1 U3942 ( .A1(n3145), .A2(n3146), .ZN(n3189) );
  INV_X1 U3943 ( .A(n3145), .ZN(n3148) );
  INV_X1 U3944 ( .A(n3146), .ZN(n3147) );
  NAND2_X1 U3945 ( .A1(n3148), .A2(n3147), .ZN(n3191) );
  NAND2_X1 U3946 ( .A1(n3189), .A2(n3191), .ZN(n3154) );
  NOR2_X1 U3947 ( .A1(n3150), .A2(n3149), .ZN(n3151) );
  XOR2_X1 U3948 ( .A(n3154), .B(n3190), .Z(n3161) );
  NAND2_X1 U3949 ( .A1(REG3_REG_8__SCAN_IN), .A2(U3149), .ZN(n4446) );
  INV_X1 U3950 ( .A(n4446), .ZN(n3155) );
  AOI21_X1 U3951 ( .B1(n4390), .B2(n3787), .A(n3155), .ZN(n3158) );
  AOI22_X1 U3952 ( .A1(n3622), .A2(n3789), .B1(n3621), .B2(n3156), .ZN(n3157)
         );
  OAI211_X1 U3953 ( .C1(n4401), .C2(n3159), .A(n3158), .B(n3157), .ZN(n3160)
         );
  AOI21_X1 U3954 ( .B1(n3161), .B2(n4396), .A(n3160), .ZN(n3162) );
  INV_X1 U3955 ( .A(n3162), .ZN(U3218) );
  NAND2_X1 U3956 ( .A1(n3221), .A2(n3219), .ZN(n3644) );
  INV_X1 U3957 ( .A(n3163), .ZN(n3164) );
  AOI21_X1 U3958 ( .B1(n3177), .B2(n3165), .A(n3164), .ZN(n3222) );
  XOR2_X1 U3959 ( .A(n3644), .B(n3222), .Z(n3169) );
  NOR2_X1 U3960 ( .A1(n3296), .A2(n4215), .ZN(n3166) );
  AOI21_X1 U3961 ( .B1(n4218), .B2(n4194), .A(n3166), .ZN(n3168) );
  NAND2_X1 U3962 ( .A1(n3785), .A2(n4219), .ZN(n3167) );
  OAI211_X1 U3963 ( .C1(n3169), .C2(n4199), .A(n3168), .B(n3167), .ZN(n3237)
         );
  INV_X1 U3964 ( .A(n3237), .ZN(n3175) );
  XNOR2_X1 U3965 ( .A(n3170), .B(n3644), .ZN(n3238) );
  OAI21_X1 U3966 ( .B1(n2229), .B2(n3296), .A(n2326), .ZN(n3243) );
  NOR2_X1 U3967 ( .A1(n3243), .A2(n4204), .ZN(n3173) );
  INV_X1 U3968 ( .A(REG2_REG_12__SCAN_IN), .ZN(n3171) );
  OAI22_X1 U3969 ( .A1(n4207), .A2(n3171), .B1(n3537), .B2(n4231), .ZN(n3172)
         );
  AOI211_X1 U3970 ( .C1(n3238), .C2(n3951), .A(n3173), .B(n3172), .ZN(n3174)
         );
  OAI21_X1 U3971 ( .B1(n3175), .B2(n4564), .A(n3174), .ZN(U3278) );
  XNOR2_X1 U3972 ( .A(n3176), .B(n3656), .ZN(n3178) );
  INV_X1 U3973 ( .A(n3178), .ZN(n4625) );
  XNOR2_X1 U3974 ( .A(n3177), .B(n3656), .ZN(n3184) );
  NAND2_X1 U3975 ( .A1(n3178), .A2(n3213), .ZN(n3183) );
  OAI22_X1 U3976 ( .A1(n3180), .A2(n4216), .B1(n4215), .B2(n3179), .ZN(n3181)
         );
  AOI21_X1 U3977 ( .B1(n4219), .B2(n3786), .A(n3181), .ZN(n3182) );
  OAI211_X1 U3978 ( .C1(n4199), .C2(n3184), .A(n3183), .B(n3182), .ZN(n4626)
         );
  NAND2_X1 U3979 ( .A1(n4626), .A2(n4207), .ZN(n3188) );
  AOI21_X1 U3980 ( .B1(n3286), .B2(n3204), .A(n2229), .ZN(n4628) );
  INV_X1 U3981 ( .A(REG2_REG_11__SCAN_IN), .ZN(n3185) );
  OAI22_X1 U3982 ( .A1(n4207), .A2(n3185), .B1(n3289), .B2(n4231), .ZN(n3186)
         );
  AOI21_X1 U3983 ( .B1(n4628), .B2(n4569), .A(n3186), .ZN(n3187) );
  OAI211_X1 U3984 ( .C1(n4625), .C2(n4237), .A(n3188), .B(n3187), .ZN(U3279)
         );
  NAND2_X1 U3985 ( .A1(n3190), .A2(n3189), .ZN(n3192) );
  NAND2_X1 U3986 ( .A1(n3192), .A2(n3191), .ZN(n3257) );
  NAND2_X1 U3987 ( .A1(n3787), .A2(n3381), .ZN(n3194) );
  NAND2_X1 U3988 ( .A1(n3197), .A2(n3438), .ZN(n3193) );
  NAND2_X1 U3989 ( .A1(n3194), .A2(n3193), .ZN(n3195) );
  XNOR2_X1 U3990 ( .A(n3195), .B(n3332), .ZN(n3258) );
  OAI22_X1 U3991 ( .A1(n3208), .A2(n3445), .B1(n3448), .B2(n3196), .ZN(n3259)
         );
  XOR2_X1 U3992 ( .A(n3258), .B(n3259), .Z(n3256) );
  XNOR2_X1 U3993 ( .A(n3257), .B(n3256), .ZN(n3202) );
  AND2_X1 U3994 ( .A1(U3149), .A2(REG3_REG_9__SCAN_IN), .ZN(n4462) );
  AOI21_X1 U3995 ( .B1(n4390), .B2(n3786), .A(n4462), .ZN(n3199) );
  AOI22_X1 U3996 ( .A1(n3622), .A2(n3788), .B1(n3621), .B2(n3197), .ZN(n3198)
         );
  OAI211_X1 U3997 ( .C1(n4401), .C2(n3200), .A(n3199), .B(n3198), .ZN(n3201)
         );
  AOI21_X1 U3998 ( .B1(n3202), .B2(n4396), .A(n3201), .ZN(n3203) );
  INV_X1 U3999 ( .A(n3203), .ZN(U3228) );
  OAI21_X1 U4000 ( .B1(n3205), .B2(n3254), .A(n3204), .ZN(n4551) );
  INV_X1 U4001 ( .A(REG1_REG_10__SCAN_IN), .ZN(n3215) );
  NAND2_X1 U4002 ( .A1(n3733), .A2(n3736), .ZN(n3643) );
  XOR2_X1 U4003 ( .A(n3643), .B(n3206), .Z(n4553) );
  XNOR2_X1 U4004 ( .A(n3207), .B(n3643), .ZN(n3211) );
  OAI22_X1 U4005 ( .A1(n3208), .A2(n4158), .B1(n3254), .B2(n4215), .ZN(n3209)
         );
  AOI21_X1 U4006 ( .B1(n4194), .B2(n3785), .A(n3209), .ZN(n3210) );
  OAI21_X1 U4007 ( .B1(n3211), .B2(n4199), .A(n3210), .ZN(n3212) );
  AOI21_X1 U4008 ( .B1(n4553), .B2(n3213), .A(n3212), .ZN(n4556) );
  INV_X1 U4009 ( .A(n4556), .ZN(n3214) );
  AOI21_X1 U4010 ( .B1(n4618), .B2(n4553), .A(n3214), .ZN(n3217) );
  MUX2_X1 U4011 ( .A(n3215), .B(n3217), .S(n4646), .Z(n3216) );
  OAI21_X1 U4012 ( .B1(n4551), .B2(n4309), .A(n3216), .ZN(U3528) );
  MUX2_X1 U4013 ( .A(n2582), .B(n3217), .S(n4631), .Z(n3218) );
  OAI21_X1 U4014 ( .B1(n4551), .B2(n4371), .A(n3218), .ZN(U3487) );
  INV_X1 U4015 ( .A(n3219), .ZN(n3220) );
  AOI21_X1 U4016 ( .B1(n3222), .B2(n3221), .A(n3220), .ZN(n3224) );
  AND2_X1 U4017 ( .A1(n3223), .A2(n4186), .ZN(n3645) );
  XNOR2_X1 U4018 ( .A(n3224), .B(n3645), .ZN(n3227) );
  AOI22_X1 U4019 ( .A1(n4196), .A2(n4194), .B1(n4244), .B2(n3308), .ZN(n3226)
         );
  NAND2_X1 U4020 ( .A1(n3784), .A2(n4219), .ZN(n3225) );
  OAI211_X1 U4021 ( .C1(n3227), .C2(n4199), .A(n3226), .B(n3225), .ZN(n3244)
         );
  INV_X1 U4022 ( .A(n3244), .ZN(n3236) );
  XOR2_X1 U4023 ( .A(n3645), .B(n3228), .Z(n3245) );
  NOR2_X1 U4024 ( .A1(n3230), .A2(n3229), .ZN(n3231) );
  NOR2_X1 U4025 ( .A1(n3250), .A2(n4204), .ZN(n3234) );
  INV_X1 U4026 ( .A(REG2_REG_13__SCAN_IN), .ZN(n3232) );
  OAI22_X1 U4027 ( .A1(n4207), .A2(n3232), .B1(n3311), .B2(n4231), .ZN(n3233)
         );
  AOI211_X1 U4028 ( .C1(n3245), .C2(n3951), .A(n3234), .B(n3233), .ZN(n3235)
         );
  OAI21_X1 U4029 ( .B1(n4564), .B2(n3236), .A(n3235), .ZN(U3277) );
  INV_X1 U4030 ( .A(REG1_REG_12__SCAN_IN), .ZN(n3239) );
  AOI21_X1 U4031 ( .B1(n4622), .B2(n3238), .A(n3237), .ZN(n3241) );
  MUX2_X1 U4032 ( .A(n3239), .B(n3241), .S(n4646), .Z(n3240) );
  OAI21_X1 U4033 ( .B1(n3243), .B2(n4309), .A(n3240), .ZN(U3530) );
  MUX2_X1 U4034 ( .A(n2602), .B(n3241), .S(n4631), .Z(n3242) );
  OAI21_X1 U4035 ( .B1(n3243), .B2(n4371), .A(n3242), .ZN(U3491) );
  AOI21_X1 U4036 ( .B1(n3245), .B2(n4622), .A(n3244), .ZN(n3247) );
  MUX2_X1 U4037 ( .A(n3866), .B(n3247), .S(n4646), .Z(n3246) );
  OAI21_X1 U4038 ( .B1(n4309), .B2(n3250), .A(n3246), .ZN(U3531) );
  MUX2_X1 U4039 ( .A(n3248), .B(n3247), .S(n4631), .Z(n3249) );
  OAI21_X1 U4040 ( .B1(n3250), .B2(n4371), .A(n3249), .ZN(U3493) );
  NAND2_X1 U4041 ( .A1(n3786), .A2(n3381), .ZN(n3252) );
  NAND2_X1 U4042 ( .A1(n3269), .A2(n3438), .ZN(n3251) );
  NAND2_X1 U40430 ( .A1(n3252), .A2(n3251), .ZN(n3253) );
  XNOR2_X1 U4044 ( .A(n3253), .B(n3332), .ZN(n3276) );
  NOR2_X1 U4045 ( .A1(n3254), .A2(n3448), .ZN(n3255) );
  AOI21_X1 U4046 ( .B1(n3786), .B2(n3282), .A(n3255), .ZN(n3274) );
  XOR2_X1 U4047 ( .A(n3276), .B(n3274), .Z(n3267) );
  NAND2_X1 U4048 ( .A1(n3257), .A2(n3256), .ZN(n3263) );
  INV_X1 U4049 ( .A(n3258), .ZN(n3261) );
  NAND2_X1 U4050 ( .A1(n3261), .A2(n3260), .ZN(n3262) );
  NAND2_X1 U4051 ( .A1(n3263), .A2(n3262), .ZN(n3266) );
  INV_X1 U4052 ( .A(n3266), .ZN(n3265) );
  NAND2_X1 U4053 ( .A1(n3265), .A2(n3264), .ZN(n3278) );
  AOI211_X1 U4054 ( .C1(n3267), .C2(n3266), .A(n3616), .B(n2385), .ZN(n3273)
         );
  NAND2_X1 U4055 ( .A1(REG3_REG_10__SCAN_IN), .A2(U3149), .ZN(n4467) );
  INV_X1 U4056 ( .A(n4467), .ZN(n3268) );
  AOI21_X1 U4057 ( .B1(n3622), .B2(n3787), .A(n3268), .ZN(n3271) );
  AOI22_X1 U4058 ( .A1(n4390), .A2(n3785), .B1(n3621), .B2(n3269), .ZN(n3270)
         );
  OAI211_X1 U4059 ( .C1(n4401), .C2(n4549), .A(n3271), .B(n3270), .ZN(n3272)
         );
  OR2_X1 U4060 ( .A1(n3273), .A2(n3272), .ZN(U3214) );
  INV_X1 U4061 ( .A(n3274), .ZN(n3275) );
  NAND2_X1 U4062 ( .A1(n3276), .A2(n3275), .ZN(n3277) );
  NAND2_X1 U4063 ( .A1(n3785), .A2(n3381), .ZN(n3280) );
  NAND2_X1 U4064 ( .A1(n3286), .A2(n3438), .ZN(n3279) );
  NAND2_X1 U4065 ( .A1(n3280), .A2(n3279), .ZN(n3281) );
  XNOR2_X1 U4066 ( .A(n3281), .B(n3332), .ZN(n3525) );
  NAND2_X1 U4067 ( .A1(n3785), .A2(n3042), .ZN(n3284) );
  NAND2_X1 U4068 ( .A1(n3286), .A2(n3381), .ZN(n3283) );
  NAND2_X1 U4069 ( .A1(n3284), .A2(n3283), .ZN(n3527) );
  INV_X1 U4070 ( .A(n3527), .ZN(n3524) );
  XNOR2_X1 U4071 ( .A(n3525), .B(n3524), .ZN(n3285) );
  XNOR2_X1 U4072 ( .A(n3299), .B(n3285), .ZN(n3291) );
  AND2_X1 U4073 ( .A1(U3149), .A2(REG3_REG_11__SCAN_IN), .ZN(n4483) );
  AOI21_X1 U4074 ( .B1(n3622), .B2(n3786), .A(n4483), .ZN(n3288) );
  AOI22_X1 U4075 ( .A1(n4390), .A2(n3784), .B1(n3621), .B2(n3286), .ZN(n3287)
         );
  OAI211_X1 U4076 ( .C1(n4401), .C2(n3289), .A(n3288), .B(n3287), .ZN(n3290)
         );
  AOI21_X1 U4077 ( .B1(n3291), .B2(n4396), .A(n3290), .ZN(n3292) );
  INV_X1 U4078 ( .A(n3292), .ZN(U3233) );
  NAND2_X1 U4079 ( .A1(n3784), .A2(n3381), .ZN(n3294) );
  NAND2_X1 U4080 ( .A1(n3534), .A2(n3438), .ZN(n3293) );
  NAND2_X1 U4081 ( .A1(n3294), .A2(n3293), .ZN(n3295) );
  XNOR2_X1 U4082 ( .A(n3295), .B(n3431), .ZN(n3300) );
  NOR2_X1 U4083 ( .A1(n3296), .A2(n3448), .ZN(n3297) );
  AOI21_X1 U4084 ( .B1(n3784), .B2(n3042), .A(n3297), .ZN(n3301) );
  NOR2_X1 U4085 ( .A1(n3300), .A2(n3301), .ZN(n3530) );
  AOI21_X1 U4086 ( .B1(n3527), .B2(n3525), .A(n3530), .ZN(n3298) );
  NOR3_X1 U4087 ( .A1(n3530), .A2(n3527), .A3(n3525), .ZN(n3304) );
  INV_X1 U4088 ( .A(n3300), .ZN(n3303) );
  INV_X1 U4089 ( .A(n3301), .ZN(n3302) );
  NOR2_X1 U4090 ( .A1(n3303), .A2(n3302), .ZN(n3529) );
  NOR2_X1 U4091 ( .A1(n3304), .A2(n3529), .ZN(n3305) );
  AOI22_X1 U4092 ( .A1(n4218), .A2(n3042), .B1(n3381), .B2(n3308), .ZN(n3317)
         );
  AOI22_X1 U4093 ( .A1(n4218), .A2(n3381), .B1(n3438), .B2(n3308), .ZN(n3306)
         );
  XNOR2_X1 U4094 ( .A(n3306), .B(n3332), .ZN(n3321) );
  XOR2_X1 U4095 ( .A(n3317), .B(n3321), .Z(n3307) );
  XNOR2_X1 U4096 ( .A(n3320), .B(n3307), .ZN(n3313) );
  NOR2_X1 U4097 ( .A1(STATE_REG_SCAN_IN), .A2(n2613), .ZN(n4501) );
  AOI21_X1 U4098 ( .B1(n3622), .B2(n3784), .A(n4501), .ZN(n3310) );
  AOI22_X1 U4099 ( .A1(n4390), .A2(n4196), .B1(n3621), .B2(n3308), .ZN(n3309)
         );
  OAI211_X1 U4100 ( .C1(n4401), .C2(n3311), .A(n3310), .B(n3309), .ZN(n3312)
         );
  AOI21_X1 U4101 ( .B1(n3313), .B2(n4396), .A(n3312), .ZN(n3314) );
  INV_X1 U4102 ( .A(n3314), .ZN(U3231) );
  OAI22_X1 U4103 ( .A1(n3316), .A2(n3448), .B1(n2352), .B2(n4068), .ZN(n3315)
         );
  XNOR2_X1 U4104 ( .A(n3315), .B(n3332), .ZN(n3410) );
  OAI22_X1 U4105 ( .A1(n3316), .A2(n3445), .B1(n3448), .B2(n4068), .ZN(n3409)
         );
  XNOR2_X1 U4106 ( .A(n3410), .B(n3409), .ZN(n3390) );
  NAND2_X1 U4107 ( .A1(n3319), .A2(n3318), .ZN(n3324) );
  NAND2_X1 U4108 ( .A1(n4196), .A2(n3381), .ZN(n3326) );
  NAND2_X1 U4109 ( .A1(n3488), .A2(n3438), .ZN(n3325) );
  NAND2_X1 U4110 ( .A1(n3326), .A2(n3325), .ZN(n3327) );
  XNOR2_X1 U4111 ( .A(n3327), .B(n3431), .ZN(n3330) );
  NOR2_X1 U4112 ( .A1(n4229), .A2(n3448), .ZN(n3328) );
  AOI21_X1 U4113 ( .B1(n4196), .B2(n3042), .A(n3328), .ZN(n3329) );
  NOR2_X1 U4114 ( .A1(n3330), .A2(n3329), .ZN(n3484) );
  NAND2_X1 U4115 ( .A1(n3330), .A2(n3329), .ZN(n3485) );
  OAI22_X1 U4116 ( .A1(n4385), .A2(n3448), .B1(n2352), .B2(n4202), .ZN(n3331)
         );
  NAND2_X1 U4117 ( .A1(n4171), .A2(n3042), .ZN(n3334) );
  NAND2_X1 U4118 ( .A1(n3620), .A2(n3381), .ZN(n3333) );
  NAND2_X1 U4119 ( .A1(n3334), .A2(n3333), .ZN(n4392) );
  NAND2_X1 U4120 ( .A1(n4195), .A2(n3381), .ZN(n3336) );
  NAND2_X1 U4121 ( .A1(n4176), .A2(n3438), .ZN(n3335) );
  NAND2_X1 U4122 ( .A1(n3336), .A2(n3335), .ZN(n3337) );
  XNOR2_X1 U4123 ( .A(n3337), .B(n3332), .ZN(n3341) );
  NAND2_X1 U4124 ( .A1(n4195), .A2(n3282), .ZN(n3339) );
  NAND2_X1 U4125 ( .A1(n4176), .A2(n3381), .ZN(n3338) );
  NAND2_X1 U4126 ( .A1(n3339), .A2(n3338), .ZN(n3340) );
  NOR2_X1 U4127 ( .A1(n3341), .A2(n3340), .ZN(n3343) );
  AND2_X1 U4128 ( .A1(n2247), .A2(n3485), .ZN(n3342) );
  INV_X1 U4129 ( .A(n3343), .ZN(n3344) );
  NAND2_X1 U4130 ( .A1(n3345), .A2(n3344), .ZN(n3556) );
  NAND2_X1 U4131 ( .A1(n4389), .A2(n3381), .ZN(n3347) );
  NAND2_X1 U4132 ( .A1(n3558), .A2(n3438), .ZN(n3346) );
  NAND2_X1 U4133 ( .A1(n3347), .A2(n3346), .ZN(n3348) );
  XNOR2_X1 U4134 ( .A(n3348), .B(n3332), .ZN(n3351) );
  NAND2_X1 U4135 ( .A1(n4389), .A2(n3042), .ZN(n3350) );
  NAND2_X1 U4136 ( .A1(n3558), .A2(n3381), .ZN(n3349) );
  NAND2_X1 U4137 ( .A1(n3350), .A2(n3349), .ZN(n3352) );
  NAND2_X1 U4138 ( .A1(n3351), .A2(n3352), .ZN(n3555) );
  NAND2_X1 U4139 ( .A1(n3556), .A2(n3555), .ZN(n3355) );
  INV_X1 U4140 ( .A(n3351), .ZN(n3354) );
  INV_X1 U4141 ( .A(n3352), .ZN(n3353) );
  NAND2_X1 U4142 ( .A1(n3354), .A2(n3353), .ZN(n3554) );
  NAND2_X1 U4143 ( .A1(n3355), .A2(n3554), .ZN(n3595) );
  NAND2_X1 U4144 ( .A1(n4155), .A2(n3381), .ZN(n3357) );
  NAND2_X1 U4145 ( .A1(n4135), .A2(n3438), .ZN(n3356) );
  NAND2_X1 U4146 ( .A1(n3357), .A2(n3356), .ZN(n3358) );
  XNOR2_X1 U4147 ( .A(n3358), .B(n3332), .ZN(n3361) );
  NAND2_X1 U4148 ( .A1(n4155), .A2(n3282), .ZN(n3360) );
  NAND2_X1 U4149 ( .A1(n4135), .A2(n3381), .ZN(n3359) );
  NAND2_X1 U4150 ( .A1(n3360), .A2(n3359), .ZN(n3362) );
  NAND2_X1 U4151 ( .A1(n3361), .A2(n3362), .ZN(n3597) );
  INV_X1 U4152 ( .A(n3361), .ZN(n3364) );
  INV_X1 U4153 ( .A(n3362), .ZN(n3363) );
  NAND2_X1 U4154 ( .A1(n3364), .A2(n3363), .ZN(n3596) );
  OAI22_X1 U4155 ( .A1(n4103), .A2(n3445), .B1(n3448), .B2(n4126), .ZN(n3369)
         );
  NAND2_X1 U4156 ( .A1(n4136), .A2(n3381), .ZN(n3366) );
  NAND2_X1 U4157 ( .A1(n3506), .A2(n3438), .ZN(n3365) );
  NAND2_X1 U4158 ( .A1(n3366), .A2(n3365), .ZN(n3367) );
  XNOR2_X1 U4159 ( .A(n3367), .B(n3332), .ZN(n3368) );
  XOR2_X1 U4160 ( .A(n3369), .B(n3368), .Z(n3503) );
  INV_X1 U4161 ( .A(n3368), .ZN(n3371) );
  INV_X1 U4162 ( .A(n3369), .ZN(n3370) );
  NAND2_X1 U4163 ( .A1(n4122), .A2(n3381), .ZN(n3373) );
  NAND2_X1 U4164 ( .A1(n4107), .A2(n3438), .ZN(n3372) );
  NAND2_X1 U4165 ( .A1(n3373), .A2(n3372), .ZN(n3374) );
  XNOR2_X1 U4166 ( .A(n3374), .B(n3332), .ZN(n3377) );
  NAND2_X1 U4167 ( .A1(n4122), .A2(n3042), .ZN(n3376) );
  NAND2_X1 U4168 ( .A1(n4107), .A2(n3381), .ZN(n3375) );
  NAND2_X1 U4169 ( .A1(n3376), .A2(n3375), .ZN(n3378) );
  NAND2_X1 U4170 ( .A1(n3377), .A2(n3378), .ZN(n3585) );
  NAND2_X1 U4171 ( .A1(n3584), .A2(n3585), .ZN(n3583) );
  INV_X1 U4172 ( .A(n3377), .ZN(n3380) );
  INV_X1 U4173 ( .A(n3378), .ZN(n3379) );
  NAND2_X1 U4174 ( .A1(n3380), .A2(n3379), .ZN(n3587) );
  NAND2_X1 U4175 ( .A1(n4101), .A2(n3381), .ZN(n3383) );
  NAND2_X1 U4176 ( .A1(n3518), .A2(n3438), .ZN(n3382) );
  NAND2_X1 U4177 ( .A1(n3383), .A2(n3382), .ZN(n3384) );
  XNOR2_X1 U4178 ( .A(n3384), .B(n3332), .ZN(n3512) );
  NAND2_X1 U4179 ( .A1(n4101), .A2(n3282), .ZN(n3386) );
  NAND2_X1 U4180 ( .A1(n3518), .A2(n3381), .ZN(n3385) );
  NAND2_X1 U4181 ( .A1(n3386), .A2(n3385), .ZN(n3513) );
  NOR2_X1 U4182 ( .A1(n3512), .A2(n3513), .ZN(n3388) );
  NAND2_X1 U4183 ( .A1(n3512), .A2(n3513), .ZN(n3387) );
  AOI21_X1 U4184 ( .B1(n3390), .B2(n3389), .A(n2233), .ZN(n3396) );
  INV_X1 U4185 ( .A(n4069), .ZN(n3394) );
  INV_X1 U4186 ( .A(REG3_REG_22__SCAN_IN), .ZN(n3391) );
  OAI22_X1 U4187 ( .A1(n4384), .A2(n4065), .B1(STATE_REG_SCAN_IN), .B2(n3391), 
        .ZN(n3393) );
  OAI22_X1 U4188 ( .A1(n4387), .A2(n4068), .B1(n4022), .B2(n3610), .ZN(n3392)
         );
  AOI211_X1 U4189 ( .C1(n3614), .C2(n3394), .A(n3393), .B(n3392), .ZN(n3395)
         );
  OAI21_X1 U4190 ( .B1(n3396), .B2(n3616), .A(n3395), .ZN(U3232) );
  INV_X1 U4191 ( .A(n3397), .ZN(n3399) );
  NOR3_X1 U4192 ( .A1(n3401), .A2(n3400), .A3(n2795), .ZN(n3402) );
  AOI21_X1 U4193 ( .B1(n4575), .B2(n3403), .A(n3402), .ZN(U3459) );
  INV_X1 U4194 ( .A(n4374), .ZN(n3404) );
  AND2_X1 U4195 ( .A1(n3404), .A2(n4588), .ZN(n3406) );
  AOI22_X1 U4196 ( .A1(n4575), .A2(n4791), .B1(n3406), .B2(n3405), .ZN(U3458)
         );
  NOR2_X1 U4197 ( .A1(n4048), .A2(n3448), .ZN(n3407) );
  AOI21_X1 U4198 ( .B1(n4062), .B2(n3042), .A(n3407), .ZN(n3414) );
  OAI22_X1 U4199 ( .A1(n4022), .A2(n3448), .B1(n2352), .B2(n4048), .ZN(n3408)
         );
  XNOR2_X1 U4200 ( .A(n3408), .B(n3332), .ZN(n3413) );
  XOR2_X1 U4201 ( .A(n3414), .B(n3413), .Z(n3494) );
  NOR2_X1 U4202 ( .A1(n3410), .A2(n3409), .ZN(n3495) );
  NOR2_X1 U4203 ( .A1(n3494), .A2(n3495), .ZN(n3411) );
  NOR2_X1 U4204 ( .A1(n4027), .A2(n3448), .ZN(n3412) );
  AOI21_X1 U4205 ( .B1(n4004), .B2(n3042), .A(n3412), .ZN(n3418) );
  INV_X1 U4206 ( .A(n3413), .ZN(n3415) );
  OR2_X1 U4207 ( .A1(n3415), .A2(n3414), .ZN(n3417) );
  NAND3_X1 U4208 ( .A1(n3496), .A2(n3418), .A3(n3417), .ZN(n3564) );
  OAI22_X1 U4209 ( .A1(n4044), .A2(n3448), .B1(n2352), .B2(n4027), .ZN(n3416)
         );
  XNOR2_X1 U4210 ( .A(n3416), .B(n3332), .ZN(n3566) );
  NAND2_X1 U4211 ( .A1(n3564), .A2(n3566), .ZN(n3421) );
  NAND2_X1 U4212 ( .A1(n3496), .A2(n3417), .ZN(n3420) );
  INV_X1 U4213 ( .A(n3418), .ZN(n3419) );
  NAND2_X1 U4214 ( .A1(n3420), .A2(n3419), .ZN(n3565) );
  NAND2_X1 U4215 ( .A1(n3421), .A2(n3565), .ZN(n3545) );
  NAND2_X1 U4216 ( .A1(n4024), .A2(n3381), .ZN(n3423) );
  NAND2_X1 U4217 ( .A1(n4003), .A2(n3438), .ZN(n3422) );
  NAND2_X1 U4218 ( .A1(n3423), .A2(n3422), .ZN(n3424) );
  XNOR2_X1 U4219 ( .A(n3424), .B(n3431), .ZN(n3427) );
  NOR2_X1 U4220 ( .A1(n4010), .A2(n3448), .ZN(n3425) );
  AOI21_X1 U4221 ( .B1(n4024), .B2(n3282), .A(n3425), .ZN(n3426) );
  NAND2_X1 U4222 ( .A1(n3427), .A2(n3426), .ZN(n3542) );
  NOR2_X1 U4223 ( .A1(n3427), .A2(n3426), .ZN(n3541) );
  NAND2_X1 U4224 ( .A1(n4002), .A2(n3381), .ZN(n3430) );
  NAND2_X1 U4225 ( .A1(n3428), .A2(n3438), .ZN(n3429) );
  NAND2_X1 U4226 ( .A1(n3430), .A2(n3429), .ZN(n3432) );
  XNOR2_X1 U4227 ( .A(n3432), .B(n3431), .ZN(n3437) );
  INV_X1 U4228 ( .A(n3437), .ZN(n3435) );
  NOR2_X1 U4229 ( .A1(n3988), .A2(n3448), .ZN(n3433) );
  AOI21_X1 U4230 ( .B1(n4002), .B2(n3042), .A(n3433), .ZN(n3436) );
  INV_X1 U4231 ( .A(n3436), .ZN(n3434) );
  NAND2_X1 U4232 ( .A1(n3435), .A2(n3434), .ZN(n3605) );
  NAND2_X1 U4233 ( .A1(n3983), .A2(n3381), .ZN(n3441) );
  NAND2_X1 U4234 ( .A1(n3439), .A2(n3438), .ZN(n3440) );
  NAND2_X1 U4235 ( .A1(n3441), .A2(n3440), .ZN(n3442) );
  XNOR2_X1 U4236 ( .A(n3442), .B(n3332), .ZN(n3451) );
  NOR2_X1 U4237 ( .A1(n3971), .A2(n3448), .ZN(n3443) );
  AOI21_X1 U4238 ( .B1(n3983), .B2(n3042), .A(n3443), .ZN(n3452) );
  XNOR2_X1 U4239 ( .A(n3451), .B(n3452), .ZN(n3476) );
  OAI22_X1 U4240 ( .A1(n3479), .A2(n3445), .B1(n3448), .B2(n3447), .ZN(n3446)
         );
  XNOR2_X1 U4241 ( .A(n3446), .B(n3332), .ZN(n3450) );
  OAI22_X1 U4242 ( .A1(n3479), .A2(n3448), .B1(n2352), .B2(n3447), .ZN(n3449)
         );
  XNOR2_X1 U4243 ( .A(n3450), .B(n3449), .ZN(n3455) );
  NAND2_X1 U4244 ( .A1(n3455), .A2(n4396), .ZN(n3466) );
  INV_X1 U4245 ( .A(n3451), .ZN(n3453) );
  NOR2_X1 U4246 ( .A1(n3453), .A2(n3452), .ZN(n3456) );
  NOR3_X1 U4247 ( .A1(n3455), .A2(n3456), .A3(n3616), .ZN(n3454) );
  INV_X1 U4248 ( .A(n3455), .ZN(n3458) );
  INV_X1 U4249 ( .A(n3456), .ZN(n3457) );
  NOR3_X1 U4250 ( .A1(n3458), .A2(n3616), .A3(n3457), .ZN(n3463) );
  AOI22_X1 U4251 ( .A1(n3983), .A2(n3622), .B1(REG3_REG_28__SCAN_IN), .B2(
        U3149), .ZN(n3461) );
  AOI22_X1 U4252 ( .A1(n3783), .A2(n4390), .B1(n3459), .B2(n3621), .ZN(n3460)
         );
  OAI211_X1 U4253 ( .C1(n4401), .C2(n3469), .A(n3461), .B(n3460), .ZN(n3462)
         );
  NOR2_X1 U4254 ( .A1(n3463), .A2(n3462), .ZN(n3464) );
  OAI211_X1 U4255 ( .C1(n3467), .C2(n3466), .A(n3465), .B(n3464), .ZN(U3217)
         );
  INV_X1 U4256 ( .A(n4251), .ZN(n3473) );
  INV_X1 U4257 ( .A(REG2_REG_28__SCAN_IN), .ZN(n3468) );
  OAI22_X1 U4258 ( .A1(n3469), .A2(n4231), .B1(n3468), .B2(n4207), .ZN(n3472)
         );
  NOR2_X1 U4259 ( .A1(n3470), .A2(n4564), .ZN(n3471) );
  AOI211_X1 U4260 ( .C1(n4569), .C2(n3473), .A(n3472), .B(n3471), .ZN(n3474)
         );
  OAI21_X1 U4261 ( .B1(n3475), .B2(n4211), .A(n3474), .ZN(U3262) );
  XNOR2_X1 U4262 ( .A(n3477), .B(n3476), .ZN(n3483) );
  INV_X1 U4263 ( .A(n3478), .ZN(n3972) );
  OAI22_X1 U4264 ( .A1(n3964), .A2(n4384), .B1(n4387), .B2(n3971), .ZN(n3481)
         );
  OAI22_X1 U4265 ( .A1(n3479), .A2(n3610), .B1(STATE_REG_SCAN_IN), .B2(n4957), 
        .ZN(n3480) );
  AOI211_X1 U4266 ( .C1(n3972), .C2(n3614), .A(n3481), .B(n3480), .ZN(n3482)
         );
  OAI21_X1 U4267 ( .B1(n3483), .B2(n3616), .A(n3482), .ZN(U3211) );
  NAND2_X1 U4268 ( .A1(n2348), .A2(n3485), .ZN(n3486) );
  XNOR2_X1 U4269 ( .A(n3487), .B(n3486), .ZN(n3492) );
  AND2_X1 U4270 ( .A1(REG3_REG_14__SCAN_IN), .A2(U3149), .ZN(n4511) );
  AOI21_X1 U4271 ( .B1(n4390), .B2(n4171), .A(n4511), .ZN(n3490) );
  AOI22_X1 U4272 ( .A1(n3622), .A2(n4218), .B1(n3621), .B2(n3488), .ZN(n3489)
         );
  OAI211_X1 U4273 ( .C1(n4401), .C2(n4232), .A(n3490), .B(n3489), .ZN(n3491)
         );
  AOI21_X1 U4274 ( .B1(n3492), .B2(n4396), .A(n3491), .ZN(n3493) );
  INV_X1 U4275 ( .A(n3493), .ZN(U3212) );
  OAI21_X1 U4276 ( .B1(n2233), .B2(n3495), .A(n3494), .ZN(n3497) );
  NAND3_X1 U4277 ( .A1(n3497), .A2(n4396), .A3(n3496), .ZN(n3502) );
  AOI22_X1 U4278 ( .A1(n4390), .A2(n4004), .B1(REG3_REG_23__SCAN_IN), .B2(
        U3149), .ZN(n3501) );
  AOI22_X1 U4279 ( .A1(n3622), .A2(n4081), .B1(n3621), .B2(n3498), .ZN(n3500)
         );
  OR2_X1 U4280 ( .A1(n4401), .A2(n4051), .ZN(n3499) );
  NAND4_X1 U4281 ( .A1(n3502), .A2(n3501), .A3(n3500), .A4(n3499), .ZN(U3213)
         );
  XNOR2_X1 U4282 ( .A(n3504), .B(n3503), .ZN(n3510) );
  NAND2_X1 U4283 ( .A1(U3149), .A2(REG3_REG_19__SCAN_IN), .ZN(n3940) );
  INV_X1 U4284 ( .A(n3940), .ZN(n3505) );
  AOI21_X1 U4285 ( .B1(n3622), .B2(n4155), .A(n3505), .ZN(n3508) );
  AOI22_X1 U4286 ( .A1(n4390), .A2(n4122), .B1(n3621), .B2(n3506), .ZN(n3507)
         );
  OAI211_X1 U4287 ( .C1(n4401), .C2(n4127), .A(n3508), .B(n3507), .ZN(n3509)
         );
  AOI21_X1 U4288 ( .B1(n3510), .B2(n4396), .A(n3509), .ZN(n3511) );
  INV_X1 U4289 ( .A(n3511), .ZN(U3216) );
  XOR2_X1 U4290 ( .A(n3513), .B(n3512), .Z(n3514) );
  XNOR2_X1 U4291 ( .A(n3515), .B(n3514), .ZN(n3522) );
  NOR2_X1 U4292 ( .A1(n3516), .A2(STATE_REG_SCAN_IN), .ZN(n3517) );
  AOI21_X1 U4293 ( .B1(n4390), .B2(n4081), .A(n3517), .ZN(n3520) );
  AOI22_X1 U4294 ( .A1(n3622), .A2(n4122), .B1(n3621), .B2(n3518), .ZN(n3519)
         );
  OAI211_X1 U4295 ( .C1(n4401), .C2(n4088), .A(n3520), .B(n3519), .ZN(n3521)
         );
  AOI21_X1 U4296 ( .B1(n3522), .B2(n4396), .A(n3521), .ZN(n3523) );
  INV_X1 U4297 ( .A(n3523), .ZN(U3220) );
  INV_X1 U4298 ( .A(n3299), .ZN(n3528) );
  NAND2_X1 U4299 ( .A1(n3299), .A2(n3524), .ZN(n3526) );
  AOI22_X1 U4300 ( .A1(n3528), .A2(n3527), .B1(n3526), .B2(n3525), .ZN(n3532)
         );
  NOR2_X1 U4301 ( .A1(n3530), .A2(n3529), .ZN(n3531) );
  XNOR2_X1 U4302 ( .A(n3532), .B(n3531), .ZN(n3539) );
  NAND2_X1 U4303 ( .A1(REG3_REG_12__SCAN_IN), .A2(U3149), .ZN(n4488) );
  INV_X1 U4304 ( .A(n4488), .ZN(n3533) );
  AOI21_X1 U4305 ( .B1(n3622), .B2(n3785), .A(n3533), .ZN(n3536) );
  AOI22_X1 U4306 ( .A1(n4390), .A2(n4218), .B1(n3621), .B2(n3534), .ZN(n3535)
         );
  OAI211_X1 U4307 ( .C1(n4401), .C2(n3537), .A(n3536), .B(n3535), .ZN(n3538)
         );
  AOI21_X1 U4308 ( .B1(n3539), .B2(n4396), .A(n3538), .ZN(n3540) );
  INV_X1 U4309 ( .A(n3540), .ZN(U3221) );
  INV_X1 U4310 ( .A(n3541), .ZN(n3543) );
  NAND2_X1 U4311 ( .A1(n3543), .A2(n3542), .ZN(n3544) );
  XNOR2_X1 U4312 ( .A(n3545), .B(n3544), .ZN(n3552) );
  INV_X1 U4313 ( .A(n4012), .ZN(n3550) );
  NOR2_X1 U4314 ( .A1(n3546), .A2(STATE_REG_SCAN_IN), .ZN(n3547) );
  AOI21_X1 U4315 ( .B1(n3622), .B2(n4004), .A(n3547), .ZN(n3549) );
  AOI22_X1 U4316 ( .A1(n4002), .A2(n4390), .B1(n4003), .B2(n3621), .ZN(n3548)
         );
  OAI211_X1 U4317 ( .C1(n4401), .C2(n3550), .A(n3549), .B(n3548), .ZN(n3551)
         );
  AOI21_X1 U4318 ( .B1(n3552), .B2(n4396), .A(n3551), .ZN(n3553) );
  INV_X1 U4319 ( .A(n3553), .ZN(U3222) );
  NAND2_X1 U4320 ( .A1(n3555), .A2(n3554), .ZN(n3557) );
  XOR2_X1 U4321 ( .A(n3557), .B(n3556), .Z(n3562) );
  INV_X1 U4322 ( .A(REG3_REG_17__SCAN_IN), .ZN(n4954) );
  NOR2_X1 U4323 ( .A1(STATE_REG_SCAN_IN), .A2(n4954), .ZN(n4540) );
  AOI21_X1 U4324 ( .B1(n3622), .B2(n4195), .A(n4540), .ZN(n3560) );
  AOI22_X1 U4325 ( .A1(n4390), .A2(n4155), .B1(n3621), .B2(n3558), .ZN(n3559)
         );
  OAI211_X1 U4326 ( .C1(n4401), .C2(n4163), .A(n3560), .B(n3559), .ZN(n3561)
         );
  AOI21_X1 U4327 ( .B1(n3562), .B2(n4396), .A(n3561), .ZN(n3563) );
  INV_X1 U4328 ( .A(n3563), .ZN(U3225) );
  NAND2_X1 U4329 ( .A1(n3565), .A2(n3564), .ZN(n3567) );
  XNOR2_X1 U4330 ( .A(n3567), .B(n3566), .ZN(n3572) );
  AOI22_X1 U4331 ( .A1(n3622), .A2(n4062), .B1(REG3_REG_24__SCAN_IN), .B2(
        U3149), .ZN(n3570) );
  AOI22_X1 U4332 ( .A1(n4390), .A2(n4024), .B1(n3621), .B2(n3568), .ZN(n3569)
         );
  OAI211_X1 U4333 ( .C1(n4401), .C2(n4030), .A(n3570), .B(n3569), .ZN(n3571)
         );
  AOI21_X1 U4334 ( .B1(n3572), .B2(n4396), .A(n3571), .ZN(n3573) );
  INV_X1 U4335 ( .A(n3573), .ZN(U3226) );
  OAI211_X1 U4336 ( .C1(n3576), .C2(n3575), .A(n3574), .B(n4396), .ZN(n3582)
         );
  AND2_X1 U4337 ( .A1(U3149), .A2(REG3_REG_4__SCAN_IN), .ZN(n3849) );
  AOI21_X1 U4338 ( .B1(n4390), .B2(n3791), .A(n3849), .ZN(n3581) );
  AOI22_X1 U4339 ( .A1(n3622), .A2(n3793), .B1(n3621), .B2(n3577), .ZN(n3580)
         );
  OR2_X1 U4340 ( .A1(n4401), .A2(n3578), .ZN(n3579) );
  NAND4_X1 U4341 ( .A1(n3582), .A2(n3581), .A3(n3580), .A4(n3579), .ZN(U3227)
         );
  INV_X1 U4342 ( .A(n3583), .ZN(n3588) );
  AOI21_X1 U4343 ( .B1(n3587), .B2(n3585), .A(n3584), .ZN(n3586) );
  AOI21_X1 U4344 ( .B1(n3588), .B2(n3587), .A(n3586), .ZN(n3593) );
  AOI22_X1 U4345 ( .A1(n4390), .A2(n4101), .B1(REG3_REG_20__SCAN_IN), .B2(
        U3149), .ZN(n3590) );
  AOI22_X1 U4346 ( .A1(n3622), .A2(n4136), .B1(n3621), .B2(n4107), .ZN(n3589)
         );
  OAI211_X1 U4347 ( .C1(n4401), .C2(n4110), .A(n3590), .B(n3589), .ZN(n3591)
         );
  INV_X1 U4348 ( .A(n3591), .ZN(n3592) );
  OAI21_X1 U4349 ( .B1(n3593), .B2(n3616), .A(n3592), .ZN(U3230) );
  NOR2_X1 U4350 ( .A1(n3594), .A2(n2360), .ZN(n3599) );
  AOI21_X1 U4351 ( .B1(n3597), .B2(n3596), .A(n3595), .ZN(n3598) );
  OAI21_X1 U4352 ( .B1(n3599), .B2(n3598), .A(n4396), .ZN(n3604) );
  NAND2_X1 U4353 ( .A1(n3621), .A2(n4135), .ZN(n3600) );
  OAI21_X1 U4354 ( .B1(n4103), .B2(n3610), .A(n3600), .ZN(n3602) );
  INV_X1 U4355 ( .A(REG3_REG_18__SCAN_IN), .ZN(n3924) );
  OAI22_X1 U4356 ( .A1(n4138), .A2(n4384), .B1(STATE_REG_SCAN_IN), .B2(n3924), 
        .ZN(n3601) );
  NOR2_X1 U4357 ( .A1(n3602), .A2(n3601), .ZN(n3603) );
  OAI211_X1 U4358 ( .C1(n4401), .C2(n4141), .A(n3604), .B(n3603), .ZN(U3235)
         );
  NAND2_X1 U4359 ( .A1(n2249), .A2(n3605), .ZN(n3606) );
  XNOR2_X1 U4360 ( .A(n3607), .B(n3606), .ZN(n3617) );
  OAI22_X1 U4361 ( .A1(n3609), .A2(n4384), .B1(STATE_REG_SCAN_IN), .B2(n3608), 
        .ZN(n3613) );
  OAI22_X1 U4362 ( .A1(n3611), .A2(n3610), .B1(n4387), .B2(n3988), .ZN(n3612)
         );
  AOI211_X1 U4363 ( .C1(n3990), .C2(n3614), .A(n3613), .B(n3612), .ZN(n3615)
         );
  OAI21_X1 U4364 ( .B1(n3617), .B2(n3616), .A(n3615), .ZN(U3237) );
  NAND2_X1 U4365 ( .A1(n3618), .A2(n4391), .ZN(n3619) );
  XNOR2_X1 U4366 ( .A(n3619), .B(n4392), .ZN(n3626) );
  AND2_X1 U4367 ( .A1(U3149), .A2(REG3_REG_15__SCAN_IN), .ZN(n4520) );
  AOI21_X1 U4368 ( .B1(n4390), .B2(n4195), .A(n4520), .ZN(n3624) );
  AOI22_X1 U4369 ( .A1(n3622), .A2(n4196), .B1(n3621), .B2(n3620), .ZN(n3623)
         );
  OAI211_X1 U4370 ( .C1(n4401), .C2(n4205), .A(n3624), .B(n3623), .ZN(n3625)
         );
  AOI21_X1 U4371 ( .B1(n3626), .B2(n4396), .A(n3625), .ZN(n3627) );
  INV_X1 U4372 ( .A(n3627), .ZN(U3238) );
  INV_X1 U4373 ( .A(n3766), .ZN(n3629) );
  NOR2_X1 U4374 ( .A1(n3629), .A2(n3628), .ZN(n3980) );
  INV_X1 U4375 ( .A(n3980), .ZN(n3635) );
  INV_X1 U4376 ( .A(REG0_REG_31__SCAN_IN), .ZN(n4310) );
  NAND2_X1 U4377 ( .A1(n2219), .A2(REG2_REG_31__SCAN_IN), .ZN(n3631) );
  NAND2_X1 U4378 ( .A1(n2502), .A2(REG1_REG_31__SCAN_IN), .ZN(n3630) );
  OAI211_X1 U4379 ( .C1(n3632), .C2(n4310), .A(n3631), .B(n3630), .ZN(n3947)
         );
  NAND2_X1 U4380 ( .A1(n2659), .A2(DATAI_31_), .ZN(n3948) );
  NAND2_X1 U4381 ( .A1(n2659), .A2(DATAI_30_), .ZN(n3689) );
  NAND2_X1 U4382 ( .A1(n3782), .A2(n3689), .ZN(n3693) );
  OAI21_X1 U4383 ( .B1(n3947), .B2(n3948), .A(n3693), .ZN(n3771) );
  NAND2_X1 U4384 ( .A1(n3947), .A2(n3948), .ZN(n3770) );
  OR2_X1 U4385 ( .A1(n3782), .A2(n3689), .ZN(n3633) );
  AND2_X1 U4386 ( .A1(n3770), .A2(n3633), .ZN(n3690) );
  INV_X1 U4387 ( .A(n3690), .ZN(n3634) );
  NOR4_X1 U4388 ( .A1(n3636), .A2(n3635), .A3(n3771), .A4(n3634), .ZN(n3648)
         );
  INV_X1 U4389 ( .A(n3637), .ZN(n3639) );
  NAND2_X1 U4390 ( .A1(n3639), .A2(n3638), .ZN(n4036) );
  INV_X1 U4391 ( .A(n4036), .ZN(n4042) );
  NAND2_X1 U4392 ( .A1(n3641), .A2(n3640), .ZN(n4120) );
  NOR3_X1 U4393 ( .A1(n3962), .A2(n4042), .A3(n4120), .ZN(n3647) );
  NAND2_X1 U4394 ( .A1(n3642), .A2(n3996), .ZN(n4020) );
  NOR4_X1 U4395 ( .A1(n4020), .A2(n3645), .A3(n3644), .A4(n3643), .ZN(n3646)
         );
  NAND3_X1 U4396 ( .A1(n3648), .A2(n3647), .A3(n3646), .ZN(n3670) );
  INV_X1 U4397 ( .A(n3649), .ZN(n3650) );
  XNOR2_X1 U4398 ( .A(n4122), .B(n3651), .ZN(n4099) );
  OR4_X1 U4399 ( .A1(n3999), .A2(n3652), .A3(n4191), .A4(n4099), .ZN(n3668) );
  INV_X1 U4400 ( .A(n3756), .ZN(n3653) );
  INV_X1 U4401 ( .A(n4075), .ZN(n4077) );
  NAND2_X1 U4402 ( .A1(n2293), .A2(n4095), .ZN(n4151) );
  NOR4_X1 U4403 ( .A1(n4077), .A2(n4151), .A3(n3655), .A4(n3654), .ZN(n3666)
         );
  NOR4_X1 U4404 ( .A1(n3658), .A2(n3657), .A3(n4143), .A4(n3656), .ZN(n3665)
         );
  NOR4_X1 U4405 ( .A1(n3661), .A2(n3660), .A3(n3659), .A4(n2743), .ZN(n3664)
         );
  INV_X1 U4406 ( .A(n4180), .ZN(n4169) );
  NOR4_X1 U4407 ( .A1(n4169), .A2(n4058), .A3(n3716), .A4(n3662), .ZN(n3663)
         );
  NAND4_X1 U4408 ( .A1(n3666), .A2(n3665), .A3(n3664), .A4(n3663), .ZN(n3667)
         );
  NOR4_X1 U4409 ( .A1(n3670), .A2(n3669), .A3(n3668), .A4(n3667), .ZN(n3699)
         );
  NAND2_X1 U4410 ( .A1(n4190), .A2(n3673), .ZN(n3740) );
  NAND2_X1 U4411 ( .A1(n3672), .A2(n3671), .ZN(n3731) );
  NAND2_X1 U4412 ( .A1(n3731), .A2(n3673), .ZN(n3739) );
  OAI21_X1 U4413 ( .B1(n4221), .B2(n3740), .A(n3739), .ZN(n3675) );
  NAND3_X1 U4414 ( .A1(n4098), .A2(n3747), .A3(n2293), .ZN(n3674) );
  AOI21_X1 U4415 ( .B1(n3675), .B2(n3745), .A(n3674), .ZN(n3677) );
  INV_X1 U4416 ( .A(n3676), .ZN(n3753) );
  OAI21_X1 U4417 ( .B1(n3677), .B2(n3753), .A(n3754), .ZN(n3678) );
  NAND2_X1 U4418 ( .A1(n3678), .A2(n3755), .ZN(n3680) );
  INV_X1 U4419 ( .A(n3679), .ZN(n3758) );
  AOI21_X1 U4420 ( .B1(n3681), .B2(n3680), .A(n3758), .ZN(n3682) );
  OAI21_X1 U4421 ( .B1(n3682), .B2(n3762), .A(n3761), .ZN(n3684) );
  INV_X1 U4422 ( .A(n3962), .ZN(n3683) );
  AND3_X1 U4423 ( .A1(n3684), .A2(n3683), .A3(n3766), .ZN(n3688) );
  NAND2_X1 U4424 ( .A1(n3686), .A2(n3685), .ZN(n3768) );
  AOI21_X1 U4425 ( .B1(n3783), .B2(n3691), .A(n3687), .ZN(n3769) );
  OAI21_X1 U4426 ( .B1(n3688), .B2(n3768), .A(n3769), .ZN(n3697) );
  INV_X1 U4427 ( .A(n3947), .ZN(n3692) );
  OAI21_X1 U4428 ( .B1(n3783), .B2(n3691), .A(n3690), .ZN(n3767) );
  AOI21_X1 U4429 ( .B1(n4245), .B2(n3692), .A(n3767), .ZN(n3696) );
  INV_X1 U4430 ( .A(n3948), .ZN(n3695) );
  NAND2_X1 U4431 ( .A1(n3693), .A2(n3947), .ZN(n3694) );
  AOI22_X1 U4432 ( .A1(n3697), .A2(n3696), .B1(n3695), .B2(n3694), .ZN(n3698)
         );
  MUX2_X1 U4433 ( .A(n3699), .B(n3698), .S(n3703), .Z(n3776) );
  INV_X1 U4434 ( .A(n3700), .ZN(n3704) );
  OAI211_X1 U4435 ( .C1(n3704), .C2(n3703), .A(n3702), .B(n3701), .ZN(n3706)
         );
  NAND3_X1 U4436 ( .A1(n3706), .A2(n3705), .A3(n2744), .ZN(n3709) );
  NAND3_X1 U4437 ( .A1(n3709), .A2(n3708), .A3(n3707), .ZN(n3712) );
  NAND3_X1 U4438 ( .A1(n3712), .A2(n3711), .A3(n3710), .ZN(n3715) );
  NAND4_X1 U4439 ( .A1(n3715), .A2(n3714), .A3(n3713), .A4(n3725), .ZN(n3719)
         );
  INV_X1 U4440 ( .A(n3716), .ZN(n3718) );
  NAND3_X1 U4441 ( .A1(n3719), .A2(n3718), .A3(n3717), .ZN(n3720) );
  NAND3_X1 U4442 ( .A1(n3720), .A2(n3727), .A3(n3726), .ZN(n3723) );
  AND3_X1 U4443 ( .A1(n3723), .A2(n3722), .A3(n3721), .ZN(n3732) );
  INV_X1 U4444 ( .A(n3739), .ZN(n3730) );
  INV_X1 U4445 ( .A(n3724), .ZN(n3728) );
  NAND4_X1 U4446 ( .A1(n3728), .A2(n3727), .A3(n3726), .A4(n3725), .ZN(n3729)
         );
  OAI22_X1 U4447 ( .A1(n3732), .A2(n3731), .B1(n3730), .B2(n3729), .ZN(n3735)
         );
  AOI22_X1 U4448 ( .A1(n3735), .A2(n3734), .B1(n2295), .B2(n3739), .ZN(n3744)
         );
  NAND2_X1 U4449 ( .A1(n3737), .A2(n3736), .ZN(n3743) );
  INV_X1 U4450 ( .A(n3738), .ZN(n3741) );
  OAI21_X1 U4451 ( .B1(n3741), .B2(n3740), .A(n3739), .ZN(n3742) );
  OAI21_X1 U4452 ( .B1(n3744), .B2(n3743), .A(n3742), .ZN(n3748) );
  INV_X1 U4453 ( .A(n3745), .ZN(n3746) );
  AOI21_X1 U4454 ( .B1(n3748), .B2(n3747), .A(n3746), .ZN(n3751) );
  INV_X1 U4455 ( .A(n3754), .ZN(n3750) );
  NOR4_X1 U4456 ( .A1(n3751), .A2(n3750), .A3(n4096), .A4(n3749), .ZN(n3752)
         );
  AOI21_X1 U4457 ( .B1(n3754), .B2(n3753), .A(n3752), .ZN(n3757) );
  OAI21_X1 U4458 ( .B1(n3757), .B2(n3756), .A(n3755), .ZN(n3759) );
  AOI21_X1 U4459 ( .B1(n3760), .B2(n3759), .A(n3758), .ZN(n3763) );
  OAI21_X1 U4460 ( .B1(n3763), .B2(n3762), .A(n3761), .ZN(n3764) );
  NAND4_X1 U4461 ( .A1(n3769), .A2(n3766), .A3(n3765), .A4(n3764), .ZN(n3773)
         );
  AOI21_X1 U4462 ( .B1(n3769), .B2(n3768), .A(n3767), .ZN(n3772) );
  AOI22_X1 U4463 ( .A1(n3773), .A2(n3772), .B1(n3771), .B2(n3770), .ZN(n3775)
         );
  MUX2_X1 U4464 ( .A(n3776), .B(n3775), .S(n3774), .Z(n3777) );
  XNOR2_X1 U4465 ( .A(n3777), .B(n4377), .ZN(n3781) );
  INV_X1 U4466 ( .A(n4406), .ZN(n3809) );
  NOR2_X1 U4467 ( .A1(n4382), .A2(n3809), .ZN(n3811) );
  NAND2_X1 U4468 ( .A1(n3811), .A2(n2432), .ZN(n3778) );
  OAI211_X1 U4469 ( .C1(n4375), .C2(n3780), .A(n3778), .B(B_REG_SCAN_IN), .ZN(
        n3779) );
  OAI21_X1 U4470 ( .B1(n3781), .B2(n3780), .A(n3779), .ZN(U3239) );
  MUX2_X1 U4471 ( .A(DATAO_REG_31__SCAN_IN), .B(n3947), .S(U4043), .Z(U3581)
         );
  MUX2_X1 U4472 ( .A(DATAO_REG_30__SCAN_IN), .B(n3782), .S(U4043), .Z(U3580)
         );
  MUX2_X1 U4473 ( .A(n3783), .B(DATAO_REG_29__SCAN_IN), .S(n3795), .Z(U3579)
         );
  MUX2_X1 U4474 ( .A(n3966), .B(DATAO_REG_28__SCAN_IN), .S(n3795), .Z(U3578)
         );
  MUX2_X1 U4475 ( .A(n3983), .B(DATAO_REG_27__SCAN_IN), .S(n3795), .Z(U3577)
         );
  MUX2_X1 U4476 ( .A(n4002), .B(DATAO_REG_26__SCAN_IN), .S(n3795), .Z(U3576)
         );
  MUX2_X1 U4477 ( .A(n4024), .B(DATAO_REG_25__SCAN_IN), .S(n3795), .Z(U3575)
         );
  MUX2_X1 U4478 ( .A(n4004), .B(DATAO_REG_24__SCAN_IN), .S(n3795), .Z(U3574)
         );
  MUX2_X1 U4479 ( .A(n4062), .B(DATAO_REG_23__SCAN_IN), .S(n3795), .Z(U3573)
         );
  MUX2_X1 U4480 ( .A(n4081), .B(DATAO_REG_22__SCAN_IN), .S(n3795), .Z(U3572)
         );
  MUX2_X1 U4481 ( .A(n4101), .B(DATAO_REG_21__SCAN_IN), .S(n3795), .Z(U3571)
         );
  MUX2_X1 U4482 ( .A(n4122), .B(DATAO_REG_20__SCAN_IN), .S(n3795), .Z(U3570)
         );
  MUX2_X1 U4483 ( .A(n4136), .B(DATAO_REG_19__SCAN_IN), .S(n3795), .Z(U3569)
         );
  MUX2_X1 U4484 ( .A(n4155), .B(DATAO_REG_18__SCAN_IN), .S(n3795), .Z(U3568)
         );
  MUX2_X1 U4485 ( .A(n4389), .B(DATAO_REG_17__SCAN_IN), .S(n3795), .Z(U3567)
         );
  MUX2_X1 U4486 ( .A(n4195), .B(DATAO_REG_16__SCAN_IN), .S(n3795), .Z(U3566)
         );
  MUX2_X1 U4487 ( .A(n4171), .B(DATAO_REG_15__SCAN_IN), .S(n3795), .Z(U3565)
         );
  MUX2_X1 U4488 ( .A(n4196), .B(DATAO_REG_14__SCAN_IN), .S(n3795), .Z(U3564)
         );
  MUX2_X1 U4489 ( .A(n4218), .B(DATAO_REG_13__SCAN_IN), .S(n3795), .Z(U3563)
         );
  MUX2_X1 U4490 ( .A(n3784), .B(DATAO_REG_12__SCAN_IN), .S(n3795), .Z(U3562)
         );
  MUX2_X1 U4491 ( .A(n3785), .B(DATAO_REG_11__SCAN_IN), .S(n3795), .Z(U3561)
         );
  MUX2_X1 U4492 ( .A(n3786), .B(DATAO_REG_10__SCAN_IN), .S(n3795), .Z(U3560)
         );
  MUX2_X1 U4493 ( .A(n3787), .B(DATAO_REG_9__SCAN_IN), .S(n3795), .Z(U3559) );
  MUX2_X1 U4494 ( .A(n3788), .B(DATAO_REG_8__SCAN_IN), .S(n3795), .Z(U3558) );
  MUX2_X1 U4495 ( .A(n3789), .B(DATAO_REG_7__SCAN_IN), .S(n3795), .Z(U3557) );
  MUX2_X1 U4496 ( .A(n3790), .B(DATAO_REG_6__SCAN_IN), .S(n3795), .Z(U3556) );
  MUX2_X1 U4497 ( .A(n3791), .B(DATAO_REG_5__SCAN_IN), .S(n3795), .Z(U3555) );
  MUX2_X1 U4498 ( .A(n3792), .B(DATAO_REG_4__SCAN_IN), .S(n3795), .Z(U3554) );
  MUX2_X1 U4499 ( .A(n3793), .B(DATAO_REG_3__SCAN_IN), .S(n3795), .Z(U3553) );
  MUX2_X1 U4500 ( .A(n3794), .B(DATAO_REG_2__SCAN_IN), .S(n3795), .Z(U3552) );
  MUX2_X1 U4501 ( .A(n2887), .B(DATAO_REG_1__SCAN_IN), .S(n3795), .Z(U3551) );
  MUX2_X1 U4502 ( .A(n3796), .B(DATAO_REG_0__SCAN_IN), .S(n3795), .Z(U3550) );
  XNOR2_X1 U4503 ( .A(n3804), .B(REG1_REG_1__SCAN_IN), .ZN(n3801) );
  AND2_X1 U4504 ( .A1(IR_REG_0__SCAN_IN), .A2(REG1_REG_0__SCAN_IN), .ZN(n3800)
         );
  INV_X1 U4505 ( .A(n3797), .ZN(n3799) );
  NAND2_X1 U4506 ( .A1(n3801), .A2(n3800), .ZN(n3830) );
  OAI211_X1 U4507 ( .C1(n3801), .C2(n3800), .A(n4542), .B(n3830), .ZN(n3808)
         );
  AND2_X1 U4508 ( .A1(IR_REG_0__SCAN_IN), .A2(REG2_REG_0__SCAN_IN), .ZN(n3810)
         );
  INV_X1 U4509 ( .A(REG2_REG_1__SCAN_IN), .ZN(n3802) );
  MUX2_X1 U4510 ( .A(n3802), .B(REG2_REG_1__SCAN_IN), .S(n3804), .Z(n3803) );
  OAI211_X1 U4511 ( .C1(n3810), .C2(n3803), .A(n4496), .B(n3826), .ZN(n3807)
         );
  INV_X1 U4512 ( .A(n4548), .ZN(n3840) );
  NAND2_X1 U4513 ( .A1(n3840), .A2(n2482), .ZN(n3806) );
  AOI22_X1 U4514 ( .A1(n4541), .A2(ADDR_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(U3149), .ZN(n3805) );
  NAND4_X1 U4515 ( .A1(n3808), .A2(n3807), .A3(n3806), .A4(n3805), .ZN(U3241)
         );
  NAND2_X1 U4516 ( .A1(n3814), .A2(n3809), .ZN(n3817) );
  AOI21_X1 U4517 ( .B1(n3811), .B2(n3810), .A(n3795), .ZN(n3816) );
  INV_X1 U4518 ( .A(REG2_REG_0__SCAN_IN), .ZN(n3812) );
  NAND2_X1 U4519 ( .A1(n4406), .A2(n3812), .ZN(n3813) );
  NAND2_X1 U4520 ( .A1(n3814), .A2(n3813), .ZN(n4407) );
  NAND2_X1 U4521 ( .A1(n4407), .A2(n2395), .ZN(n3815) );
  OAI211_X1 U4522 ( .C1(n3818), .C2(n3817), .A(n3816), .B(n3815), .ZN(n3864)
         );
  AOI22_X1 U4523 ( .A1(n4541), .A2(ADDR_REG_2__SCAN_IN), .B1(
        REG3_REG_2__SCAN_IN), .B2(U3149), .ZN(n3819) );
  OAI21_X1 U4524 ( .B1(n4548), .B2(n3836), .A(n3819), .ZN(n3820) );
  INV_X1 U4525 ( .A(n3820), .ZN(n3835) );
  NAND2_X1 U4526 ( .A1(n2482), .A2(REG2_REG_1__SCAN_IN), .ZN(n3825) );
  NAND2_X1 U4527 ( .A1(n3826), .A2(n3825), .ZN(n3823) );
  INV_X1 U4528 ( .A(REG2_REG_2__SCAN_IN), .ZN(n3821) );
  MUX2_X1 U4529 ( .A(n3821), .B(REG2_REG_2__SCAN_IN), .S(n3836), .Z(n3822) );
  NAND2_X1 U4530 ( .A1(n3823), .A2(n3822), .ZN(n3842) );
  MUX2_X1 U4531 ( .A(REG2_REG_2__SCAN_IN), .B(n3821), .S(n3836), .Z(n3824) );
  NAND3_X1 U4532 ( .A1(n3826), .A2(n3825), .A3(n3824), .ZN(n3827) );
  NAND3_X1 U4533 ( .A1(n4496), .A2(n3842), .A3(n3827), .ZN(n3834) );
  INV_X1 U4534 ( .A(REG1_REG_2__SCAN_IN), .ZN(n3828) );
  MUX2_X1 U4535 ( .A(n3828), .B(REG1_REG_2__SCAN_IN), .S(n3836), .Z(n3832) );
  NAND2_X1 U4536 ( .A1(n2482), .A2(REG1_REG_1__SCAN_IN), .ZN(n3829) );
  NAND2_X1 U4537 ( .A1(n3830), .A2(n3829), .ZN(n3831) );
  NAND2_X1 U4538 ( .A1(n3831), .A2(n3832), .ZN(n3838) );
  OAI211_X1 U4539 ( .C1(n3832), .C2(n3831), .A(n4542), .B(n3838), .ZN(n3833)
         );
  NAND4_X1 U4540 ( .A1(n3864), .A2(n3835), .A3(n3834), .A4(n3833), .ZN(U3242)
         );
  INV_X1 U4541 ( .A(n3836), .ZN(n4381) );
  NAND2_X1 U4542 ( .A1(n4381), .A2(REG1_REG_2__SCAN_IN), .ZN(n3837) );
  NAND2_X1 U4543 ( .A1(n3838), .A2(n3837), .ZN(n3852) );
  INV_X1 U4544 ( .A(n4380), .ZN(n3843) );
  XNOR2_X1 U4545 ( .A(n3852), .B(n3843), .ZN(n3839) );
  NAND2_X1 U4546 ( .A1(n3839), .A2(REG1_REG_3__SCAN_IN), .ZN(n3854) );
  OAI211_X1 U4547 ( .C1(REG1_REG_3__SCAN_IN), .C2(n3839), .A(n4542), .B(n3854), 
        .ZN(n3848) );
  NAND2_X1 U4548 ( .A1(n3840), .A2(n4380), .ZN(n3847) );
  AOI22_X1 U4549 ( .A1(n4541), .A2(ADDR_REG_3__SCAN_IN), .B1(
        REG3_REG_3__SCAN_IN), .B2(U3149), .ZN(n3846) );
  NAND2_X1 U4550 ( .A1(n4381), .A2(REG2_REG_2__SCAN_IN), .ZN(n3841) );
  NAND2_X1 U4551 ( .A1(n3842), .A2(n3841), .ZN(n3857) );
  XOR2_X1 U4552 ( .A(REG2_REG_3__SCAN_IN), .B(n3856), .Z(n3844) );
  NAND2_X1 U4553 ( .A1(n4496), .A2(n3844), .ZN(n3845) );
  NAND4_X1 U4554 ( .A1(n3848), .A2(n3847), .A3(n3846), .A4(n3845), .ZN(U3243)
         );
  AOI21_X1 U4555 ( .B1(n4541), .B2(ADDR_REG_4__SCAN_IN), .A(n3849), .ZN(n3850)
         );
  OAI21_X1 U4556 ( .B1(n4548), .B2(n3898), .A(n3850), .ZN(n3851) );
  INV_X1 U4557 ( .A(n3851), .ZN(n3863) );
  NAND2_X1 U4558 ( .A1(n3852), .A2(n4380), .ZN(n3853) );
  NAND2_X1 U4559 ( .A1(n3854), .A2(n3853), .ZN(n3868) );
  XNOR2_X1 U4560 ( .A(n3868), .B(n3898), .ZN(n3855) );
  OAI211_X1 U4561 ( .C1(REG1_REG_4__SCAN_IN), .C2(n3855), .A(n4542), .B(n3867), 
        .ZN(n3862) );
  NAND2_X1 U4562 ( .A1(n3856), .A2(REG2_REG_3__SCAN_IN), .ZN(n3859) );
  NAND2_X1 U4563 ( .A1(n3857), .A2(n4380), .ZN(n3858) );
  NAND2_X1 U4564 ( .A1(n3859), .A2(n3858), .ZN(n3897) );
  INV_X1 U4565 ( .A(n3898), .ZN(n4379) );
  XNOR2_X1 U4566 ( .A(n3897), .B(n4379), .ZN(n3901) );
  XNOR2_X1 U4567 ( .A(n3901), .B(REG2_REG_4__SCAN_IN), .ZN(n3860) );
  NAND2_X1 U4568 ( .A1(n4496), .A2(n3860), .ZN(n3861) );
  NAND4_X1 U4569 ( .A1(n3864), .A2(n3863), .A3(n3862), .A4(n3861), .ZN(U3244)
         );
  XNOR2_X1 U4570 ( .A(n3927), .B(REG1_REG_18__SCAN_IN), .ZN(n3930) );
  NOR2_X1 U4571 ( .A1(n3922), .A2(REG1_REG_17__SCAN_IN), .ZN(n3887) );
  NAND2_X1 U4572 ( .A1(REG1_REG_15__SCAN_IN), .A2(n3919), .ZN(n3882) );
  INV_X1 U4573 ( .A(n3919), .ZN(n4591) );
  INV_X1 U4574 ( .A(REG1_REG_15__SCAN_IN), .ZN(n3865) );
  AOI22_X1 U4575 ( .A1(REG1_REG_15__SCAN_IN), .A2(n3919), .B1(n4591), .B2(
        n3865), .ZN(n4523) );
  NAND2_X1 U4576 ( .A1(n3915), .A2(REG1_REG_13__SCAN_IN), .ZN(n3878) );
  INV_X1 U4577 ( .A(REG1_REG_13__SCAN_IN), .ZN(n3866) );
  INV_X1 U4578 ( .A(n3915), .ZN(n4593) );
  AOI22_X1 U4579 ( .A1(n3915), .A2(REG1_REG_13__SCAN_IN), .B1(n3866), .B2(
        n4593), .ZN(n4504) );
  INV_X1 U4580 ( .A(REG1_REG_11__SCAN_IN), .ZN(n4644) );
  AOI22_X1 U4581 ( .A1(REG1_REG_11__SCAN_IN), .A2(n3891), .B1(n4595), .B2(
        n4644), .ZN(n4476) );
  NAND2_X1 U4582 ( .A1(n3893), .A2(REG1_REG_9__SCAN_IN), .ZN(n3873) );
  INV_X1 U4583 ( .A(n3893), .ZN(n4596) );
  AOI22_X1 U4584 ( .A1(n3893), .A2(REG1_REG_9__SCAN_IN), .B1(n3109), .B2(n4596), .ZN(n4455) );
  NAND2_X1 U4585 ( .A1(n3896), .A2(REG1_REG_5__SCAN_IN), .ZN(n3869) );
  OAI21_X1 U4586 ( .B1(n3896), .B2(REG1_REG_5__SCAN_IN), .A(n3869), .ZN(n4413)
         );
  AOI21_X1 U4587 ( .B1(REG1_REG_5__SCAN_IN), .B2(n3896), .A(n4412), .ZN(n3870)
         );
  INV_X1 U4588 ( .A(n3903), .ZN(n4598) );
  XNOR2_X1 U4589 ( .A(n3870), .B(n4598), .ZN(n4424) );
  INV_X1 U4590 ( .A(REG1_REG_7__SCAN_IN), .ZN(n4641) );
  NAND2_X1 U4591 ( .A1(n4443), .A2(n3871), .ZN(n3872) );
  NAND2_X1 U4592 ( .A1(REG1_REG_8__SCAN_IN), .A2(n4450), .ZN(n4449) );
  NAND2_X1 U4593 ( .A1(n4464), .A2(n3874), .ZN(n3875) );
  NAND2_X1 U4594 ( .A1(REG1_REG_10__SCAN_IN), .A2(n4471), .ZN(n4470) );
  NAND2_X1 U4595 ( .A1(n4485), .A2(n3876), .ZN(n3877) );
  NAND2_X1 U4596 ( .A1(REG1_REG_12__SCAN_IN), .A2(n4492), .ZN(n4491) );
  NAND2_X1 U4597 ( .A1(n3879), .A2(n3880), .ZN(n3881) );
  NAND2_X1 U4598 ( .A1(REG1_REG_14__SCAN_IN), .A2(n4513), .ZN(n4512) );
  NAND2_X1 U4599 ( .A1(n3881), .A2(n4512), .ZN(n4522) );
  NAND2_X1 U4600 ( .A1(n4523), .A2(n4522), .ZN(n4521) );
  NOR2_X1 U4601 ( .A1(n3883), .A2(n3884), .ZN(n3885) );
  INV_X1 U4602 ( .A(REG1_REG_17__SCAN_IN), .ZN(n3886) );
  AOI22_X1 U4603 ( .A1(n3922), .A2(n3886), .B1(REG1_REG_17__SCAN_IN), .B2(
        n4589), .ZN(n4543) );
  NOR2_X1 U4604 ( .A1(n4544), .A2(n4543), .ZN(n4545) );
  NOR2_X1 U4605 ( .A1(n3887), .A2(n4545), .ZN(n3931) );
  XOR2_X1 U4606 ( .A(n3930), .B(n3931), .Z(n3929) );
  INV_X1 U4607 ( .A(n3927), .ZN(n4378) );
  INV_X1 U4608 ( .A(REG2_REG_18__SCAN_IN), .ZN(n3889) );
  NOR2_X1 U4609 ( .A1(n4378), .A2(n3889), .ZN(n3888) );
  AOI21_X1 U4610 ( .B1(n4378), .B2(n3889), .A(n3888), .ZN(n3923) );
  NOR2_X1 U4611 ( .A1(n3922), .A2(REG2_REG_17__SCAN_IN), .ZN(n3890) );
  AOI21_X1 U4612 ( .B1(REG2_REG_17__SCAN_IN), .B2(n3922), .A(n3890), .ZN(n4538) );
  NOR2_X1 U4613 ( .A1(n4593), .A2(n3232), .ZN(n4495) );
  NAND2_X1 U4614 ( .A1(REG2_REG_11__SCAN_IN), .A2(n3891), .ZN(n3912) );
  AOI22_X1 U4615 ( .A1(REG2_REG_11__SCAN_IN), .A2(n3891), .B1(n4595), .B2(
        n3185), .ZN(n4479) );
  NAND2_X1 U4616 ( .A1(n3893), .A2(REG2_REG_9__SCAN_IN), .ZN(n3909) );
  AOI22_X1 U4617 ( .A1(n3893), .A2(REG2_REG_9__SCAN_IN), .B1(n3892), .B2(n4596), .ZN(n4458) );
  NAND2_X1 U4618 ( .A1(n4432), .A2(REG2_REG_7__SCAN_IN), .ZN(n3906) );
  AOI22_X1 U4619 ( .A1(n4432), .A2(REG2_REG_7__SCAN_IN), .B1(n3894), .B2(n4597), .ZN(n4440) );
  NAND2_X1 U4620 ( .A1(n3896), .A2(REG2_REG_5__SCAN_IN), .ZN(n3902) );
  INV_X1 U4621 ( .A(n3896), .ZN(n4600) );
  AOI22_X1 U4622 ( .A1(n3896), .A2(REG2_REG_5__SCAN_IN), .B1(n3895), .B2(n4600), .ZN(n4419) );
  INV_X1 U4623 ( .A(REG2_REG_4__SCAN_IN), .ZN(n3900) );
  INV_X1 U4624 ( .A(n3897), .ZN(n3899) );
  NAND2_X1 U4625 ( .A1(n3903), .A2(n3904), .ZN(n3905) );
  NAND2_X1 U4626 ( .A1(REG2_REG_6__SCAN_IN), .A2(n4429), .ZN(n4428) );
  NAND2_X1 U4627 ( .A1(n4443), .A2(n3907), .ZN(n3908) );
  NAND2_X1 U4628 ( .A1(REG2_REG_8__SCAN_IN), .A2(n4445), .ZN(n4444) );
  NAND2_X1 U4629 ( .A1(n4464), .A2(n3910), .ZN(n3911) );
  NAND2_X1 U4630 ( .A1(REG2_REG_10__SCAN_IN), .A2(n4466), .ZN(n4465) );
  NAND2_X1 U4631 ( .A1(n4485), .A2(n3913), .ZN(n3914) );
  NAND2_X1 U4632 ( .A1(REG2_REG_12__SCAN_IN), .A2(n4487), .ZN(n4486) );
  NOR2_X1 U4633 ( .A1(n4592), .A2(n3916), .ZN(n3917) );
  INV_X1 U4634 ( .A(REG2_REG_14__SCAN_IN), .ZN(n4509) );
  NAND2_X1 U4635 ( .A1(REG2_REG_15__SCAN_IN), .A2(n3919), .ZN(n3918) );
  OAI21_X1 U4636 ( .B1(REG2_REG_15__SCAN_IN), .B2(n3919), .A(n3918), .ZN(n4517) );
  NAND2_X1 U4637 ( .A1(n3920), .A2(n4590), .ZN(n3921) );
  INV_X1 U4638 ( .A(REG2_REG_16__SCAN_IN), .ZN(n4526) );
  NAND2_X1 U4639 ( .A1(n3921), .A2(n4527), .ZN(n4536) );
  NAND2_X1 U4640 ( .A1(n4538), .A2(n4536), .ZN(n4537) );
  INV_X1 U4641 ( .A(n4496), .ZN(n4535) );
  NOR2_X1 U4642 ( .A1(STATE_REG_SCAN_IN), .A2(n3924), .ZN(n3925) );
  AOI21_X1 U4643 ( .B1(n4541), .B2(ADDR_REG_18__SCAN_IN), .A(n3925), .ZN(n3926) );
  OAI21_X1 U4644 ( .B1(n4548), .B2(n3927), .A(n3926), .ZN(n3928) );
  AOI22_X1 U4645 ( .A1(n3931), .A2(n3930), .B1(n4378), .B2(
        REG1_REG_18__SCAN_IN), .ZN(n3934) );
  INV_X1 U4646 ( .A(REG1_REG_19__SCAN_IN), .ZN(n3932) );
  MUX2_X1 U4647 ( .A(n3932), .B(REG1_REG_19__SCAN_IN), .S(n4377), .Z(n3933) );
  XNOR2_X1 U4648 ( .A(n3934), .B(n3933), .ZN(n3945) );
  INV_X1 U4649 ( .A(n4542), .ZN(n4422) );
  INV_X1 U4650 ( .A(REG2_REG_19__SCAN_IN), .ZN(n3936) );
  MUX2_X1 U4651 ( .A(REG2_REG_19__SCAN_IN), .B(n3936), .S(n4377), .Z(n3937) );
  XNOR2_X1 U4652 ( .A(n3938), .B(n3937), .ZN(n3943) );
  NAND2_X1 U4653 ( .A1(n4541), .A2(ADDR_REG_19__SCAN_IN), .ZN(n3939) );
  OAI211_X1 U4654 ( .C1(n4548), .C2(n3941), .A(n3940), .B(n3939), .ZN(n3942)
         );
  AOI21_X1 U4655 ( .B1(n3943), .B2(n4496), .A(n3942), .ZN(n3944) );
  OAI21_X1 U4656 ( .B1(n3945), .B2(n4422), .A(n3944), .ZN(U3259) );
  XNOR2_X1 U4657 ( .A(n4240), .B(n3948), .ZN(n4314) );
  NAND2_X1 U4658 ( .A1(n3947), .A2(n3946), .ZN(n4242) );
  OAI21_X1 U4659 ( .B1(n3948), .B2(n4215), .A(n4242), .ZN(n4312) );
  NAND2_X1 U4660 ( .A1(n4312), .A2(n4207), .ZN(n3950) );
  NAND2_X1 U4661 ( .A1(n4564), .A2(REG2_REG_31__SCAN_IN), .ZN(n3949) );
  OAI211_X1 U4662 ( .C1(n4314), .C2(n4204), .A(n3950), .B(n3949), .ZN(U3260)
         );
  NAND2_X1 U4663 ( .A1(n3952), .A2(n3951), .ZN(n3958) );
  OAI22_X1 U4664 ( .A1(n3954), .A2(n4204), .B1(n3953), .B2(n4231), .ZN(n3955)
         );
  OAI21_X1 U4665 ( .B1(n3956), .B2(n3955), .A(n4207), .ZN(n3957) );
  OAI211_X1 U4666 ( .C1(n4207), .C2(n3959), .A(n3958), .B(n3957), .ZN(U3354)
         );
  XNOR2_X1 U4667 ( .A(n3960), .B(n3962), .ZN(n4253) );
  INV_X1 U4668 ( .A(n4253), .ZN(n3976) );
  AOI21_X1 U4669 ( .B1(n3963), .B2(n3962), .A(n3961), .ZN(n3968) );
  OAI22_X1 U4670 ( .A1(n3964), .A2(n4158), .B1(n4215), .B2(n3971), .ZN(n3965)
         );
  AOI21_X1 U4671 ( .B1(n3966), .B2(n4194), .A(n3965), .ZN(n3967) );
  OAI21_X1 U4672 ( .B1(n3968), .B2(n4199), .A(n3967), .ZN(n4252) );
  INV_X1 U4673 ( .A(n3969), .ZN(n3970) );
  OAI21_X1 U4674 ( .B1(n3987), .B2(n3971), .A(n3970), .ZN(n4320) );
  AOI22_X1 U4675 ( .A1(n3972), .A2(n4565), .B1(REG2_REG_27__SCAN_IN), .B2(
        n4564), .ZN(n3973) );
  OAI21_X1 U4676 ( .B1(n4320), .B2(n4204), .A(n3973), .ZN(n3974) );
  AOI21_X1 U4677 ( .B1(n4252), .B2(n4207), .A(n3974), .ZN(n3975) );
  OAI21_X1 U4678 ( .B1(n3976), .B2(n4211), .A(n3975), .ZN(U3263) );
  XOR2_X1 U4679 ( .A(n3980), .B(n3977), .Z(n4257) );
  INV_X1 U4680 ( .A(n4257), .ZN(n3994) );
  NOR2_X1 U4681 ( .A1(n3979), .A2(n3978), .ZN(n3981) );
  XNOR2_X1 U4682 ( .A(n3981), .B(n3980), .ZN(n3986) );
  NOR2_X1 U4683 ( .A1(n3988), .A2(n4215), .ZN(n3982) );
  AOI21_X1 U4684 ( .B1(n3983), .B2(n4194), .A(n3982), .ZN(n3985) );
  NAND2_X1 U4685 ( .A1(n4024), .A2(n4219), .ZN(n3984) );
  OAI211_X1 U4686 ( .C1(n3986), .C2(n4199), .A(n3985), .B(n3984), .ZN(n4256)
         );
  INV_X1 U4687 ( .A(n4009), .ZN(n3989) );
  OAI21_X1 U4688 ( .B1(n3989), .B2(n3988), .A(n2329), .ZN(n4324) );
  AOI22_X1 U4689 ( .A1(n4564), .A2(REG2_REG_26__SCAN_IN), .B1(n3990), .B2(
        n4565), .ZN(n3991) );
  OAI21_X1 U4690 ( .B1(n4324), .B2(n4204), .A(n3991), .ZN(n3992) );
  AOI21_X1 U4691 ( .B1(n4256), .B2(n4207), .A(n3992), .ZN(n3993) );
  OAI21_X1 U4692 ( .B1(n3994), .B2(n4211), .A(n3993), .ZN(U3264) );
  XOR2_X1 U4693 ( .A(n3999), .B(n3995), .Z(n4261) );
  INV_X1 U4694 ( .A(n4261), .ZN(n4016) );
  INV_X1 U4695 ( .A(n3996), .ZN(n3997) );
  OR2_X1 U4696 ( .A1(n3998), .A2(n3997), .ZN(n4000) );
  XNOR2_X1 U4697 ( .A(n4000), .B(n3999), .ZN(n4001) );
  NAND2_X1 U4698 ( .A1(n4001), .A2(n4223), .ZN(n4008) );
  NAND2_X1 U4699 ( .A1(n4002), .A2(n4194), .ZN(n4006) );
  AOI22_X1 U4700 ( .A1(n4004), .A2(n4219), .B1(n4003), .B2(n4244), .ZN(n4005)
         );
  AND2_X1 U4701 ( .A1(n4006), .A2(n4005), .ZN(n4007) );
  NAND2_X1 U4702 ( .A1(n4008), .A2(n4007), .ZN(n4260) );
  INV_X1 U4703 ( .A(n4029), .ZN(n4011) );
  OAI21_X1 U4704 ( .B1(n4011), .B2(n4010), .A(n4009), .ZN(n4328) );
  AOI22_X1 U4705 ( .A1(n4564), .A2(REG2_REG_25__SCAN_IN), .B1(n4012), .B2(
        n4565), .ZN(n4013) );
  OAI21_X1 U4706 ( .B1(n4328), .B2(n4204), .A(n4013), .ZN(n4014) );
  AOI21_X1 U4707 ( .B1(n4260), .B2(n4207), .A(n4014), .ZN(n4015) );
  OAI21_X1 U4708 ( .B1(n4016), .B2(n4211), .A(n4015), .ZN(U3265) );
  XNOR2_X1 U4709 ( .A(n4017), .B(n4020), .ZN(n4265) );
  INV_X1 U4710 ( .A(n4265), .ZN(n4035) );
  NAND2_X1 U4711 ( .A1(n4019), .A2(n4018), .ZN(n4021) );
  XNOR2_X1 U4712 ( .A(n4021), .B(n4020), .ZN(n4026) );
  OAI22_X1 U4713 ( .A1(n4022), .A2(n4158), .B1(n4215), .B2(n4027), .ZN(n4023)
         );
  AOI21_X1 U4714 ( .B1(n4194), .B2(n4024), .A(n4023), .ZN(n4025) );
  OAI21_X1 U4715 ( .B1(n4026), .B2(n4199), .A(n4025), .ZN(n4264) );
  OR2_X1 U4716 ( .A1(n4050), .A2(n4027), .ZN(n4028) );
  NAND2_X1 U4717 ( .A1(n4029), .A2(n4028), .ZN(n4332) );
  INV_X1 U4718 ( .A(n4030), .ZN(n4031) );
  AOI22_X1 U4719 ( .A1(n4564), .A2(REG2_REG_24__SCAN_IN), .B1(n4031), .B2(
        n4565), .ZN(n4032) );
  OAI21_X1 U4720 ( .B1(n4332), .B2(n4204), .A(n4032), .ZN(n4033) );
  AOI21_X1 U4721 ( .B1(n4264), .B2(n4207), .A(n4033), .ZN(n4034) );
  OAI21_X1 U4722 ( .B1(n4035), .B2(n4211), .A(n4034), .ZN(U3266) );
  XNOR2_X1 U4723 ( .A(n4037), .B(n4036), .ZN(n4269) );
  INV_X1 U4724 ( .A(n4269), .ZN(n4056) );
  INV_X1 U4725 ( .A(n4078), .ZN(n4040) );
  INV_X1 U4726 ( .A(n4038), .ZN(n4039) );
  AOI21_X1 U4727 ( .B1(n4040), .B2(n4075), .A(n4039), .ZN(n4059) );
  OAI21_X1 U4728 ( .B1(n4059), .B2(n4058), .A(n4041), .ZN(n4043) );
  XNOR2_X1 U4729 ( .A(n4043), .B(n4042), .ZN(n4047) );
  OAI22_X1 U4730 ( .A1(n4044), .A2(n4216), .B1(n4048), .B2(n4215), .ZN(n4045)
         );
  AOI21_X1 U4731 ( .B1(n4219), .B2(n4081), .A(n4045), .ZN(n4046) );
  OAI21_X1 U4732 ( .B1(n4047), .B2(n4199), .A(n4046), .ZN(n4268) );
  NOR2_X1 U4733 ( .A1(n4066), .A2(n4048), .ZN(n4049) );
  INV_X1 U4734 ( .A(n4051), .ZN(n4052) );
  AOI22_X1 U4735 ( .A1(n4564), .A2(REG2_REG_23__SCAN_IN), .B1(n4052), .B2(
        n4565), .ZN(n4053) );
  OAI21_X1 U4736 ( .B1(n4336), .B2(n4204), .A(n4053), .ZN(n4054) );
  AOI21_X1 U4737 ( .B1(n4268), .B2(n4207), .A(n4054), .ZN(n4055) );
  OAI21_X1 U4738 ( .B1(n4056), .B2(n4211), .A(n4055), .ZN(U3267) );
  AOI21_X1 U4739 ( .B1(n2414), .B2(n4057), .A(n2238), .ZN(n4273) );
  INV_X1 U4740 ( .A(n4273), .ZN(n4074) );
  XNOR2_X1 U4741 ( .A(n4059), .B(n4058), .ZN(n4060) );
  NAND2_X1 U4742 ( .A1(n4060), .A2(n4223), .ZN(n4064) );
  NOR2_X1 U4743 ( .A1(n4068), .A2(n4215), .ZN(n4061) );
  AOI21_X1 U4744 ( .B1(n4062), .B2(n4194), .A(n4061), .ZN(n4063) );
  OAI211_X1 U4745 ( .C1(n4065), .C2(n4158), .A(n4064), .B(n4063), .ZN(n4272)
         );
  INV_X1 U4746 ( .A(n4066), .ZN(n4067) );
  OAI21_X1 U4747 ( .B1(n4084), .B2(n4068), .A(n4067), .ZN(n4340) );
  NOR2_X1 U4748 ( .A1(n4340), .A2(n4204), .ZN(n4072) );
  INV_X1 U4749 ( .A(REG2_REG_22__SCAN_IN), .ZN(n4070) );
  OAI22_X1 U4750 ( .A1(n4207), .A2(n4070), .B1(n4069), .B2(n4231), .ZN(n4071)
         );
  AOI211_X1 U4751 ( .C1(n4272), .C2(n4207), .A(n4072), .B(n4071), .ZN(n4073)
         );
  OAI21_X1 U4752 ( .B1(n4074), .B2(n4211), .A(n4073), .ZN(U3268) );
  XNOR2_X1 U4753 ( .A(n4076), .B(n4075), .ZN(n4277) );
  INV_X1 U4754 ( .A(n4277), .ZN(n4093) );
  XNOR2_X1 U4755 ( .A(n4078), .B(n4077), .ZN(n4079) );
  NAND2_X1 U4756 ( .A1(n4079), .A2(n4223), .ZN(n4083) );
  NOR2_X1 U4757 ( .A1(n4086), .A2(n4215), .ZN(n4080) );
  AOI21_X1 U4758 ( .B1(n4081), .B2(n4194), .A(n4080), .ZN(n4082) );
  OAI211_X1 U4759 ( .C1(n2270), .C2(n4158), .A(n4083), .B(n4082), .ZN(n4276)
         );
  INV_X1 U4760 ( .A(n4109), .ZN(n4087) );
  INV_X1 U4761 ( .A(n4084), .ZN(n4085) );
  OAI21_X1 U4762 ( .B1(n4087), .B2(n4086), .A(n4085), .ZN(n4344) );
  NOR2_X1 U4763 ( .A1(n4344), .A2(n4204), .ZN(n4091) );
  INV_X1 U4764 ( .A(REG2_REG_21__SCAN_IN), .ZN(n4089) );
  OAI22_X1 U4765 ( .A1(n4207), .A2(n4089), .B1(n4088), .B2(n4231), .ZN(n4090)
         );
  AOI211_X1 U4766 ( .C1(n4276), .C2(n4207), .A(n4091), .B(n4090), .ZN(n4092)
         );
  OAI21_X1 U4767 ( .B1(n4093), .B2(n4211), .A(n4092), .ZN(U3269) );
  XNOR2_X1 U4768 ( .A(n4094), .B(n4099), .ZN(n4280) );
  OAI21_X1 U4769 ( .B1(n4152), .B2(n4096), .A(n4095), .ZN(n4134) );
  AOI21_X1 U4770 ( .B1(n4134), .B2(n4098), .A(n4097), .ZN(n4100) );
  XNOR2_X1 U4771 ( .A(n4100), .B(n4099), .ZN(n4105) );
  AOI22_X1 U4772 ( .A1(n4101), .A2(n4194), .B1(n4244), .B2(n4107), .ZN(n4102)
         );
  OAI21_X1 U4773 ( .B1(n4103), .B2(n4158), .A(n4102), .ZN(n4104) );
  AOI21_X1 U4774 ( .B1(n4105), .B2(n4223), .A(n4104), .ZN(n4106) );
  OAI21_X1 U4775 ( .B1(n4280), .B2(n4227), .A(n4106), .ZN(n4281) );
  NAND2_X1 U4776 ( .A1(n4281), .A2(n4207), .ZN(n4115) );
  NAND2_X1 U4777 ( .A1(n2225), .A2(n4107), .ZN(n4108) );
  NAND2_X1 U4778 ( .A1(n4109), .A2(n4108), .ZN(n4348) );
  INV_X1 U4779 ( .A(n4348), .ZN(n4113) );
  INV_X1 U4780 ( .A(REG2_REG_20__SCAN_IN), .ZN(n4111) );
  OAI22_X1 U4781 ( .A1(n4207), .A2(n4111), .B1(n4110), .B2(n4231), .ZN(n4112)
         );
  AOI21_X1 U4782 ( .B1(n4113), .B2(n4569), .A(n4112), .ZN(n4114) );
  OAI211_X1 U4783 ( .C1(n4280), .C2(n4237), .A(n4115), .B(n4114), .ZN(U3270)
         );
  XNOR2_X1 U4784 ( .A(n4116), .B(n4120), .ZN(n4286) );
  INV_X1 U4785 ( .A(n4286), .ZN(n4131) );
  OAI21_X1 U4786 ( .B1(n4134), .B2(n4118), .A(n4117), .ZN(n4119) );
  XOR2_X1 U4787 ( .A(n4120), .B(n4119), .Z(n4125) );
  NOR2_X1 U4788 ( .A1(n4126), .A2(n4215), .ZN(n4121) );
  AOI21_X1 U4789 ( .B1(n4122), .B2(n4194), .A(n4121), .ZN(n4124) );
  NAND2_X1 U4790 ( .A1(n4155), .A2(n4219), .ZN(n4123) );
  OAI211_X1 U4791 ( .C1(n4125), .C2(n4199), .A(n4124), .B(n4123), .ZN(n4285)
         );
  OAI21_X1 U4792 ( .B1(n2330), .B2(n4126), .A(n2225), .ZN(n4352) );
  NOR2_X1 U4793 ( .A1(n4352), .A2(n4204), .ZN(n4129) );
  OAI22_X1 U4794 ( .A1(n4207), .A2(n3936), .B1(n4127), .B2(n4231), .ZN(n4128)
         );
  AOI211_X1 U4795 ( .C1(n4285), .C2(n4207), .A(n4129), .B(n4128), .ZN(n4130)
         );
  OAI21_X1 U4796 ( .B1(n4131), .B2(n4211), .A(n4130), .ZN(U3271) );
  OAI211_X1 U4797 ( .C1(n4160), .C2(n4133), .A(n4629), .B(n4132), .ZN(n4288)
         );
  XOR2_X1 U4798 ( .A(n4143), .B(n4134), .Z(n4140) );
  AOI22_X1 U4799 ( .A1(n4136), .A2(n4194), .B1(n4135), .B2(n4244), .ZN(n4137)
         );
  OAI21_X1 U4800 ( .B1(n4138), .B2(n4158), .A(n4137), .ZN(n4139) );
  AOI21_X1 U4801 ( .B1(n4140), .B2(n4223), .A(n4139), .ZN(n4289) );
  OAI21_X1 U4802 ( .B1(n4377), .B2(n4288), .A(n4289), .ZN(n4148) );
  OAI22_X1 U4803 ( .A1(n4207), .A2(n3889), .B1(n4141), .B2(n4231), .ZN(n4147)
         );
  OAI21_X1 U4804 ( .B1(n4144), .B2(n4143), .A(n4142), .ZN(n4145) );
  INV_X1 U4805 ( .A(n4145), .ZN(n4290) );
  NOR2_X1 U4806 ( .A1(n4290), .A2(n4211), .ZN(n4146) );
  AOI211_X1 U4807 ( .C1(n4207), .C2(n4148), .A(n4147), .B(n4146), .ZN(n4149)
         );
  INV_X1 U4808 ( .A(n4149), .ZN(U3272) );
  XOR2_X1 U4809 ( .A(n4151), .B(n4150), .Z(n4292) );
  INV_X1 U4810 ( .A(n4292), .ZN(n4168) );
  XNOR2_X1 U4811 ( .A(n4152), .B(n4151), .ZN(n4153) );
  NAND2_X1 U4812 ( .A1(n4153), .A2(n4223), .ZN(n4157) );
  NOR2_X1 U4813 ( .A1(n4162), .A2(n4215), .ZN(n4154) );
  AOI21_X1 U4814 ( .B1(n4155), .B2(n4194), .A(n4154), .ZN(n4156) );
  OAI211_X1 U4815 ( .C1(n4159), .C2(n4158), .A(n4157), .B(n4156), .ZN(n4291)
         );
  INV_X1 U4816 ( .A(n4160), .ZN(n4161) );
  OAI21_X1 U4817 ( .B1(n4178), .B2(n4162), .A(n4161), .ZN(n4357) );
  NOR2_X1 U4818 ( .A1(n4357), .A2(n4204), .ZN(n4166) );
  INV_X1 U4819 ( .A(REG2_REG_17__SCAN_IN), .ZN(n4164) );
  OAI22_X1 U4820 ( .A1(n4207), .A2(n4164), .B1(n4163), .B2(n4231), .ZN(n4165)
         );
  AOI211_X1 U4821 ( .C1(n4291), .C2(n4207), .A(n4166), .B(n4165), .ZN(n4167)
         );
  OAI21_X1 U4822 ( .B1(n4168), .B2(n4211), .A(n4167), .ZN(U3273) );
  XNOR2_X1 U4823 ( .A(n4170), .B(n4169), .ZN(n4175) );
  NAND2_X1 U4824 ( .A1(n4171), .A2(n4219), .ZN(n4173) );
  NAND2_X1 U4825 ( .A1(n4389), .A2(n4194), .ZN(n4172) );
  OAI211_X1 U4826 ( .C1(n4215), .C2(n4386), .A(n4173), .B(n4172), .ZN(n4174)
         );
  AOI21_X1 U4827 ( .B1(n4175), .B2(n4223), .A(n4174), .ZN(n4296) );
  AND2_X1 U4828 ( .A1(n4201), .A2(n4176), .ZN(n4177) );
  NOR2_X1 U4829 ( .A1(n4178), .A2(n4177), .ZN(n4358) );
  OAI22_X1 U4830 ( .A1(n4207), .A2(n4526), .B1(n4400), .B2(n4231), .ZN(n4184)
         );
  NAND2_X1 U4831 ( .A1(n4181), .A2(n4180), .ZN(n4182) );
  NAND2_X1 U4832 ( .A1(n4179), .A2(n4182), .ZN(n4295) );
  NOR2_X1 U4833 ( .A1(n4295), .A2(n4211), .ZN(n4183) );
  AOI211_X1 U4834 ( .C1(n4358), .C2(n4569), .A(n4184), .B(n4183), .ZN(n4185)
         );
  OAI21_X1 U4835 ( .B1(n4564), .B2(n4296), .A(n4185), .ZN(U3274) );
  NAND2_X1 U4836 ( .A1(n4187), .A2(n4186), .ZN(n4214) );
  NOR2_X1 U4837 ( .A1(n4214), .A2(n4222), .ZN(n4213) );
  NOR2_X1 U4838 ( .A1(n4213), .A2(n4188), .ZN(n4189) );
  XOR2_X1 U4839 ( .A(n4191), .B(n4189), .Z(n4302) );
  INV_X1 U4840 ( .A(n4302), .ZN(n4212) );
  NAND2_X1 U4841 ( .A1(n4220), .A2(n4190), .ZN(n4192) );
  XNOR2_X1 U4842 ( .A(n4192), .B(n4191), .ZN(n4200) );
  NOR2_X1 U4843 ( .A1(n4202), .A2(n4215), .ZN(n4193) );
  AOI21_X1 U4844 ( .B1(n4195), .B2(n4194), .A(n4193), .ZN(n4198) );
  NAND2_X1 U4845 ( .A1(n4196), .A2(n4219), .ZN(n4197) );
  OAI211_X1 U4846 ( .C1(n4200), .C2(n4199), .A(n4198), .B(n4197), .ZN(n4301)
         );
  INV_X1 U4847 ( .A(n4228), .ZN(n4203) );
  OAI21_X1 U4848 ( .B1(n4203), .B2(n4202), .A(n4201), .ZN(n4367) );
  NOR2_X1 U4849 ( .A1(n4367), .A2(n4204), .ZN(n4209) );
  INV_X1 U4850 ( .A(REG2_REG_15__SCAN_IN), .ZN(n4206) );
  OAI22_X1 U4851 ( .A1(n4207), .A2(n4206), .B1(n4205), .B2(n4231), .ZN(n4208)
         );
  AOI211_X1 U4852 ( .C1(n4301), .C2(n4207), .A(n4209), .B(n4208), .ZN(n4210)
         );
  OAI21_X1 U4853 ( .B1(n4212), .B2(n4211), .A(n4210), .ZN(U3275) );
  AOI21_X1 U4854 ( .B1(n4222), .B2(n4214), .A(n4213), .ZN(n4304) );
  OAI22_X1 U4855 ( .A1(n4385), .A2(n4216), .B1(n4215), .B2(n4229), .ZN(n4217)
         );
  AOI21_X1 U4856 ( .B1(n4219), .B2(n4218), .A(n4217), .ZN(n4226) );
  OAI21_X1 U4857 ( .B1(n4222), .B2(n4221), .A(n4220), .ZN(n4224) );
  NAND2_X1 U4858 ( .A1(n4224), .A2(n4223), .ZN(n4225) );
  OAI211_X1 U4859 ( .C1(n4304), .C2(n4227), .A(n4226), .B(n4225), .ZN(n4305)
         );
  NAND2_X1 U4860 ( .A1(n4305), .A2(n4207), .ZN(n4236) );
  OAI21_X1 U4861 ( .B1(n4230), .B2(n4229), .A(n4228), .ZN(n4372) );
  INV_X1 U4862 ( .A(n4372), .ZN(n4234) );
  OAI22_X1 U4863 ( .A1(n4207), .A2(n4509), .B1(n4232), .B2(n4231), .ZN(n4233)
         );
  AOI21_X1 U4864 ( .B1(n4234), .B2(n4569), .A(n4233), .ZN(n4235) );
  OAI211_X1 U4865 ( .C1(n4304), .C2(n4237), .A(n4236), .B(n4235), .ZN(U3276)
         );
  NAND2_X1 U4866 ( .A1(n4312), .A2(n4646), .ZN(n4239) );
  NAND2_X1 U4867 ( .A1(n4643), .A2(REG1_REG_31__SCAN_IN), .ZN(n4238) );
  OAI211_X1 U4868 ( .C1(n4314), .C2(n4309), .A(n4239), .B(n4238), .ZN(U3549)
         );
  AOI21_X1 U4869 ( .B1(n4245), .B2(n4241), .A(n4240), .ZN(n4402) );
  INV_X1 U4870 ( .A(n4402), .ZN(n4316) );
  INV_X1 U4871 ( .A(REG1_REG_30__SCAN_IN), .ZN(n4246) );
  INV_X1 U4872 ( .A(n4242), .ZN(n4243) );
  AOI21_X1 U4873 ( .B1(n4245), .B2(n4244), .A(n4243), .ZN(n4404) );
  MUX2_X1 U4874 ( .A(n4246), .B(n4404), .S(n4646), .Z(n4247) );
  OAI21_X1 U4875 ( .B1(n4316), .B2(n4309), .A(n4247), .ZN(U3548) );
  INV_X1 U4876 ( .A(n4249), .ZN(n4250) );
  OAI21_X1 U4877 ( .B1(n4309), .B2(n4251), .A(n4250), .ZN(U3546) );
  INV_X1 U4878 ( .A(REG1_REG_27__SCAN_IN), .ZN(n4254) );
  AOI21_X1 U4879 ( .B1(n4253), .B2(n4622), .A(n4252), .ZN(n4317) );
  MUX2_X1 U4880 ( .A(n4254), .B(n4317), .S(n4646), .Z(n4255) );
  OAI21_X1 U4881 ( .B1(n4309), .B2(n4320), .A(n4255), .ZN(U3545) );
  INV_X1 U4882 ( .A(REG1_REG_26__SCAN_IN), .ZN(n4258) );
  AOI21_X1 U4883 ( .B1(n4257), .B2(n4622), .A(n4256), .ZN(n4321) );
  MUX2_X1 U4884 ( .A(n4258), .B(n4321), .S(n4646), .Z(n4259) );
  OAI21_X1 U4885 ( .B1(n4309), .B2(n4324), .A(n4259), .ZN(U3544) );
  INV_X1 U4886 ( .A(REG1_REG_25__SCAN_IN), .ZN(n4262) );
  AOI21_X1 U4887 ( .B1(n4261), .B2(n4622), .A(n4260), .ZN(n4325) );
  MUX2_X1 U4888 ( .A(n4262), .B(n4325), .S(n4646), .Z(n4263) );
  OAI21_X1 U4889 ( .B1(n4309), .B2(n4328), .A(n4263), .ZN(U3543) );
  INV_X1 U4890 ( .A(REG1_REG_24__SCAN_IN), .ZN(n4266) );
  AOI21_X1 U4891 ( .B1(n4265), .B2(n4622), .A(n4264), .ZN(n4329) );
  MUX2_X1 U4892 ( .A(n4266), .B(n4329), .S(n4646), .Z(n4267) );
  OAI21_X1 U4893 ( .B1(n4309), .B2(n4332), .A(n4267), .ZN(U3542) );
  INV_X1 U4894 ( .A(REG1_REG_23__SCAN_IN), .ZN(n4270) );
  AOI21_X1 U4895 ( .B1(n4269), .B2(n4622), .A(n4268), .ZN(n4333) );
  MUX2_X1 U4896 ( .A(n4270), .B(n4333), .S(n4646), .Z(n4271) );
  OAI21_X1 U4897 ( .B1(n4309), .B2(n4336), .A(n4271), .ZN(U3541) );
  INV_X1 U4898 ( .A(REG1_REG_22__SCAN_IN), .ZN(n4274) );
  AOI21_X1 U4899 ( .B1(n4273), .B2(n4622), .A(n4272), .ZN(n4337) );
  MUX2_X1 U4900 ( .A(n4274), .B(n4337), .S(n4646), .Z(n4275) );
  OAI21_X1 U4901 ( .B1(n4309), .B2(n4340), .A(n4275), .ZN(U3540) );
  INV_X1 U4902 ( .A(REG1_REG_21__SCAN_IN), .ZN(n4278) );
  AOI21_X1 U4903 ( .B1(n4277), .B2(n4622), .A(n4276), .ZN(n4341) );
  MUX2_X1 U4904 ( .A(n4278), .B(n4341), .S(n4646), .Z(n4279) );
  OAI21_X1 U4905 ( .B1(n4309), .B2(n4344), .A(n4279), .ZN(U3539) );
  INV_X1 U4906 ( .A(REG1_REG_20__SCAN_IN), .ZN(n4283) );
  INV_X1 U4907 ( .A(n4280), .ZN(n4282) );
  AOI21_X1 U4908 ( .B1(n4618), .B2(n4282), .A(n4281), .ZN(n4345) );
  MUX2_X1 U4909 ( .A(n4283), .B(n4345), .S(n4646), .Z(n4284) );
  OAI21_X1 U4910 ( .B1(n4309), .B2(n4348), .A(n4284), .ZN(U3538) );
  AOI21_X1 U4911 ( .B1(n4286), .B2(n4622), .A(n4285), .ZN(n4349) );
  MUX2_X1 U4912 ( .A(n3932), .B(n4349), .S(n4646), .Z(n4287) );
  OAI21_X1 U4913 ( .B1(n4309), .B2(n4352), .A(n4287), .ZN(U3537) );
  OAI211_X1 U4914 ( .C1(n4290), .C2(n4294), .A(n4289), .B(n4288), .ZN(n4353)
         );
  MUX2_X1 U4915 ( .A(REG1_REG_18__SCAN_IN), .B(n4353), .S(n4646), .Z(U3536) );
  AOI21_X1 U4916 ( .B1(n4292), .B2(n4622), .A(n4291), .ZN(n4354) );
  MUX2_X1 U4917 ( .A(n3886), .B(n4354), .S(n4646), .Z(n4293) );
  OAI21_X1 U4918 ( .B1(n4309), .B2(n4357), .A(n4293), .ZN(U3535) );
  OR2_X1 U4919 ( .A1(n4295), .A2(n4294), .ZN(n4297) );
  NAND2_X1 U4920 ( .A1(n4297), .A2(n4296), .ZN(n4359) );
  MUX2_X1 U4921 ( .A(REG1_REG_16__SCAN_IN), .B(n4359), .S(n4646), .Z(n4298) );
  AOI21_X1 U4922 ( .B1(n4299), .B2(n4358), .A(n4298), .ZN(n4300) );
  INV_X1 U4923 ( .A(n4300), .ZN(U3534) );
  AOI21_X1 U4924 ( .B1(n4302), .B2(n4622), .A(n4301), .ZN(n4364) );
  MUX2_X1 U4925 ( .A(n3865), .B(n4364), .S(n4646), .Z(n4303) );
  OAI21_X1 U4926 ( .B1(n4309), .B2(n4367), .A(n4303), .ZN(U3533) );
  INV_X1 U4927 ( .A(REG1_REG_14__SCAN_IN), .ZN(n4307) );
  INV_X1 U4928 ( .A(n4304), .ZN(n4306) );
  AOI21_X1 U4929 ( .B1(n4618), .B2(n4306), .A(n4305), .ZN(n4368) );
  MUX2_X1 U4930 ( .A(n4307), .B(n4368), .S(n4646), .Z(n4308) );
  OAI21_X1 U4931 ( .B1(n4309), .B2(n4372), .A(n4308), .ZN(U3532) );
  NOR2_X1 U4932 ( .A1(n4631), .A2(n4310), .ZN(n4311) );
  AOI21_X1 U4933 ( .B1(n4631), .B2(n4312), .A(n4311), .ZN(n4313) );
  OAI21_X1 U4934 ( .B1(n4314), .B2(n4371), .A(n4313), .ZN(U3517) );
  MUX2_X1 U4935 ( .A(n2823), .B(n4404), .S(n4631), .Z(n4315) );
  OAI21_X1 U4936 ( .B1(n4316), .B2(n4371), .A(n4315), .ZN(U3516) );
  INV_X1 U4937 ( .A(REG0_REG_27__SCAN_IN), .ZN(n4318) );
  MUX2_X1 U4938 ( .A(n4318), .B(n4317), .S(n4631), .Z(n4319) );
  OAI21_X1 U4939 ( .B1(n4320), .B2(n4371), .A(n4319), .ZN(U3513) );
  INV_X1 U4940 ( .A(REG0_REG_26__SCAN_IN), .ZN(n4322) );
  MUX2_X1 U4941 ( .A(n4322), .B(n4321), .S(n4631), .Z(n4323) );
  OAI21_X1 U4942 ( .B1(n4324), .B2(n4371), .A(n4323), .ZN(U3512) );
  MUX2_X1 U4943 ( .A(n4326), .B(n4325), .S(n4631), .Z(n4327) );
  OAI21_X1 U4944 ( .B1(n4328), .B2(n4371), .A(n4327), .ZN(U3511) );
  MUX2_X1 U4945 ( .A(n4330), .B(n4329), .S(n4631), .Z(n4331) );
  OAI21_X1 U4946 ( .B1(n4332), .B2(n4371), .A(n4331), .ZN(U3510) );
  MUX2_X1 U4947 ( .A(n4334), .B(n4333), .S(n4631), .Z(n4335) );
  OAI21_X1 U4948 ( .B1(n4336), .B2(n4371), .A(n4335), .ZN(U3509) );
  MUX2_X1 U4949 ( .A(n4338), .B(n4337), .S(n4631), .Z(n4339) );
  OAI21_X1 U4950 ( .B1(n4340), .B2(n4371), .A(n4339), .ZN(U3508) );
  MUX2_X1 U4951 ( .A(n4342), .B(n4341), .S(n4631), .Z(n4343) );
  OAI21_X1 U4952 ( .B1(n4344), .B2(n4371), .A(n4343), .ZN(U3507) );
  MUX2_X1 U4953 ( .A(n4346), .B(n4345), .S(n4631), .Z(n4347) );
  OAI21_X1 U4954 ( .B1(n4348), .B2(n4371), .A(n4347), .ZN(U3506) );
  MUX2_X1 U4955 ( .A(n4350), .B(n4349), .S(n4631), .Z(n4351) );
  OAI21_X1 U4956 ( .B1(n4352), .B2(n4371), .A(n4351), .ZN(U3505) );
  MUX2_X1 U4957 ( .A(REG0_REG_18__SCAN_IN), .B(n4353), .S(n4631), .Z(U3503) );
  MUX2_X1 U4958 ( .A(n4355), .B(n4354), .S(n4631), .Z(n4356) );
  OAI21_X1 U4959 ( .B1(n4357), .B2(n4371), .A(n4356), .ZN(U3501) );
  INV_X1 U4960 ( .A(n4358), .ZN(n4363) );
  INV_X1 U4961 ( .A(n4359), .ZN(n4361) );
  MUX2_X1 U4962 ( .A(n4361), .B(n4360), .S(n4630), .Z(n4362) );
  OAI21_X1 U4963 ( .B1(n4363), .B2(n4371), .A(n4362), .ZN(U3499) );
  MUX2_X1 U4964 ( .A(n4365), .B(n4364), .S(n4631), .Z(n4366) );
  OAI21_X1 U4965 ( .B1(n4367), .B2(n4371), .A(n4366), .ZN(U3497) );
  MUX2_X1 U4966 ( .A(n4369), .B(n4368), .S(n4631), .Z(n4370) );
  OAI21_X1 U4967 ( .B1(n4372), .B2(n4371), .A(n4370), .ZN(U3495) );
  MUX2_X1 U4968 ( .A(DATAI_30_), .B(n4373), .S(STATE_REG_SCAN_IN), .Z(U3322)
         );
  MUX2_X1 U4969 ( .A(n2795), .B(DATAI_26_), .S(U3149), .Z(U3326) );
  MUX2_X1 U4970 ( .A(n4374), .B(DATAI_24_), .S(U3149), .Z(U3328) );
  MUX2_X1 U4971 ( .A(DATAI_22_), .B(n4375), .S(STATE_REG_SCAN_IN), .Z(U3330)
         );
  MUX2_X1 U4972 ( .A(DATAI_20_), .B(n4376), .S(STATE_REG_SCAN_IN), .Z(U3332)
         );
  MUX2_X1 U4973 ( .A(n4377), .B(DATAI_19_), .S(U3149), .Z(U3333) );
  MUX2_X1 U4974 ( .A(n4378), .B(DATAI_18_), .S(U3149), .Z(U3334) );
  MUX2_X1 U4975 ( .A(DATAI_4_), .B(n4379), .S(STATE_REG_SCAN_IN), .Z(U3348) );
  MUX2_X1 U4976 ( .A(DATAI_3_), .B(n4380), .S(STATE_REG_SCAN_IN), .Z(U3349) );
  MUX2_X1 U4977 ( .A(n4381), .B(DATAI_2_), .S(U3149), .Z(U3350) );
  MUX2_X1 U4978 ( .A(n2482), .B(DATAI_1_), .S(U3149), .Z(U3351) );
  INV_X1 U4979 ( .A(DATAI_28_), .ZN(n4720) );
  AOI22_X1 U4980 ( .A1(STATE_REG_SCAN_IN), .A2(n4382), .B1(n4720), .B2(U3149), 
        .ZN(U3324) );
  NOR2_X1 U4981 ( .A1(STATE_REG_SCAN_IN), .A2(n4383), .ZN(n4530) );
  OAI22_X1 U4982 ( .A1(n4387), .A2(n4386), .B1(n4385), .B2(n4384), .ZN(n4388)
         );
  AOI211_X1 U4983 ( .C1(n4390), .C2(n4389), .A(n4530), .B(n4388), .ZN(n4399)
         );
  INV_X1 U4984 ( .A(n3618), .ZN(n4393) );
  OAI21_X1 U4985 ( .B1(n4393), .B2(n4392), .A(n4391), .ZN(n4395) );
  XNOR2_X1 U4986 ( .A(n4395), .B(n4394), .ZN(n4397) );
  NAND2_X1 U4987 ( .A1(n4397), .A2(n4396), .ZN(n4398) );
  OAI211_X1 U4988 ( .C1(n4401), .C2(n4400), .A(n4399), .B(n4398), .ZN(U3223)
         );
  AOI22_X1 U4989 ( .A1(n4402), .A2(n4569), .B1(REG2_REG_30__SCAN_IN), .B2(
        n4564), .ZN(n4403) );
  OAI21_X1 U4990 ( .B1(n4564), .B2(n4404), .A(n4403), .ZN(U3261) );
  INV_X1 U4991 ( .A(n4407), .ZN(n4405) );
  OAI211_X1 U4992 ( .C1(REG1_REG_0__SCAN_IN), .C2(n4406), .A(n4405), .B(n4408), 
        .ZN(n4411) );
  AOI22_X1 U4993 ( .A1(n4408), .A2(n4407), .B1(n4542), .B2(n2863), .ZN(n4410)
         );
  AOI22_X1 U4994 ( .A1(ADDR_REG_0__SCAN_IN), .A2(n4541), .B1(
        REG3_REG_0__SCAN_IN), .B2(U3149), .ZN(n4409) );
  OAI221_X1 U4995 ( .B1(IR_REG_0__SCAN_IN), .B2(n4411), .C1(n2395), .C2(n4410), 
        .A(n4409), .ZN(U3240) );
  AOI211_X1 U4996 ( .C1(n4414), .C2(n4413), .A(n4412), .B(n4422), .ZN(n4416)
         );
  AOI211_X1 U4997 ( .C1(n4541), .C2(ADDR_REG_5__SCAN_IN), .A(n4416), .B(n4415), 
        .ZN(n4421) );
  OAI211_X1 U4998 ( .C1(n4419), .C2(n4418), .A(n4496), .B(n4417), .ZN(n4420)
         );
  OAI211_X1 U4999 ( .C1(n4548), .C2(n4600), .A(n4421), .B(n4420), .ZN(U3245)
         );
  AOI211_X1 U5000 ( .C1(n4425), .C2(n4424), .A(n4423), .B(n4422), .ZN(n4427)
         );
  AOI211_X1 U5001 ( .C1(n4541), .C2(ADDR_REG_6__SCAN_IN), .A(n4427), .B(n4426), 
        .ZN(n4431) );
  OAI211_X1 U5002 ( .C1(REG2_REG_6__SCAN_IN), .C2(n4429), .A(n4496), .B(n4428), 
        .ZN(n4430) );
  OAI211_X1 U5003 ( .C1(n4548), .C2(n4598), .A(n4431), .B(n4430), .ZN(U3246)
         );
  AOI22_X1 U5004 ( .A1(n4432), .A2(n4641), .B1(REG1_REG_7__SCAN_IN), .B2(n4597), .ZN(n4434) );
  OAI21_X1 U5005 ( .B1(n4435), .B2(n4434), .A(n4542), .ZN(n4433) );
  AOI21_X1 U5006 ( .B1(n4435), .B2(n4434), .A(n4433), .ZN(n4437) );
  AOI211_X1 U5007 ( .C1(n4541), .C2(ADDR_REG_7__SCAN_IN), .A(n4437), .B(n4436), 
        .ZN(n4442) );
  OAI211_X1 U5008 ( .C1(n4440), .C2(n4439), .A(n4496), .B(n4438), .ZN(n4441)
         );
  OAI211_X1 U5009 ( .C1(n4548), .C2(n4597), .A(n4442), .B(n4441), .ZN(U3247)
         );
  OAI211_X1 U5010 ( .C1(REG2_REG_8__SCAN_IN), .C2(n4445), .A(n4496), .B(n4444), 
        .ZN(n4447) );
  NAND2_X1 U5011 ( .A1(n4447), .A2(n4446), .ZN(n4448) );
  AOI21_X1 U5012 ( .B1(n4541), .B2(ADDR_REG_8__SCAN_IN), .A(n4448), .ZN(n4452)
         );
  OAI211_X1 U5013 ( .C1(REG1_REG_8__SCAN_IN), .C2(n4450), .A(n4542), .B(n4449), 
        .ZN(n4451) );
  OAI211_X1 U5014 ( .C1(n4548), .C2(n2279), .A(n4452), .B(n4451), .ZN(U3248)
         );
  OAI211_X1 U5015 ( .C1(n4455), .C2(n4454), .A(n4542), .B(n4453), .ZN(n4460)
         );
  OAI211_X1 U5016 ( .C1(n4458), .C2(n4457), .A(n4496), .B(n4456), .ZN(n4459)
         );
  OAI211_X1 U5017 ( .C1(n4548), .C2(n4596), .A(n4460), .B(n4459), .ZN(n4461)
         );
  AOI211_X1 U5018 ( .C1(n4541), .C2(ADDR_REG_9__SCAN_IN), .A(n4462), .B(n4461), 
        .ZN(n4463) );
  INV_X1 U5019 ( .A(n4463), .ZN(U3249) );
  OAI211_X1 U5020 ( .C1(REG2_REG_10__SCAN_IN), .C2(n4466), .A(n4496), .B(n4465), .ZN(n4468) );
  NAND2_X1 U5021 ( .A1(n4468), .A2(n4467), .ZN(n4469) );
  AOI21_X1 U5022 ( .B1(n4541), .B2(ADDR_REG_10__SCAN_IN), .A(n4469), .ZN(n4473) );
  OAI211_X1 U5023 ( .C1(REG1_REG_10__SCAN_IN), .C2(n4471), .A(n4542), .B(n4470), .ZN(n4472) );
  OAI211_X1 U5024 ( .C1(n4548), .C2(n2281), .A(n4473), .B(n4472), .ZN(U3250)
         );
  OAI211_X1 U5025 ( .C1(n4476), .C2(n4475), .A(n4542), .B(n4474), .ZN(n4481)
         );
  OAI211_X1 U5026 ( .C1(n4479), .C2(n4478), .A(n4496), .B(n4477), .ZN(n4480)
         );
  OAI211_X1 U5027 ( .C1(n4548), .C2(n4595), .A(n4481), .B(n4480), .ZN(n4482)
         );
  AOI211_X1 U5028 ( .C1(n4541), .C2(ADDR_REG_11__SCAN_IN), .A(n4483), .B(n4482), .ZN(n4484) );
  INV_X1 U5029 ( .A(n4484), .ZN(U3251) );
  OAI211_X1 U5030 ( .C1(REG2_REG_12__SCAN_IN), .C2(n4487), .A(n4496), .B(n4486), .ZN(n4489) );
  NAND2_X1 U5031 ( .A1(n4489), .A2(n4488), .ZN(n4490) );
  AOI21_X1 U5032 ( .B1(n4541), .B2(ADDR_REG_12__SCAN_IN), .A(n4490), .ZN(n4494) );
  OAI211_X1 U5033 ( .C1(REG1_REG_12__SCAN_IN), .C2(n4492), .A(n4542), .B(n4491), .ZN(n4493) );
  OAI211_X1 U5034 ( .C1(n4548), .C2(n2280), .A(n4494), .B(n4493), .ZN(U3252)
         );
  AOI21_X1 U5035 ( .B1(n4593), .B2(n3232), .A(n4495), .ZN(n4499) );
  OAI21_X1 U5036 ( .B1(n4499), .B2(n4498), .A(n4496), .ZN(n4497) );
  AOI21_X1 U5037 ( .B1(n4499), .B2(n4498), .A(n4497), .ZN(n4500) );
  AOI211_X1 U5038 ( .C1(n4541), .C2(ADDR_REG_13__SCAN_IN), .A(n4501), .B(n4500), .ZN(n4506) );
  OAI211_X1 U5039 ( .C1(n4504), .C2(n4503), .A(n4542), .B(n4502), .ZN(n4505)
         );
  OAI211_X1 U5040 ( .C1(n4548), .C2(n4593), .A(n4506), .B(n4505), .ZN(U3253)
         );
  AOI211_X1 U5041 ( .C1(n4509), .C2(n4508), .A(n4507), .B(n4535), .ZN(n4510)
         );
  AOI211_X1 U5042 ( .C1(n4541), .C2(ADDR_REG_14__SCAN_IN), .A(n4511), .B(n4510), .ZN(n4515) );
  OAI211_X1 U5043 ( .C1(REG1_REG_14__SCAN_IN), .C2(n4513), .A(n4542), .B(n4512), .ZN(n4514) );
  OAI211_X1 U5044 ( .C1(n4548), .C2(n4592), .A(n4515), .B(n4514), .ZN(U3254)
         );
  AOI211_X1 U5045 ( .C1(n4518), .C2(n4517), .A(n4516), .B(n4535), .ZN(n4519)
         );
  AOI211_X1 U5046 ( .C1(n4541), .C2(ADDR_REG_15__SCAN_IN), .A(n4520), .B(n4519), .ZN(n4525) );
  OAI211_X1 U5047 ( .C1(n4523), .C2(n4522), .A(n4542), .B(n4521), .ZN(n4524)
         );
  OAI211_X1 U5048 ( .C1(n4548), .C2(n4591), .A(n4525), .B(n4524), .ZN(U3255)
         );
  AOI221_X1 U5049 ( .B1(n4528), .B2(n4527), .C1(n4526), .C2(n4527), .A(n4535), 
        .ZN(n4529) );
  AOI211_X1 U5050 ( .C1(n4541), .C2(ADDR_REG_16__SCAN_IN), .A(n4530), .B(n4529), .ZN(n4534) );
  OAI221_X1 U5051 ( .B1(n4532), .B2(REG1_REG_16__SCAN_IN), .C1(n4532), .C2(
        n4531), .A(n4542), .ZN(n4533) );
  OAI211_X1 U5052 ( .C1(n4548), .C2(n4590), .A(n4534), .B(n4533), .ZN(U3256)
         );
  AOI221_X1 U5053 ( .B1(n4538), .B2(n4537), .C1(n4536), .C2(n4537), .A(n4535), 
        .ZN(n4539) );
  AOI211_X1 U5054 ( .C1(n4541), .C2(ADDR_REG_17__SCAN_IN), .A(n4540), .B(n4539), .ZN(n4547) );
  OAI221_X1 U5055 ( .B1(n4545), .B2(n4544), .C1(n4545), .C2(n4543), .A(n4542), 
        .ZN(n4546) );
  OAI211_X1 U5056 ( .C1(n4548), .C2(n4589), .A(n4547), .B(n4546), .ZN(U3257)
         );
  INV_X1 U5057 ( .A(n4549), .ZN(n4550) );
  AOI22_X1 U5058 ( .A1(n4550), .A2(n4565), .B1(REG2_REG_10__SCAN_IN), .B2(
        n4564), .ZN(n4555) );
  INV_X1 U5059 ( .A(n4551), .ZN(n4552) );
  AOI22_X1 U5060 ( .A1(n4553), .A2(n4570), .B1(n4569), .B2(n4552), .ZN(n4554)
         );
  OAI211_X1 U5061 ( .C1(n4564), .C2(n4556), .A(n4555), .B(n4554), .ZN(U3280)
         );
  AOI22_X1 U5062 ( .A1(n4557), .A2(n4565), .B1(REG2_REG_8__SCAN_IN), .B2(n4564), .ZN(n4562) );
  INV_X1 U5063 ( .A(n4558), .ZN(n4559) );
  AOI22_X1 U5064 ( .A1(n4560), .A2(n4570), .B1(n4569), .B2(n4559), .ZN(n4561)
         );
  OAI211_X1 U5065 ( .C1(n4564), .C2(n4563), .A(n4562), .B(n4561), .ZN(U3282)
         );
  AOI22_X1 U5066 ( .A1(n4566), .A2(n4565), .B1(REG2_REG_6__SCAN_IN), .B2(n4564), .ZN(n4573) );
  INV_X1 U5067 ( .A(n4567), .ZN(n4568) );
  AOI22_X1 U5068 ( .A1(n4571), .A2(n4570), .B1(n4569), .B2(n4568), .ZN(n4572)
         );
  OAI211_X1 U5069 ( .C1(n4564), .C2(n4574), .A(n4573), .B(n4572), .ZN(U3284)
         );
  INV_X1 U5070 ( .A(D_REG_31__SCAN_IN), .ZN(n4733) );
  NOR2_X1 U5071 ( .A1(n4587), .A2(n4733), .ZN(U3291) );
  INV_X1 U5072 ( .A(D_REG_30__SCAN_IN), .ZN(n4988) );
  NOR2_X1 U5073 ( .A1(n4587), .A2(n4988), .ZN(U3292) );
  INV_X1 U5074 ( .A(D_REG_29__SCAN_IN), .ZN(n4890) );
  NOR2_X1 U5075 ( .A1(n4587), .A2(n4890), .ZN(U3293) );
  INV_X1 U5076 ( .A(D_REG_28__SCAN_IN), .ZN(n4920) );
  NOR2_X1 U5077 ( .A1(n4587), .A2(n4920), .ZN(U3294) );
  INV_X1 U5078 ( .A(D_REG_27__SCAN_IN), .ZN(n4910) );
  NOR2_X1 U5079 ( .A1(n4587), .A2(n4910), .ZN(U3295) );
  INV_X1 U5080 ( .A(D_REG_26__SCAN_IN), .ZN(n4576) );
  NOR2_X1 U5081 ( .A1(n4587), .A2(n4576), .ZN(U3296) );
  INV_X1 U5082 ( .A(D_REG_25__SCAN_IN), .ZN(n4898) );
  NOR2_X1 U5083 ( .A1(n4587), .A2(n4898), .ZN(U3297) );
  INV_X1 U5084 ( .A(D_REG_24__SCAN_IN), .ZN(n4577) );
  NOR2_X1 U5085 ( .A1(n4587), .A2(n4577), .ZN(U3298) );
  INV_X1 U5086 ( .A(D_REG_23__SCAN_IN), .ZN(n4965) );
  NOR2_X1 U5087 ( .A1(n4587), .A2(n4965), .ZN(U3299) );
  INV_X1 U5088 ( .A(D_REG_22__SCAN_IN), .ZN(n4726) );
  NOR2_X1 U5089 ( .A1(n4587), .A2(n4726), .ZN(U3300) );
  INV_X1 U5090 ( .A(D_REG_21__SCAN_IN), .ZN(n4951) );
  NOR2_X1 U5091 ( .A1(n4587), .A2(n4951), .ZN(U3301) );
  INV_X1 U5092 ( .A(D_REG_20__SCAN_IN), .ZN(n4578) );
  NOR2_X1 U5093 ( .A1(n4587), .A2(n4578), .ZN(U3302) );
  INV_X1 U5094 ( .A(D_REG_19__SCAN_IN), .ZN(n4779) );
  NOR2_X1 U5095 ( .A1(n4587), .A2(n4779), .ZN(U3303) );
  INV_X1 U5096 ( .A(D_REG_18__SCAN_IN), .ZN(n4579) );
  NOR2_X1 U5097 ( .A1(n4587), .A2(n4579), .ZN(U3304) );
  INV_X1 U5098 ( .A(D_REG_17__SCAN_IN), .ZN(n4580) );
  NOR2_X1 U5099 ( .A1(n4587), .A2(n4580), .ZN(U3305) );
  INV_X1 U5100 ( .A(D_REG_16__SCAN_IN), .ZN(n4753) );
  NOR2_X1 U5101 ( .A1(n4587), .A2(n4753), .ZN(U3306) );
  INV_X1 U5102 ( .A(D_REG_15__SCAN_IN), .ZN(n4581) );
  NOR2_X1 U5103 ( .A1(n4587), .A2(n4581), .ZN(U3307) );
  INV_X1 U5104 ( .A(D_REG_14__SCAN_IN), .ZN(n4582) );
  NOR2_X1 U5105 ( .A1(n4587), .A2(n4582), .ZN(U3308) );
  INV_X1 U5106 ( .A(D_REG_13__SCAN_IN), .ZN(n4734) );
  NOR2_X1 U5107 ( .A1(n4587), .A2(n4734), .ZN(U3309) );
  INV_X1 U5108 ( .A(D_REG_12__SCAN_IN), .ZN(n4975) );
  NOR2_X1 U5109 ( .A1(n4587), .A2(n4975), .ZN(U3310) );
  INV_X1 U5110 ( .A(D_REG_11__SCAN_IN), .ZN(n4583) );
  NOR2_X1 U5111 ( .A1(n4587), .A2(n4583), .ZN(U3311) );
  INV_X1 U5112 ( .A(D_REG_10__SCAN_IN), .ZN(n4925) );
  NOR2_X1 U5113 ( .A1(n4587), .A2(n4925), .ZN(U3312) );
  INV_X1 U5114 ( .A(D_REG_9__SCAN_IN), .ZN(n4941) );
  NOR2_X1 U5115 ( .A1(n4587), .A2(n4941), .ZN(U3313) );
  INV_X1 U5116 ( .A(D_REG_8__SCAN_IN), .ZN(n4752) );
  NOR2_X1 U5117 ( .A1(n4587), .A2(n4752), .ZN(U3314) );
  INV_X1 U5118 ( .A(D_REG_7__SCAN_IN), .ZN(n4992) );
  NOR2_X1 U5119 ( .A1(n4587), .A2(n4992), .ZN(U3315) );
  INV_X1 U5120 ( .A(D_REG_6__SCAN_IN), .ZN(n4584) );
  NOR2_X1 U5121 ( .A1(n4587), .A2(n4584), .ZN(U3316) );
  INV_X1 U5122 ( .A(D_REG_5__SCAN_IN), .ZN(n4585) );
  NOR2_X1 U5123 ( .A1(n4587), .A2(n4585), .ZN(U3317) );
  INV_X1 U5124 ( .A(D_REG_4__SCAN_IN), .ZN(n4907) );
  NOR2_X1 U5125 ( .A1(n4587), .A2(n4907), .ZN(U3318) );
  INV_X1 U5126 ( .A(D_REG_3__SCAN_IN), .ZN(n4932) );
  NOR2_X1 U5127 ( .A1(n4587), .A2(n4932), .ZN(U3319) );
  INV_X1 U5128 ( .A(D_REG_2__SCAN_IN), .ZN(n4586) );
  NOR2_X1 U5129 ( .A1(n4587), .A2(n4586), .ZN(U3320) );
  INV_X1 U5130 ( .A(DATAI_23_), .ZN(n4893) );
  AOI21_X1 U5131 ( .B1(U3149), .B2(n4893), .A(n4588), .ZN(U3329) );
  AOI22_X1 U5132 ( .A1(STATE_REG_SCAN_IN), .A2(n4589), .B1(n2660), .B2(U3149), 
        .ZN(U3335) );
  AOI22_X1 U5133 ( .A1(STATE_REG_SCAN_IN), .A2(n4590), .B1(n4989), .B2(U3149), 
        .ZN(U3336) );
  INV_X1 U5134 ( .A(DATAI_15_), .ZN(n4909) );
  AOI22_X1 U5135 ( .A1(STATE_REG_SCAN_IN), .A2(n4591), .B1(n4909), .B2(U3149), 
        .ZN(U3337) );
  AOI22_X1 U5136 ( .A1(STATE_REG_SCAN_IN), .A2(n4592), .B1(n4980), .B2(U3149), 
        .ZN(U3338) );
  INV_X1 U5137 ( .A(DATAI_13_), .ZN(n4894) );
  AOI22_X1 U5138 ( .A1(STATE_REG_SCAN_IN), .A2(n4593), .B1(n4894), .B2(U3149), 
        .ZN(U3339) );
  INV_X1 U5139 ( .A(DATAI_12_), .ZN(n4594) );
  AOI22_X1 U5140 ( .A1(STATE_REG_SCAN_IN), .A2(n2280), .B1(n4594), .B2(U3149), 
        .ZN(U3340) );
  AOI22_X1 U5141 ( .A1(STATE_REG_SCAN_IN), .A2(n4595), .B1(n2600), .B2(U3149), 
        .ZN(U3341) );
  INV_X1 U5142 ( .A(DATAI_10_), .ZN(n4967) );
  AOI22_X1 U5143 ( .A1(STATE_REG_SCAN_IN), .A2(n2281), .B1(n4967), .B2(U3149), 
        .ZN(U3342) );
  INV_X1 U5144 ( .A(DATAI_9_), .ZN(n4769) );
  AOI22_X1 U5145 ( .A1(STATE_REG_SCAN_IN), .A2(n4596), .B1(n4769), .B2(U3149), 
        .ZN(U3343) );
  INV_X1 U5146 ( .A(DATAI_8_), .ZN(n4991) );
  AOI22_X1 U5147 ( .A1(STATE_REG_SCAN_IN), .A2(n2279), .B1(n4991), .B2(U3149), 
        .ZN(U3344) );
  AOI22_X1 U5148 ( .A1(STATE_REG_SCAN_IN), .A2(n4597), .B1(n2552), .B2(U3149), 
        .ZN(U3345) );
  INV_X1 U5149 ( .A(DATAI_6_), .ZN(n4904) );
  AOI22_X1 U5150 ( .A1(STATE_REG_SCAN_IN), .A2(n4598), .B1(n4904), .B2(U3149), 
        .ZN(U3346) );
  INV_X1 U5151 ( .A(DATAI_5_), .ZN(n4599) );
  AOI22_X1 U5152 ( .A1(STATE_REG_SCAN_IN), .A2(n4600), .B1(n4599), .B2(U3149), 
        .ZN(U3347) );
  OAI211_X1 U5153 ( .C1(n4603), .C2(n4624), .A(n4602), .B(n4601), .ZN(n4604)
         );
  INV_X1 U5154 ( .A(n4604), .ZN(n4632) );
  AOI22_X1 U5155 ( .A1(n4631), .A2(n4632), .B1(n2484), .B2(n4630), .ZN(U3467)
         );
  OAI22_X1 U5156 ( .A1(n4607), .A2(n4624), .B1(n4606), .B2(n4605), .ZN(n4608)
         );
  NOR2_X1 U5157 ( .A1(n4609), .A2(n4608), .ZN(n4634) );
  AOI22_X1 U5158 ( .A1(n4631), .A2(n4634), .B1(n2470), .B2(n4630), .ZN(U3469)
         );
  AOI21_X1 U5159 ( .B1(n4618), .B2(n4611), .A(n4610), .ZN(n4638) );
  OAI22_X1 U5160 ( .A1(n4371), .A2(n4635), .B1(n4631), .B2(n4612), .ZN(n4613)
         );
  INV_X1 U5161 ( .A(n4613), .ZN(n4614) );
  OAI21_X1 U5162 ( .B1(n4638), .B2(n4630), .A(n4614), .ZN(U3471) );
  INV_X1 U5163 ( .A(n4615), .ZN(n4617) );
  AOI211_X1 U5164 ( .C1(n4619), .C2(n4618), .A(n4617), .B(n4616), .ZN(n4640)
         );
  AOI22_X1 U5165 ( .A1(n4631), .A2(n4640), .B1(n2511), .B2(n4630), .ZN(U3475)
         );
  AOI211_X1 U5166 ( .C1(n4623), .C2(n4622), .A(n4621), .B(n4620), .ZN(n4642)
         );
  AOI22_X1 U5167 ( .A1(n4631), .A2(n4642), .B1(n2544), .B2(n4630), .ZN(U3481)
         );
  NOR2_X1 U5168 ( .A1(n4625), .A2(n4624), .ZN(n4627) );
  AOI211_X1 U5169 ( .C1(n4629), .C2(n4628), .A(n4627), .B(n4626), .ZN(n4645)
         );
  AOI22_X1 U5170 ( .A1(n4631), .A2(n4645), .B1(n2591), .B2(n4630), .ZN(U3489)
         );
  AOI22_X1 U5171 ( .A1(n4646), .A2(n4632), .B1(n2863), .B2(n4643), .ZN(U3518)
         );
  INV_X1 U5172 ( .A(REG1_REG_1__SCAN_IN), .ZN(n4633) );
  AOI22_X1 U5173 ( .A1(n4646), .A2(n4634), .B1(n4633), .B2(n4643), .ZN(U3519)
         );
  OAI22_X1 U5174 ( .A1(n4309), .A2(n4635), .B1(n4646), .B2(n3828), .ZN(n4636)
         );
  INV_X1 U5175 ( .A(n4636), .ZN(n4637) );
  OAI21_X1 U5176 ( .B1(n4638), .B2(n4643), .A(n4637), .ZN(U3520) );
  INV_X1 U5177 ( .A(REG1_REG_4__SCAN_IN), .ZN(n4639) );
  AOI22_X1 U5178 ( .A1(n4646), .A2(n4640), .B1(n4639), .B2(n4643), .ZN(U3522)
         );
  AOI22_X1 U5179 ( .A1(n4646), .A2(n4642), .B1(n4641), .B2(n4643), .ZN(U3525)
         );
  AOI22_X1 U5180 ( .A1(n4646), .A2(n4645), .B1(n4644), .B2(n4643), .ZN(U3529)
         );
  OAI22_X1 U5181 ( .A1(DATAI_25_), .A2(keyinput_g6), .B1(DATAI_8_), .B2(
        keyinput_g23), .ZN(n4647) );
  AOI221_X1 U5182 ( .B1(DATAI_25_), .B2(keyinput_g6), .C1(keyinput_g23), .C2(
        DATAI_8_), .A(n4647), .ZN(n4654) );
  OAI22_X1 U5183 ( .A1(D_REG_26__SCAN_IN), .A2(keyinput_g113), .B1(keyinput_g9), .B2(DATAI_22_), .ZN(n4648) );
  AOI221_X1 U5184 ( .B1(D_REG_26__SCAN_IN), .B2(keyinput_g113), .C1(DATAI_22_), 
        .C2(keyinput_g9), .A(n4648), .ZN(n4653) );
  OAI22_X1 U5185 ( .A1(IR_REG_1__SCAN_IN), .A2(keyinput_g56), .B1(
        keyinput_g102), .B2(D_REG_15__SCAN_IN), .ZN(n4649) );
  AOI221_X1 U5186 ( .B1(IR_REG_1__SCAN_IN), .B2(keyinput_g56), .C1(
        D_REG_15__SCAN_IN), .C2(keyinput_g102), .A(n4649), .ZN(n4652) );
  OAI22_X1 U5187 ( .A1(DATAI_19_), .A2(keyinput_g12), .B1(DATAI_14_), .B2(
        keyinput_g17), .ZN(n4650) );
  AOI221_X1 U5188 ( .B1(DATAI_19_), .B2(keyinput_g12), .C1(keyinput_g17), .C2(
        DATAI_14_), .A(n4650), .ZN(n4651) );
  NAND4_X1 U5189 ( .A1(n4654), .A2(n4653), .A3(n4652), .A4(n4651), .ZN(n4682)
         );
  OAI22_X1 U5190 ( .A1(REG3_REG_16__SCAN_IN), .A2(keyinput_g46), .B1(
        REG3_REG_10__SCAN_IN), .B2(keyinput_g37), .ZN(n4655) );
  AOI221_X1 U5191 ( .B1(REG3_REG_16__SCAN_IN), .B2(keyinput_g46), .C1(
        keyinput_g37), .C2(REG3_REG_10__SCAN_IN), .A(n4655), .ZN(n4662) );
  OAI22_X1 U5192 ( .A1(D_REG_18__SCAN_IN), .A2(keyinput_g105), .B1(
        REG3_REG_23__SCAN_IN), .B2(keyinput_g36), .ZN(n4656) );
  AOI221_X1 U5193 ( .B1(D_REG_18__SCAN_IN), .B2(keyinput_g105), .C1(
        keyinput_g36), .C2(REG3_REG_23__SCAN_IN), .A(n4656), .ZN(n4661) );
  OAI22_X1 U5194 ( .A1(D_REG_17__SCAN_IN), .A2(keyinput_g104), .B1(
        IR_REG_30__SCAN_IN), .B2(keyinput_g85), .ZN(n4657) );
  AOI221_X1 U5195 ( .B1(D_REG_17__SCAN_IN), .B2(keyinput_g104), .C1(
        keyinput_g85), .C2(IR_REG_30__SCAN_IN), .A(n4657), .ZN(n4660) );
  OAI22_X1 U5196 ( .A1(D_REG_11__SCAN_IN), .A2(keyinput_g98), .B1(DATAI_31_), 
        .B2(keyinput_g0), .ZN(n4658) );
  AOI221_X1 U5197 ( .B1(D_REG_11__SCAN_IN), .B2(keyinput_g98), .C1(keyinput_g0), .C2(DATAI_31_), .A(n4658), .ZN(n4659) );
  NAND4_X1 U5198 ( .A1(n4662), .A2(n4661), .A3(n4660), .A4(n4659), .ZN(n4681)
         );
  OAI22_X1 U5199 ( .A1(D_REG_1__SCAN_IN), .A2(keyinput_g88), .B1(keyinput_g107), .B2(D_REG_20__SCAN_IN), .ZN(n4663) );
  AOI221_X1 U5200 ( .B1(D_REG_1__SCAN_IN), .B2(keyinput_g88), .C1(
        D_REG_20__SCAN_IN), .C2(keyinput_g107), .A(n4663), .ZN(n4670) );
  OAI22_X1 U5201 ( .A1(D_REG_23__SCAN_IN), .A2(keyinput_g110), .B1(
        keyinput_g127), .B2(REG0_REG_8__SCAN_IN), .ZN(n4664) );
  AOI221_X1 U5202 ( .B1(D_REG_23__SCAN_IN), .B2(keyinput_g110), .C1(
        REG0_REG_8__SCAN_IN), .C2(keyinput_g127), .A(n4664), .ZN(n4669) );
  OAI22_X1 U5203 ( .A1(REG3_REG_9__SCAN_IN), .A2(keyinput_g51), .B1(DATAI_7_), 
        .B2(keyinput_g24), .ZN(n4665) );
  AOI221_X1 U5204 ( .B1(REG3_REG_9__SCAN_IN), .B2(keyinput_g51), .C1(
        keyinput_g24), .C2(DATAI_7_), .A(n4665), .ZN(n4668) );
  OAI22_X1 U5205 ( .A1(REG3_REG_27__SCAN_IN), .A2(keyinput_g34), .B1(
        REG3_REG_17__SCAN_IN), .B2(keyinput_g48), .ZN(n4666) );
  AOI221_X1 U5206 ( .B1(REG3_REG_27__SCAN_IN), .B2(keyinput_g34), .C1(
        keyinput_g48), .C2(REG3_REG_17__SCAN_IN), .A(n4666), .ZN(n4667) );
  NAND4_X1 U5207 ( .A1(n4670), .A2(n4669), .A3(n4668), .A4(n4667), .ZN(n4680)
         );
  OAI22_X1 U5208 ( .A1(D_REG_14__SCAN_IN), .A2(keyinput_g101), .B1(
        D_REG_6__SCAN_IN), .B2(keyinput_g93), .ZN(n4671) );
  AOI221_X1 U5209 ( .B1(D_REG_14__SCAN_IN), .B2(keyinput_g101), .C1(
        keyinput_g93), .C2(D_REG_6__SCAN_IN), .A(n4671), .ZN(n4678) );
  OAI22_X1 U5210 ( .A1(IR_REG_21__SCAN_IN), .A2(keyinput_g76), .B1(
        keyinput_g19), .B2(DATAI_12_), .ZN(n4672) );
  AOI221_X1 U5211 ( .B1(IR_REG_21__SCAN_IN), .B2(keyinput_g76), .C1(DATAI_12_), 
        .C2(keyinput_g19), .A(n4672), .ZN(n4677) );
  OAI22_X1 U5212 ( .A1(REG3_REG_25__SCAN_IN), .A2(keyinput_g45), .B1(DATAI_18_), .B2(keyinput_g13), .ZN(n4673) );
  AOI221_X1 U5213 ( .B1(REG3_REG_25__SCAN_IN), .B2(keyinput_g45), .C1(
        keyinput_g13), .C2(DATAI_18_), .A(n4673), .ZN(n4676) );
  OAI22_X1 U5214 ( .A1(n4846), .A2(keyinput_g27), .B1(keyinput_g32), .B2(
        STATE_REG_SCAN_IN), .ZN(n4674) );
  AOI221_X1 U5215 ( .B1(n4846), .B2(keyinput_g27), .C1(STATE_REG_SCAN_IN), 
        .C2(keyinput_g32), .A(n4674), .ZN(n4675) );
  NAND4_X1 U5216 ( .A1(n4678), .A2(n4677), .A3(n4676), .A4(n4675), .ZN(n4679)
         );
  NOR4_X1 U5217 ( .A1(n4682), .A2(n4681), .A3(n4680), .A4(n4679), .ZN(n5016)
         );
  OAI22_X1 U5218 ( .A1(D_REG_24__SCAN_IN), .A2(keyinput_g111), .B1(
        keyinput_g16), .B2(DATAI_15_), .ZN(n4683) );
  AOI221_X1 U5219 ( .B1(D_REG_24__SCAN_IN), .B2(keyinput_g111), .C1(DATAI_15_), 
        .C2(keyinput_g16), .A(n4683), .ZN(n4690) );
  OAI22_X1 U5220 ( .A1(D_REG_5__SCAN_IN), .A2(keyinput_g92), .B1(
        D_REG_2__SCAN_IN), .B2(keyinput_g89), .ZN(n4684) );
  AOI221_X1 U5221 ( .B1(D_REG_5__SCAN_IN), .B2(keyinput_g92), .C1(keyinput_g89), .C2(D_REG_2__SCAN_IN), .A(n4684), .ZN(n4689) );
  OAI22_X1 U5222 ( .A1(IR_REG_18__SCAN_IN), .A2(keyinput_g73), .B1(
        IR_REG_17__SCAN_IN), .B2(keyinput_g72), .ZN(n4685) );
  AOI221_X1 U5223 ( .B1(IR_REG_18__SCAN_IN), .B2(keyinput_g73), .C1(
        keyinput_g72), .C2(IR_REG_17__SCAN_IN), .A(n4685), .ZN(n4688) );
  OAI22_X1 U5224 ( .A1(IR_REG_14__SCAN_IN), .A2(keyinput_g69), .B1(DATAI_5_), 
        .B2(keyinput_g26), .ZN(n4686) );
  AOI221_X1 U5225 ( .B1(IR_REG_14__SCAN_IN), .B2(keyinput_g69), .C1(
        keyinput_g26), .C2(DATAI_5_), .A(n4686), .ZN(n4687) );
  NAND4_X1 U5226 ( .A1(n4690), .A2(n4689), .A3(n4688), .A4(n4687), .ZN(n4817)
         );
  OAI22_X1 U5227 ( .A1(DATAI_2_), .A2(keyinput_g29), .B1(DATAI_24_), .B2(
        keyinput_g7), .ZN(n4691) );
  AOI221_X1 U5228 ( .B1(DATAI_2_), .B2(keyinput_g29), .C1(keyinput_g7), .C2(
        DATAI_24_), .A(n4691), .ZN(n4716) );
  OAI22_X1 U5229 ( .A1(IR_REG_0__SCAN_IN), .A2(keyinput_g55), .B1(keyinput_g42), .B2(REG3_REG_1__SCAN_IN), .ZN(n4692) );
  AOI221_X1 U5230 ( .B1(IR_REG_0__SCAN_IN), .B2(keyinput_g55), .C1(
        REG3_REG_1__SCAN_IN), .C2(keyinput_g42), .A(n4692), .ZN(n4695) );
  OAI22_X1 U5231 ( .A1(DATAI_23_), .A2(keyinput_g8), .B1(keyinput_g52), .B2(
        REG3_REG_0__SCAN_IN), .ZN(n4693) );
  AOI221_X1 U5232 ( .B1(DATAI_23_), .B2(keyinput_g8), .C1(REG3_REG_0__SCAN_IN), 
        .C2(keyinput_g52), .A(n4693), .ZN(n4694) );
  OAI211_X1 U5233 ( .C1(n2660), .C2(keyinput_g14), .A(n4695), .B(n4694), .ZN(
        n4696) );
  AOI21_X1 U5234 ( .B1(n2660), .B2(keyinput_g14), .A(n4696), .ZN(n4715) );
  AOI22_X1 U5235 ( .A1(IR_REG_2__SCAN_IN), .A2(keyinput_g57), .B1(
        IR_REG_10__SCAN_IN), .B2(keyinput_g65), .ZN(n4697) );
  OAI221_X1 U5236 ( .B1(IR_REG_2__SCAN_IN), .B2(keyinput_g57), .C1(
        IR_REG_10__SCAN_IN), .C2(keyinput_g65), .A(n4697), .ZN(n4704) );
  AOI22_X1 U5237 ( .A1(IR_REG_5__SCAN_IN), .A2(keyinput_g60), .B1(
        IR_REG_6__SCAN_IN), .B2(keyinput_g61), .ZN(n4698) );
  OAI221_X1 U5238 ( .B1(IR_REG_5__SCAN_IN), .B2(keyinput_g60), .C1(
        IR_REG_6__SCAN_IN), .C2(keyinput_g61), .A(n4698), .ZN(n4703) );
  AOI22_X1 U5239 ( .A1(IR_REG_8__SCAN_IN), .A2(keyinput_g63), .B1(
        IR_REG_7__SCAN_IN), .B2(keyinput_g62), .ZN(n4699) );
  OAI221_X1 U5240 ( .B1(IR_REG_8__SCAN_IN), .B2(keyinput_g63), .C1(
        IR_REG_7__SCAN_IN), .C2(keyinput_g62), .A(n4699), .ZN(n4702) );
  AOI22_X1 U5241 ( .A1(DATAI_11_), .A2(keyinput_g20), .B1(IR_REG_9__SCAN_IN), 
        .B2(keyinput_g64), .ZN(n4700) );
  OAI221_X1 U5242 ( .B1(DATAI_11_), .B2(keyinput_g20), .C1(IR_REG_9__SCAN_IN), 
        .C2(keyinput_g64), .A(n4700), .ZN(n4701) );
  NOR4_X1 U5243 ( .A1(n4704), .A2(n4703), .A3(n4702), .A4(n4701), .ZN(n4714)
         );
  AOI22_X1 U5244 ( .A1(IR_REG_13__SCAN_IN), .A2(keyinput_g68), .B1(
        IR_REG_19__SCAN_IN), .B2(keyinput_g74), .ZN(n4705) );
  OAI221_X1 U5245 ( .B1(IR_REG_13__SCAN_IN), .B2(keyinput_g68), .C1(
        IR_REG_19__SCAN_IN), .C2(keyinput_g74), .A(n4705), .ZN(n4712) );
  AOI22_X1 U5246 ( .A1(D_REG_21__SCAN_IN), .A2(keyinput_g108), .B1(
        D_REG_25__SCAN_IN), .B2(keyinput_g112), .ZN(n4706) );
  OAI221_X1 U5247 ( .B1(D_REG_21__SCAN_IN), .B2(keyinput_g108), .C1(
        D_REG_25__SCAN_IN), .C2(keyinput_g112), .A(n4706), .ZN(n4711) );
  AOI22_X1 U5248 ( .A1(D_REG_27__SCAN_IN), .A2(keyinput_g114), .B1(
        D_REG_29__SCAN_IN), .B2(keyinput_g116), .ZN(n4707) );
  OAI221_X1 U5249 ( .B1(D_REG_27__SCAN_IN), .B2(keyinput_g114), .C1(
        D_REG_29__SCAN_IN), .C2(keyinput_g116), .A(n4707), .ZN(n4710) );
  AOI22_X1 U5250 ( .A1(DATAI_20_), .A2(keyinput_g11), .B1(DATAI_29_), .B2(
        keyinput_g2), .ZN(n4708) );
  OAI221_X1 U5251 ( .B1(DATAI_20_), .B2(keyinput_g11), .C1(DATAI_29_), .C2(
        keyinput_g2), .A(n4708), .ZN(n4709) );
  NOR4_X1 U5252 ( .A1(n4712), .A2(n4711), .A3(n4710), .A4(n4709), .ZN(n4713)
         );
  NAND4_X1 U5253 ( .A1(n4716), .A2(n4715), .A3(n4714), .A4(n4713), .ZN(n4816)
         );
  INV_X1 U5254 ( .A(DATAI_26_), .ZN(n4906) );
  AOI22_X1 U5255 ( .A1(n4907), .A2(keyinput_g91), .B1(keyinput_g5), .B2(n4906), 
        .ZN(n4717) );
  OAI221_X1 U5256 ( .B1(n4907), .B2(keyinput_g91), .C1(n4906), .C2(keyinput_g5), .A(n4717), .ZN(n4725) );
  AOI22_X1 U5257 ( .A1(n4894), .A2(keyinput_g18), .B1(n4896), .B2(keyinput_g71), .ZN(n4718) );
  OAI221_X1 U5258 ( .B1(n4894), .B2(keyinput_g18), .C1(n4896), .C2(
        keyinput_g71), .A(n4718), .ZN(n4724) );
  AOI22_X1 U5259 ( .A1(n4904), .A2(keyinput_g25), .B1(n4720), .B2(keyinput_g3), 
        .ZN(n4719) );
  OAI221_X1 U5260 ( .B1(n4904), .B2(keyinput_g25), .C1(n4720), .C2(keyinput_g3), .A(n4719), .ZN(n4723) );
  XNOR2_X1 U5261 ( .A(n4721), .B(keyinput_g77), .ZN(n4722) );
  NOR4_X1 U5262 ( .A1(n4725), .A2(n4724), .A3(n4723), .A4(n4722), .ZN(n4728)
         );
  XOR2_X1 U5263 ( .A(keyinput_g109), .B(n4726), .Z(n4727) );
  AND2_X1 U5264 ( .A1(n4728), .A2(n4727), .ZN(n4765) );
  AOI22_X1 U5265 ( .A1(n2446), .A2(keyinput_g84), .B1(keyinput_g122), .B2(
        n2503), .ZN(n4729) );
  OAI221_X1 U5266 ( .B1(n2446), .B2(keyinput_g84), .C1(n2503), .C2(
        keyinput_g122), .A(n4729), .ZN(n4740) );
  INV_X1 U5267 ( .A(REG3_REG_19__SCAN_IN), .ZN(n4731) );
  AOI22_X1 U5268 ( .A1(n4731), .A2(keyinput_g39), .B1(n4920), .B2(
        keyinput_g115), .ZN(n4730) );
  OAI221_X1 U5269 ( .B1(n4731), .B2(keyinput_g39), .C1(n4920), .C2(
        keyinput_g115), .A(n4730), .ZN(n4739) );
  AOI22_X1 U5270 ( .A1(n4734), .A2(keyinput_g100), .B1(n4733), .B2(
        keyinput_g118), .ZN(n4732) );
  OAI221_X1 U5271 ( .B1(n4734), .B2(keyinput_g100), .C1(n4733), .C2(
        keyinput_g118), .A(n4732), .ZN(n4738) );
  XOR2_X1 U5272 ( .A(n4919), .B(keyinput_g81), .Z(n4736) );
  XNOR2_X1 U5273 ( .A(REG3_REG_3__SCAN_IN), .B(keyinput_g38), .ZN(n4735) );
  NAND2_X1 U5274 ( .A1(n4736), .A2(n4735), .ZN(n4737) );
  NOR4_X1 U5275 ( .A1(n4740), .A2(n4739), .A3(n4738), .A4(n4737), .ZN(n4764)
         );
  AOI22_X1 U5276 ( .A1(n4941), .A2(keyinput_g96), .B1(keyinput_g43), .B2(n3516), .ZN(n4741) );
  OAI221_X1 U5277 ( .B1(n4941), .B2(keyinput_g96), .C1(n3516), .C2(
        keyinput_g43), .A(n4741), .ZN(n4750) );
  INV_X1 U5278 ( .A(DATAI_3_), .ZN(n4939) );
  AOI22_X1 U5279 ( .A1(n4925), .A2(keyinput_g97), .B1(keyinput_g28), .B2(n4939), .ZN(n4742) );
  OAI221_X1 U5280 ( .B1(n4925), .B2(keyinput_g97), .C1(n4939), .C2(
        keyinput_g28), .A(n4742), .ZN(n4749) );
  AOI22_X1 U5281 ( .A1(n4744), .A2(keyinput_g35), .B1(n4932), .B2(keyinput_g90), .ZN(n4743) );
  OAI221_X1 U5282 ( .B1(n4744), .B2(keyinput_g35), .C1(n4932), .C2(
        keyinput_g90), .A(n4743), .ZN(n4748) );
  XOR2_X1 U5283 ( .A(n4917), .B(keyinput_g10), .Z(n4746) );
  XNOR2_X1 U5284 ( .A(IR_REG_12__SCAN_IN), .B(keyinput_g67), .ZN(n4745) );
  NAND2_X1 U5285 ( .A1(n4746), .A2(n4745), .ZN(n4747) );
  NOR4_X1 U5286 ( .A1(n4750), .A2(n4749), .A3(n4748), .A4(n4747), .ZN(n4763)
         );
  AOI22_X1 U5287 ( .A1(n4752), .A2(keyinput_g95), .B1(keyinput_g40), .B2(n2728), .ZN(n4751) );
  OAI221_X1 U5288 ( .B1(n4752), .B2(keyinput_g95), .C1(n2728), .C2(
        keyinput_g40), .A(n4751), .ZN(n4761) );
  XNOR2_X1 U5289 ( .A(n4753), .B(keyinput_g103), .ZN(n4760) );
  INV_X1 U5290 ( .A(DATAI_30_), .ZN(n4934) );
  XNOR2_X1 U5291 ( .A(n4934), .B(keyinput_g1), .ZN(n4759) );
  INV_X1 U5292 ( .A(DATAI_0_), .ZN(n4950) );
  XOR2_X1 U5293 ( .A(n4950), .B(keyinput_g31), .Z(n4757) );
  XNOR2_X1 U5294 ( .A(IR_REG_25__SCAN_IN), .B(keyinput_g80), .ZN(n4756) );
  XNOR2_X1 U5295 ( .A(IR_REG_27__SCAN_IN), .B(keyinput_g82), .ZN(n4755) );
  XNOR2_X1 U5296 ( .A(IR_REG_23__SCAN_IN), .B(keyinput_g78), .ZN(n4754) );
  NAND4_X1 U5297 ( .A1(n4757), .A2(n4756), .A3(n4755), .A4(n4754), .ZN(n4758)
         );
  NOR4_X1 U5298 ( .A1(n4761), .A2(n4760), .A3(n4759), .A4(n4758), .ZN(n4762)
         );
  NAND4_X1 U5299 ( .A1(n4765), .A2(n4764), .A3(n4763), .A4(n4762), .ZN(n4815)
         );
  AOI22_X1 U5300 ( .A1(n2511), .A2(keyinput_g123), .B1(n4767), .B2(keyinput_g4), .ZN(n4766) );
  OAI221_X1 U5301 ( .B1(n2511), .B2(keyinput_g123), .C1(n4767), .C2(
        keyinput_g4), .A(n4766), .ZN(n4775) );
  AOI22_X1 U5302 ( .A1(n4955), .A2(keyinput_g44), .B1(keyinput_g22), .B2(n4769), .ZN(n4768) );
  OAI221_X1 U5303 ( .B1(n4955), .B2(keyinput_g44), .C1(n4769), .C2(
        keyinput_g22), .A(n4768), .ZN(n4774) );
  AOI22_X1 U5304 ( .A1(n4612), .A2(keyinput_g121), .B1(n2613), .B2(
        keyinput_g54), .ZN(n4770) );
  OAI221_X1 U5305 ( .B1(n4612), .B2(keyinput_g121), .C1(n2613), .C2(
        keyinput_g54), .A(n4770), .ZN(n4773) );
  AOI22_X1 U5306 ( .A1(n4958), .A2(keyinput_g41), .B1(n2646), .B2(keyinput_g70), .ZN(n4771) );
  OAI221_X1 U5307 ( .B1(n4958), .B2(keyinput_g41), .C1(n2646), .C2(
        keyinput_g70), .A(n4771), .ZN(n4772) );
  NOR4_X1 U5308 ( .A1(n4775), .A2(n4774), .A3(n4773), .A4(n4772), .ZN(n4813)
         );
  AOI22_X1 U5309 ( .A1(n2525), .A2(keyinput_g124), .B1(n4777), .B2(
        keyinput_g53), .ZN(n4776) );
  OAI221_X1 U5310 ( .B1(n2525), .B2(keyinput_g124), .C1(n4777), .C2(
        keyinput_g53), .A(n4776), .ZN(n4787) );
  AOI22_X1 U5311 ( .A1(n4779), .A2(keyinput_g106), .B1(keyinput_g21), .B2(
        n4967), .ZN(n4778) );
  OAI221_X1 U5312 ( .B1(n4779), .B2(keyinput_g106), .C1(n4967), .C2(
        keyinput_g21), .A(n4778), .ZN(n4786) );
  XOR2_X1 U5313 ( .A(n2484), .B(keyinput_g119), .Z(n4784) );
  XOR2_X1 U5314 ( .A(n4780), .B(keyinput_g47), .Z(n4783) );
  XNOR2_X1 U5315 ( .A(IR_REG_3__SCAN_IN), .B(keyinput_g58), .ZN(n4782) );
  XNOR2_X1 U5316 ( .A(IR_REG_24__SCAN_IN), .B(keyinput_g79), .ZN(n4781) );
  NAND4_X1 U5317 ( .A1(n4784), .A2(n4783), .A3(n4782), .A4(n4781), .ZN(n4785)
         );
  NOR3_X1 U5318 ( .A1(n4787), .A2(n4786), .A3(n4785), .ZN(n4812) );
  AOI22_X1 U5319 ( .A1(n4789), .A2(keyinput_g33), .B1(keyinput_g126), .B2(
        n2544), .ZN(n4788) );
  OAI221_X1 U5320 ( .B1(n4789), .B2(keyinput_g33), .C1(n2544), .C2(
        keyinput_g126), .A(n4788), .ZN(n4798) );
  INV_X1 U5321 ( .A(D_REG_0__SCAN_IN), .ZN(n4791) );
  AOI22_X1 U5322 ( .A1(n4791), .A2(keyinput_g87), .B1(keyinput_g49), .B2(n4977), .ZN(n4790) );
  OAI221_X1 U5323 ( .B1(n4791), .B2(keyinput_g87), .C1(n4977), .C2(
        keyinput_g49), .A(n4790), .ZN(n4797) );
  XNOR2_X1 U5324 ( .A(n4975), .B(keyinput_g99), .ZN(n4796) );
  XNOR2_X1 U5325 ( .A(IR_REG_31__SCAN_IN), .B(keyinput_g86), .ZN(n4794) );
  XNOR2_X1 U5326 ( .A(REG3_REG_4__SCAN_IN), .B(keyinput_g50), .ZN(n4793) );
  XNOR2_X1 U5327 ( .A(IR_REG_11__SCAN_IN), .B(keyinput_g66), .ZN(n4792) );
  NAND3_X1 U5328 ( .A1(n4794), .A2(n4793), .A3(n4792), .ZN(n4795) );
  NOR4_X1 U5329 ( .A1(n4798), .A2(n4797), .A3(n4796), .A4(n4795), .ZN(n4811)
         );
  AOI22_X1 U5330 ( .A1(n4989), .A2(keyinput_g15), .B1(keyinput_g120), .B2(
        n2470), .ZN(n4799) );
  OAI221_X1 U5331 ( .B1(n4989), .B2(keyinput_g15), .C1(n2470), .C2(
        keyinput_g120), .A(n4799), .ZN(n4805) );
  XNOR2_X1 U5332 ( .A(n4988), .B(keyinput_g117), .ZN(n4804) );
  XNOR2_X1 U5333 ( .A(n4800), .B(keyinput_g59), .ZN(n4803) );
  XNOR2_X1 U5334 ( .A(n4801), .B(keyinput_g83), .ZN(n4802) );
  OR4_X1 U5335 ( .A1(n4805), .A2(n4804), .A3(n4803), .A4(n4802), .ZN(n4809) );
  AOI22_X1 U5336 ( .A1(n2739), .A2(keyinput_g75), .B1(keyinput_g30), .B2(n2480), .ZN(n4806) );
  OAI221_X1 U5337 ( .B1(n2739), .B2(keyinput_g75), .C1(n2480), .C2(
        keyinput_g30), .A(n4806), .ZN(n4808) );
  XNOR2_X1 U5338 ( .A(n4992), .B(keyinput_g94), .ZN(n4807) );
  NOR3_X1 U5339 ( .A1(n4809), .A2(n4808), .A3(n4807), .ZN(n4810) );
  NAND4_X1 U5340 ( .A1(n4813), .A2(n4812), .A3(n4811), .A4(n4810), .ZN(n4814)
         );
  NOR4_X1 U5341 ( .A1(n4817), .A2(n4816), .A3(n4815), .A4(n4814), .ZN(n5015)
         );
  OAI22_X1 U5342 ( .A1(IR_REG_11__SCAN_IN), .A2(keyinput_f66), .B1(
        keyinput_f102), .B2(D_REG_15__SCAN_IN), .ZN(n4818) );
  AOI221_X1 U5343 ( .B1(IR_REG_11__SCAN_IN), .B2(keyinput_f66), .C1(
        D_REG_15__SCAN_IN), .C2(keyinput_f102), .A(n4818), .ZN(n4825) );
  OAI22_X1 U5344 ( .A1(D_REG_0__SCAN_IN), .A2(keyinput_f87), .B1(keyinput_f12), 
        .B2(DATAI_19_), .ZN(n4819) );
  AOI221_X1 U5345 ( .B1(D_REG_0__SCAN_IN), .B2(keyinput_f87), .C1(DATAI_19_), 
        .C2(keyinput_f12), .A(n4819), .ZN(n4824) );
  OAI22_X1 U5346 ( .A1(REG3_REG_16__SCAN_IN), .A2(keyinput_f46), .B1(
        keyinput_f33), .B2(REG3_REG_7__SCAN_IN), .ZN(n4820) );
  AOI221_X1 U5347 ( .B1(REG3_REG_16__SCAN_IN), .B2(keyinput_f46), .C1(
        REG3_REG_7__SCAN_IN), .C2(keyinput_f33), .A(n4820), .ZN(n4823) );
  OAI22_X1 U5348 ( .A1(REG3_REG_23__SCAN_IN), .A2(keyinput_f36), .B1(
        keyinput_f47), .B2(REG3_REG_5__SCAN_IN), .ZN(n4821) );
  AOI221_X1 U5349 ( .B1(REG3_REG_23__SCAN_IN), .B2(keyinput_f36), .C1(
        REG3_REG_5__SCAN_IN), .C2(keyinput_f47), .A(n4821), .ZN(n4822) );
  NAND4_X1 U5350 ( .A1(n4825), .A2(n4824), .A3(n4823), .A4(n4822), .ZN(n4854)
         );
  OAI22_X1 U5351 ( .A1(IR_REG_24__SCAN_IN), .A2(keyinput_f79), .B1(
        keyinput_f105), .B2(D_REG_18__SCAN_IN), .ZN(n4826) );
  AOI221_X1 U5352 ( .B1(IR_REG_24__SCAN_IN), .B2(keyinput_f79), .C1(
        D_REG_18__SCAN_IN), .C2(keyinput_f105), .A(n4826), .ZN(n4833) );
  OAI22_X1 U5353 ( .A1(IR_REG_3__SCAN_IN), .A2(keyinput_f58), .B1(
        keyinput_f104), .B2(D_REG_17__SCAN_IN), .ZN(n4827) );
  AOI221_X1 U5354 ( .B1(IR_REG_3__SCAN_IN), .B2(keyinput_f58), .C1(
        D_REG_17__SCAN_IN), .C2(keyinput_f104), .A(n4827), .ZN(n4832) );
  OAI22_X1 U5355 ( .A1(D_REG_20__SCAN_IN), .A2(keyinput_f107), .B1(
        D_REG_11__SCAN_IN), .B2(keyinput_f98), .ZN(n4828) );
  AOI221_X1 U5356 ( .B1(D_REG_20__SCAN_IN), .B2(keyinput_f107), .C1(
        keyinput_f98), .C2(D_REG_11__SCAN_IN), .A(n4828), .ZN(n4831) );
  OAI22_X1 U5357 ( .A1(D_REG_19__SCAN_IN), .A2(keyinput_f106), .B1(
        keyinput_f53), .B2(REG3_REG_20__SCAN_IN), .ZN(n4829) );
  AOI221_X1 U5358 ( .B1(D_REG_19__SCAN_IN), .B2(keyinput_f106), .C1(
        REG3_REG_20__SCAN_IN), .C2(keyinput_f53), .A(n4829), .ZN(n4830) );
  NAND4_X1 U5359 ( .A1(n4833), .A2(n4832), .A3(n4831), .A4(n4830), .ZN(n4853)
         );
  OAI22_X1 U5360 ( .A1(D_REG_1__SCAN_IN), .A2(keyinput_f88), .B1(keyinput_f51), 
        .B2(REG3_REG_9__SCAN_IN), .ZN(n4834) );
  AOI221_X1 U5361 ( .B1(D_REG_1__SCAN_IN), .B2(keyinput_f88), .C1(
        REG3_REG_9__SCAN_IN), .C2(keyinput_f51), .A(n4834), .ZN(n4841) );
  OAI22_X1 U5362 ( .A1(REG3_REG_13__SCAN_IN), .A2(keyinput_f54), .B1(
        REG0_REG_2__SCAN_IN), .B2(keyinput_f121), .ZN(n4835) );
  AOI221_X1 U5363 ( .B1(REG3_REG_13__SCAN_IN), .B2(keyinput_f54), .C1(
        keyinput_f121), .C2(REG0_REG_2__SCAN_IN), .A(n4835), .ZN(n4840) );
  OAI22_X1 U5364 ( .A1(D_REG_14__SCAN_IN), .A2(keyinput_f101), .B1(DATAI_9_), 
        .B2(keyinput_f22), .ZN(n4836) );
  AOI221_X1 U5365 ( .B1(D_REG_14__SCAN_IN), .B2(keyinput_f101), .C1(
        keyinput_f22), .C2(DATAI_9_), .A(n4836), .ZN(n4839) );
  OAI22_X1 U5366 ( .A1(D_REG_6__SCAN_IN), .A2(keyinput_f93), .B1(keyinput_f4), 
        .B2(DATAI_27_), .ZN(n4837) );
  AOI221_X1 U5367 ( .B1(D_REG_6__SCAN_IN), .B2(keyinput_f93), .C1(DATAI_27_), 
        .C2(keyinput_f4), .A(n4837), .ZN(n4838) );
  NAND4_X1 U5368 ( .A1(n4841), .A2(n4840), .A3(n4839), .A4(n4838), .ZN(n4852)
         );
  OAI22_X1 U5369 ( .A1(IR_REG_21__SCAN_IN), .A2(keyinput_f76), .B1(
        keyinput_f19), .B2(DATAI_12_), .ZN(n4842) );
  AOI221_X1 U5370 ( .B1(IR_REG_21__SCAN_IN), .B2(keyinput_f76), .C1(DATAI_12_), 
        .C2(keyinput_f19), .A(n4842), .ZN(n4850) );
  OAI22_X1 U5371 ( .A1(REG3_REG_25__SCAN_IN), .A2(keyinput_f45), .B1(
        REG0_REG_4__SCAN_IN), .B2(keyinput_f123), .ZN(n4843) );
  AOI221_X1 U5372 ( .B1(REG3_REG_25__SCAN_IN), .B2(keyinput_f45), .C1(
        keyinput_f123), .C2(REG0_REG_4__SCAN_IN), .A(n4843), .ZN(n4849) );
  OAI22_X1 U5373 ( .A1(STATE_REG_SCAN_IN), .A2(keyinput_f32), .B1(DATAI_18_), 
        .B2(keyinput_f13), .ZN(n4844) );
  AOI221_X1 U5374 ( .B1(STATE_REG_SCAN_IN), .B2(keyinput_f32), .C1(
        keyinput_f13), .C2(DATAI_18_), .A(n4844), .ZN(n4848) );
  OAI22_X1 U5375 ( .A1(n4846), .A2(keyinput_f27), .B1(keyinput_f95), .B2(
        D_REG_8__SCAN_IN), .ZN(n4845) );
  AOI221_X1 U5376 ( .B1(n4846), .B2(keyinput_f27), .C1(D_REG_8__SCAN_IN), .C2(
        keyinput_f95), .A(n4845), .ZN(n4847) );
  NAND4_X1 U5377 ( .A1(n4850), .A2(n4849), .A3(n4848), .A4(n4847), .ZN(n4851)
         );
  NOR4_X1 U5378 ( .A1(n4854), .A2(n4853), .A3(n4852), .A4(n4851), .ZN(n5009)
         );
  OAI22_X1 U5379 ( .A1(D_REG_24__SCAN_IN), .A2(keyinput_f111), .B1(
        D_REG_5__SCAN_IN), .B2(keyinput_f92), .ZN(n4855) );
  AOI221_X1 U5380 ( .B1(D_REG_24__SCAN_IN), .B2(keyinput_f111), .C1(
        keyinput_f92), .C2(D_REG_5__SCAN_IN), .A(n4855), .ZN(n4862) );
  OAI22_X1 U5381 ( .A1(IR_REG_31__SCAN_IN), .A2(keyinput_f86), .B1(
        keyinput_f89), .B2(D_REG_2__SCAN_IN), .ZN(n4856) );
  AOI221_X1 U5382 ( .B1(IR_REG_31__SCAN_IN), .B2(keyinput_f86), .C1(
        D_REG_2__SCAN_IN), .C2(keyinput_f89), .A(n4856), .ZN(n4861) );
  OAI22_X1 U5383 ( .A1(IR_REG_18__SCAN_IN), .A2(keyinput_f73), .B1(DATAI_5_), 
        .B2(keyinput_f26), .ZN(n4857) );
  AOI221_X1 U5384 ( .B1(IR_REG_18__SCAN_IN), .B2(keyinput_f73), .C1(
        keyinput_f26), .C2(DATAI_5_), .A(n4857), .ZN(n4860) );
  OAI22_X1 U5385 ( .A1(IR_REG_10__SCAN_IN), .A2(keyinput_f65), .B1(
        keyinput_f83), .B2(IR_REG_28__SCAN_IN), .ZN(n4858) );
  AOI221_X1 U5386 ( .B1(IR_REG_10__SCAN_IN), .B2(keyinput_f65), .C1(
        IR_REG_28__SCAN_IN), .C2(keyinput_f83), .A(n4858), .ZN(n4859) );
  NAND4_X1 U5387 ( .A1(n4862), .A2(n4861), .A3(n4860), .A4(n4859), .ZN(n5007)
         );
  OAI22_X1 U5388 ( .A1(DATAI_25_), .A2(keyinput_f6), .B1(keyinput_f29), .B2(
        DATAI_2_), .ZN(n4863) );
  AOI221_X1 U5389 ( .B1(DATAI_25_), .B2(keyinput_f6), .C1(DATAI_2_), .C2(
        keyinput_f29), .A(n4863), .ZN(n4888) );
  OAI22_X1 U5390 ( .A1(D_REG_26__SCAN_IN), .A2(keyinput_f113), .B1(
        keyinput_f35), .B2(REG3_REG_14__SCAN_IN), .ZN(n4864) );
  AOI221_X1 U5391 ( .B1(D_REG_26__SCAN_IN), .B2(keyinput_f113), .C1(
        REG3_REG_14__SCAN_IN), .C2(keyinput_f35), .A(n4864), .ZN(n4867) );
  OAI22_X1 U5392 ( .A1(DATAI_28_), .A2(keyinput_f3), .B1(REG3_REG_1__SCAN_IN), 
        .B2(keyinput_f42), .ZN(n4865) );
  AOI221_X1 U5393 ( .B1(DATAI_28_), .B2(keyinput_f3), .C1(keyinput_f42), .C2(
        REG3_REG_1__SCAN_IN), .A(n4865), .ZN(n4866) );
  OAI211_X1 U5394 ( .C1(n2660), .C2(keyinput_f14), .A(n4867), .B(n4866), .ZN(
        n4868) );
  AOI21_X1 U5395 ( .B1(n2660), .B2(keyinput_f14), .A(n4868), .ZN(n4887) );
  AOI22_X1 U5396 ( .A1(REG0_REG_1__SCAN_IN), .A2(keyinput_f120), .B1(
        IR_REG_7__SCAN_IN), .B2(keyinput_f62), .ZN(n4869) );
  OAI221_X1 U5397 ( .B1(REG0_REG_1__SCAN_IN), .B2(keyinput_f120), .C1(
        IR_REG_7__SCAN_IN), .C2(keyinput_f62), .A(n4869), .ZN(n4876) );
  AOI22_X1 U5398 ( .A1(IR_REG_8__SCAN_IN), .A2(keyinput_f63), .B1(
        IR_REG_12__SCAN_IN), .B2(keyinput_f67), .ZN(n4870) );
  OAI221_X1 U5399 ( .B1(IR_REG_8__SCAN_IN), .B2(keyinput_f63), .C1(
        IR_REG_12__SCAN_IN), .C2(keyinput_f67), .A(n4870), .ZN(n4875) );
  AOI22_X1 U5400 ( .A1(IR_REG_20__SCAN_IN), .A2(keyinput_f75), .B1(
        IR_REG_19__SCAN_IN), .B2(keyinput_f74), .ZN(n4871) );
  OAI221_X1 U5401 ( .B1(IR_REG_20__SCAN_IN), .B2(keyinput_f75), .C1(
        IR_REG_19__SCAN_IN), .C2(keyinput_f74), .A(n4871), .ZN(n4874) );
  AOI22_X1 U5402 ( .A1(D_REG_22__SCAN_IN), .A2(keyinput_f109), .B1(
        IR_REG_22__SCAN_IN), .B2(keyinput_f77), .ZN(n4872) );
  OAI221_X1 U5403 ( .B1(D_REG_22__SCAN_IN), .B2(keyinput_f109), .C1(
        IR_REG_22__SCAN_IN), .C2(keyinput_f77), .A(n4872), .ZN(n4873) );
  NOR4_X1 U5404 ( .A1(n4876), .A2(n4875), .A3(n4874), .A4(n4873), .ZN(n4886)
         );
  AOI22_X1 U5405 ( .A1(D_REG_31__SCAN_IN), .A2(keyinput_f118), .B1(
        D_REG_16__SCAN_IN), .B2(keyinput_f103), .ZN(n4877) );
  OAI221_X1 U5406 ( .B1(D_REG_31__SCAN_IN), .B2(keyinput_f118), .C1(
        D_REG_16__SCAN_IN), .C2(keyinput_f103), .A(n4877), .ZN(n4884) );
  AOI22_X1 U5407 ( .A1(IR_REG_29__SCAN_IN), .A2(keyinput_f84), .B1(
        D_REG_13__SCAN_IN), .B2(keyinput_f100), .ZN(n4878) );
  OAI221_X1 U5408 ( .B1(IR_REG_29__SCAN_IN), .B2(keyinput_f84), .C1(
        D_REG_13__SCAN_IN), .C2(keyinput_f100), .A(n4878), .ZN(n4883) );
  AOI22_X1 U5409 ( .A1(IR_REG_27__SCAN_IN), .A2(keyinput_f82), .B1(
        IR_REG_23__SCAN_IN), .B2(keyinput_f78), .ZN(n4879) );
  OAI221_X1 U5410 ( .B1(IR_REG_27__SCAN_IN), .B2(keyinput_f82), .C1(
        IR_REG_23__SCAN_IN), .C2(keyinput_f78), .A(n4879), .ZN(n4882) );
  AOI22_X1 U5411 ( .A1(REG3_REG_19__SCAN_IN), .A2(keyinput_f39), .B1(
        IR_REG_25__SCAN_IN), .B2(keyinput_f80), .ZN(n4880) );
  OAI221_X1 U5412 ( .B1(REG3_REG_19__SCAN_IN), .B2(keyinput_f39), .C1(
        IR_REG_25__SCAN_IN), .C2(keyinput_f80), .A(n4880), .ZN(n4881) );
  NOR4_X1 U5413 ( .A1(n4884), .A2(n4883), .A3(n4882), .A4(n4881), .ZN(n4885)
         );
  NAND4_X1 U5414 ( .A1(n4888), .A2(n4887), .A3(n4886), .A4(n4885), .ZN(n5006)
         );
  INV_X1 U5415 ( .A(DATAI_20_), .ZN(n4891) );
  AOI22_X1 U5416 ( .A1(n4891), .A2(keyinput_f11), .B1(n4890), .B2(
        keyinput_f116), .ZN(n4889) );
  OAI221_X1 U5417 ( .B1(n4891), .B2(keyinput_f11), .C1(n4890), .C2(
        keyinput_f116), .A(n4889), .ZN(n4902) );
  AOI22_X1 U5418 ( .A1(n4894), .A2(keyinput_f18), .B1(n4893), .B2(keyinput_f8), 
        .ZN(n4892) );
  OAI221_X1 U5419 ( .B1(n4894), .B2(keyinput_f18), .C1(n4893), .C2(keyinput_f8), .A(n4892), .ZN(n4901) );
  AOI22_X1 U5420 ( .A1(n4896), .A2(keyinput_f71), .B1(keyinput_f52), .B2(n2880), .ZN(n4895) );
  OAI221_X1 U5421 ( .B1(n4896), .B2(keyinput_f71), .C1(n2880), .C2(
        keyinput_f52), .A(n4895), .ZN(n4900) );
  AOI22_X1 U5422 ( .A1(n4898), .A2(keyinput_f112), .B1(n2421), .B2(
        keyinput_f72), .ZN(n4897) );
  OAI221_X1 U5423 ( .B1(n4898), .B2(keyinput_f112), .C1(n2421), .C2(
        keyinput_f72), .A(n4897), .ZN(n4899) );
  NOR4_X1 U5424 ( .A1(n4902), .A2(n4901), .A3(n4900), .A4(n4899), .ZN(n4948)
         );
  AOI22_X1 U5425 ( .A1(n4904), .A2(keyinput_f25), .B1(keyinput_f20), .B2(n2600), .ZN(n4903) );
  OAI221_X1 U5426 ( .B1(n4904), .B2(keyinput_f25), .C1(n2600), .C2(
        keyinput_f20), .A(n4903), .ZN(n4915) );
  AOI22_X1 U5427 ( .A1(n4907), .A2(keyinput_f91), .B1(keyinput_f5), .B2(n4906), 
        .ZN(n4905) );
  OAI221_X1 U5428 ( .B1(n4907), .B2(keyinput_f91), .C1(n4906), .C2(keyinput_f5), .A(n4905), .ZN(n4914) );
  AOI22_X1 U5429 ( .A1(n4910), .A2(keyinput_f114), .B1(keyinput_f16), .B2(
        n4909), .ZN(n4908) );
  OAI221_X1 U5430 ( .B1(n4910), .B2(keyinput_f114), .C1(n4909), .C2(
        keyinput_f16), .A(n4908), .ZN(n4913) );
  AOI22_X1 U5431 ( .A1(n2424), .A2(keyinput_f69), .B1(keyinput_f122), .B2(
        n2503), .ZN(n4911) );
  OAI221_X1 U5432 ( .B1(n2424), .B2(keyinput_f69), .C1(n2503), .C2(
        keyinput_f122), .A(n4911), .ZN(n4912) );
  NOR4_X1 U5433 ( .A1(n4915), .A2(n4914), .A3(n4913), .A4(n4912), .ZN(n4947)
         );
  AOI22_X1 U5434 ( .A1(n2395), .A2(keyinput_f55), .B1(keyinput_f10), .B2(n4917), .ZN(n4916) );
  OAI221_X1 U5435 ( .B1(n2395), .B2(keyinput_f55), .C1(n4917), .C2(
        keyinput_f10), .A(n4916), .ZN(n4929) );
  AOI22_X1 U5436 ( .A1(n4920), .A2(keyinput_f115), .B1(n4919), .B2(
        keyinput_f81), .ZN(n4918) );
  OAI221_X1 U5437 ( .B1(n4920), .B2(keyinput_f115), .C1(n4919), .C2(
        keyinput_f81), .A(n4918), .ZN(n4928) );
  XOR2_X1 U5438 ( .A(n4921), .B(keyinput_f2), .Z(n4924) );
  XNOR2_X1 U5439 ( .A(REG3_REG_3__SCAN_IN), .B(keyinput_f38), .ZN(n4923) );
  XNOR2_X1 U5440 ( .A(IR_REG_5__SCAN_IN), .B(keyinput_f60), .ZN(n4922) );
  NAND3_X1 U5441 ( .A1(n4924), .A2(n4923), .A3(n4922), .ZN(n4927) );
  XNOR2_X1 U5442 ( .A(n4925), .B(keyinput_f97), .ZN(n4926) );
  NOR4_X1 U5443 ( .A1(n4929), .A2(n4928), .A3(n4927), .A4(n4926), .ZN(n4946)
         );
  INV_X1 U5444 ( .A(DATAI_24_), .ZN(n4931) );
  AOI22_X1 U5445 ( .A1(n4932), .A2(keyinput_f90), .B1(keyinput_f7), .B2(n4931), 
        .ZN(n4930) );
  OAI221_X1 U5446 ( .B1(n4932), .B2(keyinput_f90), .C1(n4931), .C2(keyinput_f7), .A(n4930), .ZN(n4937) );
  XNOR2_X1 U5447 ( .A(n4933), .B(keyinput_f64), .ZN(n4936) );
  XNOR2_X1 U5448 ( .A(n4934), .B(keyinput_f1), .ZN(n4935) );
  OR3_X1 U5449 ( .A1(n4937), .A2(n4936), .A3(n4935), .ZN(n4944) );
  AOI22_X1 U5450 ( .A1(n4939), .A2(keyinput_f28), .B1(n3516), .B2(keyinput_f43), .ZN(n4938) );
  OAI221_X1 U5451 ( .B1(n4939), .B2(keyinput_f28), .C1(n3516), .C2(
        keyinput_f43), .A(n4938), .ZN(n4943) );
  AOI22_X1 U5452 ( .A1(n4941), .A2(keyinput_f96), .B1(n2498), .B2(keyinput_f57), .ZN(n4940) );
  OAI221_X1 U5453 ( .B1(n4941), .B2(keyinput_f96), .C1(n2498), .C2(
        keyinput_f57), .A(n4940), .ZN(n4942) );
  NOR3_X1 U5454 ( .A1(n4944), .A2(n4943), .A3(n4942), .ZN(n4945) );
  NAND4_X1 U5455 ( .A1(n4948), .A2(n4947), .A3(n4946), .A4(n4945), .ZN(n5005)
         );
  AOI22_X1 U5456 ( .A1(n4951), .A2(keyinput_f108), .B1(keyinput_f31), .B2(
        n4950), .ZN(n4949) );
  OAI221_X1 U5457 ( .B1(n4951), .B2(keyinput_f108), .C1(n4950), .C2(
        keyinput_f31), .A(n4949), .ZN(n4962) );
  AOI22_X1 U5458 ( .A1(n2574), .A2(keyinput_f61), .B1(keyinput_f40), .B2(n2728), .ZN(n4952) );
  OAI221_X1 U5459 ( .B1(n2574), .B2(keyinput_f61), .C1(n2728), .C2(
        keyinput_f40), .A(n4952), .ZN(n4961) );
  AOI22_X1 U5460 ( .A1(n4955), .A2(keyinput_f44), .B1(n4954), .B2(keyinput_f48), .ZN(n4953) );
  OAI221_X1 U5461 ( .B1(n4955), .B2(keyinput_f44), .C1(n4954), .C2(
        keyinput_f48), .A(n4953), .ZN(n4960) );
  AOI22_X1 U5462 ( .A1(n4958), .A2(keyinput_f41), .B1(n4957), .B2(keyinput_f34), .ZN(n4956) );
  OAI221_X1 U5463 ( .B1(n4958), .B2(keyinput_f41), .C1(n4957), .C2(
        keyinput_f34), .A(n4956), .ZN(n4959) );
  NOR4_X1 U5464 ( .A1(n4962), .A2(n4961), .A3(n4960), .A4(n4959), .ZN(n5003)
         );
  AOI22_X1 U5465 ( .A1(n2552), .A2(keyinput_f24), .B1(n2525), .B2(
        keyinput_f124), .ZN(n4963) );
  OAI221_X1 U5466 ( .B1(n2552), .B2(keyinput_f24), .C1(n2525), .C2(
        keyinput_f124), .A(n4963), .ZN(n4973) );
  AOI22_X1 U5467 ( .A1(n4965), .A2(keyinput_f110), .B1(n2646), .B2(
        keyinput_f70), .ZN(n4964) );
  OAI221_X1 U5468 ( .B1(n4965), .B2(keyinput_f110), .C1(n2646), .C2(
        keyinput_f70), .A(n4964), .ZN(n4972) );
  AOI22_X1 U5469 ( .A1(n2556), .A2(keyinput_f127), .B1(n4967), .B2(
        keyinput_f21), .ZN(n4966) );
  OAI221_X1 U5470 ( .B1(n2556), .B2(keyinput_f127), .C1(n4967), .C2(
        keyinput_f21), .A(n4966), .ZN(n4971) );
  AOI22_X1 U5471 ( .A1(n4969), .A2(keyinput_f0), .B1(n2836), .B2(keyinput_f85), 
        .ZN(n4968) );
  OAI221_X1 U5472 ( .B1(n4969), .B2(keyinput_f0), .C1(n2836), .C2(keyinput_f85), .A(n4968), .ZN(n4970) );
  NOR4_X1 U5473 ( .A1(n4973), .A2(n4972), .A3(n4971), .A4(n4970), .ZN(n5002)
         );
  AOI22_X1 U5474 ( .A1(n2484), .A2(keyinput_f119), .B1(n4975), .B2(
        keyinput_f99), .ZN(n4974) );
  OAI221_X1 U5475 ( .B1(n2484), .B2(keyinput_f119), .C1(n4975), .C2(
        keyinput_f99), .A(n4974), .ZN(n4986) );
  AOI22_X1 U5476 ( .A1(n2544), .A2(keyinput_f126), .B1(n4977), .B2(
        keyinput_f49), .ZN(n4976) );
  OAI221_X1 U5477 ( .B1(n2544), .B2(keyinput_f126), .C1(n4977), .C2(
        keyinput_f49), .A(n4976), .ZN(n4985) );
  INV_X1 U5478 ( .A(DATAI_22_), .ZN(n4979) );
  AOI22_X1 U5479 ( .A1(n4980), .A2(keyinput_f17), .B1(n4979), .B2(keyinput_f9), 
        .ZN(n4978) );
  OAI221_X1 U5480 ( .B1(n4980), .B2(keyinput_f17), .C1(n4979), .C2(keyinput_f9), .A(n4978), .ZN(n4984) );
  XNOR2_X1 U5481 ( .A(REG3_REG_4__SCAN_IN), .B(keyinput_f50), .ZN(n4982) );
  XNOR2_X1 U5482 ( .A(REG3_REG_10__SCAN_IN), .B(keyinput_f37), .ZN(n4981) );
  NAND2_X1 U5483 ( .A1(n4982), .A2(n4981), .ZN(n4983) );
  NOR4_X1 U5484 ( .A1(n4986), .A2(n4985), .A3(n4984), .A4(n4983), .ZN(n5001)
         );
  AOI22_X1 U5485 ( .A1(n4989), .A2(keyinput_f15), .B1(n4988), .B2(
        keyinput_f117), .ZN(n4987) );
  OAI221_X1 U5486 ( .B1(n4989), .B2(keyinput_f15), .C1(n4988), .C2(
        keyinput_f117), .A(n4987), .ZN(n4999) );
  AOI22_X1 U5487 ( .A1(n2394), .A2(keyinput_f56), .B1(keyinput_f23), .B2(n4991), .ZN(n4990) );
  OAI221_X1 U5488 ( .B1(n2394), .B2(keyinput_f56), .C1(n4991), .C2(
        keyinput_f23), .A(n4990), .ZN(n4998) );
  XNOR2_X1 U5489 ( .A(n4992), .B(keyinput_f94), .ZN(n4997) );
  XNOR2_X1 U5490 ( .A(IR_REG_4__SCAN_IN), .B(keyinput_f59), .ZN(n4995) );
  XNOR2_X1 U5491 ( .A(IR_REG_13__SCAN_IN), .B(keyinput_f68), .ZN(n4994) );
  XNOR2_X1 U5492 ( .A(keyinput_f30), .B(DATAI_1_), .ZN(n4993) );
  NAND3_X1 U5493 ( .A1(n4995), .A2(n4994), .A3(n4993), .ZN(n4996) );
  NOR4_X1 U5494 ( .A1(n4999), .A2(n4998), .A3(n4997), .A4(n4996), .ZN(n5000)
         );
  NAND4_X1 U5495 ( .A1(n5003), .A2(n5002), .A3(n5001), .A4(n5000), .ZN(n5004)
         );
  NOR4_X1 U5496 ( .A1(n5007), .A2(n5006), .A3(n5005), .A4(n5004), .ZN(n5008)
         );
  NAND2_X1 U5497 ( .A1(n5009), .A2(n5008), .ZN(n5011) );
  AOI21_X1 U5498 ( .B1(keyinput_f125), .B2(n5011), .A(keyinput_g125), .ZN(
        n5013) );
  INV_X1 U5499 ( .A(keyinput_f125), .ZN(n5010) );
  AOI21_X1 U5500 ( .B1(n5011), .B2(n5010), .A(REG0_REG_6__SCAN_IN), .ZN(n5012)
         );
  AOI22_X1 U5501 ( .A1(REG0_REG_6__SCAN_IN), .A2(n5013), .B1(keyinput_g125), 
        .B2(n5012), .ZN(n5014) );
  AOI21_X1 U5502 ( .B1(n5016), .B2(n5015), .A(n5014), .ZN(n5018) );
  AOI22_X1 U5503 ( .A1(STATE_REG_SCAN_IN), .A2(IR_REG_0__SCAN_IN), .B1(
        DATAI_0_), .B2(U3149), .ZN(n5017) );
  XNOR2_X1 U5504 ( .A(n5018), .B(n5017), .ZN(U3352) );
  CLKBUF_X1 U2463 ( .A(n3282), .Z(n3042) );
  CLKBUF_X1 U2465 ( .A(n2943), .Z(n3448) );
  CLKBUF_X1 U2466 ( .A(n2485), .Z(n2219) );
  CLKBUF_X1 U2874 ( .A(n2492), .Z(n3632) );
endmodule

