

module b21_C_SARLock_k_64_8 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3, 
        keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, 
        keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, 
        keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, 
        keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, 
        keyinput28, keyinput29, keyinput30, keyinput31, keyinput32, keyinput33, 
        keyinput34, keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, 
        keyinput40, keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, 
        keyinput46, keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, 
        keyinput52, keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, 
        keyinput58, keyinput59, keyinput60, keyinput61, keyinput62, keyinput63, 
        ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58, 
        ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63, 
        ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51, 
        ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46, 
        U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, 
        P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, 
        P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, 
        P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, 
        P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440, P1_U3441, 
        P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, 
        P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, 
        P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, 
        P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, 
        P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463, P1_U3466, 
        P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484, P1_U3487, 
        P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505, P1_U3508, 
        P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, 
        P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, 
        P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, 
        P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, 
        P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, 
        P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, 
        P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289, P1_U3288, 
        P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, 
        P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, 
        P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, 
        P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262, P1_U3261, 
        P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, 
        P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, 
        P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241, P1_U3555, 
        P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, 
        P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, 
        P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, 
        P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, 
        P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238, P1_U3237, 
        P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, 
        P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, 
        P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, 
        P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084, P1_U3083, 
        P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354, P2_U3353, 
        P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347, P2_U3346, 
        P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340, P2_U3339, 
        P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333, P2_U3332, 
        P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437, P2_U3438, 
        P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321, P2_U3320, 
        P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314, P2_U3313, 
        P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307, P2_U3306, 
        P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300, P2_U3299, 
        P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, 
        P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, 
        P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502, P2_U3505, 
        P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, 
        P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, 
        P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, 
        P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533, P2_U3534, 
        P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540, P2_U3541, 
        P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547, P2_U3548, 
        P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294, P2_U3293, 
        P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, 
        P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, 
        P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, 
        P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, 
        P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, 
        P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, 
        P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3552, 
        P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, 
        P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565, P2_U3566, 
        P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572, P2_U3573, 
        P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579, P2_U3580, 
        P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152, P2_U3151, 
        P2_U3966 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4262, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4272, n4273,
         n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283,
         n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293,
         n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303,
         n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313,
         n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323,
         n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333,
         n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343,
         n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353,
         n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363,
         n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373,
         n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383,
         n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393,
         n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403,
         n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413,
         n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423,
         n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433,
         n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443,
         n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453,
         n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463,
         n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473,
         n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483,
         n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493,
         n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503,
         n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513,
         n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523,
         n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533,
         n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543,
         n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553,
         n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563,
         n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573,
         n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583,
         n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593,
         n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603,
         n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613,
         n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623,
         n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633,
         n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643,
         n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653,
         n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663,
         n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673,
         n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683,
         n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693,
         n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703,
         n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713,
         n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723,
         n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733,
         n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743,
         n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753,
         n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763,
         n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773,
         n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783,
         n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793,
         n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803,
         n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813,
         n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823,
         n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833,
         n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843,
         n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853,
         n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863,
         n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873,
         n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883,
         n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893,
         n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903,
         n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913,
         n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923,
         n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933,
         n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943,
         n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953,
         n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963,
         n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973,
         n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983,
         n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993,
         n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003,
         n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013,
         n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023,
         n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033,
         n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043,
         n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053,
         n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063,
         n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073,
         n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083,
         n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093,
         n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103,
         n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113,
         n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123,
         n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133,
         n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143,
         n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153,
         n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163,
         n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173,
         n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183,
         n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193,
         n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203,
         n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213,
         n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223,
         n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233,
         n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243,
         n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253,
         n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263,
         n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273,
         n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283,
         n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293,
         n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303,
         n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313,
         n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323,
         n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333,
         n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343,
         n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353,
         n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363,
         n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373,
         n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383,
         n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393,
         n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403,
         n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413,
         n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423,
         n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433,
         n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443,
         n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453,
         n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463,
         n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473,
         n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483,
         n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493,
         n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503,
         n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513,
         n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523,
         n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533,
         n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543,
         n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553,
         n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563,
         n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573,
         n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583,
         n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593,
         n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603,
         n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613,
         n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623,
         n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633,
         n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643,
         n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653,
         n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663,
         n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673,
         n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683,
         n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693,
         n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703,
         n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713,
         n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723,
         n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733,
         n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743,
         n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753,
         n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763,
         n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773,
         n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783,
         n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793,
         n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803,
         n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813,
         n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823,
         n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833,
         n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843,
         n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853,
         n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863,
         n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873,
         n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883,
         n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893,
         n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903,
         n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913,
         n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923,
         n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933,
         n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943,
         n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953,
         n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963,
         n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973,
         n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983,
         n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993,
         n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003,
         n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013,
         n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023,
         n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033,
         n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043,
         n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053,
         n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063,
         n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073,
         n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083,
         n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093,
         n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103,
         n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113,
         n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123,
         n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133,
         n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143,
         n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153,
         n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163,
         n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173,
         n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183,
         n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193,
         n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203,
         n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213,
         n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223,
         n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233,
         n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243,
         n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253,
         n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263,
         n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273,
         n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283,
         n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293,
         n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303,
         n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313,
         n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323,
         n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333,
         n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343,
         n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353,
         n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363,
         n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373,
         n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383,
         n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393,
         n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403,
         n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413,
         n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423,
         n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433,
         n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443,
         n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453,
         n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463,
         n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473,
         n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483,
         n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493,
         n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503,
         n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513,
         n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523,
         n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533,
         n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543,
         n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553,
         n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563,
         n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573,
         n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583,
         n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593,
         n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603,
         n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613,
         n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623,
         n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633,
         n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643,
         n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653,
         n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663,
         n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673,
         n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683,
         n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693,
         n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703,
         n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713,
         n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723,
         n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733,
         n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743,
         n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753,
         n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763,
         n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773,
         n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783,
         n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793,
         n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803,
         n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813,
         n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823,
         n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833,
         n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843,
         n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853,
         n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863,
         n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873,
         n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883,
         n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893,
         n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903,
         n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913,
         n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923,
         n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933,
         n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943,
         n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953,
         n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963,
         n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973,
         n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983,
         n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993,
         n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003,
         n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013,
         n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023,
         n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033,
         n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043,
         n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053,
         n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063,
         n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073,
         n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083,
         n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093,
         n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103,
         n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113,
         n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123,
         n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133,
         n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143,
         n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153,
         n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163,
         n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173,
         n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183,
         n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193,
         n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203,
         n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213,
         n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223,
         n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233,
         n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243,
         n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253,
         n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263,
         n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273,
         n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283,
         n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293,
         n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303,
         n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313,
         n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323,
         n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333,
         n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343,
         n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353,
         n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363,
         n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373,
         n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383,
         n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393,
         n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403,
         n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413,
         n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423,
         n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433,
         n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443,
         n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453,
         n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463,
         n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473,
         n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483,
         n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493,
         n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503,
         n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513,
         n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523,
         n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533,
         n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543,
         n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553,
         n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563,
         n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573,
         n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583,
         n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593,
         n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603,
         n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613,
         n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623,
         n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633,
         n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643,
         n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653,
         n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663,
         n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673,
         n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683,
         n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693,
         n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703,
         n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713,
         n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723,
         n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733,
         n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743,
         n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753,
         n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763,
         n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773,
         n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783,
         n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793,
         n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803,
         n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813,
         n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823,
         n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833,
         n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843,
         n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853,
         n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863,
         n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873,
         n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883,
         n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893,
         n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903,
         n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913,
         n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923,
         n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933,
         n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943,
         n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953,
         n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963,
         n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973,
         n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983,
         n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993,
         n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003,
         n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013,
         n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023,
         n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033,
         n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043,
         n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053,
         n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063,
         n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073,
         n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083,
         n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093,
         n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103,
         n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113,
         n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123,
         n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133,
         n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143,
         n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153,
         n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163,
         n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173,
         n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183,
         n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193,
         n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203,
         n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213,
         n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223,
         n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233,
         n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243,
         n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253,
         n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263,
         n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273,
         n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283,
         n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293,
         n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303,
         n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313,
         n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323,
         n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333,
         n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343,
         n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353,
         n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363,
         n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373,
         n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383,
         n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393,
         n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403,
         n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413,
         n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423,
         n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433,
         n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443,
         n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453,
         n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463,
         n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473,
         n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483,
         n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493,
         n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503,
         n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513,
         n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523,
         n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533,
         n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543,
         n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553,
         n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563,
         n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573,
         n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583,
         n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593,
         n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603,
         n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613,
         n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623,
         n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633,
         n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643,
         n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653,
         n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663,
         n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673,
         n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683,
         n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693,
         n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703,
         n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713,
         n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723,
         n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733,
         n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743,
         n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753,
         n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763,
         n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773,
         n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783,
         n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793,
         n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803,
         n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813,
         n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823,
         n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833,
         n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843,
         n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853,
         n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863,
         n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873,
         n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883,
         n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893,
         n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903,
         n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913,
         n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923,
         n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933,
         n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943,
         n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953,
         n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963,
         n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973,
         n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983,
         n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993,
         n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003,
         n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013,
         n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023,
         n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033,
         n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043,
         n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053,
         n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063,
         n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073,
         n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083,
         n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093,
         n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103,
         n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113,
         n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123,
         n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133,
         n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143,
         n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153,
         n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163,
         n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173,
         n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183,
         n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193,
         n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203,
         n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213,
         n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223,
         n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233,
         n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243,
         n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253,
         n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263,
         n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273,
         n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283,
         n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293,
         n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303,
         n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313,
         n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323,
         n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333,
         n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343,
         n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353,
         n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363,
         n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373,
         n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383,
         n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393,
         n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403,
         n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413,
         n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423,
         n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433,
         n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443,
         n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453,
         n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463,
         n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473,
         n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483,
         n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493,
         n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503,
         n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513,
         n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523,
         n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533,
         n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543,
         n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553,
         n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563,
         n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573,
         n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583,
         n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593,
         n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603,
         n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613,
         n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623,
         n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633,
         n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643,
         n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653,
         n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663,
         n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673,
         n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683,
         n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693,
         n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703,
         n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713,
         n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723,
         n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733,
         n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743,
         n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753,
         n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763,
         n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773,
         n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783,
         n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793,
         n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803,
         n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813,
         n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823,
         n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833,
         n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843,
         n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853,
         n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863,
         n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873,
         n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883,
         n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893,
         n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903,
         n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913,
         n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923,
         n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933,
         n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943,
         n9944, n9945, n9946, n9947, n9949;

  OAI21_X1 U4768 ( .B1(n5699), .B2(n4595), .A(n4594), .ZN(n4599) );
  CLKBUF_X1 U4769 ( .A(n6309), .Z(n9949) );
  NAND2_X1 U4770 ( .A1(n7073), .A2(n7072), .ZN(n7166) );
  BUF_X2 U4771 ( .A(n5820), .Z(n6210) );
  NAND2_X1 U4772 ( .A1(n8687), .A2(n8688), .ZN(n6882) );
  INV_X1 U4773 ( .A(n8477), .ZN(n9596) );
  BUF_X1 U4774 ( .A(n4865), .Z(n4272) );
  CLKBUF_X2 U4775 ( .A(n4991), .Z(n5640) );
  CLKBUF_X2 U4777 ( .A(n7898), .Z(n4266) );
  XNOR2_X1 U4778 ( .A(n5798), .B(P2_IR_REG_29__SCAN_IN), .ZN(n5804) );
  INV_X1 U4779 ( .A(n4990), .ZN(n5070) );
  NAND2_X2 U4780 ( .A1(n7524), .A2(n7535), .ZN(n4989) );
  INV_X1 U4781 ( .A(n9949), .ZN(n4262) );
  INV_X1 U4782 ( .A(n4262), .ZN(P2_U3152) );
  INV_X1 U4783 ( .A(n4262), .ZN(n4264) );
  INV_X1 U4784 ( .A(n4266), .ZN(n4745) );
  OR2_X1 U4785 ( .A1(n9159), .A2(n9264), .ZN(n9160) );
  INV_X1 U4786 ( .A(n4971), .ZN(n8563) );
  BUF_X1 U4787 ( .A(n8694), .Z(n4267) );
  AND2_X1 U4788 ( .A1(n5800), .A2(n5804), .ZN(n5837) );
  NAND2_X1 U4789 ( .A1(n8150), .A2(n4507), .ZN(n8152) );
  NAND2_X1 U4790 ( .A1(n6505), .A2(n4266), .ZN(n9677) );
  INV_X2 U4791 ( .A(n7090), .ZN(n5032) );
  AND2_X1 U4792 ( .A1(n8933), .A2(n8932), .ZN(n8934) );
  NAND2_X1 U4793 ( .A1(n8739), .A2(n8771), .ZN(n7027) );
  INV_X1 U4794 ( .A(n7196), .ZN(n6891) );
  INV_X1 U4795 ( .A(n6505), .ZN(n6250) );
  OAI22_X1 U4796 ( .A1(n8231), .A2(n8052), .B1(n8236), .B2(n8254), .ZN(n8217)
         );
  CLKBUF_X2 U4797 ( .A(n4990), .Z(n4273) );
  NAND2_X1 U4798 ( .A1(n5070), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n4919) );
  INV_X1 U4799 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n4897) );
  INV_X1 U4800 ( .A(n7698), .ZN(n5793) );
  NAND4_X1 U4801 ( .A1(n5840), .A2(n5842), .A3(n5841), .A4(n5843), .ZN(n7916)
         );
  AOI211_X1 U4802 ( .C1(n9647), .C2(n8310), .A(n8090), .B(n8089), .ZN(n8091)
         );
  INV_X1 U4803 ( .A(n4989), .ZN(n4865) );
  NAND2_X1 U4804 ( .A1(n7524), .A2(n4868), .ZN(n4990) );
  NAND2_X2 U4805 ( .A1(n7234), .A2(n5663), .ZN(n7026) );
  NAND2_X2 U4806 ( .A1(n7236), .A2(n7235), .ZN(n7234) );
  NAND2_X2 U4807 ( .A1(n5621), .A2(n7151), .ZN(n4916) );
  NOR3_X2 U4808 ( .A1(n8288), .A2(n8358), .A3(n4472), .ZN(n4470) );
  NAND2_X2 U4809 ( .A1(n8163), .A2(n8162), .ZN(n8336) );
  BUF_X2 U4810 ( .A(n5620), .Z(n4265) );
  INV_X1 U4811 ( .A(n6695), .ZN(n6792) );
  OAI21_X2 U4812 ( .B1(n7166), .B2(n7878), .A(n7165), .ZN(n7167) );
  AND2_X1 U4814 ( .A1(n7525), .A2(n5804), .ZN(n6124) );
  INV_X1 U4815 ( .A(n7242), .ZN(n4268) );
  INV_X1 U4816 ( .A(n4268), .ZN(n4269) );
  NAND2_X1 U4818 ( .A1(n7015), .A2(n7743), .ZN(n7052) );
  OAI21_X2 U4819 ( .B1(n4714), .B2(n7167), .A(n4710), .ZN(n7427) );
  INV_X2 U4820 ( .A(n5838), .ZN(n6329) );
  NAND2_X1 U4821 ( .A1(n8192), .A2(n4665), .ZN(n8150) );
  NAND2_X1 U4822 ( .A1(n8194), .A2(n8193), .ZN(n8192) );
  AND2_X1 U4823 ( .A1(n7595), .A2(n6033), .ZN(n4740) );
  AND2_X1 U4824 ( .A1(n5719), .A2(n5717), .ZN(n8810) );
  INV_X1 U4825 ( .A(n7158), .ZN(n7209) );
  NAND2_X2 U4826 ( .A1(n6920), .A2(n7732), .ZN(n7866) );
  NAND4_X1 U4827 ( .A1(n4967), .A2(n4966), .A3(n4965), .A4(n4964), .ZN(n8848)
         );
  INV_X1 U4828 ( .A(n6919), .ZN(n9683) );
  INV_X1 U4829 ( .A(n7916), .ZN(n4698) );
  INV_X2 U4830 ( .A(n6968), .ZN(n4361) );
  NAND2_X1 U4831 ( .A1(n5057), .A2(n5056), .ZN(n5082) );
  INV_X1 U4832 ( .A(n7510), .ZN(n9590) );
  NAND2_X1 U4833 ( .A1(n4916), .A2(n6287), .ZN(n5485) );
  CLKBUF_X2 U4834 ( .A(n4992), .Z(n5241) );
  NAND2_X1 U4835 ( .A1(n5800), .A2(n7531), .ZN(n5838) );
  CLKBUF_X1 U4836 ( .A(P2_IR_REG_0__SCAN_IN), .Z(n9638) );
  NAND2_X1 U4837 ( .A1(n4815), .A2(n4814), .ZN(n4813) );
  AND3_X1 U4838 ( .A1(n4371), .A2(n4370), .A3(n8826), .ZN(n8837) );
  NAND2_X1 U4839 ( .A1(n4752), .A2(n6181), .ZN(n7651) );
  OR2_X1 U4840 ( .A1(n7863), .A2(n7862), .ZN(n4616) );
  NAND2_X1 U4841 ( .A1(n4496), .A2(n4499), .ZN(n7650) );
  NAND2_X1 U4842 ( .A1(n4799), .A2(n4797), .ZN(n8443) );
  NAND2_X1 U4843 ( .A1(n5346), .A2(n4299), .ZN(n4799) );
  NAND2_X1 U4844 ( .A1(n4577), .A2(n4575), .ZN(n9053) );
  AND2_X1 U4845 ( .A1(n9167), .A2(n9170), .ZN(n9281) );
  NAND2_X1 U4846 ( .A1(n4775), .A2(n5324), .ZN(n8484) );
  AND2_X1 U4847 ( .A1(n4454), .A2(n4327), .ZN(n4453) );
  NAND2_X1 U4848 ( .A1(n4352), .A2(n4351), .ZN(n9050) );
  OR3_X1 U4849 ( .A1(n8637), .A2(n4364), .A3(n4363), .ZN(n8628) );
  NAND2_X1 U4850 ( .A1(n5674), .A2(n4278), .ZN(n4593) );
  NAND2_X1 U4851 ( .A1(n7456), .A2(n4303), .ZN(n7482) );
  NAND2_X1 U4852 ( .A1(n6021), .A2(n6020), .ZN(n4741) );
  NAND2_X1 U4853 ( .A1(n4353), .A2(n4276), .ZN(n4539) );
  AND2_X1 U4854 ( .A1(n9401), .A2(n8595), .ZN(n7468) );
  NAND2_X1 U4855 ( .A1(n7441), .A2(n4569), .ZN(n9401) );
  NAND2_X1 U4856 ( .A1(n4790), .A2(n4792), .ZN(n7127) );
  OR2_X1 U4857 ( .A1(n5371), .A2(n4798), .ZN(n4797) );
  AND2_X1 U4858 ( .A1(n7225), .A2(n5662), .ZN(n7236) );
  NAND2_X1 U4859 ( .A1(n4765), .A2(n4763), .ZN(n7065) );
  OR2_X1 U4860 ( .A1(n9558), .A2(n9373), .ZN(n9425) );
  AND2_X1 U4861 ( .A1(n8700), .A2(n5664), .ZN(n4607) );
  AOI21_X2 U4862 ( .B1(n9652), .B2(n9661), .A(n9648), .ZN(n6895) );
  INV_X2 U4863 ( .A(n9661), .ZN(n8278) );
  INV_X2 U4864 ( .A(n9625), .ZN(n4270) );
  NAND2_X2 U4865 ( .A1(n6960), .A2(n8142), .ZN(n9661) );
  OAI21_X1 U4866 ( .B1(n6312), .B2(n4971), .A(n4567), .ZN(n7158) );
  AND2_X1 U4867 ( .A1(n8691), .A2(n8689), .ZN(n7230) );
  INV_X1 U4868 ( .A(n6716), .ZN(n7008) );
  AND3_X1 U4869 ( .A1(n5864), .A2(n5863), .A3(n5862), .ZN(n6979) );
  NAND4_X1 U4870 ( .A1(n4996), .A2(n4995), .A3(n4994), .A4(n4993), .ZN(n8847)
         );
  NAND2_X1 U4871 ( .A1(n7724), .A2(n7728), .ZN(n7867) );
  CLKBUF_X1 U4872 ( .A(n5070), .Z(n5585) );
  AND2_X2 U4873 ( .A1(n4900), .A2(n4899), .ZN(n5594) );
  AND2_X1 U4874 ( .A1(n4922), .A2(n4920), .ZN(n4573) );
  AND3_X1 U4875 ( .A1(n5825), .A2(n5826), .A3(n5824), .ZN(n6968) );
  AND2_X2 U4876 ( .A1(n4916), .A2(n5712), .ZN(n7090) );
  BUF_X2 U4877 ( .A(n5932), .Z(n7701) );
  NAND2_X1 U4878 ( .A1(n4869), .A2(n4868), .ZN(n4991) );
  CLKBUF_X3 U4879 ( .A(n6124), .Z(n7677) );
  BUF_X2 U4880 ( .A(n4866), .Z(n7524) );
  CLKBUF_X3 U4881 ( .A(n5838), .Z(n6266) );
  OR2_X2 U4882 ( .A1(n7864), .A2(n7895), .ZN(n7709) );
  AND2_X1 U4883 ( .A1(n7525), .A2(n7531), .ZN(n5839) );
  XNOR2_X1 U4884 ( .A(n4864), .B(n4863), .ZN(n4867) );
  XNOR2_X1 U4885 ( .A(n5777), .B(n5776), .ZN(n7865) );
  NAND2_X2 U4886 ( .A1(n5636), .A2(n5742), .ZN(n6346) );
  XNOR2_X1 U4887 ( .A(n5788), .B(n5796), .ZN(n6260) );
  NAND2_X1 U4888 ( .A1(n4950), .A2(n4949), .ZN(n4973) );
  XNOR2_X1 U4889 ( .A(n4907), .B(n4906), .ZN(n5636) );
  XNOR2_X1 U4890 ( .A(n4910), .B(n4909), .ZN(n5742) );
  OR2_X1 U4891 ( .A1(n4862), .A2(n9330), .ZN(n4864) );
  NAND2_X1 U4892 ( .A1(n4908), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4910) );
  NAND2_X1 U4893 ( .A1(n5792), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5788) );
  XNOR2_X1 U4894 ( .A(n4948), .B(n4927), .ZN(n4947) );
  NAND2_X1 U4895 ( .A1(n4925), .A2(n4926), .ZN(n4948) );
  NAND2_X2 U4896 ( .A1(n7698), .A2(n4264), .ZN(n8414) );
  NAND2_X2 U4897 ( .A1(n7698), .A2(P1_U3084), .ZN(n9340) );
  NOR2_X1 U4898 ( .A1(n4772), .A2(n4774), .ZN(n4771) );
  AND2_X1 U4899 ( .A1(n4851), .A2(n4793), .ZN(n4608) );
  NOR2_X1 U4900 ( .A1(n5785), .A2(n5784), .ZN(n5786) );
  NOR2_X1 U4901 ( .A1(n4310), .A2(n4804), .ZN(n4803) );
  NAND2_X1 U4902 ( .A1(n4663), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n4661) );
  NAND2_X1 U4903 ( .A1(n4852), .A2(n4795), .ZN(n4794) );
  INV_X1 U4904 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5259) );
  INV_X1 U4905 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n4795) );
  INV_X1 U4906 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5353) );
  NOR2_X1 U4907 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(P2_IR_REG_6__SCAN_IN), .ZN(
        n5763) );
  INV_X1 U4908 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n4881) );
  INV_X1 U4909 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n5138) );
  INV_X1 U4910 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n4877) );
  INV_X1 U4911 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n4848) );
  NOR2_X1 U4912 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5822) );
  NOR2_X2 U4913 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .ZN(
        n4847) );
  INV_X4 U4914 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  INV_X1 U4915 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n6225) );
  INV_X1 U4916 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n6246) );
  INV_X1 U4917 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n6222) );
  INV_X1 U4918 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n5782) );
  NOR2_X1 U4919 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(P1_IR_REG_6__SCAN_IN), .ZN(
        n4787) );
  NAND2_X1 U4920 ( .A1(n6346), .A2(n7698), .ZN(n5000) );
  NAND4_X1 U4921 ( .A1(n4873), .A2(n4872), .A3(n4871), .A4(n4870), .ZN(n5653)
         );
  INV_X2 U4922 ( .A(n7352), .ZN(n7423) );
  NAND2_X2 U4923 ( .A1(n5683), .A2(n5682), .ZN(n9099) );
  MUX2_X2 U4924 ( .A(n9182), .B(n9288), .S(n4270), .Z(n9183) );
  OAI21_X2 U4925 ( .B1(n7026), .B2(n4606), .A(n4605), .ZN(n9557) );
  XNOR2_X2 U4926 ( .A(n8802), .B(n8849), .ZN(n5713) );
  NAND3_X4 U4927 ( .A1(n4573), .A2(n4921), .A3(n4919), .ZN(n8849) );
  INV_X1 U4928 ( .A(n6217), .ZN(n5789) );
  AND4_X1 U4929 ( .A1(n5767), .A2(n5766), .A3(n5765), .A4(n5892), .ZN(n5768)
         );
  OR2_X1 U4930 ( .A1(n9215), .A2(n8437), .ZN(n8638) );
  NAND2_X1 U4931 ( .A1(n5559), .A2(n5558), .ZN(n5581) );
  OAI21_X1 U4932 ( .B1(n5303), .B2(n5302), .A(n5301), .ZN(n5326) );
  OR2_X1 U4933 ( .A1(n8321), .A2(n8122), .ZN(n8113) );
  NAND2_X1 U4934 ( .A1(n4366), .A2(n4365), .ZN(n8637) );
  NAND2_X1 U4935 ( .A1(n8626), .A2(n8679), .ZN(n4366) );
  AND2_X1 U4936 ( .A1(n4438), .A2(n7824), .ZN(n4437) );
  OR2_X1 U4937 ( .A1(n7823), .A2(n4439), .ZN(n4438) );
  NOR2_X1 U4938 ( .A1(n8162), .A2(n7819), .ZN(n4439) );
  NAND2_X1 U4939 ( .A1(n4392), .A2(n4391), .ZN(n4390) );
  NOR2_X1 U4940 ( .A1(n8629), .A2(n8679), .ZN(n4391) );
  NAND2_X1 U4941 ( .A1(n8630), .A2(n8638), .ZN(n4392) );
  INV_X1 U4942 ( .A(n4652), .ZN(n4651) );
  OAI21_X1 U4943 ( .B1(n5580), .B2(n4653), .A(n5701), .ZN(n4652) );
  AND2_X1 U4944 ( .A1(n5374), .A2(n4622), .ZN(n4618) );
  INV_X1 U4945 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n5232) );
  INV_X1 U4946 ( .A(n7641), .ZN(n4756) );
  NAND2_X1 U4947 ( .A1(n8372), .A2(n8050), .ZN(n4727) );
  OR2_X1 U4948 ( .A1(n8287), .A2(n7683), .ZN(n7786) );
  OR2_X1 U4949 ( .A1(n7780), .A2(n7907), .ZN(n8048) );
  NAND2_X1 U4950 ( .A1(n4838), .A2(n4773), .ZN(n4772) );
  INV_X1 U4951 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n4773) );
  INV_X1 U4952 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5783) );
  INV_X1 U4953 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n5892) );
  INV_X1 U4954 ( .A(n5149), .ZN(n4786) );
  AND2_X1 U4955 ( .A1(n7407), .A2(n4785), .ZN(n4784) );
  OR2_X1 U4956 ( .A1(n7378), .A2(n4786), .ZN(n4785) );
  NOR2_X1 U4957 ( .A1(n4604), .A2(n5691), .ZN(n4603) );
  INV_X1 U4958 ( .A(n5690), .ZN(n4604) );
  AND2_X1 U4959 ( .A1(n4579), .A2(n4578), .ZN(n4574) );
  INV_X1 U4960 ( .A(n5687), .ZN(n4578) );
  OR2_X1 U4961 ( .A1(n8456), .A2(n9069), .ZN(n8729) );
  OR2_X1 U4962 ( .A1(n9228), .A2(n9087), .ZN(n8627) );
  NAND2_X1 U4963 ( .A1(n4369), .A2(n4367), .ZN(n8600) );
  NOR2_X1 U4964 ( .A1(n9139), .A2(n4368), .ZN(n4367) );
  INV_X1 U4965 ( .A(n5330), .ZN(n4368) );
  OR2_X1 U4966 ( .A1(n9444), .A2(n9413), .ZN(n8608) );
  AOI21_X1 U4967 ( .B1(n4659), .B2(n4657), .A(n4656), .ZN(n4655) );
  INV_X1 U4968 ( .A(n4659), .ZN(n4658) );
  INV_X1 U4969 ( .A(n5490), .ZN(n4656) );
  NAND2_X1 U4970 ( .A1(n5427), .A2(n5426), .ZN(n4647) );
  NAND2_X1 U4971 ( .A1(n5402), .A2(n5401), .ZN(n5427) );
  OR2_X1 U4972 ( .A1(n5400), .A2(n5399), .ZN(n5402) );
  AOI21_X1 U4973 ( .B1(n4642), .B2(n4644), .A(n4319), .ZN(n4641) );
  NAND2_X1 U4974 ( .A1(n4901), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n4663) );
  INV_X1 U4975 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4901) );
  NAND2_X1 U4976 ( .A1(n7622), .A2(n4742), .ZN(n7555) );
  AND2_X1 U4977 ( .A1(n6131), .A2(n4743), .ZN(n4742) );
  INV_X1 U4978 ( .A(n6141), .ZN(n4743) );
  AND2_X1 U4979 ( .A1(n7538), .A2(n4329), .ZN(n4750) );
  NAND2_X1 U4980 ( .A1(n4498), .A2(n4291), .ZN(n4749) );
  NAND2_X1 U4981 ( .A1(n5778), .A2(n6503), .ZN(n5820) );
  NOR2_X1 U4982 ( .A1(n6505), .A2(n4745), .ZN(n4744) );
  OR2_X1 U4983 ( .A1(n7065), .A2(n5954), .ZN(n4480) );
  OAI21_X1 U4984 ( .B1(n8304), .B2(n7692), .A(n7850), .ZN(n4508) );
  INV_X1 U4985 ( .A(n6324), .ZN(n6363) );
  NAND2_X1 U4986 ( .A1(n4407), .A2(n4406), .ZN(n6521) );
  INV_X1 U4987 ( .A(n6437), .ZN(n4406) );
  AND2_X1 U4988 ( .A1(n8079), .A2(n8070), .ZN(n8068) );
  NAND2_X1 U4989 ( .A1(n4685), .A2(n4274), .ZN(n8107) );
  AND2_X1 U4990 ( .A1(n4510), .A2(n7811), .ZN(n8194) );
  OR2_X1 U4991 ( .A1(n8219), .A2(n4325), .ZN(n4510) );
  OR2_X1 U4992 ( .A1(n8361), .A2(n8254), .ZN(n8218) );
  INV_X1 U4993 ( .A(n4715), .ZN(n4714) );
  INV_X1 U4994 ( .A(n4711), .ZN(n4710) );
  OAI21_X1 U4995 ( .B1(n7315), .B2(n4712), .A(n4322), .ZN(n4711) );
  NAND2_X1 U4996 ( .A1(n9639), .A2(n4302), .ZN(n7073) );
  NAND2_X1 U4997 ( .A1(n6507), .A2(n7708), .ZN(n8213) );
  INV_X1 U4998 ( .A(n8285), .ZN(n9656) );
  NAND2_X1 U4999 ( .A1(n6170), .A2(n6169), .ZN(n8321) );
  NAND2_X1 U5000 ( .A1(n5789), .A2(n5787), .ZN(n5792) );
  NAND2_X1 U5001 ( .A1(n6005), .A2(n4356), .ZN(n6217) );
  AND2_X1 U5002 ( .A1(n5786), .A2(n4330), .ZN(n4356) );
  INV_X1 U5003 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n4691) );
  CLKBUF_X1 U5004 ( .A(n5889), .Z(n5890) );
  INV_X1 U5005 ( .A(n5300), .ZN(n4418) );
  OR2_X1 U5006 ( .A1(n5507), .A2(n5508), .ZN(n4812) );
  NAND2_X1 U5007 ( .A1(n4377), .A2(n4375), .ZN(n4374) );
  AND2_X1 U5008 ( .A1(n8678), .A2(n4376), .ZN(n4375) );
  NAND2_X1 U5009 ( .A1(n8668), .A2(n4378), .ZN(n4377) );
  NAND2_X1 U5010 ( .A1(n8568), .A2(n8674), .ZN(n4376) );
  NOR2_X1 U5011 ( .A1(n8932), .A2(n4598), .ZN(n4597) );
  AND2_X1 U5012 ( .A1(n5694), .A2(n5693), .ZN(n4590) );
  NAND2_X1 U5013 ( .A1(n8986), .A2(n8995), .ZN(n4591) );
  AND2_X1 U5014 ( .A1(n5732), .A2(n4556), .ZN(n4555) );
  NAND2_X1 U5015 ( .A1(n4558), .A2(n4557), .ZN(n4556) );
  INV_X1 U5016 ( .A(n5685), .ZN(n4583) );
  NAND2_X1 U5017 ( .A1(n9119), .A2(n8600), .ZN(n9097) );
  NAND2_X1 U5018 ( .A1(n4539), .A2(n4284), .ZN(n9117) );
  OR2_X1 U5019 ( .A1(n9254), .A2(n5678), .ZN(n9116) );
  AND2_X1 U5020 ( .A1(n5675), .A2(n4844), .ZN(n4592) );
  INV_X1 U5021 ( .A(n5000), .ZN(n5381) );
  NAND2_X1 U5022 ( .A1(n5715), .A2(n5714), .ZN(n8804) );
  AOI21_X1 U5023 ( .B1(n5746), .B2(n9550), .A(n5745), .ZN(n8922) );
  AND2_X1 U5024 ( .A1(n8841), .A2(n8911), .ZN(n5745) );
  INV_X1 U5025 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n4906) );
  NAND2_X1 U5026 ( .A1(n4859), .A2(n4803), .ZN(n4908) );
  XNOR2_X1 U5027 ( .A(n4884), .B(P1_IR_REG_26__SCAN_IN), .ZN(n5601) );
  OR2_X1 U5028 ( .A1(n4878), .A2(n4877), .ZN(n4879) );
  NAND2_X1 U5029 ( .A1(n4633), .A2(n4634), .ZN(n5204) );
  OR2_X1 U5030 ( .A1(n5152), .A2(n4637), .ZN(n4633) );
  NAND2_X1 U5031 ( .A1(n6184), .A2(n6183), .ZN(n8314) );
  NAND2_X1 U5032 ( .A1(n6209), .A2(n6208), .ZN(n8100) );
  INV_X1 U5033 ( .A(n6346), .ZN(n6290) );
  NOR2_X1 U5034 ( .A1(n7731), .A2(n4432), .ZN(n4431) );
  NAND2_X1 U5035 ( .A1(n4433), .A2(n6800), .ZN(n4432) );
  NAND2_X1 U5036 ( .A1(n7722), .A2(n7721), .ZN(n4433) );
  INV_X1 U5037 ( .A(n7823), .ZN(n4441) );
  INV_X1 U5038 ( .A(n7847), .ZN(n4455) );
  NOR2_X1 U5039 ( .A1(n7849), .A2(n7857), .ZN(n4457) );
  NOR2_X1 U5040 ( .A1(n7846), .A2(n4459), .ZN(n4458) );
  INV_X1 U5041 ( .A(n7849), .ZN(n4459) );
  NAND2_X1 U5042 ( .A1(n8640), .A2(n8679), .ZN(n4393) );
  NOR2_X1 U5043 ( .A1(n4557), .A2(n4389), .ZN(n4388) );
  NAND2_X1 U5044 ( .A1(n8645), .A2(n4333), .ZN(n4389) );
  AOI21_X1 U5045 ( .B1(n4453), .B2(n4456), .A(n4452), .ZN(n4451) );
  INV_X1 U5046 ( .A(n4458), .ZN(n4456) );
  INV_X1 U5047 ( .A(n7851), .ZN(n4452) );
  INV_X1 U5048 ( .A(n4644), .ZN(n4643) );
  INV_X1 U5049 ( .A(n4487), .ZN(n4484) );
  INV_X1 U5050 ( .A(n7579), .ZN(n4501) );
  OAI21_X1 U5051 ( .B1(n7821), .B2(n4436), .A(n4434), .ZN(n4442) );
  INV_X1 U5052 ( .A(n4451), .ZN(n4450) );
  AOI21_X1 U5053 ( .B1(n4451), .B2(n4449), .A(n7893), .ZN(n4448) );
  INV_X1 U5054 ( .A(n4453), .ZN(n4449) );
  OR2_X1 U5055 ( .A1(n9414), .A2(n9373), .ZN(n8755) );
  NOR2_X1 U5056 ( .A1(n9228), .A2(n9231), .ZN(n4531) );
  OAI21_X1 U5057 ( .B1(n7523), .B2(n7522), .A(n7521), .ZN(n7696) );
  INV_X1 U5058 ( .A(n5582), .ZN(n4653) );
  INV_X1 U5059 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n5329) );
  INV_X1 U5060 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n5256) );
  INV_X1 U5061 ( .A(SI_12_), .ZN(n5205) );
  INV_X1 U5062 ( .A(n6049), .ZN(n4762) );
  OR2_X1 U5063 ( .A1(n7580), .A2(n4501), .ZN(n4499) );
  AND2_X1 U5064 ( .A1(n4732), .A2(n8092), .ZN(n4730) );
  NAND2_X1 U5065 ( .A1(n8118), .A2(n8059), .ZN(n4738) );
  NOR2_X1 U5066 ( .A1(n8334), .A2(n8341), .ZN(n4463) );
  AND2_X1 U5067 ( .A1(n7822), .A2(n8136), .ZN(n7818) );
  AND2_X1 U5068 ( .A1(n8176), .A2(n8177), .ZN(n4665) );
  OR2_X1 U5069 ( .A1(n8341), .A2(n8056), .ZN(n7820) );
  AND2_X1 U5070 ( .A1(n7792), .A2(n4677), .ZN(n4676) );
  NOR2_X1 U5071 ( .A1(n8266), .A2(n4678), .ZN(n4677) );
  INV_X1 U5072 ( .A(n7786), .ZN(n4678) );
  NOR2_X1 U5073 ( .A1(n7780), .A2(n4522), .ZN(n4521) );
  NOR2_X1 U5074 ( .A1(n4518), .A2(n4521), .ZN(n4517) );
  INV_X1 U5075 ( .A(n4519), .ZN(n4518) );
  NAND2_X1 U5076 ( .A1(n7884), .A2(n7776), .ZN(n4514) );
  NOR2_X1 U5077 ( .A1(n7883), .A2(n4520), .ZN(n4519) );
  AND2_X1 U5078 ( .A1(n7168), .A2(n4671), .ZN(n4670) );
  NAND2_X1 U5079 ( .A1(n4672), .A2(n7756), .ZN(n4671) );
  NAND2_X1 U5080 ( .A1(n4506), .A2(n7753), .ZN(n7075) );
  NAND2_X1 U5081 ( .A1(n7074), .A2(n7758), .ZN(n4506) );
  AND2_X1 U5082 ( .A1(n4326), .A2(n7872), .ZN(n4704) );
  NAND2_X1 U5083 ( .A1(n8036), .A2(n9386), .ZN(n8286) );
  NOR2_X1 U5084 ( .A1(n7393), .A2(n8378), .ZN(n8036) );
  INV_X1 U5085 ( .A(n9677), .ZN(n6241) );
  NOR2_X2 U5086 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), .ZN(
        n5781) );
  OR2_X1 U5087 ( .A1(n7494), .A2(n7493), .ZN(n4833) );
  INV_X1 U5088 ( .A(n4833), .ZN(n4824) );
  INV_X1 U5089 ( .A(n8498), .ZN(n4779) );
  NAND2_X1 U5090 ( .A1(n8498), .A2(n4778), .ZN(n4777) );
  INV_X1 U5091 ( .A(n5398), .ZN(n4778) );
  INV_X1 U5092 ( .A(n4823), .ZN(n4822) );
  OAI21_X1 U5093 ( .B1(n4830), .B2(n4824), .A(n5275), .ZN(n4823) );
  INV_X1 U5094 ( .A(n4821), .ZN(n4820) );
  AOI21_X1 U5095 ( .B1(n4822), .B2(n4824), .A(n4332), .ZN(n4821) );
  AOI21_X1 U5096 ( .B1(n4827), .B2(n5253), .A(n4826), .ZN(n4825) );
  INV_X1 U5097 ( .A(n8424), .ZN(n4826) );
  NOR2_X1 U5098 ( .A1(n8973), .A2(n8990), .ZN(n4538) );
  OR2_X1 U5099 ( .A1(n8973), .A2(n8654), .ZN(n8736) );
  NOR2_X1 U5100 ( .A1(n4582), .A2(n5687), .ZN(n4576) );
  NAND2_X1 U5101 ( .A1(n9098), .A2(n8623), .ZN(n4566) );
  INV_X1 U5102 ( .A(n8772), .ZN(n4562) );
  INV_X1 U5103 ( .A(n8623), .ZN(n4563) );
  OR2_X1 U5104 ( .A1(n9444), .A2(n9451), .ZN(n4534) );
  INV_X1 U5105 ( .A(n4916), .ZN(n5710) );
  AND2_X1 U5106 ( .A1(n8749), .A2(n8689), .ZN(n5719) );
  NOR2_X1 U5107 ( .A1(n9105), .A2(n9231), .ZN(n9089) );
  INV_X1 U5108 ( .A(n4587), .ZN(n4586) );
  OAI21_X1 U5109 ( .B1(n5668), .B2(n4588), .A(n8706), .ZN(n4587) );
  NAND2_X1 U5110 ( .A1(n4589), .A2(n5668), .ZN(n9418) );
  INV_X1 U5111 ( .A(n9415), .ZN(n4589) );
  INV_X1 U5112 ( .A(n7402), .ZN(n5616) );
  XNOR2_X1 U5113 ( .A(n7696), .B(n7695), .ZN(n7694) );
  AND2_X1 U5114 ( .A1(n5582), .A2(n5563), .ZN(n5580) );
  OAI21_X1 U5115 ( .B1(n5535), .B2(n5534), .A(n5533), .ZN(n5557) );
  AND2_X1 U5116 ( .A1(n5558), .A2(n5539), .ZN(n5556) );
  NAND2_X1 U5117 ( .A1(n4858), .A2(n4890), .ZN(n4804) );
  NAND2_X1 U5118 ( .A1(n4876), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4878) );
  AOI21_X1 U5119 ( .B1(n5308), .B2(P1_IR_REG_31__SCAN_IN), .A(n4426), .ZN(
        n4425) );
  NAND2_X1 U5120 ( .A1(n4427), .A2(n4881), .ZN(n4426) );
  AOI21_X1 U5121 ( .B1(n5374), .B2(n4620), .A(n4340), .ZN(n4619) );
  INV_X1 U5122 ( .A(n5350), .ZN(n4620) );
  INV_X1 U5123 ( .A(SI_16_), .ZN(n5304) );
  NOR2_X1 U5124 ( .A1(n5209), .A2(n4794), .ZN(n5257) );
  INV_X1 U5125 ( .A(SI_13_), .ZN(n5233) );
  NAND2_X1 U5126 ( .A1(n5231), .A2(n5230), .ZN(n5254) );
  NAND2_X1 U5127 ( .A1(n4399), .A2(n4396), .ZN(n5231) );
  AOI21_X1 U5128 ( .B1(n4631), .B2(n4637), .A(n4318), .ZN(n4630) );
  NAND2_X1 U5129 ( .A1(n5152), .A2(n4631), .ZN(n4399) );
  NAND2_X1 U5130 ( .A1(n4495), .A2(n4754), .ZN(n4494) );
  NAND3_X1 U5131 ( .A1(n4741), .A2(n4740), .A3(n4754), .ZN(n4493) );
  XNOR2_X1 U5132 ( .A(n4502), .B(n7003), .ZN(n5808) );
  AND2_X1 U5133 ( .A1(n7918), .A2(n6783), .ZN(n5809) );
  NAND2_X1 U5134 ( .A1(n7554), .A2(n4476), .ZN(n6152) );
  OR2_X1 U5135 ( .A1(n6098), .A2(n7617), .ZN(n6112) );
  OR2_X1 U5136 ( .A1(n6122), .A2(n7626), .ZN(n6134) );
  AND2_X1 U5137 ( .A1(n4481), .A2(n7633), .ZN(n4275) );
  OR2_X1 U5138 ( .A1(n7064), .A2(n5954), .ZN(n4481) );
  NOR2_X1 U5139 ( .A1(n5808), .A2(n5809), .ZN(n5818) );
  AND2_X1 U5140 ( .A1(n7865), .A2(n7895), .ZN(n6258) );
  OR2_X1 U5141 ( .A1(n7405), .A2(n6244), .ZN(n6360) );
  OR2_X1 U5142 ( .A1(n5913), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n5939) );
  NAND2_X1 U5143 ( .A1(n8128), .A2(n4274), .ZN(n4683) );
  INV_X1 U5144 ( .A(n4469), .ZN(n4467) );
  NAND2_X1 U5145 ( .A1(n4733), .A2(n4738), .ZN(n4732) );
  INV_X1 U5146 ( .A(n4736), .ZN(n4733) );
  AOI21_X1 U5147 ( .B1(n4737), .B2(n4689), .A(n4688), .ZN(n4736) );
  NAND2_X1 U5148 ( .A1(n4737), .A2(n4738), .ZN(n4734) );
  NAND2_X1 U5149 ( .A1(n4686), .A2(n4689), .ZN(n4685) );
  OR2_X1 U5150 ( .A1(n8325), .A2(n7686), .ZN(n7828) );
  NOR2_X1 U5151 ( .A1(n8329), .A2(n8154), .ZN(n4739) );
  INV_X1 U5152 ( .A(n7890), .ZN(n8137) );
  NOR2_X2 U5153 ( .A1(n8135), .A2(n8137), .ZN(n8134) );
  OR2_X1 U5154 ( .A1(n8191), .A2(n8180), .ZN(n4837) );
  AOI21_X1 U5155 ( .B1(n8201), .B2(n8208), .A(n8054), .ZN(n8187) );
  AND2_X1 U5156 ( .A1(n8351), .A2(n8196), .ZN(n8054) );
  NOR2_X1 U5157 ( .A1(n8224), .A2(n8351), .ZN(n8202) );
  OR2_X1 U5158 ( .A1(n6075), .A2(n6074), .ZN(n6086) );
  NOR2_X1 U5159 ( .A1(n8221), .A2(n7798), .ZN(n4511) );
  NAND2_X1 U5160 ( .A1(n4323), .A2(n4727), .ZN(n4720) );
  NAND2_X1 U5161 ( .A1(n8279), .A2(n4722), .ZN(n4721) );
  NAND2_X1 U5162 ( .A1(n4666), .A2(n4519), .ZN(n4523) );
  INV_X1 U5163 ( .A(n4523), .ZN(n7432) );
  NAND2_X1 U5164 ( .A1(n7075), .A2(n4670), .ZN(n4667) );
  AOI21_X1 U5165 ( .B1(n4670), .B2(n7759), .A(n4669), .ZN(n4668) );
  INV_X1 U5166 ( .A(n7769), .ZN(n4669) );
  NOR2_X1 U5167 ( .A1(n7315), .A2(n4713), .ZN(n4715) );
  NAND2_X1 U5168 ( .A1(n7167), .A2(n7881), .ZN(n7313) );
  AND2_X1 U5169 ( .A1(n7758), .A2(n7753), .ZN(n7877) );
  NAND2_X1 U5170 ( .A1(n7045), .A2(n7874), .ZN(n9639) );
  NAND2_X1 U5171 ( .A1(n6911), .A2(n6795), .ZN(n6796) );
  NAND2_X1 U5172 ( .A1(n6796), .A2(n7872), .ZN(n6982) );
  AND2_X1 U5173 ( .A1(n7865), .A2(n5807), .ZN(n7897) );
  INV_X1 U5174 ( .A(n8284), .ZN(n9653) );
  INV_X1 U5175 ( .A(n8213), .ZN(n9660) );
  NAND2_X1 U5176 ( .A1(n6363), .A2(n7528), .ZN(n8284) );
  AND2_X1 U5177 ( .A1(n6504), .A2(n7895), .ZN(n9652) );
  INV_X1 U5178 ( .A(n8379), .ZN(n9727) );
  NAND2_X1 U5179 ( .A1(n5836), .A2(n4696), .ZN(n6695) );
  INV_X1 U5180 ( .A(n4697), .ZN(n4696) );
  OAI21_X1 U5181 ( .B1(n6300), .B2(n5911), .A(n5835), .ZN(n4697) );
  AND2_X1 U5182 ( .A1(n6241), .A2(n7901), .ZN(n8379) );
  INV_X1 U5183 ( .A(n9728), .ZN(n8380) );
  NAND2_X1 U5184 ( .A1(n4768), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6223) );
  AND2_X1 U5185 ( .A1(n4771), .A2(n5782), .ZN(n4769) );
  NAND2_X1 U5186 ( .A1(n5770), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5774) );
  AND2_X1 U5187 ( .A1(n4770), .A2(n4279), .ZN(n4444) );
  INV_X1 U5188 ( .A(n4772), .ZN(n4770) );
  NAND2_X1 U5189 ( .A1(n6034), .A2(n4838), .ZN(n6070) );
  AND2_X1 U5190 ( .A1(n4828), .A2(n4833), .ZN(n4827) );
  INV_X1 U5191 ( .A(n5275), .ZN(n4828) );
  INV_X1 U5192 ( .A(n5253), .ZN(n4830) );
  XNOR2_X1 U5193 ( .A(n4981), .B(n5032), .ZN(n4984) );
  NAND2_X1 U5194 ( .A1(n5445), .A2(n5444), .ZN(n5464) );
  NAND2_X1 U5195 ( .A1(n8450), .A2(n8452), .ZN(n5445) );
  AOI21_X1 U5196 ( .B1(n4784), .B2(n4786), .A(n4305), .ZN(n4781) );
  INV_X1 U5197 ( .A(n5522), .ZN(n5542) );
  NAND2_X1 U5198 ( .A1(n5487), .A2(n4814), .ZN(n4806) );
  AND2_X1 U5199 ( .A1(n7151), .A2(n9123), .ZN(n8832) );
  NAND2_X1 U5200 ( .A1(n5601), .A2(n4892), .ZN(n6287) );
  NAND2_X1 U5201 ( .A1(n4865), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n4873) );
  NOR2_X1 U5202 ( .A1(n8892), .A2(n4359), .ZN(n9527) );
  AND2_X1 U5203 ( .A1(n8897), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n4359) );
  AND2_X1 U5204 ( .A1(n8722), .A2(n8783), .ZN(n8932) );
  AND2_X1 U5205 ( .A1(n5477), .A2(n5476), .ZN(n5731) );
  NAND2_X1 U5206 ( .A1(n9022), .A2(n9021), .ZN(n9020) );
  INV_X1 U5207 ( .A(n9054), .ZN(n4351) );
  INV_X1 U5208 ( .A(n9038), .ZN(n9069) );
  AOI21_X1 U5209 ( .B1(n4580), .B2(n4582), .A(n4312), .ZN(n4579) );
  AND2_X1 U5210 ( .A1(n8624), .A2(n8772), .ZN(n9082) );
  OR2_X1 U5211 ( .A1(n9097), .A2(n9098), .ZN(n9095) );
  NAND2_X1 U5212 ( .A1(n5729), .A2(n9125), .ZN(n9119) );
  AOI21_X1 U5213 ( .B1(n4542), .B2(n4276), .A(n4541), .ZN(n4540) );
  INV_X1 U5214 ( .A(n8709), .ZN(n4542) );
  NAND2_X1 U5215 ( .A1(n7468), .A2(n8709), .ZN(n7467) );
  NAND2_X1 U5216 ( .A1(n5725), .A2(n4571), .ZN(n7441) );
  NOR2_X1 U5217 ( .A1(n8706), .A2(n4572), .ZN(n4571) );
  INV_X1 U5218 ( .A(n8606), .ZN(n4572) );
  NOR2_X1 U5219 ( .A1(n9425), .A2(n9451), .ZN(n9428) );
  NAND2_X1 U5220 ( .A1(n7026), .A2(n7027), .ZN(n7025) );
  INV_X1 U5221 ( .A(n4267), .ZN(n5656) );
  NAND2_X1 U5222 ( .A1(n4265), .A2(n8801), .ZN(n7089) );
  NAND2_X1 U5223 ( .A1(n8565), .A2(n8564), .ZN(n8908) );
  NAND2_X1 U5224 ( .A1(n5736), .A2(n5735), .ZN(n9550) );
  INV_X1 U5225 ( .A(n9550), .ZN(n9399) );
  INV_X1 U5226 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n4863) );
  AND2_X1 U5227 ( .A1(n5490), .A2(n5475), .ZN(n5488) );
  XNOR2_X1 U5228 ( .A(n5618), .B(n4858), .ZN(n7374) );
  NAND2_X1 U5229 ( .A1(n4647), .A2(n5428), .ZN(n5446) );
  NAND2_X1 U5230 ( .A1(n4839), .A2(n4430), .ZN(n4429) );
  NOR2_X1 U5231 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), .ZN(
        n4430) );
  NAND2_X1 U5232 ( .A1(n4621), .A2(n5350), .ZN(n5375) );
  NAND2_X1 U5233 ( .A1(n5328), .A2(n4622), .ZN(n4621) );
  AOI21_X1 U5234 ( .B1(n5103), .B2(n4627), .A(n4317), .ZN(n4626) );
  INV_X1 U5235 ( .A(n5085), .ZN(n4627) );
  NOR2_X1 U5236 ( .A1(n4628), .A2(n4625), .ZN(n4624) );
  INV_X1 U5237 ( .A(n5103), .ZN(n4628) );
  INV_X1 U5238 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n4953) );
  NAND2_X1 U5239 ( .A1(n4490), .A2(n4300), .ZN(n4489) );
  NAND2_X1 U5240 ( .A1(n6710), .A2(n4492), .ZN(n4491) );
  INV_X1 U5241 ( .A(n4753), .ZN(n4490) );
  NAND2_X1 U5242 ( .A1(n7651), .A2(n6182), .ZN(n7539) );
  NAND2_X1 U5243 ( .A1(n6873), .A2(n4766), .ZN(n4765) );
  AND2_X1 U5244 ( .A1(n4277), .A2(n6872), .ZN(n4766) );
  NAND2_X1 U5245 ( .A1(n7065), .A2(n7064), .ZN(n7063) );
  NAND2_X1 U5246 ( .A1(n6873), .A2(n6872), .ZN(n6871) );
  INV_X1 U5247 ( .A(n7673), .ZN(n7631) );
  NAND2_X1 U5248 ( .A1(n5959), .A2(n5958), .ZN(n7636) );
  NAND2_X1 U5249 ( .A1(n6019), .A2(n6018), .ZN(n8287) );
  NAND2_X1 U5250 ( .A1(n4611), .A2(n4308), .ZN(n4525) );
  INV_X1 U5251 ( .A(n7856), .ZN(n7853) );
  OAI22_X1 U5252 ( .A1(n4509), .A2(n4508), .B1(n7693), .B2(n7854), .ZN(n7706)
         );
  NAND2_X1 U5253 ( .A1(n6360), .A2(n9675), .ZN(n9669) );
  INV_X1 U5254 ( .A(n6258), .ZN(n7901) );
  NAND2_X1 U5255 ( .A1(n6363), .A2(n6261), .ZN(n8285) );
  NAND2_X1 U5256 ( .A1(n6191), .A2(n6190), .ZN(n8087) );
  OR2_X1 U5257 ( .A1(n6434), .A2(n4408), .ZN(n4407) );
  AND2_X1 U5258 ( .A1(n6445), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n4408) );
  OR2_X1 U5259 ( .A1(n6529), .A2(n6528), .ZN(n4402) );
  NAND2_X1 U5260 ( .A1(n6368), .A2(n7528), .ZN(n9628) );
  INV_X1 U5261 ( .A(n9629), .ZN(n9627) );
  NAND2_X1 U5262 ( .A1(n7704), .A2(n7703), .ZN(n8298) );
  NAND2_X1 U5263 ( .A1(n4321), .A2(n4469), .ZN(n4468) );
  AOI21_X1 U5264 ( .B1(n8100), .B2(n9656), .A(n4693), .ZN(n4692) );
  NAND2_X1 U5265 ( .A1(n4695), .A2(n8213), .ZN(n4694) );
  AND2_X1 U5266 ( .A1(n8067), .A2(n8066), .ZN(n4693) );
  AND2_X1 U5267 ( .A1(n6321), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9675) );
  NAND2_X1 U5269 ( .A1(n6217), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5790) );
  OR2_X1 U5270 ( .A1(n5894), .A2(n5893), .ZN(n6522) );
  AND2_X1 U5271 ( .A1(n5086), .A2(n4328), .ZN(n4567) );
  NAND2_X1 U5272 ( .A1(n5263), .A2(n5262), .ZN(n8430) );
  AND2_X1 U5273 ( .A1(n5627), .A2(n8475), .ZN(n5623) );
  OR2_X1 U5274 ( .A1(n6317), .A2(n4971), .ZN(n5112) );
  NAND2_X1 U5275 ( .A1(n7456), .A2(n5200), .ZN(n7484) );
  NAND2_X1 U5276 ( .A1(n4424), .A2(n4812), .ZN(n4423) );
  NAND2_X1 U5277 ( .A1(n4810), .A2(n4813), .ZN(n4424) );
  INV_X1 U5278 ( .A(n8459), .ZN(n4422) );
  NAND2_X1 U5279 ( .A1(n8541), .A2(n4417), .ZN(n4775) );
  NOR2_X1 U5280 ( .A1(n4418), .A2(n8466), .ZN(n4417) );
  NAND2_X1 U5281 ( .A1(n5492), .A2(n5491), .ZN(n9204) );
  NAND2_X1 U5282 ( .A1(n5457), .A2(n5456), .ZN(n9215) );
  INV_X1 U5283 ( .A(n8475), .ZN(n8554) );
  NAND2_X1 U5284 ( .A1(n4374), .A2(n8682), .ZN(n4370) );
  NAND2_X1 U5285 ( .A1(n4373), .A2(n4372), .ZN(n4371) );
  INV_X1 U5286 ( .A(n5620), .ZN(n8558) );
  INV_X1 U5287 ( .A(n9201), .ZN(n9039) );
  INV_X1 U5288 ( .A(n4599), .ZN(n5709) );
  NAND2_X1 U5289 ( .A1(n7183), .A2(n7182), .ZN(n9162) );
  NAND2_X1 U5290 ( .A1(n6346), .A2(n4282), .ZN(n4929) );
  INV_X1 U5291 ( .A(n8908), .ZN(n9284) );
  AOI21_X1 U5292 ( .B1(n7723), .B2(n7709), .A(n4431), .ZN(n7740) );
  INV_X1 U5293 ( .A(n4437), .ZN(n4436) );
  AOI21_X1 U5294 ( .B1(n4437), .B2(n4440), .A(n4435), .ZN(n4434) );
  INV_X1 U5295 ( .A(n7826), .ZN(n4435) );
  NAND2_X1 U5296 ( .A1(n4441), .A2(n7820), .ZN(n4440) );
  NAND2_X1 U5297 ( .A1(n4455), .A2(n4458), .ZN(n4454) );
  INV_X1 U5298 ( .A(n8648), .ZN(n4386) );
  OR2_X1 U5299 ( .A1(n8305), .A2(n7691), .ZN(n7849) );
  NAND2_X1 U5300 ( .A1(n6792), .A2(n4466), .ZN(n6798) );
  NAND2_X1 U5301 ( .A1(n4531), .A2(n9305), .ZN(n4530) );
  AND2_X1 U5302 ( .A1(n4660), .A2(n5488), .ZN(n4659) );
  INV_X1 U5303 ( .A(n5470), .ZN(n4657) );
  INV_X1 U5304 ( .A(n4794), .ZN(n4793) );
  NAND2_X1 U5305 ( .A1(n4429), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4427) );
  INV_X1 U5306 ( .A(n5228), .ZN(n4398) );
  AND2_X1 U5307 ( .A1(n4639), .A2(n4395), .ZN(n4394) );
  NOR2_X1 U5308 ( .A1(n4643), .A2(n4640), .ZN(n4639) );
  NAND2_X1 U5309 ( .A1(n4396), .A2(n4632), .ZN(n4395) );
  INV_X1 U5310 ( .A(n5230), .ZN(n4640) );
  NOR2_X1 U5311 ( .A1(n5279), .A2(n4645), .ZN(n4644) );
  INV_X1 U5312 ( .A(n5255), .ZN(n4645) );
  INV_X1 U5313 ( .A(n4841), .ZN(n4642) );
  OR2_X1 U5314 ( .A1(n4384), .A2(n5130), .ZN(n4383) );
  NAND2_X1 U5315 ( .A1(n7595), .A2(n4309), .ZN(n4495) );
  INV_X1 U5316 ( .A(n4761), .ZN(n4757) );
  NAND2_X1 U5317 ( .A1(n4500), .A2(n4499), .ZN(n4497) );
  NAND2_X1 U5318 ( .A1(n4280), .A2(n4484), .ZN(n4483) );
  NAND2_X1 U5319 ( .A1(n4486), .A2(n4280), .ZN(n4482) );
  AND2_X1 U5320 ( .A1(n7580), .A2(n4501), .ZN(n4500) );
  NAND2_X1 U5321 ( .A1(n4447), .A2(n4446), .ZN(n7861) );
  AOI21_X1 U5322 ( .B1(n4448), .B2(n4450), .A(n4307), .ZN(n4446) );
  AOI21_X1 U5323 ( .B1(n8085), .B2(n8077), .A(n7687), .ZN(n8065) );
  NAND2_X1 U5324 ( .A1(n8065), .A2(n8064), .ZN(n8063) );
  AND2_X1 U5325 ( .A1(n7849), .A2(n7850), .ZN(n8064) );
  NAND2_X1 U5326 ( .A1(n4274), .A2(n8121), .ZN(n4684) );
  NOR2_X1 U5327 ( .A1(n8092), .A2(n7827), .ZN(n4687) );
  OR2_X1 U5328 ( .A1(n8083), .A2(n8100), .ZN(n7842) );
  NAND2_X1 U5329 ( .A1(n4473), .A2(n8236), .ZN(n4472) );
  INV_X1 U5330 ( .A(n4474), .ZN(n4473) );
  NAND2_X1 U5331 ( .A1(n4726), .A2(n4475), .ZN(n4474) );
  NAND2_X1 U5332 ( .A1(n4726), .A2(n8241), .ZN(n4725) );
  NOR2_X1 U5333 ( .A1(n4681), .A2(n4723), .ZN(n4717) );
  NAND2_X1 U5334 ( .A1(n5993), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n6026) );
  NAND2_X1 U5335 ( .A1(n7168), .A2(n7312), .ZN(n4712) );
  INV_X1 U5336 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n5975) );
  OR2_X1 U5337 ( .A1(n5976), .A2(n5975), .ZN(n5995) );
  NAND2_X1 U5338 ( .A1(n4698), .A2(n6695), .ZN(n6920) );
  NAND3_X1 U5339 ( .A1(n4703), .A2(n5806), .A3(n5805), .ZN(n7725) );
  NOR2_X1 U5340 ( .A1(n8288), .A2(n8372), .ZN(n8272) );
  OAI21_X1 U5341 ( .B1(n7052), .B2(n7744), .A(n7746), .ZN(n9651) );
  INV_X1 U5342 ( .A(SI_15_), .ZN(n9826) );
  INV_X1 U5343 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n4690) );
  NAND2_X1 U5344 ( .A1(n6224), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6247) );
  INV_X1 U5345 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n4445) );
  OR2_X1 U5346 ( .A1(n5939), .A2(P2_IR_REG_9__SCAN_IN), .ZN(n5956) );
  CLKBUF_X1 U5347 ( .A(n5848), .Z(n5849) );
  INV_X1 U5348 ( .A(n4379), .ZN(n4378) );
  OAI21_X1 U5349 ( .B1(n8670), .B2(n8669), .A(n8790), .ZN(n4379) );
  INV_X1 U5350 ( .A(n9176), .ZN(n5697) );
  AND2_X1 U5351 ( .A1(n4538), .A2(n4537), .ZN(n4536) );
  OR2_X1 U5352 ( .A1(n8990), .A2(n9200), .ZN(n8737) );
  INV_X1 U5353 ( .A(n9007), .ZN(n4560) );
  NOR2_X1 U5354 ( .A1(n7238), .A2(n7158), .ZN(n7031) );
  OR2_X1 U5355 ( .A1(n9601), .A2(n7209), .ZN(n8739) );
  OR2_X1 U5356 ( .A1(n8848), .A2(n9590), .ZN(n8686) );
  NOR2_X1 U5357 ( .A1(n9105), .A2(n4529), .ZN(n9070) );
  INV_X1 U5358 ( .A(n4531), .ZN(n4529) );
  OR2_X1 U5359 ( .A1(n8430), .A2(n4534), .ZN(n4533) );
  INV_X1 U5360 ( .A(SI_30_), .ZN(n4610) );
  AOI21_X1 U5361 ( .B1(n4651), .B2(n4653), .A(n4345), .ZN(n4649) );
  AND2_X1 U5362 ( .A1(n4803), .A2(n4909), .ZN(n4526) );
  NAND2_X1 U5363 ( .A1(n5515), .A2(n5514), .ZN(n5535) );
  OR2_X1 U5364 ( .A1(n5511), .A2(n5510), .ZN(n5515) );
  NOR2_X1 U5365 ( .A1(n5351), .A2(n4623), .ZN(n4622) );
  INV_X1 U5366 ( .A(n5327), .ZN(n4623) );
  AOI21_X1 U5367 ( .B1(n4835), .B2(n4636), .A(n4635), .ZN(n4634) );
  INV_X1 U5368 ( .A(n5178), .ZN(n4635) );
  INV_X1 U5369 ( .A(n5151), .ZN(n4636) );
  NAND2_X1 U5370 ( .A1(n4382), .A2(n4380), .ZN(n5150) );
  INV_X1 U5371 ( .A(n4381), .ZN(n4380) );
  OR2_X1 U5372 ( .A1(n5082), .A2(n4383), .ZN(n4382) );
  OAI21_X1 U5373 ( .B1(n4383), .B2(n4624), .A(n5132), .ZN(n4381) );
  AND2_X1 U5374 ( .A1(n4300), .A2(n6709), .ZN(n4492) );
  NOR2_X1 U5375 ( .A1(n7547), .A2(n4747), .ZN(n4746) );
  INV_X1 U5376 ( .A(n6004), .ZN(n4747) );
  NAND2_X1 U5377 ( .A1(n7338), .A2(n7339), .ZN(n4748) );
  INV_X1 U5378 ( .A(n6302), .ZN(n4504) );
  NOR2_X1 U5379 ( .A1(n7615), .A2(n6096), .ZN(n4488) );
  OR2_X1 U5380 ( .A1(n6953), .A2(n5926), .ZN(n4764) );
  NAND2_X1 U5381 ( .A1(n4524), .A2(n6900), .ZN(n6506) );
  NAND2_X1 U5382 ( .A1(n6111), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n6122) );
  OR2_X1 U5383 ( .A1(n5946), .A2(n5945), .ZN(n5961) );
  OR2_X1 U5384 ( .A1(n7601), .A2(n4762), .ZN(n4761) );
  INV_X1 U5385 ( .A(n4759), .ZN(n4758) );
  OAI21_X1 U5386 ( .B1(n7601), .B2(n4760), .A(n6069), .ZN(n4759) );
  OR2_X1 U5387 ( .A1(n4762), .A2(n7594), .ZN(n4760) );
  NAND2_X1 U5388 ( .A1(n7593), .A2(n7595), .ZN(n6045) );
  NAND2_X1 U5389 ( .A1(n4740), .A2(n4741), .ZN(n7593) );
  NAND2_X1 U5390 ( .A1(n7897), .A2(n6250), .ZN(n4613) );
  NAND2_X1 U5391 ( .A1(n6507), .A2(n9677), .ZN(n7864) );
  INV_X1 U5392 ( .A(n8063), .ZN(n4509) );
  NAND2_X1 U5393 ( .A1(n8298), .A2(n4654), .ZN(n7856) );
  INV_X1 U5394 ( .A(n5839), .ZN(n5853) );
  INV_X1 U5395 ( .A(n6185), .ZN(n6262) );
  NAND2_X1 U5396 ( .A1(n6329), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n5828) );
  OR2_X1 U5397 ( .A1(n6431), .A2(n4404), .ZN(n7935) );
  NOR2_X1 U5398 ( .A1(n6432), .A2(n6914), .ZN(n4404) );
  NAND2_X1 U5399 ( .A1(n6521), .A2(n4337), .ZN(n7950) );
  NAND2_X1 U5400 ( .A1(n7950), .A2(n7949), .ZN(n7948) );
  NAND2_X1 U5401 ( .A1(n4400), .A2(n6742), .ZN(n6746) );
  NAND2_X1 U5402 ( .A1(n6741), .A2(n6740), .ZN(n4400) );
  OR2_X1 U5403 ( .A1(n6986), .A2(n6985), .ZN(n6987) );
  NOR2_X1 U5404 ( .A1(n8008), .A2(n8024), .ZN(n8021) );
  NOR2_X1 U5405 ( .A1(n8309), .A2(n8314), .ZN(n4469) );
  OAI21_X1 U5406 ( .B1(n8064), .B2(n8065), .A(n8063), .ZN(n4695) );
  INV_X1 U5407 ( .A(n8077), .ZN(n8084) );
  AND2_X1 U5408 ( .A1(n7842), .A2(n7838), .ZN(n8077) );
  NAND2_X1 U5409 ( .A1(n4729), .A2(n4728), .ZN(n8078) );
  AOI21_X1 U5410 ( .B1(n4730), .B2(n4734), .A(n4315), .ZN(n4728) );
  NOR2_X1 U5411 ( .A1(n8325), .A2(n4462), .ZN(n4460) );
  NAND2_X1 U5412 ( .A1(n8168), .A2(n4463), .ZN(n8156) );
  INV_X1 U5413 ( .A(n7818), .ZN(n8162) );
  AND2_X1 U5414 ( .A1(n7818), .A2(n7820), .ZN(n4507) );
  NAND2_X1 U5415 ( .A1(n8168), .A2(n8175), .ZN(n8169) );
  AND2_X1 U5416 ( .A1(n7820), .A2(n7816), .ZN(n8176) );
  AND2_X1 U5417 ( .A1(n7810), .A2(n8177), .ZN(n8193) );
  INV_X1 U5418 ( .A(n6086), .ZN(n6084) );
  NAND2_X1 U5419 ( .A1(n4286), .A2(n7792), .ZN(n4675) );
  NOR2_X1 U5420 ( .A1(n8288), .A2(n4474), .ZN(n8255) );
  NAND2_X1 U5421 ( .A1(n4716), .A2(n4718), .ZN(n8231) );
  INV_X1 U5422 ( .A(n4719), .ZN(n4718) );
  NAND2_X1 U5423 ( .A1(n8279), .A2(n4717), .ZN(n4716) );
  OAI21_X1 U5424 ( .B1(n4720), .B2(n4681), .A(n4725), .ZN(n4719) );
  OR3_X1 U5425 ( .A1(n6026), .A2(n6025), .A3(n6024), .ZN(n6039) );
  NAND2_X1 U5426 ( .A1(n4679), .A2(n7786), .ZN(n8265) );
  NAND2_X1 U5427 ( .A1(n4516), .A2(n4513), .ZN(n8281) );
  NAND2_X1 U5428 ( .A1(n4515), .A2(n4514), .ZN(n4513) );
  INV_X1 U5429 ( .A(n4521), .ZN(n4515) );
  NAND2_X1 U5430 ( .A1(n4465), .A2(n4464), .ZN(n7393) );
  AND2_X1 U5431 ( .A1(n7075), .A2(n7878), .ZN(n7169) );
  NAND2_X1 U5432 ( .A1(n4705), .A2(n4706), .ZN(n7041) );
  AOI21_X1 U5433 ( .B1(n4313), .B2(n7017), .A(n4707), .ZN(n4706) );
  AND2_X1 U5434 ( .A1(n4708), .A2(n7008), .ZN(n4707) );
  NAND2_X1 U5435 ( .A1(n6364), .A2(n7698), .ZN(n5911) );
  AOI21_X1 U5436 ( .B1(n9668), .B2(n9673), .A(n9674), .ZN(n6779) );
  NAND2_X1 U5437 ( .A1(n7868), .A2(n6502), .ZN(n6554) );
  NAND2_X1 U5438 ( .A1(n6093), .A2(n6092), .ZN(n8358) );
  AOI22_X1 U5439 ( .A1(n7702), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n5807), .B2(
        n6322), .ZN(n6092) );
  OR2_X1 U5440 ( .A1(n9677), .A2(n7862), .ZN(n9728) );
  INV_X1 U5441 ( .A(n6701), .ZN(n6778) );
  NOR2_X1 U5442 ( .A1(P2_IR_REG_27__SCAN_IN), .A2(P2_IR_REG_28__SCAN_IN), .ZN(
        n4709) );
  NAND2_X1 U5443 ( .A1(n5797), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5798) );
  NAND2_X1 U5444 ( .A1(n5786), .A2(n6005), .ZN(n6219) );
  NAND2_X1 U5445 ( .A1(n6247), .A2(n6246), .ZN(n6245) );
  INV_X1 U5446 ( .A(n5781), .ZN(n4774) );
  NAND2_X1 U5447 ( .A1(n6005), .A2(n5783), .ZN(n6016) );
  NOR2_X1 U5448 ( .A1(n5360), .A2(n5359), .ZN(n5384) );
  AND2_X1 U5449 ( .A1(n5384), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n5409) );
  INV_X1 U5450 ( .A(n5345), .ZN(n4796) );
  AND2_X1 U5451 ( .A1(n4777), .A2(n5425), .ZN(n4776) );
  INV_X1 U5452 ( .A(n8491), .ZN(n4811) );
  INV_X1 U5453 ( .A(n4790), .ZN(n4789) );
  NAND2_X1 U5454 ( .A1(n5312), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n5332) );
  NAND2_X1 U5455 ( .A1(n5467), .A2(n5466), .ZN(n8507) );
  NOR2_X1 U5456 ( .A1(n5639), .A2(n5741), .ZN(n8523) );
  NAND2_X1 U5457 ( .A1(n5035), .A2(n5034), .ZN(n4792) );
  INV_X1 U5458 ( .A(n5036), .ZN(n5034) );
  NOR2_X1 U5459 ( .A1(n5264), .A2(n8425), .ZN(n5289) );
  NOR2_X1 U5460 ( .A1(n4825), .A2(n4822), .ZN(n4819) );
  AOI21_X1 U5461 ( .B1(n4825), .B2(n4818), .A(n4820), .ZN(n4817) );
  INV_X1 U5462 ( .A(n4827), .ZN(n4818) );
  NAND2_X1 U5463 ( .A1(n8421), .A2(n4832), .ZN(n4419) );
  NAND2_X1 U5464 ( .A1(n4816), .A2(n4825), .ZN(n4832) );
  INV_X1 U5465 ( .A(n4374), .ZN(n4373) );
  NAND2_X1 U5466 ( .A1(n8681), .A2(n9074), .ZN(n4372) );
  NOR2_X1 U5467 ( .A1(n9486), .A2(n9485), .ZN(n9484) );
  OR2_X1 U5468 ( .A1(n6569), .A2(n4360), .ZN(n6595) );
  NOR2_X1 U5469 ( .A1(n6420), .A2(n5041), .ZN(n4360) );
  AND2_X1 U5470 ( .A1(n6403), .A2(n6402), .ZN(n6486) );
  AOI21_X1 U5471 ( .B1(n6487), .B2(P1_REG2_REG_10__SCAN_IN), .A(n6486), .ZN(
        n6489) );
  AND2_X1 U5472 ( .A1(n8882), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n4358) );
  AND2_X1 U5473 ( .A1(n8898), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n4357) );
  INV_X1 U5474 ( .A(n4597), .ZN(n4595) );
  AOI21_X1 U5475 ( .B1(n4597), .B2(n8964), .A(n4846), .ZN(n4594) );
  OR2_X1 U5476 ( .A1(n9186), .A2(n5697), .ZN(n8937) );
  NAND2_X1 U5477 ( .A1(n9008), .A2(n4536), .ZN(n8957) );
  NAND2_X1 U5478 ( .A1(n9008), .A2(n4538), .ZN(n8971) );
  AND2_X1 U5479 ( .A1(n8736), .A2(n8779), .ZN(n8979) );
  NAND2_X1 U5480 ( .A1(n9008), .A2(n9299), .ZN(n8987) );
  AOI21_X1 U5481 ( .B1(n4603), .B2(n4324), .A(n4285), .ZN(n4601) );
  NOR2_X1 U5482 ( .A1(n9042), .A2(n9210), .ZN(n9026) );
  NOR2_X1 U5483 ( .A1(n5478), .A2(n8436), .ZN(n5493) );
  OR2_X1 U5484 ( .A1(n5458), .A2(n8513), .ZN(n5478) );
  NAND2_X1 U5485 ( .A1(n9050), .A2(n5730), .ZN(n9036) );
  AOI21_X1 U5486 ( .B1(n4579), .B2(n4576), .A(n4336), .ZN(n4575) );
  INV_X1 U5487 ( .A(n4565), .ZN(n4564) );
  AOI21_X1 U5488 ( .B1(n4565), .B2(n4563), .A(n4562), .ZN(n4561) );
  AND2_X1 U5489 ( .A1(n4566), .A2(n9082), .ZN(n4565) );
  AND2_X1 U5490 ( .A1(n8597), .A2(n8600), .ZN(n9125) );
  OR2_X1 U5491 ( .A1(n5243), .A2(n5242), .ZN(n5264) );
  NAND2_X1 U5492 ( .A1(n7441), .A2(n8594), .ZN(n9398) );
  NOR2_X1 U5493 ( .A1(n9397), .A2(n4570), .ZN(n4569) );
  INV_X1 U5494 ( .A(n8594), .ZN(n4570) );
  NOR2_X1 U5495 ( .A1(n9425), .A2(n4534), .ZN(n9408) );
  OR2_X1 U5496 ( .A1(n5164), .A2(n5163), .ZN(n5185) );
  INV_X1 U5497 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n5184) );
  NOR2_X1 U5498 ( .A1(n5185), .A2(n5184), .ZN(n5213) );
  INV_X1 U5499 ( .A(n9548), .ZN(n9414) );
  NAND2_X1 U5500 ( .A1(n4548), .A2(n8702), .ZN(n4551) );
  INV_X1 U5501 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n5121) );
  OR2_X1 U5502 ( .A1(n5122), .A2(n5121), .ZN(n5164) );
  AND2_X1 U5503 ( .A1(n8702), .A2(n8701), .ZN(n9556) );
  AND2_X1 U5504 ( .A1(n7031), .A2(n7423), .ZN(n9560) );
  NAND2_X1 U5505 ( .A1(n4552), .A2(n8740), .ZN(n9545) );
  INV_X1 U5506 ( .A(n7347), .ZN(n4552) );
  AND2_X1 U5507 ( .A1(n5720), .A2(n8692), .ZN(n8813) );
  NAND2_X1 U5508 ( .A1(n7215), .A2(n9596), .ZN(n7237) );
  NAND2_X1 U5509 ( .A1(n4527), .A2(n4268), .ZN(n7238) );
  INV_X1 U5510 ( .A(n7237), .ZN(n4527) );
  AND3_X1 U5511 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n5040) );
  NOR2_X1 U5512 ( .A1(n7513), .A2(n7196), .ZN(n7215) );
  OR2_X1 U5513 ( .A1(n7089), .A2(n8797), .ZN(n9158) );
  INV_X1 U5514 ( .A(n9158), .ZN(n9559) );
  MUX2_X1 U5515 ( .A(n6352), .B(n9345), .S(n6346), .Z(n7100) );
  NAND2_X1 U5516 ( .A1(n8562), .A2(n8561), .ZN(n8916) );
  NAND2_X1 U5517 ( .A1(n9418), .A2(n5669), .ZN(n7444) );
  OR2_X1 U5518 ( .A1(n8680), .A2(n5741), .ZN(n9440) );
  INV_X1 U5519 ( .A(n9612), .ZN(n9452) );
  INV_X1 U5520 ( .A(n9440), .ZN(n9600) );
  INV_X1 U5521 ( .A(n9615), .ZN(n9273) );
  OR2_X1 U5522 ( .A1(n7088), .A2(n5751), .ZN(n5756) );
  OAI22_X1 U5523 ( .A1(n9576), .A2(P1_D_REG_0__SCAN_IN), .B1(n5601), .B2(n5616), .ZN(n7181) );
  XNOR2_X1 U5524 ( .A(n4609), .B(n7700), .ZN(n8405) );
  OAI21_X1 U5525 ( .B1(n7694), .B2(n4610), .A(n7697), .ZN(n4609) );
  INV_X1 U5526 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n4860) );
  NAND2_X1 U5527 ( .A1(n9329), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4861) );
  XNOR2_X1 U5528 ( .A(n5702), .B(n5701), .ZN(n7527) );
  NAND2_X1 U5529 ( .A1(n4650), .A2(n5582), .ZN(n5702) );
  XNOR2_X1 U5530 ( .A(n5581), .B(n5580), .ZN(n8412) );
  OR2_X1 U5531 ( .A1(n4882), .A2(n9330), .ZN(n4885) );
  INV_X1 U5532 ( .A(n4804), .ZN(n4802) );
  NAND2_X1 U5533 ( .A1(n4885), .A2(n4883), .ZN(n4887) );
  INV_X1 U5534 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n4883) );
  NAND2_X1 U5535 ( .A1(n5451), .A2(n5450), .ZN(n5469) );
  NAND2_X1 U5536 ( .A1(n5328), .A2(n5327), .ZN(n5352) );
  NAND2_X1 U5537 ( .A1(n4646), .A2(n5255), .ZN(n5280) );
  NAND2_X1 U5538 ( .A1(n5254), .A2(n4841), .ZN(n4646) );
  NAND2_X1 U5539 ( .A1(n4851), .A2(n5048), .ZN(n5209) );
  NAND2_X1 U5540 ( .A1(n4399), .A2(n4630), .ZN(n5229) );
  CLKBUF_X1 U5541 ( .A(n5048), .Z(n5049) );
  NAND2_X1 U5542 ( .A1(n5027), .A2(n5026), .ZN(n5053) );
  XNOR2_X1 U5543 ( .A(n4974), .B(n4951), .ZN(n4972) );
  NAND2_X1 U5544 ( .A1(n4748), .A2(n6004), .ZN(n7546) );
  NAND2_X1 U5545 ( .A1(n6133), .A2(n6132), .ZN(n8334) );
  INV_X1 U5546 ( .A(n8051), .ZN(n8254) );
  NOR2_X1 U5547 ( .A1(n5818), .A2(n4306), .ZN(n6635) );
  NAND2_X1 U5548 ( .A1(n5817), .A2(n5816), .ZN(n6634) );
  NAND2_X1 U5549 ( .A1(n5815), .A2(n6900), .ZN(n5817) );
  INV_X1 U5550 ( .A(n4485), .ZN(n7573) );
  AOI21_X1 U5551 ( .B1(n7564), .B2(n4488), .A(n4487), .ZN(n4485) );
  NAND2_X1 U5552 ( .A1(n6110), .A2(n6109), .ZN(n8346) );
  AOI21_X1 U5553 ( .B1(n4275), .B2(n5954), .A(n4320), .ZN(n4478) );
  NAND2_X1 U5554 ( .A1(n6156), .A2(n6155), .ZN(n7582) );
  NAND2_X1 U5555 ( .A1(n7592), .A2(n6049), .ZN(n7602) );
  INV_X1 U5556 ( .A(n8139), .ZN(n8181) );
  XNOR2_X1 U5557 ( .A(n6152), .B(n6153), .ZN(n7608) );
  AND2_X1 U5558 ( .A1(n5846), .A2(n5845), .ZN(n5847) );
  NAND2_X1 U5559 ( .A1(n6871), .A2(n5927), .ZN(n6952) );
  NAND2_X1 U5560 ( .A1(n6105), .A2(n6104), .ZN(n8351) );
  INV_X1 U5561 ( .A(n7643), .ZN(n7666) );
  INV_X1 U5562 ( .A(n7657), .ZN(n7665) );
  NOR2_X1 U5563 ( .A1(n7655), .A2(n8285), .ZN(n7643) );
  NAND2_X1 U5564 ( .A1(n7063), .A2(n5955), .ZN(n7634) );
  NAND2_X1 U5565 ( .A1(n4480), .A2(n4275), .ZN(n7632) );
  INV_X1 U5566 ( .A(n8210), .ZN(n8240) );
  OAI21_X1 U5567 ( .B1(n6045), .B2(n4761), .A(n4758), .ZN(n7642) );
  NAND2_X1 U5568 ( .A1(n6073), .A2(n6072), .ZN(n8361) );
  INV_X1 U5569 ( .A(n7650), .ZN(n4752) );
  NAND2_X1 U5570 ( .A1(n6259), .A2(n6252), .ZN(n7673) );
  NAND2_X1 U5571 ( .A1(n4741), .A2(n7595), .ZN(n7662) );
  NOR2_X1 U5572 ( .A1(n7655), .A2(n8284), .ZN(n7669) );
  INV_X1 U5573 ( .A(n7660), .ZN(n7670) );
  NAND2_X1 U5574 ( .A1(n9353), .A2(n9354), .ZN(n9352) );
  NOR2_X1 U5575 ( .A1(n4405), .A2(n4295), .ZN(n6367) );
  INV_X1 U5576 ( .A(n7920), .ZN(n4405) );
  NOR2_X1 U5577 ( .A1(n6367), .A2(n6366), .ZN(n6431) );
  AND2_X1 U5578 ( .A1(n5914), .A2(n5939), .ZN(n7953) );
  AND2_X1 U5579 ( .A1(n4402), .A2(n4401), .ZN(n6741) );
  NAND2_X1 U5580 ( .A1(n6658), .A2(n6527), .ZN(n4401) );
  NOR2_X1 U5581 ( .A1(n8009), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n8022) );
  OR2_X1 U5582 ( .A1(n4403), .A2(n8021), .ZN(n8009) );
  AND2_X1 U5583 ( .A1(n8008), .A2(n8024), .ZN(n4403) );
  OAI211_X1 U5584 ( .C1(n8034), .C2(n8033), .A(n9628), .B(n8032), .ZN(n4413)
         );
  NAND2_X1 U5585 ( .A1(n4412), .A2(n4411), .ZN(n4410) );
  INV_X1 U5586 ( .A(n8035), .ZN(n4411) );
  NAND2_X1 U5587 ( .A1(n9633), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n4412) );
  AND2_X1 U5588 ( .A1(n7676), .A2(n7675), .ZN(n8304) );
  NAND2_X1 U5589 ( .A1(n8107), .A2(n7832), .ZN(n8099) );
  NAND2_X1 U5590 ( .A1(n4731), .A2(n4732), .ZN(n8093) );
  OR2_X1 U5591 ( .A1(n8134), .A2(n4734), .ZN(n4731) );
  AND2_X1 U5592 ( .A1(n6202), .A2(n6172), .ZN(n8115) );
  NAND2_X1 U5593 ( .A1(n4685), .A2(n7828), .ZN(n8109) );
  NAND2_X1 U5594 ( .A1(n4735), .A2(n4737), .ZN(n8106) );
  NAND2_X1 U5595 ( .A1(n8134), .A2(n8121), .ZN(n4735) );
  NAND2_X1 U5596 ( .A1(n8249), .A2(n8248), .ZN(n8247) );
  NAND2_X1 U5597 ( .A1(n4721), .A2(n4720), .ZN(n8249) );
  AND2_X1 U5598 ( .A1(n4724), .A2(n4297), .ZN(n8264) );
  NAND2_X1 U5599 ( .A1(n8279), .A2(n8280), .ZN(n4724) );
  AND2_X1 U5600 ( .A1(n4523), .A2(n7776), .ZN(n7682) );
  NAND2_X1 U5601 ( .A1(n5992), .A2(n5991), .ZN(n8378) );
  NAND2_X1 U5602 ( .A1(n4666), .A2(n7771), .ZN(n7389) );
  NAND2_X1 U5603 ( .A1(n4667), .A2(n4668), .ZN(n7388) );
  NAND2_X1 U5604 ( .A1(n7313), .A2(n4715), .ZN(n4836) );
  NAND2_X1 U5605 ( .A1(n9639), .A2(n7046), .ZN(n7048) );
  INV_X1 U5606 ( .A(n8290), .ZN(n9647) );
  NAND2_X1 U5607 ( .A1(n6982), .A2(n6981), .ZN(n7009) );
  NOR2_X1 U5608 ( .A1(n8278), .A2(n5807), .ZN(n8257) );
  INV_X1 U5609 ( .A(n7000), .ZN(n8293) );
  AND2_X2 U5610 ( .A1(n6702), .A2(n6701), .ZN(n9752) );
  OAI21_X1 U5611 ( .B1(n8308), .B2(n9678), .A(n4354), .ZN(n8390) );
  NOR2_X1 U5612 ( .A1(n4311), .A2(n4355), .ZN(n4354) );
  INV_X1 U5613 ( .A(n8307), .ZN(n4355) );
  INV_X1 U5614 ( .A(n9670), .ZN(n9926) );
  INV_X1 U5615 ( .A(n5804), .ZN(n7531) );
  NAND2_X1 U5616 ( .A1(n6217), .A2(n6218), .ZN(n8419) );
  INV_X1 U5617 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n9829) );
  XNOR2_X1 U5618 ( .A(n6226), .B(n6225), .ZN(n7405) );
  NAND2_X1 U5619 ( .A1(n6245), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6226) );
  INV_X1 U5620 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7163) );
  INV_X1 U5621 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5776) );
  INV_X1 U5622 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7022) );
  INV_X1 U5623 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n6839) );
  INV_X1 U5624 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n6812) );
  INV_X1 U5625 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n6775) );
  INV_X1 U5626 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n9885) );
  INV_X1 U5627 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6550) );
  INV_X1 U5628 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6339) );
  INV_X1 U5629 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n9814) );
  INV_X1 U5630 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6328) );
  INV_X1 U5631 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6318) );
  INV_X1 U5632 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6310) );
  INV_X1 U5633 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6306) );
  INV_X1 U5634 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6297) );
  INV_X1 U5635 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6294) );
  XNOR2_X1 U5636 ( .A(n5794), .B(P2_IR_REG_1__SCAN_IN), .ZN(n9351) );
  NAND2_X1 U5637 ( .A1(n4829), .A2(n4827), .ZN(n8422) );
  NAND2_X1 U5638 ( .A1(n4831), .A2(n4830), .ZN(n4829) );
  NAND2_X1 U5639 ( .A1(n7377), .A2(n7378), .ZN(n4783) );
  NAND2_X1 U5640 ( .A1(n5161), .A2(n5160), .ZN(n9373) );
  CLKBUF_X1 U5641 ( .A(n8450), .Z(n8451) );
  NAND2_X1 U5642 ( .A1(n5430), .A2(n5429), .ZN(n8456) );
  NAND2_X1 U5643 ( .A1(n4813), .A2(n8433), .ZN(n8490) );
  NAND2_X1 U5644 ( .A1(n5395), .A2(n5394), .ZN(n4780) );
  INV_X1 U5645 ( .A(n8443), .ZN(n5395) );
  AND2_X1 U5646 ( .A1(n4421), .A2(n4781), .ZN(n4420) );
  INV_X1 U5647 ( .A(n7455), .ZN(n4421) );
  INV_X1 U5648 ( .A(n7411), .ZN(n8548) );
  INV_X1 U5649 ( .A(n8545), .ZN(n8534) );
  NAND2_X2 U5650 ( .A1(n4956), .A2(n4955), .ZN(n7186) );
  AND2_X1 U5651 ( .A1(n4954), .A2(n4843), .ZN(n4956) );
  NAND2_X1 U5652 ( .A1(n5346), .A2(n5345), .ZN(n4801) );
  AND2_X1 U5653 ( .A1(n5635), .A2(n5622), .ZN(n8475) );
  AOI21_X1 U5654 ( .B1(n8459), .B2(n4808), .A(n4338), .ZN(n4807) );
  INV_X1 U5655 ( .A(n4812), .ZN(n4808) );
  NAND2_X1 U5656 ( .A1(n5541), .A2(n5540), .ZN(n8973) );
  NAND2_X1 U5657 ( .A1(n6287), .A2(n5619), .ZN(n8556) );
  OR3_X1 U5658 ( .A1(n5437), .A2(n5436), .A3(n5435), .ZN(n9038) );
  OR2_X1 U5659 ( .A1(n4992), .A2(n4941), .ZN(n4943) );
  OR2_X1 U5660 ( .A1(n4989), .A2(n4940), .ZN(n4945) );
  OR2_X1 U5661 ( .A1(n4991), .A2(n9566), .ZN(n4870) );
  NOR2_X1 U5662 ( .A1(n7284), .A2(n7285), .ZN(n7288) );
  NAND2_X1 U5663 ( .A1(n6400), .A2(n6383), .ZN(n9533) );
  AND2_X1 U5664 ( .A1(n4596), .A2(n4597), .ZN(n8935) );
  NAND2_X1 U5665 ( .A1(n9020), .A2(n8734), .ZN(n9005) );
  INV_X1 U5666 ( .A(n5731), .ZN(n9210) );
  NAND2_X1 U5667 ( .A1(n4600), .A2(n5690), .ZN(n9019) );
  OR2_X1 U5668 ( .A1(n9032), .A2(n4324), .ZN(n4600) );
  OAI21_X1 U5669 ( .B1(n9099), .B2(n4581), .A(n4579), .ZN(n9065) );
  NAND2_X1 U5670 ( .A1(n9095), .A2(n8623), .ZN(n9080) );
  NAND2_X1 U5671 ( .A1(n9099), .A2(n9098), .ZN(n4584) );
  NAND2_X1 U5672 ( .A1(n5383), .A2(n5382), .ZN(n9231) );
  NAND2_X1 U5673 ( .A1(n5358), .A2(n5357), .ZN(n9241) );
  NAND2_X1 U5674 ( .A1(n4369), .A2(n5330), .ZN(n9126) );
  NAND2_X1 U5675 ( .A1(n4539), .A2(n4540), .ZN(n9130) );
  NAND2_X1 U5676 ( .A1(n5311), .A2(n5310), .ZN(n9254) );
  NAND2_X1 U5677 ( .A1(n5288), .A2(n5287), .ZN(n9264) );
  NAND2_X1 U5678 ( .A1(n7467), .A2(n8612), .ZN(n9147) );
  NAND2_X1 U5679 ( .A1(n5725), .A2(n8606), .ZN(n7440) );
  NAND2_X1 U5680 ( .A1(n5182), .A2(n5181), .ZN(n9451) );
  NAND2_X1 U5681 ( .A1(n7025), .A2(n4607), .ZN(n7348) );
  NAND2_X1 U5682 ( .A1(n6878), .A2(n5660), .ZN(n7227) );
  INV_X1 U5683 ( .A(n9162), .ZN(n9562) );
  INV_X1 U5684 ( .A(n9060), .ZN(n9554) );
  OR2_X1 U5685 ( .A1(n5756), .A2(n7181), .ZN(n9625) );
  INV_X1 U5686 ( .A(n8916), .ZN(n9287) );
  NAND2_X1 U5687 ( .A1(n8922), .A2(n4349), .ZN(n5748) );
  AND2_X1 U5688 ( .A1(n8924), .A2(n4350), .ZN(n4349) );
  NAND2_X1 U5689 ( .A1(n8965), .A2(n9603), .ZN(n4350) );
  INV_X1 U5690 ( .A(n8456), .ZN(n9305) );
  INV_X1 U5691 ( .A(n9578), .ZN(n9579) );
  INV_X1 U5692 ( .A(n8556), .ZN(n9577) );
  INV_X1 U5693 ( .A(n7181), .ZN(n9328) );
  BUF_X1 U5694 ( .A(n4867), .Z(n7535) );
  CLKBUF_X1 U5695 ( .A(n5636), .Z(n5637) );
  CLKBUF_X1 U5696 ( .A(n5742), .Z(n9337) );
  XNOR2_X1 U5697 ( .A(n4891), .B(n4890), .ZN(n7402) );
  INV_X1 U5698 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7311) );
  NAND2_X1 U5699 ( .A1(n4893), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4895) );
  INV_X1 U5700 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7249) );
  INV_X1 U5701 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7152) );
  XNOR2_X1 U5702 ( .A(n4880), .B(n4881), .ZN(n7151) );
  INV_X1 U5703 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7024) );
  INV_X1 U5704 ( .A(n4839), .ZN(n4428) );
  INV_X1 U5705 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n9903) );
  INV_X1 U5706 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n6552) );
  INV_X1 U5707 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n9828) );
  INV_X1 U5708 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n6316) );
  NAND2_X1 U5709 ( .A1(n4385), .A2(n4626), .ZN(n5131) );
  NAND2_X1 U5710 ( .A1(n5082), .A2(n4624), .ZN(n4385) );
  XNOR2_X1 U5711 ( .A(n4568), .B(n5103), .ZN(n6312) );
  NAND2_X1 U5712 ( .A1(n4629), .A2(n5085), .ZN(n4568) );
  INV_X1 U5713 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6313) );
  INV_X1 U5714 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6308) );
  INV_X1 U5715 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6299) );
  INV_X1 U5716 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6296) );
  XNOR2_X1 U5717 ( .A(n4970), .B(n4969), .ZN(n8850) );
  XNOR2_X1 U5718 ( .A(n4924), .B(n4923), .ZN(n6582) );
  NOR2_X1 U5719 ( .A1(n7275), .A2(n9939), .ZN(n9780) );
  AOI21_X1 U5720 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n9778), .ZN(n9777) );
  NOR2_X1 U5721 ( .A1(n9777), .A2(n9776), .ZN(n9775) );
  AOI21_X1 U5722 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n9775), .ZN(n9774) );
  OAI21_X1 U5723 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n9772), .ZN(n9770) );
  AOI21_X1 U5724 ( .B1(n7900), .B2(n7899), .A(n4525), .ZN(n7905) );
  INV_X1 U5725 ( .A(n4407), .ZN(n6438) );
  INV_X1 U5726 ( .A(n4402), .ZN(n6657) );
  NAND2_X1 U5727 ( .A1(n4414), .A2(n4409), .ZN(P2_U3264) );
  NAND2_X1 U5728 ( .A1(n4415), .A2(n7895), .ZN(n4414) );
  AOI21_X1 U5729 ( .B1(n4413), .B2(n5807), .A(n4410), .ZN(n4409) );
  OAI22_X1 U5730 ( .A1(n8030), .A2(n8029), .B1(n8031), .B2(n9629), .ZN(n4415)
         );
  INV_X1 U5731 ( .A(n8298), .ZN(n8040) );
  NOR2_X1 U5732 ( .A1(n6341), .A2(P1_U3084), .ZN(P1_U4006) );
  CLKBUF_X1 U5733 ( .A(n6931), .Z(n6932) );
  XNOR2_X1 U5734 ( .A(n4423), .B(n4422), .ZN(n8464) );
  MUX2_X1 U5735 ( .A(n9168), .B(n9281), .S(n4270), .Z(n9169) );
  MUX2_X1 U5736 ( .A(n9282), .B(n9281), .S(n9619), .Z(n9283) );
  INV_X1 U5737 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n7280) );
  AND2_X1 U5738 ( .A1(n4688), .A2(n7828), .ZN(n4274) );
  INV_X1 U5739 ( .A(n4992), .ZN(n5162) );
  AND2_X1 U5740 ( .A1(n8612), .A2(n4543), .ZN(n4276) );
  OR2_X1 U5741 ( .A1(n5938), .A2(n5937), .ZN(n4277) );
  OAI21_X1 U5742 ( .B1(n4758), .B2(n4756), .A(n4314), .ZN(n4755) );
  NAND2_X1 U5743 ( .A1(n8430), .A2(n9266), .ZN(n4278) );
  AND2_X1 U5744 ( .A1(n5783), .A2(n4445), .ZN(n4279) );
  INV_X1 U5745 ( .A(n9098), .ZN(n4580) );
  OR2_X1 U5746 ( .A1(n6119), .A2(n6118), .ZN(n4280) );
  XNOR2_X1 U5747 ( .A(n4861), .B(n4860), .ZN(n4866) );
  INV_X1 U5748 ( .A(n8280), .ZN(n4680) );
  NAND4_X2 U5749 ( .A1(n5830), .A2(n5829), .A3(n5828), .A4(n5827), .ZN(n7917)
         );
  INV_X1 U5750 ( .A(n7917), .ZN(n4362) );
  AND2_X1 U5751 ( .A1(n9547), .A2(n7352), .ZN(n4281) );
  NAND2_X1 U5752 ( .A1(n6008), .A2(n6007), .ZN(n7780) );
  AND2_X1 U5753 ( .A1(n7698), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n4282) );
  NAND2_X1 U5754 ( .A1(n6056), .A2(n6055), .ZN(n8368) );
  INV_X1 U5755 ( .A(n8368), .ZN(n4726) );
  OR2_X1 U5756 ( .A1(n4779), .A2(n8444), .ZN(n4283) );
  AND2_X1 U5757 ( .A1(n4540), .A2(n8767), .ZN(n4284) );
  NAND2_X1 U5758 ( .A1(n6158), .A2(n6157), .ZN(n8325) );
  INV_X1 U5759 ( .A(n8702), .ZN(n4554) );
  INV_X1 U5760 ( .A(n7312), .ZN(n4713) );
  NOR2_X1 U5761 ( .A1(n5731), .A2(n9201), .ZN(n4285) );
  AOI21_X1 U5762 ( .B1(n8121), .B2(n4739), .A(n4316), .ZN(n4737) );
  NAND2_X1 U5763 ( .A1(n4681), .A2(n7790), .ZN(n4286) );
  AND2_X1 U5764 ( .A1(n4536), .A2(n4535), .ZN(n4287) );
  NAND3_X1 U5765 ( .A1(n4811), .A2(n8459), .A3(n4806), .ZN(n4288) );
  XNOR2_X1 U5766 ( .A(n4895), .B(n4894), .ZN(n5620) );
  OR3_X1 U5767 ( .A1(n9425), .A2(n9407), .A3(n4534), .ZN(n4289) );
  OR2_X1 U5768 ( .A1(n9105), .A2(n4530), .ZN(n4290) );
  AND2_X1 U5769 ( .A1(n6182), .A2(n4497), .ZN(n4291) );
  OR2_X1 U5770 ( .A1(n5209), .A2(P1_IR_REG_12__SCAN_IN), .ZN(n4292) );
  INV_X1 U5771 ( .A(n7387), .ZN(n4464) );
  INV_X1 U5772 ( .A(n5820), .ZN(n4502) );
  OR2_X1 U5773 ( .A1(n8113), .A2(n4468), .ZN(n4293) );
  INV_X1 U5774 ( .A(n6783), .ZN(n6032) );
  NAND2_X2 U5775 ( .A1(n6241), .A2(n6258), .ZN(n6783) );
  XNOR2_X1 U5776 ( .A(n5772), .B(n5782), .ZN(n7898) );
  OAI211_X1 U5777 ( .C1(n6346), .C2(n6420), .A(n5059), .B(n5058), .ZN(n7242)
         );
  INV_X1 U5778 ( .A(n6900), .ZN(n9676) );
  AND2_X1 U5779 ( .A1(n9020), .A2(n4558), .ZN(n4294) );
  NAND2_X1 U5780 ( .A1(n5239), .A2(n5238), .ZN(n9407) );
  INV_X1 U5781 ( .A(n7874), .ZN(n9650) );
  AND2_X1 U5782 ( .A1(n6373), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n4295) );
  NAND4_X1 U5783 ( .A1(n5813), .A2(n5812), .A3(n5811), .A4(n5810), .ZN(n7919)
         );
  INV_X1 U5784 ( .A(n7919), .ZN(n4524) );
  NAND2_X1 U5785 ( .A1(n4591), .A2(n5693), .ZN(n8970) );
  NAND2_X1 U5786 ( .A1(n7690), .A2(n7689), .ZN(n8305) );
  OR2_X1 U5787 ( .A1(n8368), .A2(n8241), .ZN(n7792) );
  NAND2_X1 U5788 ( .A1(n4584), .A2(n5685), .ZN(n9081) );
  NAND2_X1 U5789 ( .A1(n4780), .A2(n5398), .ZN(n8497) );
  NOR2_X1 U5790 ( .A1(n8134), .A2(n4739), .ZN(n4296) );
  INV_X1 U5791 ( .A(n7771), .ZN(n4520) );
  NAND2_X1 U5792 ( .A1(n5521), .A2(n5520), .ZN(n8990) );
  NAND2_X1 U5793 ( .A1(n4869), .A2(n4867), .ZN(n4992) );
  NAND2_X1 U5794 ( .A1(n5212), .A2(n5211), .ZN(n9444) );
  INV_X1 U5795 ( .A(n8121), .ZN(n4689) );
  OR2_X1 U5796 ( .A1(n8287), .A2(n8268), .ZN(n4297) );
  NAND2_X1 U5797 ( .A1(n6143), .A2(n6142), .ZN(n8329) );
  INV_X1 U5798 ( .A(n5485), .ZN(n4900) );
  AND2_X1 U5799 ( .A1(n8937), .A2(n8780), .ZN(n8964) );
  AND2_X1 U5800 ( .A1(n6197), .A2(n6196), .ZN(n8083) );
  OR2_X1 U5801 ( .A1(n6681), .A2(n7090), .ZN(n4298) );
  AND2_X1 U5802 ( .A1(n8642), .A2(n8734), .ZN(n9021) );
  INV_X1 U5803 ( .A(n9021), .ZN(n4557) );
  NAND2_X1 U5804 ( .A1(n5408), .A2(n5407), .ZN(n9228) );
  NAND2_X1 U5805 ( .A1(n6121), .A2(n6120), .ZN(n8341) );
  NOR2_X1 U5806 ( .A1(n4800), .A2(n4796), .ZN(n4299) );
  INV_X1 U5807 ( .A(n4582), .ZN(n4581) );
  NOR2_X1 U5808 ( .A1(n5686), .A2(n4583), .ZN(n4582) );
  NAND2_X1 U5809 ( .A1(n5888), .A2(n5887), .ZN(n4300) );
  NAND2_X1 U5810 ( .A1(n8168), .A2(n4461), .ZN(n4301) );
  AND2_X1 U5811 ( .A1(n7047), .A2(n7046), .ZN(n4302) );
  AND2_X1 U5812 ( .A1(n5224), .A2(n5200), .ZN(n4303) );
  AND2_X1 U5813 ( .A1(n5114), .A2(n5094), .ZN(n4304) );
  AND2_X1 U5814 ( .A1(n5176), .A2(n5175), .ZN(n4305) );
  INV_X1 U5815 ( .A(n4755), .ZN(n4754) );
  AND2_X1 U5816 ( .A1(n5809), .A2(n5808), .ZN(n4306) );
  INV_X1 U5817 ( .A(n4632), .ZN(n4631) );
  NAND2_X1 U5818 ( .A1(n4634), .A2(n5201), .ZN(n4632) );
  AND2_X1 U5819 ( .A1(n7893), .A2(n7857), .ZN(n4307) );
  OR2_X1 U5820 ( .A1(n4616), .A2(n7864), .ZN(n4308) );
  AND2_X1 U5821 ( .A1(n4757), .A2(n7641), .ZN(n4309) );
  OR2_X1 U5822 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(P1_IR_REG_25__SCAN_IN), .ZN(
        n4310) );
  NAND2_X1 U5823 ( .A1(n4694), .A2(n4692), .ZN(n4311) );
  INV_X1 U5824 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5787) );
  NOR2_X1 U5825 ( .A1(n9231), .A2(n9242), .ZN(n4312) );
  OR2_X1 U5826 ( .A1(n4708), .A2(n7008), .ZN(n4313) );
  INV_X1 U5827 ( .A(n6981), .ZN(n4708) );
  NAND2_X1 U5828 ( .A1(n6082), .A2(n6083), .ZN(n4314) );
  INV_X1 U5829 ( .A(n4723), .ZN(n4722) );
  NAND2_X1 U5830 ( .A1(n4727), .A2(n8280), .ZN(n4723) );
  INV_X1 U5831 ( .A(n4462), .ZN(n4461) );
  NAND2_X1 U5832 ( .A1(n4463), .A2(n8146), .ZN(n4462) );
  NOR2_X1 U5833 ( .A1(n8314), .A2(n8087), .ZN(n4315) );
  NOR2_X1 U5834 ( .A1(n8325), .A2(n8140), .ZN(n4316) );
  INV_X1 U5835 ( .A(n4512), .ZN(n8237) );
  OR2_X1 U5836 ( .A1(n8239), .A2(n8238), .ZN(n4512) );
  OR2_X1 U5837 ( .A1(n8505), .A2(n5487), .ZN(n4815) );
  AND2_X1 U5838 ( .A1(n5105), .A2(SI_7_), .ZN(n4317) );
  AND2_X1 U5839 ( .A1(n5203), .A2(SI_11_), .ZN(n4318) );
  AND2_X1 U5840 ( .A1(n5278), .A2(SI_14_), .ZN(n4319) );
  AND2_X1 U5841 ( .A1(n5967), .A2(n5969), .ZN(n4320) );
  AND2_X1 U5842 ( .A1(n8304), .A2(n8070), .ZN(n4321) );
  OR2_X1 U5843 ( .A1(n7387), .A2(n7909), .ZN(n4322) );
  OAI21_X1 U5844 ( .B1(n4488), .B2(n4487), .A(n7572), .ZN(n4486) );
  NAND2_X1 U5845 ( .A1(n8266), .A2(n4297), .ZN(n4323) );
  AND2_X1 U5846 ( .A1(n9215), .A2(n9218), .ZN(n4324) );
  OR2_X1 U5847 ( .A1(n8208), .A2(n8207), .ZN(n4325) );
  OR2_X1 U5848 ( .A1(n7008), .A2(n7017), .ZN(n4326) );
  NOR2_X1 U5849 ( .A1(n7852), .A2(n4457), .ZN(n4327) );
  OR2_X1 U5850 ( .A1(n6346), .A2(n6311), .ZN(n4328) );
  INV_X1 U5851 ( .A(n5669), .ZN(n4588) );
  INV_X1 U5852 ( .A(n7824), .ZN(n4443) );
  OR2_X1 U5853 ( .A1(n6181), .A2(n4751), .ZN(n4329) );
  OR2_X1 U5854 ( .A1(n8351), .A2(n8223), .ZN(n7811) );
  AND2_X1 U5855 ( .A1(n4691), .A2(n4690), .ZN(n4330) );
  AND2_X1 U5856 ( .A1(n4684), .A2(n4687), .ZN(n4331) );
  INV_X1 U5857 ( .A(n4559), .ZN(n4558) );
  NAND2_X1 U5858 ( .A1(n4560), .A2(n8734), .ZN(n4559) );
  INV_X1 U5859 ( .A(n4397), .ZN(n4396) );
  NAND2_X1 U5860 ( .A1(n4630), .A2(n4398), .ZN(n4397) );
  INV_X1 U5861 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n4416) );
  CLKBUF_X3 U5862 ( .A(n6050), .Z(n7702) );
  NAND2_X1 U5863 ( .A1(n5584), .A2(n5583), .ZN(n8945) );
  INV_X1 U5864 ( .A(n8945), .ZN(n4535) );
  NAND2_X1 U5865 ( .A1(n5565), .A2(n5564), .ZN(n9186) );
  INV_X1 U5866 ( .A(n9186), .ZN(n4537) );
  INV_X1 U5867 ( .A(n8248), .ZN(n4681) );
  INV_X1 U5868 ( .A(n7907), .ZN(n4522) );
  INV_X1 U5869 ( .A(n8765), .ZN(n4543) );
  XOR2_X1 U5870 ( .A(n5297), .B(n7090), .Z(n4332) );
  INV_X1 U5871 ( .A(n8744), .ZN(n4541) );
  NAND2_X1 U5872 ( .A1(n4593), .A2(n5675), .ZN(n9149) );
  NAND2_X1 U5873 ( .A1(n5300), .A2(n8541), .ZN(n8465) );
  OR2_X1 U5874 ( .A1(n9204), .A2(n8641), .ZN(n4333) );
  INV_X1 U5875 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n9330) );
  NAND2_X1 U5876 ( .A1(n6045), .A2(n7594), .ZN(n7592) );
  AND2_X1 U5877 ( .A1(n4679), .A2(n4677), .ZN(n4334) );
  OAI21_X1 U5878 ( .B1(n7492), .B2(n4819), .A(n4817), .ZN(n8540) );
  OR2_X1 U5879 ( .A1(n4535), .A2(n9326), .ZN(n4335) );
  NOR3_X1 U5880 ( .A1(n9105), .A2(n9215), .A3(n4530), .ZN(n4528) );
  AND2_X1 U5881 ( .A1(n9228), .A2(n9232), .ZN(n4336) );
  INV_X1 U5882 ( .A(n8786), .ZN(n8926) );
  NAND2_X1 U5883 ( .A1(n5707), .A2(n5706), .ZN(n8786) );
  OR2_X1 U5884 ( .A1(n6522), .A2(n6435), .ZN(n4337) );
  AND2_X1 U5885 ( .A1(n5532), .A2(n5531), .ZN(n4338) );
  INV_X1 U5886 ( .A(n4471), .ZN(n8232) );
  NOR2_X1 U5887 ( .A1(n8288), .A2(n4472), .ZN(n4471) );
  OR2_X1 U5888 ( .A1(n5308), .A2(P1_IR_REG_16__SCAN_IN), .ZN(n4339) );
  AND2_X1 U5889 ( .A1(n5376), .A2(SI_18_), .ZN(n4340) );
  INV_X1 U5890 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n4852) );
  INV_X1 U5891 ( .A(n6182), .ZN(n4751) );
  AND2_X1 U5892 ( .A1(n5447), .A2(n5428), .ZN(n4341) );
  AND2_X1 U5893 ( .A1(n7025), .A2(n5664), .ZN(n4342) );
  INV_X1 U5894 ( .A(n8434), .ZN(n4814) );
  AND2_X1 U5895 ( .A1(n4879), .A2(n4893), .ZN(n5621) );
  NAND2_X1 U5896 ( .A1(n4479), .A2(n4478), .ZN(n7303) );
  NAND2_X1 U5897 ( .A1(n4783), .A2(n5149), .ZN(n7406) );
  AND2_X1 U5898 ( .A1(n7757), .A2(n7756), .ZN(n7878) );
  INV_X1 U5899 ( .A(n7878), .ZN(n4672) );
  INV_X1 U5900 ( .A(n8039), .ZN(n4654) );
  NAND2_X1 U5901 ( .A1(n4789), .A2(n4792), .ZN(n8472) );
  NAND2_X1 U5902 ( .A1(n4782), .A2(n4781), .ZN(n7454) );
  NAND2_X1 U5903 ( .A1(n6830), .A2(n6829), .ZN(n6828) );
  OR2_X1 U5904 ( .A1(n6219), .A2(P2_IR_REG_25__SCAN_IN), .ZN(n4343) );
  NOR3_X1 U5905 ( .A1(n9425), .A2(n4533), .A3(n9407), .ZN(n4532) );
  NAND2_X1 U5906 ( .A1(n4788), .A2(n4304), .ZN(n7326) );
  NOR2_X1 U5907 ( .A1(n7319), .A2(n7636), .ZN(n4465) );
  AND2_X1 U5908 ( .A1(n7313), .A2(n7312), .ZN(n4344) );
  AND2_X1 U5909 ( .A1(n5704), .A2(n5703), .ZN(n4345) );
  AND2_X1 U5910 ( .A1(n4753), .A2(n6708), .ZN(n4346) );
  AND2_X1 U5911 ( .A1(n4767), .A2(n6871), .ZN(n4347) );
  INV_X1 U5912 ( .A(n4551), .ZN(n4553) );
  NOR2_X1 U5913 ( .A1(n7089), .A2(n7151), .ZN(n4348) );
  XNOR2_X1 U5914 ( .A(n6223), .B(n6222), .ZN(n6505) );
  NAND2_X1 U5915 ( .A1(n5807), .A2(n6250), .ZN(n6507) );
  NAND2_X1 U5916 ( .A1(n6037), .A2(n6036), .ZN(n8372) );
  INV_X1 U5917 ( .A(n8372), .ZN(n4475) );
  INV_X1 U5918 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n4858) );
  NAND2_X1 U5919 ( .A1(n6968), .A2(n6556), .ZN(n6694) );
  INV_X1 U5920 ( .A(n6694), .ZN(n4466) );
  XNOR2_X1 U5921 ( .A(n5774), .B(P2_IR_REG_19__SCAN_IN), .ZN(n5807) );
  INV_X1 U5922 ( .A(n5807), .ZN(n7895) );
  INV_X1 U5923 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n6051) );
  INV_X1 U5924 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n4894) );
  INV_X1 U5925 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n4664) );
  NAND2_X1 U5926 ( .A1(n8963), .A2(n8964), .ZN(n8936) );
  INV_X1 U5927 ( .A(n7468), .ZN(n4353) );
  OAI21_X1 U5928 ( .B1(n9022), .B2(n4559), .A(n4555), .ZN(n8997) );
  INV_X1 U5929 ( .A(n9052), .ZN(n4352) );
  NAND2_X1 U5930 ( .A1(n5724), .A2(n8741), .ZN(n9412) );
  NAND2_X1 U5931 ( .A1(n9290), .A2(n4335), .ZN(P1_U3519) );
  NAND2_X4 U5932 ( .A1(n4661), .A2(n4662), .ZN(n7698) );
  INV_X1 U5933 ( .A(n8956), .ZN(n5699) );
  INV_X1 U5934 ( .A(n4607), .ZN(n4606) );
  AOI22_X1 U5935 ( .A1(n8078), .A2(n8084), .B1(n8060), .B2(n8083), .ZN(n8062)
         );
  AOI22_X1 U5936 ( .A1(n8167), .A2(n8057), .B1(n8175), .B2(n8056), .ZN(n8163)
         );
  OAI21_X1 U5937 ( .B1(n8228), .B2(n8240), .A(n8053), .ZN(n8201) );
  NAND2_X1 U5938 ( .A1(n7431), .A2(n7430), .ZN(n8049) );
  NAND3_X1 U5939 ( .A1(n4701), .A2(n4699), .A3(n7725), .ZN(n7868) );
  NAND3_X1 U5940 ( .A1(n4505), .A2(n4503), .A3(n5795), .ZN(n4703) );
  NAND2_X1 U5941 ( .A1(n8686), .A2(n6880), .ZN(n7503) );
  NOR2_X2 U5942 ( .A1(n8935), .A2(n8934), .ZN(n9181) );
  NAND2_X1 U5943 ( .A1(n9519), .A2(n9518), .ZN(n9517) );
  XNOR2_X1 U5944 ( .A(n7137), .B(n9513), .ZN(n9519) );
  NOR2_X1 U5945 ( .A1(n9526), .A2(n4357), .ZN(n8895) );
  NOR2_X1 U5946 ( .A1(n8878), .A2(n4358), .ZN(n8880) );
  NOR2_X1 U5947 ( .A1(n6650), .A2(n6651), .ZN(n6764) );
  NOR2_X1 U5948 ( .A1(n6571), .A2(n6570), .ZN(n6569) );
  NOR2_X1 U5949 ( .A1(n6768), .A2(n6767), .ZN(n7135) );
  NOR2_X1 U5950 ( .A1(n6394), .A2(n6593), .ZN(n6461) );
  NAND2_X2 U5952 ( .A1(n8049), .A2(n8048), .ZN(n8279) );
  INV_X1 U5953 ( .A(n8627), .ZN(n4363) );
  INV_X1 U5954 ( .A(n8729), .ZN(n4364) );
  NAND4_X1 U5955 ( .A1(n8622), .A2(n8631), .A3(n8772), .A4(n8674), .ZN(n4365)
         );
  NAND2_X1 U5956 ( .A1(n6826), .A2(n8563), .ZN(n4369) );
  INV_X1 U5957 ( .A(n4626), .ZN(n4384) );
  AND2_X1 U5958 ( .A1(n4387), .A2(n4386), .ZN(n8660) );
  NAND3_X1 U5959 ( .A1(n4393), .A2(n4390), .A3(n4388), .ZN(n4387) );
  OAI21_X1 U5960 ( .B1(n5152), .B2(n4397), .A(n4394), .ZN(n4638) );
  MUX2_X1 U5961 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n4416), .S(n9351), .Z(n9353)
         );
  AND4_X2 U5962 ( .A1(n4847), .A2(n4952), .A3(n4848), .A4(n4787), .ZN(n5048)
         );
  NAND2_X2 U5963 ( .A1(n4419), .A2(n4332), .ZN(n8541) );
  OAI21_X2 U5964 ( .B1(n8443), .B2(n4283), .A(n4776), .ZN(n8450) );
  NAND2_X2 U5965 ( .A1(n4782), .A2(n4420), .ZN(n7456) );
  OAI21_X1 U5966 ( .B1(n5308), .B2(n4429), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n4880) );
  INV_X1 U5967 ( .A(n4425), .ZN(n4876) );
  OR3_X1 U5968 ( .A1(n5308), .A2(n4428), .A3(P1_IR_REG_16__SCAN_IN), .ZN(n4896) );
  MUX2_X1 U5969 ( .A(n7713), .B(n7714), .S(n7857), .Z(n7731) );
  AOI21_X1 U5970 ( .B1(n4442), .B2(n7836), .A(n7835), .ZN(n7844) );
  NAND2_X1 U5971 ( .A1(n4444), .A2(n6005), .ZN(n5770) );
  AND2_X1 U5972 ( .A1(n6005), .A2(n4279), .ZN(n6034) );
  NAND2_X1 U5973 ( .A1(n7848), .A2(n4448), .ZN(n4447) );
  NAND2_X1 U5974 ( .A1(n8168), .A2(n4460), .ZN(n8122) );
  AND2_X1 U5975 ( .A1(n7003), .A2(n9676), .ZN(n6556) );
  OAI21_X2 U5976 ( .B1(P1_RD_REG_SCAN_IN), .B2(P2_ADDR_REG_19__SCAN_IN), .A(
        n4664), .ZN(n4662) );
  NOR2_X1 U5977 ( .A1(n8113), .A2(n8314), .ZN(n8094) );
  NOR2_X1 U5978 ( .A1(n8113), .A2(n4467), .ZN(n8079) );
  INV_X1 U5979 ( .A(n4470), .ZN(n8224) );
  NAND2_X1 U5980 ( .A1(n7555), .A2(n7556), .ZN(n4476) );
  NAND2_X1 U5981 ( .A1(n4477), .A2(n6141), .ZN(n7554) );
  NAND2_X1 U5982 ( .A1(n7622), .A2(n6131), .ZN(n4477) );
  NAND2_X1 U5983 ( .A1(n7065), .A2(n4275), .ZN(n4479) );
  XNOR2_X1 U5984 ( .A(n6130), .B(n6128), .ZN(n7624) );
  OAI21_X2 U5985 ( .B1(n7564), .B2(n4483), .A(n4482), .ZN(n6130) );
  NAND2_X1 U5986 ( .A1(n7564), .A2(n6097), .ZN(n7616) );
  NOR2_X1 U5987 ( .A1(n6108), .A2(n6107), .ZN(n4487) );
  NAND2_X1 U5988 ( .A1(n4491), .A2(n4489), .ZN(n6830) );
  AOI21_X2 U5989 ( .B1(n6721), .B2(n6723), .A(n6722), .ZN(n6710) );
  NAND2_X1 U5990 ( .A1(n4493), .A2(n4494), .ZN(n7566) );
  OR2_X1 U5991 ( .A1(n7582), .A2(n4500), .ZN(n4496) );
  NAND2_X1 U5992 ( .A1(n7582), .A2(n4499), .ZN(n4498) );
  NAND3_X1 U5993 ( .A1(n6364), .A2(n7698), .A3(n4504), .ZN(n4503) );
  NAND2_X2 U5994 ( .A1(n6260), .A2(n8413), .ZN(n6364) );
  INV_X2 U5995 ( .A(n6364), .ZN(n6322) );
  NAND3_X1 U5996 ( .A1(n7528), .A2(n8413), .A3(n9351), .ZN(n4505) );
  AND2_X2 U5997 ( .A1(n5889), .A2(n5768), .ZN(n6005) );
  OAI21_X2 U5998 ( .B1(n9651), .B2(n7874), .A(n7750), .ZN(n7074) );
  AOI21_X2 U5999 ( .B1(n8152), .B2(n7685), .A(n7710), .ZN(n8128) );
  AND2_X2 U6000 ( .A1(n4512), .A2(n4511), .ZN(n8219) );
  NAND2_X1 U6001 ( .A1(n4666), .A2(n4517), .ZN(n4516) );
  NAND2_X1 U6002 ( .A1(n6970), .A2(n6971), .ZN(n7015) );
  OAI21_X1 U6003 ( .B1(n6969), .B2(n7736), .A(n7715), .ZN(n6970) );
  MUX2_X1 U6004 ( .A(n9638), .B(n8420), .S(n6364), .Z(n6900) );
  NAND2_X1 U6005 ( .A1(n4859), .A2(n4526), .ZN(n4905) );
  INV_X2 U6006 ( .A(n5617), .ZN(n4859) );
  INV_X1 U6007 ( .A(n4528), .ZN(n9042) );
  INV_X1 U6008 ( .A(n4532), .ZN(n9159) );
  AND2_X2 U6009 ( .A1(n9008), .A2(n4287), .ZN(n8942) );
  NAND2_X1 U6010 ( .A1(n4976), .A2(n4975), .ZN(n5002) );
  NAND3_X1 U6011 ( .A1(n4546), .A2(n4544), .A3(n5022), .ZN(n5027) );
  NAND2_X1 U6012 ( .A1(n5005), .A2(n4545), .ZN(n4544) );
  INV_X1 U6013 ( .A(n5001), .ZN(n4545) );
  NAND3_X1 U6014 ( .A1(n5005), .A2(n4976), .A3(n4975), .ZN(n4546) );
  NAND2_X1 U6015 ( .A1(n4547), .A2(n5005), .ZN(n5023) );
  NAND2_X1 U6016 ( .A1(n5002), .A2(n5001), .ZN(n4547) );
  OR2_X1 U6017 ( .A1(n8756), .A2(n4554), .ZN(n4550) );
  NAND2_X1 U6018 ( .A1(n8756), .A2(n5722), .ZN(n4548) );
  NAND2_X1 U6019 ( .A1(n4549), .A2(n4553), .ZN(n7359) );
  NAND2_X1 U6020 ( .A1(n7347), .A2(n8756), .ZN(n4549) );
  OAI211_X1 U6021 ( .C1(n4551), .C2(n7347), .A(n8704), .B(n4550), .ZN(n5724)
         );
  OAI21_X1 U6022 ( .B1(n9097), .B2(n4564), .A(n4561), .ZN(n9067) );
  NAND2_X2 U6023 ( .A1(P1_U3084), .A2(n5793), .ZN(n9343) );
  MUX2_X1 U6024 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(P1_DATAO_REG_2__SCAN_IN), 
        .S(n7698), .Z(n4974) );
  MUX2_X1 U6025 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(P1_DATAO_REG_1__SCAN_IN), 
        .S(n7698), .Z(n4946) );
  MUX2_X1 U6026 ( .A(n6301), .B(n6293), .S(n7698), .Z(n5003) );
  MUX2_X1 U6027 ( .A(n6296), .B(n6294), .S(n7698), .Z(n5024) );
  MUX2_X1 U6028 ( .A(n6299), .B(n6297), .S(n7698), .Z(n5054) );
  MUX2_X1 U6029 ( .A(n6308), .B(n6306), .S(n7698), .Z(n5083) );
  MUX2_X1 U6030 ( .A(n6313), .B(n6310), .S(n7698), .Z(n5104) );
  MUX2_X1 U6031 ( .A(n6316), .B(n6318), .S(n7698), .Z(n5107) );
  MUX2_X1 U6032 ( .A(n5133), .B(n6328), .S(n7698), .Z(n5135) );
  MUX2_X1 U6033 ( .A(n6336), .B(n9814), .S(n7698), .Z(n5154) );
  MUX2_X1 U6034 ( .A(n9828), .B(n6339), .S(n7698), .Z(n5202) );
  MUX2_X1 U6035 ( .A(n6552), .B(n6550), .S(n7698), .Z(n5206) );
  MUX2_X1 U6036 ( .A(n9339), .B(n8415), .S(n7698), .Z(n5561) );
  NAND2_X2 U6037 ( .A1(n6346), .A2(n5793), .ZN(n4971) );
  NAND2_X1 U6038 ( .A1(n4982), .A2(n8849), .ZN(n4931) );
  NAND2_X1 U6039 ( .A1(n9099), .A2(n4574), .ZN(n4577) );
  NAND2_X1 U6040 ( .A1(n4585), .A2(n4586), .ZN(n7443) );
  NAND2_X1 U6041 ( .A1(n9415), .A2(n5669), .ZN(n4585) );
  NAND2_X1 U6042 ( .A1(n4591), .A2(n4590), .ZN(n5696) );
  NAND2_X1 U6043 ( .A1(n4593), .A2(n4592), .ZN(n5677) );
  NAND2_X1 U6044 ( .A1(n5699), .A2(n5698), .ZN(n4596) );
  NAND2_X1 U6045 ( .A1(n4596), .A2(n5700), .ZN(n8933) );
  INV_X1 U6046 ( .A(n5700), .ZN(n4598) );
  NAND3_X1 U6047 ( .A1(n6878), .A2(n5661), .A3(n5660), .ZN(n7225) );
  NAND2_X2 U6048 ( .A1(n6879), .A2(n6882), .ZN(n6878) );
  NAND2_X1 U6049 ( .A1(n9032), .A2(n4603), .ZN(n4602) );
  NAND3_X1 U6051 ( .A1(n4857), .A2(n5048), .A3(n4608), .ZN(n5617) );
  NOR2_X2 U6053 ( .A1(n9642), .A2(n7056), .ZN(n9643) );
  NAND2_X1 U6054 ( .A1(n4612), .A2(n4616), .ZN(n4611) );
  NAND2_X1 U6055 ( .A1(n4614), .A2(n4613), .ZN(n4612) );
  NAND2_X1 U6056 ( .A1(n4615), .A2(n4266), .ZN(n4614) );
  XNOR2_X1 U6057 ( .A(n7896), .B(n7895), .ZN(n4615) );
  NAND2_X1 U6058 ( .A1(n5328), .A2(n4618), .ZN(n4617) );
  NAND2_X1 U6059 ( .A1(n4617), .A2(n4619), .ZN(n5400) );
  NAND2_X1 U6060 ( .A1(n5082), .A2(n5081), .ZN(n4629) );
  INV_X1 U6061 ( .A(n5081), .ZN(n4625) );
  NAND2_X1 U6062 ( .A1(n5152), .A2(n5151), .ZN(n5177) );
  INV_X1 U6063 ( .A(n4835), .ZN(n4637) );
  NAND2_X1 U6064 ( .A1(n4638), .A2(n4641), .ZN(n5303) );
  NAND2_X1 U6065 ( .A1(n4647), .A2(n4341), .ZN(n5451) );
  NAND2_X1 U6066 ( .A1(n5581), .A2(n4651), .ZN(n4648) );
  NAND2_X1 U6067 ( .A1(n4648), .A2(n4649), .ZN(n7523) );
  NAND2_X1 U6068 ( .A1(n5581), .A2(n5580), .ZN(n4650) );
  OAI21_X1 U6069 ( .B1(n5469), .B2(n4658), .A(n4655), .ZN(n5511) );
  OAI21_X1 U6070 ( .B1(n5469), .B2(n5468), .A(n5470), .ZN(n5489) );
  NAND2_X1 U6071 ( .A1(n5468), .A2(n5470), .ZN(n4660) );
  NAND3_X1 U6072 ( .A1(n4662), .A2(n4661), .A3(n4903), .ZN(n4926) );
  NAND3_X1 U6073 ( .A1(n7315), .A2(n4668), .A3(n4667), .ZN(n4666) );
  OAI21_X1 U6074 ( .B1(n7075), .B2(n7759), .A(n4670), .ZN(n7316) );
  NAND2_X1 U6075 ( .A1(n4673), .A2(n4675), .ZN(n8239) );
  NAND2_X1 U6076 ( .A1(n4679), .A2(n4676), .ZN(n4673) );
  NAND2_X1 U6077 ( .A1(n4674), .A2(n4680), .ZN(n4679) );
  INV_X1 U6078 ( .A(n8281), .ZN(n4674) );
  INV_X1 U6079 ( .A(n8110), .ZN(n4688) );
  INV_X1 U6080 ( .A(n8128), .ZN(n4686) );
  NAND2_X1 U6081 ( .A1(n4682), .A2(n7837), .ZN(n8085) );
  NAND2_X1 U6082 ( .A1(n4331), .A2(n4683), .ZN(n4682) );
  INV_X2 U6083 ( .A(n4703), .ZN(n7003) );
  INV_X1 U6084 ( .A(n5806), .ZN(n4702) );
  NAND2_X1 U6085 ( .A1(n7918), .A2(n7003), .ZN(n7718) );
  NAND2_X1 U6086 ( .A1(n5806), .A2(n5805), .ZN(n7918) );
  NAND2_X1 U6087 ( .A1(n4700), .A2(n7003), .ZN(n4699) );
  INV_X1 U6088 ( .A(n5805), .ZN(n4700) );
  NAND2_X1 U6089 ( .A1(n4702), .A2(n7003), .ZN(n4701) );
  NAND2_X1 U6090 ( .A1(n6796), .A2(n4704), .ZN(n4705) );
  NAND2_X1 U6091 ( .A1(n5789), .A2(n4709), .ZN(n5797) );
  NAND2_X1 U6092 ( .A1(n4730), .A2(n8134), .ZN(n4729) );
  NAND2_X2 U6093 ( .A1(n6023), .A2(n6022), .ZN(n7595) );
  NAND2_X1 U6094 ( .A1(n7624), .A2(n7623), .ZN(n7622) );
  NAND2_X1 U6095 ( .A1(n6507), .A2(n4744), .ZN(n5778) );
  NAND2_X1 U6096 ( .A1(n4748), .A2(n4746), .ZN(n7544) );
  NAND2_X1 U6097 ( .A1(n4749), .A2(n4750), .ZN(n7537) );
  NAND2_X1 U6098 ( .A1(n6710), .A2(n6709), .ZN(n6708) );
  NAND2_X1 U6099 ( .A1(n6708), .A2(n5875), .ZN(n6713) );
  NOR2_X1 U6100 ( .A1(n6714), .A2(n5874), .ZN(n4753) );
  INV_X1 U6101 ( .A(n4764), .ZN(n4767) );
  NAND2_X1 U6102 ( .A1(n4764), .A2(n4277), .ZN(n4763) );
  NAND2_X1 U6103 ( .A1(n6034), .A2(n4771), .ZN(n5771) );
  NAND2_X1 U6104 ( .A1(n6034), .A2(n4769), .ZN(n4768) );
  NAND2_X1 U6105 ( .A1(n7377), .A2(n4784), .ZN(n4782) );
  NAND4_X1 U6106 ( .A1(n4847), .A2(n4952), .A3(n4848), .A4(n4953), .ZN(n5046)
         );
  NAND3_X1 U6107 ( .A1(n4952), .A2(n4847), .A3(n4953), .ZN(n5020) );
  NAND2_X1 U6108 ( .A1(n7153), .A2(n7154), .ZN(n4788) );
  NAND2_X1 U6109 ( .A1(n4788), .A2(n5094), .ZN(n5119) );
  NAND2_X1 U6110 ( .A1(n5037), .A2(n5036), .ZN(n4791) );
  AND2_X1 U6111 ( .A1(n4792), .A2(n4791), .ZN(n8473) );
  NAND2_X1 U6112 ( .A1(n4791), .A2(n8474), .ZN(n4790) );
  NAND2_X1 U6113 ( .A1(n4801), .A2(n5371), .ZN(n8519) );
  OR2_X1 U6114 ( .A1(n4801), .A2(n5371), .ZN(n8520) );
  INV_X1 U6115 ( .A(n8522), .ZN(n4798) );
  NOR2_X1 U6116 ( .A1(n5372), .A2(n8522), .ZN(n4800) );
  AND2_X1 U6117 ( .A1(n4859), .A2(n4802), .ZN(n4882) );
  NAND2_X1 U6118 ( .A1(n4859), .A2(n4858), .ZN(n4889) );
  NAND2_X1 U6119 ( .A1(n8433), .A2(n4805), .ZN(n4809) );
  AOI21_X1 U6120 ( .B1(n8505), .B2(n4814), .A(n4288), .ZN(n4805) );
  AND2_X1 U6121 ( .A1(n8433), .A2(n4811), .ZN(n4810) );
  AND2_X2 U6122 ( .A1(n4809), .A2(n4807), .ZN(n8533) );
  INV_X1 U6123 ( .A(n7492), .ZN(n4831) );
  NAND2_X1 U6124 ( .A1(n7492), .A2(n4827), .ZN(n4816) );
  OAI21_X2 U6125 ( .B1(n4831), .B2(n4824), .A(n4822), .ZN(n8421) );
  XNOR2_X1 U6126 ( .A(n7523), .B(n5705), .ZN(n7688) );
  NAND2_X1 U6127 ( .A1(n6329), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n5803) );
  NOR2_X2 U6128 ( .A1(n9160), .A2(n9254), .ZN(n9111) );
  INV_X1 U6129 ( .A(n7427), .ZN(n7428) );
  XNOR2_X1 U6130 ( .A(n7694), .B(SI_30_), .ZN(n8559) );
  NOR2_X1 U6131 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .ZN(
        n5761) );
  NAND2_X1 U6132 ( .A1(n6223), .A2(n6222), .ZN(n6224) );
  OR2_X2 U6133 ( .A1(n4989), .A2(n4918), .ZN(n4921) );
  INV_X1 U6134 ( .A(n5800), .ZN(n7525) );
  AOI21_X1 U6135 ( .B1(n5653), .B2(n5594), .A(n4911), .ZN(n6683) );
  INV_X1 U6136 ( .A(n4866), .ZN(n4869) );
  NAND2_X1 U6137 ( .A1(n7482), .A2(n5227), .ZN(n7492) );
  INV_X2 U6138 ( .A(n9572), .ZN(n9575) );
  OR2_X1 U6139 ( .A1(n5756), .A2(n9328), .ZN(n9617) );
  INV_X2 U6140 ( .A(n9617), .ZN(n9619) );
  AND2_X1 U6141 ( .A1(n6273), .A2(n6272), .ZN(n4834) );
  INV_X1 U6142 ( .A(P2_STATE_REG_SCAN_IN), .ZN(n6309) );
  AND2_X1 U6143 ( .A1(n5178), .A2(n5156), .ZN(n4835) );
  INV_X1 U6144 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n5072) );
  AND2_X1 U6145 ( .A1(n6051), .A2(n5769), .ZN(n4838) );
  AND2_X1 U6146 ( .A1(n5353), .A2(n4875), .ZN(n4839) );
  AND2_X1 U6147 ( .A1(n5151), .A2(n5137), .ZN(n4840) );
  AND2_X1 U6148 ( .A1(n5255), .A2(n5236), .ZN(n4841) );
  INV_X1 U6149 ( .A(n7230), .ZN(n5661) );
  AND2_X1 U6150 ( .A1(n8378), .A2(n7908), .ZN(n4842) );
  OR2_X1 U6151 ( .A1(n6346), .A2(n9470), .ZN(n4843) );
  INV_X1 U6152 ( .A(n5911), .ZN(n5932) );
  INV_X1 U6153 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5880) );
  INV_X1 U6154 ( .A(n7877), .ZN(n7047) );
  OR2_X1 U6155 ( .A1(n9264), .A2(n9255), .ZN(n4844) );
  XNOR2_X1 U6156 ( .A(n4959), .B(n7090), .ZN(n4960) );
  AND3_X1 U6157 ( .A1(n5628), .A2(n8475), .A3(n5627), .ZN(n4845) );
  AND2_X1 U6158 ( .A1(n8945), .A2(n8965), .ZN(n4846) );
  INV_X1 U6159 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n4854) );
  INV_X1 U6160 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n4849) );
  INV_X1 U6161 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n5769) );
  INV_X1 U6162 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n6024) );
  INV_X1 U6163 ( .A(n5118), .ZN(n5114) );
  OAI22_X1 U6164 ( .A1(n7100), .A2(n5485), .B1(n4912), .B2(n6287), .ZN(n4913)
         );
  INV_X1 U6165 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n4875) );
  INV_X1 U6166 ( .A(n6112), .ZN(n6111) );
  INV_X1 U6167 ( .A(n5995), .ZN(n5993) );
  NAND2_X1 U6168 ( .A1(n4980), .A2(n4979), .ZN(n4981) );
  OAI22_X1 U6169 ( .A1(n6942), .A2(n5012), .B1(n6939), .B2(n6940), .ZN(n5037)
         );
  CLKBUF_X3 U6170 ( .A(n4982), .Z(n5574) );
  INV_X1 U6171 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n5163) );
  INV_X1 U6172 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n5242) );
  INV_X1 U6173 ( .A(SI_22_), .ZN(n5452) );
  INV_X1 U6174 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n5157) );
  AND2_X1 U6175 ( .A1(P2_REG3_REG_7__SCAN_IN), .A2(P2_REG3_REG_6__SCAN_IN), 
        .ZN(n5897) );
  NAND2_X1 U6176 ( .A1(n5820), .A2(n9676), .ZN(n5816) );
  OR2_X1 U6177 ( .A1(n6134), .A2(n7558), .ZN(n6145) );
  NAND2_X1 U6178 ( .A1(n6084), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n6098) );
  INV_X1 U6179 ( .A(n6034), .ZN(n6035) );
  OR2_X1 U6180 ( .A1(n5432), .A2(n5431), .ZN(n5458) );
  AND2_X1 U6181 ( .A1(n5289), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n5312) );
  INV_X1 U6182 ( .A(n4867), .ZN(n4868) );
  OR2_X1 U6183 ( .A1(n5332), .A2(n5331), .ZN(n5360) );
  OAI22_X1 U6184 ( .A1(n9557), .A2(n5665), .B1(n8845), .B2(n9555), .ZN(n7361)
         );
  NAND2_X1 U6185 ( .A1(n9602), .A2(n9596), .ZN(n8689) );
  NAND2_X1 U6186 ( .A1(n4887), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4884) );
  OR2_X1 U6187 ( .A1(n6048), .A2(n6047), .ZN(n6049) );
  INV_X1 U6188 ( .A(n7669), .ZN(n7645) );
  OR2_X1 U6189 ( .A1(n6171), .A2(n7654), .ZN(n6202) );
  OR2_X1 U6190 ( .A1(n6370), .A2(n6369), .ZN(n9629) );
  AND2_X1 U6191 ( .A1(n7766), .A2(n7769), .ZN(n7168) );
  OR2_X1 U6192 ( .A1(n9669), .A2(n6781), .ZN(n8142) );
  INV_X1 U6193 ( .A(n8050), .ZN(n8283) );
  INV_X1 U6194 ( .A(n7780), .ZN(n9386) );
  INV_X1 U6195 ( .A(n7908), .ZN(n7434) );
  INV_X1 U6196 ( .A(n8419), .ZN(n6243) );
  INV_X1 U6197 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5796) );
  NAND2_X1 U6198 ( .A1(n8558), .A2(n5621), .ZN(n8680) );
  XNOR2_X1 U6199 ( .A(n4984), .B(n4985), .ZN(n6930) );
  AND2_X1 U6200 ( .A1(n5634), .A2(n6679), .ZN(n8550) );
  INV_X1 U6201 ( .A(n5640), .ZN(n5495) );
  INV_X1 U6202 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n8425) );
  AND2_X1 U6203 ( .A1(n6344), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6400) );
  AND2_X1 U6204 ( .A1(n8612), .A2(n8614), .ZN(n8709) );
  INV_X1 U6205 ( .A(n8843), .ZN(n9413) );
  INV_X1 U6206 ( .A(n5723), .ZN(n8704) );
  INV_X1 U6207 ( .A(n9123), .ZN(n9074) );
  OR2_X1 U6208 ( .A1(n8765), .A2(n4541), .ZN(n9150) );
  OR2_X1 U6209 ( .A1(n7089), .A2(n8832), .ZN(n9612) );
  NAND2_X1 U6210 ( .A1(n5630), .A2(n9577), .ZN(n7088) );
  INV_X1 U6211 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n4909) );
  AND2_X1 U6212 ( .A1(n5428), .A2(n5406), .ZN(n5426) );
  AND2_X1 U6213 ( .A1(n5327), .A2(n5307), .ZN(n5325) );
  AND2_X1 U6214 ( .A1(n6270), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7657) );
  INV_X1 U6215 ( .A(n6249), .ZN(n6259) );
  OR2_X1 U6216 ( .A1(n6271), .A2(n6262), .ZN(n6209) );
  AND4_X1 U6217 ( .A1(n6031), .A2(n6030), .A3(n6029), .A4(n6028), .ZN(n7683)
         );
  INV_X1 U6218 ( .A(n8029), .ZN(n9632) );
  INV_X1 U6219 ( .A(n8064), .ZN(n8061) );
  INV_X1 U6220 ( .A(n7168), .ZN(n7881) );
  INV_X1 U6221 ( .A(n8142), .ZN(n9665) );
  AND2_X1 U6222 ( .A1(n9661), .A2(n6788), .ZN(n9648) );
  NOR2_X1 U6223 ( .A1(n9672), .A2(n6239), .ZN(n6701) );
  NOR2_X2 U6224 ( .A1(n9652), .A2(n9715), .ZN(n9678) );
  AND2_X1 U6225 ( .A1(n7897), .A2(n6505), .ZN(n9715) );
  INV_X1 U6226 ( .A(n9678), .ZN(n9733) );
  AND2_X1 U6227 ( .A1(n6243), .A2(n6228), .ZN(n9668) );
  INV_X1 U6228 ( .A(n7464), .ZN(n8552) );
  AOI21_X1 U6229 ( .B1(n5484), .B2(n5495), .A(n5483), .ZN(n9201) );
  OR2_X1 U6230 ( .A1(n5640), .A2(n5014), .ZN(n5019) );
  AND2_X1 U6231 ( .A1(n6400), .A2(n6399), .ZN(n9530) );
  INV_X1 U6232 ( .A(n9533), .ZN(n9514) );
  INV_X1 U6233 ( .A(n9525), .ZN(n9539) );
  INV_X1 U6234 ( .A(n9079), .ZN(n9563) );
  INV_X1 U6235 ( .A(n9438), .ZN(n9603) );
  NAND2_X1 U6236 ( .A1(n9419), .A2(n9582), .ZN(n9615) );
  INV_X1 U6237 ( .A(n9419), .ZN(n9587) );
  NAND2_X1 U6238 ( .A1(n5601), .A2(n5603), .ZN(n9576) );
  AND2_X1 U6239 ( .A1(n5261), .A2(n5284), .ZN(n9513) );
  NAND2_X1 U6240 ( .A1(n6326), .A2(n6325), .ZN(n9633) );
  NAND2_X1 U6241 ( .A1(n6617), .A2(n6248), .ZN(n7660) );
  OR2_X1 U6242 ( .A1(n6360), .A2(n6286), .ZN(n7906) );
  OR2_X1 U6243 ( .A1(n8033), .A2(n7528), .ZN(n8029) );
  NAND2_X1 U6244 ( .A1(n9661), .A2(n6782), .ZN(n9649) );
  INV_X1 U6245 ( .A(n9752), .ZN(n9750) );
  INV_X1 U6246 ( .A(n9736), .ZN(n9734) );
  AND2_X2 U6247 ( .A1(n6702), .A2(n6778), .ZN(n9736) );
  NOR2_X1 U6248 ( .A1(n9669), .A2(n9668), .ZN(n9670) );
  NAND2_X1 U6249 ( .A1(n5792), .A2(n5791), .ZN(n8413) );
  INV_X1 U6250 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7251) );
  INV_X1 U6251 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6626) );
  OR2_X1 U6252 ( .A1(n6287), .A2(n6288), .ZN(n6341) );
  NOR2_X1 U6253 ( .A1(n4845), .A2(n5649), .ZN(n5650) );
  INV_X1 U6254 ( .A(n9555), .ZN(n9613) );
  NAND2_X1 U6255 ( .A1(n6679), .A2(n5629), .ZN(n7464) );
  NAND2_X1 U6256 ( .A1(n5501), .A2(n5500), .ZN(n9023) );
  INV_X1 U6257 ( .A(n9530), .ZN(n9503) );
  OR2_X1 U6258 ( .A1(P1_U3083), .A2(n6342), .ZN(n9525) );
  NAND2_X1 U6259 ( .A1(n9572), .A2(n4348), .ZN(n9060) );
  NAND2_X1 U6260 ( .A1(n9572), .A2(n7092), .ZN(n9079) );
  NAND2_X1 U6261 ( .A1(n4270), .A2(n9452), .ZN(n9280) );
  INV_X1 U6262 ( .A(n8990), .ZN(n9299) );
  NAND2_X1 U6263 ( .A1(n9619), .A2(n9452), .ZN(n9326) );
  AND2_X1 U6264 ( .A1(n9577), .A2(n9576), .ZN(n9578) );
  INV_X1 U6265 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n9341) );
  INV_X1 U6266 ( .A(n5621), .ZN(n8801) );
  INV_X1 U6267 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n6810) );
  INV_X1 U6268 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n6336) );
  NOR2_X1 U6269 ( .A1(n9780), .A2(n9779), .ZN(n9778) );
  OAI21_X1 U6270 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n9769), .ZN(n9767) );
  INV_X2 U6271 ( .A(n7906), .ZN(P2_U3966) );
  NOR2_X4 U6272 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n4952) );
  NOR2_X2 U6273 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n4850) );
  AND4_X2 U6274 ( .A1(n4850), .A2(n4849), .A3(n5138), .A4(n5157), .ZN(n4851)
         );
  NOR2_X1 U6275 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n4853) );
  NAND4_X1 U6276 ( .A1(n4853), .A2(n4877), .A3(n4881), .A4(n4897), .ZN(n4856)
         );
  NAND4_X1 U6277 ( .A1(n4894), .A2(n5259), .A3(n5353), .A4(n4854), .ZN(n4855)
         );
  NOR2_X1 U6278 ( .A1(n4856), .A2(n4855), .ZN(n4857) );
  NOR2_X2 U6279 ( .A1(n4905), .A2(P1_IR_REG_28__SCAN_IN), .ZN(n4862) );
  NAND2_X1 U6280 ( .A1(n4862), .A2(n4863), .ZN(n9329) );
  NAND2_X1 U6281 ( .A1(n5070), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n4872) );
  NAND2_X1 U6282 ( .A1(n5162), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n4871) );
  INV_X1 U6283 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n9566) );
  NOR2_X1 U6284 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n4874) );
  NAND2_X1 U6285 ( .A1(n5257), .A2(n4874), .ZN(n5308) );
  NAND2_X1 U6286 ( .A1(n4878), .A2(n4877), .ZN(n4893) );
  INV_X1 U6287 ( .A(n4885), .ZN(n4886) );
  NAND2_X1 U6288 ( .A1(n4886), .A2(P1_IR_REG_25__SCAN_IN), .ZN(n4888) );
  NAND2_X1 U6289 ( .A1(n4888), .A2(n4887), .ZN(n7478) );
  NAND2_X1 U6290 ( .A1(n4889), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4891) );
  INV_X1 U6291 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n4890) );
  NOR2_X1 U6292 ( .A1(n7478), .A2(n7402), .ZN(n4892) );
  NAND2_X1 U6293 ( .A1(n4896), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4898) );
  XNOR2_X2 U6294 ( .A(n4898), .B(n4897), .ZN(n9123) );
  NAND2_X1 U6295 ( .A1(n4265), .A2(n8832), .ZN(n4899) );
  INV_X1 U6296 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n6352) );
  INV_X1 U6297 ( .A(SI_0_), .ZN(n9835) );
  INV_X1 U6298 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n4902) );
  OAI21_X1 U6299 ( .B1(n7698), .B2(n9835), .A(n4902), .ZN(n4904) );
  AND2_X1 U6300 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n4903) );
  NAND2_X1 U6301 ( .A1(n4904), .A2(n4926), .ZN(n9345) );
  NAND2_X1 U6302 ( .A1(n4905), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4907) );
  NAND2_X1 U6303 ( .A1(n5710), .A2(n6287), .ZN(n5577) );
  OAI22_X1 U6304 ( .A1(n7100), .A2(n5577), .B1(n6352), .B2(n6287), .ZN(n4911)
         );
  INV_X2 U6305 ( .A(n5577), .ZN(n4982) );
  NAND2_X1 U6306 ( .A1(n5653), .A2(n4982), .ZN(n4915) );
  INV_X1 U6307 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n4912) );
  INV_X1 U6308 ( .A(n4913), .ZN(n4914) );
  NAND2_X1 U6309 ( .A1(n4915), .A2(n4914), .ZN(n6681) );
  NAND2_X1 U6310 ( .A1(n6683), .A2(n6681), .ZN(n6682) );
  NAND2_X1 U6311 ( .A1(n8558), .A2(n9123), .ZN(n5712) );
  NAND2_X1 U6312 ( .A1(n6682), .A2(n4298), .ZN(n4935) );
  INV_X1 U6313 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n4917) );
  OR2_X1 U6314 ( .A1(n4992), .A2(n4917), .ZN(n4922) );
  INV_X1 U6315 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n4918) );
  INV_X1 U6316 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n7101) );
  OR2_X1 U6317 ( .A1(n4991), .A2(n7101), .ZN(n4920) );
  INV_X1 U6318 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n4924) );
  NAND2_X1 U6319 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n4923) );
  INV_X1 U6320 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6303) );
  NAND3_X1 U6321 ( .A1(n7698), .A2(SI_0_), .A3(P1_DATAO_REG_0__SCAN_IN), .ZN(
        n4925) );
  INV_X1 U6322 ( .A(SI_1_), .ZN(n4927) );
  XNOR2_X1 U6323 ( .A(n4947), .B(n4946), .ZN(n6302) );
  OR2_X1 U6324 ( .A1(n4971), .A2(n6302), .ZN(n4928) );
  OAI211_X2 U6325 ( .C1(n6346), .C2(n6582), .A(n4929), .B(n4928), .ZN(n7103)
         );
  INV_X2 U6326 ( .A(n5485), .ZN(n5598) );
  NAND2_X1 U6327 ( .A1(n7103), .A2(n5598), .ZN(n4930) );
  NAND2_X1 U6328 ( .A1(n4931), .A2(n4930), .ZN(n4932) );
  XNOR2_X1 U6329 ( .A(n4932), .B(n7090), .ZN(n4936) );
  NAND2_X1 U6330 ( .A1(n4935), .A2(n4936), .ZN(n6857) );
  NAND2_X1 U6331 ( .A1(n8849), .A2(n5594), .ZN(n4934) );
  NAND2_X1 U6332 ( .A1(n7103), .A2(n4982), .ZN(n4933) );
  NAND2_X1 U6333 ( .A1(n4934), .A2(n4933), .ZN(n6860) );
  NAND2_X1 U6334 ( .A1(n6857), .A2(n6860), .ZN(n4939) );
  INV_X1 U6335 ( .A(n4935), .ZN(n4938) );
  INV_X1 U6336 ( .A(n4936), .ZN(n4937) );
  NAND2_X1 U6337 ( .A1(n4938), .A2(n4937), .ZN(n6858) );
  NAND2_X1 U6338 ( .A1(n4939), .A2(n6858), .ZN(n6865) );
  INV_X1 U6339 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n4940) );
  NAND2_X1 U6340 ( .A1(n5070), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n4944) );
  INV_X1 U6341 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n4941) );
  INV_X1 U6342 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n9469) );
  OR2_X1 U6343 ( .A1(n4991), .A2(n9469), .ZN(n4942) );
  NAND4_X2 U6344 ( .A1(n4945), .A2(n4944), .A3(n4943), .A4(n4942), .ZN(n5655)
         );
  NAND2_X1 U6345 ( .A1(n5655), .A2(n4982), .ZN(n4958) );
  NAND2_X1 U6346 ( .A1(n4947), .A2(n4946), .ZN(n4950) );
  NAND2_X1 U6347 ( .A1(n4948), .A2(SI_1_), .ZN(n4949) );
  INV_X1 U6348 ( .A(SI_2_), .ZN(n4951) );
  XNOR2_X1 U6349 ( .A(n4973), .B(n4972), .ZN(n6304) );
  OR2_X1 U6350 ( .A1(n4971), .A2(n6304), .ZN(n4954) );
  OR2_X1 U6351 ( .A1(n4952), .A2(n9330), .ZN(n4998) );
  NAND2_X1 U6352 ( .A1(n4998), .A2(n4953), .ZN(n4968) );
  OAI21_X1 U6353 ( .B1(n4998), .B2(n4953), .A(n4968), .ZN(n9470) );
  INV_X1 U6354 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6305) );
  OR2_X1 U6355 ( .A1(n5000), .A2(n6305), .ZN(n4955) );
  NAND2_X1 U6356 ( .A1(n7186), .A2(n5598), .ZN(n4957) );
  NAND2_X1 U6357 ( .A1(n4958), .A2(n4957), .ZN(n4959) );
  AOI22_X1 U6358 ( .A1(n5655), .A2(n5594), .B1(n4982), .B2(n7186), .ZN(n4961)
         );
  XNOR2_X1 U6359 ( .A(n4960), .B(n4961), .ZN(n6866) );
  NAND2_X1 U6360 ( .A1(n4960), .A2(n4961), .ZN(n4962) );
  OAI21_X1 U6361 ( .B1(n6865), .B2(n6866), .A(n4962), .ZN(n6931) );
  NAND2_X1 U6362 ( .A1(n5070), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n4967) );
  INV_X1 U6363 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n6389) );
  OR2_X1 U6364 ( .A1(n4992), .A2(n6389), .ZN(n4966) );
  INV_X1 U6365 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n4963) );
  OR2_X1 U6366 ( .A1(n4989), .A2(n4963), .ZN(n4965) );
  OR2_X1 U6367 ( .A1(n4991), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n4964) );
  NAND2_X1 U6368 ( .A1(n8848), .A2(n4982), .ZN(n4980) );
  NAND2_X1 U6369 ( .A1(n4968), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4970) );
  INV_X1 U6370 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n4969) );
  INV_X1 U6371 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6301) );
  OR2_X1 U6372 ( .A1(n5000), .A2(n6301), .ZN(n4978) );
  NAND2_X1 U6373 ( .A1(n4973), .A2(n4972), .ZN(n4976) );
  NAND2_X1 U6374 ( .A1(n4974), .A2(SI_2_), .ZN(n4975) );
  INV_X1 U6375 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6293) );
  XNOR2_X1 U6376 ( .A(n5003), .B(SI_3_), .ZN(n5001) );
  XNOR2_X1 U6377 ( .A(n5002), .B(n5001), .ZN(n6300) );
  OR2_X1 U6378 ( .A1(n4971), .A2(n6300), .ZN(n4977) );
  OAI211_X1 U6379 ( .C1(n6346), .C2(n8850), .A(n4978), .B(n4977), .ZN(n7510)
         );
  NAND2_X1 U6380 ( .A1(n7510), .A2(n5598), .ZN(n4979) );
  AND2_X1 U6381 ( .A1(n7510), .A2(n4982), .ZN(n4983) );
  AOI21_X1 U6382 ( .B1(n8848), .B2(n5594), .A(n4983), .ZN(n4985) );
  NAND2_X1 U6383 ( .A1(n6931), .A2(n6930), .ZN(n4988) );
  INV_X1 U6384 ( .A(n4984), .ZN(n4986) );
  NAND2_X1 U6385 ( .A1(n4986), .A2(n4985), .ZN(n4987) );
  NAND2_X1 U6386 ( .A1(n4988), .A2(n4987), .ZN(n6942) );
  NAND2_X1 U6387 ( .A1(n4272), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n4996) );
  INV_X1 U6388 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n6416) );
  OR2_X1 U6389 ( .A1(n4273), .A2(n6416), .ZN(n4995) );
  XNOR2_X1 U6390 ( .A(P1_REG3_REG_3__SCAN_IN), .B(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n7194) );
  OR2_X1 U6391 ( .A1(n5640), .A2(n7194), .ZN(n4994) );
  INV_X1 U6392 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6391) );
  OR2_X1 U6393 ( .A1(n5241), .A2(n6391), .ZN(n4993) );
  NAND2_X1 U6394 ( .A1(n8847), .A2(n4982), .ZN(n5009) );
  OAI21_X1 U6395 ( .B1(P1_IR_REG_2__SCAN_IN), .B2(P1_IR_REG_3__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n4997) );
  NAND2_X1 U6396 ( .A1(n4998), .A2(n4997), .ZN(n4999) );
  XNOR2_X1 U6397 ( .A(n4999), .B(P1_IR_REG_4__SCAN_IN), .ZN(n9483) );
  OR2_X1 U6398 ( .A1(n5000), .A2(n6296), .ZN(n5007) );
  INV_X1 U6399 ( .A(n5003), .ZN(n5004) );
  NAND2_X1 U6400 ( .A1(n5004), .A2(SI_3_), .ZN(n5005) );
  XNOR2_X1 U6401 ( .A(n5024), .B(SI_4_), .ZN(n5022) );
  XNOR2_X1 U6402 ( .A(n5023), .B(n5022), .ZN(n6295) );
  OR2_X1 U6403 ( .A1(n4971), .A2(n6295), .ZN(n5006) );
  OAI211_X1 U6404 ( .C1(n9483), .C2(n6346), .A(n5007), .B(n5006), .ZN(n7196)
         );
  NAND2_X1 U6405 ( .A1(n7196), .A2(n5598), .ZN(n5008) );
  NAND2_X1 U6406 ( .A1(n5009), .A2(n5008), .ZN(n5010) );
  XNOR2_X1 U6407 ( .A(n5010), .B(n7090), .ZN(n6939) );
  AND2_X1 U6408 ( .A1(n7196), .A2(n5574), .ZN(n5011) );
  AOI21_X1 U6409 ( .B1(n8847), .B2(n5594), .A(n5011), .ZN(n6940) );
  AND2_X1 U6410 ( .A1(n6939), .A2(n6940), .ZN(n5012) );
  INV_X1 U6411 ( .A(n5037), .ZN(n5035) );
  AOI21_X1 U6412 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(P1_REG3_REG_5__SCAN_IN), .ZN(n5013) );
  NOR2_X1 U6413 ( .A1(n5013), .A2(n5040), .ZN(n8478) );
  INV_X1 U6414 ( .A(n8478), .ZN(n5014) );
  INV_X1 U6415 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n5015) );
  OR2_X1 U6416 ( .A1(n4989), .A2(n5015), .ZN(n5018) );
  INV_X1 U6417 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n6418) );
  OR2_X1 U6418 ( .A1(n4273), .A2(n6418), .ZN(n5017) );
  INV_X1 U6419 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n7224) );
  OR2_X1 U6420 ( .A1(n5241), .A2(n7224), .ZN(n5016) );
  NAND4_X1 U6421 ( .A1(n5019), .A2(n5018), .A3(n5017), .A4(n5016), .ZN(n9602)
         );
  NAND2_X1 U6422 ( .A1(n9602), .A2(n4982), .ZN(n5031) );
  NAND2_X1 U6423 ( .A1(n5020), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5021) );
  XNOR2_X1 U6424 ( .A(n5021), .B(n4848), .ZN(n8863) );
  OR2_X1 U6425 ( .A1(n5000), .A2(n6299), .ZN(n5029) );
  INV_X1 U6426 ( .A(n5024), .ZN(n5025) );
  NAND2_X1 U6427 ( .A1(n5025), .A2(SI_4_), .ZN(n5026) );
  XNOR2_X1 U6428 ( .A(n5054), .B(SI_5_), .ZN(n5052) );
  XNOR2_X1 U6429 ( .A(n5053), .B(n5052), .ZN(n6298) );
  OR2_X1 U6430 ( .A1(n4971), .A2(n6298), .ZN(n5028) );
  OAI211_X1 U6431 ( .C1(n6346), .C2(n8863), .A(n5029), .B(n5028), .ZN(n8477)
         );
  NAND2_X1 U6432 ( .A1(n8477), .A2(n5598), .ZN(n5030) );
  NAND2_X1 U6433 ( .A1(n5031), .A2(n5030), .ZN(n5033) );
  XNOR2_X1 U6434 ( .A(n5033), .B(n5032), .ZN(n5036) );
  AND2_X1 U6435 ( .A1(n8477), .A2(n5574), .ZN(n5038) );
  AOI21_X1 U6436 ( .B1(n9602), .B2(n5594), .A(n5038), .ZN(n8474) );
  NAND2_X1 U6437 ( .A1(n4272), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5045) );
  INV_X1 U6438 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n5039) );
  OR2_X1 U6439 ( .A1(n4273), .A2(n5039), .ZN(n5044) );
  NAND2_X1 U6440 ( .A1(n5040), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5073) );
  OAI21_X1 U6441 ( .B1(n5040), .B2(P1_REG3_REG_6__SCAN_IN), .A(n5073), .ZN(
        n7240) );
  OR2_X1 U6442 ( .A1(n5640), .A2(n7240), .ZN(n5043) );
  INV_X1 U6443 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n5041) );
  OR2_X1 U6444 ( .A1(n5241), .A2(n5041), .ZN(n5042) );
  NAND4_X1 U6445 ( .A1(n5045), .A2(n5044), .A3(n5043), .A4(n5042), .ZN(n8846)
         );
  NAND2_X1 U6446 ( .A1(n8846), .A2(n5574), .ZN(n5061) );
  NAND2_X1 U6447 ( .A1(n5046), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5047) );
  MUX2_X1 U6448 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5047), .S(
        P1_IR_REG_6__SCAN_IN), .Z(n5051) );
  INV_X1 U6449 ( .A(n5049), .ZN(n5050) );
  NAND2_X1 U6450 ( .A1(n5051), .A2(n5050), .ZN(n6420) );
  OR2_X1 U6451 ( .A1(n5000), .A2(n6308), .ZN(n5059) );
  NAND2_X1 U6452 ( .A1(n5053), .A2(n5052), .ZN(n5057) );
  INV_X1 U6453 ( .A(n5054), .ZN(n5055) );
  NAND2_X1 U6454 ( .A1(n5055), .A2(SI_5_), .ZN(n5056) );
  XNOR2_X1 U6455 ( .A(n5083), .B(SI_6_), .ZN(n5081) );
  XNOR2_X1 U6456 ( .A(n5082), .B(n5081), .ZN(n6307) );
  OR2_X1 U6457 ( .A1(n4971), .A2(n6307), .ZN(n5058) );
  NAND2_X1 U6458 ( .A1(n4269), .A2(n5598), .ZN(n5060) );
  NAND2_X1 U6459 ( .A1(n5061), .A2(n5060), .ZN(n5062) );
  XNOR2_X1 U6460 ( .A(n5062), .B(n5032), .ZN(n5065) );
  NAND2_X1 U6461 ( .A1(n8846), .A2(n5594), .ZN(n5064) );
  NAND2_X1 U6462 ( .A1(n4269), .A2(n5574), .ZN(n5063) );
  NAND2_X1 U6463 ( .A1(n5064), .A2(n5063), .ZN(n5066) );
  NAND2_X1 U6464 ( .A1(n5065), .A2(n5066), .ZN(n7126) );
  NAND2_X1 U6465 ( .A1(n7127), .A2(n7126), .ZN(n5069) );
  INV_X1 U6466 ( .A(n5065), .ZN(n5068) );
  INV_X1 U6467 ( .A(n5066), .ZN(n5067) );
  NAND2_X1 U6468 ( .A1(n5068), .A2(n5067), .ZN(n7125) );
  NAND2_X1 U6469 ( .A1(n5069), .A2(n7125), .ZN(n7153) );
  NAND2_X1 U6470 ( .A1(n5585), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5079) );
  INV_X1 U6471 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n5071) );
  OR2_X1 U6472 ( .A1(n5241), .A2(n5071), .ZN(n5078) );
  AND2_X1 U6473 ( .A1(n5073), .A2(n5072), .ZN(n5074) );
  NOR2_X1 U6474 ( .A1(n5073), .A2(n5072), .ZN(n5095) );
  OR2_X1 U6475 ( .A1(n5074), .A2(n5095), .ZN(n7157) );
  OR2_X1 U6476 ( .A1(n5640), .A2(n7157), .ZN(n5077) );
  INV_X1 U6477 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n5075) );
  OR2_X1 U6478 ( .A1(n4989), .A2(n5075), .ZN(n5076) );
  NAND4_X1 U6479 ( .A1(n5079), .A2(n5078), .A3(n5077), .A4(n5076), .ZN(n9601)
         );
  NAND2_X1 U6480 ( .A1(n9601), .A2(n5574), .ZN(n5088) );
  OR2_X1 U6481 ( .A1(n5049), .A2(n9330), .ZN(n5080) );
  XNOR2_X1 U6482 ( .A(n5080), .B(P1_IR_REG_7__SCAN_IN), .ZN(n6603) );
  INV_X1 U6483 ( .A(n6603), .ZN(n6311) );
  INV_X1 U6484 ( .A(n5083), .ZN(n5084) );
  NAND2_X1 U6485 ( .A1(n5084), .A2(SI_6_), .ZN(n5085) );
  XNOR2_X1 U6486 ( .A(n5104), .B(SI_7_), .ZN(n5103) );
  OR2_X1 U6487 ( .A1(n5000), .A2(n6313), .ZN(n5086) );
  NAND2_X1 U6488 ( .A1(n7158), .A2(n5598), .ZN(n5087) );
  NAND2_X1 U6489 ( .A1(n5088), .A2(n5087), .ZN(n5089) );
  XNOR2_X1 U6490 ( .A(n5089), .B(n5032), .ZN(n5091) );
  AND2_X1 U6491 ( .A1(n7158), .A2(n5574), .ZN(n5090) );
  AOI21_X1 U6492 ( .B1(n9601), .B2(n5594), .A(n5090), .ZN(n5092) );
  XNOR2_X1 U6493 ( .A(n5091), .B(n5092), .ZN(n7154) );
  INV_X1 U6494 ( .A(n5091), .ZN(n5093) );
  NAND2_X1 U6495 ( .A1(n5093), .A2(n5092), .ZN(n5094) );
  NAND2_X1 U6496 ( .A1(n4272), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n5100) );
  INV_X1 U6497 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n6407) );
  OR2_X1 U6498 ( .A1(n4273), .A2(n6407), .ZN(n5099) );
  NAND2_X1 U6499 ( .A1(n5095), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5122) );
  OR2_X1 U6500 ( .A1(n5095), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5096) );
  NAND2_X1 U6501 ( .A1(n5122), .A2(n5096), .ZN(n7353) );
  OR2_X1 U6502 ( .A1(n5640), .A2(n7353), .ZN(n5098) );
  INV_X1 U6503 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n6395) );
  OR2_X1 U6504 ( .A1(n5241), .A2(n6395), .ZN(n5097) );
  NAND4_X1 U6505 ( .A1(n5100), .A2(n5099), .A3(n5098), .A4(n5097), .ZN(n9547)
         );
  INV_X1 U6506 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n5101) );
  AND2_X1 U6507 ( .A1(n5049), .A2(n5101), .ZN(n5139) );
  OR2_X1 U6508 ( .A1(n5139), .A2(n9330), .ZN(n5102) );
  XNOR2_X1 U6509 ( .A(n5102), .B(P1_IR_REG_8__SCAN_IN), .ZN(n6456) );
  INV_X1 U6510 ( .A(n6456), .ZN(n6463) );
  INV_X1 U6511 ( .A(n5104), .ZN(n5105) );
  INV_X1 U6512 ( .A(SI_8_), .ZN(n5106) );
  NAND2_X1 U6513 ( .A1(n5107), .A2(n5106), .ZN(n5132) );
  INV_X1 U6514 ( .A(n5107), .ZN(n5108) );
  NAND2_X1 U6515 ( .A1(n5108), .A2(SI_8_), .ZN(n5109) );
  NAND2_X1 U6516 ( .A1(n5132), .A2(n5109), .ZN(n5130) );
  INV_X1 U6517 ( .A(n5130), .ZN(n5110) );
  XNOR2_X1 U6518 ( .A(n5131), .B(n5110), .ZN(n6317) );
  OR2_X1 U6519 ( .A1(n5000), .A2(n6316), .ZN(n5111) );
  OAI211_X1 U6520 ( .C1(n6346), .C2(n6463), .A(n5112), .B(n5111), .ZN(n7352)
         );
  AND2_X1 U6521 ( .A1(n7352), .A2(n5574), .ZN(n5113) );
  AOI21_X1 U6522 ( .B1(n9547), .B2(n5594), .A(n5113), .ZN(n5118) );
  NAND2_X1 U6523 ( .A1(n9547), .A2(n5574), .ZN(n5116) );
  NAND2_X1 U6524 ( .A1(n7352), .A2(n5598), .ZN(n5115) );
  NAND2_X1 U6525 ( .A1(n5116), .A2(n5115), .ZN(n5117) );
  XNOR2_X1 U6526 ( .A(n5117), .B(n7090), .ZN(n7328) );
  NAND2_X1 U6527 ( .A1(n7326), .A2(n7328), .ZN(n5120) );
  NAND2_X1 U6528 ( .A1(n5119), .A2(n5118), .ZN(n7327) );
  NAND2_X1 U6529 ( .A1(n5120), .A2(n7327), .ZN(n7377) );
  NAND2_X1 U6530 ( .A1(n4272), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5129) );
  NAND2_X1 U6531 ( .A1(n5122), .A2(n5121), .ZN(n5123) );
  NAND2_X1 U6532 ( .A1(n5164), .A2(n5123), .ZN(n9551) );
  OR2_X1 U6533 ( .A1(n5640), .A2(n9551), .ZN(n5128) );
  INV_X1 U6534 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n5124) );
  OR2_X1 U6535 ( .A1(n4273), .A2(n5124), .ZN(n5127) );
  INV_X1 U6536 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n5125) );
  OR2_X1 U6537 ( .A1(n5241), .A2(n5125), .ZN(n5126) );
  NAND4_X1 U6538 ( .A1(n5129), .A2(n5128), .A3(n5127), .A4(n5126), .ZN(n8845)
         );
  NAND2_X1 U6539 ( .A1(n8845), .A2(n5574), .ZN(n5144) );
  INV_X1 U6540 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n5133) );
  INV_X1 U6541 ( .A(SI_9_), .ZN(n5134) );
  NAND2_X1 U6542 ( .A1(n5135), .A2(n5134), .ZN(n5151) );
  INV_X1 U6543 ( .A(n5135), .ZN(n5136) );
  NAND2_X1 U6544 ( .A1(n5136), .A2(SI_9_), .ZN(n5137) );
  XNOR2_X1 U6545 ( .A(n5150), .B(n4840), .ZN(n6319) );
  NAND2_X1 U6546 ( .A1(n6319), .A2(n8563), .ZN(n5142) );
  AND2_X1 U6547 ( .A1(n5139), .A2(n5138), .ZN(n5158) );
  OR2_X1 U6548 ( .A1(n5158), .A2(n9330), .ZN(n5140) );
  XNOR2_X1 U6549 ( .A(n5140), .B(P1_IR_REG_9__SCAN_IN), .ZN(n9499) );
  AOI22_X1 U6550 ( .A1(n5381), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n6290), .B2(
        n9499), .ZN(n5141) );
  NAND2_X1 U6551 ( .A1(n5142), .A2(n5141), .ZN(n9555) );
  NAND2_X1 U6552 ( .A1(n9555), .A2(n5598), .ZN(n5143) );
  NAND2_X1 U6553 ( .A1(n5144), .A2(n5143), .ZN(n5145) );
  XNOR2_X1 U6554 ( .A(n5145), .B(n5032), .ZN(n5146) );
  AOI22_X1 U6555 ( .A1(n8845), .A2(n5594), .B1(n9555), .B2(n4982), .ZN(n5147)
         );
  XNOR2_X1 U6556 ( .A(n5146), .B(n5147), .ZN(n7378) );
  INV_X1 U6557 ( .A(n5146), .ZN(n5148) );
  NAND2_X1 U6558 ( .A1(n5148), .A2(n5147), .ZN(n5149) );
  NAND2_X1 U6559 ( .A1(n5150), .A2(n4840), .ZN(n5152) );
  INV_X1 U6560 ( .A(SI_10_), .ZN(n5153) );
  NAND2_X1 U6561 ( .A1(n5154), .A2(n5153), .ZN(n5178) );
  INV_X1 U6562 ( .A(n5154), .ZN(n5155) );
  NAND2_X1 U6563 ( .A1(n5155), .A2(SI_10_), .ZN(n5156) );
  XNOR2_X1 U6564 ( .A(n5177), .B(n4835), .ZN(n6335) );
  NAND2_X1 U6565 ( .A1(n6335), .A2(n8563), .ZN(n5161) );
  NAND2_X1 U6566 ( .A1(n5158), .A2(n5157), .ZN(n5179) );
  NAND2_X1 U6567 ( .A1(n5179), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5159) );
  XNOR2_X1 U6568 ( .A(n5159), .B(P1_IR_REG_10__SCAN_IN), .ZN(n6487) );
  AOI22_X1 U6569 ( .A1(n5381), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n6290), .B2(
        n6487), .ZN(n5160) );
  NAND2_X1 U6570 ( .A1(n9373), .A2(n5598), .ZN(n5172) );
  NAND2_X1 U6571 ( .A1(n5162), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n5170) );
  INV_X1 U6572 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n6422) );
  OR2_X1 U6573 ( .A1(n4273), .A2(n6422), .ZN(n5169) );
  NAND2_X1 U6574 ( .A1(n5164), .A2(n5163), .ZN(n5165) );
  NAND2_X1 U6575 ( .A1(n5185), .A2(n5165), .ZN(n7408) );
  OR2_X1 U6576 ( .A1(n5640), .A2(n7408), .ZN(n5168) );
  INV_X1 U6577 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n5166) );
  OR2_X1 U6578 ( .A1(n4989), .A2(n5166), .ZN(n5167) );
  NAND4_X1 U6579 ( .A1(n5170), .A2(n5169), .A3(n5168), .A4(n5167), .ZN(n9548)
         );
  NAND2_X1 U6580 ( .A1(n9548), .A2(n5574), .ZN(n5171) );
  NAND2_X1 U6581 ( .A1(n5172), .A2(n5171), .ZN(n5173) );
  XNOR2_X1 U6582 ( .A(n5173), .B(n5032), .ZN(n5174) );
  AOI22_X1 U6583 ( .A1(n9373), .A2(n5574), .B1(n9548), .B2(n5594), .ZN(n5175)
         );
  XNOR2_X1 U6584 ( .A(n5174), .B(n5175), .ZN(n7407) );
  INV_X1 U6585 ( .A(n5174), .ZN(n5176) );
  XNOR2_X1 U6586 ( .A(n5202), .B(SI_11_), .ZN(n5201) );
  XNOR2_X1 U6587 ( .A(n5204), .B(n5201), .ZN(n6338) );
  NAND2_X1 U6588 ( .A1(n6338), .A2(n8563), .ZN(n5182) );
  OAI21_X1 U6589 ( .B1(n5179), .B2(P1_IR_REG_10__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5180) );
  XNOR2_X1 U6590 ( .A(n5180), .B(P1_IR_REG_11__SCAN_IN), .ZN(n6648) );
  AOI22_X1 U6591 ( .A1(n5381), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n6290), .B2(
        n6648), .ZN(n5181) );
  NAND2_X1 U6592 ( .A1(n9451), .A2(n5598), .ZN(n5193) );
  NAND2_X1 U6593 ( .A1(n4272), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5191) );
  INV_X1 U6594 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n5183) );
  OR2_X1 U6595 ( .A1(n4273), .A2(n5183), .ZN(n5190) );
  AND2_X1 U6596 ( .A1(n5185), .A2(n5184), .ZN(n5186) );
  OR2_X1 U6597 ( .A1(n5186), .A2(n5213), .ZN(n9423) );
  OR2_X1 U6598 ( .A1(n5640), .A2(n9423), .ZN(n5189) );
  INV_X1 U6599 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n5187) );
  OR2_X1 U6600 ( .A1(n5241), .A2(n5187), .ZN(n5188) );
  NAND4_X1 U6601 ( .A1(n5191), .A2(n5190), .A3(n5189), .A4(n5188), .ZN(n8844)
         );
  NAND2_X1 U6602 ( .A1(n8844), .A2(n5574), .ZN(n5192) );
  NAND2_X1 U6603 ( .A1(n5193), .A2(n5192), .ZN(n5194) );
  XNOR2_X1 U6604 ( .A(n5194), .B(n7090), .ZN(n5196) );
  AND2_X1 U6605 ( .A1(n8844), .A2(n5594), .ZN(n5195) );
  AOI21_X1 U6606 ( .B1(n9451), .B2(n5574), .A(n5195), .ZN(n5197) );
  XNOR2_X1 U6607 ( .A(n5196), .B(n5197), .ZN(n7455) );
  INV_X1 U6608 ( .A(n5196), .ZN(n5199) );
  INV_X1 U6609 ( .A(n5197), .ZN(n5198) );
  NAND2_X1 U6610 ( .A1(n5199), .A2(n5198), .ZN(n5200) );
  INV_X1 U6611 ( .A(n5202), .ZN(n5203) );
  NAND2_X1 U6612 ( .A1(n5206), .A2(n5205), .ZN(n5230) );
  INV_X1 U6613 ( .A(n5206), .ZN(n5207) );
  NAND2_X1 U6614 ( .A1(n5207), .A2(SI_12_), .ZN(n5208) );
  NAND2_X1 U6615 ( .A1(n5230), .A2(n5208), .ZN(n5228) );
  XNOR2_X1 U6616 ( .A(n5229), .B(n5228), .ZN(n6549) );
  NAND2_X1 U6617 ( .A1(n6549), .A2(n8563), .ZN(n5212) );
  NAND2_X1 U6618 ( .A1(n5209), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5210) );
  XNOR2_X1 U6619 ( .A(n5210), .B(P1_IR_REG_12__SCAN_IN), .ZN(n6765) );
  AOI22_X1 U6620 ( .A1(n5381), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n6290), .B2(
        n6765), .ZN(n5211) );
  NAND2_X1 U6621 ( .A1(n9444), .A2(n5598), .ZN(n5221) );
  NAND2_X1 U6622 ( .A1(n5162), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n5219) );
  INV_X1 U6623 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n6641) );
  OR2_X1 U6624 ( .A1(n4273), .A2(n6641), .ZN(n5218) );
  NAND2_X1 U6625 ( .A1(n5213), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n5243) );
  OR2_X1 U6626 ( .A1(n5213), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n5214) );
  NAND2_X1 U6627 ( .A1(n5243), .A2(n5214), .ZN(n7488) );
  OR2_X1 U6628 ( .A1(n5640), .A2(n7488), .ZN(n5217) );
  INV_X1 U6629 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n5215) );
  OR2_X1 U6630 ( .A1(n4989), .A2(n5215), .ZN(n5216) );
  NAND4_X1 U6631 ( .A1(n5219), .A2(n5218), .A3(n5217), .A4(n5216), .ZN(n8843)
         );
  NAND2_X1 U6632 ( .A1(n8843), .A2(n5574), .ZN(n5220) );
  NAND2_X1 U6633 ( .A1(n5221), .A2(n5220), .ZN(n5222) );
  XNOR2_X1 U6634 ( .A(n5222), .B(n7090), .ZN(n5226) );
  AND2_X1 U6635 ( .A1(n8843), .A2(n5594), .ZN(n5223) );
  AOI21_X1 U6636 ( .B1(n9444), .B2(n5574), .A(n5223), .ZN(n5225) );
  XNOR2_X1 U6637 ( .A(n5226), .B(n5225), .ZN(n7485) );
  INV_X1 U6638 ( .A(n7485), .ZN(n5224) );
  NAND2_X1 U6639 ( .A1(n5226), .A2(n5225), .ZN(n5227) );
  MUX2_X1 U6640 ( .A(n6626), .B(n5232), .S(n5793), .Z(n5234) );
  NAND2_X1 U6641 ( .A1(n5234), .A2(n5233), .ZN(n5255) );
  INV_X1 U6642 ( .A(n5234), .ZN(n5235) );
  NAND2_X1 U6643 ( .A1(n5235), .A2(SI_13_), .ZN(n5236) );
  XNOR2_X1 U6644 ( .A(n5254), .B(n4841), .ZN(n6612) );
  NAND2_X1 U6645 ( .A1(n6612), .A2(n8563), .ZN(n5239) );
  NAND2_X1 U6646 ( .A1(n4292), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5237) );
  XNOR2_X1 U6647 ( .A(n5237), .B(P1_IR_REG_13__SCAN_IN), .ZN(n7141) );
  AOI22_X1 U6648 ( .A1(n5381), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n6290), .B2(
        n7141), .ZN(n5238) );
  NAND2_X1 U6649 ( .A1(n9407), .A2(n5598), .ZN(n5250) );
  NAND2_X1 U6650 ( .A1(n4272), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n5248) );
  INV_X1 U6651 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n6758) );
  OR2_X1 U6652 ( .A1(n4273), .A2(n6758), .ZN(n5247) );
  INV_X1 U6653 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n5240) );
  OR2_X1 U6654 ( .A1(n5241), .A2(n5240), .ZN(n5246) );
  NAND2_X1 U6655 ( .A1(n5243), .A2(n5242), .ZN(n5244) );
  NAND2_X1 U6656 ( .A1(n5264), .A2(n5244), .ZN(n9405) );
  OR2_X1 U6657 ( .A1(n5640), .A2(n9405), .ZN(n5245) );
  NAND4_X1 U6658 ( .A1(n5248), .A2(n5247), .A3(n5246), .A4(n5245), .ZN(n8842)
         );
  NAND2_X1 U6659 ( .A1(n8842), .A2(n5574), .ZN(n5249) );
  NAND2_X1 U6660 ( .A1(n5250), .A2(n5249), .ZN(n5251) );
  XNOR2_X1 U6661 ( .A(n5251), .B(n7090), .ZN(n7494) );
  AND2_X1 U6662 ( .A1(n8842), .A2(n5594), .ZN(n5252) );
  AOI21_X1 U6663 ( .B1(n9407), .B2(n5574), .A(n5252), .ZN(n7493) );
  AND2_X1 U6664 ( .A1(n7494), .A2(n7493), .ZN(n5253) );
  MUX2_X1 U6665 ( .A(n9885), .B(n5256), .S(n5793), .Z(n5277) );
  XNOR2_X1 U6666 ( .A(n5277), .B(SI_14_), .ZN(n5276) );
  XNOR2_X1 U6667 ( .A(n5280), .B(n5276), .ZN(n6623) );
  NAND2_X1 U6668 ( .A1(n6623), .A2(n8563), .ZN(n5263) );
  OR2_X1 U6669 ( .A1(n5257), .A2(n9330), .ZN(n5260) );
  INV_X1 U6670 ( .A(n5260), .ZN(n5258) );
  NAND2_X1 U6671 ( .A1(n5258), .A2(P1_IR_REG_14__SCAN_IN), .ZN(n5261) );
  NAND2_X1 U6672 ( .A1(n5260), .A2(n5259), .ZN(n5284) );
  AOI22_X1 U6673 ( .A1(n5381), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n6290), .B2(
        n9513), .ZN(n5262) );
  NAND2_X1 U6674 ( .A1(n8430), .A2(n5598), .ZN(n5271) );
  NAND2_X1 U6675 ( .A1(n5162), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n5269) );
  INV_X1 U6676 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n9884) );
  OR2_X1 U6677 ( .A1(n4989), .A2(n9884), .ZN(n5268) );
  INV_X1 U6678 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n9278) );
  OR2_X1 U6679 ( .A1(n4273), .A2(n9278), .ZN(n5267) );
  AND2_X1 U6680 ( .A1(n5264), .A2(n8425), .ZN(n5265) );
  OR2_X1 U6681 ( .A1(n5265), .A2(n5289), .ZN(n8428) );
  OR2_X1 U6682 ( .A1(n5640), .A2(n8428), .ZN(n5266) );
  NAND4_X1 U6683 ( .A1(n5269), .A2(n5268), .A3(n5267), .A4(n5266), .ZN(n9266)
         );
  NAND2_X1 U6684 ( .A1(n9266), .A2(n5574), .ZN(n5270) );
  NAND2_X1 U6685 ( .A1(n5271), .A2(n5270), .ZN(n5272) );
  XNOR2_X1 U6686 ( .A(n5272), .B(n5032), .ZN(n5275) );
  NAND2_X1 U6687 ( .A1(n8430), .A2(n5574), .ZN(n5274) );
  NAND2_X1 U6688 ( .A1(n9266), .A2(n5594), .ZN(n5273) );
  NAND2_X1 U6689 ( .A1(n5274), .A2(n5273), .ZN(n8424) );
  INV_X1 U6690 ( .A(n5276), .ZN(n5279) );
  INV_X1 U6691 ( .A(n5277), .ZN(n5278) );
  MUX2_X1 U6692 ( .A(n6775), .B(n9903), .S(n5793), .Z(n5281) );
  NAND2_X1 U6693 ( .A1(n5281), .A2(n9826), .ZN(n5301) );
  INV_X1 U6694 ( .A(n5281), .ZN(n5282) );
  NAND2_X1 U6695 ( .A1(n5282), .A2(SI_15_), .ZN(n5283) );
  NAND2_X1 U6696 ( .A1(n5301), .A2(n5283), .ZN(n5302) );
  XNOR2_X1 U6697 ( .A(n5303), .B(n5302), .ZN(n6774) );
  NAND2_X1 U6698 ( .A1(n6774), .A2(n8563), .ZN(n5288) );
  NAND2_X1 U6699 ( .A1(n5284), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5285) );
  INV_X1 U6700 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n9905) );
  XNOR2_X1 U6701 ( .A(n5285), .B(n9905), .ZN(n7290) );
  INV_X1 U6702 ( .A(n7290), .ZN(n5286) );
  AOI22_X1 U6703 ( .A1(n5381), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n6290), .B2(
        n5286), .ZN(n5287) );
  NAND2_X1 U6704 ( .A1(n9264), .A2(n5598), .ZN(n5296) );
  NAND2_X1 U6705 ( .A1(n4272), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n5294) );
  INV_X1 U6706 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n7144) );
  OR2_X1 U6707 ( .A1(n4273), .A2(n7144), .ZN(n5293) );
  INV_X1 U6708 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n9153) );
  OR2_X1 U6709 ( .A1(n5241), .A2(n9153), .ZN(n5292) );
  NOR2_X1 U6710 ( .A1(n5289), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n5290) );
  OR2_X1 U6711 ( .A1(n5312), .A2(n5290), .ZN(n9152) );
  OR2_X1 U6712 ( .A1(n5640), .A2(n9152), .ZN(n5291) );
  NAND4_X1 U6713 ( .A1(n5294), .A2(n5293), .A3(n5292), .A4(n5291), .ZN(n9255)
         );
  NAND2_X1 U6714 ( .A1(n9255), .A2(n5574), .ZN(n5295) );
  NAND2_X1 U6715 ( .A1(n5296), .A2(n5295), .ZN(n5297) );
  NAND2_X1 U6716 ( .A1(n9264), .A2(n5574), .ZN(n5299) );
  NAND2_X1 U6717 ( .A1(n9255), .A2(n5594), .ZN(n5298) );
  NAND2_X1 U6718 ( .A1(n5299), .A2(n5298), .ZN(n8543) );
  NAND2_X1 U6719 ( .A1(n8540), .A2(n8543), .ZN(n5300) );
  MUX2_X1 U6720 ( .A(n6812), .B(n6810), .S(n5793), .Z(n5305) );
  NAND2_X1 U6721 ( .A1(n5305), .A2(n5304), .ZN(n5327) );
  INV_X1 U6722 ( .A(n5305), .ZN(n5306) );
  NAND2_X1 U6723 ( .A1(n5306), .A2(SI_16_), .ZN(n5307) );
  XNOR2_X1 U6724 ( .A(n5326), .B(n5325), .ZN(n6809) );
  NAND2_X1 U6725 ( .A1(n6809), .A2(n8563), .ZN(n5311) );
  NAND2_X1 U6726 ( .A1(n5308), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5309) );
  XNOR2_X1 U6727 ( .A(n5309), .B(P1_IR_REG_16__SCAN_IN), .ZN(n8882) );
  AOI22_X1 U6728 ( .A1(n5381), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n6290), .B2(
        n8882), .ZN(n5310) );
  NAND2_X1 U6729 ( .A1(n9254), .A2(n5598), .ZN(n5319) );
  NAND2_X1 U6730 ( .A1(n5585), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n5317) );
  INV_X1 U6731 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n9134) );
  OR2_X1 U6732 ( .A1(n5241), .A2(n9134), .ZN(n5316) );
  OR2_X1 U6733 ( .A1(n5312), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n5313) );
  NAND2_X1 U6734 ( .A1(n5332), .A2(n5313), .ZN(n9133) );
  OR2_X1 U6735 ( .A1(n5640), .A2(n9133), .ZN(n5315) );
  INV_X1 U6736 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n9320) );
  OR2_X1 U6737 ( .A1(n4989), .A2(n9320), .ZN(n5314) );
  NAND4_X1 U6738 ( .A1(n5317), .A2(n5316), .A3(n5315), .A4(n5314), .ZN(n9265)
         );
  NAND2_X1 U6739 ( .A1(n9265), .A2(n5574), .ZN(n5318) );
  NAND2_X1 U6740 ( .A1(n5319), .A2(n5318), .ZN(n5320) );
  XNOR2_X1 U6741 ( .A(n5320), .B(n7090), .ZN(n5323) );
  AND2_X1 U6742 ( .A1(n9265), .A2(n5594), .ZN(n5321) );
  AOI21_X1 U6743 ( .B1(n9254), .B2(n5574), .A(n5321), .ZN(n5322) );
  XNOR2_X1 U6744 ( .A(n5323), .B(n5322), .ZN(n8466) );
  NAND2_X1 U6745 ( .A1(n5323), .A2(n5322), .ZN(n5324) );
  NAND2_X1 U6746 ( .A1(n5326), .A2(n5325), .ZN(n5328) );
  MUX2_X1 U6747 ( .A(n6839), .B(n5329), .S(n5793), .Z(n5348) );
  XNOR2_X1 U6748 ( .A(n5348), .B(SI_17_), .ZN(n5347) );
  XNOR2_X1 U6749 ( .A(n5352), .B(n5347), .ZN(n6826) );
  NAND2_X1 U6750 ( .A1(n4339), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5354) );
  XNOR2_X1 U6751 ( .A(n5354), .B(P1_IR_REG_17__SCAN_IN), .ZN(n8897) );
  AOI22_X1 U6752 ( .A1(n5381), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n6290), .B2(
        n8897), .ZN(n5330) );
  NAND2_X1 U6753 ( .A1(n9126), .A2(n5598), .ZN(n5339) );
  NAND2_X1 U6754 ( .A1(n5162), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n5337) );
  INV_X1 U6755 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9252) );
  OR2_X1 U6756 ( .A1(n4273), .A2(n9252), .ZN(n5336) );
  INV_X1 U6757 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n5331) );
  NAND2_X1 U6758 ( .A1(n5332), .A2(n5331), .ZN(n5333) );
  NAND2_X1 U6759 ( .A1(n5360), .A2(n5333), .ZN(n9114) );
  OR2_X1 U6760 ( .A1(n5640), .A2(n9114), .ZN(n5335) );
  INV_X1 U6761 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n9316) );
  OR2_X1 U6762 ( .A1(n4989), .A2(n9316), .ZN(n5334) );
  NAND4_X1 U6763 ( .A1(n5337), .A2(n5336), .A3(n5335), .A4(n5334), .ZN(n9256)
         );
  NAND2_X1 U6764 ( .A1(n9256), .A2(n5574), .ZN(n5338) );
  NAND2_X1 U6765 ( .A1(n5339), .A2(n5338), .ZN(n5340) );
  XNOR2_X1 U6766 ( .A(n5340), .B(n5032), .ZN(n5342) );
  AND2_X1 U6767 ( .A1(n9256), .A2(n5594), .ZN(n5341) );
  AOI21_X1 U6768 ( .B1(n9126), .B2(n5574), .A(n5341), .ZN(n5343) );
  XNOR2_X1 U6769 ( .A(n5342), .B(n5343), .ZN(n8483) );
  NAND2_X1 U6770 ( .A1(n8484), .A2(n8483), .ZN(n5346) );
  INV_X1 U6771 ( .A(n5342), .ZN(n5344) );
  NAND2_X1 U6772 ( .A1(n5344), .A2(n5343), .ZN(n5345) );
  INV_X1 U6773 ( .A(n5347), .ZN(n5351) );
  INV_X1 U6774 ( .A(n5348), .ZN(n5349) );
  NAND2_X1 U6775 ( .A1(n5349), .A2(SI_17_), .ZN(n5350) );
  MUX2_X1 U6776 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n5793), .Z(n5376) );
  XNOR2_X1 U6777 ( .A(n5376), .B(SI_18_), .ZN(n5373) );
  XNOR2_X1 U6778 ( .A(n5375), .B(n5373), .ZN(n6948) );
  NAND2_X1 U6779 ( .A1(n6948), .A2(n8563), .ZN(n5358) );
  NAND2_X1 U6780 ( .A1(n5354), .A2(n5353), .ZN(n5355) );
  NAND2_X1 U6781 ( .A1(n5355), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5356) );
  XNOR2_X1 U6782 ( .A(n5356), .B(P1_IR_REG_18__SCAN_IN), .ZN(n8898) );
  AOI22_X1 U6783 ( .A1(n5381), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n6290), .B2(
        n8898), .ZN(n5357) );
  NAND2_X1 U6784 ( .A1(n9241), .A2(n5598), .ZN(n5367) );
  NAND2_X1 U6785 ( .A1(n4272), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n5365) );
  INV_X1 U6786 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9851) );
  OR2_X1 U6787 ( .A1(n4273), .A2(n9851), .ZN(n5364) );
  INV_X1 U6788 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n5359) );
  AND2_X1 U6789 ( .A1(n5360), .A2(n5359), .ZN(n5361) );
  OR2_X1 U6790 ( .A1(n5361), .A2(n5384), .ZN(n9100) );
  OR2_X1 U6791 ( .A1(n5640), .A2(n9100), .ZN(n5363) );
  INV_X1 U6792 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9101) );
  OR2_X1 U6793 ( .A1(n5241), .A2(n9101), .ZN(n5362) );
  NAND4_X1 U6794 ( .A1(n5365), .A2(n5364), .A3(n5363), .A4(n5362), .ZN(n9233)
         );
  NAND2_X1 U6795 ( .A1(n9233), .A2(n5574), .ZN(n5366) );
  NAND2_X1 U6796 ( .A1(n5367), .A2(n5366), .ZN(n5368) );
  XNOR2_X1 U6797 ( .A(n5368), .B(n7090), .ZN(n5371) );
  NAND2_X1 U6798 ( .A1(n9241), .A2(n5574), .ZN(n5370) );
  NAND2_X1 U6799 ( .A1(n9233), .A2(n5594), .ZN(n5369) );
  NAND2_X1 U6800 ( .A1(n5370), .A2(n5369), .ZN(n8522) );
  INV_X1 U6801 ( .A(n5371), .ZN(n5372) );
  INV_X1 U6802 ( .A(n5373), .ZN(n5374) );
  MUX2_X1 U6803 ( .A(n7022), .B(n7024), .S(n5793), .Z(n5378) );
  INV_X1 U6804 ( .A(SI_19_), .ZN(n5377) );
  NAND2_X1 U6805 ( .A1(n5378), .A2(n5377), .ZN(n5401) );
  INV_X1 U6806 ( .A(n5378), .ZN(n5379) );
  NAND2_X1 U6807 ( .A1(n5379), .A2(SI_19_), .ZN(n5380) );
  NAND2_X1 U6808 ( .A1(n5401), .A2(n5380), .ZN(n5399) );
  XNOR2_X1 U6809 ( .A(n5400), .B(n5399), .ZN(n7021) );
  NAND2_X1 U6810 ( .A1(n7021), .A2(n8563), .ZN(n5383) );
  AOI22_X1 U6811 ( .A1(n5381), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n9074), .B2(
        n6290), .ZN(n5382) );
  NAND2_X1 U6812 ( .A1(n9231), .A2(n5598), .ZN(n5391) );
  NOR2_X1 U6813 ( .A1(n5384), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n5385) );
  OR2_X1 U6814 ( .A1(n5409), .A2(n5385), .ZN(n9083) );
  OR2_X1 U6815 ( .A1(n9083), .A2(n5640), .ZN(n5389) );
  INV_X1 U6816 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n9308) );
  OR2_X1 U6817 ( .A1(n4989), .A2(n9308), .ZN(n5388) );
  INV_X1 U6818 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n9239) );
  OR2_X1 U6819 ( .A1(n4273), .A2(n9239), .ZN(n5387) );
  INV_X1 U6820 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n9084) );
  OR2_X1 U6821 ( .A1(n5241), .A2(n9084), .ZN(n5386) );
  NAND4_X1 U6822 ( .A1(n5389), .A2(n5388), .A3(n5387), .A4(n5386), .ZN(n9242)
         );
  NAND2_X1 U6823 ( .A1(n9242), .A2(n5574), .ZN(n5390) );
  NAND2_X1 U6824 ( .A1(n5391), .A2(n5390), .ZN(n5392) );
  XNOR2_X1 U6825 ( .A(n5392), .B(n7090), .ZN(n5397) );
  AND2_X1 U6826 ( .A1(n9242), .A2(n5594), .ZN(n5393) );
  AOI21_X1 U6827 ( .B1(n9231), .B2(n5574), .A(n5393), .ZN(n5396) );
  XNOR2_X1 U6828 ( .A(n5397), .B(n5396), .ZN(n8444) );
  INV_X1 U6829 ( .A(n8444), .ZN(n5394) );
  NAND2_X1 U6830 ( .A1(n5397), .A2(n5396), .ZN(n5398) );
  MUX2_X1 U6831 ( .A(n7163), .B(n7152), .S(n5793), .Z(n5404) );
  INV_X1 U6832 ( .A(SI_20_), .ZN(n5403) );
  NAND2_X1 U6833 ( .A1(n5404), .A2(n5403), .ZN(n5428) );
  INV_X1 U6834 ( .A(n5404), .ZN(n5405) );
  NAND2_X1 U6835 ( .A1(n5405), .A2(SI_20_), .ZN(n5406) );
  XNOR2_X1 U6836 ( .A(n5427), .B(n5426), .ZN(n7150) );
  NAND2_X1 U6837 ( .A1(n7150), .A2(n8563), .ZN(n5408) );
  OR2_X1 U6838 ( .A1(n5000), .A2(n7152), .ZN(n5407) );
  NAND2_X1 U6839 ( .A1(n9228), .A2(n5598), .ZN(n5419) );
  NAND2_X1 U6840 ( .A1(n5409), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n5432) );
  OR2_X1 U6841 ( .A1(n5409), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n5410) );
  AND2_X1 U6842 ( .A1(n5432), .A2(n5410), .ZN(n9072) );
  NAND2_X1 U6843 ( .A1(n5495), .A2(n9072), .ZN(n5417) );
  INV_X1 U6844 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n5411) );
  OR2_X1 U6845 ( .A1(n4989), .A2(n5411), .ZN(n5416) );
  INV_X1 U6846 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n5412) );
  OR2_X1 U6847 ( .A1(n4273), .A2(n5412), .ZN(n5415) );
  INV_X1 U6848 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n5413) );
  OR2_X1 U6849 ( .A1(n5241), .A2(n5413), .ZN(n5414) );
  NAND4_X1 U6850 ( .A1(n5417), .A2(n5416), .A3(n5415), .A4(n5414), .ZN(n9232)
         );
  NAND2_X1 U6851 ( .A1(n9232), .A2(n5574), .ZN(n5418) );
  NAND2_X1 U6852 ( .A1(n5419), .A2(n5418), .ZN(n5420) );
  XNOR2_X1 U6853 ( .A(n5420), .B(n5032), .ZN(n5422) );
  AND2_X1 U6854 ( .A1(n9232), .A2(n5594), .ZN(n5421) );
  AOI21_X1 U6855 ( .B1(n9228), .B2(n5574), .A(n5421), .ZN(n5423) );
  XNOR2_X1 U6856 ( .A(n5422), .B(n5423), .ZN(n8498) );
  INV_X1 U6857 ( .A(n5422), .ZN(n5424) );
  NAND2_X1 U6858 ( .A1(n5424), .A2(n5423), .ZN(n5425) );
  MUX2_X1 U6859 ( .A(n7251), .B(n7249), .S(n5793), .Z(n5448) );
  XNOR2_X1 U6860 ( .A(n5448), .B(SI_21_), .ZN(n5447) );
  XNOR2_X1 U6861 ( .A(n5446), .B(n5447), .ZN(n7248) );
  NAND2_X1 U6862 ( .A1(n7248), .A2(n8563), .ZN(n5430) );
  OR2_X1 U6863 ( .A1(n5000), .A2(n7249), .ZN(n5429) );
  NAND2_X1 U6864 ( .A1(n8456), .A2(n5598), .ZN(n5439) );
  INV_X1 U6865 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n5431) );
  NAND2_X1 U6866 ( .A1(n5432), .A2(n5431), .ZN(n5433) );
  NAND2_X1 U6867 ( .A1(n5458), .A2(n5433), .ZN(n9055) );
  NOR2_X1 U6868 ( .A1(n9055), .A2(n5640), .ZN(n5437) );
  INV_X1 U6869 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n9836) );
  NAND2_X1 U6870 ( .A1(n5585), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n5434) );
  OAI21_X1 U6871 ( .B1(n9836), .B2(n4989), .A(n5434), .ZN(n5436) );
  INV_X1 U6872 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n9056) );
  NOR2_X1 U6873 ( .A1(n5241), .A2(n9056), .ZN(n5435) );
  NAND2_X1 U6874 ( .A1(n9038), .A2(n5574), .ZN(n5438) );
  NAND2_X1 U6875 ( .A1(n5439), .A2(n5438), .ZN(n5440) );
  XNOR2_X1 U6876 ( .A(n5440), .B(n5032), .ZN(n5441) );
  AOI22_X1 U6877 ( .A1(n8456), .A2(n5574), .B1(n5594), .B2(n9038), .ZN(n5442)
         );
  XNOR2_X1 U6878 ( .A(n5441), .B(n5442), .ZN(n8452) );
  INV_X1 U6879 ( .A(n5441), .ZN(n5443) );
  NAND2_X1 U6880 ( .A1(n5443), .A2(n5442), .ZN(n5444) );
  INV_X1 U6881 ( .A(n5448), .ZN(n5449) );
  NAND2_X1 U6882 ( .A1(n5449), .A2(SI_21_), .ZN(n5450) );
  INV_X1 U6883 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7533) );
  MUX2_X1 U6884 ( .A(n7533), .B(n7311), .S(n5793), .Z(n5453) );
  NAND2_X1 U6885 ( .A1(n5453), .A2(n5452), .ZN(n5470) );
  INV_X1 U6886 ( .A(n5453), .ZN(n5454) );
  NAND2_X1 U6887 ( .A1(n5454), .A2(SI_22_), .ZN(n5455) );
  NAND2_X1 U6888 ( .A1(n5470), .A2(n5455), .ZN(n5468) );
  XNOR2_X1 U6889 ( .A(n5469), .B(n5468), .ZN(n7310) );
  NAND2_X1 U6890 ( .A1(n7310), .A2(n8563), .ZN(n5457) );
  OR2_X1 U6891 ( .A1(n5000), .A2(n7311), .ZN(n5456) );
  INV_X1 U6892 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n8513) );
  NAND2_X1 U6893 ( .A1(n5458), .A2(n8513), .ZN(n5459) );
  NAND2_X1 U6894 ( .A1(n5478), .A2(n5459), .ZN(n9043) );
  AOI22_X1 U6895 ( .A1(n5585), .A2(P1_REG1_REG_22__SCAN_IN), .B1(n4272), .B2(
        P1_REG0_REG_22__SCAN_IN), .ZN(n5461) );
  NAND2_X1 U6896 ( .A1(n5162), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n5460) );
  OAI211_X1 U6897 ( .C1(n9043), .C2(n5640), .A(n5461), .B(n5460), .ZN(n9218)
         );
  AND2_X1 U6898 ( .A1(n9218), .A2(n5594), .ZN(n5462) );
  AOI21_X1 U6899 ( .B1(n9215), .B2(n4982), .A(n5462), .ZN(n5465) );
  NAND2_X1 U6900 ( .A1(n5464), .A2(n5465), .ZN(n8511) );
  AOI22_X1 U6901 ( .A1(n9215), .A2(n5598), .B1(n5574), .B2(n9218), .ZN(n5463)
         );
  XOR2_X1 U6902 ( .A(n5032), .B(n5463), .Z(n8509) );
  NAND2_X1 U6903 ( .A1(n8511), .A2(n8509), .ZN(n8506) );
  INV_X1 U6904 ( .A(n5464), .ZN(n5467) );
  INV_X1 U6905 ( .A(n5465), .ZN(n5466) );
  NAND2_X1 U6906 ( .A1(n8506), .A2(n8507), .ZN(n8505) );
  INV_X1 U6907 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n5471) );
  INV_X1 U6908 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n7376) );
  MUX2_X1 U6909 ( .A(n5471), .B(n7376), .S(n5793), .Z(n5473) );
  INV_X1 U6910 ( .A(SI_23_), .ZN(n5472) );
  NAND2_X1 U6911 ( .A1(n5473), .A2(n5472), .ZN(n5490) );
  INV_X1 U6912 ( .A(n5473), .ZN(n5474) );
  NAND2_X1 U6913 ( .A1(n5474), .A2(SI_23_), .ZN(n5475) );
  XNOR2_X1 U6914 ( .A(n5489), .B(n5488), .ZN(n7373) );
  NAND2_X1 U6915 ( .A1(n7373), .A2(n8563), .ZN(n5477) );
  OR2_X1 U6916 ( .A1(n5000), .A2(n7376), .ZN(n5476) );
  INV_X1 U6917 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n8436) );
  AND2_X1 U6918 ( .A1(n5478), .A2(n8436), .ZN(n5479) );
  OR2_X1 U6919 ( .A1(n5479), .A2(n5493), .ZN(n9027) );
  INV_X1 U6920 ( .A(n9027), .ZN(n5484) );
  INV_X1 U6921 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n5482) );
  NAND2_X1 U6922 ( .A1(n5585), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n5481) );
  NAND2_X1 U6923 ( .A1(n4272), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n5480) );
  OAI211_X1 U6924 ( .C1(n5241), .C2(n5482), .A(n5481), .B(n5480), .ZN(n5483)
         );
  OAI22_X1 U6925 ( .A1(n5731), .A2(n5485), .B1(n9201), .B2(n5577), .ZN(n5486)
         );
  XNOR2_X1 U6926 ( .A(n5486), .B(n5032), .ZN(n5487) );
  AOI22_X1 U6927 ( .A1(n9210), .A2(n5574), .B1(n5594), .B2(n9039), .ZN(n8434)
         );
  NAND2_X1 U6928 ( .A1(n8505), .A2(n5487), .ZN(n8433) );
  INV_X1 U6929 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7403) );
  INV_X1 U6930 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7401) );
  MUX2_X1 U6931 ( .A(n7403), .B(n7401), .S(n5793), .Z(n5512) );
  XNOR2_X1 U6932 ( .A(n5512), .B(SI_24_), .ZN(n5509) );
  XNOR2_X1 U6933 ( .A(n5511), .B(n5509), .ZN(n7400) );
  NAND2_X1 U6934 ( .A1(n7400), .A2(n8563), .ZN(n5492) );
  OR2_X1 U6935 ( .A1(n5000), .A2(n7401), .ZN(n5491) );
  OR2_X1 U6936 ( .A1(n5493), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n5494) );
  NAND2_X1 U6937 ( .A1(n5493), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n5522) );
  AND2_X1 U6938 ( .A1(n5494), .A2(n5522), .ZN(n9010) );
  NAND2_X1 U6939 ( .A1(n9010), .A2(n5495), .ZN(n5501) );
  INV_X1 U6940 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n5498) );
  NAND2_X1 U6941 ( .A1(n4272), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n5497) );
  NAND2_X1 U6942 ( .A1(n5162), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n5496) );
  OAI211_X1 U6943 ( .C1(n4273), .C2(n5498), .A(n5497), .B(n5496), .ZN(n5499)
         );
  INV_X1 U6944 ( .A(n5499), .ZN(n5500) );
  AND2_X1 U6945 ( .A1(n9023), .A2(n5594), .ZN(n5502) );
  AOI21_X1 U6946 ( .B1(n9204), .B2(n5574), .A(n5502), .ZN(n5506) );
  NAND2_X1 U6947 ( .A1(n9204), .A2(n5598), .ZN(n5504) );
  NAND2_X1 U6948 ( .A1(n9023), .A2(n5574), .ZN(n5503) );
  NAND2_X1 U6949 ( .A1(n5504), .A2(n5503), .ZN(n5505) );
  XNOR2_X1 U6950 ( .A(n5505), .B(n5032), .ZN(n5507) );
  XOR2_X1 U6951 ( .A(n5506), .B(n5507), .Z(n8491) );
  INV_X1 U6952 ( .A(n5506), .ZN(n5508) );
  INV_X1 U6953 ( .A(n5509), .ZN(n5510) );
  INV_X1 U6954 ( .A(n5512), .ZN(n5513) );
  NAND2_X1 U6955 ( .A1(n5513), .A2(SI_24_), .ZN(n5514) );
  INV_X1 U6956 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7479) );
  MUX2_X1 U6957 ( .A(n9829), .B(n7479), .S(n5793), .Z(n5517) );
  INV_X1 U6958 ( .A(SI_25_), .ZN(n5516) );
  NAND2_X1 U6959 ( .A1(n5517), .A2(n5516), .ZN(n5533) );
  INV_X1 U6960 ( .A(n5517), .ZN(n5518) );
  NAND2_X1 U6961 ( .A1(n5518), .A2(SI_25_), .ZN(n5519) );
  NAND2_X1 U6962 ( .A1(n5533), .A2(n5519), .ZN(n5534) );
  XNOR2_X1 U6963 ( .A(n5535), .B(n5534), .ZN(n7477) );
  NAND2_X1 U6964 ( .A1(n7477), .A2(n8563), .ZN(n5521) );
  OR2_X1 U6965 ( .A1(n5000), .A2(n7479), .ZN(n5520) );
  NAND2_X1 U6966 ( .A1(n8990), .A2(n5598), .ZN(n5528) );
  NAND2_X1 U6967 ( .A1(n5585), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n5526) );
  INV_X1 U6968 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n8992) );
  OR2_X1 U6969 ( .A1(n5241), .A2(n8992), .ZN(n5525) );
  XNOR2_X1 U6970 ( .A(P1_REG3_REG_25__SCAN_IN), .B(n5542), .ZN(n8991) );
  OR2_X1 U6971 ( .A1(n5640), .A2(n8991), .ZN(n5524) );
  INV_X1 U6972 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n9297) );
  OR2_X1 U6973 ( .A1(n4989), .A2(n9297), .ZN(n5523) );
  NAND4_X1 U6974 ( .A1(n5526), .A2(n5525), .A3(n5524), .A4(n5523), .ZN(n9013)
         );
  NAND2_X1 U6975 ( .A1(n9013), .A2(n4982), .ZN(n5527) );
  NAND2_X1 U6976 ( .A1(n5528), .A2(n5527), .ZN(n5529) );
  XNOR2_X1 U6977 ( .A(n5529), .B(n5032), .ZN(n5530) );
  AOI22_X1 U6978 ( .A1(n8990), .A2(n5574), .B1(n5594), .B2(n9013), .ZN(n5531)
         );
  XNOR2_X1 U6979 ( .A(n5530), .B(n5531), .ZN(n8459) );
  INV_X1 U6980 ( .A(n5530), .ZN(n5532) );
  INV_X1 U6981 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n8418) );
  MUX2_X1 U6982 ( .A(n8418), .B(n9341), .S(n5793), .Z(n5537) );
  INV_X1 U6983 ( .A(SI_26_), .ZN(n5536) );
  NAND2_X1 U6984 ( .A1(n5537), .A2(n5536), .ZN(n5558) );
  INV_X1 U6985 ( .A(n5537), .ZN(n5538) );
  NAND2_X1 U6986 ( .A1(n5538), .A2(SI_26_), .ZN(n5539) );
  XNOR2_X1 U6987 ( .A(n5557), .B(n5556), .ZN(n8416) );
  NAND2_X1 U6988 ( .A1(n8416), .A2(n8563), .ZN(n5541) );
  OR2_X1 U6989 ( .A1(n5000), .A2(n9341), .ZN(n5540) );
  NAND2_X1 U6990 ( .A1(n8973), .A2(n5598), .ZN(n5551) );
  NAND2_X1 U6991 ( .A1(n4272), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n5549) );
  INV_X1 U6992 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n9192) );
  OR2_X1 U6993 ( .A1(n4273), .A2(n9192), .ZN(n5548) );
  NAND3_X1 U6994 ( .A1(P1_REG3_REG_25__SCAN_IN), .A2(P1_REG3_REG_26__SCAN_IN), 
        .A3(n5542), .ZN(n5568) );
  INV_X1 U6995 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n5544) );
  NAND2_X1 U6996 ( .A1(P1_REG3_REG_25__SCAN_IN), .A2(n5542), .ZN(n5543) );
  NAND2_X1 U6997 ( .A1(n5544), .A2(n5543), .ZN(n5545) );
  NAND2_X1 U6998 ( .A1(n5568), .A2(n5545), .ZN(n8974) );
  OR2_X1 U6999 ( .A1(n5640), .A2(n8974), .ZN(n5547) );
  INV_X1 U7000 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n8975) );
  OR2_X1 U7001 ( .A1(n5241), .A2(n8975), .ZN(n5546) );
  NAND4_X1 U7002 ( .A1(n5549), .A2(n5548), .A3(n5547), .A4(n5546), .ZN(n8999)
         );
  NAND2_X1 U7003 ( .A1(n8999), .A2(n4982), .ZN(n5550) );
  NAND2_X1 U7004 ( .A1(n5551), .A2(n5550), .ZN(n5552) );
  XNOR2_X1 U7005 ( .A(n5552), .B(n7090), .ZN(n5555) );
  AND2_X1 U7006 ( .A1(n8999), .A2(n5594), .ZN(n5553) );
  AOI21_X1 U7007 ( .B1(n8973), .B2(n4982), .A(n5553), .ZN(n5554) );
  NOR2_X1 U7008 ( .A1(n5555), .A2(n5554), .ZN(n8531) );
  NAND2_X1 U7009 ( .A1(n5555), .A2(n5554), .ZN(n8529) );
  OAI21_X2 U7010 ( .B1(n8533), .B2(n8531), .A(n8529), .ZN(n6276) );
  NAND2_X1 U7011 ( .A1(n5557), .A2(n5556), .ZN(n5559) );
  INV_X1 U7012 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n8415) );
  INV_X1 U7013 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n9339) );
  INV_X1 U7014 ( .A(SI_27_), .ZN(n5560) );
  NAND2_X1 U7015 ( .A1(n5561), .A2(n5560), .ZN(n5582) );
  INV_X1 U7016 ( .A(n5561), .ZN(n5562) );
  NAND2_X1 U7017 ( .A1(n5562), .A2(SI_27_), .ZN(n5563) );
  NAND2_X1 U7018 ( .A1(n8412), .A2(n8563), .ZN(n5565) );
  OR2_X1 U7019 ( .A1(n5000), .A2(n9339), .ZN(n5564) );
  NAND2_X1 U7020 ( .A1(n5585), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n5573) );
  INV_X1 U7021 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n5566) );
  OR2_X1 U7022 ( .A1(n4989), .A2(n5566), .ZN(n5572) );
  INV_X1 U7023 ( .A(n5568), .ZN(n5567) );
  NAND2_X1 U7024 ( .A1(n5567), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n5588) );
  INV_X1 U7025 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n9880) );
  NAND2_X1 U7026 ( .A1(n5568), .A2(n9880), .ZN(n5569) );
  NAND2_X1 U7027 ( .A1(n5588), .A2(n5569), .ZN(n8959) );
  OR2_X1 U7028 ( .A1(n5640), .A2(n8959), .ZN(n5571) );
  INV_X1 U7029 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n8960) );
  OR2_X1 U7030 ( .A1(n5241), .A2(n8960), .ZN(n5570) );
  NAND4_X1 U7031 ( .A1(n5573), .A2(n5572), .A3(n5571), .A4(n5570), .ZN(n9176)
         );
  AOI22_X1 U7032 ( .A1(n9186), .A2(n4900), .B1(n5574), .B2(n9176), .ZN(n5575)
         );
  XOR2_X1 U7033 ( .A(n5032), .B(n5575), .Z(n5579) );
  INV_X1 U7034 ( .A(n5594), .ZN(n5576) );
  OAI22_X1 U7035 ( .A1(n4537), .A2(n5577), .B1(n5697), .B2(n5576), .ZN(n5578)
         );
  NOR2_X1 U7036 ( .A1(n5579), .A2(n5578), .ZN(n5628) );
  AOI21_X1 U7037 ( .B1(n5579), .B2(n5578), .A(n5628), .ZN(n6275) );
  NAND2_X1 U7038 ( .A1(n6276), .A2(n6275), .ZN(n6277) );
  INV_X1 U7039 ( .A(n6277), .ZN(n5624) );
  INV_X1 U7040 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n9336) );
  INV_X1 U7041 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n7529) );
  MUX2_X1 U7042 ( .A(n9336), .B(n7529), .S(n7698), .Z(n5704) );
  XNOR2_X1 U7043 ( .A(n5704), .B(SI_28_), .ZN(n5701) );
  NAND2_X1 U7044 ( .A1(n7527), .A2(n8563), .ZN(n5584) );
  OR2_X1 U7045 ( .A1(n5000), .A2(n9336), .ZN(n5583) );
  NAND2_X1 U7046 ( .A1(n8945), .A2(n4982), .ZN(n5596) );
  NAND2_X1 U7047 ( .A1(n5585), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n5593) );
  INV_X1 U7048 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n9289) );
  OR2_X1 U7049 ( .A1(n4989), .A2(n9289), .ZN(n5592) );
  INV_X1 U7050 ( .A(n5588), .ZN(n5586) );
  NAND2_X1 U7051 ( .A1(n5586), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n8923) );
  INV_X1 U7052 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n5587) );
  NAND2_X1 U7053 ( .A1(n5588), .A2(n5587), .ZN(n5589) );
  NAND2_X1 U7054 ( .A1(n8923), .A2(n5589), .ZN(n8946) );
  OR2_X1 U7055 ( .A1(n5640), .A2(n8946), .ZN(n5591) );
  INV_X1 U7056 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n8947) );
  OR2_X1 U7057 ( .A1(n5241), .A2(n8947), .ZN(n5590) );
  NAND4_X1 U7058 ( .A1(n5593), .A2(n5592), .A3(n5591), .A4(n5590), .ZN(n8965)
         );
  NAND2_X1 U7059 ( .A1(n8965), .A2(n5594), .ZN(n5595) );
  NAND2_X1 U7060 ( .A1(n5596), .A2(n5595), .ZN(n5597) );
  XNOR2_X1 U7061 ( .A(n5597), .B(n5032), .ZN(n5600) );
  AOI22_X1 U7062 ( .A1(n8945), .A2(n5598), .B1(n5574), .B2(n8965), .ZN(n5599)
         );
  XNOR2_X1 U7063 ( .A(n5600), .B(n5599), .ZN(n5627) );
  NAND2_X1 U7064 ( .A1(n7478), .A2(P1_B_REG_SCAN_IN), .ZN(n5602) );
  MUX2_X1 U7065 ( .A(n5602), .B(P1_B_REG_SCAN_IN), .S(n5616), .Z(n5603) );
  INV_X1 U7066 ( .A(n9576), .ZN(n5613) );
  INV_X1 U7067 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n9811) );
  INV_X1 U7068 ( .A(n5601), .ZN(n9344) );
  AND2_X1 U7069 ( .A1(n9344), .A2(n7478), .ZN(n5604) );
  AOI21_X1 U7070 ( .B1(n5613), .B2(n9811), .A(n5604), .ZN(n6314) );
  NOR4_X1 U7071 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_17__SCAN_IN), .A3(
        P1_D_REG_18__SCAN_IN), .A4(P1_D_REG_19__SCAN_IN), .ZN(n5608) );
  NOR4_X1 U7072 ( .A1(P1_D_REG_14__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_13__SCAN_IN), .A4(P1_D_REG_15__SCAN_IN), .ZN(n5607) );
  NOR4_X1 U7073 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n5606) );
  NOR4_X1 U7074 ( .A1(P1_D_REG_21__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n5605) );
  NAND4_X1 U7075 ( .A1(n5608), .A2(n5607), .A3(n5606), .A4(n5605), .ZN(n5615)
         );
  NOR2_X1 U7076 ( .A1(P1_D_REG_20__SCAN_IN), .A2(P1_D_REG_12__SCAN_IN), .ZN(
        n5612) );
  NOR4_X1 U7077 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_22__SCAN_IN), .A4(P1_D_REG_8__SCAN_IN), .ZN(n5611) );
  NOR4_X1 U7078 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_9__SCAN_IN), .A4(P1_D_REG_10__SCAN_IN), .ZN(n5610) );
  NOR4_X1 U7079 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n5609) );
  NAND4_X1 U7080 ( .A1(n5612), .A2(n5611), .A3(n5610), .A4(n5609), .ZN(n5614)
         );
  OAI21_X1 U7081 ( .B1(n5615), .B2(n5614), .A(n5613), .ZN(n5749) );
  NAND2_X1 U7082 ( .A1(n6314), .A2(n5749), .ZN(n7087) );
  OR2_X1 U7083 ( .A1(n7087), .A2(n7181), .ZN(n5631) );
  NAND2_X1 U7084 ( .A1(n5617), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5618) );
  AND2_X1 U7085 ( .A1(n7374), .A2(P1_STATE_REG_SCAN_IN), .ZN(n5619) );
  NOR2_X1 U7086 ( .A1(n5631), .A2(n8556), .ZN(n5635) );
  AND2_X1 U7087 ( .A1(n9612), .A2(n8680), .ZN(n5622) );
  NAND2_X1 U7088 ( .A1(n5624), .A2(n5623), .ZN(n5652) );
  INV_X1 U7089 ( .A(n5628), .ZN(n5626) );
  INV_X1 U7090 ( .A(n5627), .ZN(n5625) );
  NAND4_X1 U7091 ( .A1(n6277), .A2(n8475), .A3(n5626), .A4(n5625), .ZN(n5651)
         );
  NAND3_X1 U7092 ( .A1(n5631), .A2(n9577), .A3(n4348), .ZN(n6679) );
  OR2_X1 U7093 ( .A1(n8680), .A2(n8832), .ZN(n5630) );
  NOR2_X1 U7094 ( .A1(n7088), .A2(n9612), .ZN(n5629) );
  AND3_X1 U7095 ( .A1(n5630), .A2(n6287), .A3(n7374), .ZN(n5632) );
  NAND2_X1 U7096 ( .A1(n5631), .A2(n9612), .ZN(n6677) );
  NAND2_X1 U7097 ( .A1(n5632), .A2(n6677), .ZN(n5633) );
  NAND2_X1 U7098 ( .A1(n5633), .A2(P1_STATE_REG_SCAN_IN), .ZN(n5634) );
  OR2_X1 U7099 ( .A1(n5712), .A2(n4916), .ZN(n8557) );
  INV_X1 U7100 ( .A(n8557), .ZN(n7091) );
  AND2_X1 U7101 ( .A1(n5635), .A2(n7091), .ZN(n5638) );
  INV_X1 U7102 ( .A(n5637), .ZN(n5741) );
  NAND2_X1 U7103 ( .A1(n5638), .A2(n5741), .ZN(n8545) );
  AOI22_X1 U7104 ( .A1(n8534), .A2(n9176), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3084), .ZN(n5646) );
  INV_X1 U7105 ( .A(n5638), .ZN(n5639) );
  INV_X1 U7106 ( .A(n8523), .ZN(n7411) );
  NAND2_X1 U7107 ( .A1(n5162), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n5644) );
  INV_X1 U7108 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n9813) );
  OR2_X1 U7109 ( .A1(n4273), .A2(n9813), .ZN(n5643) );
  INV_X1 U7110 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n5752) );
  OR2_X1 U7111 ( .A1(n4989), .A2(n5752), .ZN(n5642) );
  OR2_X1 U7112 ( .A1(n5640), .A2(n8923), .ZN(n5641) );
  NAND4_X1 U7113 ( .A1(n5644), .A2(n5643), .A3(n5642), .A4(n5641), .ZN(n9175)
         );
  NAND2_X1 U7114 ( .A1(n8548), .A2(n9175), .ZN(n5645) );
  OAI211_X1 U7115 ( .C1(n8550), .C2(n8946), .A(n5646), .B(n5645), .ZN(n5647)
         );
  AOI21_X1 U7116 ( .B1(n8945), .B2(n8552), .A(n5647), .ZN(n5648) );
  INV_X1 U7117 ( .A(n5648), .ZN(n5649) );
  NAND3_X1 U7118 ( .A1(n5652), .A2(n5651), .A3(n5650), .ZN(P1_U3218) );
  INV_X2 U7119 ( .A(n7103), .ZN(n8802) );
  INV_X1 U7120 ( .A(n7100), .ZN(n6680) );
  AND2_X1 U7121 ( .A1(n5653), .A2(n6680), .ZN(n7094) );
  NAND2_X1 U7122 ( .A1(n5713), .A2(n7094), .ZN(n7093) );
  NAND2_X1 U7123 ( .A1(n8849), .A2(n7103), .ZN(n5654) );
  NAND2_X1 U7124 ( .A1(n7093), .A2(n5654), .ZN(n6813) );
  INV_X1 U7125 ( .A(n6813), .ZN(n5657) );
  XNOR2_X1 U7126 ( .A(n5655), .B(n7186), .ZN(n8694) );
  NAND2_X1 U7127 ( .A1(n5657), .A2(n5656), .ZN(n6814) );
  OR2_X1 U7128 ( .A1(n5655), .A2(n7186), .ZN(n5658) );
  NAND2_X1 U7129 ( .A1(n6814), .A2(n5658), .ZN(n7504) );
  NAND2_X1 U7130 ( .A1(n8848), .A2(n9590), .ZN(n6880) );
  NAND2_X1 U7131 ( .A1(n7504), .A2(n7503), .ZN(n7506) );
  OR2_X1 U7132 ( .A1(n8848), .A2(n7510), .ZN(n5659) );
  NAND2_X1 U7133 ( .A1(n7506), .A2(n5659), .ZN(n6879) );
  OR2_X1 U7134 ( .A1(n8847), .A2(n6891), .ZN(n8687) );
  NAND2_X1 U7135 ( .A1(n8847), .A2(n6891), .ZN(n8688) );
  OR2_X1 U7136 ( .A1(n8847), .A2(n7196), .ZN(n5660) );
  OR2_X1 U7137 ( .A1(n9602), .A2(n9596), .ZN(n8691) );
  NAND2_X1 U7138 ( .A1(n9602), .A2(n8477), .ZN(n5662) );
  OR2_X1 U7139 ( .A1(n8846), .A2(n4268), .ZN(n8692) );
  NAND2_X1 U7140 ( .A1(n8846), .A2(n4268), .ZN(n8749) );
  AND2_X1 U7141 ( .A1(n8692), .A2(n8749), .ZN(n8569) );
  OR2_X1 U7142 ( .A1(n8846), .A2(n4269), .ZN(n5663) );
  NAND2_X1 U7143 ( .A1(n9601), .A2(n7209), .ZN(n8771) );
  OR2_X1 U7144 ( .A1(n9601), .A2(n7158), .ZN(n5664) );
  OR2_X1 U7145 ( .A1(n9547), .A2(n7423), .ZN(n8740) );
  NAND2_X1 U7146 ( .A1(n9547), .A2(n7423), .ZN(n9544) );
  NAND2_X1 U7147 ( .A1(n8740), .A2(n9544), .ZN(n8700) );
  AND2_X1 U7148 ( .A1(n8845), .A2(n9555), .ZN(n5665) );
  NAND2_X1 U7149 ( .A1(n9414), .A2(n9373), .ZN(n8587) );
  NAND2_X1 U7150 ( .A1(n8755), .A2(n8587), .ZN(n5723) );
  NAND2_X1 U7151 ( .A1(n7361), .A2(n5723), .ZN(n5667) );
  OR2_X1 U7152 ( .A1(n9373), .A2(n9548), .ZN(n5666) );
  NAND2_X1 U7153 ( .A1(n5667), .A2(n5666), .ZN(n9415) );
  XNOR2_X1 U7154 ( .A(n9451), .B(n8844), .ZN(n9416) );
  INV_X1 U7155 ( .A(n9416), .ZN(n5668) );
  NAND2_X1 U7156 ( .A1(n9451), .A2(n8844), .ZN(n5669) );
  NAND2_X1 U7157 ( .A1(n9444), .A2(n9413), .ZN(n8607) );
  NAND2_X1 U7158 ( .A1(n8608), .A2(n8607), .ZN(n8706) );
  NAND2_X1 U7159 ( .A1(n9444), .A2(n8843), .ZN(n5670) );
  NAND2_X1 U7160 ( .A1(n7443), .A2(n5670), .ZN(n9395) );
  OR2_X1 U7161 ( .A1(n9407), .A2(n8842), .ZN(n5671) );
  NAND2_X1 U7162 ( .A1(n9395), .A2(n5671), .ZN(n5673) );
  NAND2_X1 U7163 ( .A1(n9407), .A2(n8842), .ZN(n5672) );
  NAND2_X1 U7164 ( .A1(n5673), .A2(n5672), .ZN(n7466) );
  INV_X1 U7165 ( .A(n7466), .ZN(n5674) );
  OR2_X1 U7166 ( .A1(n8430), .A2(n9266), .ZN(n5675) );
  NAND2_X1 U7167 ( .A1(n9264), .A2(n9255), .ZN(n5676) );
  NAND2_X1 U7168 ( .A1(n5677), .A2(n5676), .ZN(n9131) );
  INV_X1 U7169 ( .A(n9265), .ZN(n5678) );
  NAND2_X1 U7170 ( .A1(n9254), .A2(n5678), .ZN(n8767) );
  NAND2_X1 U7171 ( .A1(n9116), .A2(n8767), .ZN(n9132) );
  NAND2_X1 U7172 ( .A1(n9131), .A2(n9132), .ZN(n5680) );
  NAND2_X1 U7173 ( .A1(n9254), .A2(n9265), .ZN(n5679) );
  NAND2_X1 U7174 ( .A1(n5680), .A2(n5679), .ZN(n9124) );
  OR2_X1 U7175 ( .A1(n9126), .A2(n9256), .ZN(n5681) );
  NAND2_X1 U7176 ( .A1(n9124), .A2(n5681), .ZN(n5683) );
  NAND2_X1 U7177 ( .A1(n9126), .A2(n9256), .ZN(n5682) );
  INV_X1 U7178 ( .A(n9233), .ZN(n5684) );
  OR2_X1 U7179 ( .A1(n9241), .A2(n5684), .ZN(n8621) );
  NAND2_X1 U7180 ( .A1(n9241), .A2(n5684), .ZN(n8623) );
  NAND2_X1 U7181 ( .A1(n8621), .A2(n8623), .ZN(n9098) );
  NAND2_X1 U7182 ( .A1(n9241), .A2(n9233), .ZN(n5685) );
  AND2_X1 U7183 ( .A1(n9231), .A2(n9242), .ZN(n5686) );
  NOR2_X1 U7184 ( .A1(n9228), .A2(n9232), .ZN(n5687) );
  NAND2_X1 U7185 ( .A1(n8456), .A2(n9069), .ZN(n8633) );
  NAND2_X1 U7186 ( .A1(n8729), .A2(n8633), .ZN(n9054) );
  NAND2_X1 U7187 ( .A1(n9053), .A2(n9054), .ZN(n5689) );
  NAND2_X1 U7188 ( .A1(n8456), .A2(n9038), .ZN(n5688) );
  NAND2_X1 U7189 ( .A1(n5689), .A2(n5688), .ZN(n9032) );
  OR2_X1 U7190 ( .A1(n9215), .A2(n9218), .ZN(n5690) );
  AND2_X1 U7191 ( .A1(n5731), .A2(n9201), .ZN(n5691) );
  AND2_X1 U7192 ( .A1(n9204), .A2(n9023), .ZN(n5692) );
  OAI22_X1 U7193 ( .A1(n9006), .A2(n5692), .B1(n9023), .B2(n9204), .ZN(n8986)
         );
  INV_X1 U7194 ( .A(n9013), .ZN(n9200) );
  NAND2_X1 U7195 ( .A1(n8990), .A2(n9200), .ZN(n8655) );
  NAND2_X1 U7196 ( .A1(n8737), .A2(n8655), .ZN(n8995) );
  OR2_X1 U7197 ( .A1(n8990), .A2(n9013), .ZN(n5693) );
  NOR2_X1 U7198 ( .A1(n8973), .A2(n8999), .ZN(n8659) );
  INV_X1 U7199 ( .A(n8659), .ZN(n5694) );
  NAND2_X1 U7200 ( .A1(n8973), .A2(n8999), .ZN(n5695) );
  NAND2_X1 U7201 ( .A1(n5696), .A2(n5695), .ZN(n8956) );
  NAND2_X1 U7202 ( .A1(n9186), .A2(n5697), .ZN(n8780) );
  INV_X1 U7203 ( .A(n8964), .ZN(n5698) );
  OR2_X1 U7204 ( .A1(n9186), .A2(n9176), .ZN(n5700) );
  INV_X1 U7205 ( .A(n8965), .ZN(n5747) );
  OR2_X1 U7206 ( .A1(n8945), .A2(n5747), .ZN(n8722) );
  NAND2_X1 U7207 ( .A1(n8945), .A2(n5747), .ZN(n8783) );
  INV_X1 U7208 ( .A(SI_28_), .ZN(n5703) );
  INV_X1 U7209 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n7536) );
  INV_X1 U7210 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n7530) );
  MUX2_X1 U7211 ( .A(n7536), .B(n7530), .S(n7698), .Z(n7519) );
  XNOR2_X1 U7212 ( .A(n7519), .B(SI_29_), .ZN(n5705) );
  NAND2_X1 U7213 ( .A1(n7688), .A2(n8563), .ZN(n5707) );
  OR2_X1 U7214 ( .A1(n5000), .A2(n7536), .ZN(n5706) );
  XNOR2_X1 U7215 ( .A(n8786), .B(n9175), .ZN(n8716) );
  INV_X1 U7216 ( .A(n8716), .ZN(n5708) );
  XNOR2_X1 U7217 ( .A(n5709), .B(n5708), .ZN(n8921) );
  NAND2_X1 U7218 ( .A1(n4265), .A2(n9123), .ZN(n5711) );
  MUX2_X1 U7219 ( .A(n5712), .B(n5711), .S(n5710), .Z(n9419) );
  NAND2_X1 U7220 ( .A1(n7151), .A2(n9074), .ZN(n9570) );
  INV_X1 U7221 ( .A(n9570), .ZN(n8830) );
  NAND2_X1 U7222 ( .A1(n4265), .A2(n8830), .ZN(n9582) );
  OR2_X1 U7223 ( .A1(n8680), .A2(n5637), .ZN(n9438) );
  INV_X1 U7224 ( .A(n5713), .ZN(n8696) );
  NOR2_X1 U7225 ( .A1(n5653), .A2(n7100), .ZN(n7095) );
  NAND2_X1 U7226 ( .A1(n8696), .A2(n7095), .ZN(n5715) );
  OR2_X1 U7227 ( .A1(n8849), .A2(n8802), .ZN(n5714) );
  NAND2_X1 U7228 ( .A1(n8804), .A2(n4267), .ZN(n5716) );
  INV_X1 U7229 ( .A(n7186), .ZN(n8809) );
  OR2_X1 U7230 ( .A1(n5655), .A2(n8809), .ZN(n8803) );
  NAND2_X1 U7231 ( .A1(n5716), .A2(n8803), .ZN(n8747) );
  INV_X1 U7232 ( .A(n8686), .ZN(n8811) );
  OR2_X1 U7233 ( .A1(n8747), .A2(n8811), .ZN(n6881) );
  AND2_X1 U7234 ( .A1(n8688), .A2(n6880), .ZN(n5717) );
  NAND2_X1 U7235 ( .A1(n6881), .A2(n8810), .ZN(n7028) );
  NAND2_X1 U7236 ( .A1(n8691), .A2(n8687), .ZN(n5718) );
  NAND2_X1 U7237 ( .A1(n5719), .A2(n5718), .ZN(n5720) );
  NAND2_X1 U7238 ( .A1(n7028), .A2(n8813), .ZN(n5721) );
  INV_X1 U7239 ( .A(n7027), .ZN(n8695) );
  NAND2_X1 U7240 ( .A1(n5721), .A2(n8695), .ZN(n7030) );
  NAND2_X1 U7241 ( .A1(n7030), .A2(n8739), .ZN(n7347) );
  INV_X1 U7242 ( .A(n8740), .ZN(n5722) );
  NAND2_X1 U7243 ( .A1(n9613), .A2(n8845), .ZN(n8701) );
  AND2_X1 U7244 ( .A1(n8701), .A2(n9544), .ZN(n8756) );
  OR2_X1 U7245 ( .A1(n8845), .A2(n9613), .ZN(n8702) );
  NAND2_X1 U7246 ( .A1(n8587), .A2(n8702), .ZN(n8757) );
  NAND2_X1 U7247 ( .A1(n8757), .A2(n8755), .ZN(n8741) );
  NAND2_X1 U7248 ( .A1(n9412), .A2(n9416), .ZN(n5725) );
  INV_X1 U7249 ( .A(n8844), .ZN(n9439) );
  NAND2_X1 U7250 ( .A1(n9451), .A2(n9439), .ZN(n8606) );
  OR2_X1 U7251 ( .A1(n9451), .A2(n9439), .ZN(n5726) );
  NAND2_X1 U7252 ( .A1(n8608), .A2(n5726), .ZN(n5727) );
  NAND2_X1 U7253 ( .A1(n5727), .A2(n8607), .ZN(n8594) );
  INV_X1 U7254 ( .A(n8842), .ZN(n9441) );
  OR2_X1 U7255 ( .A1(n9407), .A2(n9441), .ZN(n8611) );
  NAND2_X1 U7256 ( .A1(n9407), .A2(n9441), .ZN(n8595) );
  NAND2_X1 U7257 ( .A1(n8611), .A2(n8595), .ZN(n9397) );
  INV_X1 U7258 ( .A(n9266), .ZN(n9402) );
  OR2_X1 U7259 ( .A1(n8430), .A2(n9402), .ZN(n8612) );
  NAND2_X1 U7260 ( .A1(n8430), .A2(n9402), .ZN(n8614) );
  INV_X1 U7261 ( .A(n9255), .ZN(n5728) );
  NOR2_X1 U7262 ( .A1(n9264), .A2(n5728), .ZN(n8765) );
  NAND2_X1 U7263 ( .A1(n9264), .A2(n5728), .ZN(n8744) );
  INV_X1 U7264 ( .A(n8767), .ZN(n8746) );
  NAND2_X1 U7265 ( .A1(n9117), .A2(n9116), .ZN(n5729) );
  INV_X1 U7266 ( .A(n9256), .ZN(n9139) );
  NAND2_X1 U7267 ( .A1(n9126), .A2(n9139), .ZN(n8597) );
  INV_X1 U7268 ( .A(n9242), .ZN(n9104) );
  OR2_X1 U7269 ( .A1(n9231), .A2(n9104), .ZN(n8624) );
  NAND2_X1 U7270 ( .A1(n9231), .A2(n9104), .ZN(n8772) );
  INV_X1 U7271 ( .A(n9232), .ZN(n9087) );
  NAND2_X1 U7272 ( .A1(n9228), .A2(n9087), .ZN(n8631) );
  NAND2_X1 U7273 ( .A1(n8627), .A2(n8631), .ZN(n9066) );
  OAI21_X1 U7274 ( .B1(n9067), .B2(n9066), .A(n8627), .ZN(n9052) );
  INV_X1 U7275 ( .A(n9218), .ZN(n8437) );
  NAND2_X1 U7276 ( .A1(n9215), .A2(n8437), .ZN(n8636) );
  NAND2_X1 U7277 ( .A1(n8638), .A2(n8636), .ZN(n9034) );
  INV_X1 U7278 ( .A(n8633), .ZN(n9033) );
  NOR2_X1 U7279 ( .A1(n9034), .A2(n9033), .ZN(n5730) );
  NAND2_X1 U7280 ( .A1(n9036), .A2(n8638), .ZN(n9022) );
  OR2_X1 U7281 ( .A1(n5731), .A2(n9039), .ZN(n8642) );
  NAND2_X1 U7282 ( .A1(n5731), .A2(n9039), .ZN(n8734) );
  INV_X1 U7283 ( .A(n9023), .ZN(n8641) );
  XNOR2_X1 U7284 ( .A(n9204), .B(n8641), .ZN(n9007) );
  AND2_X1 U7285 ( .A1(n9204), .A2(n8641), .ZN(n8996) );
  NOR2_X1 U7286 ( .A1(n8995), .A2(n8996), .ZN(n5732) );
  NAND2_X1 U7287 ( .A1(n8997), .A2(n8737), .ZN(n8980) );
  INV_X1 U7288 ( .A(n8999), .ZN(n8654) );
  NAND2_X1 U7289 ( .A1(n8973), .A2(n8654), .ZN(n8779) );
  NAND2_X1 U7290 ( .A1(n8980), .A2(n8979), .ZN(n8978) );
  NAND2_X1 U7291 ( .A1(n8978), .A2(n8736), .ZN(n8963) );
  INV_X1 U7292 ( .A(n8932), .ZN(n8938) );
  INV_X1 U7293 ( .A(n8937), .ZN(n8650) );
  NOR2_X1 U7294 ( .A1(n8938), .A2(n8650), .ZN(n5733) );
  NAND2_X1 U7295 ( .A1(n8936), .A2(n5733), .ZN(n8940) );
  NAND2_X1 U7296 ( .A1(n8940), .A2(n8783), .ZN(n5734) );
  XNOR2_X1 U7297 ( .A(n5734), .B(n8716), .ZN(n5746) );
  OR2_X1 U7298 ( .A1(n4265), .A2(n9123), .ZN(n5736) );
  INV_X1 U7299 ( .A(n7151), .ZN(n8797) );
  NAND2_X1 U7300 ( .A1(n5621), .A2(n8797), .ZN(n5735) );
  INV_X1 U7301 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n5740) );
  NAND2_X1 U7302 ( .A1(n5162), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n5739) );
  INV_X1 U7303 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n5737) );
  OR2_X1 U7304 ( .A1(n4989), .A2(n5737), .ZN(n5738) );
  OAI211_X1 U7305 ( .C1(n4273), .C2(n5740), .A(n5739), .B(n5738), .ZN(n8841)
         );
  INV_X1 U7306 ( .A(P1_B_REG_SCAN_IN), .ZN(n5743) );
  NOR2_X1 U7307 ( .A1(n9337), .A2(n5743), .ZN(n5744) );
  NOR2_X1 U7308 ( .A1(n9440), .A2(n5744), .ZN(n8911) );
  NAND2_X1 U7309 ( .A1(n8802), .A2(n7100), .ZN(n7099) );
  OR2_X1 U7310 ( .A1(n7099), .A2(n7186), .ZN(n7511) );
  OR2_X1 U7311 ( .A1(n7511), .A2(n7510), .ZN(n7513) );
  NAND2_X1 U7312 ( .A1(n9560), .A2(n9613), .ZN(n9558) );
  INV_X1 U7313 ( .A(n9444), .ZN(n7450) );
  INV_X1 U7314 ( .A(n9407), .ZN(n9433) );
  INV_X1 U7315 ( .A(n9126), .ZN(n9318) );
  NAND2_X1 U7316 ( .A1(n9111), .A2(n9318), .ZN(n9112) );
  OR2_X2 U7317 ( .A1(n9112), .A2(n9241), .ZN(n9105) );
  INV_X1 U7318 ( .A(n9204), .ZN(n9015) );
  AND2_X2 U7319 ( .A1(n9026), .A2(n9015), .ZN(n9008) );
  NAND2_X1 U7320 ( .A1(n8942), .A2(n8926), .ZN(n8915) );
  OAI211_X1 U7321 ( .C1(n8942), .C2(n8926), .A(n8915), .B(n9559), .ZN(n8924)
         );
  AOI21_X1 U7322 ( .B1(n8921), .B2(n9615), .A(n5748), .ZN(n5757) );
  INV_X1 U7323 ( .A(n6314), .ZN(n5750) );
  OAI211_X1 U7324 ( .C1(n7089), .C2(n9570), .A(n5750), .B(n5749), .ZN(n5751)
         );
  MUX2_X1 U7325 ( .A(n5752), .B(n5757), .S(n9619), .Z(n5755) );
  INV_X1 U7326 ( .A(n9326), .ZN(n5753) );
  NAND2_X1 U7327 ( .A1(n8786), .A2(n5753), .ZN(n5754) );
  NAND2_X1 U7328 ( .A1(n5755), .A2(n5754), .ZN(P1_U3520) );
  MUX2_X1 U7329 ( .A(n9813), .B(n5757), .S(n4270), .Z(n5760) );
  INV_X1 U7330 ( .A(n9280), .ZN(n5758) );
  NAND2_X1 U7331 ( .A1(n8786), .A2(n5758), .ZN(n5759) );
  NAND2_X1 U7332 ( .A1(n5760), .A2(n5759), .ZN(P1_U3552) );
  NAND2_X1 U7333 ( .A1(n5822), .A2(n5761), .ZN(n5848) );
  INV_X1 U7334 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5762) );
  NAND2_X1 U7335 ( .A1(n5763), .A2(n5762), .ZN(n5764) );
  NOR2_X2 U7336 ( .A1(n5848), .A2(n5764), .ZN(n5889) );
  NOR2_X1 U7337 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n5767) );
  NOR2_X1 U7338 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n5766) );
  NOR2_X1 U7339 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .ZN(
        n5765) );
  NAND2_X1 U7340 ( .A1(n5771), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5772) );
  INV_X1 U7341 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5773) );
  NAND2_X1 U7342 ( .A1(n5774), .A2(n5773), .ZN(n5775) );
  NAND2_X1 U7343 ( .A1(n5775), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5777) );
  NAND2_X1 U7344 ( .A1(n7865), .A2(n4745), .ZN(n6503) );
  NOR2_X1 U7345 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), .ZN(
        n5780) );
  NOR2_X1 U7346 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), .ZN(
        n5779) );
  NAND4_X1 U7347 ( .A1(n5781), .A2(n5780), .A3(n5779), .A4(n6225), .ZN(n5785)
         );
  NAND4_X1 U7348 ( .A1(n5783), .A2(n5782), .A3(n6222), .A4(n6246), .ZN(n5784)
         );
  MUX2_X1 U7349 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5790), .S(
        P2_IR_REG_27__SCAN_IN), .Z(n5791) );
  AND2_X2 U7350 ( .A1(n6364), .A2(n5793), .ZN(n6050) );
  NAND2_X1 U7351 ( .A1(n6050), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n5795) );
  NAND2_X1 U7352 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n9638), .ZN(n5794) );
  NOR2_X2 U7353 ( .A1(n5797), .A2(P2_IR_REG_29__SCAN_IN), .ZN(n8406) );
  OR2_X2 U7354 ( .A1(n8406), .A2(n8407), .ZN(n5799) );
  XNOR2_X2 U7355 ( .A(n5799), .B(P2_IR_REG_30__SCAN_IN), .ZN(n5800) );
  NAND2_X1 U7356 ( .A1(n5839), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n5802) );
  NAND2_X1 U7357 ( .A1(n5837), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n5801) );
  AND3_X1 U7358 ( .A1(n5803), .A2(n5802), .A3(n5801), .ZN(n5806) );
  NAND2_X1 U7359 ( .A1(n6124), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5805) );
  NAND2_X1 U7360 ( .A1(n6124), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5813) );
  NAND2_X1 U7361 ( .A1(n6329), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5812) );
  NAND2_X1 U7362 ( .A1(n5839), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5811) );
  NAND2_X1 U7363 ( .A1(n5837), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n5810) );
  NAND2_X1 U7364 ( .A1(n7919), .A2(n6783), .ZN(n5815) );
  NAND2_X1 U7365 ( .A1(n7698), .A2(SI_0_), .ZN(n5814) );
  XNOR2_X1 U7366 ( .A(n5814), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n8420) );
  NAND2_X1 U7367 ( .A1(n6635), .A2(n6634), .ZN(n6633) );
  INV_X1 U7368 ( .A(n5818), .ZN(n5819) );
  NAND2_X1 U7369 ( .A1(n6633), .A2(n5819), .ZN(n6614) );
  INV_X1 U7370 ( .A(n6304), .ZN(n5821) );
  NAND2_X1 U7371 ( .A1(n5932), .A2(n5821), .ZN(n5826) );
  NAND2_X1 U7372 ( .A1(n6050), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n5825) );
  OR2_X1 U7373 ( .A1(n5822), .A2(n8407), .ZN(n5823) );
  XNOR2_X1 U7374 ( .A(n5823), .B(P2_IR_REG_2__SCAN_IN), .ZN(n9362) );
  NAND2_X1 U7375 ( .A1(n6322), .A2(n9362), .ZN(n5824) );
  XNOR2_X1 U7376 ( .A(n6210), .B(n6968), .ZN(n5832) );
  NAND2_X1 U7377 ( .A1(n6124), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5830) );
  NAND2_X1 U7378 ( .A1(n5837), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n5829) );
  NAND2_X1 U7379 ( .A1(n5839), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5827) );
  NAND2_X1 U7380 ( .A1(n7917), .A2(n6783), .ZN(n5831) );
  XNOR2_X1 U7381 ( .A(n5832), .B(n5831), .ZN(n6615) );
  OAI22_X1 U7382 ( .A1(n6614), .A2(n6615), .B1(n5832), .B2(n5831), .ZN(n6752)
         );
  NAND2_X1 U7383 ( .A1(n7702), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n5836) );
  OR3_X1 U7384 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .A3(
        n9638), .ZN(n5833) );
  NAND2_X1 U7385 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n5833), .ZN(n5834) );
  XNOR2_X1 U7386 ( .A(n5834), .B(P2_IR_REG_3__SCAN_IN), .ZN(n6373) );
  NAND2_X1 U7387 ( .A1(n6322), .A2(n6373), .ZN(n5835) );
  XNOR2_X1 U7388 ( .A(n6210), .B(n6695), .ZN(n5845) );
  CLKBUF_X3 U7389 ( .A(n5837), .Z(n6185) );
  NAND2_X1 U7390 ( .A1(n6185), .A2(n7923), .ZN(n5843) );
  NAND2_X1 U7391 ( .A1(n6124), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5842) );
  INV_X2 U7392 ( .A(n6266), .ZN(n7678) );
  NAND2_X1 U7393 ( .A1(n7678), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n5841) );
  NAND2_X1 U7394 ( .A1(n5839), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5840) );
  NAND2_X1 U7395 ( .A1(n7916), .A2(n6783), .ZN(n5844) );
  XNOR2_X1 U7396 ( .A(n5845), .B(n5844), .ZN(n6753) );
  INV_X1 U7397 ( .A(n5844), .ZN(n5846) );
  AOI21_X1 U7398 ( .B1(n6752), .B2(n6753), .A(n5847), .ZN(n6721) );
  NAND2_X1 U7399 ( .A1(n7702), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n5852) );
  NAND2_X1 U7400 ( .A1(n5849), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5850) );
  XNOR2_X1 U7401 ( .A(n5850), .B(P2_IR_REG_4__SCAN_IN), .ZN(n6439) );
  NAND2_X1 U7402 ( .A1(n6322), .A2(n6439), .ZN(n5851) );
  OAI211_X1 U7403 ( .C1(n5911), .C2(n6295), .A(n5852), .B(n5851), .ZN(n6919)
         );
  XNOR2_X1 U7404 ( .A(n6210), .B(n6919), .ZN(n5859) );
  NAND2_X1 U7405 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n5866) );
  OAI21_X1 U7406 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(P2_REG3_REG_4__SCAN_IN), 
        .A(n5866), .ZN(n6913) );
  INV_X1 U7407 ( .A(n6913), .ZN(n6729) );
  NAND2_X1 U7408 ( .A1(n6185), .A2(n6729), .ZN(n5857) );
  NAND2_X1 U7409 ( .A1(n6124), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5856) );
  NAND2_X1 U7410 ( .A1(n7678), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5855) );
  INV_X4 U7411 ( .A(n5853), .ZN(n6263) );
  NAND2_X1 U7412 ( .A1(n6263), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n5854) );
  NAND4_X1 U7413 ( .A1(n5857), .A2(n5856), .A3(n5855), .A4(n5854), .ZN(n7915)
         );
  AND2_X1 U7414 ( .A1(n7915), .A2(n6783), .ZN(n5858) );
  NAND2_X1 U7415 ( .A1(n5859), .A2(n5858), .ZN(n6723) );
  NOR2_X1 U7416 ( .A1(n5859), .A2(n5858), .ZN(n6722) );
  INV_X1 U7417 ( .A(n6298), .ZN(n5860) );
  NAND2_X1 U7418 ( .A1(n5860), .A2(n7701), .ZN(n5864) );
  NAND2_X1 U7419 ( .A1(n7702), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n5863) );
  OR2_X1 U7420 ( .A1(n5849), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n5861) );
  NAND2_X1 U7421 ( .A1(n5861), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5881) );
  XNOR2_X1 U7422 ( .A(n5881), .B(P2_IR_REG_5__SCAN_IN), .ZN(n6444) );
  NAND2_X1 U7423 ( .A1(n6322), .A2(n6444), .ZN(n5862) );
  XNOR2_X1 U7424 ( .A(n6210), .B(n6979), .ZN(n5873) );
  NAND2_X1 U7425 ( .A1(n6263), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5871) );
  NAND2_X1 U7426 ( .A1(n7677), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n5870) );
  INV_X1 U7427 ( .A(n5866), .ZN(n5865) );
  NAND2_X1 U7428 ( .A1(n5865), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5901) );
  INV_X1 U7429 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n7937) );
  NAND2_X1 U7430 ( .A1(n5866), .A2(n7937), .ZN(n5867) );
  AND2_X1 U7431 ( .A1(n5901), .A2(n5867), .ZN(n6904) );
  NAND2_X1 U7432 ( .A1(n6185), .A2(n6904), .ZN(n5869) );
  NAND2_X1 U7433 ( .A1(n6329), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n5868) );
  NAND4_X1 U7434 ( .A1(n5871), .A2(n5870), .A3(n5869), .A4(n5868), .ZN(n7914)
         );
  NAND2_X1 U7435 ( .A1(n7914), .A2(n6783), .ZN(n5872) );
  NOR2_X1 U7436 ( .A1(n5873), .A2(n5872), .ZN(n5874) );
  AOI21_X1 U7437 ( .B1(n5873), .B2(n5872), .A(n5874), .ZN(n6709) );
  INV_X1 U7438 ( .A(n5874), .ZN(n5875) );
  NAND2_X1 U7439 ( .A1(n6263), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5879) );
  NAND2_X1 U7440 ( .A1(n6124), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5878) );
  XNOR2_X1 U7441 ( .A(n5901), .B(P2_REG3_REG_6__SCAN_IN), .ZN(n6975) );
  NAND2_X1 U7442 ( .A1(n6185), .A2(n6975), .ZN(n5877) );
  NAND2_X1 U7443 ( .A1(n6329), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n5876) );
  NAND4_X1 U7444 ( .A1(n5879), .A2(n5878), .A3(n5877), .A4(n5876), .ZN(n7913)
         );
  NAND2_X1 U7445 ( .A1(n7913), .A2(n6783), .ZN(n5887) );
  NAND2_X1 U7446 ( .A1(n5881), .A2(n5880), .ZN(n5882) );
  NAND2_X1 U7447 ( .A1(n5882), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5883) );
  XNOR2_X1 U7448 ( .A(n5883), .B(P2_IR_REG_6__SCAN_IN), .ZN(n6445) );
  AOI22_X1 U7449 ( .A1(n7702), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n6322), .B2(
        n6445), .ZN(n5885) );
  OR2_X1 U7450 ( .A1(n5911), .A2(n6307), .ZN(n5884) );
  NAND2_X1 U7451 ( .A1(n5885), .A2(n5884), .ZN(n6716) );
  XNOR2_X1 U7452 ( .A(n6210), .B(n6716), .ZN(n5886) );
  XOR2_X1 U7453 ( .A(n5887), .B(n5886), .Z(n6714) );
  INV_X1 U7454 ( .A(n5886), .ZN(n5888) );
  OR2_X1 U7455 ( .A1(n6312), .A2(n5911), .ZN(n5896) );
  INV_X1 U7456 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n8407) );
  NOR2_X1 U7457 ( .A1(n5890), .A2(n8407), .ZN(n5891) );
  MUX2_X1 U7458 ( .A(n8407), .B(n5891), .S(P2_IR_REG_7__SCAN_IN), .Z(n5894) );
  NAND2_X1 U7459 ( .A1(n5890), .A2(n5892), .ZN(n5913) );
  INV_X1 U7460 ( .A(n5913), .ZN(n5893) );
  INV_X1 U7461 ( .A(n6522), .ZN(n6530) );
  AOI22_X1 U7462 ( .A1(n7702), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n6322), .B2(
        n6530), .ZN(n5895) );
  NAND2_X1 U7463 ( .A1(n5896), .A2(n5895), .ZN(n7050) );
  XNOR2_X1 U7464 ( .A(n7050), .B(n4502), .ZN(n5908) );
  NAND2_X1 U7465 ( .A1(n6263), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5906) );
  NAND2_X1 U7466 ( .A1(n7677), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n5905) );
  INV_X1 U7467 ( .A(n5901), .ZN(n5898) );
  NAND2_X1 U7468 ( .A1(n5898), .A2(n5897), .ZN(n5918) );
  INV_X1 U7469 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n5900) );
  INV_X1 U7470 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n5899) );
  OAI21_X1 U7471 ( .B1(n5901), .B2(n5900), .A(n5899), .ZN(n5902) );
  AND2_X1 U7472 ( .A1(n5918), .A2(n5902), .ZN(n7012) );
  NAND2_X1 U7473 ( .A1(n6185), .A2(n7012), .ZN(n5904) );
  NAND2_X1 U7474 ( .A1(n7678), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n5903) );
  NAND4_X1 U7475 ( .A1(n5906), .A2(n5905), .A3(n5904), .A4(n5903), .ZN(n9655)
         );
  NAND2_X1 U7476 ( .A1(n9655), .A2(n6783), .ZN(n5907) );
  NOR2_X1 U7477 ( .A1(n5908), .A2(n5907), .ZN(n5909) );
  AOI21_X1 U7478 ( .B1(n5908), .B2(n5907), .A(n5909), .ZN(n6829) );
  INV_X1 U7479 ( .A(n5909), .ZN(n5910) );
  NAND2_X1 U7480 ( .A1(n6828), .A2(n5910), .ZN(n6873) );
  OR2_X1 U7481 ( .A1(n6317), .A2(n5911), .ZN(n5916) );
  NAND2_X1 U7482 ( .A1(n5913), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5912) );
  MUX2_X1 U7483 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5912), .S(
        P2_IR_REG_8__SCAN_IN), .Z(n5914) );
  AOI22_X1 U7484 ( .A1(n7702), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n6322), .B2(
        n7953), .ZN(n5915) );
  NAND2_X1 U7485 ( .A1(n5916), .A2(n5915), .ZN(n7056) );
  XNOR2_X1 U7486 ( .A(n7056), .B(n4502), .ZN(n5925) );
  NAND2_X1 U7487 ( .A1(n6263), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n5923) );
  NAND2_X1 U7488 ( .A1(n7677), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5922) );
  INV_X1 U7489 ( .A(n5918), .ZN(n5917) );
  NAND2_X1 U7490 ( .A1(n5917), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5946) );
  INV_X1 U7491 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n9809) );
  NAND2_X1 U7492 ( .A1(n5918), .A2(n9809), .ZN(n5919) );
  AND2_X1 U7493 ( .A1(n5946), .A2(n5919), .ZN(n9664) );
  NAND2_X1 U7494 ( .A1(n6185), .A2(n9664), .ZN(n5921) );
  NAND2_X1 U7495 ( .A1(n7678), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n5920) );
  NAND4_X1 U7496 ( .A1(n5923), .A2(n5922), .A3(n5921), .A4(n5920), .ZN(n7912)
         );
  NAND2_X1 U7497 ( .A1(n7912), .A2(n6783), .ZN(n5924) );
  NOR2_X1 U7498 ( .A1(n5925), .A2(n5924), .ZN(n5926) );
  AOI21_X1 U7499 ( .B1(n5925), .B2(n5924), .A(n5926), .ZN(n6872) );
  INV_X1 U7500 ( .A(n5926), .ZN(n5927) );
  NAND2_X1 U7501 ( .A1(n6263), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5931) );
  NAND2_X1 U7502 ( .A1(n7677), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n5930) );
  XNOR2_X1 U7503 ( .A(n5946), .B(P2_REG3_REG_9__SCAN_IN), .ZN(n7058) );
  NAND2_X1 U7504 ( .A1(n6185), .A2(n7058), .ZN(n5929) );
  NAND2_X1 U7505 ( .A1(n6329), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n5928) );
  NAND4_X1 U7506 ( .A1(n5931), .A2(n5930), .A3(n5929), .A4(n5928), .ZN(n9654)
         );
  NAND2_X1 U7507 ( .A1(n9654), .A2(n6783), .ZN(n5936) );
  NAND2_X1 U7508 ( .A1(n6319), .A2(n7701), .ZN(n5935) );
  NAND2_X1 U7509 ( .A1(n5939), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5933) );
  XNOR2_X1 U7510 ( .A(n5933), .B(P2_IR_REG_9__SCAN_IN), .ZN(n6535) );
  AOI22_X1 U7511 ( .A1(n7702), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6322), .B2(
        n6535), .ZN(n5934) );
  NAND2_X1 U7512 ( .A1(n5935), .A2(n5934), .ZN(n7071) );
  XNOR2_X1 U7513 ( .A(n7071), .B(n6210), .ZN(n5938) );
  XOR2_X1 U7514 ( .A(n5936), .B(n5938), .Z(n6953) );
  INV_X1 U7515 ( .A(n5936), .ZN(n5937) );
  NAND2_X1 U7516 ( .A1(n6335), .A2(n7701), .ZN(n5942) );
  NAND2_X1 U7517 ( .A1(n5956), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5940) );
  XNOR2_X1 U7518 ( .A(n5940), .B(P2_IR_REG_10__SCAN_IN), .ZN(n6536) );
  AOI22_X1 U7519 ( .A1(n7702), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6322), .B2(
        n6536), .ZN(n5941) );
  NAND2_X1 U7520 ( .A1(n5942), .A2(n5941), .ZN(n7164) );
  XNOR2_X1 U7521 ( .A(n7164), .B(n4502), .ZN(n5953) );
  NAND2_X1 U7522 ( .A1(n6263), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5951) );
  NAND2_X1 U7523 ( .A1(n7677), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n5950) );
  INV_X1 U7524 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5944) );
  INV_X1 U7525 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n5943) );
  OAI21_X1 U7526 ( .B1(n5946), .B2(n5944), .A(n5943), .ZN(n5947) );
  NAND2_X1 U7527 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_REG3_REG_9__SCAN_IN), 
        .ZN(n5945) );
  AND2_X1 U7528 ( .A1(n5947), .A2(n5961), .ZN(n7082) );
  NAND2_X1 U7529 ( .A1(n6185), .A2(n7082), .ZN(n5949) );
  NAND2_X1 U7530 ( .A1(n7678), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n5948) );
  NAND4_X1 U7531 ( .A1(n5951), .A2(n5950), .A3(n5949), .A4(n5948), .ZN(n7911)
         );
  NAND2_X1 U7532 ( .A1(n7911), .A2(n6783), .ZN(n5952) );
  NOR2_X1 U7533 ( .A1(n5953), .A2(n5952), .ZN(n5954) );
  AOI21_X1 U7534 ( .B1(n5953), .B2(n5952), .A(n5954), .ZN(n7064) );
  INV_X1 U7535 ( .A(n5954), .ZN(n5955) );
  NAND2_X1 U7536 ( .A1(n6338), .A2(n7701), .ZN(n5959) );
  NOR2_X1 U7537 ( .A1(n5956), .A2(P2_IR_REG_10__SCAN_IN), .ZN(n5971) );
  OR2_X1 U7538 ( .A1(n5971), .A2(n8407), .ZN(n5957) );
  XNOR2_X1 U7539 ( .A(n5957), .B(P2_IR_REG_11__SCAN_IN), .ZN(n6660) );
  AOI22_X1 U7540 ( .A1(n7702), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n6322), .B2(
        n6660), .ZN(n5958) );
  XNOR2_X1 U7541 ( .A(n7636), .B(n6210), .ZN(n5967) );
  NAND2_X1 U7542 ( .A1(n6263), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5966) );
  NAND2_X1 U7543 ( .A1(n7677), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n5965) );
  INV_X1 U7544 ( .A(n5961), .ZN(n5960) );
  NAND2_X1 U7545 ( .A1(n5960), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5976) );
  INV_X1 U7546 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n6542) );
  NAND2_X1 U7547 ( .A1(n5961), .A2(n6542), .ZN(n5962) );
  AND2_X1 U7548 ( .A1(n5976), .A2(n5962), .ZN(n7635) );
  NAND2_X1 U7549 ( .A1(n6185), .A2(n7635), .ZN(n5964) );
  NAND2_X1 U7550 ( .A1(n6329), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n5963) );
  NAND4_X1 U7551 ( .A1(n5966), .A2(n5965), .A3(n5964), .A4(n5963), .ZN(n7910)
         );
  NAND2_X1 U7552 ( .A1(n7910), .A2(n6783), .ZN(n5968) );
  XNOR2_X1 U7553 ( .A(n5967), .B(n5968), .ZN(n7633) );
  INV_X1 U7554 ( .A(n5968), .ZN(n5969) );
  NAND2_X1 U7555 ( .A1(n6549), .A2(n7701), .ZN(n5974) );
  INV_X1 U7556 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n5970) );
  NAND2_X1 U7557 ( .A1(n5971), .A2(n5970), .ZN(n5972) );
  NAND2_X1 U7558 ( .A1(n5972), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5988) );
  XNOR2_X1 U7559 ( .A(n5988), .B(P2_IR_REG_12__SCAN_IN), .ZN(n6738) );
  AOI22_X1 U7560 ( .A1(n7702), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6322), .B2(
        n6738), .ZN(n5973) );
  NAND2_X1 U7561 ( .A1(n5974), .A2(n5973), .ZN(n7387) );
  XNOR2_X1 U7562 ( .A(n7387), .B(n4502), .ZN(n5982) );
  NAND2_X1 U7563 ( .A1(n6263), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5981) );
  NAND2_X1 U7564 ( .A1(n7677), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n5980) );
  NAND2_X1 U7565 ( .A1(n5976), .A2(n5975), .ZN(n5977) );
  AND2_X1 U7566 ( .A1(n5995), .A2(n5977), .ZN(n7320) );
  NAND2_X1 U7567 ( .A1(n6185), .A2(n7320), .ZN(n5979) );
  NAND2_X1 U7568 ( .A1(n6329), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n5978) );
  NAND4_X1 U7569 ( .A1(n5981), .A2(n5980), .A3(n5979), .A4(n5978), .ZN(n7909)
         );
  NAND2_X1 U7570 ( .A1(n7909), .A2(n6783), .ZN(n5983) );
  NAND2_X1 U7571 ( .A1(n5982), .A2(n5983), .ZN(n7302) );
  NAND2_X1 U7572 ( .A1(n7303), .A2(n7302), .ZN(n5986) );
  INV_X1 U7573 ( .A(n5982), .ZN(n5985) );
  INV_X1 U7574 ( .A(n5983), .ZN(n5984) );
  NAND2_X1 U7575 ( .A1(n5985), .A2(n5984), .ZN(n7301) );
  NAND2_X1 U7576 ( .A1(n5986), .A2(n7301), .ZN(n7338) );
  NAND2_X1 U7577 ( .A1(n6612), .A2(n7701), .ZN(n5992) );
  INV_X1 U7578 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5987) );
  NAND2_X1 U7579 ( .A1(n5988), .A2(n5987), .ZN(n5989) );
  NAND2_X1 U7580 ( .A1(n5989), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5990) );
  XNOR2_X1 U7581 ( .A(n5990), .B(P2_IR_REG_13__SCAN_IN), .ZN(n6845) );
  AOI22_X1 U7582 ( .A1(n6050), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6322), .B2(
        n6845), .ZN(n5991) );
  XNOR2_X1 U7583 ( .A(n8378), .B(n6210), .ZN(n6003) );
  NAND2_X1 U7584 ( .A1(n7677), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n6000) );
  NAND2_X1 U7585 ( .A1(n7678), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n5999) );
  INV_X1 U7586 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n5994) );
  NAND2_X1 U7587 ( .A1(n5995), .A2(n5994), .ZN(n5996) );
  AND2_X1 U7588 ( .A1(n6026), .A2(n5996), .ZN(n7394) );
  NAND2_X1 U7589 ( .A1(n6185), .A2(n7394), .ZN(n5998) );
  NAND2_X1 U7590 ( .A1(n6263), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5997) );
  NAND4_X1 U7591 ( .A1(n6000), .A2(n5999), .A3(n5998), .A4(n5997), .ZN(n7908)
         );
  NAND2_X1 U7592 ( .A1(n7908), .A2(n6783), .ZN(n6001) );
  XNOR2_X1 U7593 ( .A(n6003), .B(n6001), .ZN(n7339) );
  INV_X1 U7594 ( .A(n6001), .ZN(n6002) );
  NAND2_X1 U7595 ( .A1(n6003), .A2(n6002), .ZN(n6004) );
  NAND2_X1 U7596 ( .A1(n6623), .A2(n7701), .ZN(n6008) );
  OR2_X1 U7597 ( .A1(n6005), .A2(n8407), .ZN(n6006) );
  XNOR2_X1 U7598 ( .A(n6006), .B(P2_IR_REG_14__SCAN_IN), .ZN(n6989) );
  AOI22_X1 U7599 ( .A1(n6050), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n6322), .B2(
        n6989), .ZN(n6007) );
  XNOR2_X1 U7600 ( .A(n7780), .B(n4502), .ZN(n6014) );
  XNOR2_X1 U7601 ( .A(n6026), .B(P2_REG3_REG_14__SCAN_IN), .ZN(n7548) );
  NAND2_X1 U7602 ( .A1(n6185), .A2(n7548), .ZN(n6012) );
  NAND2_X1 U7603 ( .A1(n7677), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n6011) );
  NAND2_X1 U7604 ( .A1(n7678), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n6010) );
  NAND2_X1 U7605 ( .A1(n6263), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n6009) );
  NAND4_X1 U7606 ( .A1(n6012), .A2(n6011), .A3(n6010), .A4(n6009), .ZN(n7907)
         );
  NAND2_X1 U7607 ( .A1(n7907), .A2(n6783), .ZN(n6013) );
  NAND2_X1 U7608 ( .A1(n6014), .A2(n6013), .ZN(n6015) );
  OAI21_X1 U7609 ( .B1(n6014), .B2(n6013), .A(n6015), .ZN(n7547) );
  NAND2_X1 U7610 ( .A1(n7544), .A2(n6015), .ZN(n6023) );
  INV_X1 U7611 ( .A(n6023), .ZN(n6021) );
  NAND2_X1 U7612 ( .A1(n6774), .A2(n7701), .ZN(n6019) );
  NAND2_X1 U7613 ( .A1(n6016), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6017) );
  XNOR2_X1 U7614 ( .A(n6017), .B(P2_IR_REG_15__SCAN_IN), .ZN(n7108) );
  AOI22_X1 U7615 ( .A1(n6050), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n6322), .B2(
        n7108), .ZN(n6018) );
  XOR2_X1 U7616 ( .A(n6210), .B(n8287), .Z(n6022) );
  INV_X1 U7617 ( .A(n6022), .ZN(n6020) );
  NAND2_X1 U7618 ( .A1(n6263), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n6031) );
  NAND2_X1 U7619 ( .A1(n7677), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n6030) );
  INV_X1 U7620 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n6025) );
  OAI21_X1 U7621 ( .B1(n6026), .B2(n6025), .A(n6024), .ZN(n6027) );
  AND2_X1 U7622 ( .A1(n6027), .A2(n6039), .ZN(n8291) );
  NAND2_X1 U7623 ( .A1(n6185), .A2(n8291), .ZN(n6029) );
  NAND2_X1 U7624 ( .A1(n6329), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n6028) );
  NOR2_X1 U7625 ( .A1(n7683), .A2(n6032), .ZN(n7663) );
  INV_X1 U7626 ( .A(n7663), .ZN(n6033) );
  NAND2_X1 U7627 ( .A1(n6809), .A2(n7701), .ZN(n6037) );
  NAND2_X1 U7628 ( .A1(n6035), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6052) );
  XNOR2_X1 U7629 ( .A(n6052), .B(P2_IR_REG_16__SCAN_IN), .ZN(n7996) );
  AOI22_X1 U7630 ( .A1(n6050), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n6322), .B2(
        n7996), .ZN(n6036) );
  XNOR2_X1 U7631 ( .A(n8372), .B(n6210), .ZN(n6048) );
  NAND2_X1 U7632 ( .A1(n6263), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n6044) );
  NAND2_X1 U7633 ( .A1(n7677), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n6043) );
  INV_X1 U7634 ( .A(n6039), .ZN(n6038) );
  NAND2_X1 U7635 ( .A1(n6038), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n6059) );
  INV_X1 U7636 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n9865) );
  NAND2_X1 U7637 ( .A1(n6039), .A2(n9865), .ZN(n6040) );
  AND2_X1 U7638 ( .A1(n6059), .A2(n6040), .ZN(n8273) );
  NAND2_X1 U7639 ( .A1(n6185), .A2(n8273), .ZN(n6042) );
  NAND2_X1 U7640 ( .A1(n7678), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n6041) );
  NAND4_X1 U7641 ( .A1(n6044), .A2(n6043), .A3(n6042), .A4(n6041), .ZN(n8050)
         );
  NAND2_X1 U7642 ( .A1(n8050), .A2(n6783), .ZN(n6046) );
  XNOR2_X1 U7643 ( .A(n6048), .B(n6046), .ZN(n7594) );
  INV_X1 U7644 ( .A(n6046), .ZN(n6047) );
  NAND2_X1 U7645 ( .A1(n6826), .A2(n7701), .ZN(n6056) );
  NAND2_X1 U7646 ( .A1(n6052), .A2(n6051), .ZN(n6053) );
  NAND2_X1 U7647 ( .A1(n6053), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6054) );
  XNOR2_X1 U7648 ( .A(n6054), .B(P2_IR_REG_17__SCAN_IN), .ZN(n8013) );
  AOI22_X1 U7649 ( .A1(n7702), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n6322), .B2(
        n8013), .ZN(n6055) );
  XNOR2_X1 U7650 ( .A(n8368), .B(n4502), .ZN(n6065) );
  NAND2_X1 U7651 ( .A1(n6263), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n6064) );
  NAND2_X1 U7652 ( .A1(n7677), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n6063) );
  INV_X1 U7653 ( .A(n6059), .ZN(n6057) );
  NAND2_X1 U7654 ( .A1(n6057), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n6075) );
  INV_X1 U7655 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n6058) );
  NAND2_X1 U7656 ( .A1(n6059), .A2(n6058), .ZN(n6060) );
  AND2_X1 U7657 ( .A1(n6075), .A2(n6060), .ZN(n8258) );
  NAND2_X1 U7658 ( .A1(n6185), .A2(n8258), .ZN(n6062) );
  NAND2_X1 U7659 ( .A1(n6329), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n6061) );
  NAND4_X1 U7660 ( .A1(n6064), .A2(n6063), .A3(n6062), .A4(n6061), .ZN(n8267)
         );
  NAND2_X1 U7661 ( .A1(n8267), .A2(n6783), .ZN(n6066) );
  XNOR2_X1 U7662 ( .A(n6065), .B(n6066), .ZN(n7601) );
  INV_X1 U7663 ( .A(n6065), .ZN(n6068) );
  INV_X1 U7664 ( .A(n6066), .ZN(n6067) );
  NAND2_X1 U7665 ( .A1(n6068), .A2(n6067), .ZN(n6069) );
  NAND2_X1 U7666 ( .A1(n6948), .A2(n7701), .ZN(n6073) );
  NAND2_X1 U7667 ( .A1(n6070), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6071) );
  XNOR2_X1 U7668 ( .A(n6071), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8024) );
  AOI22_X1 U7669 ( .A1(n6050), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6322), .B2(
        n8024), .ZN(n6072) );
  XNOR2_X1 U7670 ( .A(n8361), .B(n6210), .ZN(n6082) );
  NAND2_X1 U7671 ( .A1(n7677), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n6080) );
  NAND2_X1 U7672 ( .A1(n6263), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n6079) );
  INV_X1 U7673 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n6074) );
  NAND2_X1 U7674 ( .A1(n6075), .A2(n6074), .ZN(n6076) );
  AND2_X1 U7675 ( .A1(n6086), .A2(n6076), .ZN(n8234) );
  NAND2_X1 U7676 ( .A1(n6185), .A2(n8234), .ZN(n6078) );
  NAND2_X1 U7677 ( .A1(n6329), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n6077) );
  NAND4_X1 U7678 ( .A1(n6080), .A2(n6079), .A3(n6078), .A4(n6077), .ZN(n8051)
         );
  NAND2_X1 U7679 ( .A1(n8051), .A2(n6783), .ZN(n6081) );
  XNOR2_X1 U7680 ( .A(n6082), .B(n6081), .ZN(n7641) );
  INV_X1 U7681 ( .A(n6081), .ZN(n6083) );
  NAND2_X1 U7682 ( .A1(n6263), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n6091) );
  INV_X1 U7683 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n6085) );
  NAND2_X1 U7684 ( .A1(n6086), .A2(n6085), .ZN(n6087) );
  AND2_X1 U7685 ( .A1(n6098), .A2(n6087), .ZN(n8225) );
  NAND2_X1 U7686 ( .A1(n8225), .A2(n6185), .ZN(n6090) );
  NAND2_X1 U7687 ( .A1(n7677), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n6089) );
  NAND2_X1 U7688 ( .A1(n7678), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n6088) );
  NAND4_X1 U7689 ( .A1(n6091), .A2(n6090), .A3(n6089), .A4(n6088), .ZN(n8210)
         );
  AND2_X1 U7690 ( .A1(n8210), .A2(n6783), .ZN(n6095) );
  NAND2_X1 U7691 ( .A1(n7021), .A2(n7701), .ZN(n6093) );
  XNOR2_X1 U7692 ( .A(n8358), .B(n6210), .ZN(n6094) );
  NOR2_X1 U7693 ( .A1(n6094), .A2(n6095), .ZN(n6096) );
  AOI21_X1 U7694 ( .B1(n6095), .B2(n6094), .A(n6096), .ZN(n7565) );
  NAND2_X1 U7695 ( .A1(n7566), .A2(n7565), .ZN(n7564) );
  INV_X1 U7696 ( .A(n6096), .ZN(n6097) );
  INV_X1 U7697 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n7617) );
  NAND2_X1 U7698 ( .A1(n6098), .A2(n7617), .ZN(n6099) );
  NAND2_X1 U7699 ( .A1(n6112), .A2(n6099), .ZN(n8203) );
  NAND2_X1 U7700 ( .A1(n6263), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n6101) );
  NAND2_X1 U7701 ( .A1(n7677), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n6100) );
  AND2_X1 U7702 ( .A1(n6101), .A2(n6100), .ZN(n6103) );
  NAND2_X1 U7703 ( .A1(n7678), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n6102) );
  OAI211_X1 U7704 ( .C1(n8203), .C2(n6262), .A(n6103), .B(n6102), .ZN(n8196)
         );
  NAND2_X1 U7705 ( .A1(n8196), .A2(n6783), .ZN(n6107) );
  NAND2_X1 U7706 ( .A1(n7150), .A2(n7701), .ZN(n6105) );
  NAND2_X1 U7707 ( .A1(n6050), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n6104) );
  XNOR2_X1 U7708 ( .A(n8351), .B(n6210), .ZN(n6106) );
  XOR2_X1 U7709 ( .A(n6107), .B(n6106), .Z(n7615) );
  INV_X1 U7710 ( .A(n6106), .ZN(n6108) );
  NAND2_X1 U7711 ( .A1(n7248), .A2(n7701), .ZN(n6110) );
  NAND2_X1 U7712 ( .A1(n6050), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n6109) );
  XNOR2_X1 U7713 ( .A(n8346), .B(n6210), .ZN(n6117) );
  INV_X1 U7714 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n6116) );
  INV_X1 U7715 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n7574) );
  NAND2_X1 U7716 ( .A1(n6112), .A2(n7574), .ZN(n6113) );
  NAND2_X1 U7717 ( .A1(n6122), .A2(n6113), .ZN(n8188) );
  OR2_X1 U7718 ( .A1(n8188), .A2(n6262), .ZN(n6115) );
  AOI22_X1 U7719 ( .A1(n7678), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n6124), .B2(
        P2_REG1_REG_21__SCAN_IN), .ZN(n6114) );
  OAI211_X1 U7720 ( .C1(n5853), .C2(n6116), .A(n6115), .B(n6114), .ZN(n8211)
         );
  NAND2_X1 U7721 ( .A1(n8211), .A2(n6783), .ZN(n6118) );
  XNOR2_X1 U7722 ( .A(n6117), .B(n6118), .ZN(n7572) );
  INV_X1 U7723 ( .A(n6117), .ZN(n6119) );
  NAND2_X1 U7724 ( .A1(n7310), .A2(n7701), .ZN(n6121) );
  NAND2_X1 U7725 ( .A1(n6050), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n6120) );
  XNOR2_X1 U7726 ( .A(n8341), .B(n6210), .ZN(n6128) );
  INV_X1 U7727 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n6127) );
  INV_X1 U7728 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n7626) );
  NAND2_X1 U7729 ( .A1(n6122), .A2(n7626), .ZN(n6123) );
  NAND2_X1 U7730 ( .A1(n6134), .A2(n6123), .ZN(n8172) );
  OR2_X1 U7731 ( .A1(n8172), .A2(n6262), .ZN(n6126) );
  AOI22_X1 U7732 ( .A1(n6263), .A2(P2_REG0_REG_22__SCAN_IN), .B1(n6124), .B2(
        P2_REG1_REG_22__SCAN_IN), .ZN(n6125) );
  OAI211_X1 U7733 ( .C1(n6266), .C2(n6127), .A(n6126), .B(n6125), .ZN(n8195)
         );
  NAND2_X1 U7734 ( .A1(n8195), .A2(n6783), .ZN(n7623) );
  INV_X1 U7735 ( .A(n6128), .ZN(n6129) );
  NAND2_X1 U7736 ( .A1(n6130), .A2(n6129), .ZN(n6131) );
  NAND2_X1 U7737 ( .A1(n7373), .A2(n7701), .ZN(n6133) );
  NAND2_X1 U7738 ( .A1(n7702), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n6132) );
  XOR2_X1 U7739 ( .A(n6210), .B(n8334), .Z(n6141) );
  INV_X1 U7740 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n7558) );
  NAND2_X1 U7741 ( .A1(n6134), .A2(n7558), .ZN(n6135) );
  AND2_X1 U7742 ( .A1(n6145), .A2(n6135), .ZN(n8158) );
  NAND2_X1 U7743 ( .A1(n8158), .A2(n6185), .ZN(n6140) );
  INV_X1 U7744 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n9847) );
  NAND2_X1 U7745 ( .A1(n6329), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n6137) );
  NAND2_X1 U7746 ( .A1(n7677), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n6136) );
  OAI211_X1 U7747 ( .C1(n5853), .C2(n9847), .A(n6137), .B(n6136), .ZN(n6138)
         );
  INV_X1 U7748 ( .A(n6138), .ZN(n6139) );
  NAND2_X1 U7749 ( .A1(n6140), .A2(n6139), .ZN(n8139) );
  NAND2_X1 U7750 ( .A1(n8139), .A2(n6783), .ZN(n7556) );
  NAND2_X1 U7751 ( .A1(n7400), .A2(n7701), .ZN(n6143) );
  NAND2_X1 U7752 ( .A1(n7702), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n6142) );
  XNOR2_X1 U7753 ( .A(n8329), .B(n6210), .ZN(n6153) );
  INV_X1 U7754 ( .A(n6145), .ZN(n6144) );
  NAND2_X1 U7755 ( .A1(n6144), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n6161) );
  INV_X1 U7756 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n7610) );
  NAND2_X1 U7757 ( .A1(n6145), .A2(n7610), .ZN(n6146) );
  NAND2_X1 U7758 ( .A1(n6161), .A2(n6146), .ZN(n8143) );
  OR2_X1 U7759 ( .A1(n8143), .A2(n6262), .ZN(n6151) );
  INV_X1 U7760 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n8145) );
  NAND2_X1 U7761 ( .A1(n7677), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n6148) );
  NAND2_X1 U7762 ( .A1(n6263), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n6147) );
  OAI211_X1 U7763 ( .C1(n8145), .C2(n6266), .A(n6148), .B(n6147), .ZN(n6149)
         );
  INV_X1 U7764 ( .A(n6149), .ZN(n6150) );
  NAND2_X1 U7765 ( .A1(n6151), .A2(n6150), .ZN(n8154) );
  AND2_X1 U7766 ( .A1(n8154), .A2(n6783), .ZN(n7609) );
  NAND2_X1 U7767 ( .A1(n7608), .A2(n7609), .ZN(n6156) );
  INV_X1 U7768 ( .A(n6152), .ZN(n6154) );
  NAND2_X1 U7769 ( .A1(n6154), .A2(n6153), .ZN(n6155) );
  NAND2_X1 U7770 ( .A1(n7477), .A2(n7701), .ZN(n6158) );
  NAND2_X1 U7771 ( .A1(n7702), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n6157) );
  XNOR2_X1 U7772 ( .A(n8325), .B(n6210), .ZN(n7580) );
  INV_X1 U7773 ( .A(n6161), .ZN(n6159) );
  NAND2_X1 U7774 ( .A1(n6159), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n6171) );
  INV_X1 U7775 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n6160) );
  NAND2_X1 U7776 ( .A1(n6161), .A2(n6160), .ZN(n6162) );
  NAND2_X1 U7777 ( .A1(n6171), .A2(n6162), .ZN(n8124) );
  OR2_X1 U7778 ( .A1(n8124), .A2(n6262), .ZN(n6168) );
  INV_X1 U7779 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n6165) );
  NAND2_X1 U7780 ( .A1(n6263), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n6164) );
  NAND2_X1 U7781 ( .A1(n7677), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n6163) );
  OAI211_X1 U7782 ( .C1(n6165), .C2(n6266), .A(n6164), .B(n6163), .ZN(n6166)
         );
  INV_X1 U7783 ( .A(n6166), .ZN(n6167) );
  NAND2_X1 U7784 ( .A1(n6168), .A2(n6167), .ZN(n8140) );
  NAND2_X1 U7785 ( .A1(n8140), .A2(n6783), .ZN(n7579) );
  NAND2_X1 U7786 ( .A1(n8416), .A2(n7701), .ZN(n6170) );
  NAND2_X1 U7787 ( .A1(n7702), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n6169) );
  XNOR2_X1 U7788 ( .A(n8321), .B(n6210), .ZN(n6180) );
  INV_X1 U7789 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n7654) );
  NAND2_X1 U7790 ( .A1(n6171), .A2(n7654), .ZN(n6172) );
  NAND2_X1 U7791 ( .A1(n8115), .A2(n6185), .ZN(n6178) );
  INV_X1 U7792 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n6175) );
  NAND2_X1 U7793 ( .A1(n6263), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n6174) );
  NAND2_X1 U7794 ( .A1(n7677), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n6173) );
  OAI211_X1 U7795 ( .C1(n6175), .C2(n6266), .A(n6174), .B(n6173), .ZN(n6176)
         );
  INV_X1 U7796 ( .A(n6176), .ZN(n6177) );
  NAND2_X1 U7797 ( .A1(n6178), .A2(n6177), .ZN(n8101) );
  AND2_X1 U7798 ( .A1(n8101), .A2(n6783), .ZN(n6179) );
  NAND2_X1 U7799 ( .A1(n6180), .A2(n6179), .ZN(n6182) );
  OAI21_X1 U7800 ( .B1(n6180), .B2(n6179), .A(n6182), .ZN(n7649) );
  INV_X1 U7801 ( .A(n7649), .ZN(n6181) );
  NAND2_X1 U7802 ( .A1(n8412), .A2(n7701), .ZN(n6184) );
  NAND2_X1 U7803 ( .A1(n7702), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n6183) );
  XNOR2_X1 U7804 ( .A(n8314), .B(n4502), .ZN(n6193) );
  XNOR2_X1 U7805 ( .A(n6202), .B(P2_REG3_REG_27__SCAN_IN), .ZN(n8095) );
  NAND2_X1 U7806 ( .A1(n8095), .A2(n6185), .ZN(n6191) );
  INV_X1 U7807 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n6188) );
  NAND2_X1 U7808 ( .A1(n6263), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n6187) );
  NAND2_X1 U7809 ( .A1(n7677), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n6186) );
  OAI211_X1 U7810 ( .C1(n6188), .C2(n6266), .A(n6187), .B(n6186), .ZN(n6189)
         );
  INV_X1 U7811 ( .A(n6189), .ZN(n6190) );
  NAND2_X1 U7812 ( .A1(n8087), .A2(n6783), .ZN(n6192) );
  NOR2_X1 U7813 ( .A1(n6193), .A2(n6192), .ZN(n6194) );
  AOI21_X1 U7814 ( .B1(n6193), .B2(n6192), .A(n6194), .ZN(n7538) );
  INV_X1 U7815 ( .A(n6194), .ZN(n6195) );
  NAND2_X1 U7816 ( .A1(n7537), .A2(n6195), .ZN(n6256) );
  NAND2_X1 U7817 ( .A1(n7527), .A2(n7701), .ZN(n6197) );
  NAND2_X1 U7818 ( .A1(n7702), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n6196) );
  NOR2_X1 U7819 ( .A1(n8083), .A2(n8379), .ZN(n6214) );
  INV_X1 U7820 ( .A(n6214), .ZN(n6212) );
  INV_X1 U7821 ( .A(n8083), .ZN(n8309) );
  INV_X1 U7822 ( .A(n6202), .ZN(n6199) );
  AND2_X1 U7823 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(P2_REG3_REG_28__SCAN_IN), 
        .ZN(n6198) );
  NAND2_X1 U7824 ( .A1(n6199), .A2(n6198), .ZN(n8071) );
  INV_X1 U7825 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n6201) );
  INV_X1 U7826 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n6200) );
  OAI21_X1 U7827 ( .B1(n6202), .B2(n6201), .A(n6200), .ZN(n6203) );
  NAND2_X1 U7828 ( .A1(n8071), .A2(n6203), .ZN(n6271) );
  INV_X1 U7829 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n6206) );
  NAND2_X1 U7830 ( .A1(n6263), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n6205) );
  NAND2_X1 U7831 ( .A1(n7677), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n6204) );
  OAI211_X1 U7832 ( .C1(n6206), .C2(n6266), .A(n6205), .B(n6204), .ZN(n6207)
         );
  INV_X1 U7833 ( .A(n6207), .ZN(n6208) );
  NAND2_X1 U7834 ( .A1(n8100), .A2(n6783), .ZN(n6211) );
  XNOR2_X1 U7835 ( .A(n6211), .B(n6210), .ZN(n6213) );
  MUX2_X1 U7836 ( .A(n6212), .B(n8309), .S(n6213), .Z(n6255) );
  MUX2_X1 U7837 ( .A(n8083), .B(n6214), .S(n6213), .Z(n6215) );
  NAND2_X1 U7838 ( .A1(n6256), .A2(n6215), .ZN(n6254) );
  NAND2_X1 U7839 ( .A1(n4343), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6216) );
  MUX2_X1 U7840 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6216), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n6218) );
  NAND2_X1 U7841 ( .A1(n6219), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6220) );
  MUX2_X1 U7842 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6220), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n6221) );
  NAND2_X1 U7843 ( .A1(n6221), .A2(n4343), .ZN(n7480) );
  XNOR2_X1 U7844 ( .A(n7405), .B(P2_B_REG_SCAN_IN), .ZN(n6227) );
  NAND2_X1 U7845 ( .A1(n7480), .A2(n6227), .ZN(n6228) );
  INV_X1 U7846 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n9673) );
  AND2_X1 U7847 ( .A1(n7480), .A2(n8419), .ZN(n9674) );
  NOR4_X1 U7848 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_18__SCAN_IN), .A3(
        P2_D_REG_19__SCAN_IN), .A4(P2_D_REG_21__SCAN_IN), .ZN(n6232) );
  NOR4_X1 U7849 ( .A1(P2_D_REG_14__SCAN_IN), .A2(P2_D_REG_12__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_15__SCAN_IN), .ZN(n6231) );
  NOR4_X1 U7850 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n6230) );
  NOR4_X1 U7851 ( .A1(P2_D_REG_22__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n6229) );
  NAND4_X1 U7852 ( .A1(n6232), .A2(n6231), .A3(n6230), .A4(n6229), .ZN(n6238)
         );
  NOR2_X1 U7853 ( .A1(P2_D_REG_20__SCAN_IN), .A2(P2_D_REG_4__SCAN_IN), .ZN(
        n6236) );
  NOR4_X1 U7854 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_11__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n6235) );
  NOR4_X1 U7855 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_8__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_10__SCAN_IN), .ZN(n6234) );
  NOR4_X1 U7856 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_6__SCAN_IN), .ZN(n6233) );
  NAND4_X1 U7857 ( .A1(n6236), .A2(n6235), .A3(n6234), .A4(n6233), .ZN(n6237)
         );
  OAI21_X1 U7858 ( .B1(n6238), .B2(n6237), .A(n9668), .ZN(n6498) );
  AND2_X1 U7859 ( .A1(n7405), .A2(n8419), .ZN(n9672) );
  INV_X1 U7860 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n9671) );
  AND2_X1 U7861 ( .A1(n9668), .A2(n9671), .ZN(n6239) );
  AND2_X1 U7862 ( .A1(n6498), .A2(n6701), .ZN(n6240) );
  NAND2_X1 U7863 ( .A1(n6779), .A2(n6240), .ZN(n6249) );
  NAND2_X1 U7864 ( .A1(n6241), .A2(n7897), .ZN(n6781) );
  NAND2_X1 U7865 ( .A1(n6249), .A2(n6781), .ZN(n6617) );
  INV_X1 U7866 ( .A(n7480), .ZN(n6242) );
  NAND2_X1 U7867 ( .A1(n6243), .A2(n6242), .ZN(n6244) );
  OAI21_X1 U7868 ( .B1(n6247), .B2(n6246), .A(n6245), .ZN(n6321) );
  NOR2_X1 U7869 ( .A1(n9669), .A2(n9727), .ZN(n6248) );
  NAND2_X1 U7870 ( .A1(n6250), .A2(n4745), .ZN(n6324) );
  NAND2_X1 U7871 ( .A1(n9727), .A2(n6324), .ZN(n6251) );
  NOR2_X1 U7872 ( .A1(n9669), .A2(n6251), .ZN(n6252) );
  OAI21_X1 U7873 ( .B1(n8083), .B2(n7660), .A(n7673), .ZN(n6253) );
  OAI211_X1 U7874 ( .C1(n6256), .C2(n6255), .A(n6254), .B(n6253), .ZN(n6274)
         );
  INV_X1 U7875 ( .A(n9669), .ZN(n6257) );
  NAND3_X1 U7876 ( .A1(n6259), .A2(n6258), .A3(n6257), .ZN(n7655) );
  INV_X1 U7877 ( .A(n7528), .ZN(n6261) );
  AOI22_X1 U7878 ( .A1(n7643), .A2(n8087), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        n4264), .ZN(n6273) );
  OR2_X1 U7879 ( .A1(n8071), .A2(n6262), .ZN(n6269) );
  INV_X1 U7880 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n8072) );
  NAND2_X1 U7881 ( .A1(n7677), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n6265) );
  NAND2_X1 U7882 ( .A1(n6263), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n6264) );
  OAI211_X1 U7883 ( .C1(n6266), .C2(n8072), .A(n6265), .B(n6264), .ZN(n6267)
         );
  INV_X1 U7884 ( .A(n6267), .ZN(n6268) );
  NAND2_X1 U7885 ( .A1(n6269), .A2(n6268), .ZN(n8086) );
  NAND2_X1 U7886 ( .A1(n6363), .A2(n7901), .ZN(n6496) );
  NAND4_X1 U7887 ( .A1(n6617), .A2(n6360), .A3(n6321), .A4(n6496), .ZN(n6270)
         );
  INV_X1 U7888 ( .A(n6271), .ZN(n8081) );
  AOI22_X1 U7889 ( .A1(n7669), .A2(n8086), .B1(n7657), .B2(n8081), .ZN(n6272)
         );
  NAND2_X1 U7890 ( .A1(n6274), .A2(n4834), .ZN(P2_U3222) );
  OR2_X1 U7891 ( .A1(n6276), .A2(n6275), .ZN(n6278) );
  NAND2_X1 U7892 ( .A1(n6278), .A2(n6277), .ZN(n6279) );
  NAND2_X1 U7893 ( .A1(n6279), .A2(n8475), .ZN(n6285) );
  OAI22_X1 U7894 ( .A1(n8545), .A2(n8654), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9880), .ZN(n6281) );
  NOR2_X1 U7895 ( .A1(n8550), .A2(n8959), .ZN(n6280) );
  AOI211_X1 U7896 ( .C1(n8523), .C2(n8965), .A(n6281), .B(n6280), .ZN(n6282)
         );
  OAI21_X1 U7897 ( .B1(n4537), .B2(n7464), .A(n6282), .ZN(n6283) );
  INV_X1 U7898 ( .A(n6283), .ZN(n6284) );
  NAND2_X1 U7899 ( .A1(n6285), .A2(n6284), .ZN(P1_U3212) );
  INV_X1 U7900 ( .A(n9675), .ZN(n6286) );
  INV_X1 U7901 ( .A(n7374), .ZN(n6288) );
  OR2_X1 U7902 ( .A1(n8680), .A2(n6288), .ZN(n6289) );
  NAND2_X1 U7903 ( .A1(n6289), .A2(n6341), .ZN(n6343) );
  OAI21_X1 U7904 ( .B1(n6343), .B2(n6290), .A(P1_STATE_REG_SCAN_IN), .ZN(
        P1_U3083) );
  NOR2_X1 U7905 ( .A1(n7698), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8410) );
  AOI22_X1 U7906 ( .A1(n8410), .A2(P1_DATAO_REG_2__SCAN_IN), .B1(n9362), .B2(
        P2_STATE_REG_SCAN_IN), .ZN(n6291) );
  OAI21_X1 U7907 ( .B1(n6304), .B2(n8414), .A(n6291), .ZN(P2_U3356) );
  AOI22_X1 U7908 ( .A1(n8410), .A2(P1_DATAO_REG_1__SCAN_IN), .B1(n9351), .B2(
        P2_STATE_REG_SCAN_IN), .ZN(n6292) );
  OAI21_X1 U7909 ( .B1(n6302), .B2(n8414), .A(n6292), .ZN(P2_U3357) );
  INV_X2 U7910 ( .A(n8410), .ZN(n8417) );
  INV_X1 U7911 ( .A(n6373), .ZN(n7925) );
  OAI222_X1 U7912 ( .A1(n8417), .A2(n6293), .B1(n8414), .B2(n6300), .C1(n4264), 
        .C2(n7925), .ZN(P2_U3355) );
  INV_X1 U7913 ( .A(n6439), .ZN(n6432) );
  OAI222_X1 U7914 ( .A1(n8417), .A2(n6294), .B1(n8414), .B2(n6295), .C1(
        P2_U3152), .C2(n6432), .ZN(P2_U3354) );
  OAI222_X1 U7915 ( .A1(n6296), .A2(n9340), .B1(P1_U3084), .B2(n9483), .C1(
        n9343), .C2(n6295), .ZN(P1_U3349) );
  INV_X1 U7916 ( .A(n6444), .ZN(n7939) );
  OAI222_X1 U7917 ( .A1(n8417), .A2(n6297), .B1(n8414), .B2(n6298), .C1(n4264), 
        .C2(n7939), .ZN(P2_U3353) );
  OAI222_X1 U7918 ( .A1(n9340), .A2(n6299), .B1(n9343), .B2(n6298), .C1(
        P1_U3084), .C2(n8863), .ZN(P1_U3348) );
  OAI222_X1 U7919 ( .A1(n9340), .A2(n6301), .B1(n9343), .B2(n6300), .C1(
        P1_U3084), .C2(n8850), .ZN(P1_U3350) );
  INV_X1 U7920 ( .A(n9343), .ZN(n7372) );
  OAI222_X1 U7921 ( .A1(n9340), .A2(n6303), .B1(n9343), .B2(n6302), .C1(
        P1_U3084), .C2(n6582), .ZN(P1_U3352) );
  OAI222_X1 U7922 ( .A1(n9340), .A2(n6305), .B1(n9343), .B2(n6304), .C1(
        P1_U3084), .C2(n9470), .ZN(P1_U3351) );
  INV_X1 U7923 ( .A(n6445), .ZN(n6481) );
  OAI222_X1 U7924 ( .A1(n8417), .A2(n6306), .B1(n8414), .B2(n6307), .C1(
        P2_U3152), .C2(n6481), .ZN(P2_U3352) );
  OAI222_X1 U7925 ( .A1(n9340), .A2(n6308), .B1(n9343), .B2(n6307), .C1(
        P1_U3084), .C2(n6420), .ZN(P1_U3347) );
  OAI222_X1 U7926 ( .A1(n8417), .A2(n6310), .B1(n8414), .B2(n6312), .C1(n4264), 
        .C2(n6522), .ZN(P2_U3351) );
  OAI222_X1 U7927 ( .A1(n9340), .A2(n6313), .B1(n9343), .B2(n6312), .C1(
        P1_U3084), .C2(n6311), .ZN(P1_U3346) );
  NAND2_X1 U7928 ( .A1(n6314), .A2(n9577), .ZN(n6315) );
  OAI21_X1 U7929 ( .B1(n9577), .B2(n9811), .A(n6315), .ZN(P1_U3441) );
  OAI222_X1 U7930 ( .A1(n9340), .A2(n6316), .B1(n9343), .B2(n6317), .C1(
        P1_U3084), .C2(n6463), .ZN(P1_U3345) );
  INV_X1 U7931 ( .A(n7953), .ZN(n6524) );
  OAI222_X1 U7932 ( .A1(n8417), .A2(n6318), .B1(n8414), .B2(n6317), .C1(
        P2_U3152), .C2(n6524), .ZN(P2_U3350) );
  INV_X1 U7933 ( .A(n6319), .ZN(n6327) );
  INV_X1 U7934 ( .A(n9340), .ZN(n9332) );
  AOI22_X1 U7935 ( .A1(n9499), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n9332), .ZN(n6320) );
  OAI21_X1 U7936 ( .B1(n6327), .B2(n9343), .A(n6320), .ZN(P1_U3344) );
  OR2_X1 U7937 ( .A1(n6321), .A2(n6309), .ZN(n7904) );
  NAND2_X1 U7938 ( .A1(n9669), .A2(n7904), .ZN(n6323) );
  NAND2_X1 U7939 ( .A1(n6323), .A2(n6322), .ZN(n6326) );
  OR2_X1 U7940 ( .A1(n9669), .A2(n6324), .ZN(n6325) );
  NOR2_X1 U7941 ( .A1(n9633), .A2(P2_U3966), .ZN(P2_U3151) );
  INV_X1 U7942 ( .A(n6535), .ZN(n7966) );
  OAI222_X1 U7943 ( .A1(n8417), .A2(n6328), .B1(n8414), .B2(n6327), .C1(n7966), 
        .C2(n4264), .ZN(P2_U3349) );
  INV_X1 U7944 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n6334) );
  NAND2_X1 U7945 ( .A1(n6263), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n6332) );
  NAND2_X1 U7946 ( .A1(n7677), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n6331) );
  NAND2_X1 U7947 ( .A1(n6329), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n6330) );
  NAND3_X1 U7948 ( .A1(n6332), .A2(n6331), .A3(n6330), .ZN(n8039) );
  NAND2_X1 U7949 ( .A1(P2_U3966), .A2(n8039), .ZN(n6333) );
  OAI21_X1 U7950 ( .B1(P2_U3966), .B2(n6334), .A(n6333), .ZN(P2_U3583) );
  INV_X1 U7951 ( .A(n6335), .ZN(n6337) );
  INV_X1 U7952 ( .A(n6536), .ZN(n7979) );
  OAI222_X1 U7953 ( .A1(n8417), .A2(n9814), .B1(n8414), .B2(n6337), .C1(n7979), 
        .C2(P2_U3152), .ZN(P2_U3348) );
  INV_X1 U7954 ( .A(n6487), .ZN(n6405) );
  OAI222_X1 U7955 ( .A1(P1_U3084), .A2(n6405), .B1(n9343), .B2(n6337), .C1(
        n6336), .C2(n9340), .ZN(P1_U3343) );
  INV_X1 U7956 ( .A(n6660), .ZN(n6658) );
  INV_X1 U7957 ( .A(n6338), .ZN(n6340) );
  OAI222_X1 U7958 ( .A1(n4264), .A2(n6658), .B1(n8414), .B2(n6340), .C1(n6339), 
        .C2(n8417), .ZN(P2_U3347) );
  INV_X1 U7959 ( .A(n6648), .ZN(n6490) );
  OAI222_X1 U7960 ( .A1(n9340), .A2(n9828), .B1(n9343), .B2(n6340), .C1(n6490), 
        .C2(P1_U3084), .ZN(P1_U3342) );
  INV_X1 U7961 ( .A(n6341), .ZN(n6342) );
  INV_X1 U7962 ( .A(n6343), .ZN(n6344) );
  INV_X1 U7963 ( .A(n6400), .ZN(n6350) );
  NOR2_X1 U7964 ( .A1(n9337), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n6345) );
  OR2_X1 U7965 ( .A1(n6345), .A2(n5637), .ZN(n6348) );
  AOI21_X1 U7966 ( .B1(n9337), .B2(n4912), .A(P1_IR_REG_0__SCAN_IN), .ZN(n6347) );
  NAND2_X1 U7967 ( .A1(n6348), .A2(n6352), .ZN(n9461) );
  OAI211_X1 U7968 ( .C1(n6348), .C2(n6347), .A(n9461), .B(n6346), .ZN(n6349)
         );
  OAI22_X1 U7969 ( .A1(n6350), .A2(n6349), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9566), .ZN(n6354) );
  INV_X1 U7970 ( .A(n9337), .ZN(n6382) );
  OR2_X1 U7971 ( .A1(n5637), .A2(n6382), .ZN(n9467) );
  INV_X1 U7972 ( .A(n9467), .ZN(n6351) );
  NAND2_X1 U7973 ( .A1(n6400), .A2(n6351), .ZN(n9490) );
  NOR3_X1 U7974 ( .A1(n9490), .A2(P1_REG1_REG_0__SCAN_IN), .A3(n6352), .ZN(
        n6353) );
  AOI211_X1 U7975 ( .C1(P1_ADDR_REG_0__SCAN_IN), .C2(n9539), .A(n6354), .B(
        n6353), .ZN(n6355) );
  INV_X1 U7976 ( .A(n6355), .ZN(P1_U3241) );
  INV_X1 U7977 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n6356) );
  MUX2_X1 U7978 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n6356), .S(n6373), .Z(n7921)
         );
  NAND2_X1 U7979 ( .A1(n9362), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6359) );
  INV_X1 U7980 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n6357) );
  MUX2_X1 U7981 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n6357), .S(n9362), .Z(n9365)
         );
  NAND2_X1 U7982 ( .A1(n9351), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n6358) );
  NAND2_X1 U7983 ( .A1(n6358), .A2(n9352), .ZN(n9366) );
  NAND2_X1 U7984 ( .A1(n9365), .A2(n9366), .ZN(n9364) );
  NAND2_X1 U7985 ( .A1(n6359), .A2(n9364), .ZN(n7922) );
  NAND2_X1 U7986 ( .A1(n7921), .A2(n7922), .ZN(n7920) );
  INV_X1 U7987 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n6914) );
  MUX2_X1 U7988 ( .A(n6914), .B(P2_REG2_REG_4__SCAN_IN), .S(n6439), .Z(n6366)
         );
  INV_X1 U7989 ( .A(n6360), .ZN(n6361) );
  NAND2_X1 U7990 ( .A1(n6361), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6362) );
  OAI211_X1 U7991 ( .C1(n9669), .C2(n6363), .A(n7904), .B(n6362), .ZN(n6365)
         );
  NAND2_X1 U7992 ( .A1(n6365), .A2(n6364), .ZN(n6370) );
  NAND2_X1 U7993 ( .A1(n6370), .A2(n7906), .ZN(n6368) );
  INV_X1 U7994 ( .A(n8413), .ZN(n6369) );
  NAND2_X1 U7995 ( .A1(n6368), .A2(n6369), .ZN(n8033) );
  AOI211_X1 U7996 ( .C1(n6367), .C2(n6366), .A(n6431), .B(n8029), .ZN(n6381)
         );
  XNOR2_X1 U7997 ( .A(n6439), .B(P2_REG1_REG_4__SCAN_IN), .ZN(n6375) );
  INV_X1 U7998 ( .A(n9638), .ZN(n9636) );
  INV_X1 U7999 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n9737) );
  XNOR2_X1 U8000 ( .A(n9351), .B(P2_REG1_REG_1__SCAN_IN), .ZN(n9348) );
  NOR3_X1 U8001 ( .A1(n9636), .A2(n9737), .A3(n9348), .ZN(n9347) );
  AOI21_X1 U8002 ( .B1(n9351), .B2(P2_REG1_REG_1__SCAN_IN), .A(n9347), .ZN(
        n9360) );
  XNOR2_X1 U8003 ( .A(n9362), .B(P2_REG1_REG_2__SCAN_IN), .ZN(n9359) );
  NOR2_X1 U8004 ( .A1(n9360), .A2(n9359), .ZN(n9358) );
  AOI21_X1 U8005 ( .B1(n9362), .B2(P2_REG1_REG_2__SCAN_IN), .A(n9358), .ZN(
        n7928) );
  OR2_X1 U8006 ( .A1(n6373), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6372) );
  NAND2_X1 U8007 ( .A1(n6373), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6371) );
  NAND2_X1 U8008 ( .A1(n6372), .A2(n6371), .ZN(n7927) );
  NOR2_X1 U8009 ( .A1(n7928), .A2(n7927), .ZN(n7926) );
  AOI21_X1 U8010 ( .B1(n6373), .B2(P2_REG1_REG_3__SCAN_IN), .A(n7926), .ZN(
        n6374) );
  OR2_X1 U8011 ( .A1(n6375), .A2(n6374), .ZN(n6441) );
  NAND2_X1 U8012 ( .A1(n6375), .A2(n6374), .ZN(n6376) );
  NAND3_X1 U8013 ( .A1(n9627), .A2(n6441), .A3(n6376), .ZN(n6379) );
  NAND2_X1 U8014 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3152), .ZN(n6726) );
  INV_X1 U8015 ( .A(n6726), .ZN(n6377) );
  AOI21_X1 U8016 ( .B1(n9633), .B2(P2_ADDR_REG_4__SCAN_IN), .A(n6377), .ZN(
        n6378) );
  OAI211_X1 U8017 ( .C1(n9628), .C2(n6432), .A(n6379), .B(n6378), .ZN(n6380)
         );
  OR2_X1 U8018 ( .A1(n6381), .A2(n6380), .ZN(P2_U3249) );
  AND2_X1 U8019 ( .A1(n5637), .A2(n6382), .ZN(n6383) );
  INV_X1 U8020 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n7363) );
  XNOR2_X1 U8021 ( .A(n6487), .B(n7363), .ZN(n6403) );
  NAND2_X1 U8022 ( .A1(n9499), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6398) );
  NOR2_X1 U8023 ( .A1(P1_REG2_REG_7__SCAN_IN), .A2(n6603), .ZN(n6394) );
  MUX2_X1 U8024 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n5071), .S(n6603), .Z(n6384)
         );
  INV_X1 U8025 ( .A(n6384), .ZN(n6594) );
  MUX2_X1 U8026 ( .A(n6389), .B(P1_REG2_REG_3__SCAN_IN), .S(n8850), .Z(n8858)
         );
  XNOR2_X1 U8027 ( .A(n9470), .B(P1_REG2_REG_2__SCAN_IN), .ZN(n9472) );
  XNOR2_X1 U8028 ( .A(n6582), .B(P1_REG2_REG_1__SCAN_IN), .ZN(n6587) );
  AND2_X1 U8029 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n6385) );
  NAND2_X1 U8030 ( .A1(n6587), .A2(n6385), .ZN(n6586) );
  INV_X1 U8031 ( .A(n6582), .ZN(n6411) );
  NAND2_X1 U8032 ( .A1(n6411), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6386) );
  NAND2_X1 U8033 ( .A1(n6586), .A2(n6386), .ZN(n9471) );
  NAND2_X1 U8034 ( .A1(n9472), .A2(n9471), .ZN(n6388) );
  INV_X1 U8035 ( .A(n9470), .ZN(n6413) );
  NAND2_X1 U8036 ( .A1(n6413), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6387) );
  NAND2_X1 U8037 ( .A1(n6388), .A2(n6387), .ZN(n8857) );
  NAND2_X1 U8038 ( .A1(n8858), .A2(n8857), .ZN(n8856) );
  OR2_X1 U8039 ( .A1(n8850), .A2(n6389), .ZN(n6390) );
  NAND2_X1 U8040 ( .A1(n8856), .A2(n6390), .ZN(n9486) );
  MUX2_X1 U8041 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n6391), .S(n9483), .Z(n9485)
         );
  AND2_X1 U8042 ( .A1(n9483), .A2(n6391), .ZN(n8870) );
  OR2_X1 U8043 ( .A1(n9484), .A2(n8870), .ZN(n6392) );
  MUX2_X1 U8044 ( .A(n7224), .B(P1_REG2_REG_5__SCAN_IN), .S(n8863), .Z(n8871)
         );
  NAND2_X1 U8045 ( .A1(n6392), .A2(n8871), .ZN(n8869) );
  NAND2_X1 U8046 ( .A1(n8863), .A2(n7224), .ZN(n6393) );
  NAND2_X1 U8047 ( .A1(n8869), .A2(n6393), .ZN(n6571) );
  MUX2_X1 U8048 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n5041), .S(n6420), .Z(n6570)
         );
  NOR2_X1 U8049 ( .A1(n6594), .A2(n6595), .ZN(n6593) );
  NAND2_X1 U8050 ( .A1(n6463), .A2(n6395), .ZN(n6396) );
  NOR2_X1 U8051 ( .A1(n6463), .A2(n6395), .ZN(n6460) );
  AOI21_X1 U8052 ( .B1(n6461), .B2(n6396), .A(n6460), .ZN(n9506) );
  OAI21_X1 U8053 ( .B1(n9499), .B2(P1_REG2_REG_9__SCAN_IN), .A(n6398), .ZN(
        n9505) );
  NOR2_X1 U8054 ( .A1(n9506), .A2(n9505), .ZN(n9504) );
  INV_X1 U8055 ( .A(n9504), .ZN(n6397) );
  NAND2_X1 U8056 ( .A1(n6398), .A2(n6397), .ZN(n6402) );
  OR2_X1 U8057 ( .A1(n5637), .A2(n9337), .ZN(n9463) );
  INV_X1 U8058 ( .A(n9463), .ZN(n6399) );
  INV_X1 U8059 ( .A(n6486), .ZN(n6401) );
  OAI211_X1 U8060 ( .C1(n6403), .C2(n6402), .A(n9530), .B(n6401), .ZN(n6404)
         );
  NAND2_X1 U8061 ( .A1(P1_U3084), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n7409) );
  OAI211_X1 U8062 ( .C1(n9533), .C2(n6405), .A(n6404), .B(n7409), .ZN(n6406)
         );
  AOI21_X1 U8063 ( .B1(n9539), .B2(P1_ADDR_REG_10__SCAN_IN), .A(n6406), .ZN(
        n6427) );
  MUX2_X1 U8064 ( .A(n6407), .B(P1_REG1_REG_8__SCAN_IN), .S(n6456), .Z(n6465)
         );
  NOR2_X1 U8065 ( .A1(P1_REG1_REG_7__SCAN_IN), .A2(n6603), .ZN(n6408) );
  AOI21_X1 U8066 ( .B1(n6603), .B2(P1_REG1_REG_7__SCAN_IN), .A(n6408), .ZN(
        n6597) );
  INV_X1 U8067 ( .A(n6420), .ZN(n6575) );
  INV_X1 U8068 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6409) );
  OR2_X1 U8069 ( .A1(n8850), .A2(n6409), .ZN(n6415) );
  NAND2_X1 U8070 ( .A1(n8850), .A2(n6409), .ZN(n6410) );
  AND2_X1 U8071 ( .A1(n6415), .A2(n6410), .ZN(n8855) );
  XNOR2_X1 U8072 ( .A(n9470), .B(P1_REG1_REG_2__SCAN_IN), .ZN(n9475) );
  XNOR2_X1 U8073 ( .A(n6582), .B(P1_REG1_REG_1__SCAN_IN), .ZN(n6585) );
  AND2_X1 U8074 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n6584) );
  NAND2_X1 U8075 ( .A1(n6585), .A2(n6584), .ZN(n6583) );
  NAND2_X1 U8076 ( .A1(n6411), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6412) );
  NAND2_X1 U8077 ( .A1(n6583), .A2(n6412), .ZN(n9474) );
  NAND2_X1 U8078 ( .A1(n9475), .A2(n9474), .ZN(n9473) );
  NAND2_X1 U8079 ( .A1(n6413), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6414) );
  NAND2_X1 U8080 ( .A1(n9473), .A2(n6414), .ZN(n8854) );
  NAND2_X1 U8081 ( .A1(n8855), .A2(n8854), .ZN(n8853) );
  NAND2_X1 U8082 ( .A1(n8853), .A2(n6415), .ZN(n9488) );
  XNOR2_X1 U8083 ( .A(n9483), .B(n6416), .ZN(n9489) );
  NOR2_X1 U8084 ( .A1(n9488), .A2(n9489), .ZN(n9487) );
  AND2_X1 U8085 ( .A1(n9483), .A2(n6416), .ZN(n6417) );
  NOR2_X1 U8086 ( .A1(n9487), .A2(n6417), .ZN(n8867) );
  XNOR2_X1 U8087 ( .A(n8863), .B(P1_REG1_REG_5__SCAN_IN), .ZN(n8868) );
  NAND2_X1 U8088 ( .A1(n8867), .A2(n8868), .ZN(n8866) );
  OR2_X1 U8089 ( .A1(n8863), .A2(n6418), .ZN(n6419) );
  NAND2_X1 U8090 ( .A1(n8866), .A2(n6419), .ZN(n6564) );
  MUX2_X1 U8091 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n5039), .S(n6420), .Z(n6565)
         );
  OR2_X1 U8092 ( .A1(n6564), .A2(n6565), .ZN(n6566) );
  OAI21_X1 U8093 ( .B1(P1_REG1_REG_6__SCAN_IN), .B2(n6575), .A(n6566), .ZN(
        n6598) );
  NAND2_X1 U8094 ( .A1(n6597), .A2(n6598), .ZN(n6596) );
  OAI21_X1 U8095 ( .B1(n6603), .B2(P1_REG1_REG_7__SCAN_IN), .A(n6596), .ZN(
        n6466) );
  NOR2_X1 U8096 ( .A1(n6465), .A2(n6466), .ZN(n6464) );
  AOI21_X1 U8097 ( .B1(P1_REG1_REG_8__SCAN_IN), .B2(n6456), .A(n6464), .ZN(
        n9502) );
  NOR2_X1 U8098 ( .A1(n9499), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6421) );
  AOI21_X1 U8099 ( .B1(P1_REG1_REG_9__SCAN_IN), .B2(n9499), .A(n6421), .ZN(
        n9501) );
  NAND2_X1 U8100 ( .A1(n9502), .A2(n9501), .ZN(n9500) );
  OAI21_X1 U8101 ( .B1(n9499), .B2(P1_REG1_REG_9__SCAN_IN), .A(n9500), .ZN(
        n6424) );
  MUX2_X1 U8102 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n6422), .S(n6487), .Z(n6423)
         );
  NAND2_X1 U8103 ( .A1(n6424), .A2(n6423), .ZN(n6482) );
  OAI21_X1 U8104 ( .B1(n6424), .B2(n6423), .A(n6482), .ZN(n6425) );
  INV_X1 U8105 ( .A(n9490), .ZN(n9540) );
  NAND2_X1 U8106 ( .A1(n6425), .A2(n9540), .ZN(n6426) );
  NAND2_X1 U8107 ( .A1(n6427), .A2(n6426), .ZN(P1_U3251) );
  INV_X1 U8108 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n6428) );
  MUX2_X1 U8109 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n6428), .S(n6445), .Z(n6477)
         );
  NAND2_X1 U8110 ( .A1(n6444), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n6433) );
  INV_X1 U8111 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n6429) );
  MUX2_X1 U8112 ( .A(n6429), .B(P2_REG2_REG_5__SCAN_IN), .S(n6444), .Z(n6430)
         );
  INV_X1 U8113 ( .A(n6430), .ZN(n7936) );
  NAND2_X1 U8114 ( .A1(n7936), .A2(n7935), .ZN(n7934) );
  NAND2_X1 U8115 ( .A1(n6433), .A2(n7934), .ZN(n6478) );
  NAND2_X1 U8116 ( .A1(n6477), .A2(n6478), .ZN(n6476) );
  INV_X1 U8117 ( .A(n6476), .ZN(n6434) );
  INV_X1 U8118 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n6435) );
  MUX2_X1 U8119 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n6435), .S(n6522), .Z(n6437)
         );
  INV_X1 U8120 ( .A(n6521), .ZN(n6436) );
  AOI211_X1 U8121 ( .C1(n6438), .C2(n6437), .A(n6436), .B(n8029), .ZN(n6455)
         );
  XNOR2_X1 U8122 ( .A(n6522), .B(P2_REG1_REG_7__SCAN_IN), .ZN(n6450) );
  NAND2_X1 U8123 ( .A1(n6445), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6448) );
  NAND2_X1 U8124 ( .A1(n6439), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6440) );
  NAND2_X1 U8125 ( .A1(n6441), .A2(n6440), .ZN(n7942) );
  OR2_X1 U8126 ( .A1(n6444), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6443) );
  NAND2_X1 U8127 ( .A1(n6444), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6442) );
  AND2_X1 U8128 ( .A1(n6443), .A2(n6442), .ZN(n7943) );
  AND2_X1 U8129 ( .A1(n7942), .A2(n7943), .ZN(n7940) );
  AOI21_X1 U8130 ( .B1(P2_REG1_REG_5__SCAN_IN), .B2(n6444), .A(n7940), .ZN(
        n6473) );
  INV_X1 U8131 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n6446) );
  MUX2_X1 U8132 ( .A(n6446), .B(P2_REG1_REG_6__SCAN_IN), .S(n6445), .Z(n6472)
         );
  NOR2_X1 U8133 ( .A1(n6473), .A2(n6472), .ZN(n6471) );
  INV_X1 U8134 ( .A(n6471), .ZN(n6447) );
  NAND2_X1 U8135 ( .A1(n6448), .A2(n6447), .ZN(n6449) );
  NAND2_X1 U8136 ( .A1(n6450), .A2(n6449), .ZN(n6532) );
  OAI211_X1 U8137 ( .C1(n6450), .C2(n6449), .A(n9627), .B(n6532), .ZN(n6453)
         );
  NOR2_X1 U8138 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5899), .ZN(n6451) );
  AOI21_X1 U8139 ( .B1(n9633), .B2(P2_ADDR_REG_7__SCAN_IN), .A(n6451), .ZN(
        n6452) );
  OAI211_X1 U8140 ( .C1(n9628), .C2(n6522), .A(n6453), .B(n6452), .ZN(n6454)
         );
  OR2_X1 U8141 ( .A1(n6455), .A2(n6454), .ZN(P2_U3252) );
  XNOR2_X1 U8142 ( .A(n6461), .B(n6395), .ZN(n6458) );
  NOR2_X1 U8143 ( .A1(n6461), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6457) );
  MUX2_X1 U8144 ( .A(n6458), .B(n6457), .S(n6456), .Z(n6459) );
  AOI21_X1 U8145 ( .B1(n6461), .B2(n6460), .A(n6459), .ZN(n6470) );
  INV_X1 U8146 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n6462) );
  OR2_X1 U8147 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6462), .ZN(n7330) );
  OAI21_X1 U8148 ( .B1(n9533), .B2(n6463), .A(n7330), .ZN(n6468) );
  AOI211_X1 U8149 ( .C1(n6466), .C2(n6465), .A(n6464), .B(n9490), .ZN(n6467)
         );
  AOI211_X1 U8150 ( .C1(P1_ADDR_REG_8__SCAN_IN), .C2(n9539), .A(n6468), .B(
        n6467), .ZN(n6469) );
  OAI21_X1 U8151 ( .B1(n6470), .B2(n9503), .A(n6469), .ZN(P1_U3249) );
  NAND2_X1 U8152 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3152), .ZN(n6715) );
  INV_X1 U8153 ( .A(n6715), .ZN(n6475) );
  AOI211_X1 U8154 ( .C1(n6473), .C2(n6472), .A(n6471), .B(n9629), .ZN(n6474)
         );
  AOI211_X1 U8155 ( .C1(P2_ADDR_REG_6__SCAN_IN), .C2(n9633), .A(n6475), .B(
        n6474), .ZN(n6480) );
  OAI211_X1 U8156 ( .C1(n6478), .C2(n6477), .A(n9632), .B(n6476), .ZN(n6479)
         );
  OAI211_X1 U8157 ( .C1(n9628), .C2(n6481), .A(n6480), .B(n6479), .ZN(P2_U3251) );
  INV_X1 U8158 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n6495) );
  OAI21_X1 U8159 ( .B1(P1_REG1_REG_10__SCAN_IN), .B2(n6487), .A(n6482), .ZN(
        n6484) );
  AOI22_X1 U8160 ( .A1(P1_REG1_REG_11__SCAN_IN), .A2(n6648), .B1(n6490), .B2(
        n5183), .ZN(n6483) );
  NAND2_X1 U8161 ( .A1(n6483), .A2(n6484), .ZN(n6640) );
  OAI21_X1 U8162 ( .B1(n6484), .B2(n6483), .A(n6640), .ZN(n6485) );
  NAND2_X1 U8163 ( .A1(n6485), .A2(n9540), .ZN(n6494) );
  AOI22_X1 U8164 ( .A1(P1_REG2_REG_11__SCAN_IN), .A2(n6648), .B1(n6490), .B2(
        n5187), .ZN(n6488) );
  NAND2_X1 U8165 ( .A1(n6488), .A2(n6489), .ZN(n6647) );
  OAI21_X1 U8166 ( .B1(n6489), .B2(n6488), .A(n6647), .ZN(n6492) );
  NAND2_X1 U8167 ( .A1(P1_U3084), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n7458) );
  OAI21_X1 U8168 ( .B1(n9533), .B2(n6490), .A(n7458), .ZN(n6491) );
  AOI21_X1 U8169 ( .B1(n9530), .B2(n6492), .A(n6491), .ZN(n6493) );
  OAI211_X1 U8170 ( .C1(n9525), .C2(n6495), .A(n6494), .B(n6493), .ZN(P1_U3252) );
  INV_X1 U8171 ( .A(n6496), .ZN(n6497) );
  NOR2_X1 U8172 ( .A1(n9669), .A2(n6497), .ZN(n6616) );
  NAND2_X1 U8173 ( .A1(n6498), .A2(n6616), .ZN(n6777) );
  INV_X1 U8174 ( .A(n6781), .ZN(n6499) );
  NOR2_X1 U8175 ( .A1(n6777), .A2(n6499), .ZN(n6501) );
  INV_X1 U8176 ( .A(n6779), .ZN(n6500) );
  AND2_X1 U8177 ( .A1(n6501), .A2(n6500), .ZN(n6702) );
  INV_X1 U8178 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n6516) );
  NAND2_X1 U8179 ( .A1(n7919), .A2(n6900), .ZN(n6502) );
  OAI21_X1 U8180 ( .B1(n7868), .B2(n6502), .A(n6554), .ZN(n7006) );
  INV_X1 U8181 ( .A(n7006), .ZN(n6514) );
  XNOR2_X1 U8182 ( .A(n6250), .B(n6503), .ZN(n6504) );
  NAND2_X1 U8183 ( .A1(n6506), .A2(n7725), .ZN(n7719) );
  INV_X1 U8184 ( .A(n7718), .ZN(n7726) );
  INV_X1 U8185 ( .A(n6506), .ZN(n6896) );
  NAND2_X1 U8186 ( .A1(n7868), .A2(n6896), .ZN(n6508) );
  OR2_X1 U8187 ( .A1(n7865), .A2(n4266), .ZN(n7708) );
  OAI211_X1 U8188 ( .C1(n7719), .C2(n7726), .A(n6508), .B(n8213), .ZN(n6510)
         );
  AOI22_X1 U8189 ( .A1(n9656), .A2(n7919), .B1(n7917), .B2(n9653), .ZN(n6509)
         );
  NAND2_X1 U8190 ( .A1(n6510), .A2(n6509), .ZN(n6999) );
  INV_X1 U8191 ( .A(n6999), .ZN(n6513) );
  AND2_X1 U8192 ( .A1(n6900), .A2(n4703), .ZN(n6511) );
  NOR2_X1 U8193 ( .A1(n6556), .A2(n6511), .ZN(n7001) );
  INV_X1 U8194 ( .A(n7865), .ZN(n7862) );
  AOI22_X1 U8195 ( .A1(n7001), .A2(n8380), .B1(n8379), .B2(n4703), .ZN(n6512)
         );
  OAI211_X1 U8196 ( .C1(n6514), .C2(n9678), .A(n6513), .B(n6512), .ZN(n8387)
         );
  NAND2_X1 U8197 ( .A1(n9736), .A2(n8387), .ZN(n6515) );
  OAI21_X1 U8198 ( .B1(n9736), .B2(n6516), .A(n6515), .ZN(P2_U3454) );
  NAND2_X1 U8199 ( .A1(n6536), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n6526) );
  INV_X1 U8200 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n6517) );
  MUX2_X1 U8201 ( .A(n6517), .B(P2_REG2_REG_10__SCAN_IN), .S(n6536), .Z(n6518)
         );
  INV_X1 U8202 ( .A(n6518), .ZN(n7976) );
  NAND2_X1 U8203 ( .A1(n6535), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n6525) );
  INV_X1 U8204 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n6519) );
  MUX2_X1 U8205 ( .A(n6519), .B(P2_REG2_REG_9__SCAN_IN), .S(n6535), .Z(n6520)
         );
  INV_X1 U8206 ( .A(n6520), .ZN(n7962) );
  INV_X1 U8207 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n6523) );
  MUX2_X1 U8208 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n6523), .S(n7953), .Z(n7949)
         );
  OAI21_X1 U8209 ( .B1(n6524), .B2(n6523), .A(n7948), .ZN(n7963) );
  NAND2_X1 U8210 ( .A1(n7962), .A2(n7963), .ZN(n7961) );
  NAND2_X1 U8211 ( .A1(n6525), .A2(n7961), .ZN(n7977) );
  NAND2_X1 U8212 ( .A1(n7976), .A2(n7977), .ZN(n7975) );
  NAND2_X1 U8213 ( .A1(n6526), .A2(n7975), .ZN(n6529) );
  INV_X1 U8214 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n6527) );
  MUX2_X1 U8215 ( .A(n6527), .B(P2_REG2_REG_11__SCAN_IN), .S(n6660), .Z(n6528)
         );
  AOI21_X1 U8216 ( .B1(n6529), .B2(n6528), .A(n6657), .ZN(n6548) );
  INV_X1 U8217 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n9748) );
  MUX2_X1 U8218 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n9748), .S(n6660), .Z(n6541)
         );
  NAND2_X1 U8219 ( .A1(n6536), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n6539) );
  NAND2_X1 U8220 ( .A1(n6530), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6531) );
  NAND2_X1 U8221 ( .A1(n6532), .A2(n6531), .ZN(n7955) );
  INV_X1 U8222 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n9744) );
  MUX2_X1 U8223 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n9744), .S(n7953), .Z(n7956)
         );
  NAND2_X1 U8224 ( .A1(n7955), .A2(n7956), .ZN(n7954) );
  NAND2_X1 U8225 ( .A1(n7953), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n6533) );
  AND2_X1 U8226 ( .A1(n7954), .A2(n6533), .ZN(n7969) );
  INV_X1 U8227 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n6534) );
  MUX2_X1 U8228 ( .A(n6534), .B(P2_REG1_REG_9__SCAN_IN), .S(n6535), .Z(n7968)
         );
  NOR2_X1 U8229 ( .A1(n7969), .A2(n7968), .ZN(n7967) );
  AOI21_X1 U8230 ( .B1(n6535), .B2(P2_REG1_REG_9__SCAN_IN), .A(n7967), .ZN(
        n7981) );
  INV_X1 U8231 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n6537) );
  MUX2_X1 U8232 ( .A(n6537), .B(P2_REG1_REG_10__SCAN_IN), .S(n6536), .Z(n7982)
         );
  NOR2_X1 U8233 ( .A1(n7981), .A2(n7982), .ZN(n7980) );
  INV_X1 U8234 ( .A(n7980), .ZN(n6538) );
  NAND2_X1 U8235 ( .A1(n6539), .A2(n6538), .ZN(n6540) );
  NAND2_X1 U8236 ( .A1(n6541), .A2(n6540), .ZN(n6662) );
  OAI211_X1 U8237 ( .C1(n6541), .C2(n6540), .A(n9627), .B(n6662), .ZN(n6545)
         );
  NOR2_X1 U8238 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6542), .ZN(n6543) );
  AOI21_X1 U8239 ( .B1(n9633), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n6543), .ZN(
        n6544) );
  OAI211_X1 U8240 ( .C1(n9628), .C2(n6658), .A(n6545), .B(n6544), .ZN(n6546)
         );
  INV_X1 U8241 ( .A(n6546), .ZN(n6547) );
  OAI21_X1 U8242 ( .B1(n6548), .B2(n8029), .A(n6547), .ZN(P2_U3256) );
  INV_X1 U8243 ( .A(n6549), .ZN(n6551) );
  INV_X1 U8244 ( .A(n6738), .ZN(n6670) );
  OAI222_X1 U8245 ( .A1(n8417), .A2(n6550), .B1(n8414), .B2(n6551), .C1(n4264), 
        .C2(n6670), .ZN(P2_U3346) );
  INV_X1 U8246 ( .A(n6765), .ZN(n6646) );
  OAI222_X1 U8247 ( .A1(n9340), .A2(n6552), .B1(n9343), .B2(n6551), .C1(
        P1_U3084), .C2(n6646), .ZN(P1_U3341) );
  INV_X1 U8248 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n9891) );
  INV_X1 U8249 ( .A(n7918), .ZN(n6897) );
  NAND2_X1 U8250 ( .A1(n6897), .A2(n7003), .ZN(n6553) );
  NAND2_X1 U8251 ( .A1(n6554), .A2(n6553), .ZN(n6555) );
  NAND2_X1 U8252 ( .A1(n7917), .A2(n6968), .ZN(n7728) );
  NAND2_X1 U8253 ( .A1(n6555), .A2(n7867), .ZN(n6687) );
  OAI21_X1 U8254 ( .B1(n6555), .B2(n7867), .A(n6687), .ZN(n6965) );
  INV_X1 U8255 ( .A(n6965), .ZN(n6562) );
  INV_X1 U8256 ( .A(n6556), .ZN(n6557) );
  AOI211_X1 U8257 ( .C1(n4361), .C2(n6557), .A(n9728), .B(n4466), .ZN(n6958)
         );
  AOI21_X1 U8258 ( .B1(n8379), .B2(n4361), .A(n6958), .ZN(n6561) );
  NAND2_X1 U8259 ( .A1(n7719), .A2(n7718), .ZN(n6690) );
  XNOR2_X1 U8260 ( .A(n6690), .B(n7867), .ZN(n6560) );
  NAND2_X1 U8261 ( .A1(n7916), .A2(n9653), .ZN(n6559) );
  NAND2_X1 U8262 ( .A1(n7918), .A2(n9656), .ZN(n6558) );
  NAND2_X1 U8263 ( .A1(n6559), .A2(n6558), .ZN(n6618) );
  AOI21_X1 U8264 ( .B1(n6560), .B2(n8213), .A(n6618), .ZN(n6962) );
  OAI211_X1 U8265 ( .C1(n9678), .C2(n6562), .A(n6561), .B(n6962), .ZN(n8386)
         );
  NAND2_X1 U8266 ( .A1(n8386), .A2(n9736), .ZN(n6563) );
  OAI21_X1 U8267 ( .B1(n9736), .B2(n9891), .A(n6563), .ZN(P2_U3457) );
  INV_X1 U8268 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n6578) );
  INV_X1 U8269 ( .A(n6564), .ZN(n6568) );
  INV_X1 U8270 ( .A(n6565), .ZN(n6567) );
  OAI21_X1 U8271 ( .B1(n6568), .B2(n6567), .A(n6566), .ZN(n6573) );
  AOI211_X1 U8272 ( .C1(n6571), .C2(n6570), .A(n6569), .B(n9503), .ZN(n6572)
         );
  AOI21_X1 U8273 ( .B1(n9540), .B2(n6573), .A(n6572), .ZN(n6577) );
  INV_X1 U8274 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n6574) );
  NOR2_X1 U8275 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6574), .ZN(n7129) );
  AOI21_X1 U8276 ( .B1(n9514), .B2(n6575), .A(n7129), .ZN(n6576) );
  OAI211_X1 U8277 ( .C1(n9525), .C2(n6578), .A(n6577), .B(n6576), .ZN(P1_U3247) );
  NAND2_X1 U8278 ( .A1(n5653), .A2(n7100), .ZN(n8806) );
  INV_X1 U8279 ( .A(n8806), .ZN(n6579) );
  NOR2_X1 U8280 ( .A1(n7095), .A2(n6579), .ZN(n8697) );
  NAND2_X1 U8281 ( .A1(n8557), .A2(n7089), .ZN(n6580) );
  INV_X1 U8282 ( .A(n8849), .ZN(n7189) );
  OAI22_X1 U8283 ( .A1(n8697), .A2(n6580), .B1(n7189), .B2(n9440), .ZN(n9568)
         );
  NOR2_X1 U8284 ( .A1(n7100), .A2(n7089), .ZN(n9571) );
  NOR2_X1 U8285 ( .A1(n9568), .A2(n9571), .ZN(n6676) );
  NAND2_X1 U8286 ( .A1(n9625), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6581) );
  OAI21_X1 U8287 ( .B1(n6676), .B2(n9625), .A(n6581), .ZN(P1_U3523) );
  OAI22_X1 U8288 ( .A1(n9533), .A2(n6582), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n7101), .ZN(n6591) );
  OAI211_X1 U8289 ( .C1(n6585), .C2(n6584), .A(n9540), .B(n6583), .ZN(n6589)
         );
  NAND2_X1 U8290 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n9464) );
  OAI211_X1 U8291 ( .C1(n6587), .C2(n6385), .A(n9530), .B(n6586), .ZN(n6588)
         );
  NAND2_X1 U8292 ( .A1(n6589), .A2(n6588), .ZN(n6590) );
  AOI211_X1 U8293 ( .C1(n9539), .C2(P1_ADDR_REG_1__SCAN_IN), .A(n6591), .B(
        n6590), .ZN(n6592) );
  INV_X1 U8294 ( .A(n6592), .ZN(P1_U3242) );
  INV_X1 U8295 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n6605) );
  NOR2_X1 U8296 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n5072), .ZN(n7156) );
  AOI21_X1 U8297 ( .B1(n6595), .B2(n6594), .A(n6593), .ZN(n6601) );
  OAI21_X1 U8298 ( .B1(n6598), .B2(n6597), .A(n6596), .ZN(n6599) );
  NAND2_X1 U8299 ( .A1(n9540), .A2(n6599), .ZN(n6600) );
  OAI21_X1 U8300 ( .B1(n9503), .B2(n6601), .A(n6600), .ZN(n6602) );
  AOI211_X1 U8301 ( .C1(n9514), .C2(n6603), .A(n7156), .B(n6602), .ZN(n6604)
         );
  OAI21_X1 U8302 ( .B1(n9525), .B2(n6605), .A(n6604), .ZN(P1_U3248) );
  CLKBUF_X2 U8303 ( .A(P1_U4006), .Z(n9462) );
  INV_X1 U8304 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n6607) );
  NAND2_X1 U8305 ( .A1(n5653), .A2(n9462), .ZN(n6606) );
  OAI21_X1 U8306 ( .B1(n9462), .B2(n6607), .A(n6606), .ZN(P1_U3555) );
  INV_X1 U8307 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n6611) );
  INV_X1 U8308 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n9168) );
  NAND2_X1 U8309 ( .A1(n5162), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n6609) );
  INV_X1 U8310 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n9282) );
  OR2_X1 U8311 ( .A1(n4989), .A2(n9282), .ZN(n6608) );
  OAI211_X1 U8312 ( .C1(n4273), .C2(n9168), .A(n6609), .B(n6608), .ZN(n8912)
         );
  NAND2_X1 U8313 ( .A1(n8912), .A2(n9462), .ZN(n6610) );
  OAI21_X1 U8314 ( .B1(n9462), .B2(n6611), .A(n6610), .ZN(P1_U3586) );
  INV_X1 U8315 ( .A(n6612), .ZN(n6625) );
  AOI22_X1 U8316 ( .A1(n7141), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n9332), .ZN(n6613) );
  OAI21_X1 U8317 ( .B1(n6625), .B2(n9343), .A(n6613), .ZN(P1_U3340) );
  XNOR2_X1 U8318 ( .A(n6614), .B(n6615), .ZN(n6622) );
  AND2_X1 U8319 ( .A1(n6617), .A2(n6616), .ZN(n6632) );
  INV_X1 U8320 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n6959) );
  INV_X1 U8321 ( .A(n6618), .ZN(n6619) );
  OAI22_X1 U8322 ( .A1(n6632), .A2(n6959), .B1(n7655), .B2(n6619), .ZN(n6620)
         );
  AOI21_X1 U8323 ( .B1(n7670), .B2(n4361), .A(n6620), .ZN(n6621) );
  OAI21_X1 U8324 ( .B1(n6622), .B2(n7673), .A(n6621), .ZN(P2_U3239) );
  INV_X1 U8325 ( .A(n6623), .ZN(n6631) );
  AOI22_X1 U8326 ( .A1(n9513), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n9332), .ZN(n6624) );
  OAI21_X1 U8327 ( .B1(n6631), .B2(n9343), .A(n6624), .ZN(P1_U3339) );
  INV_X1 U8328 ( .A(n6845), .ZN(n6743) );
  OAI222_X1 U8329 ( .A1(n8417), .A2(n6626), .B1(n8414), .B2(n6625), .C1(n6743), 
        .C2(n4264), .ZN(P2_U3345) );
  INV_X1 U8330 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n6630) );
  AOI22_X1 U8331 ( .A1(n7669), .A2(n7918), .B1(n7670), .B2(n6900), .ZN(n6629)
         );
  NOR2_X1 U8332 ( .A1(n4524), .A2(n6900), .ZN(n7727) );
  MUX2_X1 U8333 ( .A(n6900), .B(n7727), .S(n6783), .Z(n6627) );
  OAI21_X1 U8334 ( .B1(n6896), .B2(n6627), .A(n7631), .ZN(n6628) );
  OAI211_X1 U8335 ( .C1(n6632), .C2(n6630), .A(n6629), .B(n6628), .ZN(P2_U3234) );
  INV_X1 U8336 ( .A(n6989), .ZN(n6848) );
  OAI222_X1 U8337 ( .A1(n8417), .A2(n9885), .B1(n8414), .B2(n6631), .C1(n6848), 
        .C2(P2_U3152), .ZN(P2_U3344) );
  AOI22_X1 U8338 ( .A1(n7669), .A2(n7917), .B1(n7670), .B2(n4703), .ZN(n6639)
         );
  INV_X1 U8339 ( .A(n6632), .ZN(n6637) );
  OAI21_X1 U8340 ( .B1(n6635), .B2(n6634), .A(n6633), .ZN(n6636) );
  AOI22_X1 U8341 ( .A1(n6637), .A2(P2_REG3_REG_1__SCAN_IN), .B1(n7631), .B2(
        n6636), .ZN(n6638) );
  OAI211_X1 U8342 ( .C1(n7666), .C2(n4524), .A(n6639), .B(n6638), .ZN(P2_U3224) );
  INV_X1 U8343 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n6656) );
  OAI21_X1 U8344 ( .B1(n6648), .B2(P1_REG1_REG_11__SCAN_IN), .A(n6640), .ZN(
        n6644) );
  NOR2_X1 U8345 ( .A1(n6646), .A2(n6641), .ZN(n6642) );
  AOI21_X1 U8346 ( .B1(n6641), .B2(n6646), .A(n6642), .ZN(n6643) );
  NAND2_X1 U8347 ( .A1(n6643), .A2(n6644), .ZN(n6760) );
  OAI21_X1 U8348 ( .B1(n6644), .B2(n6643), .A(n6760), .ZN(n6654) );
  NAND2_X1 U8349 ( .A1(P1_REG3_REG_12__SCAN_IN), .A2(P1_U3084), .ZN(n6645) );
  OAI21_X1 U8350 ( .B1(n9533), .B2(n6646), .A(n6645), .ZN(n6653) );
  OAI21_X1 U8351 ( .B1(n6648), .B2(P1_REG2_REG_11__SCAN_IN), .A(n6647), .ZN(
        n6651) );
  NAND2_X1 U8352 ( .A1(P1_REG2_REG_12__SCAN_IN), .A2(n6765), .ZN(n6649) );
  OAI21_X1 U8353 ( .B1(n6765), .B2(P1_REG2_REG_12__SCAN_IN), .A(n6649), .ZN(
        n6650) );
  AOI211_X1 U8354 ( .C1(n6651), .C2(n6650), .A(n6764), .B(n9503), .ZN(n6652)
         );
  AOI211_X1 U8355 ( .C1(n9540), .C2(n6654), .A(n6653), .B(n6652), .ZN(n6655)
         );
  OAI21_X1 U8356 ( .B1(n9525), .B2(n6656), .A(n6655), .ZN(P1_U3253) );
  INV_X1 U8357 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n6659) );
  MUX2_X1 U8358 ( .A(n6659), .B(P2_REG2_REG_12__SCAN_IN), .S(n6738), .Z(n6739)
         );
  XNOR2_X1 U8359 ( .A(n6741), .B(n6739), .ZN(n6672) );
  NAND2_X1 U8360 ( .A1(n6660), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n6661) );
  AND2_X1 U8361 ( .A1(n6662), .A2(n6661), .ZN(n6665) );
  INV_X1 U8362 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n6663) );
  MUX2_X1 U8363 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n6663), .S(n6738), .Z(n6664)
         );
  NAND2_X1 U8364 ( .A1(n6665), .A2(n6664), .ZN(n6733) );
  OAI21_X1 U8365 ( .B1(n6665), .B2(n6664), .A(n6733), .ZN(n6666) );
  NAND2_X1 U8366 ( .A1(n9627), .A2(n6666), .ZN(n6669) );
  NAND2_X1 U8367 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3152), .ZN(n7305) );
  INV_X1 U8368 ( .A(n7305), .ZN(n6667) );
  AOI21_X1 U8369 ( .B1(n9633), .B2(P2_ADDR_REG_12__SCAN_IN), .A(n6667), .ZN(
        n6668) );
  OAI211_X1 U8370 ( .C1(n9628), .C2(n6670), .A(n6669), .B(n6668), .ZN(n6671)
         );
  AOI21_X1 U8371 ( .B1(n6672), .B2(n9632), .A(n6671), .ZN(n6673) );
  INV_X1 U8372 ( .A(n6673), .ZN(P2_U3257) );
  INV_X1 U8373 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n6674) );
  OR2_X1 U8374 ( .A1(n9619), .A2(n6674), .ZN(n6675) );
  OAI21_X1 U8375 ( .B1(n6676), .B2(n9617), .A(n6675), .ZN(P1_U3454) );
  INV_X1 U8376 ( .A(n7088), .ZN(n6678) );
  NAND3_X1 U8377 ( .A1(n6679), .A2(n6678), .A3(n6677), .ZN(n6867) );
  AOI22_X1 U8378 ( .A1(n8552), .A2(n6680), .B1(n6867), .B2(
        P1_REG3_REG_0__SCAN_IN), .ZN(n6685) );
  OAI21_X1 U8379 ( .B1(n6683), .B2(n6681), .A(n6682), .ZN(n9468) );
  NAND2_X1 U8380 ( .A1(n9468), .A2(n8475), .ZN(n6684) );
  OAI211_X1 U8381 ( .C1(n7411), .C2(n7189), .A(n6685), .B(n6684), .ZN(P1_U3230) );
  INV_X1 U8382 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n6700) );
  NAND2_X1 U8383 ( .A1(n4362), .A2(n6968), .ZN(n6686) );
  NAND2_X1 U8384 ( .A1(n6687), .A2(n6686), .ZN(n6688) );
  NAND2_X1 U8385 ( .A1(n7916), .A2(n6792), .ZN(n7732) );
  NAND2_X1 U8386 ( .A1(n6688), .A2(n7866), .ZN(n6794) );
  OR2_X1 U8387 ( .A1(n6688), .A2(n7866), .ZN(n6689) );
  NAND2_X1 U8388 ( .A1(n6794), .A2(n6689), .ZN(n6789) );
  INV_X1 U8389 ( .A(n6789), .ZN(n6698) );
  INV_X1 U8390 ( .A(n9715), .ZN(n8384) );
  OAI21_X1 U8391 ( .B1(n6690), .B2(n7867), .A(n7724), .ZN(n6801) );
  XNOR2_X1 U8392 ( .A(n6801), .B(n7866), .ZN(n6693) );
  NAND2_X1 U8393 ( .A1(n6789), .A2(n9652), .ZN(n6692) );
  AOI22_X1 U8394 ( .A1(n9656), .A2(n7917), .B1(n7915), .B2(n9653), .ZN(n6691)
         );
  OAI211_X1 U8395 ( .C1(n9660), .C2(n6693), .A(n6692), .B(n6691), .ZN(n6787)
         );
  INV_X1 U8396 ( .A(n6787), .ZN(n6697) );
  INV_X1 U8397 ( .A(n6798), .ZN(n6916) );
  AOI21_X1 U8398 ( .B1(n6695), .B2(n6694), .A(n6916), .ZN(n6784) );
  AOI22_X1 U8399 ( .A1(n6784), .A2(n8380), .B1(n8379), .B2(n6695), .ZN(n6696)
         );
  OAI211_X1 U8400 ( .C1(n6698), .C2(n8384), .A(n6697), .B(n6696), .ZN(n6703)
         );
  NAND2_X1 U8401 ( .A1(n6703), .A2(n9736), .ZN(n6699) );
  OAI21_X1 U8402 ( .B1(n9736), .B2(n6700), .A(n6699), .ZN(P2_U3460) );
  INV_X1 U8403 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n6705) );
  NAND2_X1 U8404 ( .A1(n6703), .A2(n9752), .ZN(n6704) );
  OAI21_X1 U8405 ( .B1(n9752), .B2(n6705), .A(n6704), .ZN(P2_U3523) );
  OAI22_X1 U8406 ( .A1(n7660), .A2(n6979), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7937), .ZN(n6707) );
  INV_X1 U8407 ( .A(n7915), .ZN(n6804) );
  INV_X1 U8408 ( .A(n7913), .ZN(n7017) );
  OAI22_X1 U8409 ( .A1(n6804), .A2(n7666), .B1(n7645), .B2(n7017), .ZN(n6706)
         );
  AOI211_X1 U8410 ( .C1(n6904), .C2(n7657), .A(n6707), .B(n6706), .ZN(n6712)
         );
  OAI211_X1 U8411 ( .C1(n6710), .C2(n6709), .A(n6708), .B(n7631), .ZN(n6711)
         );
  NAND2_X1 U8412 ( .A1(n6712), .A2(n6711), .ZN(P2_U3229) );
  AOI21_X1 U8413 ( .B1(n6714), .B2(n6713), .A(n4346), .ZN(n6720) );
  INV_X1 U8414 ( .A(n9655), .ZN(n7051) );
  OAI21_X1 U8415 ( .B1(n7645), .B2(n7051), .A(n6715), .ZN(n6718) );
  INV_X1 U8416 ( .A(n7914), .ZN(n6980) );
  OAI22_X1 U8417 ( .A1(n7666), .A2(n6980), .B1(n7008), .B2(n7660), .ZN(n6717)
         );
  AOI211_X1 U8418 ( .C1(n6975), .C2(n7657), .A(n6718), .B(n6717), .ZN(n6719)
         );
  OAI21_X1 U8419 ( .B1(n6720), .B2(n7673), .A(n6719), .ZN(P2_U3241) );
  INV_X1 U8420 ( .A(n6722), .ZN(n6724) );
  NAND2_X1 U8421 ( .A1(n6724), .A2(n6723), .ZN(n6725) );
  XNOR2_X1 U8422 ( .A(n6721), .B(n6725), .ZN(n6731) );
  OAI21_X1 U8423 ( .B1(n7660), .B2(n9683), .A(n6726), .ZN(n6728) );
  OAI22_X1 U8424 ( .A1(n4698), .A2(n7666), .B1(n7645), .B2(n6980), .ZN(n6727)
         );
  AOI211_X1 U8425 ( .C1(n6729), .C2(n7657), .A(n6728), .B(n6727), .ZN(n6730)
         );
  OAI21_X1 U8426 ( .B1(n6731), .B2(n7673), .A(n6730), .ZN(P2_U3232) );
  INV_X1 U8427 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n6732) );
  AOI22_X1 U8428 ( .A1(n6845), .A2(P2_REG1_REG_13__SCAN_IN), .B1(n6732), .B2(
        n6743), .ZN(n6735) );
  OAI21_X1 U8429 ( .B1(n6738), .B2(P2_REG1_REG_12__SCAN_IN), .A(n6733), .ZN(
        n6734) );
  NAND2_X1 U8430 ( .A1(n6735), .A2(n6734), .ZN(n6840) );
  OAI21_X1 U8431 ( .B1(n6735), .B2(n6734), .A(n6840), .ZN(n6750) );
  NAND2_X1 U8432 ( .A1(n4264), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n7340) );
  INV_X1 U8433 ( .A(n7340), .ZN(n6736) );
  AOI21_X1 U8434 ( .B1(n9633), .B2(P2_ADDR_REG_13__SCAN_IN), .A(n6736), .ZN(
        n6737) );
  OAI21_X1 U8435 ( .B1(n9628), .B2(n6743), .A(n6737), .ZN(n6749) );
  NAND2_X1 U8436 ( .A1(n6738), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n6742) );
  INV_X1 U8437 ( .A(n6739), .ZN(n6740) );
  INV_X1 U8438 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n6744) );
  AOI22_X1 U8439 ( .A1(n6845), .A2(n6744), .B1(P2_REG2_REG_13__SCAN_IN), .B2(
        n6743), .ZN(n6745) );
  NOR2_X1 U8440 ( .A1(n6746), .A2(n6745), .ZN(n6846) );
  AOI21_X1 U8441 ( .B1(n6746), .B2(n6745), .A(n6846), .ZN(n6747) );
  NOR2_X1 U8442 ( .A1(n6747), .A2(n8029), .ZN(n6748) );
  AOI211_X1 U8443 ( .C1(n6750), .C2(n9627), .A(n6749), .B(n6748), .ZN(n6751)
         );
  INV_X1 U8444 ( .A(n6751), .ZN(P2_U3258) );
  XNOR2_X1 U8445 ( .A(n6752), .B(n6753), .ZN(n6757) );
  INV_X1 U8446 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n7923) );
  OAI22_X1 U8447 ( .A1(n7660), .A2(n6792), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7923), .ZN(n6755) );
  OAI22_X1 U8448 ( .A1(n4362), .A2(n7666), .B1(n7645), .B2(n6804), .ZN(n6754)
         );
  AOI211_X1 U8449 ( .C1(n7657), .C2(n7923), .A(n6755), .B(n6754), .ZN(n6756)
         );
  OAI21_X1 U8450 ( .B1(n7673), .B2(n6757), .A(n6756), .ZN(P2_U3220) );
  INV_X1 U8451 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n6773) );
  INV_X1 U8452 ( .A(n7141), .ZN(n6763) );
  NOR2_X1 U8453 ( .A1(n6763), .A2(n6758), .ZN(n6759) );
  AOI21_X1 U8454 ( .B1(n6758), .B2(n6763), .A(n6759), .ZN(n6762) );
  OAI21_X1 U8455 ( .B1(n6765), .B2(P1_REG1_REG_12__SCAN_IN), .A(n6760), .ZN(
        n6761) );
  NAND2_X1 U8456 ( .A1(n6762), .A2(n6761), .ZN(n7140) );
  OAI21_X1 U8457 ( .B1(n6762), .B2(n6761), .A(n7140), .ZN(n6771) );
  NAND2_X1 U8458 ( .A1(P1_U3084), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n7496) );
  OAI21_X1 U8459 ( .B1(n9533), .B2(n6763), .A(n7496), .ZN(n6770) );
  AOI21_X1 U8460 ( .B1(n6765), .B2(P1_REG2_REG_12__SCAN_IN), .A(n6764), .ZN(
        n6768) );
  NAND2_X1 U8461 ( .A1(P1_REG2_REG_13__SCAN_IN), .A2(n7141), .ZN(n6766) );
  OAI21_X1 U8462 ( .B1(n7141), .B2(P1_REG2_REG_13__SCAN_IN), .A(n6766), .ZN(
        n6767) );
  AOI211_X1 U8463 ( .C1(n6768), .C2(n6767), .A(n7135), .B(n9503), .ZN(n6769)
         );
  AOI211_X1 U8464 ( .C1(n9540), .C2(n6771), .A(n6770), .B(n6769), .ZN(n6772)
         );
  OAI21_X1 U8465 ( .B1(n9525), .B2(n6773), .A(n6772), .ZN(P1_U3254) );
  INV_X1 U8466 ( .A(n6774), .ZN(n6776) );
  INV_X1 U8467 ( .A(n7108), .ZN(n6994) );
  OAI222_X1 U8468 ( .A1(n8417), .A2(n6775), .B1(n8414), .B2(n6776), .C1(
        P2_U3152), .C2(n6994), .ZN(P2_U3343) );
  OAI222_X1 U8469 ( .A1(n9340), .A2(n9903), .B1(n9343), .B2(n6776), .C1(
        P1_U3084), .C2(n7290), .ZN(P1_U3338) );
  INV_X1 U8470 ( .A(n6777), .ZN(n6780) );
  NAND3_X1 U8471 ( .A1(n6780), .A2(n6779), .A3(n6778), .ZN(n6960) );
  NOR2_X1 U8472 ( .A1(n9677), .A2(n7865), .ZN(n6782) );
  OR2_X1 U8473 ( .A1(n6960), .A2(n6783), .ZN(n8290) );
  AOI22_X1 U8474 ( .A1(n9647), .A2(n6784), .B1(n9665), .B2(n7923), .ZN(n6785)
         );
  OAI21_X1 U8475 ( .B1(n6356), .B2(n9661), .A(n6785), .ZN(n6786) );
  AOI21_X1 U8476 ( .B1(n9661), .B2(n6787), .A(n6786), .ZN(n6791) );
  AND2_X1 U8477 ( .A1(n7897), .A2(n4745), .ZN(n6788) );
  NAND2_X1 U8478 ( .A1(n9648), .A2(n6789), .ZN(n6790) );
  OAI211_X1 U8479 ( .C1(n6792), .C2(n9649), .A(n6791), .B(n6790), .ZN(P2_U3293) );
  INV_X1 U8480 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n6808) );
  NAND2_X1 U8481 ( .A1(n4698), .A2(n6792), .ZN(n6793) );
  NAND2_X1 U8482 ( .A1(n6794), .A2(n6793), .ZN(n6912) );
  OR2_X1 U8483 ( .A1(n7915), .A2(n9683), .ZN(n7711) );
  NAND2_X1 U8484 ( .A1(n7915), .A2(n9683), .ZN(n7733) );
  NAND2_X1 U8485 ( .A1(n7711), .A2(n7733), .ZN(n6922) );
  NAND2_X1 U8486 ( .A1(n6912), .A2(n6922), .ZN(n6911) );
  NAND2_X1 U8487 ( .A1(n6804), .A2(n9683), .ZN(n6795) );
  OR2_X1 U8488 ( .A1(n7914), .A2(n6979), .ZN(n7715) );
  AND2_X1 U8489 ( .A1(n7914), .A2(n6979), .ZN(n7736) );
  INV_X1 U8490 ( .A(n7736), .ZN(n7712) );
  NAND2_X1 U8491 ( .A1(n7715), .A2(n7712), .ZN(n7872) );
  OAI21_X1 U8492 ( .B1(n6796), .B2(n7872), .A(n6982), .ZN(n6797) );
  INV_X1 U8493 ( .A(n6797), .ZN(n6910) );
  INV_X1 U8494 ( .A(n6979), .ZN(n6805) );
  NOR2_X1 U8495 ( .A1(n6798), .A2(n6919), .ZN(n6799) );
  INV_X1 U8496 ( .A(n6799), .ZN(n6915) );
  AOI211_X1 U8497 ( .C1(n6805), .C2(n6915), .A(n9728), .B(n6973), .ZN(n6907)
         );
  INV_X1 U8498 ( .A(n7866), .ZN(n6800) );
  NAND2_X1 U8499 ( .A1(n6801), .A2(n6800), .ZN(n6921) );
  AND2_X1 U8500 ( .A1(n7711), .A2(n6920), .ZN(n7716) );
  NAND2_X1 U8501 ( .A1(n6921), .A2(n7716), .ZN(n6802) );
  NAND2_X1 U8502 ( .A1(n6802), .A2(n7733), .ZN(n6969) );
  XOR2_X1 U8503 ( .A(n7872), .B(n6969), .Z(n6803) );
  OAI222_X1 U8504 ( .A1(n8284), .A2(n7017), .B1(n8285), .B2(n6804), .C1(n9660), 
        .C2(n6803), .ZN(n6902) );
  AOI211_X1 U8505 ( .C1(n8379), .C2(n6805), .A(n6907), .B(n6902), .ZN(n6806)
         );
  OAI21_X1 U8506 ( .B1(n9678), .B2(n6910), .A(n6806), .ZN(n6823) );
  NAND2_X1 U8507 ( .A1(n6823), .A2(n9736), .ZN(n6807) );
  OAI21_X1 U8508 ( .B1(n9736), .B2(n6808), .A(n6807), .ZN(P2_U3466) );
  INV_X1 U8509 ( .A(n6809), .ZN(n6811) );
  INV_X1 U8510 ( .A(n8882), .ZN(n7297) );
  OAI222_X1 U8511 ( .A1(n9340), .A2(n6810), .B1(n9343), .B2(n6811), .C1(n7297), 
        .C2(P1_U3084), .ZN(P1_U3337) );
  INV_X1 U8512 ( .A(n7996), .ZN(n7121) );
  OAI222_X1 U8513 ( .A1(n8417), .A2(n6812), .B1(n8414), .B2(n6811), .C1(n7121), 
        .C2(n4264), .ZN(P2_U3342) );
  INV_X1 U8514 ( .A(n6814), .ZN(n6815) );
  AOI21_X1 U8515 ( .B1(n4267), .B2(n6813), .A(n6815), .ZN(n7179) );
  AOI22_X1 U8516 ( .A1(n9603), .A2(n8849), .B1(n8848), .B2(n9600), .ZN(n6817)
         );
  AOI21_X1 U8517 ( .B1(n7099), .B2(n7186), .A(n9158), .ZN(n6816) );
  NAND2_X1 U8518 ( .A1(n6816), .A2(n7511), .ZN(n7184) );
  OAI211_X1 U8519 ( .C1(n7179), .C2(n9273), .A(n6817), .B(n7184), .ZN(n6819)
         );
  XOR2_X1 U8520 ( .A(n4267), .B(n8804), .Z(n6818) );
  NOR2_X1 U8521 ( .A1(n6818), .A2(n9399), .ZN(n7178) );
  NOR2_X1 U8522 ( .A1(n6819), .A2(n7178), .ZN(n6837) );
  INV_X1 U8523 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n6820) );
  OAI22_X1 U8524 ( .A1(n9280), .A2(n8809), .B1(n4270), .B2(n6820), .ZN(n6821)
         );
  INV_X1 U8525 ( .A(n6821), .ZN(n6822) );
  OAI21_X1 U8526 ( .B1(n6837), .B2(n9625), .A(n6822), .ZN(P1_U3525) );
  INV_X1 U8527 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n6825) );
  NAND2_X1 U8528 ( .A1(n6823), .A2(n9752), .ZN(n6824) );
  OAI21_X1 U8529 ( .B1(n9752), .B2(n6825), .A(n6824), .ZN(P2_U3525) );
  INV_X1 U8530 ( .A(n6826), .ZN(n6838) );
  AOI22_X1 U8531 ( .A1(n8897), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n9332), .ZN(n6827) );
  OAI21_X1 U8532 ( .B1(n6838), .B2(n9343), .A(n6827), .ZN(P1_U3336) );
  OAI211_X1 U8533 ( .C1(n6830), .C2(n6829), .A(n6828), .B(n7631), .ZN(n6834)
         );
  INV_X1 U8534 ( .A(n7050), .ZN(n9694) );
  OAI22_X1 U8535 ( .A1(n7660), .A2(n9694), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n5899), .ZN(n6832) );
  INV_X1 U8536 ( .A(n7912), .ZN(n7044) );
  OAI22_X1 U8537 ( .A1(n7017), .A2(n7666), .B1(n7645), .B2(n7044), .ZN(n6831)
         );
  AOI211_X1 U8538 ( .C1(n7012), .C2(n7657), .A(n6832), .B(n6831), .ZN(n6833)
         );
  NAND2_X1 U8539 ( .A1(n6834), .A2(n6833), .ZN(P2_U3215) );
  OAI22_X1 U8540 ( .A1(n9326), .A2(n8809), .B1(n9619), .B2(n4940), .ZN(n6835)
         );
  INV_X1 U8541 ( .A(n6835), .ZN(n6836) );
  OAI21_X1 U8542 ( .B1(n6837), .B2(n9617), .A(n6836), .ZN(P1_U3460) );
  INV_X1 U8543 ( .A(n8013), .ZN(n7995) );
  OAI222_X1 U8544 ( .A1(n8417), .A2(n6839), .B1(n8414), .B2(n6838), .C1(n7995), 
        .C2(P2_U3152), .ZN(P2_U3341) );
  INV_X1 U8545 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n9391) );
  AOI22_X1 U8546 ( .A1(n6989), .A2(P2_REG1_REG_14__SCAN_IN), .B1(n9391), .B2(
        n6848), .ZN(n6842) );
  OAI21_X1 U8547 ( .B1(n6845), .B2(P2_REG1_REG_13__SCAN_IN), .A(n6840), .ZN(
        n6841) );
  NAND2_X1 U8548 ( .A1(n6842), .A2(n6841), .ZN(n6991) );
  OAI21_X1 U8549 ( .B1(n6842), .B2(n6841), .A(n6991), .ZN(n6855) );
  NAND2_X1 U8550 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3152), .ZN(n7549) );
  INV_X1 U8551 ( .A(n7549), .ZN(n6843) );
  AOI21_X1 U8552 ( .B1(n9633), .B2(P2_ADDR_REG_14__SCAN_IN), .A(n6843), .ZN(
        n6844) );
  OAI21_X1 U8553 ( .B1(n9628), .B2(n6848), .A(n6844), .ZN(n6854) );
  NOR2_X1 U8554 ( .A1(n6845), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n6847) );
  NOR2_X1 U8555 ( .A1(n6847), .A2(n6846), .ZN(n6851) );
  INV_X1 U8556 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n6849) );
  AOI22_X1 U8557 ( .A1(n6989), .A2(n6849), .B1(P2_REG2_REG_14__SCAN_IN), .B2(
        n6848), .ZN(n6850) );
  NOR2_X1 U8558 ( .A1(n6851), .A2(n6850), .ZN(n6986) );
  AOI21_X1 U8559 ( .B1(n6851), .B2(n6850), .A(n6986), .ZN(n6852) );
  NOR2_X1 U8560 ( .A1(n6852), .A2(n8029), .ZN(n6853) );
  AOI211_X1 U8561 ( .C1(n6855), .C2(n9627), .A(n6854), .B(n6853), .ZN(n6856)
         );
  INV_X1 U8562 ( .A(n6856), .ZN(P2_U3259) );
  NAND2_X1 U8563 ( .A1(n6858), .A2(n6857), .ZN(n6859) );
  XOR2_X1 U8564 ( .A(n6860), .B(n6859), .Z(n6864) );
  NAND2_X1 U8565 ( .A1(n9452), .A2(n7103), .ZN(n9580) );
  NOR2_X1 U8566 ( .A1(n6867), .A2(n9580), .ZN(n6861) );
  AOI21_X1 U8567 ( .B1(P1_REG3_REG_1__SCAN_IN), .B2(n6867), .A(n6861), .ZN(
        n6863) );
  AOI22_X1 U8568 ( .A1(n8534), .A2(n5653), .B1(n8548), .B2(n5655), .ZN(n6862)
         );
  OAI211_X1 U8569 ( .C1(n6864), .C2(n8554), .A(n6863), .B(n6862), .ZN(P1_U3220) );
  XOR2_X1 U8570 ( .A(n6866), .B(n6865), .Z(n6870) );
  AOI22_X1 U8571 ( .A1(n8552), .A2(n7186), .B1(n6867), .B2(
        P1_REG3_REG_2__SCAN_IN), .ZN(n6869) );
  AOI22_X1 U8572 ( .A1(n8534), .A2(n8849), .B1(n8548), .B2(n8848), .ZN(n6868)
         );
  OAI211_X1 U8573 ( .C1(n6870), .C2(n8554), .A(n6869), .B(n6868), .ZN(P1_U3235) );
  OAI211_X1 U8574 ( .C1(n6873), .C2(n6872), .A(n6871), .B(n7631), .ZN(n6877)
         );
  INV_X1 U8575 ( .A(n9654), .ZN(n7067) );
  NAND2_X1 U8576 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(n4264), .ZN(n7951) );
  OAI21_X1 U8577 ( .B1(n7645), .B2(n7067), .A(n7951), .ZN(n6875) );
  INV_X1 U8578 ( .A(n7056), .ZN(n9700) );
  OAI22_X1 U8579 ( .A1(n7666), .A2(n7051), .B1(n9700), .B2(n7660), .ZN(n6874)
         );
  AOI211_X1 U8580 ( .C1(n9664), .C2(n7657), .A(n6875), .B(n6874), .ZN(n6876)
         );
  NAND2_X1 U8581 ( .A1(n6877), .A2(n6876), .ZN(P2_U3223) );
  OAI21_X1 U8582 ( .B1(n6879), .B2(n6882), .A(n6878), .ZN(n7201) );
  NAND2_X1 U8583 ( .A1(n7201), .A2(n9615), .ZN(n6887) );
  AOI22_X1 U8584 ( .A1(n9603), .A2(n8848), .B1(n9602), .B2(n9600), .ZN(n6886)
         );
  NAND2_X1 U8585 ( .A1(n6881), .A2(n6880), .ZN(n7217) );
  XNOR2_X1 U8586 ( .A(n7217), .B(n6882), .ZN(n6883) );
  NAND2_X1 U8587 ( .A1(n6883), .A2(n9550), .ZN(n7203) );
  INV_X1 U8588 ( .A(n7215), .ZN(n6885) );
  AOI21_X1 U8589 ( .B1(n7513), .B2(n7196), .A(n9158), .ZN(n6884) );
  NAND2_X1 U8590 ( .A1(n6885), .A2(n6884), .ZN(n7199) );
  NAND4_X1 U8591 ( .A1(n6887), .A2(n6886), .A3(n7203), .A4(n7199), .ZN(n6893)
         );
  OAI22_X1 U8592 ( .A1(n9280), .A2(n6891), .B1(n4270), .B2(n6416), .ZN(n6888)
         );
  AOI21_X1 U8593 ( .B1(n6893), .B2(n4270), .A(n6888), .ZN(n6889) );
  INV_X1 U8594 ( .A(n6889), .ZN(P1_U3527) );
  INV_X1 U8595 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n6890) );
  OAI22_X1 U8596 ( .A1(n9326), .A2(n6891), .B1(n9619), .B2(n6890), .ZN(n6892)
         );
  AOI21_X1 U8597 ( .B1(n6893), .B2(n9619), .A(n6892), .ZN(n6894) );
  INV_X1 U8598 ( .A(n6894), .ZN(P1_U3466) );
  NOR2_X1 U8599 ( .A1(n7727), .A2(n6896), .ZN(n9679) );
  NAND2_X1 U8600 ( .A1(n9649), .A2(n8290), .ZN(n6978) );
  INV_X1 U8601 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n9631) );
  OAI22_X1 U8602 ( .A1(n9679), .A2(n9660), .B1(n6897), .B2(n8284), .ZN(n9681)
         );
  AOI22_X1 U8603 ( .A1(n9661), .A2(n9681), .B1(P2_REG3_REG_0__SCAN_IN), .B2(
        n9665), .ZN(n6898) );
  OAI21_X1 U8604 ( .B1(n9631), .B2(n9661), .A(n6898), .ZN(n6899) );
  AOI21_X1 U8605 ( .B1(n6900), .B2(n6978), .A(n6899), .ZN(n6901) );
  OAI21_X1 U8606 ( .B1(n6895), .B2(n9679), .A(n6901), .ZN(P2_U3296) );
  INV_X1 U8607 ( .A(n6902), .ZN(n6903) );
  MUX2_X1 U8608 ( .A(n6429), .B(n6903), .S(n9661), .Z(n6909) );
  INV_X1 U8609 ( .A(n6904), .ZN(n6905) );
  OAI22_X1 U8610 ( .A1(n9649), .A2(n6979), .B1(n8142), .B2(n6905), .ZN(n6906)
         );
  AOI21_X1 U8611 ( .B1(n8257), .B2(n6907), .A(n6906), .ZN(n6908) );
  OAI211_X1 U8612 ( .C1(n6895), .C2(n6910), .A(n6909), .B(n6908), .ZN(P2_U3291) );
  OAI21_X1 U8613 ( .B1(n6912), .B2(n6922), .A(n6911), .ZN(n9687) );
  INV_X1 U8614 ( .A(n9687), .ZN(n6929) );
  INV_X1 U8615 ( .A(n9649), .ZN(n7000) );
  OAI22_X1 U8616 ( .A1(n6914), .A2(n9661), .B1(n6913), .B2(n8142), .ZN(n6918)
         );
  OAI21_X1 U8617 ( .B1(n9683), .B2(n6916), .A(n6915), .ZN(n9684) );
  NOR2_X1 U8618 ( .A1(n8290), .A2(n9684), .ZN(n6917) );
  AOI211_X1 U8619 ( .C1(n7000), .C2(n6919), .A(n6918), .B(n6917), .ZN(n6928)
         );
  NAND2_X1 U8620 ( .A1(n6921), .A2(n6920), .ZN(n6923) );
  INV_X1 U8621 ( .A(n6922), .ZN(n7871) );
  XNOR2_X1 U8622 ( .A(n6923), .B(n7871), .ZN(n6924) );
  NAND2_X1 U8623 ( .A1(n6924), .A2(n8213), .ZN(n6926) );
  AOI22_X1 U8624 ( .A1(n9656), .A2(n7916), .B1(n7914), .B2(n9653), .ZN(n6925)
         );
  NAND2_X1 U8625 ( .A1(n6926), .A2(n6925), .ZN(n9685) );
  NAND2_X1 U8626 ( .A1(n9685), .A2(n9661), .ZN(n6927) );
  OAI211_X1 U8627 ( .C1(n6895), .C2(n6929), .A(n6928), .B(n6927), .ZN(P2_U3292) );
  XOR2_X1 U8628 ( .A(n6930), .B(n6932), .Z(n6938) );
  INV_X1 U8629 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n6936) );
  INV_X1 U8630 ( .A(n8550), .ZN(n8499) );
  AOI22_X1 U8631 ( .A1(n8534), .A2(n5655), .B1(n8548), .B2(n8847), .ZN(n6934)
         );
  AND2_X1 U8632 ( .A1(P1_U3084), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n8851) );
  INV_X1 U8633 ( .A(n8851), .ZN(n6933) );
  OAI211_X1 U8634 ( .C1(n9590), .C2(n7464), .A(n6934), .B(n6933), .ZN(n6935)
         );
  AOI21_X1 U8635 ( .B1(n6936), .B2(n8499), .A(n6935), .ZN(n6937) );
  OAI21_X1 U8636 ( .B1(n6938), .B2(n8554), .A(n6937), .ZN(P1_U3216) );
  XOR2_X1 U8637 ( .A(n6940), .B(n6939), .Z(n6941) );
  XNOR2_X1 U8638 ( .A(n6942), .B(n6941), .ZN(n6946) );
  AOI22_X1 U8639 ( .A1(n8534), .A2(n8848), .B1(n8548), .B2(n9602), .ZN(n6944)
         );
  AND2_X1 U8640 ( .A1(P1_U3084), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n9494) );
  AOI21_X1 U8641 ( .B1(n8552), .B2(n7196), .A(n9494), .ZN(n6943) );
  OAI211_X1 U8642 ( .C1(n8550), .C2(n7194), .A(n6944), .B(n6943), .ZN(n6945)
         );
  AOI21_X1 U8643 ( .B1(n6946), .B2(n8475), .A(n6945), .ZN(n6947) );
  INV_X1 U8644 ( .A(n6947), .ZN(P1_U3228) );
  INV_X1 U8645 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n6949) );
  INV_X1 U8646 ( .A(n6948), .ZN(n6950) );
  INV_X1 U8647 ( .A(n8024), .ZN(n8020) );
  OAI222_X1 U8648 ( .A1(n8417), .A2(n6949), .B1(n8414), .B2(n6950), .C1(n4264), 
        .C2(n8020), .ZN(P2_U3340) );
  INV_X1 U8649 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n6951) );
  INV_X1 U8650 ( .A(n8898), .ZN(n9534) );
  OAI222_X1 U8651 ( .A1(n9340), .A2(n6951), .B1(n9343), .B2(n6950), .C1(
        P1_U3084), .C2(n9534), .ZN(P1_U3335) );
  AOI21_X1 U8652 ( .B1(n6953), .B2(n6952), .A(n4347), .ZN(n6957) );
  INV_X1 U8653 ( .A(n7911), .ZN(n7173) );
  AOI22_X1 U8654 ( .A1(n7643), .A2(n7912), .B1(n7657), .B2(n7058), .ZN(n6954)
         );
  NAND2_X1 U8655 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(n4264), .ZN(n7964) );
  OAI211_X1 U8656 ( .C1(n7645), .C2(n7173), .A(n6954), .B(n7964), .ZN(n6955)
         );
  AOI21_X1 U8657 ( .B1(n7670), .B2(n7071), .A(n6955), .ZN(n6956) );
  OAI21_X1 U8658 ( .B1(n6957), .B2(n7673), .A(n6956), .ZN(P2_U3233) );
  NAND2_X1 U8659 ( .A1(n6958), .A2(n7895), .ZN(n6961) );
  OAI22_X1 U8660 ( .A1(n6961), .A2(n6960), .B1(n6959), .B2(n8142), .ZN(n6964)
         );
  NOR2_X1 U8661 ( .A1(n8278), .A2(n6962), .ZN(n6963) );
  AOI211_X1 U8662 ( .C1(n8278), .C2(P2_REG2_REG_2__SCAN_IN), .A(n6964), .B(
        n6963), .ZN(n6967) );
  INV_X1 U8663 ( .A(n6895), .ZN(n8164) );
  NAND2_X1 U8664 ( .A1(n8164), .A2(n6965), .ZN(n6966) );
  OAI211_X1 U8665 ( .C1(n6968), .C2(n9649), .A(n6967), .B(n6966), .ZN(P2_U3294) );
  OR2_X1 U8666 ( .A1(n7913), .A2(n7008), .ZN(n7743) );
  NAND2_X1 U8667 ( .A1(n7008), .A2(n7913), .ZN(n7734) );
  NAND2_X1 U8668 ( .A1(n7743), .A2(n7734), .ZN(n7873) );
  INV_X1 U8669 ( .A(n7873), .ZN(n6971) );
  OAI21_X1 U8670 ( .B1(n6971), .B2(n6970), .A(n7015), .ZN(n6972) );
  AOI222_X1 U8671 ( .A1(n8213), .A2(n6972), .B1(n9655), .B2(n9653), .C1(n7914), 
        .C2(n9656), .ZN(n9689) );
  NAND2_X1 U8672 ( .A1(n6973), .A2(n7008), .ZN(n7010) );
  OAI211_X1 U8673 ( .C1(n7008), .C2(n6973), .A(n7010), .B(n8380), .ZN(n6974)
         );
  OAI21_X1 U8674 ( .B1(n7008), .B2(n9727), .A(n6974), .ZN(n9691) );
  INV_X1 U8675 ( .A(n6975), .ZN(n6976) );
  OAI22_X1 U8676 ( .A1(n9661), .A2(n6428), .B1(n6976), .B2(n8142), .ZN(n6977)
         );
  AOI21_X1 U8677 ( .B1(n9691), .B2(n6978), .A(n6977), .ZN(n6984) );
  NAND2_X1 U8678 ( .A1(n6980), .A2(n6979), .ZN(n6981) );
  XNOR2_X1 U8679 ( .A(n7009), .B(n7873), .ZN(n9692) );
  NAND2_X1 U8680 ( .A1(n8164), .A2(n9692), .ZN(n6983) );
  OAI211_X1 U8681 ( .C1(n9689), .C2(n8278), .A(n6984), .B(n6983), .ZN(P2_U3290) );
  NOR2_X1 U8682 ( .A1(n6989), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n6985) );
  NAND2_X1 U8683 ( .A1(n6987), .A2(n6994), .ZN(n7112) );
  OAI21_X1 U8684 ( .B1(n6987), .B2(n6994), .A(n7112), .ZN(n6988) );
  NOR2_X1 U8685 ( .A1(n6988), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n7114) );
  AOI21_X1 U8686 ( .B1(P2_REG2_REG_15__SCAN_IN), .B2(n6988), .A(n7114), .ZN(
        n6998) );
  INV_X1 U8687 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n9385) );
  OR2_X1 U8688 ( .A1(n6989), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n6990) );
  NAND2_X1 U8689 ( .A1(n6991), .A2(n6990), .ZN(n7106) );
  XOR2_X1 U8690 ( .A(n7108), .B(n7106), .Z(n6992) );
  NOR2_X1 U8691 ( .A1(n6992), .A2(n9385), .ZN(n7107) );
  AOI211_X1 U8692 ( .C1(n9385), .C2(n6992), .A(n9629), .B(n7107), .ZN(n6993)
         );
  INV_X1 U8693 ( .A(n6993), .ZN(n6997) );
  AND2_X1 U8694 ( .A1(P2_U3152), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n7668) );
  NOR2_X1 U8695 ( .A1(n9628), .A2(n6994), .ZN(n6995) );
  AOI211_X1 U8696 ( .C1(P2_ADDR_REG_15__SCAN_IN), .C2(n9633), .A(n7668), .B(
        n6995), .ZN(n6996) );
  OAI211_X1 U8697 ( .C1(n6998), .C2(n8029), .A(n6997), .B(n6996), .ZN(P2_U3260) );
  MUX2_X1 U8698 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n6999), .S(n9661), .Z(n7005)
         );
  AOI22_X1 U8699 ( .A1(n9647), .A2(n7001), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        n9665), .ZN(n7002) );
  OAI21_X1 U8700 ( .B1(n7003), .B2(n8293), .A(n7002), .ZN(n7004) );
  AOI211_X1 U8701 ( .C1(n8164), .C2(n7006), .A(n7005), .B(n7004), .ZN(n7007)
         );
  INV_X1 U8702 ( .A(n7007), .ZN(P2_U3295) );
  XNOR2_X1 U8703 ( .A(n7051), .B(n7050), .ZN(n7741) );
  XNOR2_X1 U8704 ( .A(n7041), .B(n7741), .ZN(n9698) );
  INV_X1 U8705 ( .A(n7010), .ZN(n7011) );
  OR2_X1 U8706 ( .A1(n7010), .A2(n7050), .ZN(n9642) );
  OAI21_X1 U8707 ( .B1(n7011), .B2(n9694), .A(n9642), .ZN(n9695) );
  INV_X1 U8708 ( .A(n9695), .ZN(n7013) );
  AOI22_X1 U8709 ( .A1(n7013), .A2(n9647), .B1(n7012), .B2(n9665), .ZN(n7014)
         );
  OAI21_X1 U8710 ( .B1(n9694), .B2(n8293), .A(n7014), .ZN(n7019) );
  XNOR2_X1 U8711 ( .A(n7052), .B(n7741), .ZN(n7016) );
  OAI222_X1 U8712 ( .A1(n8284), .A2(n7044), .B1(n8285), .B2(n7017), .C1(n9660), 
        .C2(n7016), .ZN(n9696) );
  MUX2_X1 U8713 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n9696), .S(n9661), .Z(n7018)
         );
  AOI211_X1 U8714 ( .C1(n9698), .C2(n8164), .A(n7019), .B(n7018), .ZN(n7020)
         );
  INV_X1 U8715 ( .A(n7020), .ZN(P2_U3289) );
  INV_X1 U8716 ( .A(n7021), .ZN(n7023) );
  OAI222_X1 U8717 ( .A1(n8417), .A2(n7022), .B1(n8414), .B2(n7023), .C1(n7895), 
        .C2(n4264), .ZN(P2_U3339) );
  OAI222_X1 U8718 ( .A1(n9340), .A2(n7024), .B1(n9343), .B2(n7023), .C1(
        P1_U3084), .C2(n9123), .ZN(P1_U3334) );
  OAI21_X1 U8719 ( .B1(n7026), .B2(n7027), .A(n7025), .ZN(n7204) );
  NAND3_X1 U8720 ( .A1(n7028), .A2(n8813), .A3(n7027), .ZN(n7029) );
  AND2_X1 U8721 ( .A1(n7030), .A2(n7029), .ZN(n7214) );
  AOI22_X1 U8722 ( .A1(n9603), .A2(n8846), .B1(n9547), .B2(n9600), .ZN(n7033)
         );
  INV_X1 U8723 ( .A(n7238), .ZN(n7032) );
  INV_X1 U8724 ( .A(n7031), .ZN(n7351) );
  OAI211_X1 U8725 ( .C1(n7209), .C2(n7032), .A(n7351), .B(n9559), .ZN(n7205)
         );
  OAI211_X1 U8726 ( .C1(n7214), .C2(n9399), .A(n7033), .B(n7205), .ZN(n7034)
         );
  AOI21_X1 U8727 ( .B1(n7204), .B2(n9615), .A(n7034), .ZN(n7040) );
  OAI22_X1 U8728 ( .A1(n9326), .A2(n7209), .B1(n9619), .B2(n5075), .ZN(n7035)
         );
  INV_X1 U8729 ( .A(n7035), .ZN(n7036) );
  OAI21_X1 U8730 ( .B1(n7040), .B2(n9617), .A(n7036), .ZN(P1_U3475) );
  INV_X1 U8731 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n7037) );
  OAI22_X1 U8732 ( .A1(n9280), .A2(n7209), .B1(n4270), .B2(n7037), .ZN(n7038)
         );
  INV_X1 U8733 ( .A(n7038), .ZN(n7039) );
  OAI21_X1 U8734 ( .B1(n7040), .B2(n9625), .A(n7039), .ZN(P1_U3530) );
  NAND2_X1 U8735 ( .A1(n7041), .A2(n7741), .ZN(n7043) );
  OR2_X1 U8736 ( .A1(n9655), .A2(n7050), .ZN(n7042) );
  NAND2_X1 U8737 ( .A1(n7043), .A2(n7042), .ZN(n9641) );
  INV_X1 U8738 ( .A(n9641), .ZN(n7045) );
  OR2_X1 U8739 ( .A1(n7056), .A2(n7044), .ZN(n7749) );
  NAND2_X1 U8740 ( .A1(n7056), .A2(n7044), .ZN(n7750) );
  NAND2_X1 U8741 ( .A1(n7749), .A2(n7750), .ZN(n7874) );
  NAND2_X1 U8742 ( .A1(n7056), .A2(n7912), .ZN(n7046) );
  OR2_X1 U8743 ( .A1(n7071), .A2(n7067), .ZN(n7758) );
  NAND2_X1 U8744 ( .A1(n7071), .A2(n7067), .ZN(n7753) );
  NAND2_X1 U8745 ( .A1(n7048), .A2(n7877), .ZN(n7049) );
  NAND2_X1 U8746 ( .A1(n7073), .A2(n7049), .ZN(n9709) );
  AND2_X1 U8747 ( .A1(n7051), .A2(n7050), .ZN(n7744) );
  NAND2_X1 U8748 ( .A1(n9694), .A2(n9655), .ZN(n7746) );
  XNOR2_X1 U8749 ( .A(n7074), .B(n7047), .ZN(n7054) );
  AOI22_X1 U8750 ( .A1(n9656), .A2(n7912), .B1(n7911), .B2(n9653), .ZN(n7053)
         );
  OAI21_X1 U8751 ( .B1(n7054), .B2(n9660), .A(n7053), .ZN(n7055) );
  AOI21_X1 U8752 ( .B1(n9709), .B2(n9652), .A(n7055), .ZN(n9711) );
  INV_X1 U8753 ( .A(n7071), .ZN(n9706) );
  AND2_X1 U8754 ( .A1(n9643), .A2(n9706), .ZN(n7080) );
  NOR2_X1 U8755 ( .A1(n9643), .A2(n9706), .ZN(n7057) );
  OR2_X1 U8756 ( .A1(n7080), .A2(n7057), .ZN(n9707) );
  NOR2_X1 U8757 ( .A1(n9707), .A2(n8290), .ZN(n7061) );
  AOI22_X1 U8758 ( .A1(n8278), .A2(P2_REG2_REG_9__SCAN_IN), .B1(n7058), .B2(
        n9665), .ZN(n7059) );
  OAI21_X1 U8759 ( .B1(n9706), .B2(n8293), .A(n7059), .ZN(n7060) );
  AOI211_X1 U8760 ( .C1(n9709), .C2(n9648), .A(n7061), .B(n7060), .ZN(n7062)
         );
  OAI21_X1 U8761 ( .B1(n9711), .B2(n8278), .A(n7062), .ZN(P2_U3287) );
  INV_X1 U8762 ( .A(n7164), .ZN(n9712) );
  OAI211_X1 U8763 ( .C1(n7065), .C2(n7064), .A(n7063), .B(n7631), .ZN(n7070)
         );
  AND2_X1 U8764 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(n4264), .ZN(n7978) );
  INV_X1 U8765 ( .A(n7082), .ZN(n7066) );
  OAI22_X1 U8766 ( .A1(n7666), .A2(n7067), .B1(n7665), .B2(n7066), .ZN(n7068)
         );
  AOI211_X1 U8767 ( .C1(n7669), .C2(n7910), .A(n7978), .B(n7068), .ZN(n7069)
         );
  OAI211_X1 U8768 ( .C1(n9712), .C2(n7660), .A(n7070), .B(n7069), .ZN(P2_U3219) );
  OR2_X1 U8769 ( .A1(n7071), .A2(n9654), .ZN(n7072) );
  OR2_X1 U8770 ( .A1(n7164), .A2(n7173), .ZN(n7757) );
  NAND2_X1 U8771 ( .A1(n7164), .A2(n7173), .ZN(n7756) );
  XNOR2_X1 U8772 ( .A(n7166), .B(n4672), .ZN(n9716) );
  NOR2_X1 U8773 ( .A1(n7075), .A2(n7878), .ZN(n7076) );
  OAI21_X1 U8774 ( .B1(n7169), .B2(n7076), .A(n8213), .ZN(n7078) );
  AOI22_X1 U8775 ( .A1(n9653), .A2(n7910), .B1(n9654), .B2(n9656), .ZN(n7077)
         );
  NAND2_X1 U8776 ( .A1(n7078), .A2(n7077), .ZN(n7079) );
  AOI21_X1 U8777 ( .B1(n9716), .B2(n9652), .A(n7079), .ZN(n9718) );
  NAND2_X1 U8778 ( .A1(n7080), .A2(n9712), .ZN(n7319) );
  OR2_X1 U8779 ( .A1(n7080), .A2(n9712), .ZN(n7081) );
  NAND2_X1 U8780 ( .A1(n7319), .A2(n7081), .ZN(n9713) );
  NOR2_X1 U8781 ( .A1(n9713), .A2(n8290), .ZN(n7085) );
  AOI22_X1 U8782 ( .A1(n8278), .A2(P2_REG2_REG_10__SCAN_IN), .B1(n7082), .B2(
        n9665), .ZN(n7083) );
  OAI21_X1 U8783 ( .B1(n9712), .B2(n8293), .A(n7083), .ZN(n7084) );
  AOI211_X1 U8784 ( .C1(n9716), .C2(n9648), .A(n7085), .B(n7084), .ZN(n7086)
         );
  OAI21_X1 U8785 ( .B1(n9718), .B2(n8278), .A(n7086), .ZN(P2_U3286) );
  OR2_X1 U8786 ( .A1(n7088), .A2(n7087), .ZN(n7180) );
  OR3_X2 U8787 ( .A1(n7089), .A2(n9570), .A3(n8556), .ZN(n9567) );
  OAI21_X4 U8788 ( .B1(n7180), .B2(n9328), .A(n9567), .ZN(n9572) );
  NOR2_X1 U8789 ( .A1(n7091), .A2(n7090), .ZN(n7092) );
  OAI21_X1 U8790 ( .B1(n5713), .B2(n7094), .A(n7093), .ZN(n9583) );
  INV_X1 U8791 ( .A(n5655), .ZN(n7098) );
  INV_X1 U8792 ( .A(n5653), .ZN(n7097) );
  XNOR2_X1 U8793 ( .A(n5713), .B(n7095), .ZN(n7096) );
  OAI222_X1 U8794 ( .A1(n9440), .A2(n7098), .B1(n9438), .B2(n7097), .C1(n7096), 
        .C2(n9399), .ZN(n9584) );
  OAI211_X1 U8795 ( .C1(n8802), .C2(n7100), .A(n9559), .B(n7099), .ZN(n9581)
         );
  OAI22_X1 U8796 ( .A1(n9581), .A2(n9074), .B1(n9567), .B2(n7101), .ZN(n7102)
         );
  OAI21_X1 U8797 ( .B1(n9584), .B2(n7102), .A(n9572), .ZN(n7105) );
  AOI22_X1 U8798 ( .A1(n9554), .A2(n7103), .B1(n9575), .B2(
        P1_REG2_REG_1__SCAN_IN), .ZN(n7104) );
  OAI211_X1 U8799 ( .C1(n9079), .C2(n9583), .A(n7105), .B(n7104), .ZN(P1_U3290) );
  INV_X1 U8800 ( .A(n7106), .ZN(n7109) );
  AOI21_X1 U8801 ( .B1(n7109), .B2(n7108), .A(n7107), .ZN(n7111) );
  XOR2_X1 U8802 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n7996), .Z(n7110) );
  NAND2_X1 U8803 ( .A1(n7110), .A2(n7111), .ZN(n7997) );
  OAI21_X1 U8804 ( .B1(n7111), .B2(n7110), .A(n7997), .ZN(n7123) );
  INV_X1 U8805 ( .A(n7112), .ZN(n7113) );
  NOR2_X1 U8806 ( .A1(n7114), .A2(n7113), .ZN(n7117) );
  INV_X1 U8807 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n9894) );
  NAND2_X1 U8808 ( .A1(n7996), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n7989) );
  INV_X1 U8809 ( .A(n7989), .ZN(n7115) );
  AOI21_X1 U8810 ( .B1(n9894), .B2(n7121), .A(n7115), .ZN(n7116) );
  NAND2_X1 U8811 ( .A1(n7116), .A2(n7117), .ZN(n7988) );
  OAI211_X1 U8812 ( .C1(n7117), .C2(n7116), .A(n9632), .B(n7988), .ZN(n7120)
         );
  NAND2_X1 U8813 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(n4264), .ZN(n7590) );
  INV_X1 U8814 ( .A(n7590), .ZN(n7118) );
  AOI21_X1 U8815 ( .B1(n9633), .B2(P2_ADDR_REG_16__SCAN_IN), .A(n7118), .ZN(
        n7119) );
  OAI211_X1 U8816 ( .C1(n9628), .C2(n7121), .A(n7120), .B(n7119), .ZN(n7122)
         );
  AOI21_X1 U8817 ( .B1(n7123), .B2(n9627), .A(n7122), .ZN(n7124) );
  INV_X1 U8818 ( .A(n7124), .ZN(P2_U3261) );
  NAND2_X1 U8819 ( .A1(n7126), .A2(n7125), .ZN(n7128) );
  XOR2_X1 U8820 ( .A(n7128), .B(n7127), .Z(n7133) );
  AOI22_X1 U8821 ( .A1(n8534), .A2(n9602), .B1(n8548), .B2(n9601), .ZN(n7131)
         );
  AOI21_X1 U8822 ( .B1(n8552), .B2(n4269), .A(n7129), .ZN(n7130) );
  OAI211_X1 U8823 ( .C1(n8550), .C2(n7240), .A(n7131), .B(n7130), .ZN(n7132)
         );
  AOI21_X1 U8824 ( .B1(n7133), .B2(n8475), .A(n7132), .ZN(n7134) );
  INV_X1 U8825 ( .A(n7134), .ZN(P1_U3237) );
  INV_X1 U8826 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n7149) );
  AOI21_X1 U8827 ( .B1(n7141), .B2(P1_REG2_REG_13__SCAN_IN), .A(n7135), .ZN(
        n7137) );
  INV_X1 U8828 ( .A(n9513), .ZN(n7136) );
  NAND2_X1 U8829 ( .A1(n7137), .A2(n7136), .ZN(n7138) );
  INV_X1 U8830 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n9518) );
  NAND2_X1 U8831 ( .A1(n7138), .A2(n9517), .ZN(n7283) );
  XNOR2_X1 U8832 ( .A(n7290), .B(n7283), .ZN(n7139) );
  NOR2_X1 U8833 ( .A1(n9153), .A2(n7139), .ZN(n7284) );
  AOI211_X1 U8834 ( .C1(n7139), .C2(n9153), .A(n7284), .B(n9503), .ZN(n7147)
         );
  XNOR2_X1 U8835 ( .A(n9513), .B(P1_REG1_REG_14__SCAN_IN), .ZN(n9516) );
  OAI21_X1 U8836 ( .B1(P1_REG1_REG_13__SCAN_IN), .B2(n7141), .A(n7140), .ZN(
        n7142) );
  INV_X1 U8837 ( .A(n7142), .ZN(n9515) );
  OAI22_X1 U8838 ( .A1(n9516), .A2(n9515), .B1(n9513), .B2(
        P1_REG1_REG_14__SCAN_IN), .ZN(n7289) );
  XNOR2_X1 U8839 ( .A(n7289), .B(n7290), .ZN(n7143) );
  NOR2_X1 U8840 ( .A1(n7144), .A2(n7143), .ZN(n7291) );
  AOI211_X1 U8841 ( .C1(n7144), .C2(n7143), .A(n7291), .B(n9490), .ZN(n7146)
         );
  NAND2_X1 U8842 ( .A1(P1_U3084), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n8544) );
  OAI21_X1 U8843 ( .B1(n9533), .B2(n7290), .A(n8544), .ZN(n7145) );
  NOR3_X1 U8844 ( .A1(n7147), .A2(n7146), .A3(n7145), .ZN(n7148) );
  OAI21_X1 U8845 ( .B1(n9525), .B2(n7149), .A(n7148), .ZN(P1_U3256) );
  INV_X1 U8846 ( .A(n7150), .ZN(n7162) );
  OAI222_X1 U8847 ( .A1(n9340), .A2(n7152), .B1(n9343), .B2(n7162), .C1(n7151), 
        .C2(P1_U3084), .ZN(P1_U3333) );
  XOR2_X1 U8848 ( .A(n7153), .B(n7154), .Z(n7161) );
  INV_X1 U8849 ( .A(n9547), .ZN(n7382) );
  NOR2_X1 U8850 ( .A1(n7411), .A2(n7382), .ZN(n7155) );
  AOI211_X1 U8851 ( .C1(n8534), .C2(n8846), .A(n7156), .B(n7155), .ZN(n7160)
         );
  INV_X1 U8852 ( .A(n7157), .ZN(n7206) );
  AOI22_X1 U8853 ( .A1(n8499), .A2(n7206), .B1(n8552), .B2(n7158), .ZN(n7159)
         );
  OAI211_X1 U8854 ( .C1(n7161), .C2(n8554), .A(n7160), .B(n7159), .ZN(P1_U3211) );
  OAI222_X1 U8855 ( .A1(n8417), .A2(n7163), .B1(n4264), .B2(n7865), .C1(n8414), 
        .C2(n7162), .ZN(P2_U3338) );
  NAND2_X1 U8856 ( .A1(n7164), .A2(n7911), .ZN(n7165) );
  INV_X1 U8857 ( .A(n7910), .ZN(n7318) );
  OR2_X1 U8858 ( .A1(n7636), .A2(n7318), .ZN(n7766) );
  NAND2_X1 U8859 ( .A1(n7636), .A2(n7318), .ZN(n7769) );
  OAI21_X1 U8860 ( .B1(n7167), .B2(n7881), .A(n7313), .ZN(n9720) );
  INV_X1 U8861 ( .A(n7909), .ZN(n7314) );
  INV_X1 U8862 ( .A(n7756), .ZN(n7759) );
  INV_X1 U8863 ( .A(n7316), .ZN(n7171) );
  NOR3_X1 U8864 ( .A1(n7169), .A2(n7759), .A3(n7168), .ZN(n7170) );
  NOR2_X1 U8865 ( .A1(n7171), .A2(n7170), .ZN(n7172) );
  OAI222_X1 U8866 ( .A1(n8285), .A2(n7173), .B1(n8284), .B2(n7314), .C1(n9660), 
        .C2(n7172), .ZN(n9723) );
  XNOR2_X1 U8867 ( .A(n7319), .B(n7636), .ZN(n9722) );
  NOR2_X1 U8868 ( .A1(n9722), .A2(n8290), .ZN(n7176) );
  INV_X1 U8869 ( .A(n7636), .ZN(n9721) );
  AOI22_X1 U8870 ( .A1(n8278), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n7635), .B2(
        n9665), .ZN(n7174) );
  OAI21_X1 U8871 ( .B1(n9721), .B2(n8293), .A(n7174), .ZN(n7175) );
  AOI211_X1 U8872 ( .C1(n9723), .C2(n9661), .A(n7176), .B(n7175), .ZN(n7177)
         );
  OAI21_X1 U8873 ( .B1(n6895), .B2(n9720), .A(n7177), .ZN(P2_U3285) );
  INV_X1 U8874 ( .A(n7178), .ZN(n7193) );
  INV_X1 U8875 ( .A(n7179), .ZN(n7191) );
  AND2_X1 U8876 ( .A1(n9572), .A2(n9603), .ZN(n9136) );
  INV_X1 U8877 ( .A(n9136), .ZN(n9157) );
  INV_X1 U8878 ( .A(n7180), .ZN(n7183) );
  AND2_X1 U8879 ( .A1(n7181), .A2(n9123), .ZN(n7182) );
  OAI22_X1 U8880 ( .A1(n7184), .A2(n9162), .B1(n9469), .B2(n9567), .ZN(n7185)
         );
  AOI21_X1 U8881 ( .B1(P1_REG2_REG_2__SCAN_IN), .B2(n9575), .A(n7185), .ZN(
        n7188) );
  AND2_X1 U8882 ( .A1(n9572), .A2(n9600), .ZN(n9155) );
  AOI22_X1 U8883 ( .A1(n9554), .A2(n7186), .B1(n9155), .B2(n8848), .ZN(n7187)
         );
  OAI211_X1 U8884 ( .C1(n7189), .C2(n9157), .A(n7188), .B(n7187), .ZN(n7190)
         );
  AOI21_X1 U8885 ( .B1(n7191), .B2(n9563), .A(n7190), .ZN(n7192) );
  OAI21_X1 U8886 ( .B1(n9575), .B2(n7193), .A(n7192), .ZN(P1_U3289) );
  OAI22_X1 U8887 ( .A1(n9572), .A2(n6391), .B1(n7194), .B2(n9567), .ZN(n7195)
         );
  AOI21_X1 U8888 ( .B1(n9554), .B2(n7196), .A(n7195), .ZN(n7198) );
  AOI22_X1 U8889 ( .A1(n9136), .A2(n8848), .B1(n9155), .B2(n9602), .ZN(n7197)
         );
  OAI211_X1 U8890 ( .C1(n7199), .C2(n9162), .A(n7198), .B(n7197), .ZN(n7200)
         );
  AOI21_X1 U8891 ( .B1(n7201), .B2(n9563), .A(n7200), .ZN(n7202) );
  OAI21_X1 U8892 ( .B1(n9575), .B2(n7203), .A(n7202), .ZN(P1_U3287) );
  AND2_X1 U8893 ( .A1(n9572), .A2(n9550), .ZN(n8953) );
  INV_X1 U8894 ( .A(n8953), .ZN(n9146) );
  NAND2_X1 U8895 ( .A1(n7204), .A2(n9563), .ZN(n7213) );
  INV_X1 U8896 ( .A(n7205), .ZN(n7211) );
  AOI22_X1 U8897 ( .A1(n9136), .A2(n8846), .B1(n9155), .B2(n9547), .ZN(n7208)
         );
  INV_X1 U8898 ( .A(n9567), .ZN(n9552) );
  AOI22_X1 U8899 ( .A1(n9575), .A2(P1_REG2_REG_7__SCAN_IN), .B1(n7206), .B2(
        n9552), .ZN(n7207) );
  OAI211_X1 U8900 ( .C1(n7209), .C2(n9060), .A(n7208), .B(n7207), .ZN(n7210)
         );
  AOI21_X1 U8901 ( .B1(n7211), .B2(n9562), .A(n7210), .ZN(n7212) );
  OAI211_X1 U8902 ( .C1(n7214), .C2(n9146), .A(n7213), .B(n7212), .ZN(P1_U3284) );
  OAI211_X1 U8903 ( .C1(n7215), .C2(n9596), .A(n7237), .B(n9559), .ZN(n9595)
         );
  NOR2_X1 U8904 ( .A1(n9595), .A2(n9074), .ZN(n7222) );
  INV_X1 U8905 ( .A(n8688), .ZN(n7216) );
  OR2_X1 U8906 ( .A1(n7217), .A2(n7216), .ZN(n7218) );
  NAND2_X1 U8907 ( .A1(n7218), .A2(n8687), .ZN(n8571) );
  XNOR2_X1 U8908 ( .A(n8571), .B(n7230), .ZN(n7219) );
  NAND2_X1 U8909 ( .A1(n7219), .A2(n9550), .ZN(n7221) );
  AOI22_X1 U8910 ( .A1(n9603), .A2(n8847), .B1(n8846), .B2(n9600), .ZN(n7220)
         );
  NAND2_X1 U8911 ( .A1(n7221), .A2(n7220), .ZN(n9598) );
  AOI211_X1 U8912 ( .C1(n9552), .C2(n8478), .A(n7222), .B(n9598), .ZN(n7223)
         );
  MUX2_X1 U8913 ( .A(n7224), .B(n7223), .S(n9572), .Z(n7229) );
  INV_X1 U8914 ( .A(n7225), .ZN(n7226) );
  AOI21_X1 U8915 ( .B1(n7230), .B2(n7227), .A(n7226), .ZN(n9599) );
  AOI22_X1 U8916 ( .A1(n9599), .A2(n9563), .B1(n9554), .B2(n8477), .ZN(n7228)
         );
  NAND2_X1 U8917 ( .A1(n7229), .A2(n7228), .ZN(P1_U3286) );
  NAND2_X1 U8918 ( .A1(n8571), .A2(n7230), .ZN(n7231) );
  NAND2_X1 U8919 ( .A1(n7231), .A2(n8691), .ZN(n7232) );
  INV_X1 U8920 ( .A(n8569), .ZN(n7235) );
  XNOR2_X1 U8921 ( .A(n7232), .B(n7235), .ZN(n7233) );
  NOR2_X1 U8922 ( .A1(n7233), .A2(n9399), .ZN(n9606) );
  INV_X1 U8923 ( .A(n9606), .ZN(n7247) );
  OAI21_X1 U8924 ( .B1(n7236), .B2(n7235), .A(n7234), .ZN(n9608) );
  AOI21_X1 U8925 ( .B1(n7237), .B2(n4269), .A(n9158), .ZN(n7239) );
  NAND2_X1 U8926 ( .A1(n7239), .A2(n7238), .ZN(n9605) );
  OAI22_X1 U8927 ( .A1(n9572), .A2(n5041), .B1(n7240), .B2(n9567), .ZN(n7241)
         );
  AOI21_X1 U8928 ( .B1(n9554), .B2(n4269), .A(n7241), .ZN(n7244) );
  AOI22_X1 U8929 ( .A1(n9136), .A2(n9602), .B1(n9155), .B2(n9601), .ZN(n7243)
         );
  OAI211_X1 U8930 ( .C1(n9605), .C2(n9162), .A(n7244), .B(n7243), .ZN(n7245)
         );
  AOI21_X1 U8931 ( .B1(n9608), .B2(n9563), .A(n7245), .ZN(n7246) );
  OAI21_X1 U8932 ( .B1(n9575), .B2(n7247), .A(n7246), .ZN(P1_U3285) );
  INV_X1 U8933 ( .A(n7248), .ZN(n7250) );
  OAI222_X1 U8934 ( .A1(n9340), .A2(n7249), .B1(n9343), .B2(n7250), .C1(n8801), 
        .C2(P1_U3084), .ZN(P1_U3332) );
  OAI222_X1 U8935 ( .A1(n8417), .A2(n7251), .B1(P2_U3152), .B2(n4266), .C1(
        n8414), .C2(n7250), .ZN(P2_U3337) );
  INV_X1 U8936 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n9936) );
  NOR2_X1 U8937 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n7252) );
  AOI21_X1 U8938 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n7252), .ZN(n9759) );
  NOR2_X1 U8939 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n7253) );
  AOI21_X1 U8940 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n7253), .ZN(n9762) );
  NOR2_X1 U8941 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n7254) );
  AOI21_X1 U8942 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n7254), .ZN(n9765) );
  NOR2_X1 U8943 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n7255) );
  AOI21_X1 U8944 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n7255), .ZN(n9768) );
  NOR2_X1 U8945 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n7256) );
  AOI21_X1 U8946 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n7256), .ZN(n9771) );
  NOR2_X1 U8947 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n7262) );
  XNOR2_X1 U8948 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n9947) );
  NAND2_X1 U8949 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n7260) );
  XOR2_X1 U8950 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(P2_ADDR_REG_3__SCAN_IN), .Z(
        n9945) );
  NAND2_X1 U8951 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n7258) );
  XOR2_X1 U8952 ( .A(P2_ADDR_REG_2__SCAN_IN), .B(P1_ADDR_REG_2__SCAN_IN), .Z(
        n9943) );
  AOI21_X1 U8953 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n9753) );
  INV_X1 U8954 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n9823) );
  NAND3_X1 U8955 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_1__SCAN_IN), .ZN(n9755) );
  OAI21_X1 U8956 ( .B1(n9753), .B2(n9823), .A(n9755), .ZN(n9942) );
  NAND2_X1 U8957 ( .A1(n9943), .A2(n9942), .ZN(n7257) );
  NAND2_X1 U8958 ( .A1(n7258), .A2(n7257), .ZN(n9944) );
  NAND2_X1 U8959 ( .A1(n9945), .A2(n9944), .ZN(n7259) );
  NAND2_X1 U8960 ( .A1(n7260), .A2(n7259), .ZN(n9946) );
  NOR2_X1 U8961 ( .A1(n9947), .A2(n9946), .ZN(n7261) );
  NOR2_X1 U8962 ( .A1(n7262), .A2(n7261), .ZN(n7263) );
  NOR2_X1 U8963 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n7263), .ZN(n9931) );
  AND2_X1 U8964 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n7263), .ZN(n9930) );
  NOR2_X1 U8965 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n9930), .ZN(n7264) );
  NOR2_X1 U8966 ( .A1(n9931), .A2(n7264), .ZN(n7265) );
  NAND2_X1 U8967 ( .A1(n7265), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n7267) );
  XOR2_X1 U8968 ( .A(n7265), .B(P1_ADDR_REG_6__SCAN_IN), .Z(n9929) );
  NAND2_X1 U8969 ( .A1(n9929), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n7266) );
  NAND2_X1 U8970 ( .A1(n7267), .A2(n7266), .ZN(n7268) );
  NAND2_X1 U8971 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n7268), .ZN(n7270) );
  XOR2_X1 U8972 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n7268), .Z(n9938) );
  NAND2_X1 U8973 ( .A1(n9938), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n7269) );
  NAND2_X1 U8974 ( .A1(n7270), .A2(n7269), .ZN(n7271) );
  NAND2_X1 U8975 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n7271), .ZN(n7273) );
  XOR2_X1 U8976 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(n7271), .Z(n9933) );
  NAND2_X1 U8977 ( .A1(n9933), .A2(P2_ADDR_REG_8__SCAN_IN), .ZN(n7272) );
  NAND2_X1 U8978 ( .A1(n7273), .A2(n7272), .ZN(n7274) );
  AND2_X1 U8979 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n7274), .ZN(n7275) );
  INV_X1 U8980 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n9941) );
  XNOR2_X1 U8981 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n7274), .ZN(n9940) );
  NOR2_X1 U8982 ( .A1(n9941), .A2(n9940), .ZN(n9939) );
  NAND2_X1 U8983 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n7276) );
  OAI21_X1 U8984 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n7276), .ZN(n9779) );
  NAND2_X1 U8985 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n7277) );
  OAI21_X1 U8986 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n7277), .ZN(n9776) );
  NOR2_X1 U8987 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n7278) );
  AOI21_X1 U8988 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n7278), .ZN(n9773) );
  NAND2_X1 U8989 ( .A1(n9774), .A2(n9773), .ZN(n9772) );
  NAND2_X1 U8990 ( .A1(n9771), .A2(n9770), .ZN(n9769) );
  NAND2_X1 U8991 ( .A1(n9768), .A2(n9767), .ZN(n9766) );
  OAI21_X1 U8992 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n9766), .ZN(n9764) );
  NAND2_X1 U8993 ( .A1(n9765), .A2(n9764), .ZN(n9763) );
  OAI21_X1 U8994 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n9763), .ZN(n9761) );
  NAND2_X1 U8995 ( .A1(n9762), .A2(n9761), .ZN(n9760) );
  OAI21_X1 U8996 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n9760), .ZN(n9758) );
  NAND2_X1 U8997 ( .A1(n9759), .A2(n9758), .ZN(n9757) );
  OAI21_X1 U8998 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n9757), .ZN(n9935) );
  NOR2_X1 U8999 ( .A1(n9936), .A2(n9935), .ZN(n7279) );
  NAND2_X1 U9000 ( .A1(n9936), .A2(n9935), .ZN(n9934) );
  OAI21_X1 U9001 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n7279), .A(n9934), .ZN(
        n7282) );
  XNOR2_X1 U9002 ( .A(n7280), .B(P1_ADDR_REG_19__SCAN_IN), .ZN(n7281) );
  XNOR2_X1 U9003 ( .A(n7282), .B(n7281), .ZN(ADD_1071_U4) );
  NOR2_X1 U9004 ( .A1(n7290), .A2(n7283), .ZN(n7285) );
  NAND2_X1 U9005 ( .A1(P1_REG2_REG_16__SCAN_IN), .A2(n8882), .ZN(n7286) );
  OAI21_X1 U9006 ( .B1(n8882), .B2(P1_REG2_REG_16__SCAN_IN), .A(n7286), .ZN(
        n7287) );
  NOR2_X1 U9007 ( .A1(n7288), .A2(n7287), .ZN(n8878) );
  AOI211_X1 U9008 ( .C1(n7288), .C2(n7287), .A(n8878), .B(n9503), .ZN(n7300)
         );
  NOR2_X1 U9009 ( .A1(n7290), .A2(n7289), .ZN(n7292) );
  NOR2_X1 U9010 ( .A1(n7292), .A2(n7291), .ZN(n7294) );
  XNOR2_X1 U9011 ( .A(n8882), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n7293) );
  NOR2_X1 U9012 ( .A1(n7294), .A2(n7293), .ZN(n8881) );
  AOI211_X1 U9013 ( .C1(n7294), .C2(n7293), .A(n8881), .B(n9490), .ZN(n7299)
         );
  NAND2_X1 U9014 ( .A1(n9539), .A2(P1_ADDR_REG_16__SCAN_IN), .ZN(n7296) );
  NAND2_X1 U9015 ( .A1(P1_REG3_REG_16__SCAN_IN), .A2(P1_U3084), .ZN(n7295) );
  OAI211_X1 U9016 ( .C1(n9533), .C2(n7297), .A(n7296), .B(n7295), .ZN(n7298)
         );
  OR3_X1 U9017 ( .A1(n7300), .A2(n7299), .A3(n7298), .ZN(P1_U3257) );
  NAND2_X1 U9018 ( .A1(n7302), .A2(n7301), .ZN(n7304) );
  XOR2_X1 U9019 ( .A(n7304), .B(n7303), .Z(n7309) );
  AOI22_X1 U9020 ( .A1(n7643), .A2(n7910), .B1(n7657), .B2(n7320), .ZN(n7306)
         );
  OAI211_X1 U9021 ( .C1(n7645), .C2(n7434), .A(n7306), .B(n7305), .ZN(n7307)
         );
  AOI21_X1 U9022 ( .B1(n7670), .B2(n7387), .A(n7307), .ZN(n7308) );
  OAI21_X1 U9023 ( .B1(n7309), .B2(n7673), .A(n7308), .ZN(P2_U3226) );
  INV_X1 U9024 ( .A(n7310), .ZN(n7532) );
  OAI222_X1 U9025 ( .A1(n9340), .A2(n7311), .B1(n9343), .B2(n7532), .C1(
        P1_U3084), .C2(n4265), .ZN(P1_U3331) );
  NAND2_X1 U9026 ( .A1(n7636), .A2(n7910), .ZN(n7312) );
  OR2_X1 U9027 ( .A1(n7387), .A2(n7314), .ZN(n7771) );
  NAND2_X1 U9028 ( .A1(n7387), .A2(n7314), .ZN(n7770) );
  NAND2_X1 U9029 ( .A1(n7771), .A2(n7770), .ZN(n7882) );
  INV_X1 U9030 ( .A(n7882), .ZN(n7315) );
  OAI21_X1 U9031 ( .B1(n4344), .B2(n7882), .A(n4836), .ZN(n9732) );
  INV_X1 U9032 ( .A(n9732), .ZN(n7325) );
  XNOR2_X1 U9033 ( .A(n7388), .B(n7882), .ZN(n7317) );
  OAI222_X1 U9034 ( .A1(n8284), .A2(n7434), .B1(n8285), .B2(n7318), .C1(n7317), 
        .C2(n9660), .ZN(n9730) );
  OAI21_X1 U9035 ( .B1(n4465), .B2(n4464), .A(n7393), .ZN(n9729) );
  NOR2_X1 U9036 ( .A1(n9729), .A2(n8290), .ZN(n7323) );
  AOI22_X1 U9037 ( .A1(n8278), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n7320), .B2(
        n9665), .ZN(n7321) );
  OAI21_X1 U9038 ( .B1(n4464), .B2(n8293), .A(n7321), .ZN(n7322) );
  AOI211_X1 U9039 ( .C1(n9730), .C2(n9661), .A(n7323), .B(n7322), .ZN(n7324)
         );
  OAI21_X1 U9040 ( .B1(n6895), .B2(n7325), .A(n7324), .ZN(P2_U3284) );
  NAND2_X1 U9041 ( .A1(n7326), .A2(n7327), .ZN(n7329) );
  XNOR2_X1 U9042 ( .A(n7329), .B(n7328), .ZN(n7337) );
  INV_X1 U9043 ( .A(n9601), .ZN(n7332) );
  NAND2_X1 U9044 ( .A1(n8548), .A2(n8845), .ZN(n7331) );
  OAI211_X1 U9045 ( .C1(n7332), .C2(n8545), .A(n7331), .B(n7330), .ZN(n7334)
         );
  NOR2_X1 U9046 ( .A1(n8550), .A2(n7353), .ZN(n7333) );
  NOR2_X1 U9047 ( .A1(n7334), .A2(n7333), .ZN(n7336) );
  NAND2_X1 U9048 ( .A1(n8552), .A2(n7352), .ZN(n7335) );
  OAI211_X1 U9049 ( .C1(n7337), .C2(n8554), .A(n7336), .B(n7335), .ZN(P1_U3219) );
  XNOR2_X1 U9050 ( .A(n7338), .B(n7339), .ZN(n7344) );
  AOI22_X1 U9051 ( .A1(n9656), .A2(n7909), .B1(n7907), .B2(n9653), .ZN(n7390)
         );
  NAND2_X1 U9052 ( .A1(n7657), .A2(n7394), .ZN(n7341) );
  OAI211_X1 U9053 ( .C1(n7390), .C2(n7655), .A(n7341), .B(n7340), .ZN(n7342)
         );
  AOI21_X1 U9054 ( .B1(n7670), .B2(n8378), .A(n7342), .ZN(n7343) );
  OAI21_X1 U9055 ( .B1(n7344), .B2(n7673), .A(n7343), .ZN(P2_U3236) );
  INV_X1 U9056 ( .A(n9544), .ZN(n7345) );
  NOR2_X1 U9057 ( .A1(n9545), .A2(n7345), .ZN(n7346) );
  AOI211_X1 U9058 ( .C1(n8700), .C2(n7347), .A(n9399), .B(n7346), .ZN(n7350)
         );
  OAI21_X1 U9059 ( .B1(n4342), .B2(n8700), .A(n7348), .ZN(n7419) );
  NOR2_X1 U9060 ( .A1(n7419), .A2(n9419), .ZN(n7349) );
  AOI211_X1 U9061 ( .C1(n9603), .C2(n9601), .A(n7350), .B(n7349), .ZN(n7418)
         );
  AOI211_X1 U9062 ( .C1(n7352), .C2(n7351), .A(n9158), .B(n9560), .ZN(n7416)
         );
  OAI22_X1 U9063 ( .A1(n9572), .A2(n6395), .B1(n7353), .B2(n9567), .ZN(n7354)
         );
  AOI21_X1 U9064 ( .B1(n9155), .B2(n8845), .A(n7354), .ZN(n7355) );
  OAI21_X1 U9065 ( .B1(n7423), .B2(n9060), .A(n7355), .ZN(n7357) );
  NOR2_X1 U9066 ( .A1(n7419), .A2(n9079), .ZN(n7356) );
  AOI211_X1 U9067 ( .C1(n7416), .C2(n9562), .A(n7357), .B(n7356), .ZN(n7358)
         );
  OAI21_X1 U9068 ( .B1(n7418), .B2(n9575), .A(n7358), .ZN(P1_U3283) );
  XNOR2_X1 U9069 ( .A(n7359), .B(n8704), .ZN(n7360) );
  NAND2_X1 U9070 ( .A1(n7360), .A2(n9550), .ZN(n9374) );
  XNOR2_X1 U9071 ( .A(n7361), .B(n8704), .ZN(n9376) );
  INV_X1 U9072 ( .A(n9376), .ZN(n9378) );
  NAND2_X1 U9073 ( .A1(n9378), .A2(n9563), .ZN(n7369) );
  INV_X1 U9074 ( .A(n9425), .ZN(n7362) );
  AOI211_X1 U9075 ( .C1(n9373), .C2(n9558), .A(n9158), .B(n7362), .ZN(n9371)
         );
  INV_X1 U9076 ( .A(n8845), .ZN(n9370) );
  OAI22_X1 U9077 ( .A1(n9572), .A2(n7363), .B1(n7408), .B2(n9567), .ZN(n7364)
         );
  AOI21_X1 U9078 ( .B1(n9155), .B2(n8844), .A(n7364), .ZN(n7366) );
  NAND2_X1 U9079 ( .A1(n9554), .A2(n9373), .ZN(n7365) );
  OAI211_X1 U9080 ( .C1(n9370), .C2(n9157), .A(n7366), .B(n7365), .ZN(n7367)
         );
  AOI21_X1 U9081 ( .B1(n9371), .B2(n9562), .A(n7367), .ZN(n7368) );
  OAI211_X1 U9082 ( .C1(n9575), .C2(n9374), .A(n7369), .B(n7368), .ZN(P1_U3281) );
  INV_X1 U9083 ( .A(n7373), .ZN(n7371) );
  NAND2_X1 U9084 ( .A1(n8410), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n7370) );
  OAI211_X1 U9085 ( .C1(n7371), .C2(n8414), .A(n7904), .B(n7370), .ZN(P2_U3335) );
  NAND2_X1 U9086 ( .A1(n7373), .A2(n7372), .ZN(n7375) );
  OR2_X1 U9087 ( .A1(n7374), .A2(P1_U3084), .ZN(n8829) );
  OAI211_X1 U9088 ( .C1(n7376), .C2(n9340), .A(n7375), .B(n8829), .ZN(P1_U3330) );
  XNOR2_X1 U9089 ( .A(n7377), .B(n7378), .ZN(n7379) );
  NAND2_X1 U9090 ( .A1(n7379), .A2(n8475), .ZN(n7386) );
  NAND2_X1 U9091 ( .A1(n8548), .A2(n9548), .ZN(n7381) );
  AND2_X1 U9092 ( .A1(P1_U3084), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n9508) );
  INV_X1 U9093 ( .A(n9508), .ZN(n7380) );
  OAI211_X1 U9094 ( .C1(n7382), .C2(n8545), .A(n7381), .B(n7380), .ZN(n7384)
         );
  NOR2_X1 U9095 ( .A1(n8550), .A2(n9551), .ZN(n7383) );
  NOR2_X1 U9096 ( .A1(n7384), .A2(n7383), .ZN(n7385) );
  OAI211_X1 U9097 ( .C1(n9613), .C2(n7464), .A(n7386), .B(n7385), .ZN(P1_U3229) );
  OR2_X1 U9098 ( .A1(n8378), .A2(n7434), .ZN(n7777) );
  NAND2_X1 U9099 ( .A1(n8378), .A2(n7434), .ZN(n7776) );
  NAND2_X1 U9100 ( .A1(n7777), .A2(n7776), .ZN(n7883) );
  XNOR2_X1 U9101 ( .A(n7427), .B(n7883), .ZN(n8377) );
  AOI21_X1 U9102 ( .B1(n7883), .B2(n7389), .A(n7432), .ZN(n7391) );
  OAI21_X1 U9103 ( .B1(n7391), .B2(n9660), .A(n7390), .ZN(n7392) );
  AOI21_X1 U9104 ( .B1(n9652), .B2(n8377), .A(n7392), .ZN(n8383) );
  INV_X1 U9105 ( .A(n8378), .ZN(n7397) );
  AOI21_X1 U9106 ( .B1(n8378), .B2(n7393), .A(n8036), .ZN(n8381) );
  NAND2_X1 U9107 ( .A1(n8381), .A2(n9647), .ZN(n7396) );
  AOI22_X1 U9108 ( .A1(n8278), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n7394), .B2(
        n9665), .ZN(n7395) );
  OAI211_X1 U9109 ( .C1(n7397), .C2(n9649), .A(n7396), .B(n7395), .ZN(n7398)
         );
  AOI21_X1 U9110 ( .B1(n8377), .B2(n9648), .A(n7398), .ZN(n7399) );
  OAI21_X1 U9111 ( .B1(n8383), .B2(n8278), .A(n7399), .ZN(P2_U3283) );
  INV_X1 U9112 ( .A(n7400), .ZN(n7404) );
  OAI222_X1 U9113 ( .A1(P1_U3084), .A2(n7402), .B1(n9343), .B2(n7404), .C1(
        n7401), .C2(n9340), .ZN(P1_U3329) );
  OAI222_X1 U9114 ( .A1(P2_U3152), .A2(n7405), .B1(n8414), .B2(n7404), .C1(
        n7403), .C2(n8417), .ZN(P2_U3334) );
  XOR2_X1 U9115 ( .A(n7406), .B(n7407), .Z(n7415) );
  NOR2_X1 U9116 ( .A1(n8550), .A2(n7408), .ZN(n7413) );
  NAND2_X1 U9117 ( .A1(n8534), .A2(n8845), .ZN(n7410) );
  OAI211_X1 U9118 ( .C1(n7411), .C2(n9439), .A(n7410), .B(n7409), .ZN(n7412)
         );
  AOI211_X1 U9119 ( .C1(n8552), .C2(n9373), .A(n7413), .B(n7412), .ZN(n7414)
         );
  OAI21_X1 U9120 ( .B1(n7415), .B2(n8554), .A(n7414), .ZN(P1_U3215) );
  AOI21_X1 U9121 ( .B1(n9600), .B2(n8845), .A(n7416), .ZN(n7417) );
  OAI211_X1 U9122 ( .C1(n9582), .C2(n7419), .A(n7418), .B(n7417), .ZN(n7425)
         );
  OAI22_X1 U9123 ( .A1(n9280), .A2(n7423), .B1(n4270), .B2(n6407), .ZN(n7420)
         );
  AOI21_X1 U9124 ( .B1(n7425), .B2(n4270), .A(n7420), .ZN(n7421) );
  INV_X1 U9125 ( .A(n7421), .ZN(P1_U3531) );
  INV_X1 U9126 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n7422) );
  OAI22_X1 U9127 ( .A1(n9326), .A2(n7423), .B1(n9619), .B2(n7422), .ZN(n7424)
         );
  AOI21_X1 U9128 ( .B1(n7425), .B2(n9619), .A(n7424), .ZN(n7426) );
  INV_X1 U9129 ( .A(n7426), .ZN(P1_U3478) );
  AOI21_X1 U9130 ( .B1(n7428), .B2(n7883), .A(n4842), .ZN(n7431) );
  NAND2_X1 U9131 ( .A1(n7780), .A2(n7907), .ZN(n7429) );
  NAND2_X1 U9132 ( .A1(n8048), .A2(n7429), .ZN(n7884) );
  INV_X1 U9133 ( .A(n7884), .ZN(n7430) );
  OAI21_X1 U9134 ( .B1(n7431), .B2(n7430), .A(n8049), .ZN(n9390) );
  INV_X1 U9135 ( .A(n9390), .ZN(n7439) );
  XNOR2_X1 U9136 ( .A(n7682), .B(n7884), .ZN(n7433) );
  OAI222_X1 U9137 ( .A1(n8285), .A2(n7434), .B1(n8284), .B2(n7683), .C1(n9660), 
        .C2(n7433), .ZN(n9388) );
  XNOR2_X1 U9138 ( .A(n8036), .B(n9386), .ZN(n9387) );
  NOR2_X1 U9139 ( .A1(n9387), .A2(n8290), .ZN(n7437) );
  AOI22_X1 U9140 ( .A1(n8278), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n7548), .B2(
        n9665), .ZN(n7435) );
  OAI21_X1 U9141 ( .B1(n9386), .B2(n8293), .A(n7435), .ZN(n7436) );
  AOI211_X1 U9142 ( .C1(n9388), .C2(n9661), .A(n7437), .B(n7436), .ZN(n7438)
         );
  OAI21_X1 U9143 ( .B1(n6895), .B2(n7439), .A(n7438), .ZN(P2_U3282) );
  AOI21_X1 U9144 ( .B1(n7440), .B2(n8706), .A(n9399), .ZN(n7442) );
  NAND2_X1 U9145 ( .A1(n7442), .A2(n7441), .ZN(n9445) );
  OAI21_X1 U9146 ( .B1(n7444), .B2(n8706), .A(n7443), .ZN(n9447) );
  INV_X1 U9147 ( .A(n9447), .ZN(n9449) );
  NAND2_X1 U9148 ( .A1(n9449), .A2(n9563), .ZN(n7453) );
  INV_X1 U9149 ( .A(n9428), .ZN(n7445) );
  AOI211_X1 U9150 ( .C1(n9444), .C2(n7445), .A(n9158), .B(n9408), .ZN(n9442)
         );
  INV_X1 U9151 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n7446) );
  OAI22_X1 U9152 ( .A1(n9572), .A2(n7446), .B1(n7488), .B2(n9567), .ZN(n7447)
         );
  AOI21_X1 U9153 ( .B1(n9155), .B2(n8842), .A(n7447), .ZN(n7449) );
  NAND2_X1 U9154 ( .A1(n9136), .A2(n8844), .ZN(n7448) );
  OAI211_X1 U9155 ( .C1(n7450), .C2(n9060), .A(n7449), .B(n7448), .ZN(n7451)
         );
  AOI21_X1 U9156 ( .B1(n9442), .B2(n9562), .A(n7451), .ZN(n7452) );
  OAI211_X1 U9157 ( .C1(n9575), .C2(n9445), .A(n7453), .B(n7452), .ZN(P1_U3279) );
  INV_X1 U9158 ( .A(n9451), .ZN(n7465) );
  AOI21_X1 U9159 ( .B1(n7454), .B2(n7455), .A(n8554), .ZN(n7457) );
  NAND2_X1 U9160 ( .A1(n7457), .A2(n7456), .ZN(n7463) );
  NAND2_X1 U9161 ( .A1(n8548), .A2(n8843), .ZN(n7459) );
  OAI211_X1 U9162 ( .C1(n9414), .C2(n8545), .A(n7459), .B(n7458), .ZN(n7461)
         );
  NOR2_X1 U9163 ( .A1(n8550), .A2(n9423), .ZN(n7460) );
  NOR2_X1 U9164 ( .A1(n7461), .A2(n7460), .ZN(n7462) );
  OAI211_X1 U9165 ( .C1(n7465), .C2(n7464), .A(n7463), .B(n7462), .ZN(P1_U3234) );
  XNOR2_X1 U9166 ( .A(n7466), .B(n8709), .ZN(n9277) );
  INV_X1 U9167 ( .A(n9277), .ZN(n7476) );
  OAI211_X1 U9168 ( .C1(n7468), .C2(n8709), .A(n7467), .B(n9550), .ZN(n7470)
         );
  AOI22_X1 U9169 ( .A1(n9603), .A2(n8842), .B1(n9255), .B2(n9600), .ZN(n7469)
         );
  NAND2_X1 U9170 ( .A1(n7470), .A2(n7469), .ZN(n9275) );
  INV_X1 U9171 ( .A(n8430), .ZN(n9327) );
  AOI211_X1 U9172 ( .C1(n8430), .C2(n4289), .A(n9158), .B(n4532), .ZN(n9276)
         );
  NAND2_X1 U9173 ( .A1(n9276), .A2(n9562), .ZN(n7473) );
  INV_X1 U9174 ( .A(n8428), .ZN(n7471) );
  AOI22_X1 U9175 ( .A1(n9575), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n7471), .B2(
        n9552), .ZN(n7472) );
  OAI211_X1 U9176 ( .C1(n9327), .C2(n9060), .A(n7473), .B(n7472), .ZN(n7474)
         );
  AOI21_X1 U9177 ( .B1(n9572), .B2(n9275), .A(n7474), .ZN(n7475) );
  OAI21_X1 U9178 ( .B1(n7476), .B2(n9079), .A(n7475), .ZN(P1_U3277) );
  INV_X1 U9179 ( .A(n7477), .ZN(n7481) );
  OAI222_X1 U9180 ( .A1(n9340), .A2(n7479), .B1(n9343), .B2(n7481), .C1(
        P1_U3084), .C2(n7478), .ZN(P1_U3328) );
  OAI222_X1 U9181 ( .A1(n8417), .A2(n9829), .B1(n8414), .B2(n7481), .C1(
        P2_U3152), .C2(n7480), .ZN(P2_U3333) );
  INV_X1 U9182 ( .A(n7482), .ZN(n7483) );
  AOI21_X1 U9183 ( .B1(n7485), .B2(n7484), .A(n7483), .ZN(n7491) );
  AOI22_X1 U9184 ( .A1(n8534), .A2(n8844), .B1(P1_REG3_REG_12__SCAN_IN), .B2(
        P1_U3084), .ZN(n7487) );
  NAND2_X1 U9185 ( .A1(n8548), .A2(n8842), .ZN(n7486) );
  OAI211_X1 U9186 ( .C1(n8550), .C2(n7488), .A(n7487), .B(n7486), .ZN(n7489)
         );
  AOI21_X1 U9187 ( .B1(n8552), .B2(n9444), .A(n7489), .ZN(n7490) );
  OAI21_X1 U9188 ( .B1(n7491), .B2(n8554), .A(n7490), .ZN(P1_U3222) );
  XNOR2_X1 U9189 ( .A(n7494), .B(n7493), .ZN(n7495) );
  XNOR2_X1 U9190 ( .A(n7492), .B(n7495), .ZN(n7502) );
  INV_X1 U9191 ( .A(n7496), .ZN(n7498) );
  NOR2_X1 U9192 ( .A1(n8545), .A2(n9413), .ZN(n7497) );
  AOI211_X1 U9193 ( .C1(n8548), .C2(n9266), .A(n7498), .B(n7497), .ZN(n7499)
         );
  OAI21_X1 U9194 ( .B1(n8550), .B2(n9405), .A(n7499), .ZN(n7500) );
  AOI21_X1 U9195 ( .B1(n8552), .B2(n9407), .A(n7500), .ZN(n7501) );
  OAI21_X1 U9196 ( .B1(n7502), .B2(n8554), .A(n7501), .ZN(P1_U3232) );
  XNOR2_X1 U9197 ( .A(n8747), .B(n7503), .ZN(n7509) );
  OR2_X1 U9198 ( .A1(n7504), .A2(n7503), .ZN(n7505) );
  NAND2_X1 U9199 ( .A1(n7506), .A2(n7505), .ZN(n9593) );
  NAND2_X1 U9200 ( .A1(n9593), .A2(n9587), .ZN(n7508) );
  AOI22_X1 U9201 ( .A1(n9603), .A2(n5655), .B1(n8847), .B2(n9600), .ZN(n7507)
         );
  OAI211_X1 U9202 ( .C1(n9399), .C2(n7509), .A(n7508), .B(n7507), .ZN(n9591)
         );
  MUX2_X1 U9203 ( .A(n9591), .B(P1_REG2_REG_3__SCAN_IN), .S(n9575), .Z(n7518)
         );
  NAND2_X1 U9204 ( .A1(n9593), .A2(n9563), .ZN(n7516) );
  AOI21_X1 U9205 ( .B1(n7511), .B2(n7510), .A(n9158), .ZN(n7512) );
  AND2_X1 U9206 ( .A1(n7513), .A2(n7512), .ZN(n9588) );
  NOR2_X1 U9207 ( .A1(n9567), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n7514) );
  AOI21_X1 U9208 ( .B1(n9588), .B2(n9562), .A(n7514), .ZN(n7515) );
  OAI211_X1 U9209 ( .C1(n9590), .C2(n9060), .A(n7516), .B(n7515), .ZN(n7517)
         );
  OR2_X1 U9210 ( .A1(n7518), .A2(n7517), .ZN(P1_U3288) );
  INV_X1 U9211 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n8560) );
  INV_X1 U9212 ( .A(n7519), .ZN(n7520) );
  NOR2_X1 U9213 ( .A1(n7520), .A2(SI_29_), .ZN(n7522) );
  NAND2_X1 U9214 ( .A1(n7520), .A2(SI_29_), .ZN(n7521) );
  MUX2_X1 U9215 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n7698), .Z(n7695) );
  INV_X1 U9216 ( .A(n8559), .ZN(n7526) );
  OAI222_X1 U9217 ( .A1(n9340), .A2(n8560), .B1(n9343), .B2(n7526), .C1(n7524), 
        .C2(P1_U3084), .ZN(P1_U3323) );
  INV_X1 U9218 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n9863) );
  OAI222_X1 U9219 ( .A1(n8417), .A2(n9863), .B1(n8414), .B2(n7526), .C1(n7525), 
        .C2(P2_U3152), .ZN(P2_U3328) );
  INV_X1 U9220 ( .A(n7527), .ZN(n9335) );
  OAI222_X1 U9221 ( .A1(n8417), .A2(n7529), .B1(n4264), .B2(n7528), .C1(n8414), 
        .C2(n9335), .ZN(P2_U3330) );
  INV_X1 U9222 ( .A(n7688), .ZN(n7534) );
  OAI222_X1 U9223 ( .A1(n8414), .A2(n7534), .B1(P2_U3152), .B2(n7531), .C1(
        n7530), .C2(n8417), .ZN(P2_U3329) );
  OAI222_X1 U9224 ( .A1(n8417), .A2(n7533), .B1(n8414), .B2(n7532), .C1(n6505), 
        .C2(n4264), .ZN(P2_U3336) );
  OAI222_X1 U9225 ( .A1(n9340), .A2(n7536), .B1(P1_U3084), .B2(n7535), .C1(
        n9343), .C2(n7534), .ZN(P1_U3324) );
  OAI211_X1 U9226 ( .C1(n7539), .C2(n7538), .A(n7537), .B(n7631), .ZN(n7543)
         );
  AOI22_X1 U9227 ( .A1(n7669), .A2(n8100), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        n4264), .ZN(n7542) );
  AOI22_X1 U9228 ( .A1(n7643), .A2(n8101), .B1(n7657), .B2(n8095), .ZN(n7541)
         );
  NAND2_X1 U9229 ( .A1(n8314), .A2(n7670), .ZN(n7540) );
  NAND4_X1 U9230 ( .A1(n7543), .A2(n7542), .A3(n7541), .A4(n7540), .ZN(
        P2_U3216) );
  INV_X1 U9231 ( .A(n7544), .ZN(n7545) );
  AOI21_X1 U9232 ( .B1(n7547), .B2(n7546), .A(n7545), .ZN(n7553) );
  AOI22_X1 U9233 ( .A1(n7643), .A2(n7908), .B1(n7657), .B2(n7548), .ZN(n7550)
         );
  OAI211_X1 U9234 ( .C1(n7645), .C2(n7683), .A(n7550), .B(n7549), .ZN(n7551)
         );
  AOI21_X1 U9235 ( .B1(n7670), .B2(n7780), .A(n7551), .ZN(n7552) );
  OAI21_X1 U9236 ( .B1(n7553), .B2(n7673), .A(n7552), .ZN(P2_U3217) );
  NAND2_X1 U9237 ( .A1(n7555), .A2(n7554), .ZN(n7557) );
  XNOR2_X1 U9238 ( .A(n7557), .B(n7556), .ZN(n7563) );
  INV_X1 U9239 ( .A(n8154), .ZN(n8058) );
  OAI22_X1 U9240 ( .A1(n7645), .A2(n8058), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7558), .ZN(n7561) );
  INV_X1 U9241 ( .A(n8195), .ZN(n8056) );
  INV_X1 U9242 ( .A(n8158), .ZN(n7559) );
  OAI22_X1 U9243 ( .A1(n7666), .A2(n8056), .B1(n7665), .B2(n7559), .ZN(n7560)
         );
  AOI211_X1 U9244 ( .C1(n8334), .C2(n7670), .A(n7561), .B(n7560), .ZN(n7562)
         );
  OAI21_X1 U9245 ( .B1(n7563), .B2(n7673), .A(n7562), .ZN(P2_U3218) );
  INV_X1 U9246 ( .A(n8358), .ZN(n8228) );
  OAI21_X1 U9247 ( .B1(n7566), .B2(n7565), .A(n7564), .ZN(n7567) );
  NAND2_X1 U9248 ( .A1(n7567), .A2(n7631), .ZN(n7571) );
  AND2_X1 U9249 ( .A1(n4264), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8035) );
  INV_X1 U9250 ( .A(n8225), .ZN(n7568) );
  OAI22_X1 U9251 ( .A1(n7666), .A2(n8254), .B1(n7665), .B2(n7568), .ZN(n7569)
         );
  AOI211_X1 U9252 ( .C1(n7669), .C2(n8196), .A(n8035), .B(n7569), .ZN(n7570)
         );
  OAI211_X1 U9253 ( .C1(n8228), .C2(n7660), .A(n7571), .B(n7570), .ZN(P2_U3221) );
  XNOR2_X1 U9254 ( .A(n7573), .B(n7572), .ZN(n7578) );
  OAI22_X1 U9255 ( .A1(n7645), .A2(n8056), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7574), .ZN(n7576) );
  INV_X1 U9256 ( .A(n8196), .ZN(n8223) );
  OAI22_X1 U9257 ( .A1(n7666), .A2(n8223), .B1(n7665), .B2(n8188), .ZN(n7575)
         );
  AOI211_X1 U9258 ( .C1(n8346), .C2(n7670), .A(n7576), .B(n7575), .ZN(n7577)
         );
  OAI21_X1 U9259 ( .B1(n7578), .B2(n7673), .A(n7577), .ZN(P2_U3225) );
  XNOR2_X1 U9260 ( .A(n7580), .B(n7579), .ZN(n7581) );
  XNOR2_X1 U9261 ( .A(n7582), .B(n7581), .ZN(n7589) );
  NAND2_X1 U9262 ( .A1(n8101), .A2(n9653), .ZN(n7584) );
  NAND2_X1 U9263 ( .A1(n8154), .A2(n9656), .ZN(n7583) );
  NAND2_X1 U9264 ( .A1(n7584), .A2(n7583), .ZN(n8129) );
  INV_X1 U9265 ( .A(n7655), .ZN(n7585) );
  AOI22_X1 U9266 ( .A1(n8129), .A2(n7585), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3152), .ZN(n7586) );
  OAI21_X1 U9267 ( .B1(n7665), .B2(n8124), .A(n7586), .ZN(n7587) );
  AOI21_X1 U9268 ( .B1(n8325), .B2(n7670), .A(n7587), .ZN(n7588) );
  OAI21_X1 U9269 ( .B1(n7589), .B2(n7673), .A(n7588), .ZN(P2_U3227) );
  INV_X1 U9270 ( .A(n8267), .ZN(n8241) );
  INV_X1 U9271 ( .A(n7683), .ZN(n8268) );
  AOI22_X1 U9272 ( .A1(n7643), .A2(n8268), .B1(n7657), .B2(n8273), .ZN(n7591)
         );
  OAI211_X1 U9273 ( .C1(n7645), .C2(n8241), .A(n7591), .B(n7590), .ZN(n7599)
         );
  INV_X1 U9274 ( .A(n7594), .ZN(n7596) );
  NAND3_X1 U9275 ( .A1(n7593), .A2(n7596), .A3(n7595), .ZN(n7597) );
  AOI21_X1 U9276 ( .B1(n7592), .B2(n7597), .A(n7673), .ZN(n7598) );
  AOI211_X1 U9277 ( .C1(n7670), .C2(n8372), .A(n7599), .B(n7598), .ZN(n7600)
         );
  INV_X1 U9278 ( .A(n7600), .ZN(P2_U3228) );
  XNOR2_X1 U9279 ( .A(n7602), .B(n7601), .ZN(n7607) );
  OAI22_X1 U9280 ( .A1(n7645), .A2(n8254), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6058), .ZN(n7605) );
  INV_X1 U9281 ( .A(n8258), .ZN(n7603) );
  OAI22_X1 U9282 ( .A1(n7666), .A2(n8283), .B1(n7665), .B2(n7603), .ZN(n7604)
         );
  AOI211_X1 U9283 ( .C1(n8368), .C2(n7670), .A(n7605), .B(n7604), .ZN(n7606)
         );
  OAI21_X1 U9284 ( .B1(n7607), .B2(n7673), .A(n7606), .ZN(P2_U3230) );
  XNOR2_X1 U9285 ( .A(n7608), .B(n7609), .ZN(n7614) );
  INV_X1 U9286 ( .A(n8140), .ZN(n7686) );
  OAI22_X1 U9287 ( .A1(n7645), .A2(n7686), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7610), .ZN(n7612) );
  OAI22_X1 U9288 ( .A1(n7666), .A2(n8181), .B1(n7665), .B2(n8143), .ZN(n7611)
         );
  AOI211_X1 U9289 ( .C1(n8329), .C2(n7670), .A(n7612), .B(n7611), .ZN(n7613)
         );
  OAI21_X1 U9290 ( .B1(n7614), .B2(n7673), .A(n7613), .ZN(P2_U3231) );
  XNOR2_X1 U9291 ( .A(n7616), .B(n7615), .ZN(n7621) );
  INV_X1 U9292 ( .A(n8211), .ZN(n8180) );
  OAI22_X1 U9293 ( .A1(n7645), .A2(n8180), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7617), .ZN(n7619) );
  OAI22_X1 U9294 ( .A1(n7666), .A2(n8240), .B1(n7665), .B2(n8203), .ZN(n7618)
         );
  AOI211_X1 U9295 ( .C1(n8351), .C2(n7670), .A(n7619), .B(n7618), .ZN(n7620)
         );
  OAI21_X1 U9296 ( .B1(n7621), .B2(n7673), .A(n7620), .ZN(P2_U3235) );
  OAI21_X1 U9297 ( .B1(n7624), .B2(n7623), .A(n7622), .ZN(n7625) );
  NAND2_X1 U9298 ( .A1(n7625), .A2(n7631), .ZN(n7630) );
  OAI22_X1 U9299 ( .A1(n7645), .A2(n8181), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7626), .ZN(n7628) );
  OAI22_X1 U9300 ( .A1(n7666), .A2(n8180), .B1(n7665), .B2(n8172), .ZN(n7627)
         );
  AOI211_X1 U9301 ( .C1(n8341), .C2(n7670), .A(n7628), .B(n7627), .ZN(n7629)
         );
  NAND2_X1 U9302 ( .A1(n7630), .A2(n7629), .ZN(P2_U3237) );
  OAI211_X1 U9303 ( .C1(n7634), .C2(n7633), .A(n7632), .B(n7631), .ZN(n7640)
         );
  AOI22_X1 U9304 ( .A1(n7669), .A2(n7909), .B1(P2_REG3_REG_11__SCAN_IN), .B2(
        P2_U3152), .ZN(n7639) );
  AOI22_X1 U9305 ( .A1(n7643), .A2(n7911), .B1(n7657), .B2(n7635), .ZN(n7638)
         );
  NAND2_X1 U9306 ( .A1(n7670), .A2(n7636), .ZN(n7637) );
  NAND4_X1 U9307 ( .A1(n7640), .A2(n7639), .A3(n7638), .A4(n7637), .ZN(
        P2_U3238) );
  XNOR2_X1 U9308 ( .A(n7642), .B(n7641), .ZN(n7648) );
  AOI22_X1 U9309 ( .A1(n7643), .A2(n8267), .B1(n7657), .B2(n8234), .ZN(n7644)
         );
  NAND2_X1 U9310 ( .A1(P2_U3152), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8014) );
  OAI211_X1 U9311 ( .C1(n7645), .C2(n8240), .A(n7644), .B(n8014), .ZN(n7646)
         );
  AOI21_X1 U9312 ( .B1(n8361), .B2(n7670), .A(n7646), .ZN(n7647) );
  OAI21_X1 U9313 ( .B1(n7648), .B2(n7673), .A(n7647), .ZN(P2_U3240) );
  INV_X1 U9314 ( .A(n8321), .ZN(n8118) );
  AOI21_X1 U9315 ( .B1(n7650), .B2(n7649), .A(n7673), .ZN(n7652) );
  NAND2_X1 U9316 ( .A1(n7652), .A2(n7651), .ZN(n7659) );
  AND2_X1 U9317 ( .A1(n8140), .A2(n9656), .ZN(n7653) );
  AOI21_X1 U9318 ( .B1(n8087), .B2(n9653), .A(n7653), .ZN(n8111) );
  OAI22_X1 U9319 ( .A1(n8111), .A2(n7655), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7654), .ZN(n7656) );
  AOI21_X1 U9320 ( .B1(n8115), .B2(n7657), .A(n7656), .ZN(n7658) );
  OAI211_X1 U9321 ( .C1(n8118), .C2(n7660), .A(n7659), .B(n7658), .ZN(P2_U3242) );
  INV_X1 U9322 ( .A(n7593), .ZN(n7661) );
  AOI21_X1 U9323 ( .B1(n7663), .B2(n7662), .A(n7661), .ZN(n7674) );
  INV_X1 U9324 ( .A(n8291), .ZN(n7664) );
  OAI22_X1 U9325 ( .A1(n7666), .A2(n4522), .B1(n7665), .B2(n7664), .ZN(n7667)
         );
  AOI211_X1 U9326 ( .C1(n7669), .C2(n8050), .A(n7668), .B(n7667), .ZN(n7672)
         );
  NAND2_X1 U9327 ( .A1(n8287), .A2(n7670), .ZN(n7671) );
  OAI211_X1 U9328 ( .C1(n7674), .C2(n7673), .A(n7672), .B(n7671), .ZN(P2_U3243) );
  OR2_X1 U9329 ( .A1(n8039), .A2(n4266), .ZN(n7692) );
  INV_X1 U9330 ( .A(n7692), .ZN(n7693) );
  NAND2_X1 U9331 ( .A1(n8559), .A2(n7701), .ZN(n7676) );
  NAND2_X1 U9332 ( .A1(n7702), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n7675) );
  NAND2_X1 U9333 ( .A1(n6263), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n7681) );
  NAND2_X1 U9334 ( .A1(n7677), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n7680) );
  NAND2_X1 U9335 ( .A1(n7678), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n7679) );
  NAND3_X1 U9336 ( .A1(n7681), .A2(n7680), .A3(n7679), .ZN(n8067) );
  NAND2_X1 U9337 ( .A1(n8304), .A2(n8067), .ZN(n7854) );
  NAND2_X1 U9338 ( .A1(n8287), .A2(n7683), .ZN(n7785) );
  NAND2_X1 U9339 ( .A1(n7786), .A2(n7785), .ZN(n8280) );
  OR2_X1 U9340 ( .A1(n8372), .A2(n8283), .ZN(n7793) );
  NAND2_X1 U9341 ( .A1(n8372), .A2(n8283), .ZN(n7790) );
  NAND2_X1 U9342 ( .A1(n7793), .A2(n7790), .ZN(n8266) );
  INV_X1 U9343 ( .A(n7790), .ZN(n8251) );
  NAND2_X1 U9344 ( .A1(n8368), .A2(n8241), .ZN(n7791) );
  NAND2_X1 U9345 ( .A1(n7792), .A2(n7791), .ZN(n8248) );
  NAND2_X1 U9346 ( .A1(n8361), .A2(n8254), .ZN(n7803) );
  NAND2_X1 U9347 ( .A1(n8218), .A2(n7803), .ZN(n8238) );
  INV_X1 U9348 ( .A(n8218), .ZN(n7798) );
  OR2_X1 U9349 ( .A1(n8358), .A2(n8240), .ZN(n7804) );
  NAND2_X1 U9350 ( .A1(n8358), .A2(n8240), .ZN(n7808) );
  NAND2_X1 U9351 ( .A1(n7804), .A2(n7808), .ZN(n8221) );
  INV_X1 U9352 ( .A(n7808), .ZN(n8207) );
  NAND2_X1 U9353 ( .A1(n8351), .A2(n8223), .ZN(n7807) );
  NAND2_X1 U9354 ( .A1(n7811), .A2(n7807), .ZN(n8208) );
  OR2_X1 U9355 ( .A1(n8346), .A2(n8180), .ZN(n7810) );
  NAND2_X1 U9356 ( .A1(n8346), .A2(n8180), .ZN(n8177) );
  NAND2_X1 U9357 ( .A1(n8341), .A2(n8056), .ZN(n7816) );
  OR2_X1 U9358 ( .A1(n8334), .A2(n8181), .ZN(n7822) );
  NAND2_X1 U9359 ( .A1(n8334), .A2(n8181), .ZN(n8136) );
  OR2_X1 U9360 ( .A1(n8329), .A2(n8058), .ZN(n7684) );
  NAND2_X1 U9361 ( .A1(n8329), .A2(n8058), .ZN(n7824) );
  NAND2_X1 U9362 ( .A1(n7684), .A2(n7824), .ZN(n7890) );
  INV_X1 U9363 ( .A(n8136), .ZN(n7825) );
  NOR2_X1 U9364 ( .A1(n7890), .A2(n7825), .ZN(n7685) );
  INV_X1 U9365 ( .A(n7684), .ZN(n7710) );
  NAND2_X1 U9366 ( .A1(n8325), .A2(n7686), .ZN(n7831) );
  NAND2_X1 U9367 ( .A1(n7828), .A2(n7831), .ZN(n8121) );
  INV_X1 U9368 ( .A(n8101), .ZN(n8059) );
  OR2_X1 U9369 ( .A1(n8321), .A2(n8059), .ZN(n7829) );
  NAND2_X1 U9370 ( .A1(n8321), .A2(n8059), .ZN(n7832) );
  NAND2_X1 U9371 ( .A1(n7829), .A2(n7832), .ZN(n8110) );
  INV_X1 U9372 ( .A(n8087), .ZN(n7839) );
  XNOR2_X1 U9373 ( .A(n8314), .B(n7839), .ZN(n8092) );
  INV_X1 U9374 ( .A(n8314), .ZN(n8097) );
  NAND2_X1 U9375 ( .A1(n8097), .A2(n8087), .ZN(n7837) );
  NAND2_X1 U9376 ( .A1(n8083), .A2(n8100), .ZN(n7838) );
  INV_X1 U9377 ( .A(n7838), .ZN(n7687) );
  NAND2_X1 U9378 ( .A1(n7688), .A2(n7701), .ZN(n7690) );
  NAND2_X1 U9379 ( .A1(n7702), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n7689) );
  INV_X1 U9380 ( .A(n8086), .ZN(n7691) );
  NAND2_X1 U9381 ( .A1(n8305), .A2(n7691), .ZN(n7850) );
  NAND2_X1 U9382 ( .A1(n7696), .A2(n7695), .ZN(n7697) );
  MUX2_X1 U9383 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n7698), .Z(n7699) );
  XNOR2_X1 U9384 ( .A(n7699), .B(SI_31_), .ZN(n7700) );
  NAND2_X1 U9385 ( .A1(n8405), .A2(n7701), .ZN(n7704) );
  NAND2_X1 U9386 ( .A1(n7702), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n7703) );
  OR2_X1 U9387 ( .A1(n8298), .A2(n4654), .ZN(n7858) );
  INV_X1 U9388 ( .A(n8304), .ZN(n8044) );
  INV_X1 U9389 ( .A(n8067), .ZN(n7705) );
  NAND2_X1 U9390 ( .A1(n8044), .A2(n7705), .ZN(n7851) );
  AND2_X1 U9391 ( .A1(n7858), .A2(n7851), .ZN(n7855) );
  AOI21_X1 U9392 ( .B1(n7706), .B2(n7855), .A(n7853), .ZN(n7707) );
  XNOR2_X1 U9393 ( .A(n7707), .B(n7895), .ZN(n7900) );
  NAND2_X1 U9394 ( .A1(n6783), .A2(n7708), .ZN(n7899) );
  INV_X1 U9395 ( .A(n7709), .ZN(n7857) );
  AOI211_X1 U9396 ( .C1(n7710), .C2(n7709), .A(n8121), .B(n8110), .ZN(n7836)
         );
  NAND2_X1 U9397 ( .A1(n7715), .A2(n7711), .ZN(n7714) );
  NAND2_X1 U9398 ( .A1(n7712), .A2(n7733), .ZN(n7713) );
  OAI211_X1 U9399 ( .C1(n7731), .C2(n7716), .A(n7715), .B(n7743), .ZN(n7723)
         );
  INV_X1 U9400 ( .A(n7724), .ZN(n7717) );
  NOR2_X1 U9401 ( .A1(n7717), .A2(n7857), .ZN(n7722) );
  NOR2_X1 U9402 ( .A1(n7727), .A2(n4266), .ZN(n7720) );
  OAI211_X1 U9403 ( .C1(n7720), .C2(n7719), .A(n7718), .B(n7728), .ZN(n7721)
         );
  OAI211_X1 U9404 ( .C1(n7727), .C2(n7726), .A(n7725), .B(n7724), .ZN(n7729)
         );
  NAND3_X1 U9405 ( .A1(n7729), .A2(n7857), .A3(n7728), .ZN(n7730) );
  NAND2_X1 U9406 ( .A1(n7730), .A2(n7734), .ZN(n7739) );
  AOI21_X1 U9407 ( .B1(n7733), .B2(n7732), .A(n7731), .ZN(n7737) );
  INV_X1 U9408 ( .A(n7734), .ZN(n7735) );
  NOR3_X1 U9409 ( .A1(n7737), .A2(n7736), .A3(n7735), .ZN(n7738) );
  OAI22_X1 U9410 ( .A1(n7740), .A2(n7739), .B1(n7738), .B2(n7709), .ZN(n7742)
         );
  INV_X1 U9411 ( .A(n7741), .ZN(n7876) );
  OAI211_X1 U9412 ( .C1(n7743), .C2(n7709), .A(n7742), .B(n7876), .ZN(n7748)
         );
  INV_X1 U9413 ( .A(n7744), .ZN(n7745) );
  MUX2_X1 U9414 ( .A(n7746), .B(n7745), .S(n7709), .Z(n7747) );
  NAND3_X1 U9415 ( .A1(n7748), .A2(n9650), .A3(n7747), .ZN(n7752) );
  MUX2_X1 U9416 ( .A(n7750), .B(n7749), .S(n7709), .Z(n7751) );
  AND3_X1 U9417 ( .A1(n7752), .A2(n7753), .A3(n7751), .ZN(n7765) );
  NAND2_X1 U9418 ( .A1(n7757), .A2(n7758), .ZN(n7755) );
  NAND2_X1 U9419 ( .A1(n7756), .A2(n7753), .ZN(n7754) );
  MUX2_X1 U9420 ( .A(n7755), .B(n7754), .S(n7709), .Z(n7764) );
  NAND2_X1 U9421 ( .A1(n7769), .A2(n7756), .ZN(n7761) );
  OAI211_X1 U9422 ( .C1(n7759), .C2(n7758), .A(n7766), .B(n7757), .ZN(n7760)
         );
  MUX2_X1 U9423 ( .A(n7761), .B(n7760), .S(n7709), .Z(n7762) );
  INV_X1 U9424 ( .A(n7762), .ZN(n7763) );
  OAI21_X1 U9425 ( .B1(n7765), .B2(n7764), .A(n7763), .ZN(n7768) );
  NAND2_X1 U9426 ( .A1(n7768), .A2(n7766), .ZN(n7767) );
  AOI21_X1 U9427 ( .B1(n7767), .B2(n7770), .A(n4520), .ZN(n7775) );
  INV_X1 U9428 ( .A(n7768), .ZN(n7773) );
  NAND2_X1 U9429 ( .A1(n7770), .A2(n7769), .ZN(n7772) );
  OAI21_X1 U9430 ( .B1(n7773), .B2(n7772), .A(n7771), .ZN(n7774) );
  MUX2_X1 U9431 ( .A(n7775), .B(n7774), .S(n7709), .Z(n7779) );
  MUX2_X1 U9432 ( .A(n7777), .B(n7776), .S(n7709), .Z(n7778) );
  OAI211_X1 U9433 ( .C1(n7779), .C2(n7883), .A(n7884), .B(n7778), .ZN(n7784)
         );
  NAND2_X1 U9434 ( .A1(n7907), .A2(n7709), .ZN(n7782) );
  NAND2_X1 U9435 ( .A1(n4522), .A2(n7857), .ZN(n7781) );
  MUX2_X1 U9436 ( .A(n7782), .B(n7781), .S(n7780), .Z(n7783) );
  NAND3_X1 U9437 ( .A1(n7784), .A2(n4680), .A3(n7783), .ZN(n7788) );
  INV_X1 U9438 ( .A(n8266), .ZN(n8263) );
  MUX2_X1 U9439 ( .A(n7786), .B(n7785), .S(n7709), .Z(n7787) );
  NAND3_X1 U9440 ( .A1(n7788), .A2(n8263), .A3(n7787), .ZN(n7789) );
  OAI21_X1 U9441 ( .B1(n7790), .B2(n7709), .A(n7789), .ZN(n7797) );
  INV_X1 U9442 ( .A(n7791), .ZN(n7795) );
  OAI211_X1 U9443 ( .C1(n8248), .C2(n7793), .A(n8218), .B(n7792), .ZN(n7794)
         );
  MUX2_X1 U9444 ( .A(n7795), .B(n7794), .S(n7709), .Z(n7796) );
  AOI21_X1 U9445 ( .B1(n7797), .B2(n4681), .A(n7796), .ZN(n7806) );
  INV_X1 U9446 ( .A(n7804), .ZN(n7799) );
  AOI211_X1 U9447 ( .C1(n7806), .C2(n7803), .A(n7799), .B(n7798), .ZN(n7800)
         );
  OAI21_X1 U9448 ( .B1(n7800), .B2(n8207), .A(n7811), .ZN(n7801) );
  NAND3_X1 U9449 ( .A1(n7801), .A2(n8177), .A3(n7807), .ZN(n7802) );
  NAND3_X1 U9450 ( .A1(n7802), .A2(n7857), .A3(n7810), .ZN(n7815) );
  INV_X1 U9451 ( .A(n7803), .ZN(n7805) );
  OAI21_X1 U9452 ( .B1(n7806), .B2(n7805), .A(n7804), .ZN(n7809) );
  NAND3_X1 U9453 ( .A1(n7809), .A2(n7808), .A3(n7807), .ZN(n7812) );
  NAND3_X1 U9454 ( .A1(n7812), .A2(n7811), .A3(n7810), .ZN(n7813) );
  NAND4_X1 U9455 ( .A1(n7813), .A2(n7709), .A3(n8177), .A4(n7816), .ZN(n7814)
         );
  NAND2_X1 U9456 ( .A1(n7815), .A2(n7814), .ZN(n7821) );
  INV_X1 U9457 ( .A(n7816), .ZN(n7817) );
  INV_X1 U9458 ( .A(n7820), .ZN(n8151) );
  MUX2_X1 U9459 ( .A(n7817), .B(n8151), .S(n7709), .Z(n7819) );
  AOI21_X1 U9460 ( .B1(n8137), .B2(n7822), .A(n7709), .ZN(n7823) );
  OAI21_X1 U9461 ( .B1(n4443), .B2(n7825), .A(n7709), .ZN(n7826) );
  INV_X1 U9462 ( .A(n7832), .ZN(n7827) );
  AOI21_X1 U9463 ( .B1(n7829), .B2(n7828), .A(n7827), .ZN(n7834) );
  INV_X1 U9464 ( .A(n7829), .ZN(n7830) );
  AOI21_X1 U9465 ( .B1(n7832), .B2(n7831), .A(n7830), .ZN(n7833) );
  MUX2_X1 U9466 ( .A(n7834), .B(n7833), .S(n7709), .Z(n7835) );
  AND2_X1 U9467 ( .A1(n7838), .A2(n7837), .ZN(n7841) );
  NAND2_X1 U9468 ( .A1(n8314), .A2(n7839), .ZN(n7840) );
  MUX2_X1 U9469 ( .A(n7841), .B(n7840), .S(n7709), .Z(n7843) );
  OAI211_X1 U9470 ( .C1(n7844), .C2(n8092), .A(n7843), .B(n7842), .ZN(n7848)
         );
  INV_X1 U9471 ( .A(n8100), .ZN(n8060) );
  MUX2_X1 U9472 ( .A(n8309), .B(n8100), .S(n7709), .Z(n7845) );
  OAI21_X1 U9473 ( .B1(n8060), .B2(n8083), .A(n7845), .ZN(n7847) );
  INV_X1 U9474 ( .A(n7850), .ZN(n7846) );
  NOR2_X1 U9475 ( .A1(n7850), .A2(n7709), .ZN(n7852) );
  NAND2_X1 U9476 ( .A1(n7856), .A2(n7854), .ZN(n7893) );
  INV_X1 U9477 ( .A(n7855), .ZN(n7894) );
  NAND3_X1 U9478 ( .A1(n7894), .A2(n7857), .A3(n7856), .ZN(n7860) );
  INV_X1 U9479 ( .A(n7858), .ZN(n7859) );
  AOI22_X1 U9480 ( .A1(n7861), .A2(n7860), .B1(n7859), .B2(n7709), .ZN(n7863)
         );
  INV_X1 U9481 ( .A(n8208), .ZN(n7888) );
  NOR3_X1 U9482 ( .A1(n7867), .A2(n7866), .A3(n7865), .ZN(n7870) );
  INV_X1 U9483 ( .A(n7868), .ZN(n7869) );
  NAND4_X1 U9484 ( .A1(n9679), .A2(n7871), .A3(n7870), .A4(n7869), .ZN(n7875)
         );
  NOR4_X1 U9485 ( .A1(n7875), .A2(n7874), .A3(n7873), .A4(n7872), .ZN(n7879)
         );
  NAND4_X1 U9486 ( .A1(n7879), .A2(n7878), .A3(n7877), .A4(n7876), .ZN(n7880)
         );
  NOR4_X1 U9487 ( .A1(n7883), .A2(n7882), .A3(n7881), .A4(n7880), .ZN(n7885)
         );
  NAND4_X1 U9488 ( .A1(n8263), .A2(n4680), .A3(n7885), .A4(n7884), .ZN(n7886)
         );
  NOR4_X1 U9489 ( .A1(n8221), .A2(n8238), .A3(n8248), .A4(n7886), .ZN(n7887)
         );
  NAND4_X1 U9490 ( .A1(n8176), .A2(n7888), .A3(n8193), .A4(n7887), .ZN(n7889)
         );
  NOR4_X1 U9491 ( .A1(n8121), .A2(n7890), .A3(n8162), .A4(n7889), .ZN(n7891)
         );
  INV_X1 U9492 ( .A(n8092), .ZN(n8098) );
  NAND4_X1 U9493 ( .A1(n8077), .A2(n4688), .A3(n7891), .A4(n8098), .ZN(n7892)
         );
  NOR4_X1 U9494 ( .A1(n7894), .A2(n7893), .A3(n8061), .A4(n7892), .ZN(n7896)
         );
  NOR4_X1 U9495 ( .A1(n9669), .A2(n8413), .A3(n7901), .A4(n8285), .ZN(n7903)
         );
  OAI21_X1 U9496 ( .B1(n7904), .B2(n6250), .A(P2_B_REG_SCAN_IN), .ZN(n7902) );
  OAI22_X1 U9497 ( .A1(n7905), .A2(n7904), .B1(n7903), .B2(n7902), .ZN(
        P2_U3244) );
  MUX2_X1 U9498 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n8067), .S(P2_U3966), .Z(
        P2_U3582) );
  MUX2_X1 U9499 ( .A(n8086), .B(P2_DATAO_REG_29__SCAN_IN), .S(n7906), .Z(
        P2_U3581) );
  MUX2_X1 U9500 ( .A(n8100), .B(P2_DATAO_REG_28__SCAN_IN), .S(n7906), .Z(
        P2_U3580) );
  MUX2_X1 U9501 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8087), .S(P2_U3966), .Z(
        P2_U3579) );
  MUX2_X1 U9502 ( .A(n8101), .B(P2_DATAO_REG_26__SCAN_IN), .S(n7906), .Z(
        P2_U3578) );
  MUX2_X1 U9503 ( .A(n8140), .B(P2_DATAO_REG_25__SCAN_IN), .S(n7906), .Z(
        P2_U3577) );
  MUX2_X1 U9504 ( .A(n8154), .B(P2_DATAO_REG_24__SCAN_IN), .S(n7906), .Z(
        P2_U3576) );
  MUX2_X1 U9505 ( .A(n8139), .B(P2_DATAO_REG_23__SCAN_IN), .S(n7906), .Z(
        P2_U3575) );
  MUX2_X1 U9506 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8195), .S(P2_U3966), .Z(
        P2_U3574) );
  MUX2_X1 U9507 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8211), .S(P2_U3966), .Z(
        P2_U3573) );
  MUX2_X1 U9508 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8196), .S(P2_U3966), .Z(
        P2_U3572) );
  MUX2_X1 U9509 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8210), .S(P2_U3966), .Z(
        P2_U3571) );
  MUX2_X1 U9510 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n8051), .S(P2_U3966), .Z(
        P2_U3570) );
  MUX2_X1 U9511 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8267), .S(P2_U3966), .Z(
        P2_U3569) );
  MUX2_X1 U9512 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8050), .S(P2_U3966), .Z(
        P2_U3568) );
  MUX2_X1 U9513 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n8268), .S(P2_U3966), .Z(
        P2_U3567) );
  MUX2_X1 U9514 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n7907), .S(P2_U3966), .Z(
        P2_U3566) );
  MUX2_X1 U9515 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n7908), .S(P2_U3966), .Z(
        P2_U3565) );
  MUX2_X1 U9516 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n7909), .S(P2_U3966), .Z(
        P2_U3564) );
  MUX2_X1 U9517 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n7910), .S(P2_U3966), .Z(
        P2_U3563) );
  MUX2_X1 U9518 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n7911), .S(P2_U3966), .Z(
        P2_U3562) );
  MUX2_X1 U9519 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n9654), .S(P2_U3966), .Z(
        P2_U3561) );
  MUX2_X1 U9520 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n7912), .S(P2_U3966), .Z(
        P2_U3560) );
  MUX2_X1 U9521 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n9655), .S(P2_U3966), .Z(
        P2_U3559) );
  MUX2_X1 U9522 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n7913), .S(P2_U3966), .Z(
        P2_U3558) );
  MUX2_X1 U9523 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(n7914), .S(P2_U3966), .Z(
        P2_U3557) );
  MUX2_X1 U9524 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n7915), .S(P2_U3966), .Z(
        P2_U3556) );
  MUX2_X1 U9525 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(n7916), .S(P2_U3966), .Z(
        P2_U3555) );
  MUX2_X1 U9526 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(n7917), .S(P2_U3966), .Z(
        P2_U3554) );
  MUX2_X1 U9527 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n7918), .S(P2_U3966), .Z(
        P2_U3553) );
  MUX2_X1 U9528 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n7919), .S(P2_U3966), .Z(
        P2_U3552) );
  OAI211_X1 U9529 ( .C1(n7922), .C2(n7921), .A(n9632), .B(n7920), .ZN(n7933)
         );
  NOR2_X1 U9530 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7923), .ZN(n7924) );
  AOI21_X1 U9531 ( .B1(n9633), .B2(P2_ADDR_REG_3__SCAN_IN), .A(n7924), .ZN(
        n7932) );
  OR2_X1 U9532 ( .A1(n9628), .A2(n7925), .ZN(n7931) );
  AOI21_X1 U9533 ( .B1(n7928), .B2(n7927), .A(n7926), .ZN(n7929) );
  NAND2_X1 U9534 ( .A1(n9627), .A2(n7929), .ZN(n7930) );
  NAND4_X1 U9535 ( .A1(n7933), .A2(n7932), .A3(n7931), .A4(n7930), .ZN(
        P2_U3248) );
  OAI211_X1 U9536 ( .C1(n7936), .C2(n7935), .A(n9632), .B(n7934), .ZN(n7947)
         );
  NOR2_X1 U9537 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7937), .ZN(n7938) );
  AOI21_X1 U9538 ( .B1(n9633), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n7938), .ZN(
        n7946) );
  OR2_X1 U9539 ( .A1(n9628), .A2(n7939), .ZN(n7945) );
  INV_X1 U9540 ( .A(n7940), .ZN(n7941) );
  OAI211_X1 U9541 ( .C1(n7943), .C2(n7942), .A(n9627), .B(n7941), .ZN(n7944)
         );
  NAND4_X1 U9542 ( .A1(n7947), .A2(n7946), .A3(n7945), .A4(n7944), .ZN(
        P2_U3250) );
  OAI211_X1 U9543 ( .C1(n7950), .C2(n7949), .A(n9632), .B(n7948), .ZN(n7960)
         );
  INV_X1 U9544 ( .A(n7951), .ZN(n7952) );
  AOI21_X1 U9545 ( .B1(n9633), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n7952), .ZN(
        n7959) );
  INV_X1 U9546 ( .A(n9628), .ZN(n9363) );
  NAND2_X1 U9547 ( .A1(n9363), .A2(n7953), .ZN(n7958) );
  OAI211_X1 U9548 ( .C1(n7956), .C2(n7955), .A(n9627), .B(n7954), .ZN(n7957)
         );
  NAND4_X1 U9549 ( .A1(n7960), .A2(n7959), .A3(n7958), .A4(n7957), .ZN(
        P2_U3253) );
  OAI211_X1 U9550 ( .C1(n7963), .C2(n7962), .A(n9632), .B(n7961), .ZN(n7974)
         );
  INV_X1 U9551 ( .A(n7964), .ZN(n7965) );
  AOI21_X1 U9552 ( .B1(n9633), .B2(P2_ADDR_REG_9__SCAN_IN), .A(n7965), .ZN(
        n7973) );
  OR2_X1 U9553 ( .A1(n9628), .A2(n7966), .ZN(n7972) );
  AOI21_X1 U9554 ( .B1(n7969), .B2(n7968), .A(n7967), .ZN(n7970) );
  NAND2_X1 U9555 ( .A1(n9627), .A2(n7970), .ZN(n7971) );
  NAND4_X1 U9556 ( .A1(n7974), .A2(n7973), .A3(n7972), .A4(n7971), .ZN(
        P2_U3254) );
  OAI211_X1 U9557 ( .C1(n7977), .C2(n7976), .A(n9632), .B(n7975), .ZN(n7987)
         );
  AOI21_X1 U9558 ( .B1(n9633), .B2(P2_ADDR_REG_10__SCAN_IN), .A(n7978), .ZN(
        n7986) );
  OR2_X1 U9559 ( .A1(n9628), .A2(n7979), .ZN(n7985) );
  AOI21_X1 U9560 ( .B1(n7982), .B2(n7981), .A(n7980), .ZN(n7983) );
  NAND2_X1 U9561 ( .A1(n9627), .A2(n7983), .ZN(n7984) );
  NAND4_X1 U9562 ( .A1(n7987), .A2(n7986), .A3(n7985), .A4(n7984), .ZN(
        P2_U3255) );
  NAND2_X1 U9563 ( .A1(n7989), .A2(n7988), .ZN(n7993) );
  INV_X1 U9564 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n7991) );
  NAND2_X1 U9565 ( .A1(n8013), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n8007) );
  INV_X1 U9566 ( .A(n8007), .ZN(n7990) );
  AOI21_X1 U9567 ( .B1(n7991), .B2(n7995), .A(n7990), .ZN(n7992) );
  NAND2_X1 U9568 ( .A1(n7992), .A2(n7993), .ZN(n8006) );
  OAI211_X1 U9569 ( .C1(n7993), .C2(n7992), .A(n9632), .B(n8006), .ZN(n8005)
         );
  NOR2_X1 U9570 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6058), .ZN(n7994) );
  AOI21_X1 U9571 ( .B1(n9633), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n7994), .ZN(
        n8004) );
  OR2_X1 U9572 ( .A1(n9628), .A2(n7995), .ZN(n8003) );
  XNOR2_X1 U9573 ( .A(n8013), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n8000) );
  OR2_X1 U9574 ( .A1(n7996), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n7998) );
  NAND2_X1 U9575 ( .A1(n7998), .A2(n7997), .ZN(n7999) );
  NOR2_X1 U9576 ( .A1(n8000), .A2(n7999), .ZN(n8012) );
  AOI21_X1 U9577 ( .B1(n8000), .B2(n7999), .A(n8012), .ZN(n8001) );
  NAND2_X1 U9578 ( .A1(n9627), .A2(n8001), .ZN(n8002) );
  NAND4_X1 U9579 ( .A1(n8005), .A2(n8004), .A3(n8003), .A4(n8002), .ZN(
        P2_U3262) );
  NAND2_X1 U9580 ( .A1(n8007), .A2(n8006), .ZN(n8008) );
  AOI21_X1 U9581 ( .B1(n8009), .B2(P2_REG2_REG_18__SCAN_IN), .A(n8022), .ZN(
        n8010) );
  OR2_X1 U9582 ( .A1(n8010), .A2(n8029), .ZN(n8019) );
  INV_X1 U9583 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8011) );
  XNOR2_X1 U9584 ( .A(n8024), .B(n8011), .ZN(n8027) );
  AOI21_X1 U9585 ( .B1(P2_REG1_REG_17__SCAN_IN), .B2(n8013), .A(n8012), .ZN(
        n8026) );
  XNOR2_X1 U9586 ( .A(n8027), .B(n8026), .ZN(n8017) );
  NAND2_X1 U9587 ( .A1(n9633), .A2(P2_ADDR_REG_18__SCAN_IN), .ZN(n8015) );
  NAND2_X1 U9588 ( .A1(n8015), .A2(n8014), .ZN(n8016) );
  AOI21_X1 U9589 ( .B1(n9627), .B2(n8017), .A(n8016), .ZN(n8018) );
  OAI211_X1 U9590 ( .C1(n9628), .C2(n8020), .A(n8019), .B(n8018), .ZN(P2_U3263) );
  NOR2_X1 U9591 ( .A1(n8022), .A2(n8021), .ZN(n8023) );
  INV_X1 U9592 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n9878) );
  XNOR2_X1 U9593 ( .A(n8023), .B(n9878), .ZN(n8034) );
  INV_X1 U9594 ( .A(n8034), .ZN(n8030) );
  NOR2_X1 U9595 ( .A1(n8024), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n8025) );
  AOI21_X1 U9596 ( .B1(n8027), .B2(n8026), .A(n8025), .ZN(n8028) );
  XNOR2_X1 U9597 ( .A(n8028), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n8031) );
  NAND2_X1 U9598 ( .A1(n9627), .A2(n8031), .ZN(n8032) );
  INV_X1 U9599 ( .A(n8305), .ZN(n8070) );
  INV_X1 U9600 ( .A(n8325), .ZN(n8127) );
  OR2_X2 U9601 ( .A1(n8286), .A2(n8287), .ZN(n8288) );
  INV_X1 U9602 ( .A(n8361), .ZN(n8236) );
  INV_X1 U9603 ( .A(n8346), .ZN(n8191) );
  AND2_X1 U9604 ( .A1(n8202), .A2(n8191), .ZN(n8168) );
  INV_X1 U9605 ( .A(n8341), .ZN(n8175) );
  XNOR2_X1 U9606 ( .A(n8298), .B(n4293), .ZN(n8300) );
  INV_X1 U9607 ( .A(P2_B_REG_SCAN_IN), .ZN(n8037) );
  NOR2_X1 U9608 ( .A1(n8413), .A2(n8037), .ZN(n8038) );
  NOR2_X1 U9609 ( .A1(n8284), .A2(n8038), .ZN(n8066) );
  NAND2_X1 U9610 ( .A1(n8066), .A2(n8039), .ZN(n8302) );
  NOR2_X1 U9611 ( .A1(n8278), .A2(n8302), .ZN(n8045) );
  NOR2_X1 U9612 ( .A1(n8040), .A2(n9649), .ZN(n8041) );
  AOI211_X1 U9613 ( .C1(n8278), .C2(P2_REG2_REG_31__SCAN_IN), .A(n8045), .B(
        n8041), .ZN(n8042) );
  OAI21_X1 U9614 ( .B1(n8300), .B2(n8290), .A(n8042), .ZN(P2_U3265) );
  INV_X1 U9615 ( .A(n8068), .ZN(n8043) );
  NAND2_X1 U9616 ( .A1(n8044), .A2(n8043), .ZN(n8301) );
  NAND3_X1 U9617 ( .A1(n8301), .A2(n9647), .A3(n4293), .ZN(n8047) );
  AOI21_X1 U9618 ( .B1(n8278), .B2(P2_REG2_REG_30__SCAN_IN), .A(n8045), .ZN(
        n8046) );
  OAI211_X1 U9619 ( .C1(n8304), .C2(n9649), .A(n8047), .B(n8046), .ZN(P2_U3266) );
  INV_X1 U9620 ( .A(n8329), .ZN(n8146) );
  INV_X1 U9621 ( .A(n8334), .ZN(n8160) );
  NOR2_X1 U9622 ( .A1(n8361), .A2(n8051), .ZN(n8052) );
  OAI21_X1 U9623 ( .B1(n8210), .B2(n8358), .A(n8217), .ZN(n8053) );
  NAND2_X1 U9624 ( .A1(n8187), .A2(n4837), .ZN(n8055) );
  OAI21_X1 U9625 ( .B1(n8211), .B2(n8346), .A(n8055), .ZN(n8167) );
  INV_X1 U9626 ( .A(n8176), .ZN(n8057) );
  OAI21_X1 U9627 ( .B1(n8160), .B2(n8181), .A(n8336), .ZN(n8135) );
  XNOR2_X1 U9628 ( .A(n8062), .B(n8061), .ZN(n8308) );
  NAND2_X1 U9629 ( .A1(n4311), .A2(n9661), .ZN(n8076) );
  INV_X1 U9630 ( .A(n8079), .ZN(n8069) );
  AOI21_X1 U9631 ( .B1(n8305), .B2(n8069), .A(n8068), .ZN(n8306) );
  NOR2_X1 U9632 ( .A1(n8070), .A2(n9649), .ZN(n8074) );
  OAI22_X1 U9633 ( .A1(n9661), .A2(n8072), .B1(n8071), .B2(n8142), .ZN(n8073)
         );
  AOI211_X1 U9634 ( .C1(n8306), .C2(n9647), .A(n8074), .B(n8073), .ZN(n8075)
         );
  OAI211_X1 U9635 ( .C1(n8308), .C2(n6895), .A(n8076), .B(n8075), .ZN(P2_U3267) );
  XNOR2_X1 U9636 ( .A(n8078), .B(n8077), .ZN(n8313) );
  INV_X1 U9637 ( .A(n8094), .ZN(n8080) );
  AOI21_X1 U9638 ( .B1(n8309), .B2(n8080), .A(n8079), .ZN(n8310) );
  AOI22_X1 U9639 ( .A1(n8278), .A2(P2_REG2_REG_28__SCAN_IN), .B1(n8081), .B2(
        n9665), .ZN(n8082) );
  OAI21_X1 U9640 ( .B1(n8083), .B2(n8293), .A(n8082), .ZN(n8090) );
  XNOR2_X1 U9641 ( .A(n8085), .B(n8084), .ZN(n8088) );
  AOI222_X1 U9642 ( .A1(n8213), .A2(n8088), .B1(n8087), .B2(n9656), .C1(n8086), 
        .C2(n9653), .ZN(n8312) );
  NOR2_X1 U9643 ( .A1(n8312), .A2(n8278), .ZN(n8089) );
  OAI21_X1 U9644 ( .B1(n8313), .B2(n6895), .A(n8091), .ZN(P2_U3268) );
  XNOR2_X1 U9645 ( .A(n8093), .B(n8092), .ZN(n8318) );
  AOI21_X1 U9646 ( .B1(n8314), .B2(n8113), .A(n8094), .ZN(n8315) );
  AOI22_X1 U9647 ( .A1(n8278), .A2(P2_REG2_REG_27__SCAN_IN), .B1(n8095), .B2(
        n9665), .ZN(n8096) );
  OAI21_X1 U9648 ( .B1(n8097), .B2(n9649), .A(n8096), .ZN(n8104) );
  XNOR2_X1 U9649 ( .A(n8099), .B(n8098), .ZN(n8102) );
  AOI222_X1 U9650 ( .A1(n8213), .A2(n8102), .B1(n8101), .B2(n9656), .C1(n8100), 
        .C2(n9653), .ZN(n8317) );
  NOR2_X1 U9651 ( .A1(n8317), .A2(n8278), .ZN(n8103) );
  OAI21_X1 U9652 ( .B1(n6895), .B2(n8318), .A(n8105), .ZN(P2_U3269) );
  XNOR2_X1 U9653 ( .A(n8106), .B(n4688), .ZN(n8323) );
  INV_X1 U9654 ( .A(n8107), .ZN(n8108) );
  AOI21_X1 U9655 ( .B1(n8110), .B2(n8109), .A(n8108), .ZN(n8112) );
  OAI21_X1 U9656 ( .B1(n8112), .B2(n9660), .A(n8111), .ZN(n8319) );
  INV_X1 U9657 ( .A(n8113), .ZN(n8114) );
  AOI211_X1 U9658 ( .C1(n8321), .C2(n8122), .A(n9728), .B(n8114), .ZN(n8320)
         );
  NAND2_X1 U9659 ( .A1(n8320), .A2(n8257), .ZN(n8117) );
  AOI22_X1 U9660 ( .A1(n8278), .A2(P2_REG2_REG_26__SCAN_IN), .B1(n8115), .B2(
        n9665), .ZN(n8116) );
  OAI211_X1 U9661 ( .C1(n8118), .C2(n9649), .A(n8117), .B(n8116), .ZN(n8119)
         );
  AOI21_X1 U9662 ( .B1(n8319), .B2(n9661), .A(n8119), .ZN(n8120) );
  OAI21_X1 U9663 ( .B1(n6895), .B2(n8323), .A(n8120), .ZN(P2_U3270) );
  XNOR2_X1 U9664 ( .A(n4296), .B(n8121), .ZN(n8328) );
  INV_X1 U9665 ( .A(n8122), .ZN(n8123) );
  AOI211_X1 U9666 ( .C1(n8325), .C2(n4301), .A(n9728), .B(n8123), .ZN(n8324)
         );
  INV_X1 U9667 ( .A(n8124), .ZN(n8125) );
  AOI22_X1 U9668 ( .A1(n8278), .A2(P2_REG2_REG_25__SCAN_IN), .B1(n8125), .B2(
        n9665), .ZN(n8126) );
  OAI21_X1 U9669 ( .B1(n8127), .B2(n9649), .A(n8126), .ZN(n8132) );
  XNOR2_X1 U9670 ( .A(n8128), .B(n4689), .ZN(n8130) );
  AOI21_X1 U9671 ( .B1(n8130), .B2(n8213), .A(n8129), .ZN(n8327) );
  NOR2_X1 U9672 ( .A1(n8327), .A2(n8278), .ZN(n8131) );
  AOI211_X1 U9673 ( .C1(n8257), .C2(n8324), .A(n8132), .B(n8131), .ZN(n8133)
         );
  OAI21_X1 U9674 ( .B1(n6895), .B2(n8328), .A(n8133), .ZN(P2_U3271) );
  AOI21_X1 U9675 ( .B1(n8137), .B2(n8135), .A(n8134), .ZN(n8333) );
  NAND2_X1 U9676 ( .A1(n8152), .A2(n8136), .ZN(n8138) );
  XNOR2_X1 U9677 ( .A(n8138), .B(n8137), .ZN(n8141) );
  AOI222_X1 U9678 ( .A1(n8213), .A2(n8141), .B1(n8140), .B2(n9653), .C1(n8139), 
        .C2(n9656), .ZN(n8332) );
  OAI21_X1 U9679 ( .B1(n8143), .B2(n8142), .A(n8332), .ZN(n8144) );
  NAND2_X1 U9680 ( .A1(n8144), .A2(n9661), .ZN(n8149) );
  XNOR2_X1 U9681 ( .A(n8146), .B(n8156), .ZN(n8330) );
  OAI22_X1 U9682 ( .A1(n8146), .A2(n8293), .B1(n9661), .B2(n8145), .ZN(n8147)
         );
  AOI21_X1 U9683 ( .B1(n8330), .B2(n9647), .A(n8147), .ZN(n8148) );
  OAI211_X1 U9684 ( .C1(n6895), .C2(n8333), .A(n8149), .B(n8148), .ZN(P2_U3272) );
  INV_X1 U9685 ( .A(n8150), .ZN(n8179) );
  OAI21_X1 U9686 ( .B1(n8179), .B2(n8151), .A(n8162), .ZN(n8153) );
  NAND2_X1 U9687 ( .A1(n8153), .A2(n8152), .ZN(n8155) );
  AOI222_X1 U9688 ( .A1(n8213), .A2(n8155), .B1(n8195), .B2(n9656), .C1(n8154), 
        .C2(n9653), .ZN(n8340) );
  INV_X1 U9689 ( .A(n8156), .ZN(n8157) );
  AOI21_X1 U9690 ( .B1(n8334), .B2(n8169), .A(n8157), .ZN(n8335) );
  AOI22_X1 U9691 ( .A1(n8278), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n8158), .B2(
        n9665), .ZN(n8159) );
  OAI21_X1 U9692 ( .B1(n8160), .B2(n9649), .A(n8159), .ZN(n8161) );
  AOI21_X1 U9693 ( .B1(n8335), .B2(n9647), .A(n8161), .ZN(n8166) );
  OR2_X1 U9694 ( .A1(n8163), .A2(n8162), .ZN(n8337) );
  NAND3_X1 U9695 ( .A1(n8337), .A2(n8336), .A3(n8164), .ZN(n8165) );
  OAI211_X1 U9696 ( .C1(n8340), .C2(n8278), .A(n8166), .B(n8165), .ZN(P2_U3273) );
  XNOR2_X1 U9697 ( .A(n8167), .B(n8176), .ZN(n8345) );
  INV_X1 U9698 ( .A(n8168), .ZN(n8171) );
  INV_X1 U9699 ( .A(n8169), .ZN(n8170) );
  AOI21_X1 U9700 ( .B1(n8341), .B2(n8171), .A(n8170), .ZN(n8342) );
  INV_X1 U9701 ( .A(n8172), .ZN(n8173) );
  AOI22_X1 U9702 ( .A1(n8278), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n8173), .B2(
        n9665), .ZN(n8174) );
  OAI21_X1 U9703 ( .B1(n8175), .B2(n9649), .A(n8174), .ZN(n8185) );
  AOI21_X1 U9704 ( .B1(n8192), .B2(n8177), .A(n8176), .ZN(n8178) );
  NOR3_X1 U9705 ( .A1(n8179), .A2(n8178), .A3(n9660), .ZN(n8183) );
  OAI22_X1 U9706 ( .A1(n8181), .A2(n8284), .B1(n8180), .B2(n8285), .ZN(n8182)
         );
  NOR2_X1 U9707 ( .A1(n8183), .A2(n8182), .ZN(n8344) );
  NOR2_X1 U9708 ( .A1(n8344), .A2(n8278), .ZN(n8184) );
  AOI211_X1 U9709 ( .C1(n8342), .C2(n9647), .A(n8185), .B(n8184), .ZN(n8186)
         );
  OAI21_X1 U9710 ( .B1(n6895), .B2(n8345), .A(n8186), .ZN(P2_U3274) );
  XNOR2_X1 U9711 ( .A(n8187), .B(n8193), .ZN(n8350) );
  XNOR2_X1 U9712 ( .A(n8202), .B(n8346), .ZN(n8347) );
  INV_X1 U9713 ( .A(n8188), .ZN(n8189) );
  AOI22_X1 U9714 ( .A1(n8278), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n8189), .B2(
        n9665), .ZN(n8190) );
  OAI21_X1 U9715 ( .B1(n8191), .B2(n9649), .A(n8190), .ZN(n8199) );
  OAI21_X1 U9716 ( .B1(n8194), .B2(n8193), .A(n8192), .ZN(n8197) );
  AOI222_X1 U9717 ( .A1(n8213), .A2(n8197), .B1(n8196), .B2(n9656), .C1(n8195), 
        .C2(n9653), .ZN(n8349) );
  NOR2_X1 U9718 ( .A1(n8349), .A2(n8278), .ZN(n8198) );
  AOI211_X1 U9719 ( .C1(n8347), .C2(n9647), .A(n8199), .B(n8198), .ZN(n8200)
         );
  OAI21_X1 U9720 ( .B1(n6895), .B2(n8350), .A(n8200), .ZN(P2_U3275) );
  XNOR2_X1 U9721 ( .A(n8201), .B(n8208), .ZN(n8355) );
  AOI21_X1 U9722 ( .B1(n8351), .B2(n8224), .A(n8202), .ZN(n8352) );
  INV_X1 U9723 ( .A(n8351), .ZN(n8206) );
  INV_X1 U9724 ( .A(n8203), .ZN(n8204) );
  AOI22_X1 U9725 ( .A1(n8278), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n8204), .B2(
        n9665), .ZN(n8205) );
  OAI21_X1 U9726 ( .B1(n8206), .B2(n9649), .A(n8205), .ZN(n8215) );
  NOR2_X1 U9727 ( .A1(n8219), .A2(n8207), .ZN(n8209) );
  XNOR2_X1 U9728 ( .A(n8209), .B(n8208), .ZN(n8212) );
  AOI222_X1 U9729 ( .A1(n8213), .A2(n8212), .B1(n8211), .B2(n9653), .C1(n8210), 
        .C2(n9656), .ZN(n8354) );
  NOR2_X1 U9730 ( .A1(n8354), .A2(n8278), .ZN(n8214) );
  AOI211_X1 U9731 ( .C1(n8352), .C2(n9647), .A(n8215), .B(n8214), .ZN(n8216)
         );
  OAI21_X1 U9732 ( .B1(n6895), .B2(n8355), .A(n8216), .ZN(P2_U3276) );
  XNOR2_X1 U9733 ( .A(n8217), .B(n8221), .ZN(n8360) );
  NAND2_X1 U9734 ( .A1(n4512), .A2(n8218), .ZN(n8220) );
  AOI21_X1 U9735 ( .B1(n8221), .B2(n8220), .A(n8219), .ZN(n8222) );
  OAI222_X1 U9736 ( .A1(n8284), .A2(n8223), .B1(n8285), .B2(n8254), .C1(n9660), 
        .C2(n8222), .ZN(n8356) );
  AOI211_X1 U9737 ( .C1(n8358), .C2(n8232), .A(n9728), .B(n4470), .ZN(n8357)
         );
  NAND2_X1 U9738 ( .A1(n8357), .A2(n8257), .ZN(n8227) );
  AOI22_X1 U9739 ( .A1(n8278), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n8225), .B2(
        n9665), .ZN(n8226) );
  OAI211_X1 U9740 ( .C1(n8228), .C2(n9649), .A(n8227), .B(n8226), .ZN(n8229)
         );
  AOI21_X1 U9741 ( .B1(n8356), .B2(n9661), .A(n8229), .ZN(n8230) );
  OAI21_X1 U9742 ( .B1(n6895), .B2(n8360), .A(n8230), .ZN(P2_U3277) );
  XOR2_X1 U9743 ( .A(n8231), .B(n8238), .Z(n8365) );
  INV_X1 U9744 ( .A(n8255), .ZN(n8233) );
  AOI21_X1 U9745 ( .B1(n8361), .B2(n8233), .A(n4471), .ZN(n8362) );
  AOI22_X1 U9746 ( .A1(n8278), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n8234), .B2(
        n9665), .ZN(n8235) );
  OAI21_X1 U9747 ( .B1(n8236), .B2(n9649), .A(n8235), .ZN(n8245) );
  AOI211_X1 U9748 ( .C1(n8239), .C2(n8238), .A(n9660), .B(n8237), .ZN(n8243)
         );
  OAI22_X1 U9749 ( .A1(n8241), .A2(n8285), .B1(n8240), .B2(n8284), .ZN(n8242)
         );
  NOR2_X1 U9750 ( .A1(n8243), .A2(n8242), .ZN(n8364) );
  NOR2_X1 U9751 ( .A1(n8364), .A2(n8278), .ZN(n8244) );
  AOI211_X1 U9752 ( .C1(n8362), .C2(n9647), .A(n8245), .B(n8244), .ZN(n8246)
         );
  OAI21_X1 U9753 ( .B1(n6895), .B2(n8365), .A(n8246), .ZN(P2_U3278) );
  OAI21_X1 U9754 ( .B1(n8249), .B2(n8248), .A(n8247), .ZN(n8250) );
  INV_X1 U9755 ( .A(n8250), .ZN(n8370) );
  NOR2_X1 U9756 ( .A1(n4334), .A2(n8251), .ZN(n8252) );
  XNOR2_X1 U9757 ( .A(n8252), .B(n4681), .ZN(n8253) );
  OAI222_X1 U9758 ( .A1(n8284), .A2(n8254), .B1(n8285), .B2(n8283), .C1(n8253), 
        .C2(n9660), .ZN(n8366) );
  INV_X1 U9759 ( .A(n8272), .ZN(n8256) );
  AOI211_X1 U9760 ( .C1(n8368), .C2(n8256), .A(n9728), .B(n8255), .ZN(n8367)
         );
  NAND2_X1 U9761 ( .A1(n8367), .A2(n8257), .ZN(n8260) );
  AOI22_X1 U9762 ( .A1(n8278), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n8258), .B2(
        n9665), .ZN(n8259) );
  OAI211_X1 U9763 ( .C1(n4726), .C2(n9649), .A(n8260), .B(n8259), .ZN(n8261)
         );
  AOI21_X1 U9764 ( .B1(n8366), .B2(n9661), .A(n8261), .ZN(n8262) );
  OAI21_X1 U9765 ( .B1(n6895), .B2(n8370), .A(n8262), .ZN(P2_U3279) );
  XNOR2_X1 U9766 ( .A(n8264), .B(n8263), .ZN(n8371) );
  AOI21_X1 U9767 ( .B1(n8266), .B2(n8265), .A(n4334), .ZN(n8270) );
  AOI22_X1 U9768 ( .A1(n8268), .A2(n9656), .B1(n9653), .B2(n8267), .ZN(n8269)
         );
  OAI21_X1 U9769 ( .B1(n8270), .B2(n9660), .A(n8269), .ZN(n8271) );
  AOI21_X1 U9770 ( .B1(n9652), .B2(n8371), .A(n8271), .ZN(n8375) );
  AOI21_X1 U9771 ( .B1(n8372), .B2(n8288), .A(n8272), .ZN(n8373) );
  NAND2_X1 U9772 ( .A1(n8373), .A2(n9647), .ZN(n8275) );
  AOI22_X1 U9773 ( .A1(n8278), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n8273), .B2(
        n9665), .ZN(n8274) );
  OAI211_X1 U9774 ( .C1(n4475), .C2(n9649), .A(n8275), .B(n8274), .ZN(n8276)
         );
  AOI21_X1 U9775 ( .B1(n8371), .B2(n9648), .A(n8276), .ZN(n8277) );
  OAI21_X1 U9776 ( .B1(n8375), .B2(n8278), .A(n8277), .ZN(P2_U3280) );
  XNOR2_X1 U9777 ( .A(n8279), .B(n8280), .ZN(n9384) );
  INV_X1 U9778 ( .A(n9384), .ZN(n8297) );
  XNOR2_X1 U9779 ( .A(n8281), .B(n8280), .ZN(n8282) );
  OAI222_X1 U9780 ( .A1(n8285), .A2(n4522), .B1(n8284), .B2(n8283), .C1(n9660), 
        .C2(n8282), .ZN(n9382) );
  INV_X1 U9781 ( .A(n8286), .ZN(n8289) );
  INV_X1 U9782 ( .A(n8287), .ZN(n9380) );
  OAI21_X1 U9783 ( .B1(n8289), .B2(n9380), .A(n8288), .ZN(n9381) );
  NOR2_X1 U9784 ( .A1(n9381), .A2(n8290), .ZN(n8295) );
  AOI22_X1 U9785 ( .A1(n8278), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n8291), .B2(
        n9665), .ZN(n8292) );
  OAI21_X1 U9786 ( .B1(n9380), .B2(n8293), .A(n8292), .ZN(n8294) );
  AOI211_X1 U9787 ( .C1(n9382), .C2(n9661), .A(n8295), .B(n8294), .ZN(n8296)
         );
  OAI21_X1 U9788 ( .B1(n6895), .B2(n8297), .A(n8296), .ZN(P2_U3281) );
  NAND2_X1 U9789 ( .A1(n8298), .A2(n8379), .ZN(n8299) );
  OAI211_X1 U9790 ( .C1(n8300), .C2(n9728), .A(n8299), .B(n8302), .ZN(n8388)
         );
  MUX2_X1 U9791 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n8388), .S(n9752), .Z(
        P2_U3551) );
  NAND3_X1 U9792 ( .A1(n8301), .A2(n8380), .A3(n4293), .ZN(n8303) );
  OAI211_X1 U9793 ( .C1(n8304), .C2(n9727), .A(n8303), .B(n8302), .ZN(n8389)
         );
  MUX2_X1 U9794 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n8389), .S(n9752), .Z(
        P2_U3550) );
  AOI22_X1 U9795 ( .A1(n8306), .A2(n8380), .B1(n8379), .B2(n8305), .ZN(n8307)
         );
  MUX2_X1 U9796 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n8390), .S(n9752), .Z(
        P2_U3549) );
  AOI22_X1 U9797 ( .A1(n8310), .A2(n8380), .B1(n8379), .B2(n8309), .ZN(n8311)
         );
  OAI211_X1 U9798 ( .C1(n9678), .C2(n8313), .A(n8312), .B(n8311), .ZN(n8391)
         );
  MUX2_X1 U9799 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n8391), .S(n9752), .Z(
        P2_U3548) );
  AOI22_X1 U9800 ( .A1(n8315), .A2(n8380), .B1(n8379), .B2(n8314), .ZN(n8316)
         );
  OAI211_X1 U9801 ( .C1(n9678), .C2(n8318), .A(n8317), .B(n8316), .ZN(n8392)
         );
  MUX2_X1 U9802 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n8392), .S(n9752), .Z(
        P2_U3547) );
  AOI211_X1 U9803 ( .C1(n8379), .C2(n8321), .A(n8320), .B(n8319), .ZN(n8322)
         );
  OAI21_X1 U9804 ( .B1(n9678), .B2(n8323), .A(n8322), .ZN(n8393) );
  MUX2_X1 U9805 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n8393), .S(n9752), .Z(
        P2_U3546) );
  AOI21_X1 U9806 ( .B1(n8379), .B2(n8325), .A(n8324), .ZN(n8326) );
  OAI211_X1 U9807 ( .C1(n8328), .C2(n9678), .A(n8327), .B(n8326), .ZN(n8394)
         );
  MUX2_X1 U9808 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n8394), .S(n9752), .Z(
        P2_U3545) );
  AOI22_X1 U9809 ( .A1(n8330), .A2(n8380), .B1(n8379), .B2(n8329), .ZN(n8331)
         );
  OAI211_X1 U9810 ( .C1(n9678), .C2(n8333), .A(n8332), .B(n8331), .ZN(n8395)
         );
  MUX2_X1 U9811 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n8395), .S(n9752), .Z(
        P2_U3544) );
  AOI22_X1 U9812 ( .A1(n8335), .A2(n8380), .B1(n8379), .B2(n8334), .ZN(n8339)
         );
  NAND3_X1 U9813 ( .A1(n8337), .A2(n8336), .A3(n9733), .ZN(n8338) );
  NAND3_X1 U9814 ( .A1(n8340), .A2(n8339), .A3(n8338), .ZN(n8396) );
  MUX2_X1 U9815 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n8396), .S(n9752), .Z(
        P2_U3543) );
  AOI22_X1 U9816 ( .A1(n8342), .A2(n8380), .B1(n8379), .B2(n8341), .ZN(n8343)
         );
  OAI211_X1 U9817 ( .C1(n9678), .C2(n8345), .A(n8344), .B(n8343), .ZN(n8397)
         );
  MUX2_X1 U9818 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n8397), .S(n9752), .Z(
        P2_U3542) );
  AOI22_X1 U9819 ( .A1(n8347), .A2(n8380), .B1(n8379), .B2(n8346), .ZN(n8348)
         );
  OAI211_X1 U9820 ( .C1(n9678), .C2(n8350), .A(n8349), .B(n8348), .ZN(n8398)
         );
  MUX2_X1 U9821 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n8398), .S(n9752), .Z(
        P2_U3541) );
  AOI22_X1 U9822 ( .A1(n8352), .A2(n8380), .B1(n8379), .B2(n8351), .ZN(n8353)
         );
  OAI211_X1 U9823 ( .C1(n9678), .C2(n8355), .A(n8354), .B(n8353), .ZN(n8399)
         );
  MUX2_X1 U9824 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n8399), .S(n9752), .Z(
        P2_U3540) );
  AOI211_X1 U9825 ( .C1(n8379), .C2(n8358), .A(n8357), .B(n8356), .ZN(n8359)
         );
  OAI21_X1 U9826 ( .B1(n9678), .B2(n8360), .A(n8359), .ZN(n8400) );
  MUX2_X1 U9827 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n8400), .S(n9752), .Z(
        P2_U3539) );
  AOI22_X1 U9828 ( .A1(n8362), .A2(n8380), .B1(n8379), .B2(n8361), .ZN(n8363)
         );
  OAI211_X1 U9829 ( .C1(n9678), .C2(n8365), .A(n8364), .B(n8363), .ZN(n8401)
         );
  MUX2_X1 U9830 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n8401), .S(n9752), .Z(
        P2_U3538) );
  AOI211_X1 U9831 ( .C1(n8379), .C2(n8368), .A(n8367), .B(n8366), .ZN(n8369)
         );
  OAI21_X1 U9832 ( .B1(n9678), .B2(n8370), .A(n8369), .ZN(n8402) );
  MUX2_X1 U9833 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n8402), .S(n9752), .Z(
        P2_U3537) );
  INV_X1 U9834 ( .A(n8371), .ZN(n8376) );
  AOI22_X1 U9835 ( .A1(n8373), .A2(n8380), .B1(n8379), .B2(n8372), .ZN(n8374)
         );
  OAI211_X1 U9836 ( .C1(n8376), .C2(n8384), .A(n8375), .B(n8374), .ZN(n8403)
         );
  MUX2_X1 U9837 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n8403), .S(n9752), .Z(
        P2_U3536) );
  INV_X1 U9838 ( .A(n8377), .ZN(n8385) );
  AOI22_X1 U9839 ( .A1(n8381), .A2(n8380), .B1(n8379), .B2(n8378), .ZN(n8382)
         );
  OAI211_X1 U9840 ( .C1(n8385), .C2(n8384), .A(n8383), .B(n8382), .ZN(n8404)
         );
  MUX2_X1 U9841 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n8404), .S(n9752), .Z(
        P2_U3533) );
  MUX2_X1 U9842 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n8386), .S(n9752), .Z(
        P2_U3522) );
  MUX2_X1 U9843 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n8387), .S(n9752), .Z(
        P2_U3521) );
  MUX2_X1 U9844 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n8388), .S(n9736), .Z(
        P2_U3519) );
  MUX2_X1 U9845 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n8389), .S(n9736), .Z(
        P2_U3518) );
  MUX2_X1 U9846 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n8390), .S(n9736), .Z(
        P2_U3517) );
  MUX2_X1 U9847 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n8391), .S(n9736), .Z(
        P2_U3516) );
  MUX2_X1 U9848 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n8392), .S(n9736), .Z(
        P2_U3515) );
  MUX2_X1 U9849 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n8393), .S(n9736), .Z(
        P2_U3514) );
  MUX2_X1 U9850 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n8394), .S(n9736), .Z(
        P2_U3513) );
  MUX2_X1 U9851 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n8395), .S(n9736), .Z(
        P2_U3512) );
  MUX2_X1 U9852 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n8396), .S(n9736), .Z(
        P2_U3511) );
  MUX2_X1 U9853 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n8397), .S(n9736), .Z(
        P2_U3510) );
  MUX2_X1 U9854 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n8398), .S(n9736), .Z(
        P2_U3509) );
  MUX2_X1 U9855 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n8399), .S(n9736), .Z(
        P2_U3508) );
  MUX2_X1 U9856 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n8400), .S(n9736), .Z(
        P2_U3507) );
  MUX2_X1 U9857 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n8401), .S(n9736), .Z(
        P2_U3505) );
  MUX2_X1 U9858 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n8402), .S(n9736), .Z(
        P2_U3502) );
  MUX2_X1 U9859 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n8403), .S(n9736), .Z(
        P2_U3499) );
  MUX2_X1 U9860 ( .A(P2_REG0_REG_13__SCAN_IN), .B(n8404), .S(n9736), .Z(
        P2_U3490) );
  INV_X1 U9861 ( .A(n8405), .ZN(n9334) );
  INV_X1 U9862 ( .A(n8406), .ZN(n8408) );
  NOR4_X1 U9863 ( .A1(n8408), .A2(P2_IR_REG_30__SCAN_IN), .A3(n8407), .A4(
        P2_U3152), .ZN(n8409) );
  AOI21_X1 U9864 ( .B1(n8410), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n8409), .ZN(
        n8411) );
  OAI21_X1 U9865 ( .B1(n9334), .B2(n8414), .A(n8411), .ZN(P2_U3327) );
  INV_X1 U9866 ( .A(n8412), .ZN(n9338) );
  OAI222_X1 U9867 ( .A1(n8417), .A2(n8415), .B1(n8414), .B2(n9338), .C1(n8413), 
        .C2(P2_U3152), .ZN(P2_U3331) );
  INV_X1 U9868 ( .A(n8416), .ZN(n9342) );
  OAI222_X1 U9869 ( .A1(n4264), .A2(n8419), .B1(n8414), .B2(n9342), .C1(n8418), 
        .C2(n8417), .ZN(P2_U3332) );
  MUX2_X1 U9870 ( .A(n8420), .B(n9638), .S(P2_STATE_REG_SCAN_IN), .Z(P2_U3358)
         );
  NAND2_X1 U9871 ( .A1(n8422), .A2(n8421), .ZN(n8423) );
  XOR2_X1 U9872 ( .A(n8424), .B(n8423), .Z(n8432) );
  NOR2_X1 U9873 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n8425), .ZN(n9512) );
  NOR2_X1 U9874 ( .A1(n8545), .A2(n9441), .ZN(n8426) );
  AOI211_X1 U9875 ( .C1(n8523), .C2(n9255), .A(n9512), .B(n8426), .ZN(n8427)
         );
  OAI21_X1 U9876 ( .B1(n8550), .B2(n8428), .A(n8427), .ZN(n8429) );
  AOI21_X1 U9877 ( .B1(n8552), .B2(n8430), .A(n8429), .ZN(n8431) );
  OAI21_X1 U9878 ( .B1(n8432), .B2(n8554), .A(n8431), .ZN(P1_U3213) );
  NAND2_X1 U9879 ( .A1(n4815), .A2(n8433), .ZN(n8435) );
  XNOR2_X1 U9880 ( .A(n8435), .B(n8434), .ZN(n8442) );
  OAI22_X1 U9881 ( .A1(n8545), .A2(n8437), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8436), .ZN(n8438) );
  AOI21_X1 U9882 ( .B1(n8548), .B2(n9023), .A(n8438), .ZN(n8439) );
  OAI21_X1 U9883 ( .B1(n8550), .B2(n9027), .A(n8439), .ZN(n8440) );
  AOI21_X1 U9884 ( .B1(n9210), .B2(n8552), .A(n8440), .ZN(n8441) );
  OAI21_X1 U9885 ( .B1(n8442), .B2(n8554), .A(n8441), .ZN(P1_U3214) );
  XOR2_X1 U9886 ( .A(n8443), .B(n8444), .Z(n8449) );
  AOI22_X1 U9887 ( .A1(n8523), .A2(n9232), .B1(P1_REG3_REG_19__SCAN_IN), .B2(
        P1_U3084), .ZN(n8446) );
  NAND2_X1 U9888 ( .A1(n8534), .A2(n9233), .ZN(n8445) );
  OAI211_X1 U9889 ( .C1(n8550), .C2(n9083), .A(n8446), .B(n8445), .ZN(n8447)
         );
  AOI21_X1 U9890 ( .B1(n9231), .B2(n8552), .A(n8447), .ZN(n8448) );
  OAI21_X1 U9891 ( .B1(n8449), .B2(n8554), .A(n8448), .ZN(P1_U3217) );
  XOR2_X1 U9892 ( .A(n8452), .B(n8451), .Z(n8458) );
  AOI22_X1 U9893 ( .A1(n8523), .A2(n9218), .B1(P1_REG3_REG_21__SCAN_IN), .B2(
        P1_U3084), .ZN(n8454) );
  NAND2_X1 U9894 ( .A1(n8534), .A2(n9232), .ZN(n8453) );
  OAI211_X1 U9895 ( .C1(n8550), .C2(n9055), .A(n8454), .B(n8453), .ZN(n8455)
         );
  AOI21_X1 U9896 ( .B1(n8456), .B2(n8552), .A(n8455), .ZN(n8457) );
  OAI21_X1 U9897 ( .B1(n8458), .B2(n8554), .A(n8457), .ZN(P1_U3221) );
  AOI22_X1 U9898 ( .A1(n8523), .A2(n8999), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3084), .ZN(n8461) );
  NAND2_X1 U9899 ( .A1(n9023), .A2(n8534), .ZN(n8460) );
  OAI211_X1 U9900 ( .C1(n8991), .C2(n8550), .A(n8461), .B(n8460), .ZN(n8462)
         );
  AOI21_X1 U9901 ( .B1(n8990), .B2(n8552), .A(n8462), .ZN(n8463) );
  OAI21_X1 U9902 ( .B1(n8464), .B2(n8554), .A(n8463), .ZN(P1_U3223) );
  XOR2_X1 U9903 ( .A(n8465), .B(n8466), .Z(n8471) );
  AOI22_X1 U9904 ( .A1(n8523), .A2(n9256), .B1(P1_REG3_REG_16__SCAN_IN), .B2(
        P1_U3084), .ZN(n8468) );
  NAND2_X1 U9905 ( .A1(n8534), .A2(n9255), .ZN(n8467) );
  OAI211_X1 U9906 ( .C1(n8550), .C2(n9133), .A(n8468), .B(n8467), .ZN(n8469)
         );
  AOI21_X1 U9907 ( .B1(n9254), .B2(n8552), .A(n8469), .ZN(n8470) );
  OAI21_X1 U9908 ( .B1(n8471), .B2(n8554), .A(n8470), .ZN(P1_U3224) );
  OAI21_X1 U9909 ( .B1(n8474), .B2(n8473), .A(n8472), .ZN(n8476) );
  NAND2_X1 U9910 ( .A1(n8476), .A2(n8475), .ZN(n8482) );
  AND2_X1 U9911 ( .A1(P1_U3084), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n8864) );
  AOI21_X1 U9912 ( .B1(n8552), .B2(n8477), .A(n8864), .ZN(n8481) );
  AOI22_X1 U9913 ( .A1(n8534), .A2(n8847), .B1(n8548), .B2(n8846), .ZN(n8480)
         );
  NAND2_X1 U9914 ( .A1(n8499), .A2(n8478), .ZN(n8479) );
  NAND4_X1 U9915 ( .A1(n8482), .A2(n8481), .A3(n8480), .A4(n8479), .ZN(
        P1_U3225) );
  XOR2_X1 U9916 ( .A(n8484), .B(n8483), .Z(n8489) );
  AOI22_X1 U9917 ( .A1(n8523), .A2(n9233), .B1(P1_REG3_REG_17__SCAN_IN), .B2(
        P1_U3084), .ZN(n8486) );
  NAND2_X1 U9918 ( .A1(n8534), .A2(n9265), .ZN(n8485) );
  OAI211_X1 U9919 ( .C1(n8550), .C2(n9114), .A(n8486), .B(n8485), .ZN(n8487)
         );
  AOI21_X1 U9920 ( .B1(n9126), .B2(n8552), .A(n8487), .ZN(n8488) );
  OAI21_X1 U9921 ( .B1(n8489), .B2(n8554), .A(n8488), .ZN(P1_U3226) );
  XOR2_X1 U9922 ( .A(n8491), .B(n8490), .Z(n8496) );
  AOI22_X1 U9923 ( .A1(n8523), .A2(n9013), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3084), .ZN(n8493) );
  NAND2_X1 U9924 ( .A1(n8499), .A2(n9010), .ZN(n8492) );
  OAI211_X1 U9925 ( .C1(n9201), .C2(n8545), .A(n8493), .B(n8492), .ZN(n8494)
         );
  AOI21_X1 U9926 ( .B1(n9204), .B2(n8552), .A(n8494), .ZN(n8495) );
  OAI21_X1 U9927 ( .B1(n8496), .B2(n8554), .A(n8495), .ZN(P1_U3227) );
  XOR2_X1 U9928 ( .A(n8497), .B(n8498), .Z(n8504) );
  AOI22_X1 U9929 ( .A1(n8523), .A2(n9038), .B1(P1_REG3_REG_20__SCAN_IN), .B2(
        P1_U3084), .ZN(n8501) );
  NAND2_X1 U9930 ( .A1(n8499), .A2(n9072), .ZN(n8500) );
  OAI211_X1 U9931 ( .C1(n9104), .C2(n8545), .A(n8501), .B(n8500), .ZN(n8502)
         );
  AOI21_X1 U9932 ( .B1(n9228), .B2(n8552), .A(n8502), .ZN(n8503) );
  OAI21_X1 U9933 ( .B1(n8504), .B2(n8554), .A(n8503), .ZN(P1_U3231) );
  INV_X1 U9934 ( .A(n8505), .ZN(n8512) );
  INV_X1 U9935 ( .A(n8506), .ZN(n8508) );
  NAND2_X1 U9936 ( .A1(n8508), .A2(n8507), .ZN(n8510) );
  AOI22_X1 U9937 ( .A1(n8512), .A2(n8511), .B1(n8510), .B2(n8509), .ZN(n8518)
         );
  OAI22_X1 U9938 ( .A1(n8545), .A2(n9069), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8513), .ZN(n8514) );
  AOI21_X1 U9939 ( .B1(n9039), .B2(n8548), .A(n8514), .ZN(n8515) );
  OAI21_X1 U9940 ( .B1(n8550), .B2(n9043), .A(n8515), .ZN(n8516) );
  AOI21_X1 U9941 ( .B1(n9215), .B2(n8552), .A(n8516), .ZN(n8517) );
  OAI21_X1 U9942 ( .B1(n8518), .B2(n8554), .A(n8517), .ZN(P1_U3233) );
  NAND2_X1 U9943 ( .A1(n8520), .A2(n8519), .ZN(n8521) );
  XOR2_X1 U9944 ( .A(n8522), .B(n8521), .Z(n8528) );
  NOR2_X1 U9945 ( .A1(n8550), .A2(n9100), .ZN(n8526) );
  NAND2_X1 U9946 ( .A1(n8523), .A2(n9242), .ZN(n8524) );
  NAND2_X1 U9947 ( .A1(P1_U3084), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9531) );
  OAI211_X1 U9948 ( .C1(n9139), .C2(n8545), .A(n8524), .B(n9531), .ZN(n8525)
         );
  AOI211_X1 U9949 ( .C1(n9241), .C2(n8552), .A(n8526), .B(n8525), .ZN(n8527)
         );
  OAI21_X1 U9950 ( .B1(n8528), .B2(n8554), .A(n8527), .ZN(P1_U3236) );
  INV_X1 U9951 ( .A(n8529), .ZN(n8530) );
  NOR2_X1 U9952 ( .A1(n8531), .A2(n8530), .ZN(n8532) );
  XNOR2_X1 U9953 ( .A(n8533), .B(n8532), .ZN(n8539) );
  AOI22_X1 U9954 ( .A1(n8534), .A2(n9013), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3084), .ZN(n8536) );
  NAND2_X1 U9955 ( .A1(n8548), .A2(n9176), .ZN(n8535) );
  OAI211_X1 U9956 ( .C1(n8550), .C2(n8974), .A(n8536), .B(n8535), .ZN(n8537)
         );
  AOI21_X1 U9957 ( .B1(n8973), .B2(n8552), .A(n8537), .ZN(n8538) );
  OAI21_X1 U9958 ( .B1(n8539), .B2(n8554), .A(n8538), .ZN(P1_U3238) );
  NAND2_X1 U9959 ( .A1(n8540), .A2(n8541), .ZN(n8542) );
  XOR2_X1 U9960 ( .A(n8543), .B(n8542), .Z(n8555) );
  INV_X1 U9961 ( .A(n8544), .ZN(n8547) );
  NOR2_X1 U9962 ( .A1(n8545), .A2(n9402), .ZN(n8546) );
  AOI211_X1 U9963 ( .C1(n8548), .C2(n9265), .A(n8547), .B(n8546), .ZN(n8549)
         );
  OAI21_X1 U9964 ( .B1(n8550), .B2(n9152), .A(n8549), .ZN(n8551) );
  AOI21_X1 U9965 ( .B1(n8552), .B2(n9264), .A(n8551), .ZN(n8553) );
  OAI21_X1 U9966 ( .B1(n8555), .B2(n8554), .A(n8553), .ZN(P1_U3239) );
  NOR3_X1 U9967 ( .A1(n8557), .A2(n8556), .A3(n9463), .ZN(n8840) );
  OAI21_X1 U9968 ( .B1(n8558), .B2(n8829), .A(P1_B_REG_SCAN_IN), .ZN(n8839) );
  AND2_X1 U9969 ( .A1(n4265), .A2(n9074), .ZN(n8674) );
  INV_X1 U9970 ( .A(n8674), .ZN(n8679) );
  NAND2_X1 U9971 ( .A1(n8559), .A2(n8563), .ZN(n8562) );
  OR2_X1 U9972 ( .A1(n5000), .A2(n8560), .ZN(n8561) );
  INV_X1 U9973 ( .A(n8841), .ZN(n8685) );
  OR2_X1 U9974 ( .A1(n8916), .A2(n8685), .ZN(n8683) );
  NAND2_X1 U9975 ( .A1(n8683), .A2(n8912), .ZN(n8566) );
  NAND2_X1 U9976 ( .A1(n8405), .A2(n8563), .ZN(n8565) );
  OR2_X1 U9977 ( .A1(n5000), .A2(n6334), .ZN(n8564) );
  AND2_X1 U9978 ( .A1(n8566), .A2(n8908), .ZN(n8568) );
  INV_X1 U9979 ( .A(n8568), .ZN(n8793) );
  NOR2_X1 U9980 ( .A1(n8568), .A2(n8926), .ZN(n8567) );
  MUX2_X1 U9981 ( .A(n9175), .B(n8567), .S(n8679), .Z(n8670) );
  NOR3_X1 U9982 ( .A1(n8568), .A2(n8786), .A3(n9175), .ZN(n8669) );
  INV_X1 U9983 ( .A(n8691), .ZN(n8570) );
  OAI211_X1 U9984 ( .C1(n8571), .C2(n8570), .A(n8569), .B(n8689), .ZN(n8572)
         );
  NAND2_X1 U9985 ( .A1(n8572), .A2(n8692), .ZN(n8575) );
  INV_X1 U9986 ( .A(n8739), .ZN(n8573) );
  AOI21_X1 U9987 ( .B1(n8575), .B2(n8771), .A(n8573), .ZN(n8574) );
  MUX2_X1 U9988 ( .A(n8771), .B(n8574), .S(n8679), .Z(n8578) );
  INV_X1 U9989 ( .A(n8575), .ZN(n8576) );
  NAND3_X1 U9990 ( .A1(n8576), .A2(n8674), .A3(n8739), .ZN(n8577) );
  NAND2_X1 U9991 ( .A1(n8578), .A2(n8577), .ZN(n8581) );
  NAND2_X1 U9992 ( .A1(n8581), .A2(n9544), .ZN(n8579) );
  NAND3_X1 U9993 ( .A1(n8579), .A2(n8740), .A3(n8702), .ZN(n8580) );
  NAND3_X1 U9994 ( .A1(n8580), .A2(n8755), .A3(n8701), .ZN(n8586) );
  NAND2_X1 U9995 ( .A1(n8581), .A2(n8740), .ZN(n8582) );
  NAND2_X1 U9996 ( .A1(n8582), .A2(n8756), .ZN(n8584) );
  INV_X1 U9997 ( .A(n8757), .ZN(n8583) );
  NAND2_X1 U9998 ( .A1(n8584), .A2(n8583), .ZN(n8585) );
  MUX2_X1 U9999 ( .A(n8586), .B(n8585), .S(n8674), .Z(n8593) );
  INV_X1 U10000 ( .A(n8587), .ZN(n8589) );
  NAND2_X1 U10001 ( .A1(n8608), .A2(n8755), .ZN(n8588) );
  MUX2_X1 U10002 ( .A(n8589), .B(n8588), .S(n8674), .Z(n8591) );
  NAND2_X1 U10003 ( .A1(n8607), .A2(n9416), .ZN(n8590) );
  NOR2_X1 U10004 ( .A1(n8591), .A2(n8590), .ZN(n8592) );
  NAND2_X1 U10005 ( .A1(n8593), .A2(n8592), .ZN(n8610) );
  AND2_X1 U10006 ( .A1(n8611), .A2(n8594), .ZN(n8761) );
  NAND2_X1 U10007 ( .A1(n8614), .A2(n8595), .ZN(n8605) );
  AOI21_X1 U10008 ( .B1(n8610), .B2(n8761), .A(n8605), .ZN(n8596) );
  INV_X1 U10009 ( .A(n8612), .ZN(n8762) );
  NOR2_X1 U10010 ( .A1(n8596), .A2(n8762), .ZN(n8620) );
  NAND4_X1 U10011 ( .A1(n9125), .A2(n8767), .A3(n8744), .A4(n8679), .ZN(n8619)
         );
  NAND2_X1 U10012 ( .A1(n8623), .A2(n8597), .ZN(n8770) );
  INV_X1 U10013 ( .A(n9125), .ZN(n9115) );
  NAND3_X1 U10014 ( .A1(n8767), .A2(n8674), .A3(n8744), .ZN(n8598) );
  OAI21_X1 U10015 ( .B1(n9116), .B2(n8679), .A(n8598), .ZN(n8603) );
  NOR2_X1 U10016 ( .A1(n8765), .A2(n8674), .ZN(n8599) );
  AOI22_X1 U10017 ( .A1(n8746), .A2(n8679), .B1(n8599), .B2(n9116), .ZN(n8601)
         );
  NAND2_X1 U10018 ( .A1(n8621), .A2(n8600), .ZN(n8725) );
  AOI21_X1 U10019 ( .B1(n9125), .B2(n8601), .A(n8725), .ZN(n8602) );
  AOI211_X1 U10020 ( .C1(n8674), .C2(n9115), .A(n8603), .B(n8602), .ZN(n8604)
         );
  AOI21_X1 U10021 ( .B1(n8674), .B2(n8770), .A(n8604), .ZN(n8618) );
  INV_X1 U10022 ( .A(n8605), .ZN(n8764) );
  NAND2_X1 U10023 ( .A1(n8607), .A2(n8606), .ZN(n8754) );
  NAND2_X1 U10024 ( .A1(n8754), .A2(n8608), .ZN(n8609) );
  NAND3_X1 U10025 ( .A1(n8610), .A2(n8764), .A3(n8609), .ZN(n8616) );
  NAND2_X1 U10026 ( .A1(n8612), .A2(n8611), .ZN(n8613) );
  AOI211_X1 U10027 ( .C1(n8614), .C2(n8613), .A(n8679), .B(n8765), .ZN(n8615)
         );
  NAND4_X1 U10028 ( .A1(n8616), .A2(n9125), .A3(n8615), .A4(n9116), .ZN(n8617)
         );
  OAI211_X1 U10029 ( .C1(n8620), .C2(n8619), .A(n8618), .B(n8617), .ZN(n8625)
         );
  NAND3_X1 U10030 ( .A1(n8625), .A2(n8621), .A3(n8624), .ZN(n8622) );
  AND2_X1 U10031 ( .A1(n8772), .A2(n8623), .ZN(n8726) );
  NAND2_X1 U10032 ( .A1(n8627), .A2(n8624), .ZN(n8727) );
  AOI21_X1 U10033 ( .B1(n8625), .B2(n8726), .A(n8727), .ZN(n8626) );
  NAND2_X1 U10034 ( .A1(n8628), .A2(n8633), .ZN(n8630) );
  INV_X1 U10035 ( .A(n8636), .ZN(n8629) );
  INV_X1 U10036 ( .A(n8631), .ZN(n8632) );
  NAND2_X1 U10037 ( .A1(n8729), .A2(n8632), .ZN(n8634) );
  AND2_X1 U10038 ( .A1(n8634), .A2(n8633), .ZN(n8635) );
  NAND2_X1 U10039 ( .A1(n8636), .A2(n8635), .ZN(n8724) );
  AOI21_X1 U10040 ( .B1(n8637), .B2(n8729), .A(n8724), .ZN(n8639) );
  INV_X1 U10041 ( .A(n8638), .ZN(n8732) );
  NOR2_X1 U10042 ( .A1(n8639), .A2(n8732), .ZN(n8640) );
  INV_X1 U10043 ( .A(n8996), .ZN(n8645) );
  INV_X1 U10044 ( .A(n8642), .ZN(n8643) );
  NAND2_X1 U10045 ( .A1(n4333), .A2(n8643), .ZN(n8644) );
  NAND3_X1 U10046 ( .A1(n8655), .A2(n8645), .A3(n8644), .ZN(n8775) );
  AND2_X1 U10047 ( .A1(n4333), .A2(n8734), .ZN(n8646) );
  OAI21_X1 U10048 ( .B1(n8646), .B2(n8996), .A(n8737), .ZN(n8647) );
  MUX2_X1 U10049 ( .A(n8775), .B(n8647), .S(n8679), .Z(n8648) );
  INV_X1 U10050 ( .A(n8780), .ZN(n8649) );
  AOI21_X1 U10051 ( .B1(n8973), .B2(n8737), .A(n8649), .ZN(n8652) );
  AOI21_X1 U10052 ( .B1(n8999), .B2(n8655), .A(n8650), .ZN(n8651) );
  MUX2_X1 U10053 ( .A(n8652), .B(n8651), .S(n8679), .Z(n8653) );
  AOI21_X1 U10054 ( .B1(n8660), .B2(n8964), .A(n8653), .ZN(n8663) );
  OAI21_X1 U10055 ( .B1(n8973), .B2(n8737), .A(n8654), .ZN(n8657) );
  INV_X1 U10056 ( .A(n8973), .ZN(n9295) );
  OAI21_X1 U10057 ( .B1(n8999), .B2(n8655), .A(n9295), .ZN(n8656) );
  MUX2_X1 U10058 ( .A(n8657), .B(n8656), .S(n8679), .Z(n8658) );
  AOI21_X1 U10059 ( .B1(n8660), .B2(n8659), .A(n8658), .ZN(n8662) );
  MUX2_X1 U10060 ( .A(n8937), .B(n8780), .S(n8679), .Z(n8661) );
  OAI21_X1 U10061 ( .B1(n8663), .B2(n8662), .A(n8661), .ZN(n8664) );
  NAND2_X1 U10062 ( .A1(n8664), .A2(n8932), .ZN(n8666) );
  MUX2_X1 U10063 ( .A(n8783), .B(n8722), .S(n8674), .Z(n8665) );
  NAND2_X1 U10064 ( .A1(n8666), .A2(n8665), .ZN(n8668) );
  NAND2_X1 U10065 ( .A1(n8841), .A2(n8912), .ZN(n8667) );
  NAND2_X1 U10066 ( .A1(n8916), .A2(n8667), .ZN(n8790) );
  INV_X1 U10067 ( .A(n8790), .ZN(n8673) );
  INV_X1 U10068 ( .A(n9175), .ZN(n8785) );
  NOR2_X1 U10069 ( .A1(n8786), .A2(n8785), .ZN(n8721) );
  NOR3_X1 U10070 ( .A1(n8926), .A2(n8674), .A3(n9175), .ZN(n8671) );
  AOI21_X1 U10071 ( .B1(n8674), .B2(n8721), .A(n8671), .ZN(n8672) );
  NOR2_X1 U10072 ( .A1(n8673), .A2(n8672), .ZN(n8677) );
  NOR2_X1 U10073 ( .A1(n8790), .A2(n8674), .ZN(n8676) );
  INV_X1 U10074 ( .A(n8912), .ZN(n8675) );
  NAND2_X1 U10075 ( .A1(n8908), .A2(n8675), .ZN(n8684) );
  AOI22_X1 U10076 ( .A1(n8677), .A2(n8793), .B1(n8676), .B2(n8684), .ZN(n8678)
         );
  NAND2_X1 U10077 ( .A1(n4265), .A2(n5621), .ZN(n8682) );
  AND2_X1 U10078 ( .A1(n9284), .A2(n8912), .ZN(n8794) );
  INV_X1 U10079 ( .A(n8680), .ZN(n8681) );
  NAND2_X1 U10080 ( .A1(n8684), .A2(n8683), .ZN(n8827) );
  AND2_X1 U10081 ( .A1(n8916), .A2(n8685), .ZN(n8822) );
  INV_X1 U10082 ( .A(n8822), .ZN(n8718) );
  INV_X1 U10083 ( .A(n9034), .ZN(n9037) );
  INV_X1 U10084 ( .A(n9397), .ZN(n9396) );
  NAND2_X1 U10085 ( .A1(n8687), .A2(n8686), .ZN(n8690) );
  NAND3_X1 U10086 ( .A1(n8690), .A2(n8689), .A3(n8688), .ZN(n8693) );
  AND3_X1 U10087 ( .A1(n8693), .A2(n8692), .A3(n8691), .ZN(n8748) );
  NAND3_X1 U10088 ( .A1(n8748), .A2(n8695), .A3(n4267), .ZN(n8699) );
  NAND3_X1 U10089 ( .A1(n8810), .A2(n8697), .A3(n8696), .ZN(n8698) );
  NOR2_X1 U10090 ( .A1(n8699), .A2(n8698), .ZN(n8705) );
  INV_X1 U10091 ( .A(n8700), .ZN(n8703) );
  NAND4_X1 U10092 ( .A1(n8705), .A2(n8704), .A3(n8703), .A4(n9556), .ZN(n8707)
         );
  NOR2_X1 U10093 ( .A1(n8707), .A2(n8706), .ZN(n8708) );
  NAND4_X1 U10094 ( .A1(n8709), .A2(n9396), .A3(n8708), .A4(n9416), .ZN(n8710)
         );
  NOR3_X1 U10095 ( .A1(n9132), .A2(n9150), .A3(n8710), .ZN(n8711) );
  NAND4_X1 U10096 ( .A1(n9082), .A2(n4580), .A3(n9125), .A4(n8711), .ZN(n8712)
         );
  NOR3_X1 U10097 ( .A1(n9054), .A2(n9066), .A3(n8712), .ZN(n8713) );
  NAND3_X1 U10098 ( .A1(n9021), .A2(n9037), .A3(n8713), .ZN(n8714) );
  NOR3_X1 U10099 ( .A1(n8995), .A2(n9007), .A3(n8714), .ZN(n8715) );
  AND4_X1 U10100 ( .A1(n8932), .A2(n8964), .A3(n8979), .A4(n8715), .ZN(n8717)
         );
  NAND3_X1 U10101 ( .A1(n8718), .A2(n8717), .A3(n8716), .ZN(n8719) );
  OR3_X1 U10102 ( .A1(n8794), .A2(n8827), .A3(n8719), .ZN(n8720) );
  NAND2_X1 U10103 ( .A1(n8720), .A2(n8801), .ZN(n8799) );
  INV_X1 U10104 ( .A(n8721), .ZN(n8723) );
  NAND2_X1 U10105 ( .A1(n8723), .A2(n8722), .ZN(n8800) );
  INV_X1 U10106 ( .A(n8724), .ZN(n8773) );
  INV_X1 U10107 ( .A(n8725), .ZN(n8731) );
  INV_X1 U10108 ( .A(n8726), .ZN(n8730) );
  INV_X1 U10109 ( .A(n8727), .ZN(n8728) );
  OAI211_X1 U10110 ( .C1(n8731), .C2(n8730), .A(n8729), .B(n8728), .ZN(n8733)
         );
  AOI21_X1 U10111 ( .B1(n8773), .B2(n8733), .A(n8732), .ZN(n8735) );
  AND3_X1 U10112 ( .A1(n4333), .A2(n8735), .A3(n8734), .ZN(n8738) );
  OAI211_X1 U10113 ( .C1(n8775), .C2(n8738), .A(n8737), .B(n8736), .ZN(n8819)
         );
  INV_X1 U10114 ( .A(n8819), .ZN(n8778) );
  NAND3_X1 U10115 ( .A1(n8741), .A2(n8740), .A3(n8739), .ZN(n8742) );
  NOR2_X1 U10116 ( .A1(n8754), .A2(n8742), .ZN(n8743) );
  NAND3_X1 U10117 ( .A1(n8744), .A2(n8764), .A3(n8743), .ZN(n8745) );
  OR3_X1 U10118 ( .A1(n8770), .A2(n8746), .A3(n8745), .ZN(n8818) );
  NAND2_X1 U10119 ( .A1(n8747), .A2(n8810), .ZN(n8752) );
  INV_X1 U10120 ( .A(n8748), .ZN(n8750) );
  NAND2_X1 U10121 ( .A1(n8750), .A2(n8749), .ZN(n8751) );
  NAND2_X1 U10122 ( .A1(n8752), .A2(n8751), .ZN(n8753) );
  NOR2_X1 U10123 ( .A1(n8818), .A2(n8753), .ZN(n8776) );
  INV_X1 U10124 ( .A(n8754), .ZN(n8759) );
  OAI21_X1 U10125 ( .B1(n8757), .B2(n8756), .A(n8755), .ZN(n8758) );
  NAND2_X1 U10126 ( .A1(n8759), .A2(n8758), .ZN(n8760) );
  NAND2_X1 U10127 ( .A1(n8761), .A2(n8760), .ZN(n8763) );
  AOI21_X1 U10128 ( .B1(n8764), .B2(n8763), .A(n8762), .ZN(n8766) );
  OAI211_X1 U10129 ( .C1(n8766), .C2(n4541), .A(n9116), .B(n4543), .ZN(n8768)
         );
  NAND2_X1 U10130 ( .A1(n8768), .A2(n8767), .ZN(n8769) );
  OAI22_X1 U10131 ( .A1(n8818), .A2(n8771), .B1(n8770), .B2(n8769), .ZN(n8815)
         );
  NAND2_X1 U10132 ( .A1(n8773), .A2(n8772), .ZN(n8774) );
  NOR2_X1 U10133 ( .A1(n8775), .A2(n8774), .ZN(n8821) );
  OAI21_X1 U10134 ( .B1(n8776), .B2(n8815), .A(n8821), .ZN(n8777) );
  NAND3_X1 U10135 ( .A1(n8778), .A2(n8777), .A3(n8937), .ZN(n8791) );
  NAND2_X1 U10136 ( .A1(n8780), .A2(n8779), .ZN(n8781) );
  NAND2_X1 U10137 ( .A1(n8781), .A2(n8937), .ZN(n8782) );
  AND2_X1 U10138 ( .A1(n8783), .A2(n8782), .ZN(n8784) );
  OR2_X1 U10139 ( .A1(n8800), .A2(n8784), .ZN(n8788) );
  NAND2_X1 U10140 ( .A1(n8786), .A2(n8785), .ZN(n8787) );
  NAND2_X1 U10141 ( .A1(n8788), .A2(n8787), .ZN(n8823) );
  INV_X1 U10142 ( .A(n8823), .ZN(n8789) );
  OAI211_X1 U10143 ( .C1(n8800), .C2(n8791), .A(n8790), .B(n8789), .ZN(n8792)
         );
  NAND2_X1 U10144 ( .A1(n8793), .A2(n8792), .ZN(n8795) );
  INV_X1 U10145 ( .A(n8794), .ZN(n8826) );
  NAND3_X1 U10146 ( .A1(n8795), .A2(n5621), .A3(n8826), .ZN(n8796) );
  NAND3_X1 U10147 ( .A1(n8799), .A2(n9123), .A3(n8796), .ZN(n8798) );
  OAI211_X1 U10148 ( .C1(n8799), .C2(n9123), .A(n8798), .B(n8797), .ZN(n8836)
         );
  INV_X1 U10149 ( .A(n8800), .ZN(n8825) );
  AOI21_X1 U10150 ( .B1(n8849), .B2(n8802), .A(n8801), .ZN(n8807) );
  INV_X1 U10151 ( .A(n8803), .ZN(n8805) );
  AOI211_X1 U10152 ( .C1(n8807), .C2(n8806), .A(n8805), .B(n8804), .ZN(n8808)
         );
  AOI21_X1 U10153 ( .B1(n8809), .B2(n5655), .A(n8808), .ZN(n8812) );
  OAI21_X1 U10154 ( .B1(n8812), .B2(n8811), .A(n8810), .ZN(n8814) );
  NAND2_X1 U10155 ( .A1(n8814), .A2(n8813), .ZN(n8817) );
  INV_X1 U10156 ( .A(n8815), .ZN(n8816) );
  OAI21_X1 U10157 ( .B1(n8818), .B2(n8817), .A(n8816), .ZN(n8820) );
  AOI211_X1 U10158 ( .C1(n8821), .C2(n8820), .A(n8819), .B(n5698), .ZN(n8824)
         );
  AOI211_X1 U10159 ( .C1(n8825), .C2(n8824), .A(n8823), .B(n8822), .ZN(n8828)
         );
  OAI21_X1 U10160 ( .B1(n8828), .B2(n8827), .A(n8826), .ZN(n8831) );
  AOI21_X1 U10161 ( .B1(n8831), .B2(n8830), .A(n8829), .ZN(n8835) );
  INV_X1 U10162 ( .A(n8831), .ZN(n8833) );
  NAND2_X1 U10163 ( .A1(n8833), .A2(n8832), .ZN(n8834) );
  OAI211_X1 U10164 ( .C1(n8837), .C2(n8836), .A(n8835), .B(n8834), .ZN(n8838)
         );
  OAI21_X1 U10165 ( .B1(n8840), .B2(n8839), .A(n8838), .ZN(P1_U3240) );
  MUX2_X1 U10166 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n8841), .S(n9462), .Z(
        P1_U3585) );
  MUX2_X1 U10167 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n9175), .S(n9462), .Z(
        P1_U3584) );
  MUX2_X1 U10168 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n8965), .S(n9462), .Z(
        P1_U3583) );
  MUX2_X1 U10169 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9176), .S(n9462), .Z(
        P1_U3582) );
  MUX2_X1 U10170 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n8999), .S(n9462), .Z(
        P1_U3581) );
  MUX2_X1 U10171 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9013), .S(n9462), .Z(
        P1_U3580) );
  MUX2_X1 U10172 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9023), .S(n9462), .Z(
        P1_U3579) );
  MUX2_X1 U10173 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9039), .S(n9462), .Z(
        P1_U3578) );
  MUX2_X1 U10174 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9218), .S(n9462), .Z(
        P1_U3577) );
  MUX2_X1 U10175 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9038), .S(n9462), .Z(
        P1_U3576) );
  MUX2_X1 U10176 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9232), .S(n9462), .Z(
        P1_U3575) );
  MUX2_X1 U10177 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9242), .S(n9462), .Z(
        P1_U3574) );
  MUX2_X1 U10178 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9233), .S(n9462), .Z(
        P1_U3573) );
  MUX2_X1 U10179 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9256), .S(P1_U4006), .Z(
        P1_U3572) );
  MUX2_X1 U10180 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9265), .S(P1_U4006), .Z(
        P1_U3571) );
  MUX2_X1 U10181 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9255), .S(P1_U4006), .Z(
        P1_U3570) );
  MUX2_X1 U10182 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n9266), .S(P1_U4006), .Z(
        P1_U3569) );
  MUX2_X1 U10183 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n8842), .S(P1_U4006), .Z(
        P1_U3568) );
  MUX2_X1 U10184 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n8843), .S(P1_U4006), .Z(
        P1_U3567) );
  MUX2_X1 U10185 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n8844), .S(P1_U4006), .Z(
        P1_U3566) );
  MUX2_X1 U10186 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n9548), .S(P1_U4006), .Z(
        P1_U3565) );
  MUX2_X1 U10187 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n8845), .S(n9462), .Z(
        P1_U3564) );
  MUX2_X1 U10188 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9547), .S(n9462), .Z(
        P1_U3563) );
  MUX2_X1 U10189 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n9601), .S(n9462), .Z(
        P1_U3562) );
  MUX2_X1 U10190 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n8846), .S(P1_U4006), .Z(
        P1_U3561) );
  MUX2_X1 U10191 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n9602), .S(n9462), .Z(
        P1_U3560) );
  MUX2_X1 U10192 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n8847), .S(n9462), .Z(
        P1_U3559) );
  MUX2_X1 U10193 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n8848), .S(n9462), .Z(
        P1_U3558) );
  MUX2_X1 U10194 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n5655), .S(n9462), .Z(
        P1_U3557) );
  MUX2_X1 U10195 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n8849), .S(n9462), .Z(
        P1_U3556) );
  INV_X1 U10196 ( .A(n8850), .ZN(n8852) );
  AOI21_X1 U10197 ( .B1(n9514), .B2(n8852), .A(n8851), .ZN(n8862) );
  NAND2_X1 U10198 ( .A1(n9539), .A2(P1_ADDR_REG_3__SCAN_IN), .ZN(n8861) );
  OAI211_X1 U10199 ( .C1(n8855), .C2(n8854), .A(n9540), .B(n8853), .ZN(n8860)
         );
  OAI211_X1 U10200 ( .C1(n8858), .C2(n8857), .A(n9530), .B(n8856), .ZN(n8859)
         );
  NAND4_X1 U10201 ( .A1(n8862), .A2(n8861), .A3(n8860), .A4(n8859), .ZN(
        P1_U3244) );
  INV_X1 U10202 ( .A(n8863), .ZN(n8865) );
  AOI21_X1 U10203 ( .B1(n9514), .B2(n8865), .A(n8864), .ZN(n8877) );
  NAND2_X1 U10204 ( .A1(n9539), .A2(P1_ADDR_REG_5__SCAN_IN), .ZN(n8876) );
  OAI211_X1 U10205 ( .C1(n8868), .C2(n8867), .A(n9540), .B(n8866), .ZN(n8875)
         );
  INV_X1 U10206 ( .A(n8869), .ZN(n8873) );
  NOR3_X1 U10207 ( .A1(n9484), .A2(n8871), .A3(n8870), .ZN(n8872) );
  OAI21_X1 U10208 ( .B1(n8873), .B2(n8872), .A(n9530), .ZN(n8874) );
  NAND4_X1 U10209 ( .A1(n8877), .A2(n8876), .A3(n8875), .A4(n8874), .ZN(
        P1_U3246) );
  INV_X1 U10210 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n8891) );
  XNOR2_X1 U10211 ( .A(n8897), .B(P1_REG2_REG_17__SCAN_IN), .ZN(n8879) );
  NOR2_X1 U10212 ( .A1(n8880), .A2(n8879), .ZN(n8892) );
  AOI211_X1 U10213 ( .C1(n8880), .C2(n8879), .A(n8892), .B(n9503), .ZN(n8889)
         );
  AOI21_X1 U10214 ( .B1(n8882), .B2(P1_REG1_REG_16__SCAN_IN), .A(n8881), .ZN(
        n8884) );
  XNOR2_X1 U10215 ( .A(n8897), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n8883) );
  NOR2_X1 U10216 ( .A1(n8884), .A2(n8883), .ZN(n8896) );
  AOI211_X1 U10217 ( .C1(n8884), .C2(n8883), .A(n8896), .B(n9490), .ZN(n8888)
         );
  INV_X1 U10218 ( .A(n8897), .ZN(n8886) );
  NAND2_X1 U10219 ( .A1(P1_REG3_REG_17__SCAN_IN), .A2(P1_U3084), .ZN(n8885) );
  OAI21_X1 U10220 ( .B1(n9533), .B2(n8886), .A(n8885), .ZN(n8887) );
  NOR3_X1 U10221 ( .A1(n8889), .A2(n8888), .A3(n8887), .ZN(n8890) );
  OAI21_X1 U10222 ( .B1(n9525), .B2(n8891), .A(n8890), .ZN(P1_U3258) );
  OR2_X1 U10223 ( .A1(n8898), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n8894) );
  NAND2_X1 U10224 ( .A1(P1_REG2_REG_18__SCAN_IN), .A2(n8898), .ZN(n8893) );
  NAND2_X1 U10225 ( .A1(n8894), .A2(n8893), .ZN(n9528) );
  NOR2_X1 U10226 ( .A1(n9527), .A2(n9528), .ZN(n9526) );
  XNOR2_X1 U10227 ( .A(P1_REG2_REG_19__SCAN_IN), .B(n8895), .ZN(n8903) );
  INV_X1 U10228 ( .A(n8903), .ZN(n8901) );
  AOI22_X1 U10229 ( .A1(P1_REG1_REG_18__SCAN_IN), .A2(n8898), .B1(n9534), .B2(
        n9851), .ZN(n9538) );
  AOI21_X1 U10230 ( .B1(n8897), .B2(P1_REG1_REG_17__SCAN_IN), .A(n8896), .ZN(
        n9537) );
  NAND2_X1 U10231 ( .A1(n9538), .A2(n9537), .ZN(n9536) );
  OAI21_X1 U10232 ( .B1(P1_REG1_REG_18__SCAN_IN), .B2(n8898), .A(n9536), .ZN(
        n8899) );
  XNOR2_X1 U10233 ( .A(n8899), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n8902) );
  OAI21_X1 U10234 ( .B1(n8902), .B2(n9490), .A(n9533), .ZN(n8900) );
  AOI21_X1 U10235 ( .B1(n8901), .B2(n9530), .A(n8900), .ZN(n8905) );
  AOI22_X1 U10236 ( .A1(n8903), .A2(n9530), .B1(n9540), .B2(n8902), .ZN(n8904)
         );
  MUX2_X1 U10237 ( .A(n8905), .B(n8904), .S(n9123), .Z(n8907) );
  NAND2_X1 U10238 ( .A1(P1_REG3_REG_19__SCAN_IN), .A2(P1_U3084), .ZN(n8906) );
  OAI211_X1 U10239 ( .C1(n4664), .C2(n9525), .A(n8907), .B(n8906), .ZN(
        P1_U3260) );
  NOR2_X1 U10240 ( .A1(n8916), .A2(n8915), .ZN(n8909) );
  XNOR2_X1 U10241 ( .A(n8909), .B(n8908), .ZN(n8910) );
  NAND2_X1 U10242 ( .A1(n8910), .A2(n9559), .ZN(n9167) );
  NAND2_X1 U10243 ( .A1(n8912), .A2(n8911), .ZN(n9170) );
  NOR2_X1 U10244 ( .A1(n9575), .A2(n9170), .ZN(n8918) );
  NOR2_X1 U10245 ( .A1(n9284), .A2(n9060), .ZN(n8913) );
  AOI211_X1 U10246 ( .C1(n9575), .C2(P1_REG2_REG_31__SCAN_IN), .A(n8918), .B(
        n8913), .ZN(n8914) );
  OAI21_X1 U10247 ( .B1(n9162), .B2(n9167), .A(n8914), .ZN(P1_U3261) );
  XNOR2_X1 U10248 ( .A(n8916), .B(n8915), .ZN(n8917) );
  NOR2_X1 U10249 ( .A1(n8917), .A2(n9158), .ZN(n9172) );
  NAND2_X1 U10250 ( .A1(n9172), .A2(n9562), .ZN(n8920) );
  AOI21_X1 U10251 ( .B1(n9575), .B2(P1_REG2_REG_30__SCAN_IN), .A(n8918), .ZN(
        n8919) );
  OAI211_X1 U10252 ( .C1(n9287), .C2(n9060), .A(n8920), .B(n8919), .ZN(
        P1_U3262) );
  INV_X1 U10253 ( .A(n8921), .ZN(n8931) );
  OAI21_X1 U10254 ( .B1(n8923), .B2(n9567), .A(n8922), .ZN(n8929) );
  NOR2_X1 U10255 ( .A1(n8924), .A2(n9162), .ZN(n8928) );
  AOI22_X1 U10256 ( .A1(n9136), .A2(n8965), .B1(n9575), .B2(
        P1_REG2_REG_29__SCAN_IN), .ZN(n8925) );
  OAI21_X1 U10257 ( .B1(n8926), .B2(n9060), .A(n8925), .ZN(n8927) );
  AOI211_X1 U10258 ( .C1(n8929), .C2(n9572), .A(n8928), .B(n8927), .ZN(n8930)
         );
  OAI21_X1 U10259 ( .B1(n8931), .B2(n9079), .A(n8930), .ZN(P1_U3355) );
  INV_X1 U10260 ( .A(n9181), .ZN(n8955) );
  NAND2_X1 U10261 ( .A1(n8936), .A2(n8937), .ZN(n8939) );
  NAND2_X1 U10262 ( .A1(n8939), .A2(n8938), .ZN(n8941) );
  NAND2_X1 U10263 ( .A1(n8941), .A2(n8940), .ZN(n9174) );
  INV_X1 U10264 ( .A(n8942), .ZN(n8944) );
  AOI21_X1 U10265 ( .B1(n8957), .B2(n8945), .A(n9158), .ZN(n8943) );
  NAND2_X1 U10266 ( .A1(n8944), .A2(n8943), .ZN(n9177) );
  NOR2_X1 U10267 ( .A1(n9177), .A2(n9162), .ZN(n8952) );
  OAI22_X1 U10268 ( .A1(n9572), .A2(n8947), .B1(n8946), .B2(n9567), .ZN(n8948)
         );
  AOI21_X1 U10269 ( .B1(n9136), .B2(n9176), .A(n8948), .ZN(n8950) );
  NAND2_X1 U10270 ( .A1(n9155), .A2(n9175), .ZN(n8949) );
  OAI211_X1 U10271 ( .C1(n4535), .C2(n9060), .A(n8950), .B(n8949), .ZN(n8951)
         );
  AOI211_X1 U10272 ( .C1(n9174), .C2(n8953), .A(n8952), .B(n8951), .ZN(n8954)
         );
  OAI21_X1 U10273 ( .B1(n8955), .B2(n9079), .A(n8954), .ZN(P1_U3263) );
  XOR2_X1 U10274 ( .A(n8964), .B(n8956), .Z(n9188) );
  INV_X1 U10275 ( .A(n8957), .ZN(n8958) );
  AOI211_X1 U10276 ( .C1(n9186), .C2(n8971), .A(n9158), .B(n8958), .ZN(n9185)
         );
  NOR2_X1 U10277 ( .A1(n4537), .A2(n9060), .ZN(n8962) );
  OAI22_X1 U10278 ( .A1(n9572), .A2(n8960), .B1(n8959), .B2(n9567), .ZN(n8961)
         );
  AOI211_X1 U10279 ( .C1(n9185), .C2(n9562), .A(n8962), .B(n8961), .ZN(n8969)
         );
  OAI211_X1 U10280 ( .C1(n8964), .C2(n8963), .A(n8936), .B(n9550), .ZN(n8967)
         );
  AOI22_X1 U10281 ( .A1(n9603), .A2(n8999), .B1(n8965), .B2(n9600), .ZN(n8966)
         );
  NAND2_X1 U10282 ( .A1(n8967), .A2(n8966), .ZN(n9184) );
  NAND2_X1 U10283 ( .A1(n9184), .A2(n9572), .ZN(n8968) );
  OAI211_X1 U10284 ( .C1(n9188), .C2(n9079), .A(n8969), .B(n8968), .ZN(
        P1_U3264) );
  XOR2_X1 U10285 ( .A(n8979), .B(n8970), .Z(n9191) );
  INV_X1 U10286 ( .A(n9191), .ZN(n8985) );
  INV_X1 U10287 ( .A(n8971), .ZN(n8972) );
  AOI211_X1 U10288 ( .C1(n8973), .C2(n8987), .A(n9158), .B(n8972), .ZN(n9190)
         );
  NOR2_X1 U10289 ( .A1(n9295), .A2(n9060), .ZN(n8977) );
  OAI22_X1 U10290 ( .A1(n9572), .A2(n8975), .B1(n8974), .B2(n9567), .ZN(n8976)
         );
  AOI211_X1 U10291 ( .C1(n9190), .C2(n9562), .A(n8977), .B(n8976), .ZN(n8984)
         );
  OAI211_X1 U10292 ( .C1(n8980), .C2(n8979), .A(n8978), .B(n9550), .ZN(n8982)
         );
  AOI22_X1 U10293 ( .A1(n9603), .A2(n9013), .B1(n9176), .B2(n9600), .ZN(n8981)
         );
  NAND2_X1 U10294 ( .A1(n8982), .A2(n8981), .ZN(n9189) );
  NAND2_X1 U10295 ( .A1(n9189), .A2(n9572), .ZN(n8983) );
  OAI211_X1 U10296 ( .C1(n8985), .C2(n9079), .A(n8984), .B(n8983), .ZN(
        P1_U3265) );
  XNOR2_X1 U10297 ( .A(n8986), .B(n8995), .ZN(n9196) );
  INV_X1 U10298 ( .A(n9196), .ZN(n9004) );
  INV_X1 U10299 ( .A(n9008), .ZN(n8989) );
  INV_X1 U10300 ( .A(n8987), .ZN(n8988) );
  AOI211_X1 U10301 ( .C1(n8990), .C2(n8989), .A(n9158), .B(n8988), .ZN(n9195)
         );
  NOR2_X1 U10302 ( .A1(n9299), .A2(n9060), .ZN(n8994) );
  OAI22_X1 U10303 ( .A1(n9572), .A2(n8992), .B1(n8991), .B2(n9567), .ZN(n8993)
         );
  AOI211_X1 U10304 ( .C1(n9195), .C2(n9562), .A(n8994), .B(n8993), .ZN(n9003)
         );
  OAI21_X1 U10305 ( .B1(n4294), .B2(n8996), .A(n8995), .ZN(n8998) );
  NAND3_X1 U10306 ( .A1(n8998), .A2(n9550), .A3(n8997), .ZN(n9001) );
  AOI22_X1 U10307 ( .A1(n9023), .A2(n9603), .B1(n9600), .B2(n8999), .ZN(n9000)
         );
  NAND2_X1 U10308 ( .A1(n9001), .A2(n9000), .ZN(n9194) );
  NAND2_X1 U10309 ( .A1(n9194), .A2(n9572), .ZN(n9002) );
  OAI211_X1 U10310 ( .C1(n9004), .C2(n9079), .A(n9003), .B(n9002), .ZN(
        P1_U3266) );
  AOI21_X1 U10311 ( .B1(n9007), .B2(n9005), .A(n4294), .ZN(n9207) );
  XOR2_X1 U10312 ( .A(n9007), .B(n9006), .Z(n9199) );
  NAND2_X1 U10313 ( .A1(n9199), .A2(n9563), .ZN(n9018) );
  INV_X1 U10314 ( .A(n9026), .ZN(n9009) );
  AOI211_X1 U10315 ( .C1(n9204), .C2(n9009), .A(n9158), .B(n9008), .ZN(n9202)
         );
  AOI22_X1 U10316 ( .A1(P1_REG2_REG_24__SCAN_IN), .A2(n9575), .B1(n9010), .B2(
        n9552), .ZN(n9011) );
  OAI21_X1 U10317 ( .B1(n9201), .B2(n9157), .A(n9011), .ZN(n9012) );
  AOI21_X1 U10318 ( .B1(n9155), .B2(n9013), .A(n9012), .ZN(n9014) );
  OAI21_X1 U10319 ( .B1(n9015), .B2(n9060), .A(n9014), .ZN(n9016) );
  AOI21_X1 U10320 ( .B1(n9202), .B2(n9562), .A(n9016), .ZN(n9017) );
  OAI211_X1 U10321 ( .C1(n9207), .C2(n9146), .A(n9018), .B(n9017), .ZN(
        P1_U3267) );
  XNOR2_X1 U10322 ( .A(n9019), .B(n9021), .ZN(n9212) );
  AOI22_X1 U10323 ( .A1(n9210), .A2(n9554), .B1(n9575), .B2(
        P1_REG2_REG_23__SCAN_IN), .ZN(n9031) );
  OAI211_X1 U10324 ( .C1(n9022), .C2(n9021), .A(n9020), .B(n9550), .ZN(n9025)
         );
  AOI22_X1 U10325 ( .A1(n9023), .A2(n9600), .B1(n9603), .B2(n9218), .ZN(n9024)
         );
  NAND2_X1 U10326 ( .A1(n9025), .A2(n9024), .ZN(n9208) );
  AOI211_X1 U10327 ( .C1(n9210), .C2(n9042), .A(n9158), .B(n9026), .ZN(n9209)
         );
  INV_X1 U10328 ( .A(n9209), .ZN(n9028) );
  OAI22_X1 U10329 ( .A1(n9028), .A2(n9074), .B1(n9567), .B2(n9027), .ZN(n9029)
         );
  OAI21_X1 U10330 ( .B1(n9208), .B2(n9029), .A(n9572), .ZN(n9030) );
  OAI211_X1 U10331 ( .C1(n9212), .C2(n9079), .A(n9031), .B(n9030), .ZN(
        P1_U3268) );
  XNOR2_X1 U10332 ( .A(n9032), .B(n9034), .ZN(n9217) );
  AOI21_X1 U10333 ( .B1(n9034), .B2(n9033), .A(n9399), .ZN(n9035) );
  OAI211_X1 U10334 ( .C1(n9050), .C2(n9037), .A(n9036), .B(n9035), .ZN(n9041)
         );
  AOI22_X1 U10335 ( .A1(n9039), .A2(n9600), .B1(n9603), .B2(n9038), .ZN(n9040)
         );
  NAND2_X1 U10336 ( .A1(n9041), .A2(n9040), .ZN(n9213) );
  INV_X1 U10337 ( .A(n9215), .ZN(n9047) );
  AOI211_X1 U10338 ( .C1(n9215), .C2(n4290), .A(n9158), .B(n4528), .ZN(n9214)
         );
  NAND2_X1 U10339 ( .A1(n9214), .A2(n9562), .ZN(n9046) );
  INV_X1 U10340 ( .A(n9043), .ZN(n9044) );
  AOI22_X1 U10341 ( .A1(n9575), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n9044), .B2(
        n9552), .ZN(n9045) );
  OAI211_X1 U10342 ( .C1(n9047), .C2(n9060), .A(n9046), .B(n9045), .ZN(n9048)
         );
  AOI21_X1 U10343 ( .B1(n9213), .B2(n9572), .A(n9048), .ZN(n9049) );
  OAI21_X1 U10344 ( .B1(n9217), .B2(n9079), .A(n9049), .ZN(P1_U3269) );
  INV_X1 U10345 ( .A(n9050), .ZN(n9051) );
  AOI21_X1 U10346 ( .B1(n9054), .B2(n9052), .A(n9051), .ZN(n9221) );
  XOR2_X1 U10347 ( .A(n9053), .B(n9054), .Z(n9223) );
  NAND2_X1 U10348 ( .A1(n9223), .A2(n9563), .ZN(n9064) );
  OAI211_X1 U10349 ( .C1(n9070), .C2(n9305), .A(n9559), .B(n4290), .ZN(n9219)
         );
  INV_X1 U10350 ( .A(n9219), .ZN(n9062) );
  OAI22_X1 U10351 ( .A1(n9572), .A2(n9056), .B1(n9055), .B2(n9567), .ZN(n9058)
         );
  NOR2_X1 U10352 ( .A1(n9157), .A2(n9087), .ZN(n9057) );
  AOI211_X1 U10353 ( .C1(n9155), .C2(n9218), .A(n9058), .B(n9057), .ZN(n9059)
         );
  OAI21_X1 U10354 ( .B1(n9305), .B2(n9060), .A(n9059), .ZN(n9061) );
  AOI21_X1 U10355 ( .B1(n9062), .B2(n9562), .A(n9061), .ZN(n9063) );
  OAI211_X1 U10356 ( .C1(n9221), .C2(n9146), .A(n9064), .B(n9063), .ZN(
        P1_U3270) );
  XOR2_X1 U10357 ( .A(n9065), .B(n9066), .Z(n9230) );
  AOI22_X1 U10358 ( .A1(n9228), .A2(n9554), .B1(P1_REG2_REG_20__SCAN_IN), .B2(
        n9575), .ZN(n9078) );
  XNOR2_X1 U10359 ( .A(n9067), .B(n9066), .ZN(n9068) );
  OAI222_X1 U10360 ( .A1(n9440), .A2(n9069), .B1(n9438), .B2(n9104), .C1(n9068), .C2(n9399), .ZN(n9226) );
  INV_X1 U10361 ( .A(n9089), .ZN(n9071) );
  AOI211_X1 U10362 ( .C1(n9228), .C2(n9071), .A(n9158), .B(n9070), .ZN(n9227)
         );
  INV_X1 U10363 ( .A(n9227), .ZN(n9075) );
  INV_X1 U10364 ( .A(n9072), .ZN(n9073) );
  OAI22_X1 U10365 ( .A1(n9075), .A2(n9074), .B1(n9567), .B2(n9073), .ZN(n9076)
         );
  OAI21_X1 U10366 ( .B1(n9226), .B2(n9076), .A(n9572), .ZN(n9077) );
  OAI211_X1 U10367 ( .C1(n9230), .C2(n9079), .A(n9078), .B(n9077), .ZN(
        P1_U3271) );
  XOR2_X1 U10368 ( .A(n9082), .B(n9080), .Z(n9236) );
  XNOR2_X1 U10369 ( .A(n9081), .B(n9082), .ZN(n9238) );
  NAND2_X1 U10370 ( .A1(n9238), .A2(n9563), .ZN(n9094) );
  INV_X1 U10371 ( .A(n9155), .ZN(n9138) );
  OAI22_X1 U10372 ( .A1(n9572), .A2(n9084), .B1(n9083), .B2(n9567), .ZN(n9085)
         );
  AOI21_X1 U10373 ( .B1(n9136), .B2(n9233), .A(n9085), .ZN(n9086) );
  OAI21_X1 U10374 ( .B1(n9087), .B2(n9138), .A(n9086), .ZN(n9092) );
  NAND2_X1 U10375 ( .A1(n9105), .A2(n9231), .ZN(n9088) );
  NAND2_X1 U10376 ( .A1(n9088), .A2(n9559), .ZN(n9090) );
  OR2_X1 U10377 ( .A1(n9090), .A2(n9089), .ZN(n9234) );
  NOR2_X1 U10378 ( .A1(n9234), .A2(n9162), .ZN(n9091) );
  AOI211_X1 U10379 ( .C1(n9554), .C2(n9231), .A(n9092), .B(n9091), .ZN(n9093)
         );
  OAI211_X1 U10380 ( .C1(n9236), .C2(n9146), .A(n9094), .B(n9093), .ZN(
        P1_U3272) );
  INV_X1 U10381 ( .A(n9095), .ZN(n9096) );
  AOI21_X1 U10382 ( .B1(n9098), .B2(n9097), .A(n9096), .ZN(n9245) );
  XNOR2_X1 U10383 ( .A(n9099), .B(n4580), .ZN(n9247) );
  NAND2_X1 U10384 ( .A1(n9247), .A2(n9563), .ZN(n9110) );
  OAI22_X1 U10385 ( .A1(n9572), .A2(n9101), .B1(n9100), .B2(n9567), .ZN(n9102)
         );
  AOI21_X1 U10386 ( .B1(n9136), .B2(n9256), .A(n9102), .ZN(n9103) );
  OAI21_X1 U10387 ( .B1(n9104), .B2(n9138), .A(n9103), .ZN(n9108) );
  AOI21_X1 U10388 ( .B1(n9112), .B2(n9241), .A(n9158), .ZN(n9106) );
  NAND2_X1 U10389 ( .A1(n9106), .A2(n9105), .ZN(n9243) );
  NOR2_X1 U10390 ( .A1(n9243), .A2(n9162), .ZN(n9107) );
  AOI211_X1 U10391 ( .C1(n9554), .C2(n9241), .A(n9108), .B(n9107), .ZN(n9109)
         );
  OAI211_X1 U10392 ( .C1(n9245), .C2(n9146), .A(n9110), .B(n9109), .ZN(
        P1_U3273) );
  INV_X1 U10393 ( .A(n9111), .ZN(n9141) );
  INV_X1 U10394 ( .A(n9112), .ZN(n9113) );
  AOI211_X1 U10395 ( .C1(n9126), .C2(n9141), .A(n9158), .B(n9113), .ZN(n9250)
         );
  NOR2_X1 U10396 ( .A1(n9567), .A2(n9114), .ZN(n9122) );
  NAND3_X1 U10397 ( .A1(n9117), .A2(n9116), .A3(n9115), .ZN(n9118) );
  NAND3_X1 U10398 ( .A1(n9119), .A2(n9550), .A3(n9118), .ZN(n9121) );
  AOI22_X1 U10399 ( .A1(n9603), .A2(n9265), .B1(n9233), .B2(n9600), .ZN(n9120)
         );
  NAND2_X1 U10400 ( .A1(n9121), .A2(n9120), .ZN(n9249) );
  AOI211_X1 U10401 ( .C1(n9250), .C2(n9123), .A(n9122), .B(n9249), .ZN(n9129)
         );
  XNOR2_X1 U10402 ( .A(n9124), .B(n9125), .ZN(n9251) );
  NAND2_X1 U10403 ( .A1(n9251), .A2(n9563), .ZN(n9128) );
  AOI22_X1 U10404 ( .A1(n9126), .A2(n9554), .B1(P1_REG2_REG_17__SCAN_IN), .B2(
        n9575), .ZN(n9127) );
  OAI211_X1 U10405 ( .C1(n9575), .C2(n9129), .A(n9128), .B(n9127), .ZN(
        P1_U3274) );
  XNOR2_X1 U10406 ( .A(n9130), .B(n9132), .ZN(n9259) );
  XOR2_X1 U10407 ( .A(n9131), .B(n9132), .Z(n9261) );
  NAND2_X1 U10408 ( .A1(n9261), .A2(n9563), .ZN(n9145) );
  OAI22_X1 U10409 ( .A1(n9572), .A2(n9134), .B1(n9133), .B2(n9567), .ZN(n9135)
         );
  AOI21_X1 U10410 ( .B1(n9136), .B2(n9255), .A(n9135), .ZN(n9137) );
  OAI21_X1 U10411 ( .B1(n9139), .B2(n9138), .A(n9137), .ZN(n9143) );
  AOI21_X1 U10412 ( .B1(n9160), .B2(n9254), .A(n9158), .ZN(n9140) );
  NAND2_X1 U10413 ( .A1(n9141), .A2(n9140), .ZN(n9257) );
  NOR2_X1 U10414 ( .A1(n9257), .A2(n9162), .ZN(n9142) );
  AOI211_X1 U10415 ( .C1(n9554), .C2(n9254), .A(n9143), .B(n9142), .ZN(n9144)
         );
  OAI211_X1 U10416 ( .C1(n9259), .C2(n9146), .A(n9145), .B(n9144), .ZN(
        P1_U3275) );
  XNOR2_X1 U10417 ( .A(n9147), .B(n9150), .ZN(n9148) );
  NAND2_X1 U10418 ( .A1(n9148), .A2(n9550), .ZN(n9271) );
  XOR2_X1 U10419 ( .A(n9149), .B(n9150), .Z(n9274) );
  INV_X1 U10420 ( .A(n9274), .ZN(n9151) );
  NAND2_X1 U10421 ( .A1(n9151), .A2(n9563), .ZN(n9166) );
  OAI22_X1 U10422 ( .A1(n9572), .A2(n9153), .B1(n9152), .B2(n9567), .ZN(n9154)
         );
  AOI21_X1 U10423 ( .B1(n9155), .B2(n9265), .A(n9154), .ZN(n9156) );
  OAI21_X1 U10424 ( .B1(n9402), .B2(n9157), .A(n9156), .ZN(n9164) );
  AOI21_X1 U10425 ( .B1(n9159), .B2(n9264), .A(n9158), .ZN(n9161) );
  NAND2_X1 U10426 ( .A1(n9161), .A2(n9160), .ZN(n9268) );
  NOR2_X1 U10427 ( .A1(n9268), .A2(n9162), .ZN(n9163) );
  AOI211_X1 U10428 ( .C1(n9554), .C2(n9264), .A(n9164), .B(n9163), .ZN(n9165)
         );
  OAI211_X1 U10429 ( .C1(n9575), .C2(n9271), .A(n9166), .B(n9165), .ZN(
        P1_U3276) );
  OAI21_X1 U10430 ( .B1(n9284), .B2(n9280), .A(n9169), .ZN(P1_U3554) );
  INV_X1 U10431 ( .A(n9170), .ZN(n9171) );
  NOR2_X1 U10432 ( .A1(n9172), .A2(n9171), .ZN(n9285) );
  MUX2_X1 U10433 ( .A(n5740), .B(n9285), .S(n4270), .Z(n9173) );
  OAI21_X1 U10434 ( .B1(n9287), .B2(n9280), .A(n9173), .ZN(P1_U3553) );
  INV_X1 U10435 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n9182) );
  NAND2_X1 U10436 ( .A1(n9174), .A2(n9550), .ZN(n9179) );
  AOI22_X1 U10437 ( .A1(n9603), .A2(n9176), .B1(n9175), .B2(n9600), .ZN(n9178)
         );
  NAND3_X1 U10438 ( .A1(n9179), .A2(n9178), .A3(n9177), .ZN(n9180) );
  AOI21_X1 U10439 ( .B1(n9181), .B2(n9615), .A(n9180), .ZN(n9288) );
  OAI21_X1 U10440 ( .B1(n4535), .B2(n9280), .A(n9183), .ZN(P1_U3551) );
  AOI211_X1 U10441 ( .C1(n9452), .C2(n9186), .A(n9185), .B(n9184), .ZN(n9187)
         );
  OAI21_X1 U10442 ( .B1(n9188), .B2(n9273), .A(n9187), .ZN(n9291) );
  MUX2_X1 U10443 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9291), .S(n4270), .Z(
        P1_U3550) );
  AOI211_X1 U10444 ( .C1(n9191), .C2(n9615), .A(n9190), .B(n9189), .ZN(n9292)
         );
  MUX2_X1 U10445 ( .A(n9192), .B(n9292), .S(n4270), .Z(n9193) );
  OAI21_X1 U10446 ( .B1(n9295), .B2(n9280), .A(n9193), .ZN(P1_U3549) );
  INV_X1 U10447 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n9197) );
  AOI211_X1 U10448 ( .C1(n9196), .C2(n9615), .A(n9195), .B(n9194), .ZN(n9296)
         );
  MUX2_X1 U10449 ( .A(n9197), .B(n9296), .S(n4270), .Z(n9198) );
  OAI21_X1 U10450 ( .B1(n9299), .B2(n9280), .A(n9198), .ZN(P1_U3548) );
  NAND2_X1 U10451 ( .A1(n9199), .A2(n9615), .ZN(n9206) );
  OAI22_X1 U10452 ( .A1(n9201), .A2(n9438), .B1(n9200), .B2(n9440), .ZN(n9203)
         );
  AOI211_X1 U10453 ( .C1(n9452), .C2(n9204), .A(n9203), .B(n9202), .ZN(n9205)
         );
  OAI211_X1 U10454 ( .C1(n9399), .C2(n9207), .A(n9206), .B(n9205), .ZN(n9300)
         );
  MUX2_X1 U10455 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9300), .S(n4270), .Z(
        P1_U3547) );
  AOI211_X1 U10456 ( .C1(n9452), .C2(n9210), .A(n9209), .B(n9208), .ZN(n9211)
         );
  OAI21_X1 U10457 ( .B1(n9212), .B2(n9273), .A(n9211), .ZN(n9301) );
  MUX2_X1 U10458 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9301), .S(n4270), .Z(
        P1_U3546) );
  AOI211_X1 U10459 ( .C1(n9452), .C2(n9215), .A(n9214), .B(n9213), .ZN(n9216)
         );
  OAI21_X1 U10460 ( .B1(n9217), .B2(n9273), .A(n9216), .ZN(n9302) );
  MUX2_X1 U10461 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9302), .S(n4270), .Z(
        P1_U3545) );
  INV_X1 U10462 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n9224) );
  AOI22_X1 U10463 ( .A1(n9218), .A2(n9600), .B1(n9603), .B2(n9232), .ZN(n9220)
         );
  OAI211_X1 U10464 ( .C1(n9221), .C2(n9399), .A(n9220), .B(n9219), .ZN(n9222)
         );
  AOI21_X1 U10465 ( .B1(n9223), .B2(n9615), .A(n9222), .ZN(n9303) );
  MUX2_X1 U10466 ( .A(n9224), .B(n9303), .S(n4270), .Z(n9225) );
  OAI21_X1 U10467 ( .B1(n9305), .B2(n9280), .A(n9225), .ZN(P1_U3544) );
  AOI211_X1 U10468 ( .C1(n9452), .C2(n9228), .A(n9227), .B(n9226), .ZN(n9229)
         );
  OAI21_X1 U10469 ( .B1(n9230), .B2(n9273), .A(n9229), .ZN(n9306) );
  MUX2_X1 U10470 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9306), .S(n4270), .Z(
        P1_U3543) );
  INV_X1 U10471 ( .A(n9231), .ZN(n9310) );
  AOI22_X1 U10472 ( .A1(n9603), .A2(n9233), .B1(n9232), .B2(n9600), .ZN(n9235)
         );
  OAI211_X1 U10473 ( .C1(n9236), .C2(n9399), .A(n9235), .B(n9234), .ZN(n9237)
         );
  AOI21_X1 U10474 ( .B1(n9238), .B2(n9615), .A(n9237), .ZN(n9307) );
  MUX2_X1 U10475 ( .A(n9239), .B(n9307), .S(n4270), .Z(n9240) );
  OAI21_X1 U10476 ( .B1(n9310), .B2(n9280), .A(n9240), .ZN(P1_U3542) );
  INV_X1 U10477 ( .A(n9241), .ZN(n9314) );
  AOI22_X1 U10478 ( .A1(n9603), .A2(n9256), .B1(n9242), .B2(n9600), .ZN(n9244)
         );
  OAI211_X1 U10479 ( .C1(n9245), .C2(n9399), .A(n9244), .B(n9243), .ZN(n9246)
         );
  AOI21_X1 U10480 ( .B1(n9247), .B2(n9615), .A(n9246), .ZN(n9311) );
  MUX2_X1 U10481 ( .A(n9851), .B(n9311), .S(n4270), .Z(n9248) );
  OAI21_X1 U10482 ( .B1(n9314), .B2(n9280), .A(n9248), .ZN(P1_U3541) );
  AOI211_X1 U10483 ( .C1(n9251), .C2(n9615), .A(n9250), .B(n9249), .ZN(n9315)
         );
  MUX2_X1 U10484 ( .A(n9252), .B(n9315), .S(n4270), .Z(n9253) );
  OAI21_X1 U10485 ( .B1(n9318), .B2(n9280), .A(n9253), .ZN(P1_U3540) );
  INV_X1 U10486 ( .A(n9254), .ZN(n9322) );
  INV_X1 U10487 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9262) );
  AOI22_X1 U10488 ( .A1(n9600), .A2(n9256), .B1(n9255), .B2(n9603), .ZN(n9258)
         );
  OAI211_X1 U10489 ( .C1(n9259), .C2(n9399), .A(n9258), .B(n9257), .ZN(n9260)
         );
  AOI21_X1 U10490 ( .B1(n9261), .B2(n9615), .A(n9260), .ZN(n9319) );
  MUX2_X1 U10491 ( .A(n9262), .B(n9319), .S(n4270), .Z(n9263) );
  OAI21_X1 U10492 ( .B1(n9322), .B2(n9280), .A(n9263), .ZN(P1_U3539) );
  INV_X1 U10493 ( .A(n9264), .ZN(n9269) );
  AOI22_X1 U10494 ( .A1(n9603), .A2(n9266), .B1(n9265), .B2(n9600), .ZN(n9267)
         );
  OAI211_X1 U10495 ( .C1(n9269), .C2(n9612), .A(n9268), .B(n9267), .ZN(n9270)
         );
  INV_X1 U10496 ( .A(n9270), .ZN(n9272) );
  OAI211_X1 U10497 ( .C1(n9274), .C2(n9273), .A(n9272), .B(n9271), .ZN(n9323)
         );
  MUX2_X1 U10498 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n9323), .S(n4270), .Z(
        P1_U3538) );
  AOI211_X1 U10499 ( .C1(n9277), .C2(n9615), .A(n9276), .B(n9275), .ZN(n9324)
         );
  MUX2_X1 U10500 ( .A(n9278), .B(n9324), .S(n4270), .Z(n9279) );
  OAI21_X1 U10501 ( .B1(n9327), .B2(n9280), .A(n9279), .ZN(P1_U3537) );
  OAI21_X1 U10502 ( .B1(n9284), .B2(n9326), .A(n9283), .ZN(P1_U3522) );
  MUX2_X1 U10503 ( .A(n5737), .B(n9285), .S(n9619), .Z(n9286) );
  OAI21_X1 U10504 ( .B1(n9287), .B2(n9326), .A(n9286), .ZN(P1_U3521) );
  MUX2_X1 U10505 ( .A(n9289), .B(n9288), .S(n9619), .Z(n9290) );
  MUX2_X1 U10506 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9291), .S(n9619), .Z(
        P1_U3518) );
  INV_X1 U10507 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n9293) );
  MUX2_X1 U10508 ( .A(n9293), .B(n9292), .S(n9619), .Z(n9294) );
  OAI21_X1 U10509 ( .B1(n9295), .B2(n9326), .A(n9294), .ZN(P1_U3517) );
  MUX2_X1 U10510 ( .A(n9297), .B(n9296), .S(n9619), .Z(n9298) );
  OAI21_X1 U10511 ( .B1(n9299), .B2(n9326), .A(n9298), .ZN(P1_U3516) );
  MUX2_X1 U10512 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9300), .S(n9619), .Z(
        P1_U3515) );
  MUX2_X1 U10513 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9301), .S(n9619), .Z(
        P1_U3514) );
  MUX2_X1 U10514 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9302), .S(n9619), .Z(
        P1_U3513) );
  MUX2_X1 U10515 ( .A(n9836), .B(n9303), .S(n9619), .Z(n9304) );
  OAI21_X1 U10516 ( .B1(n9305), .B2(n9326), .A(n9304), .ZN(P1_U3512) );
  MUX2_X1 U10517 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9306), .S(n9619), .Z(
        P1_U3511) );
  MUX2_X1 U10518 ( .A(n9308), .B(n9307), .S(n9619), .Z(n9309) );
  OAI21_X1 U10519 ( .B1(n9310), .B2(n9326), .A(n9309), .ZN(P1_U3510) );
  INV_X1 U10520 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n9312) );
  MUX2_X1 U10521 ( .A(n9312), .B(n9311), .S(n9619), .Z(n9313) );
  OAI21_X1 U10522 ( .B1(n9314), .B2(n9326), .A(n9313), .ZN(P1_U3508) );
  MUX2_X1 U10523 ( .A(n9316), .B(n9315), .S(n9619), .Z(n9317) );
  OAI21_X1 U10524 ( .B1(n9318), .B2(n9326), .A(n9317), .ZN(P1_U3505) );
  MUX2_X1 U10525 ( .A(n9320), .B(n9319), .S(n9619), .Z(n9321) );
  OAI21_X1 U10526 ( .B1(n9322), .B2(n9326), .A(n9321), .ZN(P1_U3502) );
  MUX2_X1 U10527 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n9323), .S(n9619), .Z(
        P1_U3499) );
  MUX2_X1 U10528 ( .A(n9884), .B(n9324), .S(n9619), .Z(n9325) );
  OAI21_X1 U10529 ( .B1(n9327), .B2(n9326), .A(n9325), .ZN(P1_U3496) );
  MUX2_X1 U10530 ( .A(P1_D_REG_0__SCAN_IN), .B(n9328), .S(n9577), .Z(P1_U3440)
         );
  NOR4_X1 U10531 ( .A1(n9329), .A2(P1_IR_REG_30__SCAN_IN), .A3(n9330), .A4(
        P1_U3084), .ZN(n9331) );
  AOI21_X1 U10532 ( .B1(n9332), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9331), .ZN(
        n9333) );
  OAI21_X1 U10533 ( .B1(n9334), .B2(n9343), .A(n9333), .ZN(P1_U3322) );
  OAI222_X1 U10534 ( .A1(n9340), .A2(n9336), .B1(n9343), .B2(n9335), .C1(n5637), .C2(P1_U3084), .ZN(P1_U3325) );
  OAI222_X1 U10535 ( .A1(n9340), .A2(n9339), .B1(n9343), .B2(n9338), .C1(n9337), .C2(P1_U3084), .ZN(P1_U3326) );
  OAI222_X1 U10536 ( .A1(P1_U3084), .A2(n9344), .B1(n9343), .B2(n9342), .C1(
        n9341), .C2(n9340), .ZN(P1_U3327) );
  INV_X1 U10537 ( .A(n9345), .ZN(n9346) );
  MUX2_X1 U10538 ( .A(n9346), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3353) );
  AOI22_X1 U10539 ( .A1(n9633), .A2(P2_ADDR_REG_1__SCAN_IN), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(n4264), .ZN(n9357) );
  NAND2_X1 U10540 ( .A1(n9638), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n9349) );
  AOI211_X1 U10541 ( .C1(n9349), .C2(n9348), .A(n9347), .B(n9629), .ZN(n9350)
         );
  AOI21_X1 U10542 ( .B1(n9363), .B2(n9351), .A(n9350), .ZN(n9356) );
  AND2_X1 U10543 ( .A1(n9638), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n9354) );
  OAI211_X1 U10544 ( .C1(n9354), .C2(n9353), .A(n9632), .B(n9352), .ZN(n9355)
         );
  NAND3_X1 U10545 ( .A1(n9357), .A2(n9356), .A3(n9355), .ZN(P2_U3246) );
  AOI22_X1 U10546 ( .A1(n9633), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3152), .ZN(n9369) );
  AOI211_X1 U10547 ( .C1(n9360), .C2(n9359), .A(n9358), .B(n9629), .ZN(n9361)
         );
  AOI21_X1 U10548 ( .B1(n9363), .B2(n9362), .A(n9361), .ZN(n9368) );
  OAI211_X1 U10549 ( .C1(n9366), .C2(n9365), .A(n9632), .B(n9364), .ZN(n9367)
         );
  NAND3_X1 U10550 ( .A1(n9369), .A2(n9368), .A3(n9367), .ZN(P2_U3247) );
  OAI22_X1 U10551 ( .A1(n9370), .A2(n9438), .B1(n9439), .B2(n9440), .ZN(n9372)
         );
  AOI211_X1 U10552 ( .C1(n9452), .C2(n9373), .A(n9372), .B(n9371), .ZN(n9375)
         );
  OAI211_X1 U10553 ( .C1(n9376), .C2(n9582), .A(n9375), .B(n9374), .ZN(n9377)
         );
  AOI21_X1 U10554 ( .B1(n9587), .B2(n9378), .A(n9377), .ZN(n9379) );
  AOI22_X1 U10555 ( .A1(n9619), .A2(n9379), .B1(n5166), .B2(n9617), .ZN(
        P1_U3484) );
  AOI22_X1 U10556 ( .A1(n4270), .A2(n9379), .B1(n6422), .B2(n9625), .ZN(
        P1_U3533) );
  OAI22_X1 U10557 ( .A1(n9381), .A2(n9728), .B1(n9380), .B2(n9727), .ZN(n9383)
         );
  AOI211_X1 U10558 ( .C1(n9733), .C2(n9384), .A(n9383), .B(n9382), .ZN(n9393)
         );
  AOI22_X1 U10559 ( .A1(n9752), .A2(n9393), .B1(n9385), .B2(n9750), .ZN(
        P2_U3535) );
  OAI22_X1 U10560 ( .A1(n9387), .A2(n9728), .B1(n9386), .B2(n9727), .ZN(n9389)
         );
  AOI211_X1 U10561 ( .C1(n9733), .C2(n9390), .A(n9389), .B(n9388), .ZN(n9394)
         );
  AOI22_X1 U10562 ( .A1(n9752), .A2(n9394), .B1(n9391), .B2(n9750), .ZN(
        P2_U3534) );
  INV_X1 U10563 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n9392) );
  AOI22_X1 U10564 ( .A1(n9736), .A2(n9393), .B1(n9392), .B2(n9734), .ZN(
        P2_U3496) );
  INV_X1 U10565 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n9815) );
  AOI22_X1 U10566 ( .A1(n9736), .A2(n9394), .B1(n9815), .B2(n9734), .ZN(
        P2_U3493) );
  XNOR2_X1 U10567 ( .A(n9395), .B(n9396), .ZN(n9437) );
  NAND2_X1 U10568 ( .A1(n9398), .A2(n9397), .ZN(n9400) );
  AOI21_X1 U10569 ( .B1(n9401), .B2(n9400), .A(n9399), .ZN(n9404) );
  OAI22_X1 U10570 ( .A1(n9413), .A2(n9438), .B1(n9402), .B2(n9440), .ZN(n9403)
         );
  AOI211_X1 U10571 ( .C1(n9437), .C2(n9587), .A(n9404), .B(n9403), .ZN(n9434)
         );
  INV_X1 U10572 ( .A(n9405), .ZN(n9406) );
  AOI222_X1 U10573 ( .A1(n9407), .A2(n9554), .B1(P1_REG2_REG_13__SCAN_IN), 
        .B2(n9575), .C1(n9552), .C2(n9406), .ZN(n9411) );
  OAI211_X1 U10574 ( .C1(n9408), .C2(n9433), .A(n9559), .B(n4289), .ZN(n9432)
         );
  INV_X1 U10575 ( .A(n9432), .ZN(n9409) );
  AOI22_X1 U10576 ( .A1(n9437), .A2(n9563), .B1(n9562), .B2(n9409), .ZN(n9410)
         );
  OAI211_X1 U10577 ( .C1(n9575), .C2(n9434), .A(n9411), .B(n9410), .ZN(
        P1_U3278) );
  XNOR2_X1 U10578 ( .A(n9412), .B(n9416), .ZN(n9422) );
  OAI22_X1 U10579 ( .A1(n9414), .A2(n9438), .B1(n9413), .B2(n9440), .ZN(n9421)
         );
  NAND2_X1 U10580 ( .A1(n9415), .A2(n9416), .ZN(n9417) );
  NAND2_X1 U10581 ( .A1(n9418), .A2(n9417), .ZN(n9455) );
  NOR2_X1 U10582 ( .A1(n9455), .A2(n9419), .ZN(n9420) );
  AOI211_X1 U10583 ( .C1(n9550), .C2(n9422), .A(n9421), .B(n9420), .ZN(n9454)
         );
  INV_X1 U10584 ( .A(n9423), .ZN(n9424) );
  AOI222_X1 U10585 ( .A1(n9451), .A2(n9554), .B1(P1_REG2_REG_11__SCAN_IN), 
        .B2(n9575), .C1(n9424), .C2(n9552), .ZN(n9431) );
  INV_X1 U10586 ( .A(n9455), .ZN(n9429) );
  NAND2_X1 U10587 ( .A1(n9425), .A2(n9451), .ZN(n9426) );
  NAND2_X1 U10588 ( .A1(n9426), .A2(n9559), .ZN(n9427) );
  NOR2_X1 U10589 ( .A1(n9428), .A2(n9427), .ZN(n9450) );
  AOI22_X1 U10590 ( .A1(n9429), .A2(n9563), .B1(n9562), .B2(n9450), .ZN(n9430)
         );
  OAI211_X1 U10591 ( .C1(n9575), .C2(n9454), .A(n9431), .B(n9430), .ZN(
        P1_U3280) );
  INV_X1 U10592 ( .A(n9582), .ZN(n9594) );
  OAI21_X1 U10593 ( .B1(n9433), .B2(n9612), .A(n9432), .ZN(n9436) );
  INV_X1 U10594 ( .A(n9434), .ZN(n9435) );
  AOI211_X1 U10595 ( .C1(n9594), .C2(n9437), .A(n9436), .B(n9435), .ZN(n9457)
         );
  AOI22_X1 U10596 ( .A1(n4270), .A2(n9457), .B1(n6758), .B2(n9625), .ZN(
        P1_U3536) );
  OAI22_X1 U10597 ( .A1(n9441), .A2(n9440), .B1(n9439), .B2(n9438), .ZN(n9443)
         );
  AOI211_X1 U10598 ( .C1(n9452), .C2(n9444), .A(n9443), .B(n9442), .ZN(n9446)
         );
  OAI211_X1 U10599 ( .C1(n9447), .C2(n9582), .A(n9446), .B(n9445), .ZN(n9448)
         );
  AOI21_X1 U10600 ( .B1(n9587), .B2(n9449), .A(n9448), .ZN(n9458) );
  AOI22_X1 U10601 ( .A1(n4270), .A2(n9458), .B1(n6641), .B2(n9625), .ZN(
        P1_U3535) );
  AOI21_X1 U10602 ( .B1(n9452), .B2(n9451), .A(n9450), .ZN(n9453) );
  OAI211_X1 U10603 ( .C1(n9582), .C2(n9455), .A(n9454), .B(n9453), .ZN(n9456)
         );
  INV_X1 U10604 ( .A(n9456), .ZN(n9460) );
  AOI22_X1 U10605 ( .A1(n4270), .A2(n9460), .B1(n5183), .B2(n9625), .ZN(
        P1_U3534) );
  INV_X1 U10606 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n9914) );
  AOI22_X1 U10607 ( .A1(n9619), .A2(n9457), .B1(n9914), .B2(n9617), .ZN(
        P1_U3493) );
  AOI22_X1 U10608 ( .A1(n9619), .A2(n9458), .B1(n5215), .B2(n9617), .ZN(
        P1_U3490) );
  INV_X1 U10609 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n9459) );
  AOI22_X1 U10610 ( .A1(n9619), .A2(n9460), .B1(n9459), .B2(n9617), .ZN(
        P1_U3487) );
  XNOR2_X1 U10611 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U10612 ( .A(P2_RD_REG_SCAN_IN), .B(P1_RD_REG_SCAN_IN), .ZN(U126) );
  INV_X1 U10613 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n9482) );
  OAI211_X1 U10614 ( .C1(n9464), .C2(n9463), .A(n9462), .B(n9461), .ZN(n9465)
         );
  INV_X1 U10615 ( .A(n9465), .ZN(n9466) );
  OAI21_X1 U10616 ( .B1(n9468), .B2(n9467), .A(n9466), .ZN(n9496) );
  INV_X1 U10617 ( .A(n9496), .ZN(n9480) );
  OAI22_X1 U10618 ( .A1(n9533), .A2(n9470), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9469), .ZN(n9479) );
  XNOR2_X1 U10619 ( .A(n9472), .B(n9471), .ZN(n9477) );
  OAI211_X1 U10620 ( .C1(n9475), .C2(n9474), .A(n9540), .B(n9473), .ZN(n9476)
         );
  OAI21_X1 U10621 ( .B1(n9503), .B2(n9477), .A(n9476), .ZN(n9478) );
  NOR3_X1 U10622 ( .A1(n9480), .A2(n9479), .A3(n9478), .ZN(n9481) );
  OAI21_X1 U10623 ( .B1(n9525), .B2(n9482), .A(n9481), .ZN(P1_U3243) );
  INV_X1 U10624 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n9498) );
  INV_X1 U10625 ( .A(n9483), .ZN(n9495) );
  AOI21_X1 U10626 ( .B1(n9486), .B2(n9485), .A(n9484), .ZN(n9492) );
  AOI21_X1 U10627 ( .B1(n9489), .B2(n9488), .A(n9487), .ZN(n9491) );
  OAI22_X1 U10628 ( .A1(n9503), .A2(n9492), .B1(n9491), .B2(n9490), .ZN(n9493)
         );
  AOI211_X1 U10629 ( .C1(n9514), .C2(n9495), .A(n9494), .B(n9493), .ZN(n9497)
         );
  OAI211_X1 U10630 ( .C1(n9498), .C2(n9525), .A(n9497), .B(n9496), .ZN(
        P1_U3245) );
  AOI22_X1 U10631 ( .A1(n9539), .A2(P1_ADDR_REG_9__SCAN_IN), .B1(n9514), .B2(
        n9499), .ZN(n9511) );
  OAI21_X1 U10632 ( .B1(n9502), .B2(n9501), .A(n9500), .ZN(n9509) );
  AOI211_X1 U10633 ( .C1(n9506), .C2(n9505), .A(n9504), .B(n9503), .ZN(n9507)
         );
  AOI211_X1 U10634 ( .C1(n9540), .C2(n9509), .A(n9508), .B(n9507), .ZN(n9510)
         );
  NAND2_X1 U10635 ( .A1(n9511), .A2(n9510), .ZN(P1_U3250) );
  INV_X1 U10636 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n9524) );
  AOI21_X1 U10637 ( .B1(n9514), .B2(n9513), .A(n9512), .ZN(n9523) );
  XNOR2_X1 U10638 ( .A(n9516), .B(n9515), .ZN(n9521) );
  OAI21_X1 U10639 ( .B1(n9519), .B2(n9518), .A(n9517), .ZN(n9520) );
  AOI22_X1 U10640 ( .A1(n9540), .A2(n9521), .B1(n9530), .B2(n9520), .ZN(n9522)
         );
  OAI211_X1 U10641 ( .C1(n9525), .C2(n9524), .A(n9523), .B(n9522), .ZN(
        P1_U3255) );
  AOI21_X1 U10642 ( .B1(n9528), .B2(n9527), .A(n9526), .ZN(n9529) );
  NAND2_X1 U10643 ( .A1(n9530), .A2(n9529), .ZN(n9532) );
  OAI211_X1 U10644 ( .C1(n9534), .C2(n9533), .A(n9532), .B(n9531), .ZN(n9535)
         );
  INV_X1 U10645 ( .A(n9535), .ZN(n9543) );
  OAI21_X1 U10646 ( .B1(n9538), .B2(n9537), .A(n9536), .ZN(n9541) );
  AOI22_X1 U10647 ( .A1(n9541), .A2(n9540), .B1(n9539), .B2(
        P1_ADDR_REG_18__SCAN_IN), .ZN(n9542) );
  NAND2_X1 U10648 ( .A1(n9543), .A2(n9542), .ZN(P1_U3259) );
  NAND2_X1 U10649 ( .A1(n9545), .A2(n9544), .ZN(n9546) );
  XOR2_X1 U10650 ( .A(n9556), .B(n9546), .Z(n9549) );
  AOI222_X1 U10651 ( .A1(n9550), .A2(n9549), .B1(n9548), .B2(n9600), .C1(n9547), .C2(n9603), .ZN(n9611) );
  INV_X1 U10652 ( .A(n9551), .ZN(n9553) );
  AOI222_X1 U10653 ( .A1(n9555), .A2(n9554), .B1(P1_REG2_REG_9__SCAN_IN), .B2(
        n9575), .C1(n9553), .C2(n9552), .ZN(n9565) );
  XNOR2_X1 U10654 ( .A(n9557), .B(n9556), .ZN(n9616) );
  OAI211_X1 U10655 ( .C1(n9560), .C2(n9613), .A(n9559), .B(n9558), .ZN(n9610)
         );
  INV_X1 U10656 ( .A(n9610), .ZN(n9561) );
  AOI22_X1 U10657 ( .A1(n9616), .A2(n9563), .B1(n9562), .B2(n9561), .ZN(n9564)
         );
  OAI211_X1 U10658 ( .C1(n9575), .C2(n9611), .A(n9565), .B(n9564), .ZN(
        P1_U3282) );
  INV_X1 U10659 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n9574) );
  NOR2_X1 U10660 ( .A1(n9567), .A2(n9566), .ZN(n9569) );
  AOI211_X1 U10661 ( .C1(n9571), .C2(n9570), .A(n9569), .B(n9568), .ZN(n9573)
         );
  AOI22_X1 U10662 ( .A1(n9575), .A2(n9574), .B1(n9573), .B2(n9572), .ZN(
        P1_U3291) );
  AND2_X1 U10663 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n9579), .ZN(P1_U3292) );
  AND2_X1 U10664 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n9579), .ZN(P1_U3293) );
  AND2_X1 U10665 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n9579), .ZN(P1_U3294) );
  AND2_X1 U10666 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n9579), .ZN(P1_U3295) );
  AND2_X1 U10667 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n9579), .ZN(P1_U3296) );
  AND2_X1 U10668 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n9579), .ZN(P1_U3297) );
  AND2_X1 U10669 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n9579), .ZN(P1_U3298) );
  AND2_X1 U10670 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9579), .ZN(P1_U3299) );
  AND2_X1 U10671 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n9579), .ZN(P1_U3300) );
  INV_X1 U10672 ( .A(P1_D_REG_22__SCAN_IN), .ZN(n9913) );
  NOR2_X1 U10673 ( .A1(n9578), .A2(n9913), .ZN(P1_U3301) );
  AND2_X1 U10674 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n9579), .ZN(P1_U3302) );
  INV_X1 U10675 ( .A(P1_D_REG_20__SCAN_IN), .ZN(n9871) );
  NOR2_X1 U10676 ( .A1(n9578), .A2(n9871), .ZN(P1_U3303) );
  AND2_X1 U10677 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n9579), .ZN(P1_U3304) );
  AND2_X1 U10678 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n9579), .ZN(P1_U3305) );
  AND2_X1 U10679 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n9579), .ZN(P1_U3306) );
  AND2_X1 U10680 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n9579), .ZN(P1_U3307) );
  AND2_X1 U10681 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n9579), .ZN(P1_U3308) );
  AND2_X1 U10682 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n9579), .ZN(P1_U3309) );
  AND2_X1 U10683 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n9579), .ZN(P1_U3310) );
  INV_X1 U10684 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n9910) );
  NOR2_X1 U10685 ( .A1(n9578), .A2(n9910), .ZN(P1_U3311) );
  AND2_X1 U10686 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n9579), .ZN(P1_U3312) );
  AND2_X1 U10687 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n9579), .ZN(P1_U3313) );
  AND2_X1 U10688 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n9579), .ZN(P1_U3314) );
  INV_X1 U10689 ( .A(P1_D_REG_8__SCAN_IN), .ZN(n9904) );
  NOR2_X1 U10690 ( .A1(n9578), .A2(n9904), .ZN(P1_U3315) );
  AND2_X1 U10691 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n9579), .ZN(P1_U3316) );
  AND2_X1 U10692 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n9579), .ZN(P1_U3317) );
  AND2_X1 U10693 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n9579), .ZN(P1_U3318) );
  AND2_X1 U10694 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n9579), .ZN(P1_U3319) );
  AND2_X1 U10695 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n9579), .ZN(P1_U3320) );
  AND2_X1 U10696 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n9579), .ZN(P1_U3321) );
  INV_X1 U10697 ( .A(n9583), .ZN(n9586) );
  OAI211_X1 U10698 ( .C1(n9583), .C2(n9582), .A(n9581), .B(n9580), .ZN(n9585)
         );
  AOI211_X1 U10699 ( .C1(n9587), .C2(n9586), .A(n9585), .B(n9584), .ZN(n9621)
         );
  AOI22_X1 U10700 ( .A1(n9619), .A2(n9621), .B1(n4918), .B2(n9617), .ZN(
        P1_U3457) );
  INV_X1 U10701 ( .A(n9588), .ZN(n9589) );
  OAI21_X1 U10702 ( .B1(n9590), .B2(n9612), .A(n9589), .ZN(n9592) );
  AOI211_X1 U10703 ( .C1(n9594), .C2(n9593), .A(n9592), .B(n9591), .ZN(n9622)
         );
  AOI22_X1 U10704 ( .A1(n9619), .A2(n9622), .B1(n4963), .B2(n9617), .ZN(
        P1_U3463) );
  OAI21_X1 U10705 ( .B1(n9596), .B2(n9612), .A(n9595), .ZN(n9597) );
  AOI211_X1 U10706 ( .C1(n9599), .C2(n9615), .A(n9598), .B(n9597), .ZN(n9623)
         );
  AOI22_X1 U10707 ( .A1(n9619), .A2(n9623), .B1(n5015), .B2(n9617), .ZN(
        P1_U3469) );
  AOI22_X1 U10708 ( .A1(n9603), .A2(n9602), .B1(n9601), .B2(n9600), .ZN(n9604)
         );
  OAI211_X1 U10709 ( .C1(n4268), .C2(n9612), .A(n9605), .B(n9604), .ZN(n9607)
         );
  AOI211_X1 U10710 ( .C1(n9615), .C2(n9608), .A(n9607), .B(n9606), .ZN(n9624)
         );
  INV_X1 U10711 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n9609) );
  AOI22_X1 U10712 ( .A1(n9619), .A2(n9624), .B1(n9609), .B2(n9617), .ZN(
        P1_U3472) );
  OAI211_X1 U10713 ( .C1(n9613), .C2(n9612), .A(n9611), .B(n9610), .ZN(n9614)
         );
  AOI21_X1 U10714 ( .B1(n9616), .B2(n9615), .A(n9614), .ZN(n9626) );
  INV_X1 U10715 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n9618) );
  AOI22_X1 U10716 ( .A1(n9619), .A2(n9626), .B1(n9618), .B2(n9617), .ZN(
        P1_U3481) );
  INV_X1 U10717 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n9620) );
  AOI22_X1 U10718 ( .A1(n4270), .A2(n9621), .B1(n9620), .B2(n9625), .ZN(
        P1_U3524) );
  AOI22_X1 U10719 ( .A1(n4270), .A2(n9622), .B1(n6409), .B2(n9625), .ZN(
        P1_U3526) );
  AOI22_X1 U10720 ( .A1(n4270), .A2(n9623), .B1(n6418), .B2(n9625), .ZN(
        P1_U3528) );
  AOI22_X1 U10721 ( .A1(n4270), .A2(n9624), .B1(n5039), .B2(n9625), .ZN(
        P1_U3529) );
  AOI22_X1 U10722 ( .A1(n4270), .A2(n9626), .B1(n5124), .B2(n9625), .ZN(
        P1_U3532) );
  AOI22_X1 U10723 ( .A1(n9632), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n9627), .ZN(n9637) );
  OAI21_X1 U10724 ( .B1(n9629), .B2(P2_REG1_REG_0__SCAN_IN), .A(n9628), .ZN(
        n9630) );
  AOI21_X1 U10725 ( .B1(n9632), .B2(n9631), .A(n9630), .ZN(n9635) );
  AOI22_X1 U10726 ( .A1(n9633), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3152), .ZN(n9634) );
  OAI221_X1 U10727 ( .B1(n9638), .B2(n9637), .C1(n9636), .C2(n9635), .A(n9634), 
        .ZN(P2_U3245) );
  INV_X1 U10728 ( .A(n9639), .ZN(n9640) );
  AOI21_X1 U10729 ( .B1(n9650), .B2(n9641), .A(n9640), .ZN(n9704) );
  INV_X1 U10730 ( .A(n9642), .ZN(n9645) );
  INV_X1 U10731 ( .A(n9643), .ZN(n9644) );
  OAI21_X1 U10732 ( .B1(n9700), .B2(n9645), .A(n9644), .ZN(n9701) );
  INV_X1 U10733 ( .A(n9701), .ZN(n9646) );
  AOI22_X1 U10734 ( .A1(n9704), .A2(n9648), .B1(n9647), .B2(n9646), .ZN(n9667)
         );
  NOR2_X1 U10735 ( .A1(n9649), .A2(n9700), .ZN(n9663) );
  XNOR2_X1 U10736 ( .A(n9651), .B(n9650), .ZN(n9659) );
  NAND2_X1 U10737 ( .A1(n9704), .A2(n9652), .ZN(n9658) );
  AOI22_X1 U10738 ( .A1(n9656), .A2(n9655), .B1(n9654), .B2(n9653), .ZN(n9657)
         );
  OAI211_X1 U10739 ( .C1(n9660), .C2(n9659), .A(n9658), .B(n9657), .ZN(n9702)
         );
  MUX2_X1 U10740 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n9702), .S(n9661), .Z(n9662)
         );
  AOI211_X1 U10741 ( .C1(n9665), .C2(n9664), .A(n9663), .B(n9662), .ZN(n9666)
         );
  NAND2_X1 U10742 ( .A1(n9667), .A2(n9666), .ZN(P2_U3288) );
  AND2_X1 U10743 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n9926), .ZN(P2_U3297) );
  AND2_X1 U10744 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n9926), .ZN(P2_U3298) );
  AND2_X1 U10745 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n9926), .ZN(P2_U3299) );
  AND2_X1 U10746 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n9926), .ZN(P2_U3300) );
  AND2_X1 U10747 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n9926), .ZN(P2_U3301) );
  AND2_X1 U10748 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n9926), .ZN(P2_U3302) );
  AND2_X1 U10749 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n9926), .ZN(P2_U3303) );
  AND2_X1 U10750 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n9926), .ZN(P2_U3304) );
  AND2_X1 U10751 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n9926), .ZN(P2_U3305) );
  AND2_X1 U10752 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n9926), .ZN(P2_U3306) );
  AND2_X1 U10753 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n9926), .ZN(P2_U3307) );
  AND2_X1 U10754 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n9926), .ZN(P2_U3309) );
  AND2_X1 U10755 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n9926), .ZN(P2_U3310) );
  AND2_X1 U10756 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n9926), .ZN(P2_U3311) );
  INV_X1 U10757 ( .A(P2_D_REG_16__SCAN_IN), .ZN(n9893) );
  NOR2_X1 U10758 ( .A1(n9670), .A2(n9893), .ZN(P2_U3312) );
  AND2_X1 U10759 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n9926), .ZN(P2_U3313) );
  AND2_X1 U10760 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n9926), .ZN(P2_U3314) );
  AND2_X1 U10761 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n9926), .ZN(P2_U3315) );
  AND2_X1 U10762 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n9926), .ZN(P2_U3316) );
  INV_X1 U10763 ( .A(P2_D_REG_11__SCAN_IN), .ZN(n9867) );
  NOR2_X1 U10764 ( .A1(n9670), .A2(n9867), .ZN(P2_U3317) );
  AND2_X1 U10765 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n9926), .ZN(P2_U3318) );
  AND2_X1 U10766 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n9926), .ZN(P2_U3319) );
  AND2_X1 U10767 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n9926), .ZN(P2_U3320) );
  AND2_X1 U10768 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n9926), .ZN(P2_U3321) );
  AND2_X1 U10769 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n9926), .ZN(P2_U3322) );
  AND2_X1 U10770 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n9926), .ZN(P2_U3323) );
  INV_X1 U10771 ( .A(P2_D_REG_4__SCAN_IN), .ZN(n9852) );
  NOR2_X1 U10772 ( .A1(n9670), .A2(n9852), .ZN(P2_U3324) );
  AND2_X1 U10773 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n9926), .ZN(P2_U3325) );
  AND2_X1 U10774 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n9926), .ZN(P2_U3326) );
  AOI22_X1 U10775 ( .A1(n9675), .A2(n9672), .B1(n9671), .B2(n9926), .ZN(
        P2_U3437) );
  AOI22_X1 U10776 ( .A1(n9675), .A2(n9674), .B1(n9673), .B2(n9926), .ZN(
        P2_U3438) );
  OAI22_X1 U10777 ( .A1(n9679), .A2(n9678), .B1(n9677), .B2(n9676), .ZN(n9680)
         );
  NOR2_X1 U10778 ( .A1(n9681), .A2(n9680), .ZN(n9738) );
  INV_X1 U10779 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n9682) );
  AOI22_X1 U10780 ( .A1(n9736), .A2(n9738), .B1(n9682), .B2(n9734), .ZN(
        P2_U3451) );
  OAI22_X1 U10781 ( .A1(n9684), .A2(n9728), .B1(n9683), .B2(n9727), .ZN(n9686)
         );
  AOI211_X1 U10782 ( .C1(n9733), .C2(n9687), .A(n9686), .B(n9685), .ZN(n9740)
         );
  INV_X1 U10783 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n9688) );
  AOI22_X1 U10784 ( .A1(n9736), .A2(n9740), .B1(n9688), .B2(n9734), .ZN(
        P2_U3463) );
  INV_X1 U10785 ( .A(n9689), .ZN(n9690) );
  AOI211_X1 U10786 ( .C1(n9733), .C2(n9692), .A(n9691), .B(n9690), .ZN(n9741)
         );
  INV_X1 U10787 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n9693) );
  AOI22_X1 U10788 ( .A1(n9736), .A2(n9741), .B1(n9693), .B2(n9734), .ZN(
        P2_U3469) );
  OAI22_X1 U10789 ( .A1(n9695), .A2(n9728), .B1(n9694), .B2(n9727), .ZN(n9697)
         );
  AOI211_X1 U10790 ( .C1(n9698), .C2(n9733), .A(n9697), .B(n9696), .ZN(n9743)
         );
  INV_X1 U10791 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n9699) );
  AOI22_X1 U10792 ( .A1(n9736), .A2(n9743), .B1(n9699), .B2(n9734), .ZN(
        P2_U3472) );
  OAI22_X1 U10793 ( .A1(n9701), .A2(n9728), .B1(n9700), .B2(n9727), .ZN(n9703)
         );
  AOI211_X1 U10794 ( .C1(n9715), .C2(n9704), .A(n9703), .B(n9702), .ZN(n9745)
         );
  INV_X1 U10795 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n9705) );
  AOI22_X1 U10796 ( .A1(n9736), .A2(n9745), .B1(n9705), .B2(n9734), .ZN(
        P2_U3475) );
  OAI22_X1 U10797 ( .A1(n9707), .A2(n9728), .B1(n9706), .B2(n9727), .ZN(n9708)
         );
  AOI21_X1 U10798 ( .B1(n9709), .B2(n9715), .A(n9708), .ZN(n9710) );
  AND2_X1 U10799 ( .A1(n9711), .A2(n9710), .ZN(n9746) );
  INV_X1 U10800 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n9877) );
  AOI22_X1 U10801 ( .A1(n9736), .A2(n9746), .B1(n9877), .B2(n9734), .ZN(
        P2_U3478) );
  OAI22_X1 U10802 ( .A1(n9713), .A2(n9728), .B1(n9712), .B2(n9727), .ZN(n9714)
         );
  AOI21_X1 U10803 ( .B1(n9716), .B2(n9715), .A(n9714), .ZN(n9717) );
  AND2_X1 U10804 ( .A1(n9718), .A2(n9717), .ZN(n9747) );
  INV_X1 U10805 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n9719) );
  AOI22_X1 U10806 ( .A1(n9736), .A2(n9747), .B1(n9719), .B2(n9734), .ZN(
        P2_U3481) );
  INV_X1 U10807 ( .A(n9720), .ZN(n9725) );
  OAI22_X1 U10808 ( .A1(n9722), .A2(n9728), .B1(n9721), .B2(n9727), .ZN(n9724)
         );
  AOI211_X1 U10809 ( .C1(n9725), .C2(n9733), .A(n9724), .B(n9723), .ZN(n9749)
         );
  INV_X1 U10810 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n9726) );
  AOI22_X1 U10811 ( .A1(n9736), .A2(n9749), .B1(n9726), .B2(n9734), .ZN(
        P2_U3484) );
  OAI22_X1 U10812 ( .A1(n9729), .A2(n9728), .B1(n4464), .B2(n9727), .ZN(n9731)
         );
  AOI211_X1 U10813 ( .C1(n9733), .C2(n9732), .A(n9731), .B(n9730), .ZN(n9751)
         );
  INV_X1 U10814 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n9735) );
  AOI22_X1 U10815 ( .A1(n9736), .A2(n9751), .B1(n9735), .B2(n9734), .ZN(
        P2_U3487) );
  AOI22_X1 U10816 ( .A1(n9752), .A2(n9738), .B1(n9737), .B2(n9750), .ZN(
        P2_U3520) );
  INV_X1 U10817 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n9739) );
  AOI22_X1 U10818 ( .A1(n9752), .A2(n9740), .B1(n9739), .B2(n9750), .ZN(
        P2_U3524) );
  AOI22_X1 U10819 ( .A1(n9752), .A2(n9741), .B1(n6446), .B2(n9750), .ZN(
        P2_U3526) );
  INV_X1 U10820 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n9742) );
  AOI22_X1 U10821 ( .A1(n9752), .A2(n9743), .B1(n9742), .B2(n9750), .ZN(
        P2_U3527) );
  AOI22_X1 U10822 ( .A1(n9752), .A2(n9745), .B1(n9744), .B2(n9750), .ZN(
        P2_U3528) );
  AOI22_X1 U10823 ( .A1(n9752), .A2(n9746), .B1(n6534), .B2(n9750), .ZN(
        P2_U3529) );
  AOI22_X1 U10824 ( .A1(n9752), .A2(n9747), .B1(n6537), .B2(n9750), .ZN(
        P2_U3530) );
  AOI22_X1 U10825 ( .A1(n9752), .A2(n9749), .B1(n9748), .B2(n9750), .ZN(
        P2_U3531) );
  AOI22_X1 U10826 ( .A1(n9752), .A2(n9751), .B1(n6663), .B2(n9750), .ZN(
        P2_U3532) );
  INV_X1 U10827 ( .A(n9753), .ZN(n9754) );
  NAND2_X1 U10828 ( .A1(n9755), .A2(n9754), .ZN(n9756) );
  XNOR2_X1 U10829 ( .A(P2_ADDR_REG_1__SCAN_IN), .B(n9756), .ZN(ADD_1071_U5) );
  XOR2_X1 U10830 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1071_U46) );
  OAI21_X1 U10831 ( .B1(n9759), .B2(n9758), .A(n9757), .ZN(ADD_1071_U56) );
  OAI21_X1 U10832 ( .B1(n9762), .B2(n9761), .A(n9760), .ZN(ADD_1071_U57) );
  OAI21_X1 U10833 ( .B1(n9765), .B2(n9764), .A(n9763), .ZN(ADD_1071_U58) );
  OAI21_X1 U10834 ( .B1(n9768), .B2(n9767), .A(n9766), .ZN(ADD_1071_U59) );
  OAI21_X1 U10835 ( .B1(n9771), .B2(n9770), .A(n9769), .ZN(ADD_1071_U60) );
  OAI21_X1 U10836 ( .B1(n9774), .B2(n9773), .A(n9772), .ZN(ADD_1071_U61) );
  AOI21_X1 U10837 ( .B1(n9777), .B2(n9776), .A(n9775), .ZN(ADD_1071_U62) );
  AOI21_X1 U10838 ( .B1(n9780), .B2(n9779), .A(n9778), .ZN(ADD_1071_U63) );
  NAND3_X1 U10839 ( .A1(keyinput58), .A2(keyinput33), .A3(keyinput46), .ZN(
        n9787) );
  INV_X1 U10840 ( .A(keyinput35), .ZN(n9781) );
  NAND4_X1 U10841 ( .A1(keyinput59), .A2(keyinput27), .A3(keyinput14), .A4(
        n9781), .ZN(n9786) );
  NOR3_X1 U10842 ( .A1(keyinput55), .A2(keyinput13), .A3(keyinput2), .ZN(n9784) );
  INV_X1 U10843 ( .A(keyinput11), .ZN(n9782) );
  NOR3_X1 U10844 ( .A1(keyinput56), .A2(keyinput44), .A3(n9782), .ZN(n9783) );
  NAND4_X1 U10845 ( .A1(keyinput4), .A2(n9784), .A3(keyinput20), .A4(n9783), 
        .ZN(n9785) );
  NOR4_X1 U10846 ( .A1(keyinput60), .A2(n9787), .A3(n9786), .A4(n9785), .ZN(
        n9925) );
  NAND3_X1 U10847 ( .A1(keyinput45), .A2(keyinput63), .A3(keyinput53), .ZN(
        n9806) );
  NOR2_X1 U10848 ( .A1(keyinput36), .A2(keyinput49), .ZN(n9791) );
  NAND3_X1 U10849 ( .A1(keyinput7), .A2(keyinput41), .A3(keyinput34), .ZN(
        n9789) );
  NAND3_X1 U10850 ( .A1(keyinput54), .A2(keyinput12), .A3(keyinput10), .ZN(
        n9788) );
  NOR4_X1 U10851 ( .A1(keyinput9), .A2(keyinput1), .A3(n9789), .A4(n9788), 
        .ZN(n9790) );
  NAND4_X1 U10852 ( .A1(keyinput8), .A2(keyinput24), .A3(n9791), .A4(n9790), 
        .ZN(n9805) );
  NOR3_X1 U10853 ( .A1(keyinput52), .A2(keyinput16), .A3(keyinput39), .ZN(
        n9803) );
  NAND2_X1 U10854 ( .A1(keyinput3), .A2(keyinput37), .ZN(n9795) );
  NOR2_X1 U10855 ( .A1(keyinput38), .A2(keyinput50), .ZN(n9793) );
  NOR4_X1 U10856 ( .A1(keyinput22), .A2(keyinput25), .A3(keyinput61), .A4(
        keyinput62), .ZN(n9792) );
  NAND4_X1 U10857 ( .A1(keyinput29), .A2(keyinput18), .A3(n9793), .A4(n9792), 
        .ZN(n9794) );
  NOR4_X1 U10858 ( .A1(keyinput17), .A2(keyinput57), .A3(n9795), .A4(n9794), 
        .ZN(n9802) );
  NAND4_X1 U10859 ( .A1(keyinput21), .A2(keyinput6), .A3(keyinput28), .A4(
        keyinput23), .ZN(n9800) );
  NAND3_X1 U10860 ( .A1(keyinput30), .A2(keyinput5), .A3(keyinput42), .ZN(
        n9799) );
  NOR2_X1 U10861 ( .A1(keyinput51), .A2(keyinput47), .ZN(n9797) );
  NOR4_X1 U10862 ( .A1(keyinput19), .A2(keyinput40), .A3(keyinput31), .A4(
        keyinput32), .ZN(n9796) );
  NAND4_X1 U10863 ( .A1(keyinput26), .A2(keyinput15), .A3(n9797), .A4(n9796), 
        .ZN(n9798) );
  NOR4_X1 U10864 ( .A1(keyinput48), .A2(n9800), .A3(n9799), .A4(n9798), .ZN(
        n9801) );
  NAND4_X1 U10865 ( .A1(keyinput43), .A2(n9803), .A3(n9802), .A4(n9801), .ZN(
        n9804) );
  NOR4_X1 U10866 ( .A1(keyinput0), .A2(n9806), .A3(n9805), .A4(n9804), .ZN(
        n9924) );
  INV_X1 U10867 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n9808) );
  AOI22_X1 U10868 ( .A1(n9809), .A2(keyinput16), .B1(keyinput39), .B2(n9808), 
        .ZN(n9807) );
  OAI221_X1 U10869 ( .B1(n9809), .B2(keyinput16), .C1(n9808), .C2(keyinput39), 
        .A(n9807), .ZN(n9821) );
  AOI22_X1 U10870 ( .A1(n6051), .A2(keyinput3), .B1(n9811), .B2(keyinput37), 
        .ZN(n9810) );
  OAI221_X1 U10871 ( .B1(n6051), .B2(keyinput3), .C1(n9811), .C2(keyinput37), 
        .A(n9810), .ZN(n9820) );
  AOI22_X1 U10872 ( .A1(n9814), .A2(keyinput52), .B1(keyinput43), .B2(n9813), 
        .ZN(n9812) );
  OAI221_X1 U10873 ( .B1(n9814), .B2(keyinput52), .C1(n9813), .C2(keyinput43), 
        .A(n9812), .ZN(n9819) );
  XOR2_X1 U10874 ( .A(n9815), .B(keyinput57), .Z(n9817) );
  XNOR2_X1 U10875 ( .A(P2_IR_REG_9__SCAN_IN), .B(keyinput17), .ZN(n9816) );
  NAND2_X1 U10876 ( .A1(n9817), .A2(n9816), .ZN(n9818) );
  NOR4_X1 U10877 ( .A1(n9821), .A2(n9820), .A3(n9819), .A4(n9818), .ZN(n9861)
         );
  AOI22_X1 U10878 ( .A1(n9823), .A2(keyinput29), .B1(n5987), .B2(keyinput38), 
        .ZN(n9822) );
  OAI221_X1 U10879 ( .B1(n9823), .B2(keyinput29), .C1(n5987), .C2(keyinput38), 
        .A(n9822), .ZN(n9833) );
  AOI22_X1 U10880 ( .A1(n5041), .A2(keyinput18), .B1(keyinput50), .B2(n6188), 
        .ZN(n9824) );
  OAI221_X1 U10881 ( .B1(n5041), .B2(keyinput18), .C1(n6188), .C2(keyinput50), 
        .A(n9824), .ZN(n9832) );
  AOI22_X1 U10882 ( .A1(n6663), .A2(keyinput22), .B1(n9826), .B2(keyinput25), 
        .ZN(n9825) );
  OAI221_X1 U10883 ( .B1(n6663), .B2(keyinput22), .C1(n9826), .C2(keyinput25), 
        .A(n9825), .ZN(n9831) );
  AOI22_X1 U10884 ( .A1(n9829), .A2(keyinput61), .B1(keyinput62), .B2(n9828), 
        .ZN(n9827) );
  OAI221_X1 U10885 ( .B1(n9829), .B2(keyinput61), .C1(n9828), .C2(keyinput62), 
        .A(n9827), .ZN(n9830) );
  NOR4_X1 U10886 ( .A1(n9833), .A2(n9832), .A3(n9831), .A4(n9830), .ZN(n9860)
         );
  AOI22_X1 U10887 ( .A1(n9836), .A2(keyinput41), .B1(n9835), .B2(keyinput34), 
        .ZN(n9834) );
  OAI221_X1 U10888 ( .B1(n9836), .B2(keyinput41), .C1(n9835), .C2(keyinput34), 
        .A(n9834), .ZN(n9845) );
  XNOR2_X1 U10889 ( .A(P1_IR_REG_8__SCAN_IN), .B(keyinput63), .ZN(n9840) );
  XNOR2_X1 U10890 ( .A(SI_2_), .B(keyinput0), .ZN(n9839) );
  XNOR2_X1 U10891 ( .A(P2_IR_REG_14__SCAN_IN), .B(keyinput9), .ZN(n9838) );
  XNOR2_X1 U10892 ( .A(P2_REG1_REG_17__SCAN_IN), .B(keyinput53), .ZN(n9837) );
  NAND4_X1 U10893 ( .A1(n9840), .A2(n9839), .A3(n9838), .A4(n9837), .ZN(n9844)
         );
  XNOR2_X1 U10894 ( .A(keyinput45), .B(n5482), .ZN(n9843) );
  INV_X1 U10895 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n9841) );
  XNOR2_X1 U10896 ( .A(keyinput7), .B(n9841), .ZN(n9842) );
  NOR4_X1 U10897 ( .A1(n9845), .A2(n9844), .A3(n9843), .A4(n9842), .ZN(n9859)
         );
  INV_X1 U10898 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n9848) );
  AOI22_X1 U10899 ( .A1(n9848), .A2(keyinput36), .B1(keyinput8), .B2(n9847), 
        .ZN(n9846) );
  OAI221_X1 U10900 ( .B1(n9848), .B2(keyinput36), .C1(n9847), .C2(keyinput8), 
        .A(n9846), .ZN(n9857) );
  AOI22_X1 U10901 ( .A1(n4897), .A2(keyinput49), .B1(keyinput24), .B2(n4894), 
        .ZN(n9849) );
  OAI221_X1 U10902 ( .B1(n4897), .B2(keyinput49), .C1(n4894), .C2(keyinput24), 
        .A(n9849), .ZN(n9856) );
  AOI22_X1 U10903 ( .A1(n9852), .A2(keyinput54), .B1(n9851), .B2(keyinput12), 
        .ZN(n9850) );
  OAI221_X1 U10904 ( .B1(n9852), .B2(keyinput54), .C1(n9851), .C2(keyinput12), 
        .A(n9850), .ZN(n9855) );
  AOI22_X1 U10905 ( .A1(n5737), .A2(keyinput10), .B1(n6418), .B2(keyinput1), 
        .ZN(n9853) );
  OAI221_X1 U10906 ( .B1(n5737), .B2(keyinput10), .C1(n6418), .C2(keyinput1), 
        .A(n9853), .ZN(n9854) );
  NOR4_X1 U10907 ( .A1(n9857), .A2(n9856), .A3(n9855), .A4(n9854), .ZN(n9858)
         );
  NAND4_X1 U10908 ( .A1(n9861), .A2(n9860), .A3(n9859), .A4(n9858), .ZN(n9923)
         );
  AOI22_X1 U10909 ( .A1(n9056), .A2(keyinput11), .B1(keyinput44), .B2(n9863), 
        .ZN(n9862) );
  OAI221_X1 U10910 ( .B1(n9056), .B2(keyinput11), .C1(n9863), .C2(keyinput44), 
        .A(n9862), .ZN(n9875) );
  AOI22_X1 U10911 ( .A1(n6527), .A2(keyinput20), .B1(n9865), .B2(keyinput56), 
        .ZN(n9864) );
  OAI221_X1 U10912 ( .B1(n6527), .B2(keyinput20), .C1(n9865), .C2(keyinput56), 
        .A(n9864), .ZN(n9874) );
  INV_X1 U10913 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n9868) );
  AOI22_X1 U10914 ( .A1(n9868), .A2(keyinput27), .B1(n9867), .B2(keyinput14), 
        .ZN(n9866) );
  OAI221_X1 U10915 ( .B1(n9868), .B2(keyinput27), .C1(n9867), .C2(keyinput14), 
        .A(n9866), .ZN(n9873) );
  INV_X1 U10916 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n9870) );
  AOI22_X1 U10917 ( .A1(n9871), .A2(keyinput35), .B1(keyinput59), .B2(n9870), 
        .ZN(n9869) );
  OAI221_X1 U10918 ( .B1(n9871), .B2(keyinput35), .C1(n9870), .C2(keyinput59), 
        .A(n9869), .ZN(n9872) );
  NOR4_X1 U10919 ( .A1(n9875), .A2(n9874), .A3(n9873), .A4(n9872), .ZN(n9921)
         );
  AOI22_X1 U10920 ( .A1(n9878), .A2(keyinput33), .B1(keyinput46), .B2(n9877), 
        .ZN(n9876) );
  OAI221_X1 U10921 ( .B1(n9878), .B2(keyinput33), .C1(n9877), .C2(keyinput46), 
        .A(n9876), .ZN(n9889) );
  AOI22_X1 U10922 ( .A1(n6395), .A2(keyinput58), .B1(n9880), .B2(keyinput60), 
        .ZN(n9879) );
  OAI221_X1 U10923 ( .B1(n6395), .B2(keyinput58), .C1(n9880), .C2(keyinput60), 
        .A(n9879), .ZN(n9888) );
  INV_X1 U10924 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n9882) );
  AOI22_X1 U10925 ( .A1(n4858), .A2(keyinput2), .B1(keyinput4), .B2(n9882), 
        .ZN(n9881) );
  OAI221_X1 U10926 ( .B1(n4858), .B2(keyinput2), .C1(n9882), .C2(keyinput4), 
        .A(n9881), .ZN(n9887) );
  AOI22_X1 U10927 ( .A1(n9885), .A2(keyinput55), .B1(keyinput13), .B2(n9884), 
        .ZN(n9883) );
  OAI221_X1 U10928 ( .B1(n9885), .B2(keyinput55), .C1(n9884), .C2(keyinput13), 
        .A(n9883), .ZN(n9886) );
  NOR4_X1 U10929 ( .A1(n9889), .A2(n9888), .A3(n9887), .A4(n9886), .ZN(n9920)
         );
  AOI22_X1 U10930 ( .A1(n5072), .A2(keyinput30), .B1(keyinput5), .B2(n9891), 
        .ZN(n9890) );
  OAI221_X1 U10931 ( .B1(n5072), .B2(keyinput30), .C1(n9891), .C2(keyinput5), 
        .A(n9890), .ZN(n9901) );
  AOI22_X1 U10932 ( .A1(n9941), .A2(keyinput28), .B1(n9893), .B2(keyinput23), 
        .ZN(n9892) );
  OAI221_X1 U10933 ( .B1(n9941), .B2(keyinput28), .C1(n9893), .C2(keyinput23), 
        .A(n9892), .ZN(n9900) );
  XOR2_X1 U10934 ( .A(n9894), .B(keyinput21), .Z(n9898) );
  XNOR2_X1 U10935 ( .A(P2_IR_REG_31__SCAN_IN), .B(keyinput6), .ZN(n9897) );
  XNOR2_X1 U10936 ( .A(P2_REG3_REG_20__SCAN_IN), .B(keyinput42), .ZN(n9896) );
  XNOR2_X1 U10937 ( .A(P1_IR_REG_5__SCAN_IN), .B(keyinput48), .ZN(n9895) );
  NAND4_X1 U10938 ( .A1(n9898), .A2(n9897), .A3(n9896), .A4(n9895), .ZN(n9899)
         );
  NOR3_X1 U10939 ( .A1(n9901), .A2(n9900), .A3(n9899), .ZN(n9919) );
  AOI22_X1 U10940 ( .A1(n5166), .A2(keyinput31), .B1(n9903), .B2(keyinput32), 
        .ZN(n9902) );
  OAI221_X1 U10941 ( .B1(n5166), .B2(keyinput31), .C1(n9903), .C2(keyinput32), 
        .A(n9902), .ZN(n9908) );
  XNOR2_X1 U10942 ( .A(n9904), .B(keyinput40), .ZN(n9907) );
  XNOR2_X1 U10943 ( .A(n9905), .B(keyinput19), .ZN(n9906) );
  OR3_X1 U10944 ( .A1(n9908), .A2(n9907), .A3(n9906), .ZN(n9917) );
  INV_X1 U10945 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n9911) );
  AOI22_X1 U10946 ( .A1(n9911), .A2(keyinput51), .B1(n9910), .B2(keyinput26), 
        .ZN(n9909) );
  OAI221_X1 U10947 ( .B1(n9911), .B2(keyinput51), .C1(n9910), .C2(keyinput26), 
        .A(n9909), .ZN(n9916) );
  AOI22_X1 U10948 ( .A1(n9914), .A2(keyinput47), .B1(n9913), .B2(keyinput15), 
        .ZN(n9912) );
  OAI221_X1 U10949 ( .B1(n9914), .B2(keyinput47), .C1(n9913), .C2(keyinput15), 
        .A(n9912), .ZN(n9915) );
  NOR3_X1 U10950 ( .A1(n9917), .A2(n9916), .A3(n9915), .ZN(n9918) );
  NAND4_X1 U10951 ( .A1(n9921), .A2(n9920), .A3(n9919), .A4(n9918), .ZN(n9922)
         );
  AOI211_X1 U10952 ( .C1(n9925), .C2(n9924), .A(n9923), .B(n9922), .ZN(n9928)
         );
  NAND2_X1 U10953 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n9926), .ZN(n9927) );
  XNOR2_X1 U10954 ( .A(n9928), .B(n9927), .ZN(P2_U3308) );
  XOR2_X1 U10955 ( .A(n9929), .B(P2_ADDR_REG_6__SCAN_IN), .Z(ADD_1071_U50) );
  NOR2_X1 U10956 ( .A1(n9931), .A2(n9930), .ZN(n9932) );
  XOR2_X1 U10957 ( .A(P1_ADDR_REG_5__SCAN_IN), .B(n9932), .Z(ADD_1071_U51) );
  XOR2_X1 U10958 ( .A(n9933), .B(P2_ADDR_REG_8__SCAN_IN), .Z(ADD_1071_U48) );
  OAI21_X1 U10959 ( .B1(n9936), .B2(n9935), .A(n9934), .ZN(n9937) );
  XNOR2_X1 U10960 ( .A(n9937), .B(P1_ADDR_REG_18__SCAN_IN), .ZN(ADD_1071_U55)
         );
  XOR2_X1 U10961 ( .A(n9938), .B(P2_ADDR_REG_7__SCAN_IN), .Z(ADD_1071_U49) );
  AOI21_X1 U10962 ( .B1(n9941), .B2(n9940), .A(n9939), .ZN(ADD_1071_U47) );
  XOR2_X1 U10963 ( .A(n9943), .B(n9942), .Z(ADD_1071_U54) );
  XOR2_X1 U10964 ( .A(n9945), .B(n9944), .Z(ADD_1071_U53) );
  XNOR2_X1 U10965 ( .A(n9947), .B(n9946), .ZN(ADD_1071_U52) );
  NAND2_X1 U4813 ( .A1(n4602), .A2(n4601), .ZN(n9006) );
  AOI21_X1 U6050 ( .B1(n4607), .B2(n8695), .A(n4281), .ZN(n4605) );
  NAND2_X1 U4776 ( .A1(n4362), .A2(n4361), .ZN(n7724) );
  AND2_X1 U4817 ( .A1(n6799), .A2(n6979), .ZN(n6973) );
  AOI211_X1 U5268 ( .C1(n9647), .C2(n8315), .A(n8104), .B(n8103), .ZN(n8105)
         );
  CLKBUF_X1 U5951 ( .A(n6260), .Z(n7528) );
endmodule

