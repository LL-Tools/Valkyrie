

module b22_C_AntiSAT_k_128_9 ( P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, 
        SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65, 
        SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70, 
        SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58, 
        SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53, 
        U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, 
        P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, 
        P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, 
        P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, 
        P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446, 
        P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, 
        P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, 
        P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, 
        P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, 
        P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, 
        P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, 
        P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513, 
        P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, 
        P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, 
        P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, 
        P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, 
        P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, 
        P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556, 
        P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290, 
        P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, 
        P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, 
        P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, 
        P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, 
        P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, 
        P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, 
        P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560, 
        P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, 
        P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, 
        P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, 
        P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588, 
        P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239, 
        P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, 
        P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, 
        P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, 
        P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, 
        P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, 
        P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, 
        P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, 
        P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, 
        P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442, 
        P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, 
        P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, 
        P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492, 
        P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, 
        P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, 
        P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, 
        P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, 
        P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, 
        P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262, 
        P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, 
        P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, 
        P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531, 
        P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, 
        P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, 
        P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552, 
        P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, 
        P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211, 
        P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, 
        P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, 
        P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, 
        P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087, 
        P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290, 
        P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283, 
        P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276, 
        P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269, 
        P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377, 
        P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257, 
        P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250, 
        P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243, 
        P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236, 
        P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402, 
        P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423, 
        P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444, 
        P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452, 
        P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459, 
        P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466, 
        P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473, 
        P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480, 
        P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487, 
        P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230, 
        P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223, 
        P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216, 
        P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209, 
        P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202, 
        P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195, 
        P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188, 
        P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491, 
        P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498, 
        P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505, 
        P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512, 
        P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519, 
        P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179, 
        P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172, 
        P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165, 
        P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158, 
        P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150, 
        P3_U3897 );
  input P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput0,
         keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6,
         keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12,
         keyinput13, keyinput14, keyinput15, keyinput16, keyinput17,
         keyinput18, keyinput19, keyinput20, keyinput21, keyinput22,
         keyinput23, keyinput24, keyinput25, keyinput26, keyinput27,
         keyinput28, keyinput29, keyinput30, keyinput31, keyinput32,
         keyinput33, keyinput34, keyinput35, keyinput36, keyinput37,
         keyinput38, keyinput39, keyinput40, keyinput41, keyinput42,
         keyinput43, keyinput44, keyinput45, keyinput46, keyinput47,
         keyinput48, keyinput49, keyinput50, keyinput51, keyinput52,
         keyinput53, keyinput54, keyinput55, keyinput56, keyinput57,
         keyinput58, keyinput59, keyinput60, keyinput61, keyinput62,
         keyinput63, keyinput64, keyinput65, keyinput66, keyinput67,
         keyinput68, keyinput69, keyinput70, keyinput71, keyinput72,
         keyinput73, keyinput74, keyinput75, keyinput76, keyinput77,
         keyinput78, keyinput79, keyinput80, keyinput81, keyinput82,
         keyinput83, keyinput84, keyinput85, keyinput86, keyinput87,
         keyinput88, keyinput89, keyinput90, keyinput91, keyinput92,
         keyinput93, keyinput94, keyinput95, keyinput96, keyinput97,
         keyinput98, keyinput99, keyinput100, keyinput101, keyinput102,
         keyinput103, keyinput104, keyinput105, keyinput106, keyinput107,
         keyinput108, keyinput109, keyinput110, keyinput111, keyinput112,
         keyinput113, keyinput114, keyinput115, keyinput116, keyinput117,
         keyinput118, keyinput119, keyinput120, keyinput121, keyinput122,
         keyinput123, keyinput124, keyinput125, keyinput126, keyinput127;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488,
         n6489, n6490, n6491, n6492, n6494, n6495, n6496, n6497, n6498, n6499,
         n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509,
         n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519,
         n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529,
         n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539,
         n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549,
         n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559,
         n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569,
         n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579,
         n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589,
         n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599,
         n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609,
         n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619,
         n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629,
         n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639,
         n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649,
         n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659,
         n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669,
         n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6680,
         n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690,
         n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700,
         n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710,
         n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720,
         n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730,
         n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740,
         n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750,
         n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760,
         n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770,
         n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780,
         n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790,
         n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800,
         n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810,
         n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820,
         n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830,
         n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840,
         n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850,
         n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860,
         n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870,
         n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880,
         n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890,
         n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900,
         n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910,
         n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920,
         n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930,
         n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940,
         n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950,
         n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960,
         n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970,
         n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980,
         n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990,
         n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000,
         n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010,
         n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020,
         n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030,
         n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040,
         n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050,
         n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060,
         n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070,
         n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080,
         n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090,
         n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100,
         n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110,
         n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120,
         n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130,
         n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140,
         n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150,
         n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160,
         n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170,
         n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180,
         n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190,
         n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200,
         n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210,
         n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220,
         n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230,
         n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240,
         n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250,
         n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260,
         n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270,
         n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280,
         n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290,
         n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300,
         n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310,
         n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320,
         n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330,
         n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340,
         n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350,
         n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360,
         n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370,
         n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380,
         n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390,
         n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400,
         n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410,
         n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420,
         n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430,
         n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440,
         n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450,
         n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460,
         n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470,
         n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480,
         n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490,
         n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500,
         n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510,
         n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520,
         n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530,
         n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540,
         n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550,
         n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560,
         n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570,
         n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580,
         n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590,
         n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600,
         n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610,
         n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620,
         n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630,
         n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640,
         n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650,
         n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660,
         n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670,
         n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680,
         n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690,
         n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700,
         n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710,
         n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720,
         n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730,
         n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740,
         n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750,
         n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760,
         n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770,
         n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780,
         n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790,
         n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800,
         n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810,
         n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820,
         n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830,
         n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840,
         n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850,
         n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860,
         n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870,
         n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880,
         n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890,
         n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900,
         n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910,
         n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920,
         n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930,
         n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940,
         n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950,
         n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960,
         n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970,
         n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980,
         n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990,
         n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000,
         n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010,
         n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020,
         n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030,
         n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040,
         n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050,
         n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060,
         n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070,
         n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080,
         n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090,
         n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100,
         n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110,
         n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120,
         n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130,
         n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140,
         n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150,
         n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160,
         n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170,
         n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180,
         n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190,
         n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200,
         n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210,
         n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220,
         n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230,
         n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240,
         n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250,
         n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260,
         n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270,
         n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280,
         n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290,
         n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300,
         n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310,
         n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320,
         n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330,
         n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340,
         n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350,
         n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360,
         n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370,
         n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380,
         n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390,
         n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400,
         n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410,
         n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420,
         n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430,
         n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440,
         n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450,
         n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460,
         n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470,
         n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480,
         n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490,
         n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500,
         n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510,
         n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520,
         n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530,
         n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540,
         n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550,
         n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560,
         n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570,
         n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580,
         n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590,
         n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600,
         n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610,
         n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620,
         n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630,
         n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640,
         n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650,
         n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660,
         n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670,
         n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680,
         n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690,
         n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700,
         n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710,
         n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720,
         n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730,
         n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740,
         n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750,
         n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760,
         n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770,
         n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780,
         n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790,
         n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800,
         n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810,
         n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820,
         n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830,
         n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840,
         n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850,
         n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860,
         n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870,
         n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880,
         n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890,
         n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900,
         n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910,
         n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920,
         n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930,
         n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940,
         n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950,
         n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960,
         n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970,
         n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980,
         n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990,
         n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000,
         n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010,
         n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020,
         n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030,
         n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040,
         n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050,
         n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060,
         n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070,
         n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080,
         n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090,
         n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100,
         n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110,
         n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120,
         n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130,
         n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140,
         n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150,
         n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160,
         n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170,
         n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180,
         n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190,
         n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200,
         n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210,
         n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220,
         n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230,
         n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240,
         n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250,
         n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260,
         n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270,
         n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280,
         n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290,
         n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300,
         n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310,
         n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320,
         n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330,
         n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340,
         n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350,
         n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360,
         n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370,
         n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380,
         n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390,
         n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400,
         n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410,
         n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420,
         n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430,
         n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440,
         n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450,
         n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460,
         n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470,
         n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480,
         n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490,
         n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500,
         n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510,
         n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520,
         n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530,
         n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540,
         n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550,
         n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560,
         n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570,
         n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580,
         n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590,
         n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600,
         n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610,
         n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620,
         n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630,
         n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9639, n9640, n9641,
         n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651,
         n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661,
         n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671,
         n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681,
         n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691,
         n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701,
         n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711,
         n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721,
         n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731,
         n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741,
         n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751,
         n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761,
         n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771,
         n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781,
         n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791,
         n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801,
         n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811,
         n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821,
         n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831,
         n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841,
         n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851,
         n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861,
         n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871,
         n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881,
         n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891,
         n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901,
         n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911,
         n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921,
         n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931,
         n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941,
         n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951,
         n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961,
         n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971,
         n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981,
         n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991,
         n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
         n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
         n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296,
         n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304,
         n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
         n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320,
         n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328,
         n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336,
         n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344,
         n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352,
         n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360,
         n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368,
         n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376,
         n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384,
         n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392,
         n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400,
         n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408,
         n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416,
         n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424,
         n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432,
         n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440,
         n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448,
         n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456,
         n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464,
         n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472,
         n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480,
         n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488,
         n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496,
         n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504,
         n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512,
         n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520,
         n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528,
         n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536,
         n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544,
         n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552,
         n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560,
         n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568,
         n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576,
         n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584,
         n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592,
         n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600,
         n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608,
         n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616,
         n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624,
         n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632,
         n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640,
         n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648,
         n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656,
         n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10664,
         n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672,
         n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10680,
         n10681, n10682, n10683, n10684, n10685, n10686, n10687, n10688,
         n10689, n10690, n10691, n10692, n10693, n10694, n10695, n10696,
         n10697, n10698, n10699, n10700, n10701, n10702, n10703, n10704,
         n10705, n10706, n10707, n10708, n10709, n10710, n10711, n10712,
         n10713, n10714, n10715, n10716, n10717, n10718, n10719, n10720,
         n10721, n10722, n10723, n10724, n10725, n10726, n10727, n10728,
         n10729, n10730, n10731, n10732, n10733, n10734, n10735, n10736,
         n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10744,
         n10745, n10746, n10747, n10748, n10749, n10750, n10751, n10752,
         n10753, n10754, n10755, n10756, n10757, n10758, n10759, n10760,
         n10761, n10762, n10763, n10764, n10765, n10766, n10767, n10768,
         n10769, n10770, n10771, n10772, n10773, n10774, n10775, n10776,
         n10777, n10778, n10779, n10780, n10781, n10782, n10783, n10784,
         n10785, n10786, n10787, n10788, n10789, n10790, n10791, n10792,
         n10793, n10794, n10795, n10796, n10797, n10798, n10799, n10800,
         n10801, n10802, n10803, n10804, n10805, n10806, n10807, n10808,
         n10809, n10810, n10811, n10812, n10813, n10814, n10815, n10816,
         n10817, n10818, n10819, n10820, n10821, n10822, n10823, n10824,
         n10825, n10826, n10827, n10828, n10829, n10830, n10831, n10832,
         n10833, n10834, n10835, n10836, n10837, n10838, n10839, n10840,
         n10841, n10842, n10843, n10844, n10845, n10846, n10847, n10848,
         n10849, n10850, n10851, n10852, n10853, n10854, n10855, n10856,
         n10857, n10858, n10859, n10860, n10861, n10862, n10863, n10864,
         n10865, n10866, n10867, n10868, n10869, n10870, n10871, n10872,
         n10873, n10874, n10875, n10876, n10877, n10878, n10879, n10880,
         n10881, n10882, n10883, n10884, n10885, n10886, n10887, n10888,
         n10889, n10890, n10891, n10892, n10893, n10894, n10895, n10896,
         n10897, n10898, n10899, n10900, n10901, n10902, n10903, n10904,
         n10905, n10906, n10907, n10908, n10909, n10910, n10911, n10912,
         n10913, n10914, n10915, n10916, n10917, n10918, n10919, n10920,
         n10921, n10922, n10923, n10924, n10925, n10926, n10927, n10928,
         n10929, n10930, n10931, n10932, n10933, n10934, n10935, n10936,
         n10937, n10938, n10939, n10940, n10941, n10942, n10943, n10944,
         n10945, n10946, n10947, n10948, n10949, n10950, n10951, n10952,
         n10953, n10954, n10955, n10956, n10957, n10958, n10959, n10960,
         n10961, n10962, n10963, n10964, n10965, n10966, n10967, n10968,
         n10969, n10970, n10971, n10972, n10973, n10974, n10975, n10976,
         n10977, n10978, n10979, n10980, n10981, n10982, n10983, n10984,
         n10985, n10986, n10987, n10988, n10989, n10990, n10991, n10992,
         n10993, n10994, n10995, n10996, n10997, n10998, n10999, n11000,
         n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008,
         n11009, n11010, n11011, n11012, n11013, n11014, n11015, n11016,
         n11017, n11018, n11019, n11020, n11021, n11022, n11023, n11024,
         n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11032,
         n11033, n11034, n11035, n11036, n11037, n11038, n11039, n11040,
         n11041, n11042, n11043, n11044, n11045, n11046, n11047, n11048,
         n11049, n11050, n11051, n11052, n11053, n11054, n11055, n11056,
         n11057, n11058, n11059, n11060, n11061, n11062, n11063, n11064,
         n11065, n11066, n11067, n11068, n11069, n11070, n11071, n11072,
         n11073, n11074, n11075, n11076, n11077, n11078, n11079, n11080,
         n11081, n11082, n11083, n11084, n11085, n11086, n11087, n11088,
         n11089, n11090, n11091, n11092, n11093, n11094, n11095, n11096,
         n11097, n11098, n11099, n11100, n11101, n11102, n11103, n11104,
         n11105, n11106, n11107, n11108, n11109, n11110, n11111, n11112,
         n11113, n11114, n11115, n11116, n11117, n11118, n11119, n11120,
         n11121, n11122, n11123, n11124, n11125, n11126, n11127, n11128,
         n11129, n11130, n11131, n11132, n11133, n11134, n11135, n11136,
         n11137, n11138, n11139, n11140, n11141, n11142, n11143, n11144,
         n11145, n11146, n11147, n11148, n11149, n11150, n11151, n11152,
         n11153, n11154, n11155, n11156, n11157, n11158, n11159, n11160,
         n11161, n11162, n11163, n11164, n11165, n11166, n11167, n11168,
         n11169, n11170, n11171, n11172, n11173, n11174, n11175, n11176,
         n11177, n11178, n11179, n11180, n11181, n11182, n11183, n11184,
         n11185, n11186, n11187, n11188, n11189, n11190, n11191, n11192,
         n11193, n11194, n11195, n11196, n11197, n11198, n11199, n11200,
         n11201, n11202, n11203, n11204, n11205, n11206, n11207, n11208,
         n11209, n11210, n11211, n11212, n11213, n11214, n11215, n11216,
         n11217, n11218, n11219, n11220, n11221, n11222, n11223, n11224,
         n11225, n11226, n11227, n11228, n11229, n11230, n11231, n11232,
         n11233, n11234, n11235, n11236, n11237, n11238, n11239, n11240,
         n11241, n11242, n11243, n11244, n11245, n11246, n11247, n11248,
         n11249, n11250, n11251, n11252, n11253, n11254, n11255, n11256,
         n11257, n11258, n11259, n11260, n11261, n11262, n11263, n11264,
         n11265, n11266, n11267, n11268, n11269, n11270, n11271, n11272,
         n11273, n11274, n11275, n11276, n11277, n11278, n11279, n11280,
         n11281, n11282, n11283, n11284, n11285, n11286, n11287, n11288,
         n11289, n11290, n11291, n11292, n11293, n11294, n11295, n11296,
         n11297, n11298, n11299, n11300, n11301, n11302, n11303, n11304,
         n11305, n11306, n11307, n11308, n11309, n11310, n11311, n11312,
         n11313, n11314, n11315, n11316, n11317, n11318, n11319, n11320,
         n11321, n11322, n11323, n11324, n11325, n11326, n11327, n11328,
         n11329, n11330, n11331, n11332, n11333, n11334, n11335, n11336,
         n11337, n11338, n11339, n11340, n11341, n11342, n11343, n11344,
         n11345, n11346, n11347, n11348, n11349, n11350, n11351, n11352,
         n11353, n11354, n11355, n11356, n11357, n11358, n11359, n11360,
         n11361, n11362, n11363, n11364, n11365, n11366, n11367, n11368,
         n11369, n11370, n11371, n11372, n11373, n11374, n11375, n11376,
         n11377, n11378, n11379, n11380, n11381, n11382, n11383, n11384,
         n11385, n11386, n11387, n11388, n11389, n11390, n11391, n11392,
         n11393, n11394, n11395, n11396, n11397, n11398, n11399, n11400,
         n11401, n11402, n11403, n11404, n11405, n11406, n11407, n11408,
         n11409, n11410, n11411, n11412, n11413, n11414, n11415, n11416,
         n11417, n11418, n11419, n11420, n11421, n11422, n11423, n11424,
         n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432,
         n11433, n11434, n11435, n11436, n11437, n11438, n11439, n11440,
         n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448,
         n11449, n11450, n11451, n11452, n11453, n11454, n11455, n11456,
         n11457, n11458, n11459, n11460, n11461, n11462, n11463, n11464,
         n11465, n11466, n11467, n11468, n11469, n11470, n11471, n11472,
         n11473, n11474, n11475, n11476, n11477, n11478, n11479, n11480,
         n11481, n11482, n11483, n11484, n11485, n11486, n11487, n11488,
         n11489, n11490, n11491, n11492, n11493, n11494, n11495, n11496,
         n11497, n11498, n11499, n11500, n11501, n11502, n11503, n11504,
         n11505, n11506, n11507, n11508, n11509, n11510, n11511, n11512,
         n11513, n11514, n11515, n11516, n11517, n11518, n11519, n11520,
         n11521, n11522, n11523, n11524, n11525, n11526, n11527, n11528,
         n11529, n11530, n11531, n11532, n11533, n11534, n11535, n11536,
         n11537, n11538, n11539, n11540, n11541, n11542, n11543, n11544,
         n11545, n11546, n11547, n11548, n11549, n11550, n11551, n11552,
         n11553, n11554, n11555, n11556, n11557, n11558, n11559, n11560,
         n11561, n11562, n11563, n11564, n11565, n11566, n11567, n11568,
         n11569, n11570, n11571, n11572, n11573, n11574, n11575, n11576,
         n11577, n11578, n11579, n11580, n11581, n11582, n11583, n11584,
         n11585, n11586, n11587, n11588, n11589, n11590, n11591, n11592,
         n11593, n11594, n11595, n11596, n11597, n11598, n11599, n11600,
         n11601, n11602, n11603, n11604, n11605, n11606, n11607, n11608,
         n11609, n11610, n11611, n11612, n11613, n11614, n11615, n11616,
         n11617, n11618, n11619, n11620, n11621, n11622, n11623, n11624,
         n11625, n11626, n11627, n11628, n11629, n11630, n11631, n11632,
         n11633, n11634, n11635, n11636, n11637, n11638, n11639, n11640,
         n11641, n11642, n11643, n11644, n11645, n11646, n11647, n11648,
         n11649, n11650, n11651, n11652, n11653, n11654, n11655, n11656,
         n11657, n11658, n11659, n11660, n11661, n11662, n11663, n11664,
         n11665, n11666, n11667, n11668, n11669, n11670, n11671, n11672,
         n11673, n11674, n11675, n11676, n11677, n11678, n11679, n11680,
         n11681, n11682, n11683, n11684, n11685, n11686, n11687, n11688,
         n11689, n11690, n11691, n11692, n11693, n11694, n11695, n11696,
         n11697, n11698, n11699, n11700, n11701, n11702, n11703, n11704,
         n11705, n11706, n11707, n11708, n11709, n11710, n11711, n11712,
         n11713, n11714, n11715, n11716, n11717, n11718, n11719, n11720,
         n11721, n11722, n11723, n11724, n11725, n11726, n11727, n11728,
         n11729, n11730, n11731, n11732, n11733, n11734, n11735, n11736,
         n11737, n11738, n11739, n11740, n11741, n11742, n11743, n11744,
         n11745, n11746, n11747, n11748, n11749, n11750, n11751, n11752,
         n11753, n11754, n11755, n11756, n11757, n11758, n11759, n11760,
         n11761, n11762, n11763, n11764, n11765, n11766, n11767, n11768,
         n11769, n11770, n11771, n11772, n11773, n11774, n11775, n11776,
         n11777, n11778, n11779, n11780, n11781, n11782, n11783, n11784,
         n11785, n11786, n11787, n11788, n11789, n11790, n11791, n11792,
         n11793, n11794, n11795, n11796, n11797, n11798, n11799, n11800,
         n11801, n11802, n11803, n11804, n11805, n11806, n11807, n11808,
         n11809, n11810, n11811, n11812, n11813, n11814, n11815, n11816,
         n11817, n11818, n11819, n11820, n11821, n11822, n11823, n11824,
         n11825, n11826, n11827, n11828, n11829, n11830, n11831, n11832,
         n11833, n11834, n11835, n11836, n11837, n11838, n11839, n11840,
         n11841, n11842, n11843, n11844, n11845, n11846, n11847, n11848,
         n11849, n11850, n11851, n11852, n11853, n11854, n11855, n11856,
         n11857, n11858, n11859, n11860, n11861, n11862, n11863, n11864,
         n11865, n11866, n11867, n11868, n11869, n11870, n11871, n11872,
         n11873, n11874, n11875, n11876, n11877, n11878, n11879, n11880,
         n11881, n11882, n11883, n11884, n11885, n11886, n11887, n11888,
         n11889, n11890, n11891, n11892, n11893, n11894, n11895, n11896,
         n11897, n11898, n11899, n11900, n11901, n11902, n11903, n11904,
         n11905, n11906, n11907, n11908, n11909, n11910, n11911, n11912,
         n11913, n11914, n11915, n11916, n11917, n11918, n11919, n11920,
         n11921, n11922, n11923, n11924, n11925, n11926, n11927, n11928,
         n11929, n11930, n11931, n11932, n11933, n11934, n11935, n11936,
         n11937, n11938, n11939, n11940, n11941, n11942, n11943, n11944,
         n11945, n11946, n11947, n11948, n11949, n11950, n11951, n11952,
         n11953, n11954, n11955, n11956, n11957, n11958, n11959, n11960,
         n11961, n11962, n11963, n11964, n11965, n11966, n11967, n11968,
         n11969, n11970, n11971, n11972, n11973, n11974, n11975, n11976,
         n11977, n11978, n11979, n11980, n11981, n11982, n11983, n11984,
         n11985, n11986, n11987, n11988, n11989, n11990, n11991, n11992,
         n11993, n11994, n11995, n11996, n11997, n11998, n11999, n12000,
         n12001, n12002, n12003, n12004, n12005, n12006, n12007, n12008,
         n12009, n12010, n12011, n12012, n12013, n12014, n12015, n12016,
         n12017, n12018, n12019, n12020, n12021, n12022, n12023, n12024,
         n12025, n12026, n12027, n12028, n12029, n12030, n12031, n12032,
         n12033, n12034, n12035, n12036, n12037, n12038, n12039, n12040,
         n12041, n12042, n12043, n12044, n12045, n12046, n12047, n12048,
         n12049, n12050, n12051, n12052, n12053, n12054, n12055, n12056,
         n12057, n12058, n12059, n12060, n12061, n12062, n12063, n12064,
         n12065, n12066, n12067, n12068, n12069, n12070, n12071, n12072,
         n12073, n12074, n12075, n12076, n12077, n12078, n12079, n12080,
         n12081, n12082, n12083, n12084, n12085, n12086, n12087, n12088,
         n12089, n12090, n12091, n12092, n12093, n12094, n12095, n12096,
         n12097, n12098, n12099, n12100, n12101, n12102, n12103, n12104,
         n12105, n12106, n12107, n12108, n12109, n12110, n12111, n12112,
         n12113, n12114, n12115, n12116, n12117, n12119, n12120, n12121,
         n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129,
         n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137,
         n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145,
         n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153,
         n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161,
         n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169,
         n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177,
         n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185,
         n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193,
         n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201,
         n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209,
         n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217,
         n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225,
         n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233,
         n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241,
         n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249,
         n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257,
         n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265,
         n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273,
         n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281,
         n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289,
         n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297,
         n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305,
         n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313,
         n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321,
         n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329,
         n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337,
         n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345,
         n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353,
         n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361,
         n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369,
         n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377,
         n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385,
         n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393,
         n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401,
         n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409,
         n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417,
         n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425,
         n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433,
         n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441,
         n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449,
         n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457,
         n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465,
         n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473,
         n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481,
         n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489,
         n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497,
         n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505,
         n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513,
         n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521,
         n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529,
         n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537,
         n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545,
         n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553,
         n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561,
         n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569,
         n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577,
         n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585,
         n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593,
         n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601,
         n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609,
         n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617,
         n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625,
         n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633,
         n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641,
         n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649,
         n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657,
         n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665,
         n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673,
         n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681,
         n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689,
         n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697,
         n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705,
         n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713,
         n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721,
         n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729,
         n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737,
         n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745,
         n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753,
         n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761,
         n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769,
         n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777,
         n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785,
         n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793,
         n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801,
         n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809,
         n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817,
         n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825,
         n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833,
         n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841,
         n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849,
         n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857,
         n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865,
         n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873,
         n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881,
         n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889,
         n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897,
         n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905,
         n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913,
         n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921,
         n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929,
         n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937,
         n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945,
         n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953,
         n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961,
         n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969,
         n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977,
         n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985,
         n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993,
         n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001,
         n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009,
         n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017,
         n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025,
         n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033,
         n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041,
         n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049,
         n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057,
         n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065,
         n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073,
         n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081,
         n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089,
         n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097,
         n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105,
         n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113,
         n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121,
         n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129,
         n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137,
         n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145,
         n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153,
         n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161,
         n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169,
         n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177,
         n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185,
         n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193,
         n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201,
         n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209,
         n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217,
         n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225,
         n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233,
         n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241,
         n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249,
         n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257,
         n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265,
         n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273,
         n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281,
         n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289,
         n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297,
         n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305,
         n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313,
         n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321,
         n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329,
         n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337,
         n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345,
         n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353,
         n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361,
         n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369,
         n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377,
         n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385,
         n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393,
         n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401,
         n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409,
         n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417,
         n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425,
         n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433,
         n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441,
         n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449,
         n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457,
         n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465,
         n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473,
         n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481,
         n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489,
         n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497,
         n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505,
         n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513,
         n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521,
         n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529,
         n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537,
         n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545,
         n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553,
         n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561,
         n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569,
         n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577,
         n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585,
         n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593,
         n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601,
         n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609,
         n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617,
         n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625,
         n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633,
         n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641,
         n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649,
         n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657,
         n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665,
         n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673,
         n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681,
         n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689,
         n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697,
         n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705,
         n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713,
         n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721,
         n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729,
         n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737,
         n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745,
         n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753,
         n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761,
         n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769,
         n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777,
         n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785,
         n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793,
         n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801,
         n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809,
         n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817,
         n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825,
         n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833,
         n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841,
         n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849,
         n13850, n13851, n13852, n13853, n13854, n13855, n13856, n13857,
         n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865,
         n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873,
         n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881,
         n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889,
         n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897,
         n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905,
         n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913,
         n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921,
         n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929,
         n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937,
         n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945,
         n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953,
         n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961,
         n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969,
         n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977,
         n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985,
         n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993,
         n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001,
         n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009,
         n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017,
         n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025,
         n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033,
         n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041,
         n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049,
         n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057,
         n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065,
         n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073,
         n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081,
         n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089,
         n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097,
         n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105,
         n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113,
         n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121,
         n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129,
         n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137,
         n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145,
         n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153,
         n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161,
         n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169,
         n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177,
         n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185,
         n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193,
         n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201,
         n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209,
         n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217,
         n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225,
         n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233,
         n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241,
         n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249,
         n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257,
         n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265,
         n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273,
         n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281,
         n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289,
         n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297,
         n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305,
         n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313,
         n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321,
         n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329,
         n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337,
         n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345,
         n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353,
         n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361,
         n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369,
         n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377,
         n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385,
         n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393,
         n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401,
         n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409,
         n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417,
         n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425,
         n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433,
         n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441,
         n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449,
         n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457,
         n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465,
         n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473,
         n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14482,
         n14483, n14484, n14485, n14486, n14487, n14488, n14489, n14490,
         n14491, n14492, n14493, n14494, n14495, n14496, n14497, n14498,
         n14499, n14500, n14501, n14502, n14503, n14504, n14505, n14506,
         n14507, n14508, n14509, n14510, n14511, n14512, n14513, n14514,
         n14515, n14516, n14517, n14518, n14519, n14520, n14521, n14522,
         n14523, n14524, n14525, n14526, n14527, n14528, n14529, n14530,
         n14531, n14532, n14533, n14534, n14535, n14536, n14537, n14538,
         n14539, n14540, n14541, n14542, n14543, n14544, n14545, n14546,
         n14547, n14548, n14549, n14550, n14551, n14552, n14553, n14554,
         n14555, n14556, n14557, n14558, n14559, n14560, n14561, n14562,
         n14563, n14564, n14565, n14566, n14567, n14568, n14569, n14570,
         n14571, n14572, n14573, n14574, n14575, n14576, n14577, n14578,
         n14579, n14580, n14581, n14582, n14583, n14584, n14585, n14586,
         n14587, n14588, n14589, n14590, n14591, n14592, n14593, n14594,
         n14595, n14596, n14597, n14598, n14599, n14600, n14601, n14602,
         n14603, n14604, n14605, n14606, n14607, n14608, n14609, n14610,
         n14611, n14612, n14613, n14614, n14615, n14616, n14617, n14618,
         n14619, n14620, n14621, n14622, n14623, n14624, n14625, n14626,
         n14627, n14628, n14629, n14630, n14631, n14632, n14633, n14634,
         n14635, n14636, n14637, n14638, n14639, n14640, n14641, n14642,
         n14643, n14644, n14645, n14646, n14647, n14648, n14649, n14650,
         n14651, n14652, n14653, n14654, n14655, n14656, n14657, n14658,
         n14659, n14660, n14661, n14662, n14663, n14664, n14665, n14666,
         n14667, n14668, n14669, n14670, n14671, n14672, n14673, n14674,
         n14675, n14676, n14677, n14678, n14679, n14680, n14681, n14682,
         n14683, n14684, n14685, n14686, n14687, n14688, n14689, n14690,
         n14691, n14692, n14693, n14694, n14695, n14696, n14697, n14698,
         n14699, n14700, n14701, n14702, n14703, n14704, n14705, n14706,
         n14707, n14708, n14709, n14710, n14711, n14712, n14713, n14714,
         n14715, n14716, n14717, n14718, n14719, n14720, n14721, n14722,
         n14723, n14724, n14725, n14726, n14727, n14728, n14729, n14730,
         n14731, n14732, n14733, n14734, n14735, n14736, n14737, n14738,
         n14739, n14740, n14741, n14742, n14743, n14744, n14745, n14746,
         n14747, n14748, n14749, n14750, n14751, n14752, n14753, n14754,
         n14755, n14756, n14757, n14758, n14759, n14760, n14761, n14762,
         n14763, n14764, n14765, n14766, n14767, n14768, n14769, n14770,
         n14771, n14772, n14773, n14774, n14775, n14776, n14777, n14778,
         n14779, n14780, n14781, n14782, n14783, n14784, n14785, n14786,
         n14787, n14788, n14789, n14790, n14791, n14792, n14793, n14794,
         n14795, n14796, n14797, n14798, n14799, n14800, n14801, n14802,
         n14803, n14804, n14805, n14806, n14807, n14808, n14809, n14810,
         n14811, n14812, n14813, n14814, n14815, n14816, n14817, n14818,
         n14819, n14820, n14821, n14822, n14823, n14824, n14825, n14826,
         n14827, n14828, n14829, n14830, n14831, n14832, n14833, n14834,
         n14835, n14836, n14837, n14838, n14839, n14840, n14841, n14842,
         n14843, n14844, n14845, n14846, n14847, n14848, n14849, n14850,
         n14851, n14852, n14853, n14854, n14855, n14856, n14857, n14858,
         n14859, n14860, n14861, n14862, n14863, n14864, n14865, n14866,
         n14867, n14868, n14869, n14870, n14871, n14872, n14873, n14874,
         n14875, n14876, n14877, n14878, n14879, n14880, n14881, n14882,
         n14883, n14884, n14885, n14886, n14887, n14888, n14889, n14890,
         n14891, n14892, n14893, n14894, n14895, n14896, n14897, n14898,
         n14899, n14900, n14901, n14902, n14903, n14904, n14905, n14906,
         n14907, n14908, n14909, n14910, n14911, n14912, n14913, n14914,
         n14915, n14916, n14917, n14918, n14919, n14920, n14921, n14922,
         n14923, n14924, n14925, n14926, n14927, n14928, n14929, n14930,
         n14931, n14932, n14933, n14934, n14935, n14936, n14937, n14938,
         n14939, n14940, n14941, n14942, n14943, n14944, n14945, n14946,
         n14947, n14948, n14949, n14950, n14951, n14952, n14953, n14954,
         n14955, n14956, n14957, n14958, n14959, n14960, n14961, n14962,
         n14963, n14964, n14965, n14966, n14967, n14968, n14969, n14970,
         n14971, n14972, n14973, n14974, n14975, n14976, n14977, n14978,
         n14979, n14980, n14981, n14982, n14983, n14984, n14985, n14986,
         n14987, n14988, n14989, n14990, n14991, n14992, n14993, n14994,
         n14995, n14996, n14997, n14998, n14999, n15000, n15001, n15002,
         n15003, n15004, n15005, n15006, n15007, n15008, n15009, n15010,
         n15011, n15012, n15013, n15014, n15015, n15016, n15017, n15018,
         n15019, n15020, n15021, n15022, n15023, n15024, n15025, n15026,
         n15027, n15028, n15029, n15030, n15031, n15032, n15033, n15034,
         n15035, n15036, n15037, n15038, n15039, n15040, n15041, n15042,
         n15043, n15044, n15045, n15046, n15047, n15048, n15049, n15050,
         n15051, n15052, n15053, n15054, n15055, n15056, n15057, n15058,
         n15059, n15060, n15061, n15062, n15063, n15064, n15065, n15066,
         n15067, n15068, n15069, n15070, n15071, n15072, n15073, n15074,
         n15075, n15076, n15077, n15078, n15079, n15080, n15081, n15082,
         n15083, n15084, n15085, n15086, n15087, n15088, n15089, n15090,
         n15091, n15092, n15093, n15094, n15095, n15096, n15097, n15098,
         n15099, n15100, n15101, n15102, n15103, n15104, n15105, n15106,
         n15107, n15108, n15109, n15110, n15111, n15112, n15113, n15114,
         n15115, n15116, n15117, n15118, n15119, n15120, n15121, n15122,
         n15123, n15124, n15125, n15126, n15127, n15128, n15129, n15130,
         n15131, n15132, n15133, n15134, n15135, n15136, n15137, n15138,
         n15139, n15140, n15141, n15142, n15143, n15144, n15145, n15146,
         n15147, n15148, n15149, n15150, n15151, n15152, n15153, n15154,
         n15155, n15156, n15157, n15158, n15159, n15160, n15161, n15162,
         n15163, n15164, n15165, n15166, n15167, n15168, n15169, n15170,
         n15171, n15172, n15173, n15174, n15175, n15176, n15177, n15178,
         n15179, n15180, n15181, n15182, n15183, n15184, n15185, n15186,
         n15187, n15188, n15189, n15190, n15191, n15192, n15193, n15194,
         n15195, n15196, n15197, n15198, n15199, n15200, n15201, n15202,
         n15203, n15204, n15205, n15206, n15207, n15208, n15209, n15210,
         n15211, n15212, n15213, n15214, n15215, n15216, n15217, n15218,
         n15219, n15220, n15221, n15222, n15223, n15224, n15225, n15226,
         n15227, n15228, n15229, n15230, n15231, n15232, n15233, n15234,
         n15235, n15236, n15237, n15238, n15239, n15240, n15241, n15242,
         n15243, n15244, n15245, n15246, n15247, n15248, n15249, n15250,
         n15251, n15252, n15253, n15254, n15255, n15256, n15257, n15258,
         n15259, n15260, n15261, n15262, n15263, n15264, n15265, n15266,
         n15267, n15268, n15269, n15270, n15271, n15272, n15273, n15274,
         n15275, n15276, n15277, n15278, n15279, n15280, n15281, n15282,
         n15283, n15284, n15285, n15286, n15287, n15288, n15289, n15290,
         n15291, n15292, n15293, n15294;

  OAI222_X1 U7227 ( .A1(n13873), .A2(n13868), .B1(P2_U3088), .B2(n13867), .C1(
        n13866), .C2(n13870), .ZN(P2_U3297) );
  INV_X1 U7228 ( .A(n6479), .ZN(n11246) );
  NAND2_X1 U7229 ( .A1(n9143), .A2(n9142), .ZN(n13779) );
  NAND2_X1 U7230 ( .A1(n13400), .A2(n7439), .ZN(n12592) );
  OR2_X1 U7231 ( .A1(n12778), .A2(n6727), .ZN(n6726) );
  OR2_X1 U7232 ( .A1(n13011), .A2(n13010), .ZN(n13013) );
  NAND2_X1 U7233 ( .A1(n13021), .A2(n12306), .ZN(n13003) );
  NAND2_X1 U7234 ( .A1(n12840), .A2(n12839), .ZN(n13038) );
  AND2_X1 U7235 ( .A1(n6806), .A2(n6805), .ZN(n11461) );
  NAND2_X1 U7236 ( .A1(n7010), .A2(n7013), .ZN(n11987) );
  NAND2_X1 U7237 ( .A1(n7122), .A2(n14555), .ZN(n14558) );
  NAND2_X1 U7238 ( .A1(n11527), .A2(n12418), .ZN(n11692) );
  NAND2_X1 U7239 ( .A1(n10805), .A2(n10806), .ZN(n11113) );
  AND2_X1 U7240 ( .A1(n7334), .A2(n7333), .ZN(n11311) );
  BUF_X1 U7241 ( .A(n10389), .Z(n12611) );
  INV_X2 U7242 ( .A(n12481), .ZN(n11001) );
  NAND2_X1 U7243 ( .A1(n7284), .A2(n7283), .ZN(n7836) );
  INV_X2 U7244 ( .A(n12605), .ZN(n10086) );
  INV_X2 U7245 ( .A(n10560), .ZN(n12292) );
  OR2_X1 U7246 ( .A1(n8314), .A2(n8325), .ZN(n11878) );
  NAND2_X1 U7247 ( .A1(n6993), .A2(n10297), .ZN(n12375) );
  OAI22_X1 U7248 ( .A1(n9636), .A2(n9635), .B1(P2_DATAO_REG_9__SCAN_IN), .B2(
        n9651), .ZN(n9641) );
  AND4_X1 U7249 ( .A1(n10292), .A2(n10291), .A3(n10290), .A4(n10289), .ZN(
        n10993) );
  OR2_X1 U7250 ( .A1(n14046), .A2(n9548), .ZN(n6684) );
  XNOR2_X1 U7251 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .ZN(n9592) );
  AND2_X1 U7252 ( .A1(n12628), .A2(n7480), .ZN(n8200) );
  INV_X1 U7253 ( .A(n12108), .ZN(n9502) );
  CLKBUF_X2 U7254 ( .A(n7527), .Z(n9667) );
  INV_X1 U7255 ( .A(n9582), .ZN(n8621) );
  BUF_X1 U7256 ( .A(n7670), .Z(n7671) );
  NAND2_X1 U7257 ( .A1(n6842), .A2(n6839), .ZN(n9582) );
  NAND2_X1 U7258 ( .A1(n6843), .A2(P3_ADDR_REG_19__SCAN_IN), .ZN(n6842) );
  NOR2_X1 U7259 ( .A1(P2_IR_REG_14__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), .ZN(
        n8559) );
  AND2_X2 U7260 ( .A1(n10957), .A2(n10956), .ZN(n6479) );
  NOR2_X1 U7261 ( .A1(n10332), .A2(n7444), .ZN(n9297) );
  AOI21_X2 U7262 ( .B1(n10465), .B2(n10464), .A(n7151), .ZN(n10579) );
  NAND2_X2 U7263 ( .A1(n12951), .A2(n12950), .ZN(n12953) );
  XNOR2_X1 U7265 ( .A(n14582), .B(n14581), .ZN(n14782) );
  NAND2_X1 U7266 ( .A1(n11313), .A2(n11312), .ZN(n6481) );
  AOI21_X1 U7267 ( .B1(n12949), .B2(n12852), .A(n12851), .ZN(n6482) );
  AOI21_X1 U7268 ( .B1(n12949), .B2(n12852), .A(n12851), .ZN(n12940) );
  INV_X4 U7269 ( .A(n8215), .ZN(n8176) );
  NOR2_X1 U7270 ( .A1(n10413), .A2(n8468), .ZN(n8469) );
  NOR2_X1 U7271 ( .A1(P3_IR_REG_10__SCAN_IN), .A2(P3_IR_REG_11__SCAN_IN), .ZN(
        n8302) );
  NOR2_X1 U7272 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n8558) );
  INV_X1 U7273 ( .A(n8176), .ZN(n8150) );
  NOR2_X1 U7274 ( .A1(P3_IR_REG_5__SCAN_IN), .A2(P3_IR_REG_4__SCAN_IN), .ZN(
        n8407) );
  NAND2_X1 U7275 ( .A1(n6876), .A2(n6503), .ZN(n7117) );
  NAND2_X1 U7276 ( .A1(n7166), .A2(n10296), .ZN(n10560) );
  NOR2_X1 U7277 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), .ZN(
        n8353) );
  XNOR2_X1 U7278 ( .A(n6726), .B(n6725), .ZN(n14629) );
  AND3_X1 U7279 ( .A1(n10926), .A2(n10925), .A3(n10924), .ZN(n11020) );
  NAND2_X1 U7280 ( .A1(n8638), .A2(n10187), .ZN(n8678) );
  OR2_X1 U7281 ( .A1(n13605), .A2(n13604), .ZN(n6729) );
  INV_X1 U7282 ( .A(n9287), .ZN(n12057) );
  INV_X1 U7283 ( .A(n9287), .ZN(n12066) );
  INV_X1 U7284 ( .A(n10503), .ZN(n10509) );
  BUF_X1 U7285 ( .A(n10993), .Z(n15198) );
  NAND2_X1 U7286 ( .A1(n9920), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9921) );
  NAND2_X1 U7287 ( .A1(n9055), .A2(n9054), .ZN(n13795) );
  OR2_X1 U7288 ( .A1(n13642), .A2(n6942), .ZN(n13606) );
  AOI21_X1 U7289 ( .B1(n7394), .B2(n6748), .A(n6573), .ZN(n11547) );
  CLKBUF_X3 U7290 ( .A(n8200), .Z(n8137) );
  OR2_X1 U7291 ( .A1(n14136), .A2(n12555), .ZN(n12082) );
  NAND2_X1 U7292 ( .A1(n9506), .A2(n7569), .ZN(n10503) );
  NAND2_X1 U7293 ( .A1(n8647), .A2(n8646), .ZN(n10769) );
  NOR2_X1 U7294 ( .A1(n10333), .A2(n10334), .ZN(n10332) );
  XNOR2_X1 U7295 ( .A(n7953), .B(n7952), .ZN(n8963) );
  XNOR2_X1 U7297 ( .A(n7171), .B(n8307), .ZN(n9808) );
  NAND3_X1 U7298 ( .A1(n6733), .A2(n8567), .A3(n6732), .ZN(n13872) );
  XOR2_X1 U7299 ( .A(n14538), .B(P2_ADDR_REG_1__SCAN_IN), .Z(n15293) );
  INV_X1 U7300 ( .A(n10449), .ZN(n12165) );
  MUX2_X1 U7301 ( .A(P2_IR_REG_0__SCAN_IN), .B(n13874), .S(n8638), .Z(n14990)
         );
  NOR2_X2 U7303 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .ZN(
        n7371) );
  INV_X1 U7305 ( .A(n8678), .ZN(n9168) );
  AND2_X2 U7306 ( .A1(n8569), .A2(n13872), .ZN(n8683) );
  OAI21_X1 U7307 ( .B1(n13666), .B2(n7307), .A(n7304), .ZN(n7311) );
  NAND2_X2 U7308 ( .A1(n13683), .A2(n7295), .ZN(n13670) );
  NAND2_X1 U7309 ( .A1(n6842), .A2(n6839), .ZN(n6484) );
  AOI21_X2 U7310 ( .B1(n12810), .B2(n12809), .A(n12808), .ZN(n12812) );
  NAND3_X2 U7311 ( .A1(n6973), .A2(n6971), .A3(n6972), .ZN(n12810) );
  OAI21_X2 U7312 ( .B1(n14545), .B2(n9767), .A(n15289), .ZN(n15282) );
  XNOR2_X1 U7313 ( .A(n8464), .B(n8463), .ZN(n8510) );
  NAND2_X1 U7314 ( .A1(n7166), .A2(n10296), .ZN(n6486) );
  INV_X2 U7315 ( .A(n12292), .ZN(n12151) );
  CLKBUF_X1 U7316 ( .A(n12328), .Z(n6487) );
  NAND2_X1 U7317 ( .A1(n9922), .A2(n12119), .ZN(n12328) );
  INV_X2 U7318 ( .A(n9667), .ZN(n6753) );
  AOI22_X2 U7319 ( .A1(n10450), .A2(P3_REG2_REG_2__SCAN_IN), .B1(n8352), .B2(
        n6496), .ZN(n10418) );
  BUF_X2 U7320 ( .A(n8357), .Z(n6496) );
  NAND2_X2 U7321 ( .A1(n8567), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8566) );
  AOI21_X2 U7322 ( .B1(P3_REG1_REG_4__SCAN_IN), .B2(n9597), .A(n15112), .ZN(
        n8472) );
  NAND2_X2 U7323 ( .A1(n13867), .A2(n8568), .ZN(n6932) );
  XNOR2_X2 U7324 ( .A(n12592), .B(n12591), .ZN(n13343) );
  INV_X2 U7325 ( .A(n9230), .ZN(n8663) );
  INV_X2 U7326 ( .A(n9230), .ZN(n9035) );
  OR2_X1 U7327 ( .A1(n15026), .A2(n9230), .ZN(n8626) );
  AOI22_X2 U7328 ( .A1(n10867), .A2(n10866), .B1(n13441), .B2(n10918), .ZN(
        n10949) );
  AND2_X2 U7329 ( .A1(n7508), .A2(n7457), .ZN(n7551) );
  NOR2_X2 U7330 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n7508) );
  NAND2_X2 U7331 ( .A1(n9042), .A2(n9041), .ZN(n13806) );
  INV_X1 U7332 ( .A(n9922), .ZN(n12094) );
  AOI22_X2 U7333 ( .A1(n14167), .A2(n14171), .B1(n14147), .B2(n14366), .ZN(
        n14145) );
  OAI22_X2 U7334 ( .A1(n10085), .A2(n10084), .B1(n10083), .B2(n10082), .ZN(
        n10090) );
  NAND2_X2 U7335 ( .A1(n10052), .A2(n10051), .ZN(n10085) );
  CLKBUF_X1 U7336 ( .A(n15098), .Z(n6488) );
  BUF_X4 U7337 ( .A(n15098), .Z(n6489) );
  BUF_X4 U7338 ( .A(n15098), .Z(n6490) );
  NAND2_X2 U7339 ( .A1(n7031), .A2(n9918), .ZN(n15098) );
  XNOR2_X2 U7340 ( .A(n8469), .B(n10549), .ZN(n10436) );
  OAI21_X2 U7341 ( .B1(n9631), .B2(n8678), .A(n6953), .ZN(n6952) );
  BUF_X4 U7342 ( .A(n10288), .Z(n6491) );
  INV_X1 U7343 ( .A(n12290), .ZN(n10288) );
  AOI21_X2 U7344 ( .B1(n7836), .B2(n6861), .A(n6860), .ZN(n7883) );
  AND2_X4 U7345 ( .A1(n9275), .A2(n14326), .ZN(n9278) );
  NOR2_X2 U7347 ( .A1(n15109), .A2(P1_ADDR_REG_0__SCAN_IN), .ZN(n14537) );
  OR2_X4 U7348 ( .A1(n14989), .A2(n9207), .ZN(n12605) );
  XNOR2_X2 U7349 ( .A(n8490), .B(n14623), .ZN(n14626) );
  XNOR2_X1 U7350 ( .A(n14536), .B(n14535), .ZN(n14538) );
  XNOR2_X2 U7351 ( .A(n14488), .B(n14489), .ZN(n14531) );
  AND2_X2 U7352 ( .A1(n7116), .A2(n7115), .ZN(n14488) );
  NAND2_X1 U7353 ( .A1(n13369), .A2(n13368), .ZN(n13367) );
  OAI22_X1 U7354 ( .A1(n12117), .A2(n12115), .B1(n13871), .B2(
        P2_DATAO_REG_29__SCAN_IN), .ZN(n12316) );
  NAND2_X1 U7355 ( .A1(n8192), .A2(n8191), .ZN(n14438) );
  NAND2_X1 U7356 ( .A1(n8088), .A2(n8087), .ZN(n14374) );
  NAND2_X1 U7357 ( .A1(n11952), .A2(n11951), .ZN(n11973) );
  NAND2_X1 U7358 ( .A1(n11700), .A2(n6555), .ZN(n11952) );
  NAND2_X1 U7359 ( .A1(n11332), .A2(n11331), .ZN(n11633) );
  CLKBUF_X2 U7360 ( .A(P2_U3947), .Z(n6492) );
  INV_X1 U7361 ( .A(n10837), .ZN(n14839) );
  INV_X1 U7362 ( .A(n11031), .ZN(n12753) );
  INV_X4 U7363 ( .A(n10086), .ZN(n12610) );
  AND4_X1 U7364 ( .A1(n10934), .A2(n10933), .A3(n10932), .A4(n10931), .ZN(
        n11266) );
  INV_X4 U7365 ( .A(n9035), .ZN(n9172) );
  INV_X2 U7366 ( .A(n10769), .ZN(n6747) );
  CLKBUF_X2 U7367 ( .A(n10369), .Z(n6713) );
  INV_X1 U7368 ( .A(n9926), .ZN(n12119) );
  OR2_X2 U7369 ( .A1(n14988), .A2(n10369), .ZN(n9230) );
  INV_X1 U7370 ( .A(n15026), .ZN(n10987) );
  OAI21_X1 U7371 ( .B1(n8280), .B2(P1_IR_REG_23__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n8281) );
  NAND2_X1 U7372 ( .A1(n7593), .A2(n7594), .ZN(n7597) );
  AND3_X2 U7373 ( .A1(n8782), .A2(n6909), .A3(n6907), .ZN(n7231) );
  AND2_X1 U7374 ( .A1(n8642), .A2(n6908), .ZN(n6906) );
  NAND2_X1 U7375 ( .A1(n12885), .A2(n12497), .ZN(n12834) );
  OAI21_X1 U7376 ( .B1(n12685), .B2(n7206), .A(n7204), .ZN(n7202) );
  AND2_X1 U7377 ( .A1(n7077), .A2(n6863), .ZN(n7075) );
  NAND2_X1 U7378 ( .A1(n13367), .A2(n7241), .ZN(n13417) );
  NAND2_X1 U7379 ( .A1(n13378), .A2(n12596), .ZN(n13369) );
  NAND2_X1 U7380 ( .A1(n12698), .A2(n12697), .ZN(n12696) );
  NAND2_X1 U7381 ( .A1(n9414), .A2(n9413), .ZN(n13952) );
  NAND2_X1 U7382 ( .A1(n13895), .A2(n13896), .ZN(n9414) );
  CLKBUF_X1 U7383 ( .A(n14304), .Z(n6686) );
  INV_X1 U7384 ( .A(n12859), .ZN(n12897) );
  NOR2_X1 U7385 ( .A1(n12082), .A2(n14438), .ZN(n14119) );
  NAND2_X1 U7386 ( .A1(n8175), .A2(n8174), .ZN(n14118) );
  NAND2_X1 U7387 ( .A1(n12986), .A2(n12993), .ZN(n7323) );
  AND2_X1 U7388 ( .A1(n7278), .A2(n7277), .ZN(n12577) );
  NAND2_X1 U7389 ( .A1(n13981), .A2(n13982), .ZN(n7108) );
  NAND2_X1 U7390 ( .A1(n13542), .A2(n13541), .ZN(n13698) );
  NAND2_X1 U7391 ( .A1(n7160), .A2(n12089), .ZN(n12281) );
  NAND2_X1 U7392 ( .A1(n6797), .A2(n6796), .ZN(n13981) );
  OAI211_X1 U7393 ( .C1(n8149), .C2(n13878), .A(n6846), .B(n6845), .ZN(n14135)
         );
  NAND2_X1 U7394 ( .A1(n8149), .A2(n8148), .ZN(n14138) );
  NOR2_X1 U7395 ( .A1(n13419), .A2(n12599), .ZN(n7241) );
  CLKBUF_X1 U7396 ( .A(n11861), .Z(n6711) );
  NAND2_X2 U7397 ( .A1(n8043), .A2(n8042), .ZN(n14385) );
  NAND2_X1 U7398 ( .A1(n8106), .A2(n8105), .ZN(n14366) );
  NAND2_X1 U7399 ( .A1(n9096), .A2(n9095), .ZN(n13635) );
  NAND2_X1 U7400 ( .A1(n9077), .A2(n9076), .ZN(n13791) );
  AND2_X1 U7401 ( .A1(n7269), .A2(n11666), .ZN(n11669) );
  NAND2_X1 U7402 ( .A1(n11693), .A2(n12425), .ZN(n11694) );
  NAND2_X1 U7403 ( .A1(n7956), .A2(n7955), .ZN(n14409) );
  AND2_X1 U7404 ( .A1(n11588), .A2(n11587), .ZN(n11591) );
  OAI21_X1 U7405 ( .B1(n14626), .B2(n7052), .A(n7051), .ZN(n14652) );
  NAND2_X1 U7406 ( .A1(n8760), .A2(n8759), .ZN(n8777) );
  NAND2_X1 U7407 ( .A1(n12023), .A2(n12022), .ZN(n12021) );
  NAND2_X1 U7408 ( .A1(n11370), .A2(n11369), .ZN(n11496) );
  NOR2_X1 U7409 ( .A1(n11508), .A2(n6723), .ZN(n8541) );
  NAND2_X1 U7410 ( .A1(n11895), .A2(n9343), .ZN(n12023) );
  NAND2_X1 U7411 ( .A1(n8950), .A2(n8949), .ZN(n13745) );
  NAND2_X1 U7412 ( .A1(n7939), .A2(n7938), .ZN(n14414) );
  NAND2_X1 U7413 ( .A1(n11227), .A2(n6768), .ZN(n11739) );
  NAND2_X1 U7414 ( .A1(n7987), .A2(n7986), .ZN(n14404) );
  NAND2_X1 U7415 ( .A1(n8985), .A2(n8984), .ZN(n13822) );
  NOR2_X1 U7416 ( .A1(n11426), .A2(n11427), .ZN(n11425) );
  OAI21_X1 U7417 ( .B1(n10853), .B2(n8440), .A(n8439), .ZN(n11455) );
  NOR2_X1 U7418 ( .A1(n8488), .A2(n12765), .ZN(n12777) );
  NAND2_X1 U7419 ( .A1(n8928), .A2(n8927), .ZN(n13569) );
  NOR2_X1 U7420 ( .A1(n12766), .A2(n14673), .ZN(n12765) );
  OAI21_X2 U7421 ( .B1(n11147), .B2(n9514), .A(n9513), .ZN(n11238) );
  XNOR2_X1 U7422 ( .A(n8487), .B(n8540), .ZN(n12766) );
  NAND2_X1 U7423 ( .A1(n7891), .A2(n7890), .ZN(n14425) );
  NAND2_X1 U7424 ( .A1(n7842), .A2(n7841), .ZN(n13892) );
  NAND2_X1 U7425 ( .A1(n8915), .A2(n8914), .ZN(n11964) );
  OAI21_X1 U7426 ( .B1(n15152), .B2(n8422), .A(n8421), .ZN(n10856) );
  NAND2_X1 U7427 ( .A1(n8861), .A2(n8860), .ZN(n11638) );
  OR2_X1 U7428 ( .A1(n11448), .A2(n11447), .ZN(n11445) );
  NAND2_X1 U7429 ( .A1(n7826), .A2(n7825), .ZN(n11736) );
  NOR2_X1 U7430 ( .A1(n11434), .A2(n14684), .ZN(n11433) );
  NAND2_X1 U7431 ( .A1(n8836), .A2(n8835), .ZN(n14716) );
  AND2_X1 U7432 ( .A1(n11441), .A2(n8483), .ZN(n8484) );
  INV_X2 U7433 ( .A(n15002), .ZN(n15005) );
  NAND2_X1 U7434 ( .A1(n6880), .A2(n6879), .ZN(n11441) );
  AND2_X2 U7435 ( .A1(n10382), .A2(n10381), .ZN(n15066) );
  CLKBUF_X1 U7436 ( .A(n7816), .Z(n7794) );
  AND2_X1 U7437 ( .A1(n11008), .A2(n11007), .ZN(n11027) );
  NAND2_X1 U7438 ( .A1(n8764), .A2(n8763), .ZN(n15068) );
  NAND3_X1 U7439 ( .A1(n7746), .A2(SI_10_), .A3(n7767), .ZN(n7768) );
  AND3_X1 U7440 ( .A1(n6882), .A2(n8476), .A3(P3_REG1_REG_7__SCAN_IN), .ZN(
        n15160) );
  OR2_X1 U7441 ( .A1(n7745), .A2(n7744), .ZN(n7746) );
  NAND2_X1 U7442 ( .A1(n7745), .A2(n7744), .ZN(n7767) );
  AOI22_X1 U7443 ( .A1(n10143), .A2(n10144), .B1(n9281), .B2(n9280), .ZN(
        n10138) );
  NAND2_X1 U7444 ( .A1(n7678), .A2(n7677), .ZN(n11200) );
  XNOR2_X1 U7445 ( .A(n14551), .B(n7123), .ZN(n14597) );
  AND3_X1 U7446 ( .A1(n11086), .A2(n11085), .A3(n11084), .ZN(n11210) );
  INV_X1 U7447 ( .A(n11266), .ZN(n12751) );
  OR2_X1 U7448 ( .A1(n10400), .A2(n8475), .ZN(n8477) );
  NAND2_X2 U7449 ( .A1(n12553), .A2(n14307), .ZN(n14313) );
  AND2_X1 U7450 ( .A1(n6864), .A2(n6598), .ZN(n14551) );
  OR2_X1 U7451 ( .A1(n15126), .A2(n6985), .ZN(n6983) );
  NAND2_X1 U7452 ( .A1(n9773), .A2(n9772), .ZN(n9874) );
  NAND2_X1 U7453 ( .A1(n10346), .A2(n9991), .ZN(n10389) );
  AND3_X1 U7454 ( .A1(n10453), .A2(n10452), .A3(n10451), .ZN(n10992) );
  NAND2_X1 U7455 ( .A1(n6721), .A2(n7511), .ZN(n10623) );
  AND3_X1 U7456 ( .A1(n10800), .A2(n10799), .A3(n10798), .ZN(n11021) );
  AND3_X1 U7457 ( .A1(n10552), .A2(n10551), .A3(n10550), .ZN(n15223) );
  INV_X1 U7458 ( .A(n14041), .ZN(n10900) );
  NAND4_X2 U7459 ( .A1(n7575), .A2(n7574), .A3(n7573), .A4(n7572), .ZN(n14041)
         );
  NAND2_X2 U7460 ( .A1(n12094), .A2(n12119), .ZN(n10791) );
  CLKBUF_X1 U7461 ( .A(n10200), .Z(n10203) );
  XNOR2_X1 U7462 ( .A(n8590), .B(P2_IR_REG_22__SCAN_IN), .ZN(n10369) );
  AND2_X1 U7464 ( .A1(n11516), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n6723) );
  NAND2_X1 U7465 ( .A1(n13322), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9919) );
  INV_X1 U7466 ( .A(n7032), .ZN(n7031) );
  INV_X2 U7467 ( .A(n9669), .ZN(n8964) );
  XOR2_X1 U7468 ( .A(n9606), .B(n8522), .Z(n10434) );
  NAND2_X1 U7469 ( .A1(n7554), .A2(n7553), .ZN(n7558) );
  NAND2_X2 U7470 ( .A1(n9915), .A2(n9270), .ZN(n14326) );
  INV_X1 U7471 ( .A(n14476), .ZN(n7480) );
  NAND2_X1 U7472 ( .A1(n8179), .A2(n11493), .ZN(n9499) );
  AND2_X1 U7473 ( .A1(n6979), .A2(n6976), .ZN(n8522) );
  NAND2_X1 U7475 ( .A1(n7495), .A2(n7494), .ZN(n14059) );
  NAND2_X2 U7476 ( .A1(n7532), .A2(n8280), .ZN(n9915) );
  XNOR2_X1 U7477 ( .A(n8318), .B(n8317), .ZN(n11748) );
  OAI21_X1 U7478 ( .B1(n8322), .B2(P3_IR_REG_24__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8318) );
  XNOR2_X1 U7479 ( .A(n8460), .B(n8459), .ZN(n12345) );
  NAND2_X1 U7480 ( .A1(n8322), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7171) );
  CLKBUF_X1 U7481 ( .A(n8610), .Z(n11523) );
  NAND2_X1 U7482 ( .A1(n7493), .A2(n7492), .ZN(n7495) );
  NAND2_X1 U7483 ( .A1(n7541), .A2(n6519), .ZN(n11493) );
  XNOR2_X1 U7484 ( .A(n8281), .B(P1_IR_REG_24__SCAN_IN), .ZN(n9447) );
  NAND2_X1 U7485 ( .A1(n7538), .A2(n7209), .ZN(n11614) );
  NAND2_X1 U7486 ( .A1(n8288), .A2(n8287), .ZN(n11882) );
  NAND2_X1 U7487 ( .A1(n8285), .A2(n8284), .ZN(n12009) );
  XNOR2_X1 U7488 ( .A(n8508), .B(n8507), .ZN(n12367) );
  NAND2_X1 U7489 ( .A1(n7501), .A2(n7503), .ZN(n6838) );
  OR2_X1 U7490 ( .A1(n7500), .A2(SI_1_), .ZN(n7501) );
  NAND2_X2 U7491 ( .A1(n8621), .A2(P2_U3088), .ZN(n13870) );
  AOI21_X1 U7492 ( .B1(n6835), .B2(n7672), .A(n6635), .ZN(n6833) );
  NAND2_X1 U7493 ( .A1(n7060), .A2(n6763), .ZN(n7494) );
  NOR2_X1 U7494 ( .A1(n8311), .A2(P3_IR_REG_20__SCAN_IN), .ZN(n8505) );
  NOR2_X1 U7495 ( .A1(n7340), .A2(P3_IR_REG_26__SCAN_IN), .ZN(n7339) );
  NOR2_X1 U7496 ( .A1(n7149), .A2(n6641), .ZN(n7147) );
  NAND2_X1 U7497 ( .A1(n8346), .A2(n7078), .ZN(n6958) );
  AND2_X2 U7498 ( .A1(n8642), .A2(n7372), .ZN(n8782) );
  AND2_X1 U7499 ( .A1(n7551), .A2(n7460), .ZN(n7670) );
  INV_X1 U7500 ( .A(n8924), .ZN(n6907) );
  AND2_X1 U7501 ( .A1(n8302), .A2(n8306), .ZN(n7187) );
  AND3_X1 U7502 ( .A1(n8407), .A2(n8295), .A3(n8406), .ZN(n8298) );
  AND4_X1 U7503 ( .A1(n7887), .A2(n7468), .A3(n7467), .A4(n7466), .ZN(n6499)
         );
  AND2_X2 U7504 ( .A1(n8617), .A2(n7373), .ZN(n8642) );
  AND3_X1 U7505 ( .A1(n8301), .A2(n8300), .A3(n8299), .ZN(n8305) );
  AND4_X1 U7506 ( .A1(n7464), .A2(n7463), .A3(n7462), .A4(n7461), .ZN(n7465)
         );
  NAND2_X1 U7507 ( .A1(P1_DATAO_REG_12__SCAN_IN), .A2(n10169), .ZN(n9772) );
  XNOR2_X1 U7508 ( .A(P3_ADDR_REG_1__SCAN_IN), .B(P1_ADDR_REG_1__SCAN_IN), 
        .ZN(n6878) );
  NOR2_X1 U7509 ( .A1(P3_IR_REG_2__SCAN_IN), .A2(P3_IR_REG_3__SCAN_IN), .ZN(
        n8296) );
  INV_X4 U7510 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  INV_X1 U7511 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n7373) );
  INV_X1 U7512 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n8307) );
  INV_X1 U7513 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n13121) );
  NOR2_X1 U7514 ( .A1(P3_IR_REG_17__SCAN_IN), .A2(P3_IR_REG_15__SCAN_IN), .ZN(
        n8304) );
  NOR2_X1 U7515 ( .A1(P3_IR_REG_16__SCAN_IN), .A2(P3_IR_REG_12__SCAN_IN), .ZN(
        n8303) );
  INV_X1 U7516 ( .A(P3_IR_REG_25__SCAN_IN), .ZN(n8317) );
  NOR2_X1 U7518 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_9__SCAN_IN), .ZN(
        n8575) );
  XNOR2_X1 U7519 ( .A(n6868), .B(P3_ADDR_REG_4__SCAN_IN), .ZN(n14529) );
  INV_X1 U7520 ( .A(n6868), .ZN(n14490) );
  NAND2_X1 U7522 ( .A1(n9471), .A2(n9289), .ZN(n9506) );
  NAND2_X2 U7523 ( .A1(n7231), .A2(n7230), .ZN(n8567) );
  XNOR2_X1 U7524 ( .A(n14558), .B(n7121), .ZN(n15287) );
  INV_X1 U7525 ( .A(n7527), .ZN(n7954) );
  AND2_X1 U7526 ( .A1(n8569), .A2(n8568), .ZN(n6494) );
  OR2_X2 U7527 ( .A1(n6932), .A2(n6749), .ZN(n8573) );
  AOI21_X2 U7528 ( .B1(P3_REG1_REG_14__SCAN_IN), .B2(n12783), .A(n8489), .ZN(
        n8490) );
  NOR2_X2 U7529 ( .A1(n10720), .A2(n15068), .ZN(n6948) );
  INV_X1 U7530 ( .A(n10375), .ZN(n15042) );
  NAND2_X2 U7531 ( .A1(n8662), .A2(n8661), .ZN(n10375) );
  NAND2_X1 U7532 ( .A1(n14191), .A2(n6566), .ZN(n14167) );
  AND2_X4 U7533 ( .A1(n9922), .A2(n9926), .ZN(n10235) );
  OAI21_X2 U7534 ( .B1(n13038), .B2(n12841), .A(n12842), .ZN(n13027) );
  INV_X1 U7535 ( .A(n12290), .ZN(n6495) );
  XNOR2_X1 U7536 ( .A(n8355), .B(n8354), .ZN(n8357) );
  XNOR2_X2 U7537 ( .A(n6935), .B(n15026), .ZN(n10349) );
  AND2_X1 U7538 ( .A1(n6499), .A2(n7491), .ZN(n7367) );
  AND2_X1 U7539 ( .A1(n8282), .A2(n6539), .ZN(n7473) );
  INV_X1 U7540 ( .A(SI_15_), .ZN(n7879) );
  NAND2_X1 U7541 ( .A1(n13032), .A2(n13031), .ZN(n7030) );
  NAND2_X1 U7542 ( .A1(n6816), .A2(n6518), .ZN(n6815) );
  INV_X1 U7543 ( .A(n13993), .ZN(n6816) );
  INV_X1 U7544 ( .A(n8137), .ZN(n8036) );
  INV_X1 U7545 ( .A(n8185), .ZN(n8033) );
  BUF_X1 U7546 ( .A(n7623), .Z(n8119) );
  INV_X1 U7547 ( .A(n7608), .ZN(n7623) );
  AND2_X1 U7548 ( .A1(n11614), .A2(n11493), .ZN(n9270) );
  AOI22_X1 U7549 ( .A1(n13448), .A2(n9087), .B1(n10769), .B2(n9035), .ZN(n8654) );
  INV_X1 U7550 ( .A(n8066), .ZN(n6718) );
  INV_X1 U7551 ( .A(n8067), .ZN(n6719) );
  OAI21_X1 U7552 ( .B1(n7793), .B2(n7792), .A(n7791), .ZN(n7816) );
  AND2_X1 U7553 ( .A1(n7459), .A2(n7458), .ZN(n7460) );
  INV_X1 U7554 ( .A(n10235), .ZN(n10788) );
  OR2_X1 U7555 ( .A1(n12872), .A2(n12881), .ZN(n12508) );
  NAND2_X1 U7556 ( .A1(n12860), .A2(n7328), .ZN(n7327) );
  NAND2_X1 U7557 ( .A1(n12857), .A2(n7329), .ZN(n7328) );
  INV_X1 U7558 ( .A(n12856), .ZN(n7329) );
  OR2_X1 U7559 ( .A1(n13066), .A2(n12923), .ZN(n12349) );
  NAND2_X1 U7560 ( .A1(n11127), .A2(n12396), .ZN(n11090) );
  INV_X1 U7561 ( .A(n8372), .ZN(n8297) );
  AND2_X1 U7562 ( .A1(n6498), .A2(n6532), .ZN(n7127) );
  NAND2_X1 U7563 ( .A1(n11669), .A2(n11668), .ZN(n11861) );
  INV_X1 U7564 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n8557) );
  NAND2_X1 U7565 ( .A1(n13588), .A2(n6533), .ZN(n7303) );
  INV_X1 U7566 ( .A(n11247), .ZN(n6916) );
  AND2_X1 U7567 ( .A1(n14716), .A2(n11252), .ZN(n11248) );
  INV_X1 U7569 ( .A(n11656), .ZN(n6832) );
  INV_X1 U7570 ( .A(n14233), .ZN(n9493) );
  NOR2_X1 U7571 ( .A1(n6548), .A2(n6782), .ZN(n6781) );
  INV_X1 U7572 ( .A(n9484), .ZN(n6782) );
  NOR2_X1 U7573 ( .A1(n11767), .A2(n11663), .ZN(n6893) );
  AND2_X1 U7574 ( .A1(n9436), .A2(n9657), .ZN(n10594) );
  NAND2_X1 U7575 ( .A1(n7670), .A2(n7465), .ZN(n7852) );
  OAI21_X1 U7576 ( .B1(n8160), .B2(n8159), .A(n8163), .ZN(n8211) );
  INV_X1 U7577 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n8283) );
  AND3_X1 U7578 ( .A1(n7471), .A2(n7470), .A3(n7469), .ZN(n8282) );
  INV_X1 U7579 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n7468) );
  INV_X1 U7580 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n7467) );
  NAND2_X1 U7581 ( .A1(n7849), .A2(SI_14_), .ZN(n6861) );
  AND2_X1 U7582 ( .A1(n7850), .A2(n9877), .ZN(n6860) );
  NAND2_X1 U7583 ( .A1(n7768), .A2(n7767), .ZN(n7793) );
  NAND2_X1 U7584 ( .A1(n7558), .A2(n7557), .ZN(n7598) );
  NOR2_X1 U7585 ( .A1(n14502), .A2(n6671), .ZN(n14564) );
  AND2_X1 U7586 ( .A1(n14503), .A2(P1_ADDR_REG_8__SCAN_IN), .ZN(n6671) );
  XNOR2_X1 U7587 ( .A(n8524), .B(n15138), .ZN(n15126) );
  NAND2_X1 U7588 ( .A1(n6883), .A2(n15154), .ZN(n6882) );
  INV_X1 U7589 ( .A(n11443), .ZN(n6879) );
  AND2_X1 U7590 ( .A1(n6974), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n6971) );
  NAND2_X1 U7591 ( .A1(n12892), .A2(n12493), .ZN(n12886) );
  OR2_X1 U7592 ( .A1(n13090), .A2(n12658), .ZN(n12354) );
  AOI21_X1 U7593 ( .B1(n11989), .B2(n7001), .A(n6999), .ZN(n6998) );
  NAND2_X1 U7594 ( .A1(n7000), .A2(n13043), .ZN(n6999) );
  AOI21_X1 U7595 ( .B1(n12526), .B2(n7015), .A(n7014), .ZN(n7013) );
  INV_X1 U7596 ( .A(n12428), .ZN(n7015) );
  INV_X1 U7597 ( .A(n11392), .ZN(n12162) );
  INV_X2 U7598 ( .A(n12165), .ZN(n12311) );
  NAND2_X1 U7599 ( .A1(P1_DATAO_REG_22__SCAN_IN), .A2(n11064), .ZN(n6768) );
  NAND2_X1 U7600 ( .A1(n7140), .A2(n7138), .ZN(n11062) );
  NAND2_X1 U7601 ( .A1(P2_DATAO_REG_20__SCAN_IN), .A2(n7139), .ZN(n7138) );
  NAND2_X1 U7602 ( .A1(n10961), .A2(n10962), .ZN(n7140) );
  NAND2_X1 U7603 ( .A1(n9641), .A2(n9640), .ZN(n9643) );
  CLKBUF_X1 U7604 ( .A(n8329), .Z(n8424) );
  NAND2_X1 U7605 ( .A1(n9584), .A2(n9583), .ZN(n9586) );
  AND2_X1 U7606 ( .A1(n8395), .A2(n8403), .ZN(n8528) );
  AOI21_X1 U7607 ( .B1(n7248), .B2(n7247), .A(n6585), .ZN(n7246) );
  NOR2_X1 U7608 ( .A1(n9981), .A2(n15013), .ZN(n9989) );
  INV_X1 U7609 ( .A(n7308), .ZN(n7307) );
  AOI21_X1 U7610 ( .B1(n7306), .B2(n7308), .A(n7305), .ZN(n7304) );
  AOI21_X1 U7611 ( .B1(n7379), .B2(n7381), .A(n6569), .ZN(n7377) );
  NAND2_X1 U7612 ( .A1(n6703), .A2(n13575), .ZN(n6706) );
  NAND2_X1 U7613 ( .A1(n13734), .A2(n6709), .ZN(n6708) );
  AND2_X1 U7614 ( .A1(n13569), .A2(n13567), .ZN(n13535) );
  NAND2_X1 U7615 ( .A1(n6658), .A2(n6657), .ZN(n14704) );
  OR2_X1 U7616 ( .A1(n11638), .A2(n13437), .ZN(n6657) );
  NAND2_X1 U7617 ( .A1(n11547), .A2(n6556), .ZN(n6658) );
  INV_X2 U7618 ( .A(n8657), .ZN(n8965) );
  XNOR2_X1 U7619 ( .A(n11059), .B(n13440), .ZN(n10953) );
  OR2_X1 U7620 ( .A1(n6713), .A2(n11616), .ZN(n14989) );
  OR2_X1 U7621 ( .A1(n14989), .A2(n9986), .ZN(n15077) );
  NOR2_X1 U7622 ( .A1(P2_IR_REG_27__SCAN_IN), .A2(P2_IR_REG_26__SCAN_IN), .ZN(
        n8597) );
  NAND2_X1 U7623 ( .A1(n6813), .A2(n6809), .ZN(n6805) );
  NAND2_X1 U7624 ( .A1(n7082), .A2(n7083), .ZN(n13971) );
  AND2_X1 U7625 ( .A1(n13973), .A2(n7084), .ZN(n7083) );
  NAND2_X1 U7626 ( .A1(n13914), .A2(n9399), .ZN(n7084) );
  NOR2_X1 U7627 ( .A1(n14135), .A2(n7362), .ZN(n7361) );
  INV_X1 U7628 ( .A(n9497), .ZN(n7362) );
  NAND2_X1 U7629 ( .A1(n14300), .A2(n7354), .ZN(n7353) );
  NOR2_X1 U7630 ( .A1(n14280), .A2(n7355), .ZN(n7354) );
  INV_X1 U7631 ( .A(n9489), .ZN(n7355) );
  OAI21_X2 U7632 ( .B1(n11772), .B2(n11771), .A(n9483), .ZN(n11839) );
  AOI21_X1 U7633 ( .B1(n6774), .B2(n6776), .A(n6574), .ZN(n6773) );
  NAND2_X1 U7634 ( .A1(n14427), .A2(n9502), .ZN(n9553) );
  AND2_X1 U7635 ( .A1(n9666), .A2(n8291), .ZN(n14321) );
  NAND2_X1 U7636 ( .A1(n9667), .A2(n10187), .ZN(n7823) );
  MUX2_X1 U7637 ( .A(P1_IR_REG_31__SCAN_IN), .B(n7531), .S(
        P1_IR_REG_22__SCAN_IN), .Z(n7532) );
  OR2_X1 U7638 ( .A1(n15284), .A2(P2_ADDR_REG_5__SCAN_IN), .ZN(n6864) );
  NAND2_X1 U7639 ( .A1(n10155), .A2(n15103), .ZN(n10423) );
  XNOR2_X1 U7640 ( .A(n8498), .B(n6888), .ZN(n6887) );
  OR2_X1 U7641 ( .A1(n11815), .A2(n9249), .ZN(n9983) );
  NAND2_X1 U7642 ( .A1(n9154), .A2(n9153), .ZN(n13585) );
  OAI21_X1 U7643 ( .B1(n14239), .B2(n8119), .A(n8038), .ZN(n14249) );
  INV_X1 U7644 ( .A(n8654), .ZN(n6757) );
  INV_X1 U7645 ( .A(n7755), .ZN(n7226) );
  NOR2_X1 U7646 ( .A1(n8777), .A2(n8776), .ZN(n6735) );
  INV_X1 U7647 ( .A(n8799), .ZN(n7434) );
  NAND2_X1 U7648 ( .A1(n8873), .A2(n8872), .ZN(n7431) );
  NAND2_X1 U7649 ( .A1(n7427), .A2(n7426), .ZN(n7425) );
  INV_X1 U7650 ( .A(n8831), .ZN(n7427) );
  INV_X1 U7651 ( .A(n8962), .ZN(n7420) );
  INV_X1 U7652 ( .A(n6551), .ZN(n7421) );
  NAND2_X1 U7653 ( .A1(n8962), .A2(n6551), .ZN(n7418) );
  INV_X1 U7654 ( .A(n8026), .ZN(n6761) );
  INV_X1 U7655 ( .A(n8027), .ZN(n6762) );
  INV_X1 U7656 ( .A(n9036), .ZN(n6695) );
  NAND2_X1 U7657 ( .A1(n8089), .A2(n8091), .ZN(n7216) );
  AND4_X1 U7658 ( .A1(n14303), .A2(n8247), .A3(n14332), .A4(n11832), .ZN(n8248) );
  NAND2_X1 U7659 ( .A1(n10184), .A2(n9913), .ZN(n8238) );
  OAI21_X1 U7660 ( .B1(n7320), .B2(n6854), .A(n6852), .ZN(n8002) );
  INV_X1 U7661 ( .A(n6855), .ZN(n6854) );
  AND2_X1 U7662 ( .A1(n6853), .A2(n7982), .ZN(n6852) );
  NOR2_X1 U7663 ( .A1(n7721), .A2(n7694), .ZN(n7314) );
  INV_X1 U7664 ( .A(n7718), .ZN(n7317) );
  NAND2_X1 U7665 ( .A1(n6527), .A2(n7185), .ZN(n7184) );
  INV_X1 U7666 ( .A(n15111), .ZN(n6992) );
  INV_X1 U7667 ( .A(n11511), .ZN(n7064) );
  OR2_X1 U7668 ( .A1(n8485), .A2(n6633), .ZN(n6884) );
  NOR2_X1 U7669 ( .A1(n11941), .A2(n6728), .ZN(n6727) );
  INV_X1 U7670 ( .A(n8445), .ZN(n6728) );
  NOR2_X1 U7671 ( .A1(n14652), .A2(n6881), .ZN(n8493) );
  NOR2_X1 U7672 ( .A1(n14646), .A2(n8492), .ZN(n6881) );
  INV_X1 U7673 ( .A(n12354), .ZN(n7026) );
  OR2_X1 U7674 ( .A1(n13082), .A2(n12636), .ZN(n12465) );
  AND2_X1 U7675 ( .A1(n7332), .A2(n11214), .ZN(n7331) );
  OR2_X1 U7676 ( .A1(n12513), .A2(n7336), .ZN(n7332) );
  INV_X1 U7677 ( .A(n11069), .ZN(n7336) );
  NOR2_X1 U7678 ( .A1(n13769), .A2(n13635), .ZN(n6943) );
  NOR2_X1 U7679 ( .A1(n7380), .A2(n6557), .ZN(n7379) );
  NOR2_X1 U7680 ( .A1(n13549), .A2(n7381), .ZN(n7380) );
  INV_X1 U7681 ( .A(n7386), .ZN(n7385) );
  OAI21_X1 U7682 ( .B1(n13742), .B2(n7387), .A(n13538), .ZN(n7386) );
  INV_X1 U7683 ( .A(n13537), .ZN(n7387) );
  OR2_X1 U7684 ( .A1(n13734), .A2(n13575), .ZN(n13539) );
  INV_X1 U7685 ( .A(n10367), .ZN(n6922) );
  INV_X1 U7686 ( .A(n10569), .ZN(n6919) );
  AND2_X1 U7687 ( .A1(n10709), .A2(n13443), .ZN(n7374) );
  XNOR2_X1 U7688 ( .A(n15049), .B(n13446), .ZN(n14971) );
  NAND2_X1 U7689 ( .A1(n7093), .A2(n6575), .ZN(n7092) );
  OR2_X1 U7690 ( .A1(n7095), .A2(n7094), .ZN(n7093) );
  AOI21_X1 U7691 ( .B1(n7040), .B2(n7042), .A(n6577), .ZN(n7039) );
  INV_X1 U7692 ( .A(n9499), .ZN(n9264) );
  NAND2_X1 U7693 ( .A1(n8239), .A2(n8238), .ZN(n10171) );
  NAND2_X1 U7694 ( .A1(n10171), .A2(n10170), .ZN(n10172) );
  INV_X1 U7695 ( .A(n14171), .ZN(n7071) );
  NOR2_X1 U7696 ( .A1(n14192), .A2(n7073), .ZN(n7072) );
  INV_X1 U7697 ( .A(n9540), .ZN(n7073) );
  NAND2_X1 U7698 ( .A1(n7049), .A2(n9532), .ZN(n14284) );
  NOR2_X1 U7699 ( .A1(n14283), .A2(n7048), .ZN(n7047) );
  INV_X1 U7700 ( .A(n9532), .ZN(n7048) );
  NAND2_X1 U7701 ( .A1(n7050), .A2(n14303), .ZN(n7049) );
  INV_X1 U7702 ( .A(n6686), .ZN(n7050) );
  CLKBUF_X1 U7703 ( .A(n9277), .Z(n10177) );
  OAI21_X1 U7704 ( .B1(n8125), .B2(n11877), .A(n8124), .ZN(n8127) );
  OAI21_X1 U7705 ( .B1(n8103), .B2(n8102), .A(n8101), .ZN(n8125) );
  INV_X1 U7706 ( .A(n6850), .ZN(n6849) );
  OAI21_X1 U7707 ( .B1(n8021), .B2(n6851), .A(n8061), .ZN(n6850) );
  INV_X1 U7708 ( .A(n8054), .ZN(n6851) );
  NAND2_X1 U7709 ( .A1(n7111), .A2(n7109), .ZN(n8280) );
  AND2_X1 U7710 ( .A1(n7112), .A2(n7110), .ZN(n7109) );
  INV_X1 U7711 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n7110) );
  INV_X1 U7712 ( .A(n7533), .ZN(n7111) );
  NOR2_X1 U7713 ( .A1(n7113), .A2(P1_IR_REG_21__SCAN_IN), .ZN(n7112) );
  NAND2_X1 U7714 ( .A1(n7899), .A2(n7898), .ZN(n7320) );
  AOI21_X1 U7715 ( .B1(n7286), .B2(n7288), .A(n6590), .ZN(n7283) );
  NAND2_X1 U7716 ( .A1(n7504), .A2(SI_2_), .ZN(n7553) );
  OAI22_X1 U7717 ( .A1(n14554), .A2(n14497), .B1(P1_ADDR_REG_6__SCAN_IN), .B2(
        n14496), .ZN(n14498) );
  INV_X1 U7718 ( .A(P3_ADDR_REG_6__SCAN_IN), .ZN(n14496) );
  OAI22_X1 U7719 ( .A1(n14511), .A2(n14573), .B1(P1_ADDR_REG_13__SCAN_IN), 
        .B2(n14571), .ZN(n14518) );
  OR2_X1 U7720 ( .A1(n12012), .A2(n12017), .ZN(n7185) );
  NAND2_X1 U7721 ( .A1(n12374), .A2(n6486), .ZN(n10298) );
  NAND2_X1 U7722 ( .A1(n11591), .A2(n11590), .ZN(n11784) );
  AND2_X1 U7723 ( .A1(n11783), .A2(n11785), .ZN(n7178) );
  NOR2_X1 U7724 ( .A1(n11316), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n11399) );
  AOI21_X1 U7725 ( .B1(n12663), .B2(n7205), .A(n6593), .ZN(n7204) );
  INV_X1 U7726 ( .A(n12236), .ZN(n7205) );
  NAND2_X1 U7727 ( .A1(n12663), .A2(n7207), .ZN(n7206) );
  INV_X1 U7728 ( .A(n12237), .ZN(n7207) );
  INV_X1 U7729 ( .A(n12218), .ZN(n7196) );
  NAND2_X1 U7730 ( .A1(n15105), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n8518) );
  NOR2_X1 U7731 ( .A1(n10158), .A2(n8344), .ZN(n10157) );
  INV_X1 U7732 ( .A(n10418), .ZN(n6980) );
  NAND2_X1 U7733 ( .A1(n8523), .A2(n6992), .ZN(n6990) );
  OR2_X1 U7734 ( .A1(n10434), .A2(n6991), .ZN(n6989) );
  NAND2_X1 U7735 ( .A1(n6992), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n6991) );
  XNOR2_X1 U7736 ( .A(n8472), .B(n10923), .ZN(n15135) );
  OR2_X1 U7737 ( .A1(n15135), .A2(n8381), .ZN(n7068) );
  OR2_X1 U7738 ( .A1(n15160), .A2(n8478), .ZN(n7057) );
  OR2_X1 U7739 ( .A1(n8434), .A2(P3_IR_REG_11__SCAN_IN), .ZN(n8339) );
  AOI21_X1 U7740 ( .B1(n8443), .B2(n11516), .A(n11512), .ZN(n12761) );
  NAND2_X1 U7741 ( .A1(n12761), .A2(n12760), .ZN(n12759) );
  AOI21_X1 U7742 ( .B1(n8452), .B2(n10327), .A(n12797), .ZN(n8456) );
  NAND2_X1 U7743 ( .A1(n12861), .A2(n12857), .ZN(n7325) );
  NAND2_X1 U7744 ( .A1(n7327), .A2(n12861), .ZN(n7324) );
  INV_X1 U7745 ( .A(n7022), .ZN(n12893) );
  AOI21_X1 U7746 ( .B1(n7019), .B2(n7018), .A(n7017), .ZN(n7016) );
  INV_X1 U7747 ( .A(n12349), .ZN(n7017) );
  NAND2_X1 U7748 ( .A1(n12893), .A2(n12897), .ZN(n12892) );
  OR2_X1 U7749 ( .A1(n12266), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n12285) );
  AND2_X1 U7750 ( .A1(n12350), .A2(n12349), .ZN(n12913) );
  NAND2_X1 U7751 ( .A1(n12222), .A2(n12221), .ZN(n12241) );
  AND2_X1 U7752 ( .A1(n12207), .A2(n12637), .ZN(n12222) );
  NAND2_X1 U7753 ( .A1(n13003), .A2(n6500), .ZN(n12990) );
  AND2_X1 U7754 ( .A1(n12168), .A2(n12167), .ZN(n12179) );
  NOR2_X1 U7755 ( .A1(n13018), .A2(n7029), .ZN(n7028) );
  INV_X1 U7756 ( .A(n13010), .ZN(n13018) );
  AND2_X1 U7757 ( .A1(n13002), .A2(n12451), .ZN(n13010) );
  AND2_X1 U7758 ( .A1(n12355), .A2(n12358), .ZN(n13031) );
  AND2_X1 U7759 ( .A1(n12429), .A2(n12428), .ZN(n12525) );
  NAND2_X1 U7760 ( .A1(n11694), .A2(n12525), .ZN(n11714) );
  AOI21_X1 U7761 ( .B1(n6497), .B2(n12520), .A(n6586), .ZN(n7343) );
  AND4_X1 U7762 ( .A1(n11539), .A2(n11538), .A3(n11537), .A4(n11536), .ZN(
        n11926) );
  OR2_X1 U7763 ( .A1(n6481), .A2(n12520), .ZN(n7344) );
  AND2_X1 U7764 ( .A1(n7344), .A2(n6521), .ZN(n11398) );
  AOI21_X1 U7765 ( .B1(n7007), .B2(n7009), .A(n7006), .ZN(n7005) );
  INV_X1 U7766 ( .A(n12407), .ZN(n7006) );
  AND2_X1 U7767 ( .A1(n12396), .A2(n12398), .ZN(n12513) );
  NAND2_X1 U7768 ( .A1(n15171), .A2(n15177), .ZN(n15170) );
  NAND2_X1 U7769 ( .A1(n10482), .A2(n12347), .ZN(n15200) );
  INV_X1 U7770 ( .A(n15197), .ZN(n13040) );
  NAND2_X1 U7771 ( .A1(n10498), .A2(n10479), .ZN(n10485) );
  NAND2_X1 U7772 ( .A1(n12872), .A2(n15224), .ZN(n7023) );
  NAND2_X1 U7773 ( .A1(n12177), .A2(n12176), .ZN(n13090) );
  NAND2_X1 U7774 ( .A1(n12132), .A2(n12131), .ZN(n13106) );
  OAI22_X1 U7775 ( .A1(n12281), .A2(n12090), .B1(P1_DATAO_REG_28__SCAN_IN), 
        .B2(n12277), .ZN(n12117) );
  NAND2_X1 U7776 ( .A1(n11874), .A2(n6677), .ZN(n12085) );
  NAND2_X1 U7777 ( .A1(P1_DATAO_REG_25__SCAN_IN), .A2(n6678), .ZN(n6677) );
  XNOR2_X1 U7778 ( .A(n11742), .B(P2_DATAO_REG_24__SCAN_IN), .ZN(n12219) );
  AOI21_X1 U7779 ( .B1(n11062), .B2(n11063), .A(n7137), .ZN(n11226) );
  AND2_X1 U7780 ( .A1(n11619), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n7137) );
  AND2_X1 U7781 ( .A1(n8459), .A2(n7189), .ZN(n7188) );
  AND2_X1 U7782 ( .A1(n7187), .A2(n8305), .ZN(n7186) );
  AND2_X1 U7783 ( .A1(n8303), .A2(n8304), .ZN(n7189) );
  AND2_X1 U7784 ( .A1(n13208), .A2(P2_DATAO_REG_17__SCAN_IN), .ZN(n7151) );
  AND2_X1 U7785 ( .A1(n9875), .A2(n7145), .ZN(n7144) );
  INV_X1 U7786 ( .A(n9938), .ZN(n7145) );
  NAND2_X1 U7787 ( .A1(n9873), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n7146) );
  XNOR2_X1 U7788 ( .A(n9874), .B(P2_DATAO_REG_13__SCAN_IN), .ZN(n9873) );
  INV_X1 U7789 ( .A(n9588), .ZN(n7131) );
  INV_X1 U7790 ( .A(n7130), .ZN(n7129) );
  OAI21_X1 U7791 ( .B1(n7133), .B2(n6498), .A(n7135), .ZN(n7130) );
  NAND2_X1 U7792 ( .A1(P1_DATAO_REG_7__SCAN_IN), .A2(n7136), .ZN(n7135) );
  NOR2_X1 U7793 ( .A1(n9607), .A2(n7134), .ZN(n7133) );
  INV_X1 U7794 ( .A(n9585), .ZN(n7134) );
  NAND2_X1 U7795 ( .A1(n9581), .A2(n9580), .ZN(n9584) );
  XNOR2_X1 U7796 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .ZN(n9583) );
  INV_X1 U7797 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n8453) );
  INV_X1 U7798 ( .A(n12011), .ZN(n9969) );
  NAND2_X1 U7799 ( .A1(n10386), .A2(n10584), .ZN(n7265) );
  OR2_X1 U7800 ( .A1(n12590), .A2(n12589), .ZN(n7439) );
  AND2_X1 U7801 ( .A1(n13350), .A2(n12571), .ZN(n7281) );
  NAND2_X1 U7802 ( .A1(n7279), .A2(n7282), .ZN(n7280) );
  INV_X1 U7803 ( .A(n12609), .ZN(n7255) );
  NAND2_X1 U7804 ( .A1(n7265), .A2(n7268), .ZN(n7260) );
  INV_X1 U7805 ( .A(n7268), .ZN(n7256) );
  INV_X1 U7806 ( .A(n10629), .ZN(n7267) );
  INV_X1 U7807 ( .A(n13432), .ZN(n13556) );
  INV_X1 U7808 ( .A(n10272), .ZN(n7261) );
  INV_X1 U7809 ( .A(n11999), .ZN(n7244) );
  NAND2_X1 U7810 ( .A1(n7238), .A2(n7237), .ZN(n13378) );
  AND2_X1 U7811 ( .A1(n7239), .A2(n12595), .ZN(n7237) );
  XNOR2_X1 U7812 ( .A(n9992), .B(n10769), .ZN(n9993) );
  INV_X1 U7813 ( .A(n7280), .ZN(n13407) );
  NOR3_X1 U7814 ( .A1(n9165), .A2(n9164), .A3(n9163), .ZN(n7445) );
  INV_X1 U7815 ( .A(n8664), .ZN(n9147) );
  NAND2_X1 U7816 ( .A1(n8664), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n8651) );
  NAND2_X1 U7817 ( .A1(n8568), .A2(n6933), .ZN(n6936) );
  AND2_X1 U7818 ( .A1(n13867), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n6933) );
  NAND2_X1 U7819 ( .A1(n9170), .A2(n9169), .ZN(n13521) );
  NAND2_X1 U7820 ( .A1(n7301), .A2(n15064), .ZN(n7298) );
  NAND2_X1 U7821 ( .A1(n9117), .A2(n9116), .ZN(n13763) );
  NOR2_X1 U7822 ( .A1(n13642), .A2(n6940), .ZN(n13561) );
  NAND2_X1 U7823 ( .A1(n6943), .A2(n6941), .ZN(n6940) );
  NOR2_X1 U7824 ( .A1(n13763), .A2(n13779), .ZN(n6941) );
  XNOR2_X1 U7825 ( .A(n13779), .B(n13585), .ZN(n13617) );
  NAND2_X1 U7826 ( .A1(n6517), .A2(n13549), .ZN(n13654) );
  NOR2_X1 U7827 ( .A1(n13669), .A2(n7401), .ZN(n7400) );
  INV_X1 U7828 ( .A(n13546), .ZN(n7401) );
  XNOR2_X1 U7829 ( .A(n13806), .B(n13580), .ZN(n13669) );
  OR2_X1 U7830 ( .A1(n13811), .A2(n13579), .ZN(n7295) );
  AND2_X1 U7831 ( .A1(n6930), .A2(n6929), .ZN(n6928) );
  INV_X1 U7832 ( .A(n13706), .ZN(n6930) );
  NAND2_X1 U7833 ( .A1(n13576), .A2(n13715), .ZN(n6929) );
  NAND2_X1 U7834 ( .A1(n13714), .A2(n13576), .ZN(n6926) );
  OR2_X1 U7835 ( .A1(n8986), .A2(n13394), .ZN(n9000) );
  NOR2_X1 U7836 ( .A1(n13714), .A2(n13715), .ZN(n13713) );
  AND2_X1 U7837 ( .A1(n13745), .A2(n13573), .ZN(n6910) );
  OR2_X1 U7838 ( .A1(n13745), .A2(n13566), .ZN(n13537) );
  NAND2_X1 U7839 ( .A1(n13743), .A2(n13742), .ZN(n13741) );
  OAI21_X1 U7840 ( .B1(n7407), .B2(n7410), .A(n7409), .ZN(n7404) );
  OR2_X1 U7841 ( .A1(n11802), .A2(n13435), .ZN(n11803) );
  AOI21_X1 U7842 ( .B1(n6915), .B2(n6914), .A(n6584), .ZN(n6913) );
  INV_X1 U7843 ( .A(n11245), .ZN(n6914) );
  NAND2_X1 U7844 ( .A1(n15078), .A2(n11249), .ZN(n7393) );
  NAND2_X1 U7845 ( .A1(n6520), .A2(n10953), .ZN(n7389) );
  NAND3_X1 U7846 ( .A1(n10949), .A2(n7390), .A3(n6520), .ZN(n7394) );
  NAND2_X1 U7847 ( .A1(n8823), .A2(n8822), .ZN(n11276) );
  NOR2_X1 U7848 ( .A1(n10983), .A2(n10769), .ZN(n10768) );
  INV_X1 U7849 ( .A(n10767), .ZN(n10343) );
  NAND2_X1 U7850 ( .A1(n8998), .A2(n8997), .ZN(n13817) );
  INV_X1 U7851 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n6908) );
  XNOR2_X1 U7852 ( .A(n8582), .B(P2_IR_REG_21__SCAN_IN), .ZN(n8611) );
  NAND2_X1 U7853 ( .A1(n8587), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8582) );
  NAND2_X1 U7854 ( .A1(n6840), .A2(n7497), .ZN(n6839) );
  NAND2_X1 U7855 ( .A1(n6831), .A2(n6830), .ZN(n6829) );
  INV_X1 U7856 ( .A(n9325), .ZN(n6830) );
  INV_X1 U7857 ( .A(n11762), .ZN(n6831) );
  NOR2_X1 U7858 ( .A1(n7454), .A2(n7097), .ZN(n7096) );
  INV_X1 U7859 ( .A(n13953), .ZN(n7097) );
  NOR2_X1 U7860 ( .A1(n7092), .A2(n7090), .ZN(n7089) );
  INV_X1 U7861 ( .A(n9413), .ZN(n7090) );
  INV_X1 U7862 ( .A(n7092), .ZN(n7088) );
  INV_X1 U7863 ( .A(n11193), .ZN(n6814) );
  AND2_X1 U7864 ( .A1(n9268), .A2(n9499), .ZN(n9501) );
  OAI21_X1 U7865 ( .B1(n14007), .B2(n7081), .A(n9368), .ZN(n7080) );
  OR2_X1 U7866 ( .A1(n9367), .A2(n9366), .ZN(n9368) );
  NAND2_X1 U7867 ( .A1(n7085), .A2(n9396), .ZN(n13911) );
  INV_X1 U7868 ( .A(n13913), .ZN(n7085) );
  NAND2_X1 U7869 ( .A1(n6511), .A2(n6832), .ZN(n6823) );
  NAND2_X1 U7870 ( .A1(n11461), .A2(n9321), .ZN(n9324) );
  OAI21_X2 U7871 ( .B1(n9324), .B2(n6822), .A(n6820), .ZN(n11820) );
  INV_X1 U7872 ( .A(n6823), .ZN(n6822) );
  AOI21_X1 U7873 ( .B1(n6825), .B2(n6823), .A(n6821), .ZN(n6820) );
  INV_X1 U7874 ( .A(n11822), .ZN(n6821) );
  NOR2_X1 U7875 ( .A1(n7893), .A2(n7892), .ZN(n7940) );
  NAND2_X1 U7876 ( .A1(n6808), .A2(n6537), .ZN(n6807) );
  INV_X1 U7877 ( .A(n9301), .ZN(n6808) );
  NAND2_X1 U7878 ( .A1(n10895), .A2(n9303), .ZN(n7101) );
  NOR2_X1 U7879 ( .A1(n7105), .A2(n7104), .ZN(n7103) );
  INV_X1 U7880 ( .A(n10691), .ZN(n7104) );
  NOR2_X1 U7881 ( .A1(n9303), .A2(n10895), .ZN(n7105) );
  NAND2_X1 U7882 ( .A1(n13883), .A2(n6560), .ZN(n14008) );
  AND2_X1 U7883 ( .A1(n8217), .A2(n8263), .ZN(n6692) );
  INV_X1 U7884 ( .A(n8151), .ZN(n7218) );
  NOR2_X1 U7885 ( .A1(n8154), .A2(n8151), .ZN(n7219) );
  NOR2_X1 U7886 ( .A1(n8272), .A2(n8271), .ZN(n6715) );
  NOR2_X1 U7887 ( .A1(n8258), .A2(n6667), .ZN(n8253) );
  OR2_X1 U7888 ( .A1(n8252), .A2(n6668), .ZN(n6667) );
  AND2_X1 U7889 ( .A1(n14138), .A2(n14146), .ZN(n7363) );
  INV_X1 U7890 ( .A(n7361), .ZN(n7360) );
  NAND2_X1 U7891 ( .A1(n6895), .A2(n6571), .ZN(n14136) );
  INV_X1 U7892 ( .A(n14220), .ZN(n6895) );
  INV_X1 U7893 ( .A(n6897), .ZN(n6896) );
  AND2_X1 U7894 ( .A1(n14175), .A2(n14319), .ZN(n6770) );
  NAND2_X1 U7895 ( .A1(n14148), .A2(n9541), .ZN(n14130) );
  NAND2_X1 U7896 ( .A1(n14146), .A2(n6848), .ZN(n6845) );
  NAND2_X1 U7897 ( .A1(n8149), .A2(n6847), .ZN(n6846) );
  NOR2_X1 U7898 ( .A1(n14146), .A2(n6848), .ZN(n6847) );
  NAND2_X1 U7899 ( .A1(n14215), .A2(n7072), .ZN(n14169) );
  INV_X1 U7900 ( .A(n14174), .ZN(n14213) );
  NAND2_X1 U7901 ( .A1(n14251), .A2(n9492), .ZN(n14234) );
  AOI21_X1 U7902 ( .B1(n6781), .B2(n11832), .A(n6538), .ZN(n6779) );
  NAND2_X1 U7903 ( .A1(n11839), .A2(n11838), .ZN(n11837) );
  NAND2_X1 U7904 ( .A1(n11598), .A2(n7356), .ZN(n11640) );
  INV_X1 U7905 ( .A(n9480), .ZN(n7357) );
  AND2_X1 U7906 ( .A1(n11477), .A2(n6775), .ZN(n6774) );
  OR2_X1 U7907 ( .A1(n11413), .A2(n6776), .ZN(n6775) );
  INV_X1 U7908 ( .A(n9479), .ZN(n6776) );
  XNOR2_X1 U7909 ( .A(n11571), .B(n11352), .ZN(n11413) );
  NAND2_X1 U7910 ( .A1(n11359), .A2(n9478), .ZN(n11414) );
  NAND2_X1 U7911 ( .A1(n11413), .A2(n11414), .ZN(n11412) );
  INV_X1 U7912 ( .A(n9477), .ZN(n7352) );
  INV_X1 U7913 ( .A(n7351), .ZN(n7350) );
  OAI21_X1 U7914 ( .B1(n11231), .B2(n7352), .A(n11161), .ZN(n7351) );
  AND4_X1 U7915 ( .A1(n7717), .A2(n7716), .A3(n7715), .A4(n7714), .ZN(n11465)
         );
  INV_X1 U7916 ( .A(n14038), .ZN(n11241) );
  NAND2_X1 U7917 ( .A1(n11232), .A2(n11231), .ZN(n11230) );
  INV_X1 U7918 ( .A(n14324), .ZN(n14282) );
  NAND2_X1 U7919 ( .A1(n10597), .A2(n10596), .ZN(n12553) );
  AND2_X1 U7920 ( .A1(n9552), .A2(n6639), .ZN(n6863) );
  NAND2_X1 U7921 ( .A1(n12560), .A2(n14848), .ZN(n7077) );
  AND2_X1 U7922 ( .A1(n12558), .A2(n12552), .ZN(n9552) );
  NAND2_X1 U7923 ( .A1(n8214), .A2(n8213), .ZN(n12555) );
  AND2_X1 U7924 ( .A1(n14482), .A2(n9667), .ZN(n14394) );
  AND2_X1 U7925 ( .A1(n7559), .A2(n6751), .ZN(n6750) );
  NAND2_X1 U7926 ( .A1(n9435), .A2(n9434), .ZN(n9653) );
  AND2_X1 U7927 ( .A1(n7367), .A2(n7487), .ZN(n7059) );
  AND2_X1 U7928 ( .A1(n6836), .A2(P1_IR_REG_26__SCAN_IN), .ZN(n6835) );
  OR2_X1 U7929 ( .A1(n6530), .A2(n7672), .ZN(n6836) );
  NAND2_X1 U7930 ( .A1(n7060), .A2(n6543), .ZN(n8284) );
  AND2_X1 U7931 ( .A1(n6499), .A2(n7114), .ZN(n6837) );
  NAND2_X1 U7932 ( .A1(n8022), .A2(n8021), .ZN(n8055) );
  XNOR2_X1 U7933 ( .A(n8055), .B(n8056), .ZN(n9018) );
  XNOR2_X1 U7934 ( .A(n7793), .B(n7792), .ZN(n9932) );
  INV_X1 U7935 ( .A(n6878), .ZN(n14535) );
  NAND2_X1 U7936 ( .A1(n14597), .A2(n14596), .ZN(n7122) );
  INV_X1 U7937 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n14557) );
  INV_X1 U7938 ( .A(n6867), .ZN(n14565) );
  OAI21_X1 U7939 ( .B1(n14598), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n6540), .ZN(
        n6867) );
  NAND2_X1 U7940 ( .A1(n14564), .A2(n14563), .ZN(n14504) );
  NAND2_X1 U7941 ( .A1(n6874), .A2(n14900), .ZN(n6873) );
  INV_X1 U7942 ( .A(n14773), .ZN(n6874) );
  NAND2_X1 U7943 ( .A1(n14773), .A2(P2_ADDR_REG_13__SCAN_IN), .ZN(n6872) );
  NAND2_X1 U7944 ( .A1(n7194), .A2(n7193), .ZN(n12630) );
  AOI21_X1 U7945 ( .B1(n12218), .B2(n7203), .A(n7195), .ZN(n7194) );
  INV_X1 U7946 ( .A(n7199), .ZN(n7195) );
  INV_X1 U7947 ( .A(n12967), .ZN(n12937) );
  INV_X1 U7948 ( .A(n12960), .ZN(n13078) );
  CLKBUF_X1 U7949 ( .A(n11784), .Z(n6685) );
  AND2_X1 U7950 ( .A1(n12186), .A2(n12185), .ZN(n12658) );
  NAND2_X1 U7951 ( .A1(n12192), .A2(n12191), .ZN(n13086) );
  NAND2_X1 U7952 ( .A1(n12240), .A2(n12239), .ZN(n13070) );
  AND4_X1 U7953 ( .A1(n12145), .A2(n12144), .A3(n12143), .A4(n12142), .ZN(
        n13014) );
  INV_X1 U7954 ( .A(n12918), .ZN(n13066) );
  AND4_X1 U7955 ( .A1(n11711), .A2(n11710), .A3(n11709), .A4(n11708), .ZN(
        n12737) );
  NAND2_X1 U7956 ( .A1(n7455), .A2(n12544), .ZN(n6676) );
  NAND2_X1 U7957 ( .A1(n12542), .A2(n12541), .ZN(n12543) );
  NAND2_X1 U7958 ( .A1(n12248), .A2(n12247), .ZN(n12909) );
  NAND2_X1 U7959 ( .A1(n12200), .A2(n12199), .ZN(n12988) );
  INV_X1 U7960 ( .A(n12658), .ZN(n13000) );
  INV_X1 U7961 ( .A(n12737), .ZN(n12744) );
  OAI21_X1 U7962 ( .B1(n6490), .B2(n15099), .A(n6730), .ZN(n8350) );
  NAND2_X1 U7963 ( .A1(n6490), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n6730) );
  OR2_X1 U7964 ( .A1(n10398), .A2(n8382), .ZN(n6985) );
  INV_X1 U7965 ( .A(n10398), .ZN(n6986) );
  OR2_X1 U7966 ( .A1(n10850), .A2(n8481), .ZN(n6880) );
  AND2_X1 U7967 ( .A1(P3_U3897), .A2(n6485), .ZN(n15155) );
  NAND2_X1 U7968 ( .A1(n12812), .A2(n6724), .ZN(n6966) );
  AND2_X1 U7969 ( .A1(n8556), .A2(n6967), .ZN(n6724) );
  AOI21_X1 U7970 ( .B1(n13321), .B2(n12311), .A(n12320), .ZN(n14658) );
  XNOR2_X1 U7971 ( .A(n12834), .B(n12835), .ZN(n13056) );
  NOR2_X1 U7972 ( .A1(n12901), .A2(n6741), .ZN(n13065) );
  NAND2_X1 U7973 ( .A1(n6743), .A2(n6742), .ZN(n6741) );
  INV_X1 U7974 ( .A(n12902), .ZN(n6742) );
  NAND2_X1 U7975 ( .A1(n11943), .A2(n11942), .ZN(n14667) );
  AND3_X1 U7976 ( .A1(n11209), .A2(n11208), .A3(n11207), .ZN(n15249) );
  NAND2_X1 U7977 ( .A1(n8504), .A2(n8503), .ZN(n13053) );
  INV_X1 U7978 ( .A(n8528), .ZN(n11074) );
  MUX2_X1 U7979 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8345), .S(
        P3_IR_REG_1__SCAN_IN), .Z(n8346) );
  NAND2_X1 U7980 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(P3_IR_REG_31__SCAN_IN), .ZN(
        n8345) );
  OR2_X1 U7981 ( .A1(n9777), .A2(n8678), .ZN(n8803) );
  NAND2_X1 U7982 ( .A1(n13417), .A2(n12604), .ZN(n13337) );
  INV_X1 U7983 ( .A(n7263), .ZN(n10388) );
  AND2_X1 U7984 ( .A1(n9977), .A2(n14996), .ZN(n13415) );
  NAND4_X2 U7985 ( .A1(n8570), .A2(n8571), .A3(n8573), .A4(n8572), .ZN(n9205)
         );
  NAND2_X1 U7986 ( .A1(n8683), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n8572) );
  NAND2_X1 U7987 ( .A1(n15016), .A2(n10339), .ZN(n14996) );
  AND2_X1 U7988 ( .A1(n13771), .A2(n13770), .ZN(n13772) );
  OR2_X1 U7989 ( .A1(n13789), .A2(n15061), .ZN(n6700) );
  AND2_X1 U7990 ( .A1(n6623), .A2(n6734), .ZN(n7230) );
  XNOR2_X1 U7991 ( .A(n9241), .B(n9240), .ZN(n11815) );
  NAND2_X1 U7992 ( .A1(n9239), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9241) );
  NAND2_X1 U7993 ( .A1(n13971), .A2(n9406), .ZN(n13895) );
  NAND2_X1 U7994 ( .A1(n8006), .A2(n8005), .ZN(n14271) );
  INV_X1 U7995 ( .A(n14033), .ZN(n11824) );
  OR2_X1 U7996 ( .A1(n9371), .A2(n9370), .ZN(n6796) );
  NAND2_X1 U7997 ( .A1(n13942), .A2(n13943), .ZN(n6797) );
  INV_X1 U7998 ( .A(n6803), .ZN(n6802) );
  OAI21_X1 U7999 ( .B1(n12053), .B2(n9432), .A(n13995), .ZN(n6803) );
  NAND2_X1 U8000 ( .A1(n13923), .A2(n12051), .ZN(n6804) );
  NAND2_X1 U8001 ( .A1(n9458), .A2(n14307), .ZN(n14018) );
  OAI21_X1 U8002 ( .B1(n14272), .B2(n8119), .A(n7998), .ZN(n14248) );
  OAI21_X1 U8003 ( .B1(n14292), .B2(n8119), .A(n7975), .ZN(n14028) );
  NAND2_X1 U8004 ( .A1(n14236), .A2(n9494), .ZN(n14208) );
  INV_X1 U8005 ( .A(n14243), .ZN(n14817) );
  OR2_X1 U8006 ( .A1(n9457), .A2(n9553), .ZN(n14307) );
  NAND2_X1 U8007 ( .A1(n7728), .A2(n7727), .ZN(n11767) );
  NAND2_X1 U8008 ( .A1(n6792), .A2(n6791), .ZN(n6790) );
  INV_X1 U8009 ( .A(n14362), .ZN(n6791) );
  NAND2_X1 U8010 ( .A1(n14153), .A2(n14154), .ZN(n6794) );
  NOR2_X1 U8011 ( .A1(n6786), .A2(n14155), .ZN(n6785) );
  XNOR2_X1 U8012 ( .A(n14565), .B(n7125), .ZN(n14599) );
  INV_X1 U8013 ( .A(n14566), .ZN(n7125) );
  NOR2_X2 U8014 ( .A1(n14769), .A2(n14770), .ZN(n14768) );
  XNOR2_X1 U8015 ( .A(n6866), .B(n6865), .ZN(n14605) );
  INV_X1 U8016 ( .A(n14585), .ZN(n6865) );
  NAND2_X1 U8017 ( .A1(n6683), .A2(n6579), .ZN(n6682) );
  INV_X1 U8018 ( .A(n9504), .ZN(n6683) );
  OAI21_X1 U8019 ( .B1(n8176), .B2(n10900), .A(n6687), .ZN(n7588) );
  NAND2_X1 U8020 ( .A1(n8176), .A2(n10837), .ZN(n6687) );
  NAND2_X1 U8021 ( .A1(n8677), .A2(n8676), .ZN(n8696) );
  NAND2_X1 U8022 ( .A1(n7679), .A2(n7681), .ZN(n7221) );
  NAND2_X1 U8023 ( .A1(n6525), .A2(n8736), .ZN(n7437) );
  INV_X1 U8024 ( .A(n7754), .ZN(n7224) );
  NOR2_X1 U8025 ( .A1(n7226), .A2(n7754), .ZN(n7225) );
  NAND2_X1 U8026 ( .A1(n7435), .A2(n7434), .ZN(n7433) );
  INV_X1 U8027 ( .A(n8800), .ZN(n7435) );
  INV_X1 U8028 ( .A(n8830), .ZN(n7426) );
  INV_X1 U8029 ( .A(n8849), .ZN(n6710) );
  AND2_X1 U8030 ( .A1(n7914), .A2(n7915), .ZN(n7211) );
  NAND2_X1 U8031 ( .A1(n7213), .A2(n6531), .ZN(n7212) );
  AOI21_X1 U8032 ( .B1(n7945), .B2(n7944), .A(n7215), .ZN(n7214) );
  NAND2_X1 U8033 ( .A1(n7930), .A2(n7929), .ZN(n7215) );
  NAND2_X1 U8034 ( .A1(n6681), .A2(n6680), .ZN(n7453) );
  INV_X1 U8035 ( .A(n8907), .ZN(n6680) );
  NOR2_X1 U8036 ( .A1(n7419), .A2(n6558), .ZN(n7417) );
  AND2_X1 U8037 ( .A1(n7421), .A2(n7420), .ZN(n7419) );
  NAND2_X1 U8038 ( .A1(n8007), .A2(n8009), .ZN(n7223) );
  NAND2_X1 U8039 ( .A1(n8982), .A2(n8981), .ZN(n6694) );
  INV_X1 U8040 ( .A(n8980), .ZN(n6693) );
  NOR2_X1 U8041 ( .A1(n6526), .A2(n7424), .ZN(n7423) );
  NAND2_X1 U8042 ( .A1(n8044), .A2(n7229), .ZN(n7228) );
  NAND2_X1 U8043 ( .A1(n7414), .A2(n6549), .ZN(n7413) );
  AOI21_X1 U8044 ( .B1(n9037), .B2(n9033), .A(n6695), .ZN(n7412) );
  XNOR2_X1 U8045 ( .A(n9915), .B(n9502), .ZN(n7542) );
  NAND2_X1 U8046 ( .A1(n7542), .A2(n11614), .ZN(n8195) );
  NOR2_X1 U8047 ( .A1(n7983), .A2(n6856), .ZN(n6855) );
  INV_X1 U8048 ( .A(n7935), .ZN(n6856) );
  NAND2_X1 U8049 ( .A1(n7319), .A2(n6855), .ZN(n6853) );
  NAND2_X1 U8050 ( .A1(n6496), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n6982) );
  OR2_X1 U8051 ( .A1(n13053), .A2(n12367), .ZN(n12481) );
  INV_X1 U8052 ( .A(n13876), .ZN(n7094) );
  NAND2_X1 U8053 ( .A1(n8114), .A2(n8113), .ZN(n8135) );
  INV_X1 U8054 ( .A(n9520), .ZN(n7042) );
  INV_X1 U8055 ( .A(n7287), .ZN(n7286) );
  OAI21_X1 U8056 ( .B1(n7815), .B2(n7288), .A(n7832), .ZN(n7287) );
  INV_X1 U8057 ( .A(n7819), .ZN(n7288) );
  AOI21_X1 U8058 ( .B1(n12342), .B2(n12336), .A(n12341), .ZN(n12537) );
  AND2_X1 U8059 ( .A1(n12503), .A2(n12338), .ZN(n12339) );
  INV_X1 U8060 ( .A(n6958), .ZN(n8519) );
  NAND2_X1 U8061 ( .A1(n6989), .A2(n6987), .ZN(n8524) );
  NOR2_X1 U8062 ( .A1(n6988), .A2(n6588), .ZN(n6987) );
  INV_X1 U8063 ( .A(n6990), .ZN(n6988) );
  AOI21_X1 U8064 ( .B1(n10856), .B2(n10855), .A(n10854), .ZN(n10853) );
  INV_X1 U8065 ( .A(n12927), .ZN(n7018) );
  NAND2_X1 U8066 ( .A1(n12491), .A2(n12493), .ZN(n12859) );
  NAND2_X1 U8067 ( .A1(n7001), .A2(n12837), .ZN(n7000) );
  NOR2_X1 U8068 ( .A1(n11706), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n11945) );
  NOR2_X1 U8069 ( .A1(n11715), .A2(n7012), .ZN(n7011) );
  INV_X1 U8070 ( .A(n12525), .ZN(n7012) );
  INV_X1 U8071 ( .A(n12362), .ZN(n7014) );
  INV_X1 U8072 ( .A(P3_REG3_REG_12__SCAN_IN), .ZN(n11533) );
  OR2_X1 U8073 ( .A1(n14679), .A2(n12747), .ZN(n12425) );
  AND2_X1 U8074 ( .A1(n12425), .A2(n12424), .ZN(n12421) );
  INV_X1 U8075 ( .A(n7008), .ZN(n7007) );
  OAI21_X1 U8076 ( .B1(n12514), .B2(n7009), .A(n12408), .ZN(n7008) );
  INV_X1 U8077 ( .A(n12402), .ZN(n7009) );
  INV_X1 U8078 ( .A(P3_REG3_REG_8__SCAN_IN), .ZN(n11092) );
  INV_X1 U8079 ( .A(n12383), .ZN(n6995) );
  INV_X1 U8080 ( .A(P2_RD_REG_SCAN_IN), .ZN(n6841) );
  OR2_X1 U8081 ( .A1(n10215), .A2(n10214), .ZN(n10472) );
  OR2_X1 U8082 ( .A1(n13053), .A2(n12345), .ZN(n10482) );
  AOI21_X1 U8083 ( .B1(n7157), .B2(n7156), .A(n11741), .ZN(n11742) );
  AND2_X1 U8084 ( .A1(n11892), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n11741) );
  INV_X1 U8085 ( .A(n11740), .ZN(n7156) );
  NOR2_X1 U8086 ( .A1(n7192), .A2(P3_IR_REG_18__SCAN_IN), .ZN(n7190) );
  NAND2_X1 U8087 ( .A1(n8353), .A2(n8296), .ZN(n8372) );
  AOI21_X1 U8088 ( .B1(n7234), .B2(n7236), .A(n6510), .ZN(n7232) );
  NAND2_X1 U8089 ( .A1(n7303), .A2(n13559), .ZN(n7301) );
  INV_X1 U8090 ( .A(n6523), .ZN(n7306) );
  INV_X1 U8091 ( .A(n13583), .ZN(n7305) );
  INV_X1 U8092 ( .A(n13551), .ZN(n7381) );
  NOR2_X1 U8093 ( .A1(n13744), .A2(n13745), .ZN(n6704) );
  INV_X1 U8094 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n8790) );
  OR2_X1 U8095 ( .A1(n8791), .A2(n8790), .ZN(n8806) );
  XNOR2_X1 U8096 ( .A(n10357), .B(n10375), .ZN(n10356) );
  INV_X1 U8097 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n8574) );
  INV_X1 U8098 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n8659) );
  NOR2_X2 U8099 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n8617) );
  NAND3_X1 U8100 ( .A1(n7496), .A2(n12114), .A3(n6844), .ZN(n6843) );
  INV_X1 U8101 ( .A(P1_RD_REG_SCAN_IN), .ZN(n6844) );
  INV_X1 U8102 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n7710) );
  INV_X1 U8103 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n7654) );
  NOR2_X1 U8104 ( .A1(n11463), .A2(n6810), .ZN(n6809) );
  INV_X1 U8105 ( .A(n9314), .ZN(n6810) );
  INV_X1 U8106 ( .A(n11614), .ZN(n8179) );
  OR4_X1 U8107 ( .A1(n14192), .A2(n14210), .A3(n14252), .A4(n8249), .ZN(n8250)
         );
  XNOR2_X1 U8108 ( .A(n14438), .B(n8194), .ZN(n8252) );
  INV_X1 U8109 ( .A(n8148), .ZN(n6848) );
  OR2_X1 U8110 ( .A1(n14366), .A2(n14374), .ZN(n6898) );
  OR2_X1 U8111 ( .A1(n14158), .A2(n6898), .ZN(n6897) );
  NOR2_X1 U8112 ( .A1(n14254), .A2(n14385), .ZN(n14219) );
  NAND2_X1 U8113 ( .A1(n6779), .A2(n6780), .ZN(n6777) );
  OR2_X1 U8114 ( .A1(n14409), .A2(n14286), .ZN(n7966) );
  NOR2_X1 U8115 ( .A1(n11840), .A2(n14425), .ZN(n6903) );
  NOR2_X1 U8116 ( .A1(n11642), .A2(n13892), .ZN(n6905) );
  INV_X1 U8117 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n7807) );
  AND3_X1 U8118 ( .A1(n6892), .A2(n6891), .A3(n11233), .ZN(n11485) );
  AND2_X1 U8119 ( .A1(n11830), .A2(n6893), .ZN(n6892) );
  INV_X1 U8120 ( .A(n11360), .ZN(n9518) );
  INV_X1 U8121 ( .A(n11356), .ZN(n9519) );
  NOR2_X1 U8122 ( .A1(n11161), .A2(n7034), .ZN(n7033) );
  INV_X1 U8123 ( .A(n9516), .ZN(n7034) );
  NAND2_X1 U8124 ( .A1(n14294), .A2(n14461), .ZN(n14268) );
  NAND2_X1 U8125 ( .A1(n6753), .A2(n6752), .ZN(n6751) );
  INV_X1 U8126 ( .A(n10623), .ZN(n14834) );
  INV_X1 U8127 ( .A(n10620), .ZN(n10611) );
  NAND2_X1 U8128 ( .A1(n8083), .A2(n8082), .ZN(n8103) );
  NAND2_X1 U8129 ( .A1(n8004), .A2(n8003), .ZN(n8019) );
  OR2_X1 U8130 ( .A1(n8002), .A2(n10777), .ZN(n8003) );
  NAND2_X1 U8131 ( .A1(n7530), .A2(n7114), .ZN(n7113) );
  NAND2_X1 U8132 ( .A1(n6857), .A2(n7935), .ZN(n7984) );
  XNOR2_X1 U8133 ( .A(n7984), .B(SI_18_), .ZN(n7946) );
  OR2_X1 U8134 ( .A1(n7904), .A2(P1_IR_REG_17__SCAN_IN), .ZN(n7936) );
  INV_X1 U8135 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n7887) );
  CLKBUF_X1 U8136 ( .A(n7852), .Z(n7853) );
  OR2_X1 U8137 ( .A1(n7795), .A2(P1_IR_REG_11__SCAN_IN), .ZN(n7796) );
  NAND2_X1 U8138 ( .A1(n7313), .A2(n7315), .ZN(n7745) );
  AOI21_X1 U8139 ( .B1(n7722), .B2(n7317), .A(n7316), .ZN(n7315) );
  INV_X1 U8140 ( .A(n7742), .ZN(n7316) );
  INV_X1 U8141 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n7457) );
  NAND2_X1 U8142 ( .A1(n6484), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n6712) );
  NAND2_X1 U8143 ( .A1(n7117), .A2(n14532), .ZN(n7115) );
  INV_X1 U8144 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n14489) );
  NOR2_X1 U8145 ( .A1(n14491), .A2(n14492), .ZN(n14493) );
  XNOR2_X1 U8146 ( .A(n14493), .B(n15145), .ZN(n14548) );
  NOR2_X1 U8147 ( .A1(n14500), .A2(n14499), .ZN(n14528) );
  AOI21_X1 U8148 ( .B1(n7203), .B2(n7200), .A(n6509), .ZN(n7199) );
  INV_X1 U8149 ( .A(n7204), .ZN(n7200) );
  INV_X1 U8150 ( .A(n12260), .ZN(n7208) );
  NOR2_X1 U8151 ( .A1(n7201), .A2(n12977), .ZN(n7198) );
  NAND2_X1 U8152 ( .A1(n12495), .A2(n12497), .ZN(n12862) );
  NAND2_X1 U8153 ( .A1(n12696), .A2(n7164), .ZN(n12652) );
  NOR2_X1 U8154 ( .A1(n12655), .A2(n7165), .ZN(n7164) );
  INV_X1 U8155 ( .A(n12189), .ZN(n7165) );
  OR2_X1 U8156 ( .A1(n7178), .A2(n11915), .ZN(n7176) );
  NAND2_X1 U8157 ( .A1(n11496), .A2(n6568), .ZN(n11588) );
  OR2_X1 U8158 ( .A1(n11095), .A2(P3_REG3_REG_9__SCAN_IN), .ZN(n11316) );
  OR2_X1 U8159 ( .A1(n11675), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n11706) );
  INV_X1 U8160 ( .A(P3_REG3_REG_11__SCAN_IN), .ZN(n11431) );
  INV_X1 U8161 ( .A(n12736), .ZN(n12720) );
  AOI21_X1 U8162 ( .B1(n7183), .B2(n7182), .A(n6634), .ZN(n7181) );
  INV_X1 U8163 ( .A(n7185), .ZN(n7182) );
  NAND2_X1 U8164 ( .A1(n12504), .A2(n12505), .ZN(n7163) );
  NAND2_X1 U8165 ( .A1(n8320), .A2(n8319), .ZN(n10225) );
  OAI21_X1 U8166 ( .B1(n6490), .B2(P3_REG2_REG_1__SCAN_IN), .A(n6767), .ZN(
        n8347) );
  NAND2_X1 U8167 ( .A1(n6488), .A2(n8343), .ZN(n6767) );
  AOI22_X1 U8168 ( .A1(n10450), .A2(P3_REG1_REG_2__SCAN_IN), .B1(n8351), .B2(
        n6496), .ZN(n10414) );
  NOR2_X1 U8169 ( .A1(n10415), .A2(n10414), .ZN(n10413) );
  NOR2_X1 U8170 ( .A1(n10434), .A2(n11013), .ZN(n10433) );
  OAI21_X1 U8171 ( .B1(n10436), .B2(n7062), .A(n7061), .ZN(n15112) );
  NAND2_X1 U8172 ( .A1(n7063), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n7062) );
  NAND2_X1 U8173 ( .A1(n8470), .A2(n7063), .ZN(n7061) );
  INV_X1 U8174 ( .A(n15113), .ZN(n7063) );
  NOR2_X1 U8175 ( .A1(n10436), .A2(n8362), .ZN(n10435) );
  INV_X1 U8176 ( .A(n8473), .ZN(n7067) );
  OAI21_X1 U8177 ( .B1(n15135), .B2(n7066), .A(n7065), .ZN(n10400) );
  NAND2_X1 U8178 ( .A1(n7069), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n7066) );
  INV_X1 U8179 ( .A(n10401), .ZN(n7069) );
  INV_X1 U8180 ( .A(n10533), .ZN(n7056) );
  OAI21_X1 U8181 ( .B1(n7055), .B2(n15160), .A(n7054), .ZN(n8480) );
  NAND2_X1 U8182 ( .A1(n10533), .A2(n7058), .ZN(n7054) );
  NAND2_X1 U8183 ( .A1(n8476), .A2(n7058), .ZN(n7055) );
  NAND2_X1 U8184 ( .A1(n11206), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n7058) );
  NOR2_X1 U8185 ( .A1(n11513), .A2(n11514), .ZN(n11512) );
  OR2_X1 U8186 ( .A1(n12756), .A2(n8542), .ZN(n6957) );
  NAND2_X1 U8187 ( .A1(n12759), .A2(n6630), .ZN(n12780) );
  NOR2_X1 U8188 ( .A1(n12773), .A2(n6954), .ZN(n8543) );
  NOR2_X1 U8189 ( .A1(n11941), .A2(n6955), .ZN(n6954) );
  NAND2_X1 U8190 ( .A1(n7053), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n7052) );
  NAND2_X1 U8191 ( .A1(n8491), .A2(n7053), .ZN(n7051) );
  OR2_X1 U8192 ( .A1(n8446), .A2(P3_IR_REG_15__SCAN_IN), .ZN(n8449) );
  INV_X1 U8193 ( .A(n6726), .ZN(n8448) );
  OR2_X1 U8194 ( .A1(n14638), .A2(n6653), .ZN(n6973) );
  OAI21_X1 U8195 ( .B1(n12792), .B2(n6522), .A(n7036), .ZN(n12817) );
  INV_X1 U8196 ( .A(n7037), .ZN(n7036) );
  OAI21_X1 U8197 ( .B1(n6522), .B2(P3_REG1_REG_17__SCAN_IN), .A(n12814), .ZN(
        n7037) );
  AND2_X1 U8198 ( .A1(n12792), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n12815) );
  INV_X1 U8199 ( .A(n8497), .ZN(n6888) );
  NOR2_X1 U8200 ( .A1(n12805), .A2(n6536), .ZN(n8462) );
  NAND2_X1 U8201 ( .A1(n8550), .A2(n6970), .ZN(n6969) );
  AND2_X1 U8202 ( .A1(n12508), .A2(n12507), .ZN(n12863) );
  INV_X1 U8203 ( .A(n12862), .ZN(n12887) );
  OAI21_X1 U8204 ( .B1(n12925), .B2(n7330), .A(n7326), .ZN(n12900) );
  INV_X1 U8205 ( .A(n7327), .ZN(n7326) );
  NAND2_X1 U8206 ( .A1(n13063), .A2(n15204), .ZN(n6743) );
  AND2_X1 U8207 ( .A1(n12471), .A2(n12473), .ZN(n12939) );
  NOR2_X1 U8208 ( .A1(n12206), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n12207) );
  INV_X1 U8209 ( .A(n7025), .ZN(n7024) );
  OAI21_X1 U8210 ( .B1(n6500), .B2(n7026), .A(n12351), .ZN(n7025) );
  NOR2_X1 U8211 ( .A1(n6582), .A2(n7322), .ZN(n7321) );
  INV_X1 U8212 ( .A(n12845), .ZN(n7322) );
  AOI21_X1 U8213 ( .B1(n12441), .B2(n7003), .A(n7002), .ZN(n7001) );
  INV_X1 U8214 ( .A(n11988), .ZN(n7003) );
  INV_X1 U8215 ( .A(n12445), .ZN(n7002) );
  AND2_X1 U8216 ( .A1(n11396), .A2(n11395), .ZN(n11589) );
  AND3_X1 U8217 ( .A1(n11309), .A2(n11308), .A3(n11307), .ZN(n12413) );
  AND4_X1 U8218 ( .A1(n11099), .A2(n11098), .A3(n11097), .A4(n11096), .ZN(
        n11502) );
  NOR2_X1 U8219 ( .A1(n12405), .A2(n11213), .ZN(n6670) );
  INV_X1 U8220 ( .A(n12411), .ZN(n12412) );
  NAND2_X1 U8221 ( .A1(n11204), .A2(n12402), .ZN(n11314) );
  NAND2_X1 U8222 ( .A1(n11090), .A2(n12514), .ZN(n11204) );
  NAND2_X1 U8223 ( .A1(n11070), .A2(n11069), .ZN(n11131) );
  NAND2_X1 U8224 ( .A1(n11070), .A2(n7335), .ZN(n11215) );
  OR2_X1 U8225 ( .A1(n10929), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n11075) );
  NAND2_X1 U8226 ( .A1(n11030), .A2(n7337), .ZN(n11070) );
  AND4_X1 U8227 ( .A1(n10812), .A2(n10811), .A3(n10810), .A4(n10809), .ZN(
        n11128) );
  OR2_X1 U8228 ( .A1(n10791), .A2(n10236), .ZN(n10238) );
  OR2_X1 U8229 ( .A1(n12290), .A2(n8343), .ZN(n10237) );
  INV_X1 U8230 ( .A(n15194), .ZN(n15173) );
  INV_X1 U8231 ( .A(n12345), .ZN(n12539) );
  NAND2_X1 U8232 ( .A1(n15202), .A2(n15191), .ZN(n15193) );
  NAND2_X1 U8233 ( .A1(n12545), .A2(n11001), .ZN(n15197) );
  INV_X1 U8234 ( .A(n15200), .ZN(n15178) );
  INV_X1 U8235 ( .A(P3_ADDR_REG_8__SCAN_IN), .ZN(n14503) );
  INV_X1 U8236 ( .A(n11210), .ZN(n15244) );
  AND2_X1 U8237 ( .A1(n10225), .A2(n13318), .ZN(n13295) );
  INV_X1 U8238 ( .A(n14680), .ZN(n15214) );
  INV_X1 U8239 ( .A(n13318), .ZN(n10231) );
  NAND2_X1 U8240 ( .A1(n10202), .A2(n10201), .ZN(n10471) );
  AND2_X1 U8241 ( .A1(n6544), .A2(n7346), .ZN(n7345) );
  INV_X1 U8242 ( .A(P3_IR_REG_29__SCAN_IN), .ZN(n7346) );
  NAND2_X1 U8243 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n12088), .ZN(n12089) );
  NAND2_X1 U8244 ( .A1(n12087), .A2(n7161), .ZN(n12263) );
  NAND2_X1 U8245 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(n12008), .ZN(n7161) );
  NAND2_X1 U8246 ( .A1(n12085), .A2(n12086), .ZN(n12087) );
  INV_X1 U8247 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n8324) );
  NAND2_X1 U8248 ( .A1(n8325), .A2(n8324), .ZN(n9918) );
  INV_X1 U8249 ( .A(n7341), .ZN(n7340) );
  NOR2_X1 U8250 ( .A1(n8310), .A2(P3_IR_REG_19__SCAN_IN), .ZN(n7341) );
  INV_X1 U8251 ( .A(n7172), .ZN(n8504) );
  NAND2_X1 U8252 ( .A1(P2_DATAO_REG_19__SCAN_IN), .A2(n7142), .ZN(n7141) );
  CLKBUF_X1 U8253 ( .A(n8457), .Z(n8458) );
  AND2_X1 U8254 ( .A1(n7153), .A2(n7152), .ZN(n10465) );
  NAND2_X1 U8255 ( .A1(n10976), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n7152) );
  AND2_X1 U8256 ( .A1(n8337), .A2(n8299), .ZN(n8333) );
  NAND2_X1 U8257 ( .A1(n9643), .A2(n7150), .ZN(n7148) );
  AND2_X1 U8258 ( .A1(n6642), .A2(n9642), .ZN(n7150) );
  AOI21_X1 U8259 ( .B1(n7129), .B2(n7127), .A(n6592), .ZN(n7126) );
  CLKBUF_X1 U8260 ( .A(n8372), .Z(n8373) );
  OAI21_X1 U8261 ( .B1(n9605), .B2(n9578), .A(n9579), .ZN(n9596) );
  XNOR2_X1 U8262 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .ZN(n9595) );
  XNOR2_X1 U8263 ( .A(n9238), .B(n9237), .ZN(n9982) );
  INV_X1 U8264 ( .A(n14990), .ZN(n6945) );
  AND2_X1 U8265 ( .A1(n7235), .A2(n13360), .ZN(n7234) );
  NAND2_X1 U8266 ( .A1(n13388), .A2(n13387), .ZN(n7235) );
  INV_X1 U8267 ( .A(n13550), .ZN(n13581) );
  NAND2_X1 U8268 ( .A1(n8916), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8930) );
  INV_X1 U8269 ( .A(n8917), .ZN(n8916) );
  NAND2_X1 U8270 ( .A1(n7240), .A2(n12591), .ZN(n7239) );
  NAND2_X1 U8271 ( .A1(n13343), .A2(n13344), .ZN(n7238) );
  OR2_X1 U8272 ( .A1(n10911), .A2(n10910), .ZN(n7276) );
  NAND2_X1 U8273 ( .A1(n11632), .A2(n11631), .ZN(n7273) );
  OR2_X1 U8274 ( .A1(n11632), .A2(n11631), .ZN(n7274) );
  OR2_X1 U8275 ( .A1(n9024), .A2(n13403), .ZN(n9044) );
  OR2_X1 U8276 ( .A1(n10910), .A2(n6505), .ZN(n7275) );
  INV_X1 U8277 ( .A(n13447), .ZN(n10357) );
  NAND2_X1 U8278 ( .A1(n12568), .A2(n12567), .ZN(n13409) );
  INV_X1 U8279 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n11727) );
  NAND2_X1 U8280 ( .A1(n8611), .A2(n11523), .ZN(n9991) );
  INV_X1 U8281 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n6749) );
  NAND2_X1 U8282 ( .A1(n6494), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n8571) );
  OR2_X1 U8283 ( .A1(n8858), .A2(P2_IR_REG_13__SCAN_IN), .ZN(n8894) );
  NOR2_X1 U8284 ( .A1(n7300), .A2(n7302), .ZN(n7299) );
  INV_X1 U8285 ( .A(n7303), .ZN(n7300) );
  OAI21_X1 U8286 ( .B1(n13555), .B2(n7396), .A(n7395), .ZN(n13605) );
  INV_X1 U8287 ( .A(n7397), .ZN(n7396) );
  AOI21_X1 U8288 ( .B1(n7397), .B2(n13553), .A(n6580), .ZN(n7395) );
  NAND2_X1 U8289 ( .A1(n6943), .A2(n6944), .ZN(n6942) );
  NOR2_X1 U8290 ( .A1(n13617), .A2(n7398), .ZN(n7397) );
  INV_X1 U8291 ( .A(n13557), .ZN(n7398) );
  AND2_X1 U8292 ( .A1(n7310), .A2(n6616), .ZN(n7308) );
  NAND2_X1 U8293 ( .A1(n13666), .A2(n6523), .ZN(n7309) );
  OR2_X1 U8294 ( .A1(n13647), .A2(n13646), .ZN(n7310) );
  NAND2_X1 U8295 ( .A1(n13666), .A2(n13665), .ZN(n13664) );
  NOR2_X1 U8296 ( .A1(n6504), .A2(n13577), .ZN(n6927) );
  NAND2_X1 U8297 ( .A1(n8999), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n9024) );
  INV_X1 U8298 ( .A(n9000), .ZN(n8999) );
  NOR2_X1 U8299 ( .A1(n13729), .A2(n13822), .ZN(n13718) );
  NAND2_X1 U8300 ( .A1(n13718), .A2(n13699), .ZN(n13701) );
  NAND2_X1 U8301 ( .A1(n8968), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8986) );
  AOI21_X1 U8302 ( .B1(n7385), .B2(n7387), .A(n7383), .ZN(n7382) );
  INV_X1 U8303 ( .A(n13539), .ZN(n7383) );
  NAND2_X1 U8304 ( .A1(n6704), .A2(n6703), .ZN(n13729) );
  INV_X1 U8305 ( .A(n6704), .ZN(n13746) );
  NAND2_X1 U8306 ( .A1(n6911), .A2(n11962), .ZN(n13572) );
  NAND2_X1 U8307 ( .A1(n11804), .A2(n7407), .ZN(n7406) );
  INV_X1 U8308 ( .A(n6950), .ZN(n11797) );
  NOR2_X1 U8309 ( .A1(n14735), .A2(n13436), .ZN(n6939) );
  AND2_X1 U8310 ( .A1(n14702), .A2(n13436), .ZN(n11549) );
  NAND2_X1 U8311 ( .A1(n6951), .A2(n14735), .ZN(n14707) );
  OR2_X1 U8312 ( .A1(n8877), .A2(n11671), .ZN(n8897) );
  INV_X1 U8313 ( .A(n11548), .ZN(n14705) );
  NOR2_X1 U8314 ( .A1(n7388), .A2(n6563), .ZN(n6748) );
  OR2_X1 U8315 ( .A1(n8840), .A2(n8839), .ZN(n8864) );
  NOR2_X1 U8316 ( .A1(n10950), .A2(n11276), .ZN(n14720) );
  NAND2_X1 U8317 ( .A1(n6946), .A2(n10968), .ZN(n10950) );
  INV_X1 U8318 ( .A(n10877), .ZN(n6946) );
  NAND2_X1 U8319 ( .A1(n6948), .A2(n6947), .ZN(n10877) );
  INV_X1 U8320 ( .A(n6921), .ZN(n6920) );
  NOR2_X1 U8321 ( .A1(n10710), .A2(n6922), .ZN(n6921) );
  AND2_X1 U8322 ( .A1(n15058), .A2(n13445), .ZN(n7375) );
  NAND2_X1 U8323 ( .A1(n6702), .A2(n6701), .ZN(n14981) );
  INV_X1 U8324 ( .A(n14980), .ZN(n6702) );
  NAND2_X1 U8325 ( .A1(n15042), .A2(n10768), .ZN(n14980) );
  NAND2_X1 U8326 ( .A1(n8637), .A2(n9168), .ZN(n8647) );
  NOR2_X1 U8327 ( .A1(n9669), .A2(n9723), .ZN(n8645) );
  NAND2_X1 U8328 ( .A1(n15026), .A2(n6945), .ZN(n10983) );
  NOR2_X1 U8329 ( .A1(n14989), .A2(n10348), .ZN(n10339) );
  OR2_X1 U8330 ( .A1(n13764), .A2(n15077), .ZN(n7450) );
  NAND2_X1 U8331 ( .A1(n9023), .A2(n9022), .ZN(n13811) );
  INV_X1 U8332 ( .A(n15077), .ZN(n15069) );
  CLKBUF_X1 U8333 ( .A(n10346), .Z(n10347) );
  OR2_X1 U8334 ( .A1(n6713), .A2(n10348), .ZN(n15076) );
  AND2_X1 U8335 ( .A1(n9969), .A2(n9968), .ZN(n15006) );
  CLKBUF_X1 U8336 ( .A(n9250), .Z(n9251) );
  AND2_X1 U8337 ( .A1(n9248), .A2(n9242), .ZN(n9966) );
  NAND2_X1 U8338 ( .A1(n9228), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9238) );
  OR2_X1 U8339 ( .A1(n9227), .A2(P2_IR_REG_22__SCAN_IN), .ZN(n9228) );
  INV_X1 U8340 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n9237) );
  XNOR2_X1 U8341 ( .A(n8584), .B(n8580), .ZN(n8610) );
  NAND2_X1 U8342 ( .A1(n8583), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8584) );
  OR2_X1 U8343 ( .A1(n8925), .A2(P2_IR_REG_10__SCAN_IN), .ZN(n8832) );
  OR2_X1 U8344 ( .A1(n8725), .A2(P2_IR_REG_6__SCAN_IN), .ZN(n8761) );
  OR2_X1 U8345 ( .A1(n8697), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n8699) );
  NAND2_X1 U8346 ( .A1(n7098), .A2(n6565), .ZN(n7095) );
  NOR2_X1 U8347 ( .A1(n7808), .A2(n7807), .ZN(n7843) );
  NOR2_X1 U8348 ( .A1(n7711), .A2(n7710), .ZN(n7760) );
  INV_X1 U8349 ( .A(n14043), .ZN(n9282) );
  NAND2_X1 U8350 ( .A1(n7108), .A2(n9378), .ZN(n13904) );
  OR2_X1 U8351 ( .A1(n7655), .A2(n7654), .ZN(n7683) );
  NOR2_X1 U8352 ( .A1(n7993), .A2(n13915), .ZN(n8010) );
  NAND2_X1 U8353 ( .A1(n9300), .A2(n9299), .ZN(n9301) );
  OR2_X1 U8354 ( .A1(n7872), .A2(n7871), .ZN(n7893) );
  INV_X1 U8355 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n7892) );
  OAI211_X1 U8356 ( .C1(n9288), .C2(n9273), .A(n9272), .B(n9271), .ZN(n10133)
         );
  OR2_X1 U8357 ( .A1(n7969), .A2(n13966), .ZN(n7993) );
  OR2_X1 U8358 ( .A1(n7957), .A2(n12111), .ZN(n7969) );
  AND2_X1 U8359 ( .A1(n6542), .A2(n9378), .ZN(n7107) );
  AOI22_X1 U8360 ( .A1(n12057), .A2(n14043), .B1(n9275), .B2(n10623), .ZN(
        n9283) );
  INV_X1 U8361 ( .A(n9287), .ZN(n12061) );
  AND2_X1 U8362 ( .A1(n10594), .A2(n9562), .ZN(n9463) );
  AND2_X1 U8363 ( .A1(n7843), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n7857) );
  AND2_X1 U8364 ( .A1(n14483), .A2(n8179), .ZN(n9666) );
  NAND4_X1 U8365 ( .A1(n7521), .A2(n7519), .A3(n7520), .A4(n7522), .ZN(n9913)
         );
  OR2_X1 U8366 ( .A1(n8201), .A2(n7518), .ZN(n7521) );
  NOR2_X1 U8367 ( .A1(n14220), .A2(n6898), .ZN(n14181) );
  NOR2_X1 U8368 ( .A1(n14220), .A2(n6897), .ZN(n14156) );
  OAI21_X1 U8369 ( .B1(n14234), .B2(n7365), .A(n6587), .ZN(n14193) );
  NAND2_X1 U8370 ( .A1(n9493), .A2(n9495), .ZN(n7365) );
  INV_X1 U8371 ( .A(n9495), .ZN(n7364) );
  NOR2_X1 U8372 ( .A1(n14220), .A2(n14374), .ZN(n14194) );
  NAND2_X1 U8373 ( .A1(n14219), .A2(n14379), .ZN(n14220) );
  NAND2_X1 U8374 ( .A1(n7366), .A2(n9493), .ZN(n14236) );
  XNOR2_X1 U8375 ( .A(n14385), .B(n14249), .ZN(n14233) );
  OR2_X1 U8376 ( .A1(n14268), .A2(n14394), .ZN(n14254) );
  NAND2_X1 U8377 ( .A1(n6771), .A2(n9491), .ZN(n14253) );
  NAND2_X1 U8378 ( .A1(n7353), .A2(n6572), .ZN(n6771) );
  XNOR2_X1 U8379 ( .A(n14394), .B(n14265), .ZN(n14252) );
  AOI21_X1 U8380 ( .B1(n7045), .B2(n7047), .A(n6502), .ZN(n7044) );
  NOR2_X1 U8381 ( .A1(n14311), .A2(n14404), .ZN(n14294) );
  NAND2_X1 U8382 ( .A1(n14310), .A2(n9549), .ZN(n14311) );
  INV_X1 U8383 ( .A(n6781), .ZN(n6780) );
  NOR2_X1 U8384 ( .A1(n14327), .A2(n14414), .ZN(n14310) );
  INV_X1 U8385 ( .A(n11831), .ZN(n12035) );
  NOR2_X1 U8386 ( .A1(n12042), .A2(n12034), .ZN(n9528) );
  NAND2_X1 U8387 ( .A1(n14469), .A2(n6903), .ZN(n14327) );
  INV_X1 U8388 ( .A(n6903), .ZN(n12033) );
  NAND2_X1 U8389 ( .A1(n6905), .A2(n6904), .ZN(n11840) );
  AND2_X1 U8390 ( .A1(n8235), .A2(n8234), .ZN(n11771) );
  NAND2_X1 U8391 ( .A1(n11640), .A2(n9482), .ZN(n11772) );
  INV_X1 U8392 ( .A(n6905), .ZN(n11773) );
  NAND2_X1 U8393 ( .A1(n9519), .A2(n9518), .ZN(n11354) );
  NAND2_X1 U8394 ( .A1(n7349), .A2(n7348), .ZN(n11361) );
  AOI21_X1 U8395 ( .B1(n7350), .B2(n7352), .A(n6578), .ZN(n7348) );
  OR2_X1 U8396 ( .A1(n10658), .A2(n14002), .ZN(n11142) );
  NOR2_X1 U8397 ( .A1(n10831), .A2(n10837), .ZN(n10832) );
  NAND2_X1 U8398 ( .A1(n10832), .A2(n10668), .ZN(n10658) );
  AND2_X1 U8399 ( .A1(n9507), .A2(n8236), .ZN(n10828) );
  NAND2_X1 U8400 ( .A1(n10827), .A2(n10828), .ZN(n10826) );
  INV_X1 U8401 ( .A(n10828), .ZN(n10824) );
  CLKBUF_X1 U8402 ( .A(n10506), .Z(n10507) );
  NAND2_X1 U8403 ( .A1(n10172), .A2(n9469), .ZN(n10622) );
  AND2_X1 U8404 ( .A1(n14024), .A2(n12084), .ZN(n14351) );
  NAND2_X1 U8405 ( .A1(n7070), .A2(n6528), .ZN(n14168) );
  NAND2_X1 U8406 ( .A1(n7049), .A2(n7047), .ZN(n14290) );
  CLKBUF_X1 U8407 ( .A(n14834), .Z(n6691) );
  NAND2_X1 U8408 ( .A1(n9915), .A2(n9450), .ZN(n14843) );
  NAND2_X1 U8409 ( .A1(n14155), .A2(n10515), .ZN(n14848) );
  INV_X1 U8410 ( .A(n14843), .ZN(n14426) );
  NOR2_X1 U8411 ( .A1(n10594), .A2(n9554), .ZN(n9564) );
  INV_X1 U8412 ( .A(n14848), .ZN(n14431) );
  AND2_X1 U8413 ( .A1(n9265), .A2(n9658), .ZN(n9664) );
  XNOR2_X1 U8414 ( .A(n8190), .B(n8189), .ZN(n12626) );
  OAI21_X1 U8415 ( .B1(n8147), .B2(n8146), .A(n8145), .ZN(n8160) );
  AND2_X1 U8416 ( .A1(n7473), .A2(n7367), .ZN(n6763) );
  NAND2_X1 U8417 ( .A1(n8284), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7490) );
  XNOR2_X1 U8418 ( .A(n8147), .B(n8129), .ZN(n12047) );
  XNOR2_X1 U8419 ( .A(n8277), .B(n8276), .ZN(n9665) );
  INV_X1 U8420 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n8276) );
  NAND2_X1 U8421 ( .A1(n7111), .A2(n7112), .ZN(n7209) );
  NAND2_X1 U8422 ( .A1(n7320), .A2(n7901), .ZN(n7931) );
  NAND2_X1 U8423 ( .A1(n6859), .A2(n6858), .ZN(n7851) );
  NAND2_X1 U8424 ( .A1(n7836), .A2(n9877), .ZN(n6858) );
  NAND2_X1 U8425 ( .A1(n7285), .A2(n7819), .ZN(n7833) );
  NAND2_X1 U8426 ( .A1(n7794), .A2(n7815), .ZN(n7285) );
  XNOR2_X1 U8427 ( .A(n7794), .B(n7815), .ZN(n10167) );
  NAND2_X1 U8428 ( .A1(n7294), .A2(n7597), .ZN(n7293) );
  AND2_X1 U8429 ( .A1(n7579), .A2(n7580), .ZN(n9598) );
  OR2_X1 U8430 ( .A1(n7578), .A2(n7595), .ZN(n7579) );
  NAND2_X1 U8431 ( .A1(n7598), .A2(n7593), .ZN(n7578) );
  NAND2_X1 U8432 ( .A1(n6890), .A2(n7556), .ZN(n6889) );
  INV_X1 U8433 ( .A(n7558), .ZN(n6890) );
  OAI21_X1 U8434 ( .B1(n6838), .B2(n7523), .A(n7503), .ZN(n7507) );
  NAND2_X1 U8435 ( .A1(n7507), .A2(n7506), .ZN(n7554) );
  INV_X1 U8436 ( .A(n7117), .ZN(n14533) );
  NAND2_X1 U8437 ( .A1(n14539), .A2(n14540), .ZN(n14541) );
  XNOR2_X1 U8438 ( .A(n14548), .B(P1_ADDR_REG_5__SCAN_IN), .ZN(n14549) );
  NAND2_X1 U8439 ( .A1(n14560), .A2(n14559), .ZN(n14561) );
  NOR2_X1 U8440 ( .A1(n14506), .A2(n6672), .ZN(n14524) );
  AND2_X1 U8441 ( .A1(n14507), .A2(P1_ADDR_REG_10__SCAN_IN), .ZN(n6672) );
  AOI21_X1 U8442 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(n14509), .A(n14508), .ZN(
        n14521) );
  NOR2_X1 U8443 ( .A1(n14524), .A2(n14523), .ZN(n14508) );
  AOI21_X1 U8444 ( .B1(n12888), .B2(n10235), .A(n12291), .ZN(n12894) );
  INV_X1 U8445 ( .A(n12745), .ZN(n12017) );
  OAI21_X1 U8446 ( .B1(n12013), .B2(n6527), .A(n7185), .ZN(n12124) );
  NAND2_X1 U8447 ( .A1(n10559), .A2(n10558), .ZN(n10561) );
  AND3_X1 U8448 ( .A1(n12158), .A2(n12157), .A3(n12156), .ZN(n12648) );
  AND2_X1 U8449 ( .A1(n12630), .A2(n12275), .ZN(n12303) );
  AND4_X1 U8450 ( .A1(n11081), .A2(n11080), .A3(n11079), .A4(n11078), .ZN(
        n11371) );
  NAND2_X1 U8451 ( .A1(n12696), .A2(n12189), .ZN(n12654) );
  OAI21_X1 U8452 ( .B1(n11784), .B2(n7177), .A(n7174), .ZN(n11909) );
  NOR2_X1 U8453 ( .A1(n11786), .A2(n12747), .ZN(n7177) );
  AND2_X1 U8454 ( .A1(n7176), .A2(n7175), .ZN(n7174) );
  OR2_X1 U8455 ( .A1(n11783), .A2(n11785), .ZN(n7175) );
  OAI21_X1 U8456 ( .B1(n12685), .B2(n12237), .A(n12236), .ZN(n12662) );
  AND4_X1 U8457 ( .A1(n11950), .A2(n11949), .A3(n11948), .A4(n11947), .ZN(
        n12727) );
  NAND2_X1 U8458 ( .A1(n7170), .A2(n12133), .ZN(n12671) );
  INV_X1 U8459 ( .A(n12670), .ZN(n7170) );
  AND2_X1 U8460 ( .A1(n12678), .A2(n6637), .ZN(n7168) );
  NAND2_X1 U8461 ( .A1(n12671), .A2(n12136), .ZN(n12679) );
  AND4_X1 U8462 ( .A1(n11321), .A2(n11320), .A3(n11319), .A4(n11318), .ZN(
        n11542) );
  NAND2_X1 U8463 ( .A1(n11496), .A2(n11495), .ZN(n11499) );
  AND3_X1 U8464 ( .A1(n12172), .A2(n12171), .A3(n12170), .ZN(n13015) );
  INV_X1 U8465 ( .A(n12988), .ZN(n12846) );
  NAND2_X1 U8466 ( .A1(n12205), .A2(n12204), .ZN(n13082) );
  NAND2_X1 U8467 ( .A1(n6685), .A2(n7178), .ZN(n11904) );
  NAND2_X1 U8468 ( .A1(n7173), .A2(n11786), .ZN(n11905) );
  NAND2_X1 U8469 ( .A1(n6685), .A2(n11783), .ZN(n7173) );
  OR2_X1 U8470 ( .A1(n10542), .A2(n10541), .ZN(n12732) );
  OR2_X1 U8471 ( .A1(n11115), .A2(n11114), .ZN(n11264) );
  AND2_X1 U8472 ( .A1(n12274), .A2(n12273), .ZN(n12880) );
  INV_X1 U8473 ( .A(n7202), .ZN(n12718) );
  NAND2_X1 U8474 ( .A1(n10243), .A2(n11954), .ZN(n12739) );
  NAND2_X1 U8475 ( .A1(n7180), .A2(n7181), .ZN(n12730) );
  AND2_X1 U8476 ( .A1(n12331), .A2(n10793), .ZN(n12881) );
  INV_X1 U8477 ( .A(n12880), .ZN(n12910) );
  NAND2_X1 U8478 ( .A1(n12229), .A2(n12228), .ZN(n12954) );
  NAND2_X1 U8479 ( .A1(n10253), .A2(n10252), .ZN(n12967) );
  OR2_X1 U8480 ( .A1(n10225), .A2(n10231), .ZN(n12743) );
  INV_X1 U8481 ( .A(n12648), .ZN(n13029) );
  INV_X1 U8482 ( .A(n12727), .ZN(n13039) );
  INV_X1 U8483 ( .A(n11542), .ZN(n12748) );
  INV_X1 U8484 ( .A(n11502), .ZN(n12749) );
  INV_X1 U8485 ( .A(n11371), .ZN(n12750) );
  INV_X1 U8486 ( .A(n11128), .ZN(n12752) );
  INV_X1 U8487 ( .A(P3_ADDR_REG_0__SCAN_IN), .ZN(n15109) );
  INV_X1 U8488 ( .A(n6981), .ZN(n10419) );
  INV_X1 U8489 ( .A(P3_ADDR_REG_4__SCAN_IN), .ZN(n15125) );
  NAND2_X1 U8490 ( .A1(n6989), .A2(n6990), .ZN(n15110) );
  INV_X1 U8491 ( .A(P3_ADDR_REG_5__SCAN_IN), .ZN(n15145) );
  INV_X1 U8492 ( .A(n7068), .ZN(n15134) );
  NOR2_X1 U8493 ( .A1(n6652), .A2(n8526), .ZN(n10399) );
  INV_X1 U8494 ( .A(P3_ADDR_REG_7__SCAN_IN), .ZN(n15169) );
  NAND2_X1 U8495 ( .A1(n6882), .A2(n8476), .ZN(n15157) );
  INV_X1 U8496 ( .A(n7057), .ZN(n10534) );
  NOR2_X1 U8497 ( .A1(n11326), .A2(n10849), .ZN(n10848) );
  XNOR2_X1 U8498 ( .A(n8341), .B(n8340), .ZN(n11516) );
  NOR2_X1 U8499 ( .A1(n11425), .A2(n8538), .ZN(n11510) );
  XNOR2_X1 U8500 ( .A(n8541), .B(n8540), .ZN(n12757) );
  NOR2_X1 U8501 ( .A1(n12757), .A2(n12758), .ZN(n12756) );
  AND2_X1 U8502 ( .A1(n6957), .A2(n6956), .ZN(n12773) );
  INV_X1 U8503 ( .A(n12774), .ZN(n6956) );
  INV_X1 U8504 ( .A(n6957), .ZN(n12775) );
  INV_X1 U8505 ( .A(n15097), .ZN(n15168) );
  OAI21_X1 U8506 ( .B1(n14645), .B2(n14641), .A(n14642), .ZN(n12798) );
  NOR2_X1 U8507 ( .A1(n12798), .A2(n12799), .ZN(n12797) );
  INV_X1 U8508 ( .A(n15155), .ZN(n15131) );
  NOR2_X1 U8509 ( .A1(n8424), .A2(n7192), .ZN(n8454) );
  NOR2_X1 U8510 ( .A1(n12806), .A2(n12807), .ZN(n12805) );
  AND2_X1 U8511 ( .A1(n12252), .A2(n12251), .ZN(n12918) );
  NAND2_X1 U8512 ( .A1(n7021), .A2(n12480), .ZN(n12912) );
  NAND2_X1 U8513 ( .A1(n12928), .A2(n12927), .ZN(n7021) );
  AOI21_X1 U8514 ( .B1(n12623), .B2(n12311), .A(n12220), .ZN(n12946) );
  AND2_X1 U8515 ( .A1(n12232), .A2(n12231), .ZN(n12960) );
  NAND2_X1 U8516 ( .A1(n12990), .A2(n12354), .ZN(n12979) );
  NAND2_X1 U8517 ( .A1(n7323), .A2(n12845), .ZN(n12976) );
  OAI21_X1 U8518 ( .B1(n12166), .B2(n12165), .A(n12164), .ZN(n13097) );
  NAND2_X1 U8519 ( .A1(n7030), .A2(n12358), .ZN(n13019) );
  NAND2_X1 U8520 ( .A1(n11989), .A2(n11988), .ZN(n12304) );
  NAND2_X1 U8521 ( .A1(n11714), .A2(n12428), .ZN(n11939) );
  AND2_X1 U8522 ( .A1(n11700), .A2(n11699), .ZN(n11705) );
  INV_X1 U8523 ( .A(n12877), .ZN(n13050) );
  NAND2_X1 U8524 ( .A1(n7344), .A2(n6497), .ZN(n11540) );
  INV_X1 U8525 ( .A(n15208), .ZN(n11954) );
  NAND2_X1 U8526 ( .A1(n10995), .A2(n12512), .ZN(n11018) );
  NAND2_X1 U8527 ( .A1(n15170), .A2(n12378), .ZN(n10995) );
  NAND2_X1 U8528 ( .A1(n10485), .A2(n11954), .ZN(n15211) );
  AND2_X2 U8529 ( .A1(n10242), .A2(n15206), .ZN(n15208) );
  AND2_X2 U8530 ( .A1(n10498), .A2(n10497), .ZN(n15281) );
  AND2_X1 U8531 ( .A1(n14659), .A2(n14661), .ZN(n14685) );
  INV_X1 U8532 ( .A(n6765), .ZN(n6764) );
  OAI21_X1 U8533 ( .B1(n13056), .B2(n14680), .A(n7023), .ZN(n6765) );
  NAND2_X1 U8534 ( .A1(n13065), .A2(n13064), .ZN(n13303) );
  INV_X2 U8535 ( .A(n15268), .ZN(n15266) );
  AND2_X1 U8536 ( .A1(n10198), .A2(n10197), .ZN(n13317) );
  AND2_X1 U8537 ( .A1(n8509), .A2(P3_STATE_REG_SCAN_IN), .ZN(n13318) );
  XNOR2_X1 U8538 ( .A(n7158), .B(n12319), .ZN(n13321) );
  AOI21_X1 U8539 ( .B1(n12316), .B2(n12317), .A(n7159), .ZN(n7158) );
  NOR2_X1 U8540 ( .A1(n13866), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n7159) );
  XNOR2_X1 U8541 ( .A(n12091), .B(n12317), .ZN(n12333) );
  INV_X1 U8542 ( .A(SI_26_), .ZN(n11877) );
  XNOR2_X1 U8543 ( .A(n10217), .B(n10216), .ZN(n10779) );
  INV_X1 U8544 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n10216) );
  INV_X1 U8545 ( .A(SI_19_), .ZN(n12163) );
  INV_X1 U8546 ( .A(SI_16_), .ZN(n10152) );
  INV_X1 U8547 ( .A(n7155), .ZN(n10324) );
  NAND2_X1 U8548 ( .A1(n7146), .A2(n9875), .ZN(n9939) );
  INV_X1 U8549 ( .A(SI_13_), .ZN(n11702) );
  NOR2_X1 U8550 ( .A1(n10187), .A2(P3_STATE_REG_SCAN_IN), .ZN(n13320) );
  NAND2_X1 U8551 ( .A1(n9643), .A2(n9642), .ZN(n9661) );
  OAI21_X1 U8552 ( .B1(n9586), .B2(n6498), .A(n7129), .ZN(n9621) );
  NAND2_X1 U8553 ( .A1(n7132), .A2(n9588), .ZN(n9617) );
  NAND2_X1 U8554 ( .A1(n9586), .A2(n7133), .ZN(n7132) );
  NAND2_X1 U8555 ( .A1(n9586), .A2(n9585), .ZN(n9608) );
  NOR2_X1 U8556 ( .A1(n13335), .A2(n9594), .ZN(n6961) );
  INV_X1 U8557 ( .A(n7264), .ZN(n10631) );
  OAI21_X1 U8558 ( .B1(n10388), .B2(n7265), .A(n7268), .ZN(n7264) );
  INV_X1 U8559 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n11671) );
  NAND2_X1 U8560 ( .A1(n7280), .A2(n7281), .ZN(n13349) );
  NOR2_X1 U8561 ( .A1(n13407), .A2(n12572), .ZN(n13351) );
  INV_X1 U8562 ( .A(n12614), .ZN(n7252) );
  AOI21_X1 U8563 ( .B1(n13336), .B2(n7254), .A(n6546), .ZN(n7253) );
  NAND2_X1 U8564 ( .A1(n10628), .A2(n7267), .ZN(n7266) );
  AND2_X1 U8565 ( .A1(n10003), .A2(n10005), .ZN(n10032) );
  NAND2_X1 U8566 ( .A1(n10032), .A2(n10031), .ZN(n10030) );
  OAI21_X1 U8567 ( .B1(n12577), .B2(n7236), .A(n7234), .ZN(n13359) );
  NAND2_X1 U8568 ( .A1(n7250), .A2(n7248), .ZN(n11997) );
  AND2_X1 U8569 ( .A1(n7250), .A2(n6553), .ZN(n11863) );
  NAND2_X1 U8570 ( .A1(n6711), .A2(n11860), .ZN(n7250) );
  NAND2_X1 U8571 ( .A1(n7242), .A2(n7246), .ZN(n11998) );
  OR2_X1 U8572 ( .A1(n6711), .A2(n7249), .ZN(n7242) );
  NAND2_X1 U8573 ( .A1(n7238), .A2(n7239), .ZN(n13377) );
  INV_X1 U8574 ( .A(n12577), .ZN(n13389) );
  NOR2_X1 U8575 ( .A1(n10388), .A2(n10387), .ZN(n10585) );
  INV_X1 U8576 ( .A(n13372), .ZN(n13422) );
  INV_X1 U8577 ( .A(n13415), .ZN(n13426) );
  NAND2_X1 U8578 ( .A1(n9989), .A2(n9988), .ZN(n13428) );
  NOR4_X2 U8579 ( .A1(n9222), .A2(n9221), .A3(n13588), .A4(n9220), .ZN(n9223)
         );
  NOR2_X1 U8580 ( .A1(n7445), .A2(n9195), .ZN(n9196) );
  OR2_X1 U8581 ( .A1(n13609), .A2(n9147), .ZN(n9136) );
  NAND2_X1 U8582 ( .A1(n9105), .A2(n9104), .ZN(n13432) );
  NAND2_X1 U8583 ( .A1(n9086), .A2(n9085), .ZN(n13552) );
  OR2_X1 U8584 ( .A1(n13645), .A2(n9147), .ZN(n9086) );
  AND2_X1 U8585 ( .A1(n8651), .A2(n8650), .ZN(n6660) );
  INV_X1 U8586 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n7496) );
  NAND2_X1 U8587 ( .A1(n13523), .A2(n10086), .ZN(n13756) );
  INV_X1 U8588 ( .A(n13521), .ZN(n13759) );
  AOI21_X1 U8589 ( .B1(n13601), .B2(n13602), .A(n13600), .ZN(n13773) );
  NAND2_X1 U8590 ( .A1(n7399), .A2(n13557), .ZN(n13616) );
  NAND2_X1 U8591 ( .A1(n7399), .A2(n7397), .ZN(n13776) );
  NAND2_X1 U8592 ( .A1(n13654), .A2(n13551), .ZN(n13639) );
  NOR2_X1 U8593 ( .A1(n13713), .A2(n13577), .ZN(n13707) );
  INV_X1 U8594 ( .A(n13822), .ZN(n13722) );
  NAND2_X1 U8595 ( .A1(n13741), .A2(n13537), .ZN(n13725) );
  INV_X1 U8596 ( .A(n7406), .ZN(n11963) );
  NAND2_X1 U8597 ( .A1(n8896), .A2(n8895), .ZN(n11802) );
  NAND2_X1 U8598 ( .A1(n6912), .A2(n6913), .ZN(n11555) );
  NAND2_X1 U8599 ( .A1(n11246), .A2(n11245), .ZN(n6917) );
  NAND2_X1 U8600 ( .A1(n7391), .A2(n7394), .ZN(n14718) );
  NAND2_X1 U8601 ( .A1(n7392), .A2(n6520), .ZN(n11251) );
  NAND2_X1 U8602 ( .A1(n6923), .A2(n10367), .ZN(n10711) );
  NAND2_X1 U8603 ( .A1(n10568), .A2(n10569), .ZN(n6923) );
  AND2_X1 U8604 ( .A1(n15002), .A2(n13516), .ZN(n14722) );
  INV_X1 U8605 ( .A(n14722), .ZN(n14983) );
  AND2_X1 U8606 ( .A1(n8610), .A2(n10368), .ZN(n14992) );
  AND2_X1 U8607 ( .A1(n9983), .A2(n9567), .ZN(n15016) );
  INV_X1 U8608 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n8565) );
  NAND2_X1 U8609 ( .A1(n6734), .A2(n8783), .ZN(n6732) );
  NAND2_X1 U8610 ( .A1(n8607), .A2(n6731), .ZN(n6733) );
  NOR2_X1 U8611 ( .A1(n8783), .A2(n6734), .ZN(n6731) );
  INV_X1 U8612 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n13871) );
  NAND2_X2 U8613 ( .A1(n8599), .A2(n8598), .ZN(n13526) );
  NAND3_X1 U8614 ( .A1(n9242), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_IR_REG_27__SCAN_IN), .ZN(n8598) );
  NAND2_X1 U8615 ( .A1(n9245), .A2(n9244), .ZN(n12011) );
  INV_X1 U8616 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n11619) );
  INV_X1 U8618 ( .A(n10368), .ZN(n13516) );
  INV_X1 U8619 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n13208) );
  INV_X1 U8620 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n10783) );
  INV_X1 U8621 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n10524) );
  INV_X1 U8622 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n9936) );
  INV_X1 U8623 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n9651) );
  INV_X1 U8624 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n9646) );
  INV_X1 U8625 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n9632) );
  NAND2_X1 U8626 ( .A1(n6817), .A2(n6815), .ZN(n11194) );
  NAND2_X1 U8627 ( .A1(n7091), .A2(n7095), .ZN(n13875) );
  NAND2_X1 U8628 ( .A1(n13952), .A2(n7096), .ZN(n7091) );
  NAND2_X1 U8629 ( .A1(n12021), .A2(n9351), .ZN(n13885) );
  NAND2_X1 U8630 ( .A1(n9324), .A2(n6829), .ZN(n6826) );
  CLKBUF_X1 U8631 ( .A(n9282), .Z(n10510) );
  NAND2_X1 U8632 ( .A1(n6594), .A2(n7088), .ZN(n7087) );
  NAND2_X1 U8633 ( .A1(n6811), .A2(n9314), .ZN(n11464) );
  NAND2_X1 U8634 ( .A1(n6817), .A2(n6812), .ZN(n6811) );
  NAND2_X1 U8635 ( .A1(n11820), .A2(n7099), .ZN(n11895) );
  NOR2_X1 U8636 ( .A1(n11893), .A2(n7100), .ZN(n7099) );
  INV_X1 U8637 ( .A(n9335), .ZN(n7100) );
  NAND2_X1 U8638 ( .A1(n11820), .A2(n9335), .ZN(n11894) );
  NAND2_X1 U8639 ( .A1(n9361), .A2(n14007), .ZN(n13933) );
  NAND2_X1 U8640 ( .A1(n7079), .A2(n6798), .ZN(n13942) );
  NAND2_X1 U8641 ( .A1(n6799), .A2(n13932), .ZN(n6798) );
  INV_X1 U8642 ( .A(n9361), .ZN(n6799) );
  XNOR2_X1 U8643 ( .A(n9324), .B(n9325), .ZN(n11763) );
  INV_X1 U8644 ( .A(n11736), .ZN(n12031) );
  NAND2_X1 U8645 ( .A1(n13911), .A2(n9399), .ZN(n13972) );
  NAND2_X1 U8646 ( .A1(n6819), .A2(n6823), .ZN(n11821) );
  NAND2_X1 U8647 ( .A1(n9324), .A2(n6824), .ZN(n6819) );
  AND2_X1 U8648 ( .A1(n13999), .A2(n14319), .ZN(n14011) );
  AND2_X1 U8649 ( .A1(n9463), .A2(n10593), .ZN(n13999) );
  NAND2_X1 U8650 ( .A1(n6818), .A2(n7102), .ZN(n13994) );
  AND2_X1 U8651 ( .A1(n6807), .A2(n7101), .ZN(n6818) );
  AND2_X1 U8652 ( .A1(n9664), .A2(n9460), .ZN(n10593) );
  AND2_X1 U8653 ( .A1(n9666), .A2(n9747), .ZN(n14319) );
  AND3_X1 U8654 ( .A1(n6716), .A2(n6715), .A3(n6600), .ZN(n8273) );
  OAI21_X1 U8655 ( .B1(n13975), .B2(n8119), .A(n8016), .ZN(n14027) );
  OAI211_X1 U8656 ( .C1(n13947), .C2(n8119), .A(n7897), .B(n7896), .ZN(n14320)
         );
  INV_X1 U8657 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n12114) );
  OR2_X1 U8658 ( .A1(n12083), .A2(n14119), .ZN(n14128) );
  NAND2_X1 U8659 ( .A1(n14138), .A2(n13878), .ZN(n9542) );
  AOI21_X1 U8660 ( .B1(n7361), .B2(n14150), .A(n7363), .ZN(n7359) );
  AND2_X1 U8661 ( .A1(n14143), .A2(n7361), .ZN(n14133) );
  INV_X1 U8662 ( .A(n6769), .ZN(n6714) );
  AOI21_X1 U8663 ( .B1(n14131), .B2(n14321), .A(n6770), .ZN(n6769) );
  INV_X1 U8664 ( .A(n6794), .ZN(n6793) );
  NAND2_X1 U8665 ( .A1(n14215), .A2(n9540), .ZN(n14187) );
  NAND2_X1 U8666 ( .A1(n8063), .A2(n8062), .ZN(n14377) );
  AND2_X1 U8667 ( .A1(n14218), .A2(n14217), .ZN(n14384) );
  NAND2_X1 U8668 ( .A1(n7353), .A2(n6524), .ZN(n14267) );
  NAND2_X1 U8669 ( .A1(n11837), .A2(n9484), .ZN(n12043) );
  AND2_X1 U8670 ( .A1(n11598), .A2(n9480), .ZN(n11641) );
  CLKBUF_X1 U8671 ( .A(n11648), .Z(n11650) );
  CLKBUF_X1 U8672 ( .A(n11601), .Z(n11603) );
  OAI21_X1 U8673 ( .B1(n11414), .B2(n6776), .A(n6774), .ZN(n11476) );
  NAND2_X1 U8674 ( .A1(n11412), .A2(n9479), .ZN(n11478) );
  NAND2_X1 U8675 ( .A1(n11233), .A2(n11345), .ZN(n11351) );
  NAND2_X1 U8676 ( .A1(n11230), .A2(n9477), .ZN(n11157) );
  NAND2_X1 U8677 ( .A1(n7347), .A2(n7350), .ZN(n11156) );
  OR2_X1 U8678 ( .A1(n11232), .A2(n7352), .ZN(n7347) );
  INV_X1 U8679 ( .A(n14346), .ZN(n14823) );
  CLKBUF_X1 U8680 ( .A(n9289), .Z(n10605) );
  NAND2_X1 U8681 ( .A1(n10602), .A2(n12108), .ZN(n14243) );
  NOR2_X2 U8682 ( .A1(n14830), .A2(n10619), .ZN(n14277) );
  NOR2_X2 U8683 ( .A1(n14830), .A2(n10601), .ZN(n14346) );
  INV_X1 U8684 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n6901) );
  NAND2_X1 U8685 ( .A1(n14363), .A2(n14209), .ZN(n6795) );
  INV_X1 U8686 ( .A(n14423), .ZN(n14375) );
  INV_X1 U8687 ( .A(n14118), .ZN(n14437) );
  NAND2_X1 U8688 ( .A1(n14128), .A2(n14120), .ZN(n14439) );
  NAND2_X1 U8689 ( .A1(n9932), .A2(n8212), .ZN(n7773) );
  INV_X1 U8690 ( .A(n9289), .ZN(n10518) );
  NAND2_X1 U8691 ( .A1(n9653), .A2(n9664), .ZN(n14831) );
  AND2_X1 U8692 ( .A1(n10187), .A2(P1_U3086), .ZN(n14473) );
  MUX2_X1 U8693 ( .A(P1_IR_REG_31__SCAN_IN), .B(n7474), .S(
        P1_IR_REG_29__SCAN_IN), .Z(n7476) );
  XNOR2_X1 U8694 ( .A(n8160), .B(n8159), .ZN(n12121) );
  CLKBUF_X1 U8695 ( .A(n8290), .Z(n8291) );
  NAND2_X1 U8696 ( .A1(n6834), .A2(n6833), .ZN(n8285) );
  NAND2_X1 U8697 ( .A1(n7535), .A2(n6530), .ZN(n8287) );
  XNOR2_X1 U8698 ( .A(n8041), .B(n8040), .ZN(n11888) );
  XNOR2_X1 U8699 ( .A(n8023), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n14482) );
  INV_X1 U8700 ( .A(n9915), .ZN(n14483) );
  INV_X1 U8701 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n11123) );
  INV_X1 U8702 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n10976) );
  INV_X1 U8703 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n10781) );
  INV_X1 U8704 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n9778) );
  NAND2_X1 U8705 ( .A1(n7723), .A2(n7722), .ZN(n7743) );
  NAND2_X1 U8706 ( .A1(n7719), .A2(n7718), .ZN(n7723) );
  OAI21_X1 U8707 ( .B1(n7507), .B2(n7506), .A(n7554), .ZN(n9628) );
  XNOR2_X1 U8708 ( .A(n14541), .B(n6766), .ZN(n14595) );
  INV_X1 U8709 ( .A(n14542), .ZN(n6766) );
  INV_X1 U8710 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n7120) );
  INV_X1 U8711 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n7123) );
  INV_X1 U8712 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n7121) );
  XNOR2_X1 U8713 ( .A(n14561), .B(n14562), .ZN(n14598) );
  NAND2_X1 U8714 ( .A1(n7124), .A2(n14567), .ZN(n14602) );
  NAND2_X1 U8715 ( .A1(n14599), .A2(P2_ADDR_REG_9__SCAN_IN), .ZN(n7124) );
  NAND2_X1 U8716 ( .A1(n6659), .A2(n6870), .ZN(n14775) );
  NAND2_X1 U8717 ( .A1(n6871), .A2(n14574), .ZN(n6870) );
  INV_X1 U8718 ( .A(n6872), .ZN(n6871) );
  NOR2_X1 U8719 ( .A1(n14574), .A2(n14575), .ZN(n14776) );
  XNOR2_X1 U8720 ( .A(n7119), .B(n7118), .ZN(n14606) );
  OR2_X1 U8721 ( .A1(n12548), .A2(n12547), .ZN(n6673) );
  NAND2_X1 U8722 ( .A1(n10166), .A2(n6648), .ZN(P3_U3183) );
  NAND2_X1 U8723 ( .A1(n6983), .A2(n6984), .ZN(n10397) );
  INV_X1 U8724 ( .A(n6880), .ZN(n11444) );
  NAND2_X1 U8725 ( .A1(n8556), .A2(n15163), .ZN(n6965) );
  OAI21_X1 U8726 ( .B1(n13333), .B2(n9593), .A(n6959), .ZN(P3_U3294) );
  NOR2_X1 U8727 ( .A1(n6961), .A2(n6960), .ZN(n6959) );
  INV_X1 U8728 ( .A(n9567), .ZN(n9568) );
  INV_X1 U8729 ( .A(n6689), .ZN(n6688) );
  OAI21_X1 U8730 ( .B1(n6944), .B2(n13415), .A(n13342), .ZN(n6689) );
  NAND2_X1 U8731 ( .A1(n15094), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n6937) );
  NAND2_X1 U8732 ( .A1(n13849), .A2(n15096), .ZN(n6938) );
  NAND2_X1 U8733 ( .A1(n6699), .A2(n6698), .ZN(P2_U3493) );
  OR2_X1 U8734 ( .A1(n15066), .A2(n9102), .ZN(n6698) );
  OAI211_X1 U8735 ( .C1(n6804), .C2(n6801), .A(n6800), .B(n9468), .ZN(P1_U3240) );
  NAND2_X1 U8736 ( .A1(n6802), .A2(n9432), .ZN(n6801) );
  NAND2_X1 U8737 ( .A1(n6804), .A2(n6508), .ZN(n6800) );
  NAND2_X1 U8738 ( .A1(n6902), .A2(n6899), .ZN(P1_U3558) );
  AOI21_X1 U8739 ( .B1(n14438), .B2(n14375), .A(n6900), .ZN(n6899) );
  NAND2_X1 U8740 ( .A1(n14439), .A2(n14856), .ZN(n6902) );
  NOR2_X1 U8741 ( .A1(n14856), .A2(n6901), .ZN(n6900) );
  OAI21_X1 U8742 ( .B1(n14445), .B2(n14854), .A(n6696), .ZN(P1_U3555) );
  INV_X1 U8743 ( .A(n6697), .ZN(n6696) );
  AND2_X1 U8744 ( .A1(n6788), .A2(n6795), .ZN(n14445) );
  OAI22_X1 U8745 ( .A1(n9496), .A2(n14423), .B1(n14856), .B2(n14364), .ZN(
        n6697) );
  NAND2_X1 U8746 ( .A1(n14363), .A2(n6785), .ZN(n6787) );
  AOI21_X1 U8747 ( .B1(n6794), .B2(n14849), .A(n6789), .ZN(n6784) );
  NAND2_X1 U8748 ( .A1(n6790), .A2(n14849), .ZN(n6783) );
  NAND2_X1 U8749 ( .A1(n6629), .A2(n6739), .ZN(n14772) );
  INV_X2 U8750 ( .A(n10389), .ZN(n9992) );
  INV_X1 U8751 ( .A(n9275), .ZN(n9288) );
  NAND2_X2 U8752 ( .A1(n8967), .A2(n8966), .ZN(n13734) );
  NAND2_X1 U8753 ( .A1(n12094), .A2(n9926), .ZN(n12290) );
  INV_X1 U8754 ( .A(n8215), .ZN(n8216) );
  AND2_X1 U8755 ( .A1(n9265), .A2(n9264), .ZN(n12065) );
  INV_X1 U8756 ( .A(n12065), .ZN(n9287) );
  AND2_X1 U8757 ( .A1(n6521), .A2(n11525), .ZN(n6497) );
  OR2_X1 U8758 ( .A1(n9616), .A2(n7131), .ZN(n6498) );
  AND2_X1 U8759 ( .A1(n7027), .A2(n12457), .ZN(n6500) );
  OR2_X1 U8760 ( .A1(n14586), .A2(n14585), .ZN(n6501) );
  INV_X1 U8761 ( .A(n9543), .ZN(n6669) );
  NOR2_X1 U8762 ( .A1(n14404), .A2(n14264), .ZN(n6502) );
  NAND2_X1 U8763 ( .A1(n14487), .A2(P3_ADDR_REG_1__SCAN_IN), .ZN(n6503) );
  AND2_X1 U8764 ( .A1(n13817), .A2(n13578), .ZN(n6504) );
  AND2_X1 U8765 ( .A1(n11273), .A2(n11274), .ZN(n6505) );
  OR2_X1 U8766 ( .A1(n14582), .A2(n14581), .ZN(n6506) );
  AND2_X1 U8767 ( .A1(n7402), .A2(n13543), .ZN(n6507) );
  AND2_X1 U8768 ( .A1(n6596), .A2(n6802), .ZN(n6508) );
  AND2_X1 U8769 ( .A1(n7208), .A2(n12923), .ZN(n6509) );
  NOR2_X1 U8770 ( .A1(n12584), .A2(n12583), .ZN(n6510) );
  OR2_X1 U8771 ( .A1(n6827), .A2(n6643), .ZN(n6511) );
  AND2_X1 U8772 ( .A1(n7148), .A2(n9662), .ZN(n6512) );
  INV_X1 U8773 ( .A(n13408), .ZN(n7282) );
  AND2_X1 U8774 ( .A1(n7181), .A2(n6632), .ZN(n6513) );
  AND2_X1 U8775 ( .A1(n7337), .A2(n11214), .ZN(n6514) );
  INV_X1 U8776 ( .A(n11964), .ZN(n6949) );
  INV_X1 U8777 ( .A(n14768), .ZN(n6739) );
  OAI22_X1 U8778 ( .A1(n9496), .A2(n14468), .B1(n14849), .B2(n14446), .ZN(
        n6789) );
  INV_X1 U8779 ( .A(n6951), .ZN(n14706) );
  NAND2_X1 U8780 ( .A1(n7798), .A2(n7797), .ZN(n11488) );
  INV_X1 U8781 ( .A(n11488), .ZN(n6891) );
  NAND2_X1 U8782 ( .A1(n11233), .A2(n6893), .ZN(n6894) );
  OR2_X1 U8783 ( .A1(n14849), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n6515) );
  OR2_X1 U8784 ( .A1(n14856), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n6516) );
  INV_X4 U8785 ( .A(n10791), .ZN(n10454) );
  AND2_X1 U8786 ( .A1(n13671), .A2(n13548), .ZN(n6517) );
  NAND2_X1 U8787 ( .A1(n9309), .A2(n9308), .ZN(n6518) );
  INV_X1 U8788 ( .A(n14090), .ZN(n6752) );
  OR2_X1 U8789 ( .A1(n7533), .A2(n7113), .ZN(n6519) );
  OR2_X1 U8790 ( .A1(n10968), .A2(n10955), .ZN(n6520) );
  INV_X1 U8791 ( .A(n8683), .ZN(n8765) );
  NAND2_X1 U8792 ( .A1(n12412), .A2(n15254), .ZN(n6521) );
  OAI211_X2 U8793 ( .C1(n7749), .C2(n9631), .A(n7529), .B(n7528), .ZN(n14345)
         );
  NAND2_X1 U8794 ( .A1(n12265), .A2(n12264), .ZN(n13062) );
  NOR2_X1 U8795 ( .A1(n8493), .A2(n12802), .ZN(n6522) );
  NAND2_X1 U8796 ( .A1(n13386), .A2(n13387), .ZN(n13358) );
  AND2_X1 U8797 ( .A1(n7312), .A2(n13665), .ZN(n6523) );
  NAND2_X1 U8798 ( .A1(n14404), .A2(n14028), .ZN(n6524) );
  AND2_X1 U8799 ( .A1(n8734), .A2(n8733), .ZN(n6525) );
  AND2_X1 U8800 ( .A1(n8995), .A2(n8994), .ZN(n6526) );
  AND2_X1 U8801 ( .A1(n12012), .A2(n12017), .ZN(n6527) );
  OR2_X1 U8802 ( .A1(n14171), .A2(n14170), .ZN(n6528) );
  AND2_X1 U8803 ( .A1(n7513), .A2(n7043), .ZN(n6529) );
  NAND2_X1 U8804 ( .A1(n9447), .A2(n8289), .ZN(n9265) );
  AND2_X1 U8805 ( .A1(n8282), .A2(n8283), .ZN(n6530) );
  OR2_X1 U8806 ( .A1(n7945), .A2(n7944), .ZN(n6531) );
  OR2_X1 U8807 ( .A1(n9646), .A2(P2_DATAO_REG_8__SCAN_IN), .ZN(n6532) );
  NOR2_X1 U8808 ( .A1(n13769), .A2(n13592), .ZN(n6533) );
  AND2_X1 U8809 ( .A1(n6518), .A2(n7101), .ZN(n6534) );
  INV_X1 U8810 ( .A(n12837), .ZN(n12441) );
  NAND2_X1 U8811 ( .A1(n7291), .A2(n7293), .ZN(n7633) );
  INV_X1 U8812 ( .A(n7410), .ZN(n7405) );
  NAND2_X1 U8813 ( .A1(n8803), .A2(n8802), .ZN(n11059) );
  AND2_X1 U8814 ( .A1(n7309), .A2(n7308), .ZN(n6535) );
  AND2_X1 U8815 ( .A1(n8456), .A2(n12820), .ZN(n6536) );
  OR2_X1 U8816 ( .A1(n9303), .A2(n10895), .ZN(n6537) );
  NAND2_X1 U8817 ( .A1(n7907), .A2(n7906), .ZN(n13949) );
  AOI21_X1 U8818 ( .B1(n12333), .B2(n10449), .A(n7451), .ZN(n14662) );
  INV_X1 U8819 ( .A(n12993), .ZN(n7027) );
  NAND2_X1 U8820 ( .A1(n12577), .A2(n12576), .ZN(n13386) );
  NAND2_X1 U8821 ( .A1(n13367), .A2(n12600), .ZN(n13416) );
  NOR2_X1 U8822 ( .A1(n8458), .A2(n7340), .ZN(n8313) );
  AND2_X1 U8823 ( .A1(n13949), .A2(n14320), .ZN(n6538) );
  AND3_X1 U8824 ( .A1(n7114), .A2(n8283), .A3(n7472), .ZN(n6539) );
  NAND2_X1 U8825 ( .A1(n14193), .A2(n14192), .ZN(n14191) );
  OR2_X1 U8826 ( .A1(n14562), .A2(n14561), .ZN(n6540) );
  INV_X1 U8827 ( .A(n8045), .ZN(n7229) );
  INV_X1 U8828 ( .A(n7249), .ZN(n7248) );
  INV_X1 U8829 ( .A(n13949), .ZN(n14469) );
  OR2_X1 U8830 ( .A1(n11802), .A2(n11796), .ZN(n6541) );
  INV_X1 U8831 ( .A(n13932), .ZN(n7081) );
  INV_X1 U8832 ( .A(n9303), .ZN(n7106) );
  NOR2_X1 U8833 ( .A1(n13903), .A2(n9388), .ZN(n6542) );
  AND3_X1 U8834 ( .A1(n8282), .A2(n6539), .A3(n6499), .ZN(n6543) );
  AND2_X1 U8835 ( .A1(n8324), .A2(n8463), .ZN(n6544) );
  NOR2_X1 U8836 ( .A1(n14625), .A2(n8491), .ZN(n6545) );
  AND2_X1 U8837 ( .A1(n7255), .A2(n12614), .ZN(n6546) );
  INV_X1 U8838 ( .A(n7203), .ZN(n7201) );
  NOR2_X1 U8839 ( .A1(n6554), .A2(n12719), .ZN(n7203) );
  AND2_X1 U8840 ( .A1(n13773), .A2(n13772), .ZN(n6547) );
  NOR2_X1 U8841 ( .A1(n13949), .A2(n14320), .ZN(n6548) );
  AND2_X1 U8842 ( .A1(n9052), .A2(n9051), .ZN(n6549) );
  AND3_X1 U8843 ( .A1(n7163), .A2(n12543), .A3(n7162), .ZN(n6550) );
  AND2_X1 U8844 ( .A1(n8960), .A2(n8959), .ZN(n6551) );
  OR2_X1 U8845 ( .A1(n11392), .A2(n6958), .ZN(n6552) );
  NAND2_X1 U8846 ( .A1(n11859), .A2(n11858), .ZN(n6553) );
  AND2_X1 U8847 ( .A1(n7206), .A2(n7204), .ZN(n6554) );
  AND2_X1 U8848 ( .A1(n11715), .A2(n11699), .ZN(n6555) );
  OR2_X1 U8849 ( .A1(n14743), .A2(n11556), .ZN(n6556) );
  INV_X1 U8850 ( .A(n12857), .ZN(n7330) );
  NOR2_X1 U8851 ( .A1(n13791), .A2(n13552), .ZN(n6557) );
  NOR2_X1 U8852 ( .A1(n8944), .A2(n8943), .ZN(n6558) );
  OR2_X1 U8853 ( .A1(n13722), .A2(n13540), .ZN(n6559) );
  AND2_X1 U8854 ( .A1(n9356), .A2(n9358), .ZN(n6560) );
  AND2_X1 U8855 ( .A1(n13544), .A2(n13543), .ZN(n6561) );
  AND2_X1 U8856 ( .A1(n13688), .A2(n13546), .ZN(n6562) );
  AND2_X1 U8857 ( .A1(n14750), .A2(n11252), .ZN(n6563) );
  AND2_X1 U8858 ( .A1(n7309), .A2(n7310), .ZN(n6564) );
  NAND2_X1 U8859 ( .A1(n12051), .A2(n12052), .ZN(n6565) );
  OR2_X1 U8860 ( .A1(n14451), .A2(n14213), .ZN(n6566) );
  AND2_X1 U8861 ( .A1(n9353), .A2(n9351), .ZN(n6567) );
  AND2_X1 U8862 ( .A1(n11497), .A2(n11495), .ZN(n6568) );
  AND2_X1 U8863 ( .A1(n13791), .A2(n13552), .ZN(n6569) );
  OR2_X1 U8864 ( .A1(n8135), .A2(n8134), .ZN(n6570) );
  AND2_X1 U8865 ( .A1(n6896), .A2(n14356), .ZN(n6571) );
  AND2_X1 U8866 ( .A1(n9490), .A2(n6524), .ZN(n6572) );
  INV_X1 U8867 ( .A(n7454), .ZN(n7098) );
  NOR2_X1 U8868 ( .A1(n12056), .A2(n12055), .ZN(n7454) );
  AND2_X1 U8869 ( .A1(n12367), .A2(n10481), .ZN(n12541) );
  AND2_X1 U8870 ( .A1(n14716), .A2(n13438), .ZN(n6573) );
  NAND2_X1 U8871 ( .A1(n8131), .A2(n8130), .ZN(n14158) );
  NOR2_X1 U8872 ( .A1(n11488), .A2(n14033), .ZN(n6574) );
  NAND2_X1 U8873 ( .A1(n12064), .A2(n12063), .ZN(n6575) );
  NOR2_X1 U8874 ( .A1(n10709), .A2(n10708), .ZN(n6576) );
  NOR2_X1 U8875 ( .A1(n11571), .A2(n11352), .ZN(n6577) );
  NOR2_X1 U8876 ( .A1(n11767), .A2(n14036), .ZN(n6578) );
  AND2_X1 U8877 ( .A1(n8237), .A2(n8215), .ZN(n6579) );
  AND4_X1 U8878 ( .A1(n10546), .A2(n10545), .A3(n10544), .A4(n10543), .ZN(
        n11031) );
  AND2_X1 U8879 ( .A1(n13779), .A2(n13585), .ZN(n6580) );
  AND2_X1 U8880 ( .A1(n6926), .A2(n6928), .ZN(n6581) );
  AND2_X1 U8881 ( .A1(n13086), .A2(n12988), .ZN(n6582) );
  OR2_X1 U8882 ( .A1(n8696), .A2(n8695), .ZN(n6583) );
  NOR2_X1 U8883 ( .A1(n14716), .A2(n11252), .ZN(n6584) );
  NOR2_X1 U8884 ( .A1(n11996), .A2(n11995), .ZN(n6585) );
  AND2_X1 U8885 ( .A1(n11589), .A2(n12748), .ZN(n6586) );
  OR2_X1 U8886 ( .A1(n9494), .A2(n7364), .ZN(n6587) );
  AND2_X1 U8887 ( .A1(n9597), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n6588) );
  NAND2_X1 U8888 ( .A1(n7535), .A2(n8282), .ZN(n6589) );
  INV_X1 U8889 ( .A(P3_IR_REG_18__SCAN_IN), .ZN(n8306) );
  AND2_X1 U8890 ( .A1(n7835), .A2(n11702), .ZN(n6590) );
  OR2_X1 U8891 ( .A1(n14488), .A2(n14489), .ZN(n6591) );
  AND2_X1 U8892 ( .A1(n9646), .A2(P2_DATAO_REG_8__SCAN_IN), .ZN(n6592) );
  INV_X1 U8893 ( .A(n6825), .ZN(n6824) );
  NAND2_X1 U8894 ( .A1(n6832), .A2(n6829), .ZN(n6825) );
  INV_X1 U8895 ( .A(n13734), .ZN(n6703) );
  INV_X1 U8896 ( .A(n13388), .ZN(n12576) );
  OR2_X1 U8897 ( .A1(n13635), .A2(n13556), .ZN(n13583) );
  AND2_X1 U8898 ( .A1(n12249), .A2(n12938), .ZN(n6593) );
  INV_X1 U8899 ( .A(n6813), .ZN(n6812) );
  NAND2_X1 U8900 ( .A1(n6815), .A2(n6814), .ZN(n6813) );
  INV_X1 U8901 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n9637) );
  NAND2_X1 U8902 ( .A1(n7096), .A2(n13876), .ZN(n6594) );
  AND2_X1 U8903 ( .A1(n6873), .A2(n14574), .ZN(n6595) );
  NAND2_X1 U8904 ( .A1(n12053), .A2(n9432), .ZN(n6596) );
  AND2_X1 U8905 ( .A1(n14135), .A2(n14233), .ZN(n6597) );
  OR2_X1 U8906 ( .A1(n14550), .A2(n14549), .ZN(n6598) );
  OR2_X1 U8907 ( .A1(n11638), .A2(n11556), .ZN(n6599) );
  OR2_X1 U8908 ( .A1(n8256), .A2(n8255), .ZN(n6600) );
  OR2_X1 U8909 ( .A1(n8528), .A2(n8527), .ZN(n6601) );
  AND2_X1 U8910 ( .A1(n6913), .A2(n6599), .ZN(n6602) );
  NOR2_X1 U8911 ( .A1(n12575), .A2(n12574), .ZN(n6603) );
  AND2_X1 U8912 ( .A1(n7072), .A2(n7071), .ZN(n6604) );
  AND2_X1 U8913 ( .A1(n11052), .A2(n11275), .ZN(n6605) );
  AND2_X1 U8914 ( .A1(n6809), .A2(n6534), .ZN(n6606) );
  AND2_X1 U8915 ( .A1(n10201), .A2(n12541), .ZN(n6607) );
  NOR2_X1 U8916 ( .A1(n12614), .A2(n7255), .ZN(n7254) );
  NOR2_X1 U8917 ( .A1(n11248), .A2(n6916), .ZN(n6915) );
  NOR2_X1 U8918 ( .A1(n10375), .A2(n13447), .ZN(n6608) );
  AND2_X1 U8919 ( .A1(n9485), .A2(n6777), .ZN(n6609) );
  OR2_X1 U8920 ( .A1(n10883), .A2(n10366), .ZN(n6610) );
  AND2_X1 U8921 ( .A1(n11445), .A2(n8536), .ZN(n6611) );
  AND2_X1 U8922 ( .A1(n7129), .A2(n6532), .ZN(n6612) );
  OR2_X1 U8923 ( .A1(n8007), .A2(n8009), .ZN(n6613) );
  AND2_X1 U8924 ( .A1(n10563), .A2(n10558), .ZN(n6614) );
  OR2_X1 U8925 ( .A1(n7229), .A2(n8044), .ZN(n6615) );
  NAND2_X1 U8926 ( .A1(n13791), .A2(n13582), .ZN(n6616) );
  OR2_X1 U8927 ( .A1(n8089), .A2(n8091), .ZN(n6617) );
  OR2_X1 U8928 ( .A1(n6525), .A2(n8736), .ZN(n6618) );
  OR2_X1 U8929 ( .A1(n7679), .A2(n7681), .ZN(n6619) );
  OR2_X1 U8930 ( .A1(n9092), .A2(n9091), .ZN(n6620) );
  OR2_X1 U8931 ( .A1(n7414), .A2(n6549), .ZN(n6621) );
  OR2_X1 U8932 ( .A1(n9093), .A2(n9090), .ZN(n6622) );
  AND2_X1 U8933 ( .A1(n8597), .A2(n8564), .ZN(n6623) );
  NAND2_X1 U8934 ( .A1(n8800), .A2(n8799), .ZN(n6624) );
  NAND2_X1 U8935 ( .A1(n8830), .A2(n8831), .ZN(n6625) );
  INV_X1 U8936 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n7114) );
  INV_X1 U8937 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n7487) );
  INV_X1 U8938 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n6734) );
  OR2_X1 U8939 ( .A1(n6928), .A2(n6504), .ZN(n6626) );
  OR2_X1 U8940 ( .A1(n15058), .A2(n13445), .ZN(n6627) );
  NAND2_X1 U8941 ( .A1(n10582), .A2(n10583), .ZN(n7268) );
  INV_X1 U8942 ( .A(n7020), .ZN(n7019) );
  OR2_X1 U8943 ( .A1(n12348), .A2(n12482), .ZN(n7020) );
  OR2_X1 U8944 ( .A1(n13336), .A2(n7252), .ZN(n6628) );
  INV_X1 U8945 ( .A(n12282), .ZN(n12313) );
  INV_X1 U8946 ( .A(n12313), .ZN(n12332) );
  INV_X4 U8947 ( .A(n6932), .ZN(n8684) );
  NAND2_X1 U8948 ( .A1(n14570), .A2(n14898), .ZN(n6875) );
  INV_X1 U8949 ( .A(n11649), .ZN(n9481) );
  INV_X1 U8950 ( .A(n13779), .ZN(n6944) );
  NAND2_X1 U8951 ( .A1(n11140), .A2(n9476), .ZN(n11232) );
  NAND2_X1 U8952 ( .A1(n11354), .A2(n9520), .ZN(n11415) );
  NAND2_X1 U8953 ( .A1(n6917), .A2(n11247), .ZN(n14711) );
  AND2_X1 U8954 ( .A1(n7966), .A2(n9532), .ZN(n14303) );
  INV_X1 U8955 ( .A(n14303), .ZN(n7045) );
  AND4_X1 U8956 ( .A1(n11404), .A2(n11403), .A3(n11402), .A4(n11401), .ZN(
        n11915) );
  INV_X1 U8957 ( .A(n13387), .ZN(n7236) );
  INV_X1 U8958 ( .A(n12358), .ZN(n7029) );
  XNOR2_X1 U8959 ( .A(n13811), .B(n13545), .ZN(n13687) );
  NAND2_X1 U8960 ( .A1(n8977), .A2(n8976), .ZN(n13575) );
  INV_X1 U8961 ( .A(n13575), .ZN(n6709) );
  AND2_X1 U8962 ( .A1(n6875), .A2(n14773), .ZN(n6629) );
  OR2_X1 U8963 ( .A1(n12764), .A2(n8444), .ZN(n6630) );
  INV_X1 U8964 ( .A(n15154), .ZN(n9618) );
  AND2_X1 U8965 ( .A1(n8409), .A2(n8414), .ZN(n15154) );
  AND2_X1 U8966 ( .A1(n7406), .A2(n7405), .ZN(n6631) );
  NAND2_X1 U8967 ( .A1(n12728), .A2(n13039), .ZN(n6632) );
  INV_X1 U8968 ( .A(n9662), .ZN(n7149) );
  NAND2_X1 U8969 ( .A1(n12021), .A2(n6567), .ZN(n13883) );
  AND2_X1 U8970 ( .A1(n7184), .A2(n12123), .ZN(n7183) );
  AND2_X1 U8971 ( .A1(n11516), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n6633) );
  AND2_X1 U8972 ( .A1(n12126), .A2(n12744), .ZN(n6634) );
  AND2_X1 U8973 ( .A1(n7472), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6635) );
  INV_X1 U8974 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n7472) );
  INV_X1 U8975 ( .A(n7319), .ZN(n7318) );
  NAND2_X1 U8976 ( .A1(n7901), .A2(n7932), .ZN(n7319) );
  NOR2_X1 U8977 ( .A1(n11433), .A2(n8485), .ZN(n6636) );
  INV_X1 U8978 ( .A(n12136), .ZN(n7169) );
  OR2_X1 U8979 ( .A1(n12133), .A2(n7169), .ZN(n6637) );
  AND2_X1 U8980 ( .A1(n6739), .A2(n6875), .ZN(n6638) );
  NAND2_X1 U8981 ( .A1(n14146), .A2(n14319), .ZN(n6639) );
  INV_X1 U8982 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7139) );
  INV_X1 U8983 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7142) );
  AND2_X1 U8984 ( .A1(n6892), .A2(n11233), .ZN(n6640) );
  INV_X1 U8985 ( .A(n10323), .ZN(n7154) );
  XOR2_X1 U8986 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .Z(n6641) );
  AND2_X1 U8987 ( .A1(n9662), .A2(n9644), .ZN(n6642) );
  NAND2_X1 U8988 ( .A1(n7856), .A2(n7855), .ZN(n14019) );
  INV_X1 U8989 ( .A(n14019), .ZN(n6904) );
  OR2_X1 U8990 ( .A1(n8336), .A2(n8335), .ZN(n12783) );
  AND2_X1 U8991 ( .A1(n9331), .A2(n9330), .ZN(n6643) );
  AND2_X1 U8992 ( .A1(n8536), .A2(n8537), .ZN(n6644) );
  NAND2_X1 U8993 ( .A1(n7035), .A2(n9516), .ZN(n11158) );
  INV_X1 U8994 ( .A(n6948), .ZN(n10734) );
  INV_X1 U8995 ( .A(n12977), .ZN(n12636) );
  NAND2_X1 U8996 ( .A1(n12214), .A2(n12213), .ZN(n12977) );
  INV_X1 U8997 ( .A(n6828), .ZN(n6827) );
  NAND2_X1 U8998 ( .A1(n11762), .A2(n9325), .ZN(n6828) );
  AND2_X1 U8999 ( .A1(n7057), .A2(n7056), .ZN(n6645) );
  INV_X1 U9000 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n11813) );
  INV_X1 U9001 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n11475) );
  AND2_X1 U9002 ( .A1(n7276), .A2(n11052), .ZN(n6646) );
  AND2_X1 U9003 ( .A1(n6826), .A2(n6828), .ZN(n6647) );
  INV_X1 U9004 ( .A(n14022), .ZN(n13995) );
  INV_X1 U9005 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n6678) );
  INV_X1 U9006 ( .A(n10918), .ZN(n6947) );
  INV_X1 U9007 ( .A(n14849), .ZN(n6786) );
  AND2_X2 U9008 ( .A1(n10382), .A2(n10342), .ZN(n15096) );
  NAND2_X1 U9009 ( .A1(n8477), .A2(n9618), .ZN(n8476) );
  AND2_X2 U9010 ( .A1(n9564), .A2(n9563), .ZN(n14856) );
  INV_X1 U9011 ( .A(n10444), .ZN(n10297) );
  NAND2_X1 U9012 ( .A1(n8682), .A2(n8681), .ZN(n15049) );
  INV_X1 U9013 ( .A(n15049), .ZN(n6701) );
  OR2_X1 U9014 ( .A1(n15139), .A2(n6958), .ZN(n6648) );
  NOR2_X1 U9015 ( .A1(n10433), .A2(n8523), .ZN(n6649) );
  NOR2_X1 U9016 ( .A1(n10435), .A2(n8470), .ZN(n6650) );
  INV_X1 U9017 ( .A(n8546), .ZN(n6975) );
  AND2_X1 U9018 ( .A1(n7068), .A2(n7067), .ZN(n6651) );
  OR2_X1 U9019 ( .A1(n9501), .A2(n9500), .ZN(n14155) );
  AND2_X1 U9020 ( .A1(n12394), .A2(n12392), .ZN(n12509) );
  INV_X1 U9021 ( .A(n12509), .ZN(n7337) );
  INV_X1 U9022 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n11881) );
  AND2_X1 U9023 ( .A1(n10371), .A2(n10370), .ZN(n14997) );
  NOR2_X1 U9024 ( .A1(n15126), .A2(n8382), .ZN(n6652) );
  NAND2_X1 U9025 ( .A1(n12802), .A2(n6975), .ZN(n6653) );
  NAND2_X1 U9026 ( .A1(n13053), .A2(n12367), .ZN(n15261) );
  INV_X1 U9027 ( .A(n15261), .ZN(n15224) );
  AND2_X1 U9028 ( .A1(n6981), .A2(n6980), .ZN(n6654) );
  OR2_X1 U9029 ( .A1(n8550), .A2(n6970), .ZN(n6655) );
  AND2_X1 U9030 ( .A1(n10779), .A2(n12539), .ZN(n15206) );
  AND2_X1 U9031 ( .A1(n6655), .A2(n6969), .ZN(n6656) );
  INV_X1 U9032 ( .A(P3_REG2_REG_14__SCAN_IN), .ZN(n6955) );
  INV_X1 U9033 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n7136) );
  OAI211_X1 U9034 ( .C1(n11445), .C2(n8537), .A(n6963), .B(n6962), .ZN(n11426)
         );
  OR2_X1 U9035 ( .A1(n8536), .A2(n8537), .ZN(n6963) );
  XNOR2_X1 U9036 ( .A(n8484), .B(n8537), .ZN(n11434) );
  INV_X1 U9037 ( .A(n14623), .ZN(n6725) );
  NAND2_X1 U9038 ( .A1(n7245), .A2(n7243), .ZN(n12568) );
  NAND2_X1 U9039 ( .A1(n6553), .A2(n11862), .ZN(n7249) );
  NAND2_X1 U9040 ( .A1(n12577), .A2(n7234), .ZN(n7233) );
  NOR2_X2 U9041 ( .A1(n14703), .A2(n11549), .ZN(n11550) );
  NOR2_X2 U9042 ( .A1(n13536), .A2(n13535), .ZN(n13743) );
  AOI21_X1 U9043 ( .B1(n7376), .B2(n6627), .A(n7375), .ZN(n10567) );
  OAI21_X2 U9044 ( .B1(n14568), .B2(n14603), .A(n14600), .ZN(n14765) );
  NAND2_X1 U9045 ( .A1(n6924), .A2(n10731), .ZN(n10727) );
  NAND3_X1 U9046 ( .A1(n6875), .A2(n6739), .A3(n6595), .ZN(n6659) );
  OAI21_X2 U9047 ( .B1(n10568), .B2(n6920), .A(n6918), .ZN(n10713) );
  NAND2_X1 U9048 ( .A1(n14770), .A2(n14769), .ZN(n14570) );
  OAI21_X2 U9049 ( .B1(n14569), .B2(n14766), .A(n14763), .ZN(n14770) );
  NAND2_X1 U9050 ( .A1(n10355), .A2(n10354), .ZN(n10701) );
  NAND2_X1 U9051 ( .A1(n13726), .A2(n6708), .ZN(n6707) );
  INV_X1 U9052 ( .A(n11795), .ZN(n6705) );
  XNOR2_X1 U9053 ( .A(n6747), .B(n13448), .ZN(n10767) );
  NAND3_X2 U9054 ( .A1(n8648), .A2(n8649), .A3(n6660), .ZN(n13448) );
  NAND2_X1 U9055 ( .A1(n8615), .A2(n6661), .ZN(n8631) );
  NAND3_X1 U9056 ( .A1(n8614), .A2(n9206), .A3(n6662), .ZN(n6661) );
  NAND2_X1 U9057 ( .A1(n9230), .A2(n14990), .ZN(n6662) );
  NAND4_X2 U9058 ( .A1(n6909), .A2(n6906), .A3(n7372), .A4(n6907), .ZN(n9242)
         );
  AOI21_X1 U9059 ( .B1(n7281), .B2(n13408), .A(n6603), .ZN(n7278) );
  NAND3_X1 U9060 ( .A1(n6664), .A2(n6663), .A3(n6625), .ZN(n7428) );
  NAND2_X1 U9061 ( .A1(n8820), .A2(n8819), .ZN(n6663) );
  NAND2_X1 U9062 ( .A1(n8816), .A2(n8815), .ZN(n6664) );
  NAND2_X1 U9063 ( .A1(n6665), .A2(n6620), .ZN(n9110) );
  NAND3_X1 U9064 ( .A1(n9075), .A2(n9074), .A3(n6622), .ZN(n6665) );
  OR2_X1 U9065 ( .A1(n8254), .A2(n9454), .ZN(n6716) );
  NAND2_X1 U9066 ( .A1(n7338), .A2(n7339), .ZN(n8326) );
  NAND2_X1 U9067 ( .A1(n6666), .A2(n8279), .ZN(n8294) );
  NAND3_X1 U9068 ( .A1(n8273), .A2(n8275), .A3(n8274), .ZN(n6666) );
  OAI22_X2 U9069 ( .A1(n12999), .A2(n12844), .B1(n13015), .B2(n13097), .ZN(
        n12986) );
  NAND2_X2 U9070 ( .A1(n13013), .A2(n12843), .ZN(n12999) );
  NAND4_X1 U9071 ( .A1(n8251), .A2(n14150), .A3(n6597), .A4(n6669), .ZN(n6668)
         );
  NOR2_X1 U9072 ( .A1(n7331), .A2(n6670), .ZN(n7333) );
  NOR2_X1 U9073 ( .A1(n13588), .A2(n6533), .ZN(n7302) );
  NOR2_X1 U9074 ( .A1(n7299), .A2(n14997), .ZN(n7297) );
  NOR2_X1 U9075 ( .A1(n14780), .A2(n14779), .ZN(n14778) );
  OAI22_X1 U9076 ( .A1(P3_ADDR_REG_12__SCAN_IN), .A2(n14510), .B1(n14519), 
        .B2(n14521), .ZN(n14573) );
  NOR2_X1 U9077 ( .A1(n14495), .A2(n14494), .ZN(n14554) );
  NOR2_X1 U9078 ( .A1(n14606), .A2(P2_ADDR_REG_18__SCAN_IN), .ZN(n14610) );
  NAND3_X1 U9079 ( .A1(n6876), .A2(n6503), .A3(P1_ADDR_REG_2__SCAN_IN), .ZN(
        n6877) );
  OAI22_X2 U9080 ( .A1(n8152), .A2(n7219), .B1(n8153), .B2(n7218), .ZN(n8229)
         );
  NAND2_X1 U9081 ( .A1(n7222), .A2(n7223), .ZN(n8027) );
  INV_X1 U9082 ( .A(n7214), .ZN(n7213) );
  INV_X1 U9083 ( .A(n7927), .ZN(n7928) );
  NAND2_X1 U9084 ( .A1(n6674), .A2(n6673), .ZN(P3_U3296) );
  NAND2_X1 U9085 ( .A1(n6675), .A2(n10541), .ZN(n6674) );
  NAND2_X1 U9086 ( .A1(n6676), .A2(n6550), .ZN(n6675) );
  NAND2_X1 U9087 ( .A1(n12263), .A2(n12261), .ZN(n7160) );
  OR2_X1 U9088 ( .A1(n12504), .A2(n10997), .ZN(n7162) );
  INV_X1 U9089 ( .A(n11739), .ZN(n7157) );
  NAND2_X1 U9090 ( .A1(n7143), .A2(n9937), .ZN(n10150) );
  NAND2_X1 U9091 ( .A1(n7155), .A2(n7154), .ZN(n7153) );
  OAI21_X1 U9092 ( .B1(n9518), .B2(n7042), .A(n11416), .ZN(n7041) );
  NAND2_X1 U9093 ( .A1(n9531), .A2(n9530), .ZN(n14304) );
  AOI21_X2 U9094 ( .B1(n14262), .B2(n14266), .A(n9533), .ZN(n14247) );
  NAND2_X1 U9095 ( .A1(n11833), .A2(n11832), .ZN(n11831) );
  NAND2_X1 U9096 ( .A1(n6862), .A2(n6516), .ZN(n9566) );
  INV_X1 U9097 ( .A(n8908), .ZN(n6681) );
  NAND2_X1 U9098 ( .A1(n8893), .A2(n8892), .ZN(n8908) );
  INV_X2 U9099 ( .A(n13872), .ZN(n8568) );
  NAND2_X1 U9100 ( .A1(n7490), .A2(P1_IR_REG_27__SCAN_IN), .ZN(n7493) );
  OAI21_X1 U9101 ( .B1(n7991), .B2(n7990), .A(n6613), .ZN(n6755) );
  OAI21_X1 U9102 ( .B1(n7829), .B2(n7828), .A(n7827), .ZN(n7831) );
  NAND4_X1 U9103 ( .A1(n7567), .A2(n7568), .A3(n10509), .A4(n6682), .ZN(n6717)
         );
  OAI22_X2 U9104 ( .A1(n7756), .A2(n7225), .B1(n7755), .B2(n7224), .ZN(n7776)
         );
  NOR2_X2 U9105 ( .A1(n7486), .A2(P1_IR_REG_29__SCAN_IN), .ZN(n7477) );
  NAND2_X2 U9106 ( .A1(n6684), .A2(n10170), .ZN(n10822) );
  NAND2_X1 U9107 ( .A1(n14046), .A2(n9548), .ZN(n10170) );
  NAND2_X1 U9108 ( .A1(n7172), .A2(n13121), .ZN(n8322) );
  NAND2_X1 U9109 ( .A1(n11922), .A2(n11921), .ZN(n12013) );
  NAND2_X1 U9110 ( .A1(n12129), .A2(n12128), .ZN(n12670) );
  NAND2_X1 U9111 ( .A1(n12652), .A2(n12202), .ZN(n12217) );
  NAND2_X1 U9112 ( .A1(n7179), .A2(n7183), .ZN(n7180) );
  NAND2_X1 U9113 ( .A1(n11265), .A2(n11365), .ZN(n11368) );
  NAND2_X1 U9114 ( .A1(n12645), .A2(n12644), .ZN(n12643) );
  NAND2_X1 U9115 ( .A1(n10446), .A2(n10445), .ZN(n10556) );
  NAND2_X1 U9116 ( .A1(n7167), .A2(n7168), .ZN(n12677) );
  AOI21_X1 U9117 ( .B1(n9809), .B2(n11748), .A(n11878), .ZN(n10200) );
  AOI21_X1 U9118 ( .B1(n11113), .B2(n11112), .A(n7441), .ZN(n11115) );
  OR2_X1 U9119 ( .A1(n7488), .A2(n7443), .ZN(n7489) );
  NAND2_X1 U9120 ( .A1(n14359), .A2(n14360), .ZN(n14444) );
  OAI21_X2 U9121 ( .B1(n14168), .B2(n14149), .A(n14150), .ZN(n14148) );
  NAND2_X1 U9122 ( .A1(n6690), .A2(n6688), .ZN(P2_U3186) );
  NAND2_X1 U9123 ( .A1(n13339), .A2(n13338), .ZN(n6690) );
  INV_X1 U9124 ( .A(n7852), .ZN(n7060) );
  INV_X1 U9125 ( .A(n7852), .ZN(n6720) );
  AOI21_X1 U9126 ( .B1(n7246), .B2(n7249), .A(n7244), .ZN(n7243) );
  OAI21_X1 U9127 ( .B1(n7749), .B2(n9628), .A(n7510), .ZN(n6722) );
  INV_X1 U9128 ( .A(n11860), .ZN(n7247) );
  AND2_X2 U9129 ( .A1(n7480), .A2(n7481), .ZN(n7608) );
  NAND2_X1 U9130 ( .A1(n8218), .A2(n6692), .ZN(n8275) );
  NAND2_X1 U9131 ( .A1(n7486), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7474) );
  INV_X1 U9132 ( .A(n12013), .ZN(n7179) );
  NAND3_X1 U9133 ( .A1(n10286), .A2(n10285), .A3(n6552), .ZN(n15190) );
  NAND2_X1 U9134 ( .A1(n12292), .A2(n15202), .ZN(n10299) );
  NAND2_X1 U9135 ( .A1(n9040), .A2(n6621), .ZN(n7411) );
  NAND2_X1 U9136 ( .A1(n6694), .A2(n6693), .ZN(n6737) );
  NAND2_X1 U9137 ( .A1(n8854), .A2(n7431), .ZN(n7430) );
  NAND3_X1 U9138 ( .A1(n7290), .A2(n7289), .A3(n7634), .ZN(n7638) );
  INV_X1 U9139 ( .A(n7577), .ZN(n7595) );
  NOR2_X1 U9140 ( .A1(n6790), .A2(n6794), .ZN(n6788) );
  NAND2_X1 U9141 ( .A1(n6950), .A2(n6949), .ZN(n11966) );
  NAND2_X1 U9142 ( .A1(n13851), .A2(n15066), .ZN(n6699) );
  NAND2_X1 U9143 ( .A1(n13788), .A2(n6700), .ZN(n13851) );
  NOR2_X4 U9144 ( .A1(n13673), .A2(n13795), .ZN(n13657) );
  NAND2_X2 U9145 ( .A1(n13657), .A2(n13640), .ZN(n13642) );
  NOR2_X2 U9146 ( .A1(n14981), .A2(n15058), .ZN(n10744) );
  AOI21_X2 U9147 ( .B1(n6705), .B2(n6541), .A(n7452), .ZN(n11960) );
  NAND2_X2 U9148 ( .A1(n6707), .A2(n6706), .ZN(n13714) );
  NAND2_X1 U9149 ( .A1(n6719), .A2(n6718), .ZN(n8068) );
  NAND2_X1 U9150 ( .A1(n9488), .A2(n7045), .ZN(n14300) );
  AOI21_X1 U9151 ( .B1(n8850), .B2(n8851), .A(n6710), .ZN(n7429) );
  NOR2_X4 U9152 ( .A1(n6952), .A2(n6934), .ZN(n15026) );
  NAND2_X1 U9153 ( .A1(n8718), .A2(n8719), .ZN(n8717) );
  NAND2_X1 U9154 ( .A1(n6583), .A2(n6746), .ZN(n8718) );
  XNOR2_X1 U9155 ( .A(n8002), .B(SI_20_), .ZN(n8001) );
  NAND2_X1 U9156 ( .A1(n7262), .A2(n7261), .ZN(n7263) );
  INV_X1 U9157 ( .A(n13337), .ZN(n6740) );
  NAND2_X1 U9158 ( .A1(n11280), .A2(n11279), .ZN(n11332) );
  NOR2_X1 U9159 ( .A1(n10907), .A2(n10906), .ZN(n10911) );
  NAND2_X1 U9160 ( .A1(n7697), .A2(n7719), .ZN(n9647) );
  OAI22_X2 U9161 ( .A1(n14697), .A2(n6939), .B1(n11559), .B2(n14702), .ZN(
        n11795) );
  OAI21_X1 U9162 ( .B1(n6484), .B2(n9627), .A(n6712), .ZN(n7504) );
  NAND2_X1 U9163 ( .A1(n6479), .A2(n6915), .ZN(n6912) );
  NAND2_X1 U9164 ( .A1(n10871), .A2(n10870), .ZN(n10954) );
  AOI21_X1 U9165 ( .B1(n13572), .B2(n13571), .A(n13570), .ZN(n13740) );
  OAI22_X2 U9166 ( .A1(n7430), .A2(n7429), .B1(n8872), .B2(n8873), .ZN(n8888)
         );
  OAI21_X2 U9167 ( .B1(n7411), .B2(n7412), .A(n7413), .ZN(n9070) );
  NAND2_X1 U9168 ( .A1(n7436), .A2(n7437), .ZN(n8755) );
  NAND2_X1 U9169 ( .A1(n6736), .A2(n7422), .ZN(n9012) );
  NOR2_X1 U9170 ( .A1(n8983), .A2(n7423), .ZN(n6738) );
  NAND2_X1 U9171 ( .A1(n8755), .A2(n8756), .ZN(n8754) );
  NAND2_X1 U9172 ( .A1(n11019), .A2(n12387), .ZN(n11088) );
  INV_X1 U9173 ( .A(n13761), .ZN(n13766) );
  NAND2_X1 U9174 ( .A1(n6744), .A2(n7296), .ZN(n13761) );
  NAND3_X1 U9175 ( .A1(n7438), .A2(n8781), .A3(n6624), .ZN(n7432) );
  AND2_X4 U9176 ( .A1(n11392), .A2(n10187), .ZN(n12282) );
  NAND2_X1 U9177 ( .A1(n10993), .A2(n10992), .ZN(n12378) );
  NAND2_X1 U9178 ( .A1(n13057), .A2(n6764), .ZN(n13301) );
  OAI21_X1 U9179 ( .B1(n12928), .B2(n7020), .A(n7016), .ZN(n7022) );
  AOI22_X1 U9180 ( .A1(n13615), .A2(n13617), .B1(n13586), .B2(n13779), .ZN(
        n13598) );
  OAI21_X1 U9181 ( .B1(n8327), .B2(n8324), .A(n8328), .ZN(n7032) );
  AOI21_X1 U9182 ( .B1(n11769), .B2(n11771), .A(n9527), .ZN(n11833) );
  NAND2_X1 U9183 ( .A1(n11238), .A2(n11239), .ZN(n7035) );
  AOI21_X2 U9184 ( .B1(n14132), .B2(n14324), .A(n6714), .ZN(n14359) );
  INV_X4 U9185 ( .A(n8621), .ZN(n10187) );
  NAND2_X1 U9186 ( .A1(n6740), .A2(n12608), .ZN(n13338) );
  NAND2_X1 U9187 ( .A1(n8579), .A2(n8578), .ZN(n8583) );
  NAND2_X1 U9188 ( .A1(n7272), .A2(n7270), .ZN(n7269) );
  NOR2_X1 U9189 ( .A1(n10635), .A2(n10634), .ZN(n10907) );
  INV_X1 U9190 ( .A(n10273), .ZN(n7262) );
  OAI22_X1 U9191 ( .A1(n10911), .A2(n7275), .B1(n6505), .B2(n6605), .ZN(n11280) );
  NAND2_X1 U9192 ( .A1(n6717), .A2(n7570), .ZN(n7587) );
  NAND2_X1 U9193 ( .A1(n6762), .A2(n6761), .ZN(n8028) );
  NAND2_X1 U9194 ( .A1(n14834), .A2(n14043), .ZN(n8237) );
  NAND2_X2 U9195 ( .A1(n7527), .A2(n8621), .ZN(n7749) );
  NAND3_X1 U9196 ( .A1(n8069), .A2(n8068), .A3(n6617), .ZN(n7217) );
  INV_X1 U9197 ( .A(n8353), .ZN(n7078) );
  INV_X1 U9198 ( .A(n6722), .ZN(n6721) );
  AOI21_X1 U9199 ( .B1(n7494), .B2(P1_IR_REG_31__SCAN_IN), .A(n7487), .ZN(
        n7488) );
  NOR2_X1 U9200 ( .A1(n14622), .A2(n14621), .ZN(n14620) );
  AOI21_X1 U9201 ( .B1(P3_REG2_REG_8__SCAN_IN), .B2(n11206), .A(n10526), .ZN(
        n8533) );
  NOR2_X1 U9202 ( .A1(n8531), .A2(n15146), .ZN(n10528) );
  INV_X1 U9203 ( .A(n7231), .ZN(n9246) );
  NAND2_X1 U9204 ( .A1(n13774), .A2(n6547), .ZN(n13849) );
  AOI21_X1 U9205 ( .B1(n10697), .B2(n10356), .A(n6608), .ZN(n14970) );
  NAND2_X1 U9206 ( .A1(n9598), .A2(n6483), .ZN(n8682) );
  AND2_X4 U9207 ( .A1(n13867), .A2(n13872), .ZN(n9174) );
  XNOR2_X2 U9208 ( .A(n8566), .B(n8565), .ZN(n13867) );
  INV_X1 U9209 ( .A(n8329), .ZN(n7191) );
  NAND2_X1 U9210 ( .A1(n8517), .A2(n15155), .ZN(n6886) );
  NAND2_X1 U9211 ( .A1(n13603), .A2(n6729), .ZN(n13768) );
  NAND2_X1 U9212 ( .A1(n13605), .A2(n13604), .ZN(n13603) );
  INV_X2 U9213 ( .A(n8326), .ZN(n8325) );
  NAND2_X1 U9214 ( .A1(n8556), .A2(n6656), .ZN(n6968) );
  NOR2_X1 U9215 ( .A1(n12780), .A2(n12779), .ZN(n12778) );
  OAI22_X1 U9216 ( .A1(n14970), .A2(n14971), .B1(n15049), .B2(n13446), .ZN(
        n10743) );
  NOR2_X1 U9217 ( .A1(n14629), .A2(n14630), .ZN(n14628) );
  AOI21_X1 U9218 ( .B1(n10706), .B2(n10705), .A(n7374), .ZN(n10732) );
  INV_X1 U9219 ( .A(n8694), .ZN(n6759) );
  NAND2_X1 U9220 ( .A1(n9227), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8590) );
  BUF_X4 U9221 ( .A(n8663), .Z(n9181) );
  INV_X1 U9222 ( .A(n6745), .ZN(n6744) );
  INV_X1 U9223 ( .A(n6735), .ZN(n7438) );
  NAND2_X1 U9224 ( .A1(n6738), .A2(n6737), .ZN(n6736) );
  OAI21_X1 U9225 ( .B1(n13601), .B2(n7298), .A(n13594), .ZN(n6745) );
  NAND2_X1 U9226 ( .A1(n11479), .A2(n11480), .ZN(n9522) );
  NAND2_X1 U9227 ( .A1(n7039), .A2(n7038), .ZN(n11479) );
  INV_X1 U9228 ( .A(n7041), .ZN(n7040) );
  NAND2_X1 U9229 ( .A1(n9526), .A2(n9525), .ZN(n11769) );
  NAND2_X1 U9230 ( .A1(n7046), .A2(n7044), .ZN(n14262) );
  NAND2_X1 U9231 ( .A1(n6877), .A2(P3_ADDR_REG_2__SCAN_IN), .ZN(n7116) );
  NOR2_X1 U9232 ( .A1(n14529), .A2(P1_ADDR_REG_4__SCAN_IN), .ZN(n14491) );
  AOI21_X2 U9233 ( .B1(n14580), .B2(n14579), .A(n14778), .ZN(n14581) );
  NOR2_X2 U9234 ( .A1(n14776), .A2(n14576), .ZN(n14780) );
  NAND2_X1 U9235 ( .A1(n7233), .A2(n7232), .ZN(n12587) );
  NAND2_X1 U9236 ( .A1(n12908), .A2(n12857), .ZN(n12896) );
  OAI21_X1 U9237 ( .B1(n11028), .B2(n11027), .A(n11026), .ZN(n11029) );
  INV_X1 U9238 ( .A(n8524), .ZN(n8525) );
  NOR2_X2 U9239 ( .A1(n14640), .A2(n14639), .ZN(n14638) );
  NAND2_X1 U9240 ( .A1(n9017), .A2(n9016), .ZN(n9037) );
  NAND2_X1 U9241 ( .A1(n8909), .A2(n7453), .ZN(n8942) );
  OAI22_X2 U9242 ( .A1(n13670), .A2(n13672), .B1(n13679), .B2(n13580), .ZN(
        n13666) );
  NAND2_X1 U9243 ( .A1(n6760), .A2(n6759), .ZN(n6746) );
  OAI21_X1 U9244 ( .B1(n10869), .B2(n10868), .A(n10918), .ZN(n10871) );
  AND4_X2 U9245 ( .A1(n8563), .A2(n8562), .A3(n8561), .A4(n8575), .ZN(n6909)
         );
  INV_X1 U9246 ( .A(n10713), .ZN(n6924) );
  NAND2_X1 U9247 ( .A1(n13684), .A2(n13687), .ZN(n13683) );
  NAND2_X1 U9248 ( .A1(n7311), .A2(n13584), .ZN(n13615) );
  NAND2_X1 U9249 ( .A1(n11558), .A2(n11557), .ZN(n14697) );
  NAND2_X1 U9250 ( .A1(n11960), .A2(n11959), .ZN(n6911) );
  OAI21_X1 U9251 ( .B1(n10567), .B2(n10569), .A(n6610), .ZN(n10706) );
  NAND2_X1 U9252 ( .A1(n13698), .A2(n13706), .ZN(n13544) );
  NAND2_X1 U9253 ( .A1(n13688), .A2(n7400), .ZN(n13671) );
  AND2_X4 U9254 ( .A1(n8569), .A2(n8568), .ZN(n8664) );
  INV_X1 U9255 ( .A(n10743), .ZN(n7376) );
  OAI22_X1 U9256 ( .A1(n10732), .A2(n10731), .B1(n10730), .B2(n10729), .ZN(
        n10867) );
  NAND2_X1 U9257 ( .A1(n6938), .A2(n6937), .ZN(P2_U3527) );
  NAND2_X1 U9258 ( .A1(n7378), .A2(n7377), .ZN(n13628) );
  INV_X1 U9259 ( .A(n9998), .ZN(n6935) );
  NAND2_X1 U9260 ( .A1(n10766), .A2(n10767), .ZN(n10345) );
  NAND2_X1 U9261 ( .A1(n7384), .A2(n7382), .ZN(n13712) );
  NOR2_X1 U9262 ( .A1(n11804), .A2(n7410), .ZN(n7403) );
  NAND2_X1 U9263 ( .A1(n7428), .A2(n7425), .ZN(n8850) );
  NAND2_X1 U9264 ( .A1(n7432), .A2(n7433), .ZN(n8817) );
  NOR3_X2 U9265 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), .A3(
        P2_IR_REG_20__SCAN_IN), .ZN(n8563) );
  NAND2_X1 U9266 ( .A1(n7560), .A2(n6750), .ZN(n9289) );
  NAND2_X1 U9267 ( .A1(n7992), .A2(n6754), .ZN(n7222) );
  INV_X1 U9268 ( .A(n6755), .ZN(n6754) );
  OAI21_X1 U9269 ( .B1(n8656), .B2(n8655), .A(n6756), .ZN(n8673) );
  NAND2_X1 U9270 ( .A1(n6758), .A2(n6757), .ZN(n6756) );
  NAND2_X1 U9271 ( .A1(n8656), .A2(n8655), .ZN(n6758) );
  NAND2_X1 U9272 ( .A1(n8696), .A2(n8695), .ZN(n6760) );
  NAND2_X1 U9273 ( .A1(n7486), .A2(n7489), .ZN(n8290) );
  INV_X1 U9274 ( .A(n8229), .ZN(n8218) );
  NAND2_X1 U9275 ( .A1(n7217), .A2(n7216), .ZN(n8109) );
  NAND2_X1 U9276 ( .A1(n7227), .A2(n7228), .ZN(n8067) );
  XNOR2_X1 U9277 ( .A(n6838), .B(n7523), .ZN(n9631) );
  INV_X4 U9278 ( .A(n7749), .ZN(n8212) );
  NAND2_X1 U9279 ( .A1(n12878), .A2(n12862), .ZN(n12883) );
  INV_X1 U9280 ( .A(n6866), .ZN(n14586) );
  NAND2_X1 U9281 ( .A1(n6869), .A2(n6872), .ZN(n14575) );
  NAND2_X1 U9282 ( .A1(n7191), .A2(n7190), .ZN(n8457) );
  NAND2_X1 U9283 ( .A1(n7323), .A2(n7321), .ZN(n12965) );
  NAND2_X1 U9284 ( .A1(n12850), .A2(n12849), .ZN(n12949) );
  NAND2_X1 U9285 ( .A1(n11688), .A2(n11687), .ZN(n11690) );
  AND2_X1 U9286 ( .A1(n10422), .A2(n8349), .ZN(n10155) );
  NAND2_X1 U9287 ( .A1(n6886), .A2(n8516), .ZN(n6885) );
  NAND2_X1 U9288 ( .A1(n10776), .A2(n7141), .ZN(n10961) );
  NAND2_X1 U9289 ( .A1(n12219), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n11743) );
  NAND2_X1 U9290 ( .A1(n9577), .A2(n9576), .ZN(n9605) );
  NAND2_X1 U9291 ( .A1(n7128), .A2(n7126), .ZN(n9636) );
  NAND2_X1 U9292 ( .A1(n9596), .A2(n9595), .ZN(n9581) );
  OAI21_X2 U9293 ( .B1(n10150), .B2(n10149), .A(n10151), .ZN(n7155) );
  OAI21_X2 U9294 ( .B1(n7883), .B2(n7882), .A(n7881), .ZN(n7899) );
  NOR2_X1 U9295 ( .A1(n7595), .A2(n7596), .ZN(n7442) );
  NAND3_X2 U9296 ( .A1(n6529), .A2(n7514), .A3(n7515), .ZN(n14046) );
  INV_X1 U9297 ( .A(n14345), .ZN(n10184) );
  NAND2_X1 U9298 ( .A1(n11414), .A2(n6774), .ZN(n6772) );
  NAND2_X1 U9299 ( .A1(n6773), .A2(n6772), .ZN(n11600) );
  OAI21_X1 U9300 ( .B1(n11839), .B2(n6780), .A(n6779), .ZN(n14333) );
  NAND2_X1 U9301 ( .A1(n6778), .A2(n6609), .ZN(n9487) );
  NAND2_X1 U9302 ( .A1(n11839), .A2(n6779), .ZN(n6778) );
  NAND3_X1 U9303 ( .A1(n6787), .A2(n6784), .A3(n6783), .ZN(P1_U3523) );
  NAND2_X1 U9304 ( .A1(n6795), .A2(n6793), .ZN(n14361) );
  NAND2_X1 U9305 ( .A1(n14363), .A2(n14381), .ZN(n6792) );
  NAND3_X1 U9306 ( .A1(n7102), .A2(n6807), .A3(n6606), .ZN(n6806) );
  NAND3_X1 U9307 ( .A1(n7102), .A2(n6807), .A3(n6534), .ZN(n6817) );
  NAND2_X1 U9308 ( .A1(n7535), .A2(n6835), .ZN(n6834) );
  NAND3_X1 U9309 ( .A1(n7671), .A2(n7465), .A3(n6499), .ZN(n7533) );
  AND3_X1 U9310 ( .A1(n7671), .A2(n7465), .A3(n6837), .ZN(n7535) );
  NAND3_X1 U9311 ( .A1(n6841), .A2(P2_ADDR_REG_19__SCAN_IN), .A3(
        P1_ADDR_REG_19__SCAN_IN), .ZN(n6840) );
  OAI21_X2 U9312 ( .B1(n8022), .B2(n6851), .A(n6849), .ZN(n8080) );
  NAND2_X1 U9313 ( .A1(n8080), .A2(n8079), .ZN(n8083) );
  NAND2_X1 U9314 ( .A1(n7320), .A2(n7318), .ZN(n6857) );
  OR2_X1 U9315 ( .A1(n7836), .A2(n9877), .ZN(n6859) );
  NAND3_X1 U9316 ( .A1(n7076), .A2(n14856), .A3(n7075), .ZN(n6862) );
  OAI21_X2 U9317 ( .B1(n14605), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n6501), .ZN(
        n7119) );
  OAI21_X2 U9318 ( .B1(n14782), .B2(P2_ADDR_REG_16__SCAN_IN), .A(n6506), .ZN(
        n6866) );
  OAI21_X2 U9319 ( .B1(n14531), .B2(P1_ADDR_REG_3__SCAN_IN), .A(n6591), .ZN(
        n6868) );
  NAND3_X1 U9320 ( .A1(n6739), .A2(n6875), .A3(n6873), .ZN(n6869) );
  NAND2_X1 U9321 ( .A1(n14537), .A2(n6878), .ZN(n6876) );
  INV_X1 U9322 ( .A(n14537), .ZN(n14536) );
  INV_X1 U9323 ( .A(n8477), .ZN(n6883) );
  OAI22_X2 U9324 ( .A1(n11433), .A2(n6884), .B1(n7064), .B2(n6633), .ZN(n8487)
         );
  AOI21_X2 U9325 ( .B1(n6887), .B2(n15158), .A(n6885), .ZN(n8556) );
  NAND2_X2 U9326 ( .A1(n8290), .A2(n14059), .ZN(n7527) );
  NAND2_X1 U9327 ( .A1(n9570), .A2(n8212), .ZN(n7560) );
  AND2_X1 U9328 ( .A1(n6889), .A2(n7598), .ZN(n9570) );
  NOR2_X2 U9329 ( .A1(n11142), .A2(n11200), .ZN(n11235) );
  INV_X1 U9330 ( .A(n6894), .ZN(n11350) );
  AOI21_X2 U9331 ( .B1(n13740), .B2(n13574), .A(n6910), .ZN(n13726) );
  NAND2_X1 U9332 ( .A1(n6602), .A2(n6912), .ZN(n11558) );
  AOI21_X1 U9333 ( .B1(n6921), .B2(n6919), .A(n6576), .ZN(n6918) );
  NAND2_X1 U9334 ( .A1(n13714), .A2(n6927), .ZN(n6925) );
  NAND2_X1 U9335 ( .A1(n6925), .A2(n6626), .ZN(n13684) );
  NAND3_X2 U9336 ( .A1(n6931), .A2(n8623), .A3(n8624), .ZN(n9998) );
  AND2_X1 U9337 ( .A1(n8622), .A2(n6936), .ZN(n6931) );
  NOR2_X2 U9338 ( .A1(n8657), .A2(n9572), .ZN(n6934) );
  NOR3_X2 U9339 ( .A1(n13642), .A2(n13635), .A3(n13779), .ZN(n13620) );
  OR2_X1 U9340 ( .A1(n13635), .A2(n13642), .ZN(n13630) );
  NOR2_X2 U9341 ( .A1(n14707), .A2(n11802), .ZN(n6950) );
  NOR2_X2 U9342 ( .A1(n14719), .A2(n11638), .ZN(n6951) );
  OR2_X2 U9343 ( .A1(n13689), .A2(n13806), .ZN(n13673) );
  OR2_X2 U9344 ( .A1(n13701), .A2(n13811), .ZN(n13689) );
  NAND2_X2 U9345 ( .A1(n9250), .A2(n13526), .ZN(n8638) );
  NAND3_X1 U9346 ( .A1(n9250), .A2(n13526), .A3(n8620), .ZN(n6953) );
  OAI21_X1 U9347 ( .B1(n8466), .B2(n6958), .A(n8465), .ZN(n10160) );
  NOR2_X1 U9348 ( .A1(n6958), .A2(P3_U3151), .ZN(n6960) );
  NAND2_X1 U9349 ( .A1(n8348), .A2(n6958), .ZN(n8349) );
  NAND2_X1 U9350 ( .A1(n11445), .A2(n6644), .ZN(n6962) );
  INV_X1 U9351 ( .A(n6964), .ZN(P3_U3201) );
  OAI211_X1 U9352 ( .C1(n12812), .C2(n6968), .A(n6966), .B(n6965), .ZN(n6964)
         );
  AND2_X1 U9353 ( .A1(n6969), .A2(n8551), .ZN(n6967) );
  INV_X1 U9354 ( .A(n8551), .ZN(n6970) );
  NAND2_X1 U9355 ( .A1(n14638), .A2(n10327), .ZN(n6972) );
  NAND3_X1 U9356 ( .A1(n6973), .A2(n6974), .A3(n6972), .ZN(n12790) );
  OAI21_X1 U9357 ( .B1(n14638), .B2(n8546), .A(n10327), .ZN(n12809) );
  NAND2_X1 U9358 ( .A1(n8546), .A2(n10327), .ZN(n6974) );
  INV_X1 U9359 ( .A(n6977), .ZN(n6976) );
  OAI21_X1 U9360 ( .B1(n10418), .B2(n6978), .A(n6982), .ZN(n6977) );
  INV_X1 U9361 ( .A(n8521), .ZN(n6978) );
  NAND2_X1 U9362 ( .A1(n10157), .A2(n6980), .ZN(n6979) );
  OR2_X1 U9363 ( .A1(n10157), .A2(n8521), .ZN(n6981) );
  NAND2_X1 U9364 ( .A1(n8526), .A2(n6986), .ZN(n6984) );
  NAND3_X1 U9365 ( .A1(n6984), .A2(n6983), .A3(n6601), .ZN(n8530) );
  NAND2_X1 U9366 ( .A1(n6993), .A2(n10444), .ZN(n15176) );
  INV_X1 U9367 ( .A(n15190), .ZN(n6993) );
  OAI21_X2 U9368 ( .B1(n15170), .B2(n6997), .A(n6994), .ZN(n11041) );
  AOI21_X1 U9369 ( .B1(n12512), .B2(n6996), .A(n6995), .ZN(n6994) );
  INV_X1 U9370 ( .A(n12378), .ZN(n6996) );
  INV_X1 U9371 ( .A(n12512), .ZN(n6997) );
  OAI21_X1 U9372 ( .B1(n11989), .B2(n12837), .A(n7001), .ZN(n13044) );
  INV_X1 U9373 ( .A(n6998), .ZN(n12305) );
  NAND2_X1 U9374 ( .A1(n11090), .A2(n7007), .ZN(n7004) );
  NAND2_X1 U9375 ( .A1(n7004), .A2(n7005), .ZN(n11388) );
  NAND2_X1 U9376 ( .A1(n11694), .A2(n7011), .ZN(n7010) );
  OAI21_X2 U9377 ( .B1(n13003), .B2(n7026), .A(n7024), .ZN(n12307) );
  NAND2_X1 U9378 ( .A1(n13003), .A2(n12457), .ZN(n12992) );
  NAND2_X2 U9379 ( .A1(n7030), .A2(n7028), .ZN(n13021) );
  NAND2_X4 U9380 ( .A1(n8510), .A2(n6489), .ZN(n11392) );
  INV_X1 U9381 ( .A(n6489), .ZN(n8552) );
  NAND2_X1 U9382 ( .A1(n7035), .A2(n7033), .ZN(n11159) );
  XNOR2_X1 U9383 ( .A(n8493), .B(n10327), .ZN(n12792) );
  NAND2_X1 U9384 ( .A1(n9519), .A2(n7040), .ZN(n7038) );
  NAND2_X2 U9385 ( .A1(n12628), .A2(n14476), .ZN(n8201) );
  NAND3_X1 U9386 ( .A1(n12628), .A2(n14476), .A3(P1_REG0_REG_0__SCAN_IN), .ZN(
        n7043) );
  NOR2_X1 U9387 ( .A1(n9273), .A2(n14046), .ZN(n7561) );
  NAND2_X1 U9388 ( .A1(n14304), .A2(n7047), .ZN(n7046) );
  NOR2_X1 U9389 ( .A1(n14626), .A2(n14627), .ZN(n14625) );
  INV_X1 U9390 ( .A(n14653), .ZN(n7053) );
  XNOR2_X1 U9391 ( .A(n8480), .B(n11306), .ZN(n10851) );
  NAND2_X1 U9392 ( .A1(n8473), .A2(n7069), .ZN(n7065) );
  NAND2_X1 U9393 ( .A1(n14215), .A2(n6604), .ZN(n7070) );
  NAND2_X1 U9394 ( .A1(n9547), .A2(n14324), .ZN(n7076) );
  NAND2_X1 U9395 ( .A1(n7074), .A2(n6515), .ZN(n9561) );
  NAND3_X1 U9396 ( .A1(n7076), .A2(n14849), .A3(n7075), .ZN(n7074) );
  AND2_X1 U9397 ( .A1(n7076), .A2(n6639), .ZN(n12550) );
  NAND2_X1 U9398 ( .A1(n7078), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8355) );
  INV_X1 U9399 ( .A(n7080), .ZN(n7079) );
  NAND2_X1 U9400 ( .A1(n13913), .A2(n9399), .ZN(n7082) );
  NAND2_X1 U9401 ( .A1(n9414), .A2(n7089), .ZN(n7086) );
  NAND2_X1 U9402 ( .A1(n7086), .A2(n7087), .ZN(n12071) );
  NAND2_X1 U9403 ( .A1(n13952), .A2(n13953), .ZN(n13923) );
  NAND2_X1 U9404 ( .A1(n10692), .A2(n10691), .ZN(n10690) );
  NAND2_X1 U9405 ( .A1(n10692), .A2(n7103), .ZN(n7102) );
  NAND2_X1 U9406 ( .A1(n10690), .A2(n9301), .ZN(n10894) );
  NAND2_X1 U9407 ( .A1(n13883), .A2(n9356), .ZN(n9360) );
  NAND2_X1 U9408 ( .A1(n7108), .A2(n7107), .ZN(n13962) );
  AND2_X2 U9409 ( .A1(n9265), .A2(n9499), .ZN(n9275) );
  INV_X1 U9410 ( .A(n7119), .ZN(n14608) );
  INV_X1 U9411 ( .A(n14607), .ZN(n7118) );
  NAND2_X1 U9412 ( .A1(n15283), .A2(n15282), .ZN(n14546) );
  XNOR2_X1 U9413 ( .A(n14530), .B(n7120), .ZN(n15283) );
  XNOR2_X1 U9414 ( .A(n14529), .B(P1_ADDR_REG_4__SCAN_IN), .ZN(n14530) );
  NAND2_X1 U9415 ( .A1(n9586), .A2(n6612), .ZN(n7128) );
  NAND2_X1 U9416 ( .A1(n7146), .A2(n7144), .ZN(n7143) );
  NAND2_X1 U9417 ( .A1(n7148), .A2(n7147), .ZN(n9773) );
  NAND2_X1 U9418 ( .A1(n10559), .A2(n6614), .ZN(n10804) );
  AND2_X1 U9419 ( .A1(n10804), .A2(n10803), .ZN(n10805) );
  NAND2_X1 U9420 ( .A1(n10202), .A2(n6607), .ZN(n7166) );
  NAND2_X1 U9421 ( .A1(n12670), .A2(n12136), .ZN(n7167) );
  NOR2_X2 U9422 ( .A1(n8501), .A2(P3_IR_REG_22__SCAN_IN), .ZN(n7172) );
  NAND2_X1 U9423 ( .A1(n7180), .A2(n6513), .ZN(n12129) );
  NAND2_X1 U9424 ( .A1(n8297), .A2(n8298), .ZN(n8329) );
  NAND4_X1 U9425 ( .A1(n7188), .A2(n8298), .A3(n7186), .A4(n8297), .ZN(n8311)
         );
  NAND4_X1 U9426 ( .A1(n8305), .A2(n8302), .A3(n8303), .A4(n8304), .ZN(n7192)
         );
  NAND2_X1 U9427 ( .A1(n12703), .A2(n12636), .ZN(n7197) );
  NAND2_X1 U9428 ( .A1(n12703), .A2(n7198), .ZN(n7193) );
  AND2_X2 U9429 ( .A1(n7197), .A2(n7196), .ZN(n12685) );
  NAND2_X1 U9430 ( .A1(n7209), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7531) );
  NAND2_X1 U9431 ( .A1(n7210), .A2(n7212), .ZN(n7965) );
  NAND3_X1 U9432 ( .A1(n7916), .A2(n7211), .A3(n6531), .ZN(n7210) );
  NAND3_X1 U9433 ( .A1(n7653), .A2(n7652), .A3(n6619), .ZN(n7220) );
  NAND2_X1 U9434 ( .A1(n7220), .A2(n7221), .ZN(n7703) );
  NAND2_X1 U9435 ( .A1(n7776), .A2(n7777), .ZN(n7775) );
  NAND3_X1 U9436 ( .A1(n8029), .A2(n8028), .A3(n6615), .ZN(n7227) );
  AND2_X4 U9437 ( .A1(n8182), .A2(n7543), .ZN(n8215) );
  NAND2_X1 U9438 ( .A1(n7231), .A2(n6623), .ZN(n8607) );
  INV_X1 U9439 ( .A(n12592), .ZN(n7240) );
  NAND2_X1 U9440 ( .A1(n11861), .A2(n7246), .ZN(n7245) );
  NAND2_X1 U9441 ( .A1(n13337), .A2(n7254), .ZN(n7251) );
  OAI211_X1 U9442 ( .C1(n13337), .C2(n6628), .A(n7253), .B(n7251), .ZN(n12622)
         );
  NAND3_X1 U9443 ( .A1(n7259), .A2(n7260), .A3(n7256), .ZN(n7257) );
  NAND3_X1 U9444 ( .A1(n7258), .A2(n7257), .A3(n7266), .ZN(n10635) );
  NAND3_X1 U9445 ( .A1(n7260), .A2(n7263), .A3(n7259), .ZN(n7258) );
  INV_X1 U9446 ( .A(n10630), .ZN(n7259) );
  NAND2_X1 U9447 ( .A1(n11633), .A2(n7274), .ZN(n7272) );
  NAND2_X1 U9448 ( .A1(n7272), .A2(n7273), .ZN(n11634) );
  INV_X1 U9449 ( .A(n7269), .ZN(n11667) );
  NOR2_X1 U9450 ( .A1(n11635), .A2(n7271), .ZN(n7270) );
  INV_X1 U9451 ( .A(n7273), .ZN(n7271) );
  INV_X1 U9452 ( .A(n7276), .ZN(n11053) );
  INV_X1 U9453 ( .A(n13409), .ZN(n7279) );
  NAND2_X1 U9454 ( .A1(n13409), .A2(n7281), .ZN(n7277) );
  NAND2_X1 U9455 ( .A1(n7816), .A2(n7286), .ZN(n7284) );
  NAND3_X1 U9456 ( .A1(n7294), .A2(n7632), .A3(n7597), .ZN(n7289) );
  NAND3_X1 U9457 ( .A1(n7558), .A2(n7292), .A3(n7294), .ZN(n7290) );
  NAND3_X1 U9458 ( .A1(n7558), .A2(n7294), .A3(n7557), .ZN(n7291) );
  AND2_X1 U9459 ( .A1(n7632), .A2(n7557), .ZN(n7292) );
  INV_X1 U9460 ( .A(n7442), .ZN(n7294) );
  NAND2_X1 U9461 ( .A1(n13601), .A2(n7297), .ZN(n7296) );
  INV_X1 U9462 ( .A(n13647), .ZN(n7312) );
  NAND2_X1 U9463 ( .A1(n7696), .A2(n7695), .ZN(n7719) );
  NAND2_X1 U9464 ( .A1(n7696), .A2(n7314), .ZN(n7313) );
  NAND2_X1 U9465 ( .A1(n7746), .A2(n7767), .ZN(n7747) );
  NAND2_X1 U9466 ( .A1(n12925), .A2(n12856), .ZN(n12908) );
  OAI21_X2 U9467 ( .B1(n12925), .B2(n7325), .A(n7324), .ZN(n12878) );
  NAND2_X1 U9468 ( .A1(n11973), .A2(n11986), .ZN(n11975) );
  NAND2_X1 U9469 ( .A1(n11030), .A2(n6514), .ZN(n7334) );
  INV_X1 U9470 ( .A(n7332), .ZN(n7335) );
  INV_X1 U9471 ( .A(n8457), .ZN(n7338) );
  NAND2_X1 U9472 ( .A1(n11397), .A2(n6497), .ZN(n7342) );
  NAND2_X1 U9473 ( .A1(n7342), .A2(n7343), .ZN(n11686) );
  OAI22_X2 U9474 ( .A1(n13027), .A2(n13031), .B1(n13014), .B2(n13035), .ZN(
        n13011) );
  NAND2_X1 U9475 ( .A1(n8325), .A2(n6544), .ZN(n9920) );
  NAND2_X1 U9476 ( .A1(n8325), .A2(n7345), .ZN(n13322) );
  NAND2_X1 U9477 ( .A1(n10622), .A2(n10620), .ZN(n10621) );
  NAND2_X1 U9478 ( .A1(n11232), .A2(n7350), .ZN(n7349) );
  NAND2_X1 U9479 ( .A1(n14300), .A2(n9489), .ZN(n14281) );
  NAND2_X1 U9480 ( .A1(n11600), .A2(n11599), .ZN(n11598) );
  NOR2_X1 U9481 ( .A1(n11649), .A2(n7357), .ZN(n7356) );
  OAI21_X1 U9482 ( .B1(n14145), .B2(n7360), .A(n7359), .ZN(n7358) );
  NAND2_X1 U9483 ( .A1(n14145), .A2(n14144), .ZN(n14143) );
  INV_X1 U9484 ( .A(n7358), .ZN(n9498) );
  NAND2_X1 U9485 ( .A1(n14143), .A2(n9497), .ZN(n14134) );
  INV_X1 U9486 ( .A(n14234), .ZN(n7366) );
  XNOR2_X2 U9488 ( .A(n7368), .B(n7478), .ZN(n7481) );
  NOR2_X1 U9489 ( .A1(n7477), .A2(n7672), .ZN(n7368) );
  AND3_X2 U9490 ( .A1(n7371), .A2(n7370), .A3(n7369), .ZN(n7372) );
  NOR2_X2 U9491 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_5__SCAN_IN), .ZN(
        n7369) );
  NOR2_X2 U9492 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n7370) );
  NAND2_X1 U9493 ( .A1(n6517), .A2(n7379), .ZN(n7378) );
  NAND2_X1 U9494 ( .A1(n13743), .A2(n7385), .ZN(n7384) );
  INV_X1 U9495 ( .A(n7388), .ZN(n7391) );
  OAI21_X1 U9496 ( .B1(n11250), .B2(n7389), .A(n7393), .ZN(n7388) );
  INV_X1 U9497 ( .A(n11250), .ZN(n7390) );
  OR2_X1 U9498 ( .A1(n10949), .A2(n10953), .ZN(n7392) );
  NAND2_X1 U9499 ( .A1(n13555), .A2(n13554), .ZN(n7399) );
  NAND2_X2 U9500 ( .A1(n13544), .A2(n6507), .ZN(n13688) );
  INV_X1 U9501 ( .A(n13687), .ZN(n7402) );
  NOR2_X1 U9502 ( .A1(n7404), .A2(n7403), .ZN(n13536) );
  INV_X1 U9503 ( .A(n11965), .ZN(n7409) );
  NAND2_X1 U9504 ( .A1(n11804), .A2(n11803), .ZN(n11805) );
  NOR2_X1 U9505 ( .A1(n11959), .A2(n7408), .ZN(n7407) );
  INV_X1 U9506 ( .A(n11803), .ZN(n7408) );
  AND2_X1 U9507 ( .A1(n11964), .A2(n13434), .ZN(n7410) );
  INV_X1 U9508 ( .A(n9053), .ZN(n7414) );
  NAND2_X1 U9509 ( .A1(n8946), .A2(n7417), .ZN(n7416) );
  NAND2_X1 U9510 ( .A1(n8945), .A2(n7417), .ZN(n7415) );
  NAND3_X1 U9511 ( .A1(n7416), .A2(n7415), .A3(n7418), .ZN(n8982) );
  NAND2_X1 U9512 ( .A1(n6526), .A2(n7424), .ZN(n7422) );
  INV_X1 U9513 ( .A(n8996), .ZN(n7424) );
  NAND3_X1 U9514 ( .A1(n8723), .A2(n8722), .A3(n6618), .ZN(n7436) );
  OR2_X1 U9515 ( .A1(n9285), .A2(n9284), .ZN(n9286) );
  NAND2_X1 U9516 ( .A1(n9018), .A2(n8058), .ZN(n11810) );
  XOR2_X1 U9517 ( .A(n9283), .B(n9295), .Z(n9285) );
  AND2_X1 U9518 ( .A1(n10883), .A2(n10744), .ZN(n10572) );
  NAND2_X1 U9519 ( .A1(n7708), .A2(n7707), .ZN(n7731) );
  XNOR2_X1 U9520 ( .A(n13531), .B(n13522), .ZN(n13523) );
  NAND2_X1 U9521 ( .A1(n12340), .A2(n12339), .ZN(n12344) );
  NAND2_X1 U9522 ( .A1(n7592), .A2(n7591), .ZN(n7619) );
  XNOR2_X1 U9523 ( .A(n10389), .B(n15026), .ZN(n10002) );
  NAND2_X1 U9524 ( .A1(n9990), .A2(n13516), .ZN(n10346) );
  OR2_X1 U9525 ( .A1(n13768), .A2(n15061), .ZN(n13774) );
  NAND2_X1 U9526 ( .A1(n7806), .A2(n7805), .ZN(n7829) );
  NAND4_X2 U9527 ( .A1(n7485), .A2(n7484), .A3(n7483), .A4(n7482), .ZN(n14043)
         );
  OR2_X2 U9528 ( .A1(n8205), .A2(n9797), .ZN(n7482) );
  AND2_X1 U9529 ( .A1(n10187), .A2(P2_U3088), .ZN(n12078) );
  XNOR2_X1 U9530 ( .A(n6713), .B(n9991), .ZN(n9990) );
  OR2_X1 U9531 ( .A1(n12827), .A2(n10788), .ZN(n12331) );
  NAND2_X1 U9532 ( .A1(n9998), .A2(n12605), .ZN(n10001) );
  NAND2_X2 U9533 ( .A1(n12375), .A2(n12374), .ZN(n15202) );
  NAND2_X1 U9534 ( .A1(n12755), .A2(n15184), .ZN(n12365) );
  INV_X1 U9535 ( .A(n8817), .ZN(n8820) );
  CLKBUF_X1 U9536 ( .A(n8617), .Z(n8639) );
  INV_X1 U9537 ( .A(n9012), .ZN(n9015) );
  INV_X1 U9538 ( .A(n13867), .ZN(n8569) );
  NAND2_X1 U9539 ( .A1(n11141), .A2(n11148), .ZN(n11140) );
  CLKBUF_X1 U9540 ( .A(n9913), .Z(n14045) );
  INV_X1 U9541 ( .A(n15163), .ZN(n8555) );
  NOR2_X1 U9542 ( .A1(n8657), .A2(n9600), .ZN(n7440) );
  INV_X2 U9543 ( .A(n15211), .ZN(n15213) );
  NOR2_X1 U9544 ( .A1(n11111), .A2(n11110), .ZN(n7441) );
  AND2_X1 U9545 ( .A1(n7487), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7443) );
  AND2_X1 U9546 ( .A1(n9294), .A2(n9293), .ZN(n7444) );
  AND2_X1 U9547 ( .A1(n13766), .A2(n7449), .ZN(n7446) );
  OR2_X1 U9548 ( .A1(n9565), .A2(n14468), .ZN(n7447) );
  OR2_X1 U9549 ( .A1(n9565), .A2(n14423), .ZN(n7448) );
  AND2_X1 U9550 ( .A1(n13765), .A2(n7450), .ZN(n7449) );
  INV_X1 U9551 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n13222) );
  INV_X1 U9552 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n7497) );
  INV_X1 U9553 ( .A(SI_10_), .ZN(n11394) );
  INV_X1 U9554 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n9094) );
  INV_X1 U9555 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n11819) );
  INV_X1 U9556 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n10169) );
  INV_X1 U9557 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n7499) );
  INV_X1 U9558 ( .A(n11885), .ZN(n8279) );
  AND2_X1 U9559 ( .A1(n12332), .A2(SI_30_), .ZN(n7451) );
  INV_X1 U9560 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n12563) );
  INV_X1 U9561 ( .A(n13665), .ZN(n13549) );
  INV_X1 U9562 ( .A(n9174), .ZN(n9150) );
  INV_X1 U9563 ( .A(n13398), .ZN(n12585) );
  AND2_X1 U9564 ( .A1(n11802), .A2(n11796), .ZN(n7452) );
  INV_X1 U9565 ( .A(n14310), .ZN(n14325) );
  XOR2_X1 U9566 ( .A(n12346), .B(n12345), .Z(n7455) );
  NAND2_X1 U9567 ( .A1(n9232), .A2(n9231), .ZN(n7456) );
  NAND2_X2 U9568 ( .A1(n10678), .A2(n14996), .ZN(n15002) );
  INV_X2 U9569 ( .A(n14313), .ZN(n14830) );
  OAI211_X1 U9570 ( .C1(n6945), .C2(n8614), .A(n9205), .B(n9230), .ZN(n8615)
         );
  INV_X1 U9571 ( .A(n8632), .ZN(n8633) );
  INV_X1 U9572 ( .A(n8735), .ZN(n8736) );
  INV_X1 U9573 ( .A(n8778), .ZN(n8779) );
  INV_X1 U9574 ( .A(n8818), .ZN(n8819) );
  INV_X1 U9575 ( .A(n8851), .ZN(n8852) );
  INV_X1 U9576 ( .A(n8889), .ZN(n8890) );
  NAND2_X1 U9577 ( .A1(n7928), .A2(n13949), .ZN(n7929) );
  INV_X1 U9578 ( .A(n8939), .ZN(n8940) );
  OAI21_X1 U9579 ( .B1(n8942), .B2(n8941), .A(n8937), .ZN(n8946) );
  NAND2_X1 U9580 ( .A1(n7968), .A2(n7967), .ZN(n7991) );
  INV_X1 U9581 ( .A(n9013), .ZN(n9014) );
  INV_X2 U9582 ( .A(n8663), .ZN(n9087) );
  INV_X1 U9583 ( .A(n12826), .ZN(n12336) );
  INV_X1 U9584 ( .A(n14662), .ZN(n12337) );
  INV_X1 U9585 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n7466) );
  NAND2_X1 U9586 ( .A1(n12337), .A2(n12336), .ZN(n12338) );
  INV_X1 U9587 ( .A(n12537), .ZN(n12500) );
  INV_X1 U9588 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n8600) );
  INV_X1 U9589 ( .A(SI_12_), .ZN(n7817) );
  INV_X1 U9590 ( .A(P3_REG3_REG_15__SCAN_IN), .ZN(n11944) );
  AOI21_X1 U9591 ( .B1(n8519), .B2(n8518), .A(n8521), .ZN(n8520) );
  INV_X1 U9592 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n12088) );
  AND2_X1 U9593 ( .A1(P2_DATAO_REG_15__SCAN_IN), .A2(n10783), .ZN(n10149) );
  NOR2_X1 U9594 ( .A1(n9144), .A2(n13340), .ZN(n9129) );
  INV_X1 U9595 ( .A(n8970), .ZN(n8968) );
  INV_X1 U9596 ( .A(n11523), .ZN(n9207) );
  AND2_X1 U9597 ( .A1(n8607), .A2(n8606), .ZN(n8608) );
  INV_X1 U9598 ( .A(n9298), .ZN(n9299) );
  INV_X1 U9599 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n7871) );
  INV_X1 U9600 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n7682) );
  AND2_X1 U9601 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_REG3_REG_10__SCAN_IN), 
        .ZN(n7759) );
  INV_X1 U9602 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n7469) );
  INV_X1 U9603 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n7884) );
  INV_X1 U9604 ( .A(P3_REG3_REG_19__SCAN_IN), .ZN(n12167) );
  INV_X1 U9605 ( .A(P3_REG3_REG_20__SCAN_IN), .ZN(n12178) );
  NOR2_X1 U9606 ( .A1(n12152), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n12168) );
  OR2_X1 U9607 ( .A1(n12241), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n12253) );
  OR2_X1 U9608 ( .A1(n12193), .A2(P3_REG3_REG_21__SCAN_IN), .ZN(n12206) );
  INV_X1 U9609 ( .A(n13317), .ZN(n10495) );
  INV_X1 U9610 ( .A(P3_IR_REG_6__SCAN_IN), .ZN(n8406) );
  NAND2_X1 U9611 ( .A1(n10002), .A2(n10001), .ZN(n10005) );
  OR2_X1 U9612 ( .A1(n12566), .A2(n12565), .ZN(n12567) );
  OR2_X1 U9613 ( .A1(n9098), .A2(n9097), .ZN(n9144) );
  INV_X1 U9614 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n9043) );
  NAND2_X1 U9615 ( .A1(n8929), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n8951) );
  INV_X1 U9616 ( .A(n13361), .ZN(n13540) );
  INV_X1 U9617 ( .A(n13591), .ZN(n13420) );
  NAND2_X1 U9618 ( .A1(n9333), .A2(n9334), .ZN(n9335) );
  INV_X1 U9619 ( .A(n8070), .ZN(n8071) );
  INV_X1 U9620 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n13915) );
  OR2_X1 U9621 ( .A1(n7683), .A2(n7682), .ZN(n7711) );
  INV_X1 U9622 ( .A(n14205), .ZN(n14210) );
  INV_X1 U9623 ( .A(n14409), .ZN(n9549) );
  OR2_X1 U9624 ( .A1(n7782), .A2(n11897), .ZN(n7808) );
  INV_X1 U9625 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n7491) );
  INV_X1 U9626 ( .A(SI_22_), .ZN(n8056) );
  INV_X1 U9627 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n7530) );
  OR2_X1 U9628 ( .A1(n7725), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n7750) );
  INV_X1 U9629 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n14487) );
  INV_X1 U9630 ( .A(P3_REG3_REG_23__SCAN_IN), .ZN(n12637) );
  INV_X1 U9631 ( .A(n10562), .ZN(n10563) );
  OR2_X1 U9632 ( .A1(n11979), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n12140) );
  OR2_X1 U9633 ( .A1(n12140), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n12152) );
  NAND2_X1 U9634 ( .A1(n12179), .A2(n12178), .ZN(n12193) );
  AND2_X1 U9635 ( .A1(n11399), .A2(n11431), .ZN(n11534) );
  OR2_X1 U9636 ( .A1(n13294), .A2(n10234), .ZN(n12723) );
  OR2_X1 U9637 ( .A1(n10287), .A2(n13294), .ZN(n12736) );
  AND2_X1 U9638 ( .A1(n8316), .A2(n8315), .ZN(n8320) );
  INV_X1 U9639 ( .A(n12954), .ZN(n12922) );
  INV_X1 U9640 ( .A(n12852), .ZN(n12950) );
  AND2_X1 U9641 ( .A1(n13295), .A2(n15224), .ZN(n10242) );
  AND2_X1 U9642 ( .A1(n10472), .A2(n13295), .ZN(n10473) );
  INV_X1 U9643 ( .A(n11715), .ZN(n12526) );
  AND2_X1 U9644 ( .A1(n13054), .A2(n15262), .ZN(n14680) );
  AND2_X1 U9645 ( .A1(n11000), .A2(n10999), .ZN(n13054) );
  INV_X1 U9646 ( .A(P3_D_REG_1__SCAN_IN), .ZN(n10196) );
  INV_X1 U9647 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n8463) );
  INV_X1 U9648 ( .A(P3_IR_REG_10__SCAN_IN), .ZN(n8330) );
  INV_X1 U9649 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n13340) );
  AND2_X1 U9650 ( .A1(n10051), .A2(n9997), .ZN(n10007) );
  OR2_X1 U9651 ( .A1(n8951), .A2(n13411), .ZN(n8970) );
  AND2_X1 U9652 ( .A1(n9144), .A2(n9099), .ZN(n13632) );
  OR2_X1 U9653 ( .A1(n9044), .A2(n9043), .ZN(n9058) );
  OR2_X1 U9654 ( .A1(n8897), .A2(n11727), .ZN(n8917) );
  OR2_X1 U9655 ( .A1(n10101), .A2(n10100), .ZN(n14888) );
  INV_X1 U9656 ( .A(n13528), .ZN(n13522) );
  NAND2_X1 U9657 ( .A1(n15002), .A2(n10680), .ZN(n14968) );
  OAI21_X1 U9658 ( .B1(n9971), .B2(n9970), .A(n15006), .ZN(n10677) );
  INV_X1 U9659 ( .A(n8058), .ZN(n9019) );
  INV_X1 U9660 ( .A(n14032), .ZN(n11898) );
  INV_X1 U9661 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n13966) );
  NAND2_X1 U9662 ( .A1(n9340), .A2(n9342), .ZN(n9343) );
  INV_X1 U9663 ( .A(n9664), .ZN(n9457) );
  AND2_X1 U9664 ( .A1(n8010), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n8030) );
  INV_X1 U9665 ( .A(n8205), .ZN(n8032) );
  INV_X1 U9666 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n14485) );
  INV_X1 U9667 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n11897) );
  INV_X1 U9668 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n12111) );
  OR2_X1 U9669 ( .A1(n9667), .A2(n7526), .ZN(n7528) );
  XNOR2_X1 U9670 ( .A(n14414), .B(n14029), .ZN(n14332) );
  INV_X1 U9671 ( .A(n14326), .ZN(n14427) );
  INV_X1 U9672 ( .A(n14035), .ZN(n11418) );
  INV_X1 U9673 ( .A(n11767), .ZN(n11345) );
  NAND2_X1 U9674 ( .A1(n10825), .A2(n10824), .ZN(n10823) );
  INV_X1 U9675 ( .A(n9553), .ZN(n9554) );
  AOI21_X1 U9676 ( .B1(P3_ADDR_REG_15__SCAN_IN), .B2(n14816), .A(n14514), .ZN(
        n14584) );
  INV_X1 U9677 ( .A(n12946), .ZN(n13074) );
  INV_X1 U9678 ( .A(n12741), .ZN(n12709) );
  INV_X1 U9679 ( .A(n12723), .ZN(n12733) );
  NAND2_X1 U9680 ( .A1(n10233), .A2(n11001), .ZN(n13297) );
  AND2_X1 U9681 ( .A1(n12259), .A2(n12258), .ZN(n12923) );
  NOR2_X1 U9682 ( .A1(n8544), .A2(n14620), .ZN(n14640) );
  INV_X1 U9683 ( .A(n15139), .ZN(n15153) );
  INV_X1 U9684 ( .A(n13054), .ZN(n15204) );
  AND2_X1 U9685 ( .A1(n13021), .A2(n13020), .ZN(n13099) );
  AND2_X1 U9686 ( .A1(n11002), .A2(n11001), .ZN(n15194) );
  INV_X1 U9687 ( .A(n12421), .ZN(n12522) );
  NOR2_X1 U9688 ( .A1(n15213), .A2(n15186), .ZN(n15209) );
  AND2_X1 U9689 ( .A1(n10474), .A2(n10473), .ZN(n10498) );
  OR2_X1 U9690 ( .A1(n13298), .A2(n13297), .ZN(n13299) );
  NAND2_X1 U9691 ( .A1(n8323), .A2(n8322), .ZN(n8509) );
  INV_X1 U9692 ( .A(P3_IR_REG_21__SCAN_IN), .ZN(n8507) );
  INV_X1 U9693 ( .A(P3_IR_REG_19__SCAN_IN), .ZN(n8459) );
  AND2_X1 U9694 ( .A1(n10187), .A2(P3_U3151), .ZN(n12092) );
  INV_X1 U9695 ( .A(n13428), .ZN(n13391) );
  AND2_X1 U9696 ( .A1(n9989), .A2(n9986), .ZN(n13374) );
  INV_X1 U9697 ( .A(n14992), .ZN(n10348) );
  OR2_X1 U9698 ( .A1(n13621), .A2(n9147), .ZN(n9154) );
  AND2_X1 U9699 ( .A1(n9689), .A2(n9688), .ZN(n14961) );
  INV_X1 U9700 ( .A(n13511), .ZN(n14956) );
  INV_X1 U9701 ( .A(n14968), .ZN(n14715) );
  INV_X1 U9702 ( .A(n14996), .ZN(n14979) );
  INV_X1 U9703 ( .A(n13739), .ZN(n14723) );
  NOR2_X1 U9704 ( .A1(n10675), .A2(n15012), .ZN(n10342) );
  OR2_X1 U9705 ( .A1(n13590), .A2(n13527), .ZN(n13757) );
  INV_X1 U9706 ( .A(n15035), .ZN(n15061) );
  INV_X1 U9707 ( .A(n14997), .ZN(n15064) );
  NAND2_X1 U9708 ( .A1(n10347), .A2(n15076), .ZN(n15035) );
  AND2_X1 U9709 ( .A1(n9982), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9567) );
  INV_X1 U9710 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n9240) );
  AND2_X1 U9711 ( .A1(n8726), .A2(n8761), .ZN(n9847) );
  NAND2_X1 U9712 ( .A1(n9462), .A2(n11885), .ZN(n14016) );
  AND4_X1 U9713 ( .A1(n8209), .A2(n8208), .A3(n8207), .A4(n8206), .ZN(n12074)
         );
  OR2_X1 U9714 ( .A1(n14308), .A2(n8119), .ZN(n7964) );
  INV_X1 U9715 ( .A(n14811), .ZN(n14108) );
  AND2_X1 U9716 ( .A1(n9794), .A2(n14059), .ZN(n14102) );
  INV_X1 U9717 ( .A(n14807), .ZN(n14113) );
  OR2_X1 U9718 ( .A1(n9664), .A2(n8279), .ZN(n9744) );
  NAND2_X1 U9719 ( .A1(n9487), .A2(n9486), .ZN(n14302) );
  NAND2_X1 U9720 ( .A1(n9546), .A2(n9545), .ZN(n14324) );
  INV_X1 U9721 ( .A(n10515), .ZN(n14381) );
  XNOR2_X1 U9722 ( .A(n8172), .B(n8171), .ZN(n13861) );
  INV_X1 U9723 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n7837) );
  AND2_X1 U9724 ( .A1(n8514), .A2(n8513), .ZN(n15097) );
  INV_X1 U9725 ( .A(n12739), .ZN(n12717) );
  NAND2_X1 U9726 ( .A1(n10222), .A2(n13295), .ZN(n12741) );
  INV_X1 U9727 ( .A(n12923), .ZN(n12858) );
  INV_X1 U9728 ( .A(n13015), .ZN(n12987) );
  INV_X1 U9729 ( .A(n11915), .ZN(n12747) );
  OR2_X1 U9730 ( .A1(n8554), .A2(n8552), .ZN(n15136) );
  OR2_X1 U9731 ( .A1(n8554), .A2(n10232), .ZN(n15163) );
  INV_X1 U9732 ( .A(n15209), .ZN(n11224) );
  OR2_X1 U9733 ( .A1(n10485), .A2(n10480), .ZN(n13047) );
  INV_X1 U9734 ( .A(n15281), .ZN(n15279) );
  AND2_X1 U9735 ( .A1(n13300), .A2(n13299), .ZN(n15268) );
  CLKBUF_X1 U9736 ( .A(n9812), .Z(n9829) );
  INV_X1 U9737 ( .A(SI_28_), .ZN(n13329) );
  NAND2_X1 U9738 ( .A1(n8499), .A2(P3_STATE_REG_SCAN_IN), .ZN(n12549) );
  INV_X1 U9739 ( .A(SI_17_), .ZN(n10328) );
  INV_X1 U9740 ( .A(SI_11_), .ZN(n11530) );
  INV_X1 U9741 ( .A(n14702), .ZN(n14735) );
  INV_X1 U9742 ( .A(n13817), .ZN(n13699) );
  INV_X1 U9743 ( .A(n13374), .ZN(n13424) );
  NAND2_X1 U9744 ( .A1(n9136), .A2(n9135), .ZN(n13431) );
  OAI21_X1 U9745 ( .B1(n13675), .B2(n9147), .A(n9050), .ZN(n13580) );
  OR2_X1 U9746 ( .A1(n14870), .A2(P2_U3088), .ZN(n14894) );
  OR2_X1 U9747 ( .A1(n9689), .A2(P2_U3088), .ZN(n14901) );
  AND2_X1 U9748 ( .A1(n13686), .A2(n13685), .ZN(n13813) );
  NAND2_X1 U9749 ( .A1(n15002), .A2(n10679), .ZN(n13739) );
  INV_X1 U9750 ( .A(n15096), .ZN(n15094) );
  AND3_X1 U9751 ( .A1(n15054), .A2(n15053), .A3(n15052), .ZN(n15091) );
  NOR2_X1 U9752 ( .A1(n15013), .A2(n15006), .ZN(n15009) );
  INV_X1 U9753 ( .A(n15009), .ZN(n15010) );
  INV_X1 U9754 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n12278) );
  INV_X1 U9755 ( .A(n14903), .ZN(n13498) );
  INV_X2 U9756 ( .A(n12078), .ZN(n13873) );
  INV_X1 U9757 ( .A(n14016), .ZN(n13989) );
  INV_X1 U9758 ( .A(n14018), .ZN(n13980) );
  NAND2_X1 U9759 ( .A1(n9463), .A2(n9453), .ZN(n14022) );
  NAND4_X1 U9760 ( .A1(n8123), .A2(n8122), .A3(n8121), .A4(n8120), .ZN(n14175)
         );
  INV_X1 U9761 ( .A(n14102), .ZN(n14809) );
  NAND2_X1 U9762 ( .A1(n9794), .A2(n8291), .ZN(n14811) );
  INV_X1 U9763 ( .A(n14277), .ZN(n14334) );
  NAND2_X1 U9764 ( .A1(n14856), .A2(n14426), .ZN(n14423) );
  INV_X2 U9765 ( .A(n14856), .ZN(n14854) );
  INV_X1 U9766 ( .A(n14271), .ZN(n14461) );
  AND2_X2 U9767 ( .A1(n9564), .A2(n9559), .ZN(n14849) );
  AND2_X1 U9768 ( .A1(n9665), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9658) );
  NAND2_X1 U9769 ( .A1(n8278), .A2(P1_STATE_REG_SCAN_IN), .ZN(n11885) );
  INV_X1 U9770 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n11378) );
  INV_X1 U9771 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n10283) );
  INV_X2 U9772 ( .A(n12743), .ZN(P3_U3897) );
  NOR2_X1 U9773 ( .A1(n9983), .A2(n9568), .ZN(P2_U3947) );
  INV_X1 U9774 ( .A(n14044), .ZN(P1_U4016) );
  NOR2_X1 U9775 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_6__SCAN_IN), .ZN(
        n7459) );
  NOR2_X1 U9776 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .ZN(
        n7458) );
  NOR2_X1 U9777 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n7464) );
  NOR2_X1 U9778 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n7463) );
  NOR2_X1 U9779 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n7462) );
  NOR2_X1 U9780 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n7461) );
  NOR2_X1 U9781 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), .ZN(
        n7471) );
  NOR2_X1 U9782 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), .ZN(
        n7470) );
  INV_X1 U9784 ( .A(n7475), .ZN(n14471) );
  NAND2_X4 U9785 ( .A1(n7476), .A2(n14471), .ZN(n14476) );
  INV_X1 U9786 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n7478) );
  INV_X1 U9787 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n7479) );
  OR2_X1 U9788 ( .A1(n8201), .A2(n7479), .ZN(n7485) );
  NAND2_X1 U9789 ( .A1(n7608), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n7484) );
  NAND2_X1 U9790 ( .A1(n8200), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n7483) );
  INV_X1 U9792 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n9797) );
  NAND2_X1 U9793 ( .A1(n7491), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7492) );
  NAND2_X1 U9794 ( .A1(n9582), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n7498) );
  OAI21_X1 U9795 ( .B1(n6484), .B2(n7499), .A(n7498), .ZN(n7500) );
  NAND2_X1 U9796 ( .A1(n7500), .A2(SI_1_), .ZN(n7503) );
  MUX2_X1 U9797 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(P1_DATAO_REG_0__SCAN_IN), 
        .S(n6484), .Z(n7502) );
  NAND2_X1 U9798 ( .A1(n7502), .A2(SI_0_), .ZN(n7523) );
  OAI21_X1 U9799 ( .B1(n7504), .B2(SI_2_), .A(n7553), .ZN(n7505) );
  INV_X1 U9800 ( .A(n7505), .ZN(n7506) );
  NAND2_X1 U9801 ( .A1(n7524), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n7511) );
  INV_X1 U9802 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n7672) );
  OR2_X1 U9803 ( .A1(n7508), .A2(n7672), .ZN(n7509) );
  XNOR2_X1 U9804 ( .A(n7509), .B(P1_IR_REG_2__SCAN_IN), .ZN(n14073) );
  NAND2_X1 U9805 ( .A1(n7954), .A2(n14073), .ZN(n7510) );
  NAND2_X2 U9806 ( .A1(n9282), .A2(n10623), .ZN(n9505) );
  INV_X1 U9807 ( .A(n9505), .ZN(n7517) );
  INV_X1 U9808 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n9795) );
  OR2_X1 U9809 ( .A1(n8205), .A2(n9795), .ZN(n7515) );
  INV_X1 U9810 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n7512) );
  NAND2_X1 U9811 ( .A1(n8200), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n7514) );
  NAND2_X1 U9812 ( .A1(n7608), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n7513) );
  NOR2_X1 U9813 ( .A1(n10187), .A2(n13279), .ZN(n7516) );
  INV_X1 U9814 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n9612) );
  XNOR2_X1 U9815 ( .A(n7516), .B(n9612), .ZN(n14484) );
  MUX2_X1 U9816 ( .A(P1_IR_REG_0__SCAN_IN), .B(n14484), .S(n7527), .Z(n9548)
         );
  INV_X1 U9817 ( .A(n9548), .ZN(n9273) );
  NOR2_X1 U9818 ( .A1(n7517), .A2(n7561), .ZN(n7545) );
  INV_X1 U9819 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n14341) );
  OR2_X1 U9820 ( .A1(n8205), .A2(n14341), .ZN(n7522) );
  INV_X1 U9821 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n7518) );
  NAND2_X1 U9822 ( .A1(n8200), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n7520) );
  NAND2_X1 U9823 ( .A1(n7608), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n7519) );
  INV_X1 U9824 ( .A(n9913), .ZN(n9277) );
  AND2_X1 U9825 ( .A1(n7527), .A2(n10187), .ZN(n7524) );
  NAND2_X1 U9826 ( .A1(n7524), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n7529) );
  NAND2_X1 U9827 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n7525) );
  XNOR2_X1 U9828 ( .A(n7525), .B(P1_IR_REG_1__SCAN_IN), .ZN(n14052) );
  INV_X1 U9829 ( .A(n14052), .ZN(n7526) );
  NAND2_X1 U9830 ( .A1(n9277), .A2(n14345), .ZN(n8239) );
  NAND2_X1 U9831 ( .A1(n7533), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7534) );
  MUX2_X1 U9832 ( .A(P1_IR_REG_31__SCAN_IN), .B(n7534), .S(
        P1_IR_REG_19__SCAN_IN), .Z(n7536) );
  INV_X1 U9833 ( .A(n7535), .ZN(n7539) );
  NAND2_X2 U9834 ( .A1(n7536), .A2(n7539), .ZN(n12108) );
  NAND2_X1 U9835 ( .A1(n6519), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7537) );
  MUX2_X1 U9836 ( .A(P1_IR_REG_31__SCAN_IN), .B(n7537), .S(
        P1_IR_REG_21__SCAN_IN), .Z(n7538) );
  NAND2_X1 U9837 ( .A1(n7539), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7540) );
  MUX2_X1 U9838 ( .A(P1_IR_REG_31__SCAN_IN), .B(n7540), .S(
        P1_IR_REG_20__SCAN_IN), .Z(n7541) );
  INV_X1 U9839 ( .A(n11493), .ZN(n8181) );
  NAND2_X1 U9840 ( .A1(n8179), .A2(n8181), .ZN(n9545) );
  NAND2_X1 U9841 ( .A1(n8195), .A2(n9545), .ZN(n8182) );
  NAND2_X1 U9842 ( .A1(n7542), .A2(n8181), .ZN(n7543) );
  NAND2_X1 U9843 ( .A1(n10822), .A2(n9264), .ZN(n7544) );
  NAND4_X1 U9844 ( .A1(n7545), .A2(n8239), .A3(n8216), .A4(n7544), .ZN(n7568)
         );
  NAND2_X1 U9845 ( .A1(n8200), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n7549) );
  INV_X1 U9846 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n10600) );
  OR2_X1 U9847 ( .A1(n8205), .A2(n10600), .ZN(n7548) );
  INV_X1 U9848 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n7546) );
  OR2_X1 U9849 ( .A1(n8201), .A2(n7546), .ZN(n7547) );
  NAND4_X4 U9850 ( .A1(n7550), .A2(n7549), .A3(n7548), .A4(n7547), .ZN(n14042)
         );
  INV_X1 U9851 ( .A(n14042), .ZN(n9471) );
  OR2_X1 U9852 ( .A1(n7551), .A2(n7672), .ZN(n7552) );
  INV_X1 U9853 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n7581) );
  XNOR2_X1 U9854 ( .A(n7552), .B(n7581), .ZN(n14090) );
  MUX2_X1 U9855 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(P1_DATAO_REG_3__SCAN_IN), 
        .S(n6484), .Z(n7555) );
  NAND2_X1 U9856 ( .A1(n7555), .A2(SI_3_), .ZN(n7593) );
  OAI21_X1 U9857 ( .B1(n7555), .B2(SI_3_), .A(n7593), .ZN(n7556) );
  INV_X1 U9858 ( .A(n7556), .ZN(n7557) );
  NAND2_X1 U9859 ( .A1(n7524), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n7559) );
  NAND2_X1 U9860 ( .A1(n14042), .A2(n10518), .ZN(n7569) );
  NAND2_X1 U9861 ( .A1(n7561), .A2(n8238), .ZN(n9504) );
  OR2_X1 U9862 ( .A1(n9505), .A2(n8215), .ZN(n7566) );
  NAND3_X1 U9863 ( .A1(n6579), .A2(n9505), .A3(n8239), .ZN(n7565) );
  NAND3_X1 U9864 ( .A1(n8237), .A2(n8238), .A3(n8216), .ZN(n7564) );
  INV_X1 U9865 ( .A(n8237), .ZN(n7562) );
  NAND2_X1 U9866 ( .A1(n7562), .A2(n8215), .ZN(n7563) );
  NAND4_X1 U9867 ( .A1(n7565), .A2(n7566), .A3(n7564), .A4(n7563), .ZN(n7567)
         );
  MUX2_X1 U9868 ( .A(n9506), .B(n7569), .S(n8215), .Z(n7570) );
  NAND2_X1 U9869 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n7610) );
  OAI21_X1 U9870 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(n7610), .ZN(n10835) );
  OR2_X1 U9871 ( .A1(n7623), .A2(n10835), .ZN(n7575) );
  NAND2_X1 U9872 ( .A1(n8137), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n7574) );
  INV_X1 U9873 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n7571) );
  OR2_X1 U9874 ( .A1(n8185), .A2(n7571), .ZN(n7573) );
  INV_X1 U9875 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n10830) );
  OR2_X1 U9876 ( .A1(n8205), .A2(n10830), .ZN(n7572) );
  MUX2_X1 U9877 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(P1_DATAO_REG_4__SCAN_IN), 
        .S(n6484), .Z(n7576) );
  NAND2_X1 U9878 ( .A1(n7576), .A2(SI_4_), .ZN(n7594) );
  OAI21_X1 U9879 ( .B1(n7576), .B2(SI_4_), .A(n7594), .ZN(n7577) );
  NAND2_X1 U9880 ( .A1(n7578), .A2(n7595), .ZN(n7580) );
  NAND2_X1 U9881 ( .A1(n9598), .A2(n8212), .ZN(n7584) );
  INV_X4 U9882 ( .A(n7823), .ZN(n8173) );
  NAND2_X1 U9883 ( .A1(n7551), .A2(n7581), .ZN(n7600) );
  NAND2_X1 U9884 ( .A1(n7600), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7582) );
  XNOR2_X1 U9885 ( .A(n7582), .B(P1_IR_REG_4__SCAN_IN), .ZN(n9799) );
  AOI22_X1 U9886 ( .A1(n8173), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n6753), .B2(
        n9799), .ZN(n7583) );
  NAND2_X1 U9887 ( .A1(n7584), .A2(n7583), .ZN(n10837) );
  NAND2_X1 U9888 ( .A1(n7587), .A2(n7588), .ZN(n7586) );
  MUX2_X1 U9889 ( .A(n10837), .B(n14041), .S(n8176), .Z(n7585) );
  NAND2_X1 U9890 ( .A1(n7586), .A2(n7585), .ZN(n7592) );
  INV_X1 U9891 ( .A(n7587), .ZN(n7590) );
  INV_X1 U9892 ( .A(n7588), .ZN(n7589) );
  NAND2_X1 U9893 ( .A1(n7590), .A2(n7589), .ZN(n7591) );
  INV_X1 U9894 ( .A(n7594), .ZN(n7596) );
  MUX2_X1 U9895 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(P1_DATAO_REG_5__SCAN_IN), 
        .S(n6484), .Z(n7599) );
  NAND2_X1 U9896 ( .A1(n7599), .A2(SI_5_), .ZN(n7634) );
  OAI21_X1 U9897 ( .B1(n7599), .B2(SI_5_), .A(n7634), .ZN(n7631) );
  XNOR2_X1 U9898 ( .A(n7633), .B(n7631), .ZN(n9619) );
  NAND2_X1 U9899 ( .A1(n9619), .A2(n8212), .ZN(n7607) );
  OR2_X1 U9900 ( .A1(n7600), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n7602) );
  NAND2_X1 U9901 ( .A1(n7602), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7601) );
  MUX2_X1 U9902 ( .A(P1_IR_REG_31__SCAN_IN), .B(n7601), .S(
        P1_IR_REG_5__SCAN_IN), .Z(n7605) );
  INV_X1 U9903 ( .A(n7602), .ZN(n7604) );
  INV_X1 U9904 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n7603) );
  NAND2_X1 U9905 ( .A1(n7604), .A2(n7603), .ZN(n7640) );
  NAND2_X1 U9906 ( .A1(n7605), .A2(n7640), .ZN(n9884) );
  INV_X1 U9907 ( .A(n9884), .ZN(n9880) );
  AOI22_X1 U9908 ( .A1(n8173), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n6753), .B2(
        n9880), .ZN(n7606) );
  NAND2_X1 U9909 ( .A1(n7607), .A2(n7606), .ZN(n10897) );
  NAND2_X1 U9910 ( .A1(n8137), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n7616) );
  INV_X1 U9911 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n7609) );
  NOR2_X1 U9912 ( .A1(n7610), .A2(n7609), .ZN(n7624) );
  AND2_X1 U9913 ( .A1(n7610), .A2(n7609), .ZN(n7611) );
  NOR2_X1 U9914 ( .A1(n7624), .A2(n7611), .ZN(n10902) );
  NAND2_X1 U9915 ( .A1(n7608), .A2(n10902), .ZN(n7615) );
  INV_X1 U9916 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n7612) );
  OR2_X1 U9917 ( .A1(n8201), .A2(n7612), .ZN(n7614) );
  INV_X1 U9918 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n9883) );
  OR2_X1 U9919 ( .A1(n8205), .A2(n9883), .ZN(n7613) );
  NAND4_X1 U9920 ( .A1(n7616), .A2(n7615), .A3(n7614), .A4(n7613), .ZN(n14040)
         );
  MUX2_X1 U9921 ( .A(n10897), .B(n14040), .S(n8176), .Z(n7620) );
  NAND2_X1 U9922 ( .A1(n7619), .A2(n7620), .ZN(n7618) );
  MUX2_X1 U9923 ( .A(n14040), .B(n10897), .S(n8176), .Z(n7617) );
  NAND2_X1 U9924 ( .A1(n7618), .A2(n7617), .ZN(n7647) );
  INV_X1 U9925 ( .A(n7619), .ZN(n7622) );
  INV_X1 U9926 ( .A(n7620), .ZN(n7621) );
  NAND2_X1 U9927 ( .A1(n7622), .A2(n7621), .ZN(n7650) );
  NAND2_X1 U9928 ( .A1(n7647), .A2(n7650), .ZN(n7644) );
  NAND2_X1 U9929 ( .A1(n7624), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n7655) );
  OR2_X1 U9930 ( .A1(n7624), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n7625) );
  NAND2_X1 U9931 ( .A1(n7655), .A2(n7625), .ZN(n14000) );
  OR2_X1 U9932 ( .A1(n8119), .A2(n14000), .ZN(n7630) );
  NAND2_X1 U9933 ( .A1(n8137), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n7629) );
  INV_X1 U9934 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n7626) );
  OR2_X1 U9935 ( .A1(n8185), .A2(n7626), .ZN(n7628) );
  INV_X1 U9936 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n10942) );
  OR2_X1 U9937 ( .A1(n8205), .A2(n10942), .ZN(n7627) );
  NAND4_X1 U9938 ( .A1(n7630), .A2(n7629), .A3(n7628), .A4(n7627), .ZN(n14039)
         );
  INV_X1 U9939 ( .A(n7631), .ZN(n7632) );
  MUX2_X1 U9940 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(P1_DATAO_REG_6__SCAN_IN), 
        .S(n9582), .Z(n7635) );
  NAND2_X1 U9941 ( .A1(n7635), .A2(SI_6_), .ZN(n7663) );
  OAI21_X1 U9942 ( .B1(SI_6_), .B2(n7635), .A(n7663), .ZN(n7636) );
  INV_X1 U9943 ( .A(n7636), .ZN(n7637) );
  NAND2_X1 U9944 ( .A1(n7638), .A2(n7637), .ZN(n7664) );
  OR2_X1 U9945 ( .A1(n7638), .A2(n7637), .ZN(n7639) );
  NAND2_X1 U9946 ( .A1(n7664), .A2(n7639), .ZN(n9633) );
  OR2_X1 U9947 ( .A1(n9633), .A2(n7749), .ZN(n7643) );
  NAND2_X1 U9948 ( .A1(n7640), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7641) );
  XNOR2_X1 U9949 ( .A(n7641), .B(P1_IR_REG_6__SCAN_IN), .ZN(n9885) );
  AOI22_X1 U9950 ( .A1(n8173), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n6753), .B2(
        n9885), .ZN(n7642) );
  NAND2_X1 U9951 ( .A1(n7643), .A2(n7642), .ZN(n14002) );
  MUX2_X1 U9952 ( .A(n14039), .B(n14002), .S(n8176), .Z(n7648) );
  NAND2_X1 U9953 ( .A1(n7644), .A2(n7648), .ZN(n7646) );
  MUX2_X1 U9954 ( .A(n14002), .B(n14039), .S(n8176), .Z(n7645) );
  NAND2_X1 U9955 ( .A1(n7646), .A2(n7645), .ZN(n7653) );
  INV_X1 U9956 ( .A(n7648), .ZN(n7649) );
  AND2_X1 U9957 ( .A1(n7650), .A2(n7649), .ZN(n7651) );
  NAND2_X1 U9958 ( .A1(n7647), .A2(n7651), .ZN(n7652) );
  NAND2_X1 U9959 ( .A1(n7655), .A2(n7654), .ZN(n7656) );
  NAND2_X1 U9960 ( .A1(n7683), .A2(n7656), .ZN(n11195) );
  OR2_X1 U9961 ( .A1(n8119), .A2(n11195), .ZN(n7662) );
  NAND2_X1 U9962 ( .A1(n8137), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n7661) );
  INV_X1 U9963 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n7657) );
  OR2_X1 U9964 ( .A1(n8201), .A2(n7657), .ZN(n7660) );
  INV_X1 U9965 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n7658) );
  OR2_X1 U9966 ( .A1(n8205), .A2(n7658), .ZN(n7659) );
  NAND4_X1 U9967 ( .A1(n7662), .A2(n7661), .A3(n7660), .A4(n7659), .ZN(n14038)
         );
  NAND2_X1 U9968 ( .A1(n7664), .A2(n7663), .ZN(n7668) );
  MUX2_X1 U9969 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(P1_DATAO_REG_7__SCAN_IN), 
        .S(n10187), .Z(n7665) );
  NAND2_X1 U9970 ( .A1(n7665), .A2(SI_7_), .ZN(n7691) );
  OAI21_X1 U9971 ( .B1(n7665), .B2(SI_7_), .A(n7691), .ZN(n7666) );
  INV_X1 U9972 ( .A(n7666), .ZN(n7667) );
  NAND2_X1 U9973 ( .A1(n7668), .A2(n7667), .ZN(n7692) );
  OR2_X1 U9974 ( .A1(n7668), .A2(n7667), .ZN(n7669) );
  NAND2_X1 U9975 ( .A1(n7692), .A2(n7669), .ZN(n9639) );
  OR2_X1 U9976 ( .A1(n9639), .A2(n7749), .ZN(n7678) );
  NOR2_X1 U9977 ( .A1(n7671), .A2(n7672), .ZN(n7673) );
  MUX2_X1 U9978 ( .A(n7672), .B(n7673), .S(P1_IR_REG_7__SCAN_IN), .Z(n7676) );
  INV_X1 U9979 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n7674) );
  NAND2_X1 U9980 ( .A1(n7671), .A2(n7674), .ZN(n7725) );
  INV_X1 U9981 ( .A(n7725), .ZN(n7675) );
  NOR2_X1 U9982 ( .A1(n7676), .A2(n7675), .ZN(n10011) );
  AOI22_X1 U9983 ( .A1(n8173), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n6753), .B2(
        n10011), .ZN(n7677) );
  MUX2_X1 U9984 ( .A(n14038), .B(n11200), .S(n8215), .Z(n7680) );
  MUX2_X1 U9985 ( .A(n14038), .B(n11200), .S(n8176), .Z(n7679) );
  INV_X1 U9986 ( .A(n7680), .ZN(n7681) );
  NAND2_X1 U9987 ( .A1(n7683), .A2(n7682), .ZN(n7684) );
  NAND2_X1 U9988 ( .A1(n7711), .A2(n7684), .ZN(n11469) );
  OR2_X1 U9989 ( .A1(n8119), .A2(n11469), .ZN(n7690) );
  NAND2_X1 U9990 ( .A1(n8137), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n7689) );
  INV_X1 U9991 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n7685) );
  OR2_X1 U9992 ( .A1(n8185), .A2(n7685), .ZN(n7688) );
  INV_X1 U9993 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n7686) );
  OR2_X1 U9994 ( .A1(n8205), .A2(n7686), .ZN(n7687) );
  NAND4_X1 U9995 ( .A1(n7690), .A2(n7689), .A3(n7688), .A4(n7687), .ZN(n14037)
         );
  NAND2_X1 U9996 ( .A1(n7692), .A2(n7691), .ZN(n7696) );
  MUX2_X1 U9997 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(P1_DATAO_REG_8__SCAN_IN), 
        .S(n10187), .Z(n7693) );
  NAND2_X1 U9998 ( .A1(n7693), .A2(SI_8_), .ZN(n7718) );
  OAI21_X1 U9999 ( .B1(SI_8_), .B2(n7693), .A(n7718), .ZN(n7694) );
  INV_X1 U10000 ( .A(n7694), .ZN(n7695) );
  OR2_X1 U10001 ( .A1(n7696), .A2(n7695), .ZN(n7697) );
  OR2_X1 U10002 ( .A1(n9647), .A2(n7749), .ZN(n7700) );
  NAND2_X1 U10003 ( .A1(n7725), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7698) );
  XNOR2_X1 U10004 ( .A(n7698), .B(P1_IR_REG_8__SCAN_IN), .ZN(n10023) );
  AOI22_X1 U10005 ( .A1(n8173), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n6753), .B2(
        n10023), .ZN(n7699) );
  NAND2_X1 U10006 ( .A1(n7700), .A2(n7699), .ZN(n11471) );
  MUX2_X1 U10007 ( .A(n14037), .B(n11471), .S(n8176), .Z(n7704) );
  NAND2_X1 U10008 ( .A1(n7703), .A2(n7704), .ZN(n7702) );
  MUX2_X1 U10009 ( .A(n14037), .B(n11471), .S(n8215), .Z(n7701) );
  NAND2_X1 U10010 ( .A1(n7702), .A2(n7701), .ZN(n7708) );
  INV_X1 U10011 ( .A(n7703), .ZN(n7706) );
  INV_X1 U10012 ( .A(n7704), .ZN(n7705) );
  NAND2_X1 U10013 ( .A1(n7706), .A2(n7705), .ZN(n7707) );
  NAND2_X1 U10014 ( .A1(n8033), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n7717) );
  INV_X1 U10015 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n7709) );
  OR2_X1 U10016 ( .A1(n8036), .A2(n7709), .ZN(n7716) );
  INV_X1 U10017 ( .A(n7760), .ZN(n7713) );
  NAND2_X1 U10018 ( .A1(n7711), .A2(n7710), .ZN(n7712) );
  NAND2_X1 U10019 ( .A1(n7713), .A2(n7712), .ZN(n11166) );
  OR2_X1 U10020 ( .A1(n8119), .A2(n11166), .ZN(n7715) );
  INV_X1 U10021 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n10012) );
  OR2_X1 U10022 ( .A1(n8205), .A2(n10012), .ZN(n7714) );
  INV_X1 U10023 ( .A(n11465), .ZN(n14036) );
  MUX2_X1 U10024 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(P1_DATAO_REG_9__SCAN_IN), 
        .S(n10187), .Z(n7720) );
  NAND2_X1 U10025 ( .A1(n7720), .A2(SI_9_), .ZN(n7742) );
  OAI21_X1 U10026 ( .B1(n7720), .B2(SI_9_), .A(n7742), .ZN(n7721) );
  INV_X1 U10027 ( .A(n7721), .ZN(n7722) );
  OR2_X1 U10028 ( .A1(n7723), .A2(n7722), .ZN(n7724) );
  NAND2_X1 U10029 ( .A1(n7743), .A2(n7724), .ZN(n9652) );
  OR2_X1 U10030 ( .A1(n9652), .A2(n7749), .ZN(n7728) );
  NAND2_X1 U10031 ( .A1(n7750), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7726) );
  XNOR2_X1 U10032 ( .A(n7726), .B(P1_IR_REG_9__SCAN_IN), .ZN(n10042) );
  AOI22_X1 U10033 ( .A1(n8173), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n6753), .B2(
        n10042), .ZN(n7727) );
  MUX2_X1 U10034 ( .A(n14036), .B(n11767), .S(n8215), .Z(n7732) );
  NAND2_X1 U10035 ( .A1(n7731), .A2(n7732), .ZN(n7730) );
  MUX2_X1 U10036 ( .A(n14036), .B(n11767), .S(n8176), .Z(n7729) );
  NAND2_X1 U10037 ( .A1(n7730), .A2(n7729), .ZN(n7736) );
  INV_X1 U10038 ( .A(n7731), .ZN(n7734) );
  INV_X1 U10039 ( .A(n7732), .ZN(n7733) );
  NAND2_X1 U10040 ( .A1(n7734), .A2(n7733), .ZN(n7735) );
  NAND2_X1 U10041 ( .A1(n7736), .A2(n7735), .ZN(n7756) );
  XNOR2_X1 U10042 ( .A(n7760), .B(P1_REG3_REG_10__SCAN_IN), .ZN(n11661) );
  OR2_X1 U10043 ( .A1(n8119), .A2(n11661), .ZN(n7741) );
  NAND2_X1 U10044 ( .A1(n8137), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n7740) );
  INV_X1 U10045 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n7737) );
  OR2_X1 U10046 ( .A1(n8185), .A2(n7737), .ZN(n7739) );
  INV_X1 U10047 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n11357) );
  OR2_X1 U10048 ( .A1(n8205), .A2(n11357), .ZN(n7738) );
  NAND4_X1 U10049 ( .A1(n7741), .A2(n7740), .A3(n7739), .A4(n7738), .ZN(n14035) );
  MUX2_X1 U10050 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(P1_DATAO_REG_10__SCAN_IN), 
        .S(n10187), .Z(n7744) );
  NAND2_X1 U10051 ( .A1(n7747), .A2(n11394), .ZN(n7748) );
  NAND2_X1 U10052 ( .A1(n7768), .A2(n7748), .ZN(n9777) );
  OR2_X1 U10053 ( .A1(n9777), .A2(n7749), .ZN(n7753) );
  NOR2_X1 U10054 ( .A1(n7750), .A2(P1_IR_REG_9__SCAN_IN), .ZN(n7770) );
  OR2_X1 U10055 ( .A1(n7770), .A2(n7672), .ZN(n7751) );
  XNOR2_X1 U10056 ( .A(n7751), .B(P1_IR_REG_10__SCAN_IN), .ZN(n10120) );
  AOI22_X1 U10057 ( .A1(n8173), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n6753), 
        .B2(n10120), .ZN(n7752) );
  NAND2_X2 U10058 ( .A1(n7753), .A2(n7752), .ZN(n11663) );
  MUX2_X1 U10059 ( .A(n14035), .B(n11663), .S(n8176), .Z(n7755) );
  MUX2_X1 U10060 ( .A(n14035), .B(n11663), .S(n8150), .Z(n7754) );
  NAND2_X1 U10061 ( .A1(n7760), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n7758) );
  INV_X1 U10062 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n7757) );
  NAND2_X1 U10063 ( .A1(n7758), .A2(n7757), .ZN(n7761) );
  NAND2_X1 U10064 ( .A1(n7760), .A2(n7759), .ZN(n7782) );
  NAND2_X1 U10065 ( .A1(n7761), .A2(n7782), .ZN(n11825) );
  OR2_X1 U10066 ( .A1(n8119), .A2(n11825), .ZN(n7766) );
  NAND2_X1 U10067 ( .A1(n8137), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n7765) );
  INV_X1 U10068 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n7762) );
  OR2_X1 U10069 ( .A1(n8201), .A2(n7762), .ZN(n7764) );
  INV_X1 U10070 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n11419) );
  OR2_X1 U10071 ( .A1(n8205), .A2(n11419), .ZN(n7763) );
  NAND4_X1 U10072 ( .A1(n7766), .A2(n7765), .A3(n7764), .A4(n7763), .ZN(n14034) );
  MUX2_X1 U10073 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(P1_DATAO_REG_11__SCAN_IN), 
        .S(n10187), .Z(n7789) );
  XNOR2_X1 U10074 ( .A(n7789), .B(SI_11_), .ZN(n7792) );
  INV_X1 U10075 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n7769) );
  NAND2_X1 U10076 ( .A1(n7770), .A2(n7769), .ZN(n7795) );
  NAND2_X1 U10077 ( .A1(n7795), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7771) );
  XNOR2_X1 U10078 ( .A(n7771), .B(P1_IR_REG_11__SCAN_IN), .ZN(n14107) );
  AOI22_X1 U10079 ( .A1(n8173), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n7954), 
        .B2(n14107), .ZN(n7772) );
  NAND2_X2 U10080 ( .A1(n7773), .A2(n7772), .ZN(n11571) );
  MUX2_X1 U10081 ( .A(n14034), .B(n11571), .S(n8150), .Z(n7777) );
  MUX2_X1 U10082 ( .A(n14034), .B(n11571), .S(n8176), .Z(n7774) );
  NAND2_X1 U10083 ( .A1(n7775), .A2(n7774), .ZN(n7781) );
  INV_X1 U10084 ( .A(n7776), .ZN(n7779) );
  INV_X1 U10085 ( .A(n7777), .ZN(n7778) );
  NAND2_X1 U10086 ( .A1(n7779), .A2(n7778), .ZN(n7780) );
  NAND2_X1 U10087 ( .A1(n7781), .A2(n7780), .ZN(n7801) );
  NAND2_X1 U10088 ( .A1(n7782), .A2(n11897), .ZN(n7783) );
  NAND2_X1 U10089 ( .A1(n7808), .A2(n7783), .ZN(n11899) );
  OR2_X1 U10090 ( .A1(n8119), .A2(n11899), .ZN(n7788) );
  NAND2_X1 U10091 ( .A1(n8137), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n7787) );
  INV_X1 U10092 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n7784) );
  OR2_X1 U10093 ( .A1(n8185), .A2(n7784), .ZN(n7786) );
  INV_X1 U10094 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n11484) );
  OR2_X1 U10095 ( .A1(n8205), .A2(n11484), .ZN(n7785) );
  NAND4_X1 U10096 ( .A1(n7788), .A2(n7787), .A3(n7786), .A4(n7785), .ZN(n14033) );
  INV_X1 U10097 ( .A(n7789), .ZN(n7790) );
  NAND2_X1 U10098 ( .A1(n7790), .A2(n11530), .ZN(n7791) );
  MUX2_X1 U10099 ( .A(n10169), .B(n13222), .S(n10187), .Z(n7818) );
  XNOR2_X1 U10100 ( .A(n7818), .B(SI_12_), .ZN(n7815) );
  NAND2_X1 U10101 ( .A1(n10167), .A2(n8212), .ZN(n7798) );
  NAND2_X1 U10102 ( .A1(n7796), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7821) );
  XNOR2_X1 U10103 ( .A(n7821), .B(P1_IR_REG_12__SCAN_IN), .ZN(n10126) );
  AOI22_X1 U10104 ( .A1(n8173), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n6753), 
        .B2(n10126), .ZN(n7797) );
  MUX2_X1 U10105 ( .A(n14033), .B(n11488), .S(n8176), .Z(n7802) );
  NAND2_X1 U10106 ( .A1(n7801), .A2(n7802), .ZN(n7800) );
  MUX2_X1 U10107 ( .A(n14033), .B(n11488), .S(n8150), .Z(n7799) );
  NAND2_X1 U10108 ( .A1(n7800), .A2(n7799), .ZN(n7806) );
  INV_X1 U10109 ( .A(n7801), .ZN(n7804) );
  INV_X1 U10110 ( .A(n7802), .ZN(n7803) );
  NAND2_X1 U10111 ( .A1(n7804), .A2(n7803), .ZN(n7805) );
  INV_X1 U10112 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n10312) );
  OR2_X1 U10113 ( .A1(n8036), .A2(n10312), .ZN(n7814) );
  INV_X1 U10114 ( .A(n7843), .ZN(n7810) );
  NAND2_X1 U10115 ( .A1(n7808), .A2(n7807), .ZN(n7809) );
  NAND2_X1 U10116 ( .A1(n7810), .A2(n7809), .ZN(n12026) );
  OR2_X1 U10117 ( .A1(n8119), .A2(n12026), .ZN(n7813) );
  NAND2_X1 U10118 ( .A1(n8033), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n7812) );
  NAND2_X1 U10119 ( .A1(n8032), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n7811) );
  NAND4_X1 U10120 ( .A1(n7814), .A2(n7813), .A3(n7812), .A4(n7811), .ZN(n14032) );
  NAND2_X1 U10121 ( .A1(n7818), .A2(n7817), .ZN(n7819) );
  MUX2_X1 U10122 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(P1_DATAO_REG_13__SCAN_IN), 
        .S(n10187), .Z(n7834) );
  XNOR2_X1 U10123 ( .A(n7834), .B(n11702), .ZN(n7832) );
  XNOR2_X1 U10124 ( .A(n7833), .B(n7832), .ZN(n10280) );
  NAND2_X1 U10125 ( .A1(n10280), .A2(n8212), .ZN(n7826) );
  INV_X1 U10126 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n7820) );
  NAND2_X1 U10127 ( .A1(n7821), .A2(n7820), .ZN(n7822) );
  NAND2_X1 U10128 ( .A1(n7822), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7838) );
  XNOR2_X1 U10129 ( .A(n7838), .B(n7837), .ZN(n10316) );
  OAI22_X1 U10130 ( .A1(n10316), .A2(n9667), .B1(n7823), .B2(n10283), .ZN(
        n7824) );
  INV_X1 U10131 ( .A(n7824), .ZN(n7825) );
  MUX2_X1 U10132 ( .A(n14032), .B(n11736), .S(n8150), .Z(n7828) );
  MUX2_X1 U10133 ( .A(n11898), .B(n12031), .S(n8176), .Z(n7827) );
  NAND2_X1 U10134 ( .A1(n7829), .A2(n7828), .ZN(n7830) );
  NAND2_X1 U10135 ( .A1(n7831), .A2(n7830), .ZN(n7867) );
  INV_X1 U10136 ( .A(n7834), .ZN(n7835) );
  INV_X1 U10137 ( .A(SI_14_), .ZN(n9877) );
  MUX2_X1 U10138 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(P1_DATAO_REG_14__SCAN_IN), 
        .S(n10187), .Z(n7849) );
  XNOR2_X1 U10139 ( .A(n7851), .B(n7849), .ZN(n10522) );
  NAND2_X1 U10140 ( .A1(n10522), .A2(n8212), .ZN(n7842) );
  NAND2_X1 U10141 ( .A1(n7838), .A2(n7837), .ZN(n7839) );
  NAND2_X1 U10142 ( .A1(n7839), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7840) );
  XNOR2_X1 U10143 ( .A(n7840), .B(P1_IR_REG_14__SCAN_IN), .ZN(n11172) );
  AOI22_X1 U10144 ( .A1(n11172), .A2(n6753), .B1(n8173), .B2(
        P2_DATAO_REG_14__SCAN_IN), .ZN(n7841) );
  NOR2_X1 U10145 ( .A1(n7843), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n7844) );
  OR2_X1 U10146 ( .A1(n7857), .A2(n7844), .ZN(n13890) );
  OR2_X1 U10147 ( .A1(n8119), .A2(n13890), .ZN(n7848) );
  INV_X1 U10148 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n11183) );
  OR2_X1 U10149 ( .A1(n8036), .A2(n11183), .ZN(n7847) );
  NAND2_X1 U10150 ( .A1(n8033), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n7846) );
  NAND2_X1 U10151 ( .A1(n8032), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n7845) );
  NAND4_X1 U10152 ( .A1(n7848), .A2(n7847), .A3(n7846), .A4(n7845), .ZN(n14031) );
  XNOR2_X1 U10153 ( .A(n13892), .B(n14031), .ZN(n11649) );
  INV_X1 U10154 ( .A(n7849), .ZN(n7850) );
  MUX2_X1 U10155 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(P1_DATAO_REG_15__SCAN_IN), 
        .S(n10187), .Z(n7878) );
  XNOR2_X1 U10156 ( .A(n7878), .B(SI_15_), .ZN(n7882) );
  XNOR2_X1 U10157 ( .A(n7883), .B(n7882), .ZN(n10780) );
  NAND2_X1 U10158 ( .A1(n10780), .A2(n8212), .ZN(n7856) );
  NAND2_X1 U10159 ( .A1(n7853), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7854) );
  XNOR2_X1 U10160 ( .A(n7854), .B(P1_IR_REG_15__SCAN_IN), .ZN(n11186) );
  AOI22_X1 U10161 ( .A1(n8173), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n7954), 
        .B2(n11186), .ZN(n7855) );
  NAND2_X1 U10162 ( .A1(n8137), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n7864) );
  NAND2_X1 U10163 ( .A1(n7857), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n7872) );
  OR2_X1 U10164 ( .A1(n7857), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n7858) );
  AND2_X1 U10165 ( .A1(n7872), .A2(n7858), .ZN(n14017) );
  NAND2_X1 U10166 ( .A1(n7608), .A2(n14017), .ZN(n7863) );
  INV_X1 U10167 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n7859) );
  OR2_X1 U10168 ( .A1(n8205), .A2(n7859), .ZN(n7862) );
  INV_X1 U10169 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n7860) );
  OR2_X1 U10170 ( .A1(n8201), .A2(n7860), .ZN(n7861) );
  NAND4_X1 U10171 ( .A1(n7864), .A2(n7863), .A3(n7862), .A4(n7861), .ZN(n14030) );
  INV_X1 U10172 ( .A(n14030), .ZN(n7868) );
  NAND2_X1 U10173 ( .A1(n14019), .A2(n7868), .ZN(n8234) );
  INV_X1 U10174 ( .A(n14031), .ZN(n12025) );
  NAND2_X1 U10175 ( .A1(n13892), .A2(n12025), .ZN(n7865) );
  AOI21_X1 U10176 ( .B1(n8234), .B2(n7865), .A(n8176), .ZN(n7866) );
  AOI21_X1 U10177 ( .B1(n7867), .B2(n11649), .A(n7866), .ZN(n7870) );
  OR2_X1 U10178 ( .A1(n14019), .A2(n7868), .ZN(n8235) );
  INV_X1 U10179 ( .A(n8235), .ZN(n9527) );
  OR2_X1 U10180 ( .A1(n13892), .A2(n12025), .ZN(n9525) );
  AND2_X1 U10181 ( .A1(n8235), .A2(n9525), .ZN(n7869) );
  OAI22_X1 U10182 ( .A1(n7870), .A2(n9527), .B1(n8215), .B2(n7869), .ZN(n7916)
         );
  OR2_X1 U10183 ( .A1(n8234), .A2(n8215), .ZN(n7915) );
  NAND2_X1 U10184 ( .A1(n7872), .A2(n7871), .ZN(n7873) );
  AND2_X1 U10185 ( .A1(n7893), .A2(n7873), .ZN(n13934) );
  NAND2_X1 U10186 ( .A1(n13934), .A2(n7608), .ZN(n7877) );
  NAND2_X1 U10187 ( .A1(n8137), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n7876) );
  NAND2_X1 U10188 ( .A1(n8033), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n7875) );
  NAND2_X1 U10189 ( .A1(n8032), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n7874) );
  NAND4_X1 U10190 ( .A1(n7877), .A2(n7876), .A3(n7875), .A4(n7874), .ZN(n12038) );
  INV_X1 U10191 ( .A(n7878), .ZN(n7880) );
  NAND2_X1 U10192 ( .A1(n7880), .A2(n7879), .ZN(n7881) );
  MUX2_X1 U10193 ( .A(n10976), .B(n7884), .S(n10187), .Z(n7900) );
  XNOR2_X1 U10194 ( .A(n7900), .B(SI_16_), .ZN(n7898) );
  XNOR2_X1 U10195 ( .A(n7899), .B(n7898), .ZN(n10975) );
  NAND2_X1 U10196 ( .A1(n10975), .A2(n8212), .ZN(n7891) );
  NOR2_X1 U10197 ( .A1(n7853), .A2(P1_IR_REG_15__SCAN_IN), .ZN(n7888) );
  INV_X1 U10198 ( .A(n7888), .ZN(n7885) );
  NAND2_X1 U10199 ( .A1(n7885), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7886) );
  MUX2_X1 U10200 ( .A(P1_IR_REG_31__SCAN_IN), .B(n7886), .S(
        P1_IR_REG_16__SCAN_IN), .Z(n7889) );
  NAND2_X1 U10201 ( .A1(n7888), .A2(n7887), .ZN(n7904) );
  NAND2_X1 U10202 ( .A1(n7889), .A2(n7904), .ZN(n11289) );
  INV_X1 U10203 ( .A(n11289), .ZN(n11295) );
  AOI22_X1 U10204 ( .A1(n8173), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n6753), 
        .B2(n11295), .ZN(n7890) );
  MUX2_X1 U10205 ( .A(n12038), .B(n14425), .S(n8150), .Z(n7926) );
  AND2_X1 U10206 ( .A1(n7893), .A2(n7892), .ZN(n7894) );
  OR2_X1 U10207 ( .A1(n7894), .A2(n7940), .ZN(n13947) );
  AOI22_X1 U10208 ( .A1(n8137), .A2(P1_REG1_REG_17__SCAN_IN), .B1(n8033), .B2(
        P1_REG0_REG_17__SCAN_IN), .ZN(n7897) );
  INV_X1 U10209 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n7895) );
  OR2_X1 U10210 ( .A1(n8205), .A2(n7895), .ZN(n7896) );
  NOR2_X1 U10211 ( .A1(n8176), .A2(n12038), .ZN(n7925) );
  AOI21_X1 U10212 ( .B1(n7926), .B2(n14320), .A(n7925), .ZN(n7913) );
  NAND2_X1 U10213 ( .A1(n7900), .A2(n10152), .ZN(n7901) );
  MUX2_X1 U10214 ( .A(n11123), .B(n13208), .S(n10187), .Z(n7933) );
  XNOR2_X1 U10215 ( .A(n7933), .B(SI_17_), .ZN(n7902) );
  XNOR2_X1 U10216 ( .A(n7931), .B(n7902), .ZN(n11122) );
  NAND2_X1 U10217 ( .A1(n11122), .A2(n8212), .ZN(n7907) );
  NAND2_X1 U10218 ( .A1(n7904), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7903) );
  MUX2_X1 U10219 ( .A(P1_IR_REG_31__SCAN_IN), .B(n7903), .S(
        P1_IR_REG_17__SCAN_IN), .Z(n7905) );
  AND2_X1 U10220 ( .A1(n7905), .A2(n7936), .ZN(n11296) );
  AOI22_X1 U10221 ( .A1(n8173), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n7954), 
        .B2(n11296), .ZN(n7906) );
  NAND2_X1 U10222 ( .A1(n14320), .A2(n8176), .ZN(n7919) );
  OR2_X1 U10223 ( .A1(n14425), .A2(n7919), .ZN(n7909) );
  NOR2_X1 U10224 ( .A1(n14320), .A2(n8176), .ZN(n7924) );
  INV_X1 U10225 ( .A(n12038), .ZN(n14014) );
  NAND2_X1 U10226 ( .A1(n7924), .A2(n14014), .ZN(n7908) );
  AND2_X1 U10227 ( .A1(n7909), .A2(n7908), .ZN(n7921) );
  INV_X1 U10228 ( .A(n14320), .ZN(n13984) );
  NAND2_X1 U10229 ( .A1(n7926), .A2(n13984), .ZN(n7910) );
  OR2_X1 U10230 ( .A1(n14425), .A2(n8215), .ZN(n7917) );
  NAND2_X1 U10231 ( .A1(n7910), .A2(n7917), .ZN(n7911) );
  NAND2_X1 U10232 ( .A1(n7911), .A2(n14469), .ZN(n7912) );
  OAI211_X1 U10233 ( .C1(n7913), .C2(n14469), .A(n7921), .B(n7912), .ZN(n7914)
         );
  INV_X1 U10234 ( .A(n7917), .ZN(n7918) );
  NAND2_X1 U10235 ( .A1(n7926), .A2(n7918), .ZN(n7920) );
  NAND2_X1 U10236 ( .A1(n7920), .A2(n7919), .ZN(n7923) );
  INV_X1 U10237 ( .A(n7921), .ZN(n7922) );
  AOI22_X1 U10238 ( .A1(n7923), .A2(n14469), .B1(n7926), .B2(n7922), .ZN(n7930) );
  AOI21_X1 U10239 ( .B1(n7926), .B2(n7925), .A(n7924), .ZN(n7927) );
  NAND2_X1 U10240 ( .A1(n7933), .A2(n10328), .ZN(n7932) );
  INV_X1 U10241 ( .A(n7933), .ZN(n7934) );
  NAND2_X1 U10242 ( .A1(n7934), .A2(SI_17_), .ZN(n7935) );
  MUX2_X1 U10243 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(P1_DATAO_REG_18__SCAN_IN), 
        .S(n10187), .Z(n7977) );
  XNOR2_X1 U10244 ( .A(n7946), .B(n7977), .ZN(n11377) );
  NAND2_X1 U10245 ( .A1(n11377), .A2(n8212), .ZN(n7939) );
  NAND2_X1 U10246 ( .A1(n7936), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7937) );
  XNOR2_X1 U10247 ( .A(n7937), .B(P1_IR_REG_18__SCAN_IN), .ZN(n12100) );
  AOI22_X1 U10248 ( .A1(n8173), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n6753), 
        .B2(n12100), .ZN(n7938) );
  XNOR2_X1 U10249 ( .A(n14414), .B(n8150), .ZN(n7945) );
  NAND2_X1 U10250 ( .A1(n7940), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n7957) );
  OR2_X1 U10251 ( .A1(n7940), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n7941) );
  NAND2_X1 U10252 ( .A1(n7957), .A2(n7941), .ZN(n14328) );
  AOI22_X1 U10253 ( .A1(n8137), .A2(P1_REG1_REG_18__SCAN_IN), .B1(n8032), .B2(
        P1_REG2_REG_18__SCAN_IN), .ZN(n7943) );
  NAND2_X1 U10254 ( .A1(n8033), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n7942) );
  OAI211_X1 U10255 ( .C1(n14328), .C2(n8119), .A(n7943), .B(n7942), .ZN(n14029) );
  XNOR2_X1 U10256 ( .A(n14029), .B(n8176), .ZN(n7944) );
  INV_X1 U10257 ( .A(n7946), .ZN(n7947) );
  NAND2_X1 U10258 ( .A1(n7947), .A2(n7977), .ZN(n7949) );
  NAND2_X1 U10259 ( .A1(n7984), .A2(SI_18_), .ZN(n7948) );
  NAND2_X1 U10260 ( .A1(n7949), .A2(n7948), .ZN(n7953) );
  MUX2_X1 U10261 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(P1_DATAO_REG_19__SCAN_IN), 
        .S(n10187), .Z(n7950) );
  NAND2_X1 U10262 ( .A1(n7950), .A2(SI_19_), .ZN(n7980) );
  INV_X1 U10263 ( .A(n7950), .ZN(n7951) );
  NAND2_X1 U10264 ( .A1(n7951), .A2(n12163), .ZN(n7978) );
  NAND2_X1 U10265 ( .A1(n7980), .A2(n7978), .ZN(n7952) );
  NAND2_X1 U10266 ( .A1(n8963), .A2(n8212), .ZN(n7956) );
  AOI22_X1 U10267 ( .A1(n8173), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n7954), 
        .B2(n9502), .ZN(n7955) );
  NAND2_X1 U10268 ( .A1(n7957), .A2(n12111), .ZN(n7958) );
  NAND2_X1 U10269 ( .A1(n7969), .A2(n7958), .ZN(n14308) );
  INV_X1 U10270 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n7961) );
  NAND2_X1 U10271 ( .A1(n8033), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n7960) );
  NAND2_X1 U10272 ( .A1(n8032), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n7959) );
  OAI211_X1 U10273 ( .C1(n8036), .C2(n7961), .A(n7960), .B(n7959), .ZN(n7962)
         );
  INV_X1 U10274 ( .A(n7962), .ZN(n7963) );
  NAND2_X1 U10275 ( .A1(n7964), .A2(n7963), .ZN(n14322) );
  INV_X1 U10276 ( .A(n14322), .ZN(n14286) );
  NAND2_X1 U10277 ( .A1(n14409), .A2(n14286), .ZN(n9532) );
  NAND2_X1 U10278 ( .A1(n7965), .A2(n14303), .ZN(n7968) );
  MUX2_X1 U10279 ( .A(n9532), .B(n7966), .S(n8176), .Z(n7967) );
  NAND2_X1 U10280 ( .A1(n7969), .A2(n13966), .ZN(n7970) );
  NAND2_X1 U10281 ( .A1(n7993), .A2(n7970), .ZN(n14292) );
  INV_X1 U10282 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n7973) );
  NAND2_X1 U10283 ( .A1(n8033), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n7972) );
  NAND2_X1 U10284 ( .A1(n8032), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n7971) );
  OAI211_X1 U10285 ( .C1(n8036), .C2(n7973), .A(n7972), .B(n7971), .ZN(n7974)
         );
  INV_X1 U10286 ( .A(n7974), .ZN(n7975) );
  INV_X1 U10287 ( .A(SI_18_), .ZN(n10469) );
  INV_X1 U10288 ( .A(n7977), .ZN(n7976) );
  OAI21_X1 U10289 ( .B1(n10469), .B2(n7976), .A(n7980), .ZN(n7983) );
  NOR2_X1 U10290 ( .A1(n7977), .A2(SI_18_), .ZN(n7981) );
  INV_X1 U10291 ( .A(n7978), .ZN(n7979) );
  AOI21_X1 U10292 ( .B1(n7981), .B2(n7980), .A(n7979), .ZN(n7982) );
  INV_X1 U10293 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7985) );
  MUX2_X1 U10294 ( .A(n7985), .B(n7139), .S(n10187), .Z(n7999) );
  XNOR2_X1 U10295 ( .A(n8001), .B(n7999), .ZN(n11492) );
  NAND2_X1 U10296 ( .A1(n11492), .A2(n8212), .ZN(n7987) );
  NAND2_X1 U10297 ( .A1(n8173), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n7986) );
  MUX2_X1 U10298 ( .A(n14028), .B(n14404), .S(n8150), .Z(n7990) );
  NAND2_X1 U10299 ( .A1(n7991), .A2(n7990), .ZN(n7989) );
  MUX2_X1 U10300 ( .A(n14028), .B(n14404), .S(n8176), .Z(n7988) );
  NAND2_X1 U10301 ( .A1(n7989), .A2(n7988), .ZN(n7992) );
  AND2_X1 U10302 ( .A1(n7993), .A2(n13915), .ZN(n7994) );
  OR2_X1 U10303 ( .A1(n7994), .A2(n8010), .ZN(n14272) );
  INV_X1 U10304 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n14401) );
  NAND2_X1 U10305 ( .A1(n8033), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n7996) );
  NAND2_X1 U10306 ( .A1(n8032), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n7995) );
  OAI211_X1 U10307 ( .C1(n8036), .C2(n14401), .A(n7996), .B(n7995), .ZN(n7997)
         );
  INV_X1 U10308 ( .A(n7997), .ZN(n7998) );
  INV_X1 U10309 ( .A(n7999), .ZN(n8000) );
  NAND2_X1 U10310 ( .A1(n8001), .A2(n8000), .ZN(n8004) );
  INV_X1 U10311 ( .A(SI_20_), .ZN(n10777) );
  MUX2_X1 U10312 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(P1_DATAO_REG_21__SCAN_IN), 
        .S(n10187), .Z(n8020) );
  XNOR2_X1 U10313 ( .A(n8020), .B(SI_21_), .ZN(n8017) );
  XNOR2_X1 U10314 ( .A(n8019), .B(n8017), .ZN(n11613) );
  NAND2_X1 U10315 ( .A1(n11613), .A2(n8212), .ZN(n8006) );
  NAND2_X1 U10316 ( .A1(n8173), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n8005) );
  MUX2_X1 U10317 ( .A(n14248), .B(n14271), .S(n8176), .Z(n8008) );
  MUX2_X1 U10318 ( .A(n14248), .B(n14271), .S(n8150), .Z(n8007) );
  INV_X1 U10319 ( .A(n8008), .ZN(n8009) );
  NOR2_X1 U10320 ( .A1(n8010), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n8011) );
  OR2_X1 U10321 ( .A1(n8030), .A2(n8011), .ZN(n13975) );
  INV_X1 U10322 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n8014) );
  NAND2_X1 U10323 ( .A1(n8033), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n8013) );
  NAND2_X1 U10324 ( .A1(n8032), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n8012) );
  OAI211_X1 U10325 ( .C1(n8036), .C2(n8014), .A(n8013), .B(n8012), .ZN(n8015)
         );
  INV_X1 U10326 ( .A(n8015), .ZN(n8016) );
  INV_X1 U10327 ( .A(n8017), .ZN(n8018) );
  NAND2_X1 U10328 ( .A1(n8019), .A2(n8018), .ZN(n8022) );
  NAND2_X1 U10329 ( .A1(n8020), .A2(SI_21_), .ZN(n8021) );
  NAND2_X1 U10330 ( .A1(n9018), .A2(n8621), .ZN(n8023) );
  MUX2_X1 U10331 ( .A(n14027), .B(n14394), .S(n8150), .Z(n8026) );
  NAND2_X1 U10332 ( .A1(n8027), .A2(n8026), .ZN(n8025) );
  MUX2_X1 U10333 ( .A(n14027), .B(n14394), .S(n8176), .Z(n8024) );
  NAND2_X1 U10334 ( .A1(n8025), .A2(n8024), .ZN(n8029) );
  OR2_X1 U10335 ( .A1(n8030), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n8031) );
  NAND2_X1 U10336 ( .A1(n8030), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n8046) );
  NAND2_X1 U10337 ( .A1(n8031), .A2(n8046), .ZN(n14239) );
  INV_X1 U10338 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n14390) );
  NAND2_X1 U10339 ( .A1(n8032), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n8035) );
  NAND2_X1 U10340 ( .A1(n8033), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n8034) );
  OAI211_X1 U10341 ( .C1(n8036), .C2(n14390), .A(n8035), .B(n8034), .ZN(n8037)
         );
  INV_X1 U10342 ( .A(n8037), .ZN(n8038) );
  MUX2_X1 U10343 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(P1_DATAO_REG_22__SCAN_IN), 
        .S(n10187), .Z(n8058) );
  NAND2_X1 U10344 ( .A1(n8055), .A2(SI_22_), .ZN(n8039) );
  NAND2_X1 U10345 ( .A1(n11810), .A2(n8039), .ZN(n8041) );
  MUX2_X1 U10346 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(P1_DATAO_REG_23__SCAN_IN), 
        .S(n10187), .Z(n8059) );
  XNOR2_X1 U10347 ( .A(n8059), .B(SI_23_), .ZN(n8040) );
  NAND2_X1 U10348 ( .A1(n11888), .A2(n8212), .ZN(n8043) );
  NAND2_X1 U10349 ( .A1(n8173), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n8042) );
  MUX2_X1 U10350 ( .A(n14249), .B(n14385), .S(n8176), .Z(n8045) );
  MUX2_X1 U10351 ( .A(n14249), .B(n14385), .S(n8150), .Z(n8044) );
  INV_X1 U10352 ( .A(n8046), .ZN(n8047) );
  NAND2_X1 U10353 ( .A1(n8047), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n8070) );
  OAI21_X1 U10354 ( .B1(P1_REG3_REG_24__SCAN_IN), .B2(n8047), .A(n8070), .ZN(
        n14222) );
  OR2_X1 U10355 ( .A1(n8119), .A2(n14222), .ZN(n8052) );
  NAND2_X1 U10356 ( .A1(n8137), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n8051) );
  INV_X1 U10357 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n8048) );
  OR2_X1 U10358 ( .A1(n8185), .A2(n8048), .ZN(n8050) );
  INV_X1 U10359 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n14223) );
  OR2_X1 U10360 ( .A1(n8205), .A2(n14223), .ZN(n8049) );
  NAND4_X1 U10361 ( .A1(n8052), .A2(n8051), .A3(n8050), .A4(n8049), .ZN(n14026) );
  INV_X1 U10362 ( .A(n8059), .ZN(n8053) );
  INV_X1 U10363 ( .A(SI_23_), .ZN(n11229) );
  AOI22_X1 U10364 ( .A1(n8056), .A2(n9019), .B1(n8053), .B2(n11229), .ZN(n8054) );
  OAI21_X1 U10365 ( .B1(n9019), .B2(n8056), .A(n11229), .ZN(n8060) );
  AND2_X1 U10366 ( .A1(SI_22_), .A2(SI_23_), .ZN(n8057) );
  AOI22_X1 U10367 ( .A1(n8060), .A2(n8059), .B1(n8058), .B2(n8057), .ZN(n8061)
         );
  MUX2_X1 U10368 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(P1_DATAO_REG_24__SCAN_IN), 
        .S(n10187), .Z(n8081) );
  XNOR2_X1 U10369 ( .A(n8081), .B(SI_24_), .ZN(n8078) );
  XNOR2_X1 U10370 ( .A(n8080), .B(n8078), .ZN(n11814) );
  NAND2_X1 U10371 ( .A1(n11814), .A2(n8212), .ZN(n8063) );
  NAND2_X1 U10372 ( .A1(n8173), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n8062) );
  MUX2_X1 U10373 ( .A(n14026), .B(n14377), .S(n8150), .Z(n8066) );
  NAND2_X1 U10374 ( .A1(n8067), .A2(n8066), .ZN(n8065) );
  MUX2_X1 U10375 ( .A(n14026), .B(n14377), .S(n8176), .Z(n8064) );
  NAND2_X1 U10376 ( .A1(n8065), .A2(n8064), .ZN(n8069) );
  NAND2_X1 U10377 ( .A1(P1_REG3_REG_25__SCAN_IN), .A2(n8071), .ZN(n8093) );
  OAI21_X1 U10378 ( .B1(P1_REG3_REG_25__SCAN_IN), .B2(n8071), .A(n8093), .ZN(
        n14198) );
  OR2_X1 U10379 ( .A1(n8119), .A2(n14198), .ZN(n8077) );
  NAND2_X1 U10380 ( .A1(n8137), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n8076) );
  INV_X1 U10381 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n8072) );
  OR2_X1 U10382 ( .A1(n8201), .A2(n8072), .ZN(n8075) );
  INV_X1 U10383 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n8073) );
  OR2_X1 U10384 ( .A1(n8205), .A2(n8073), .ZN(n8074) );
  NAND4_X1 U10385 ( .A1(n8077), .A2(n8076), .A3(n8075), .A4(n8074), .ZN(n14174) );
  INV_X1 U10386 ( .A(n8078), .ZN(n8079) );
  NAND2_X1 U10387 ( .A1(n8081), .A2(SI_24_), .ZN(n8082) );
  MUX2_X1 U10388 ( .A(n6678), .B(n11881), .S(n10187), .Z(n8084) );
  INV_X1 U10389 ( .A(SI_25_), .ZN(n11747) );
  NAND2_X1 U10390 ( .A1(n8084), .A2(n11747), .ZN(n8101) );
  INV_X1 U10391 ( .A(n8084), .ZN(n8085) );
  NAND2_X1 U10392 ( .A1(n8085), .A2(SI_25_), .ZN(n8086) );
  NAND2_X1 U10393 ( .A1(n8101), .A2(n8086), .ZN(n8102) );
  XNOR2_X1 U10394 ( .A(n8103), .B(n8102), .ZN(n11879) );
  NAND2_X1 U10395 ( .A1(n11879), .A2(n8212), .ZN(n8088) );
  NAND2_X1 U10396 ( .A1(n8173), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n8087) );
  MUX2_X1 U10397 ( .A(n14174), .B(n14374), .S(n8176), .Z(n8090) );
  MUX2_X1 U10398 ( .A(n14174), .B(n14374), .S(n8150), .Z(n8089) );
  INV_X1 U10399 ( .A(n8090), .ZN(n8091) );
  INV_X1 U10400 ( .A(n8093), .ZN(n8092) );
  NAND2_X1 U10401 ( .A1(n8092), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n8117) );
  INV_X1 U10402 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n13179) );
  NAND2_X1 U10403 ( .A1(n8093), .A2(n13179), .ZN(n8094) );
  NAND2_X1 U10404 ( .A1(n8117), .A2(n8094), .ZN(n14178) );
  OR2_X1 U10405 ( .A1(n8119), .A2(n14178), .ZN(n8100) );
  NAND2_X1 U10406 ( .A1(n8137), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n8099) );
  INV_X1 U10407 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n8095) );
  OR2_X1 U10408 ( .A1(n8205), .A2(n8095), .ZN(n8098) );
  INV_X1 U10409 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n8096) );
  OR2_X1 U10410 ( .A1(n8201), .A2(n8096), .ZN(n8097) );
  NAND4_X1 U10411 ( .A1(n8100), .A2(n8099), .A3(n8098), .A4(n8097), .ZN(n14147) );
  INV_X1 U10412 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n12008) );
  MUX2_X1 U10413 ( .A(n12008), .B(n9094), .S(n10187), .Z(n8124) );
  XNOR2_X1 U10414 ( .A(n8124), .B(SI_26_), .ZN(n8104) );
  XNOR2_X1 U10415 ( .A(n8125), .B(n8104), .ZN(n12007) );
  NAND2_X1 U10416 ( .A1(n12007), .A2(n8212), .ZN(n8106) );
  NAND2_X1 U10417 ( .A1(n8173), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n8105) );
  MUX2_X1 U10418 ( .A(n14147), .B(n14366), .S(n8150), .Z(n8110) );
  NAND2_X1 U10419 ( .A1(n8109), .A2(n8110), .ZN(n8108) );
  MUX2_X1 U10420 ( .A(n14147), .B(n14366), .S(n8176), .Z(n8107) );
  NAND2_X1 U10421 ( .A1(n8108), .A2(n8107), .ZN(n8114) );
  INV_X1 U10422 ( .A(n8109), .ZN(n8112) );
  INV_X1 U10423 ( .A(n8110), .ZN(n8111) );
  NAND2_X1 U10424 ( .A1(n8112), .A2(n8111), .ZN(n8113) );
  INV_X1 U10425 ( .A(n8117), .ZN(n8115) );
  NAND2_X1 U10426 ( .A1(n8115), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n8202) );
  INV_X1 U10427 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n8116) );
  NAND2_X1 U10428 ( .A1(n8117), .A2(n8116), .ZN(n8118) );
  NAND2_X1 U10429 ( .A1(n8202), .A2(n8118), .ZN(n14159) );
  OR2_X1 U10430 ( .A1(n8119), .A2(n14159), .ZN(n8123) );
  NAND2_X1 U10431 ( .A1(n8137), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n8122) );
  INV_X1 U10432 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n14446) );
  OR2_X1 U10433 ( .A1(n8201), .A2(n14446), .ZN(n8121) );
  INV_X1 U10434 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n14160) );
  OR2_X1 U10435 ( .A1(n8205), .A2(n14160), .ZN(n8120) );
  NAND2_X1 U10436 ( .A1(n8125), .A2(n11877), .ZN(n8126) );
  NAND2_X1 U10437 ( .A1(n8127), .A2(n8126), .ZN(n8147) );
  MUX2_X1 U10438 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(P1_DATAO_REG_27__SCAN_IN), 
        .S(n10187), .Z(n8144) );
  INV_X1 U10439 ( .A(n8144), .ZN(n8128) );
  XNOR2_X1 U10440 ( .A(n8128), .B(SI_27_), .ZN(n8129) );
  NAND2_X1 U10441 ( .A1(n12047), .A2(n8212), .ZN(n8131) );
  NAND2_X1 U10442 ( .A1(n8173), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n8130) );
  MUX2_X1 U10443 ( .A(n14175), .B(n14158), .S(n8176), .Z(n8134) );
  NAND2_X1 U10444 ( .A1(n8135), .A2(n8134), .ZN(n8133) );
  MUX2_X1 U10445 ( .A(n14158), .B(n14175), .S(n8176), .Z(n8132) );
  NAND2_X1 U10446 ( .A1(n8133), .A2(n8132), .ZN(n8136) );
  NAND2_X1 U10447 ( .A1(n8136), .A2(n6570), .ZN(n8152) );
  NAND2_X1 U10448 ( .A1(n8137), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n8143) );
  XNOR2_X1 U10449 ( .A(n8202), .B(P1_REG3_REG_28__SCAN_IN), .ZN(n14137) );
  NAND2_X1 U10450 ( .A1(n7608), .A2(n14137), .ZN(n8142) );
  INV_X1 U10451 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n8138) );
  OR2_X1 U10452 ( .A1(n8185), .A2(n8138), .ZN(n8141) );
  INV_X1 U10453 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n8139) );
  OR2_X1 U10454 ( .A1(n8205), .A2(n8139), .ZN(n8140) );
  NAND4_X1 U10455 ( .A1(n8143), .A2(n8142), .A3(n8141), .A4(n8140), .ZN(n14146) );
  NOR2_X1 U10456 ( .A1(n8144), .A2(SI_27_), .ZN(n8146) );
  NAND2_X1 U10457 ( .A1(n8144), .A2(SI_27_), .ZN(n8145) );
  MUX2_X1 U10458 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(P1_DATAO_REG_28__SCAN_IN), 
        .S(n10187), .Z(n8161) );
  XNOR2_X1 U10459 ( .A(n8161), .B(SI_28_), .ZN(n8159) );
  NAND2_X1 U10460 ( .A1(n12121), .A2(n8212), .ZN(n8149) );
  NAND2_X1 U10461 ( .A1(n8173), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n8148) );
  MUX2_X1 U10462 ( .A(n14146), .B(n14138), .S(n8150), .Z(n8153) );
  MUX2_X1 U10463 ( .A(n14146), .B(n14138), .S(n8176), .Z(n8151) );
  INV_X1 U10464 ( .A(n8153), .ZN(n8154) );
  NAND2_X1 U10465 ( .A1(n8137), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n8158) );
  INV_X1 U10466 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n8155) );
  OR2_X1 U10467 ( .A1(n8205), .A2(n8155), .ZN(n8157) );
  INV_X1 U10468 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n14435) );
  OR2_X1 U10469 ( .A1(n8185), .A2(n14435), .ZN(n8156) );
  AND3_X1 U10470 ( .A1(n8158), .A2(n8157), .A3(n8156), .ZN(n8219) );
  INV_X1 U10471 ( .A(n8219), .ZN(n14024) );
  INV_X1 U10472 ( .A(n8161), .ZN(n8162) );
  NAND2_X1 U10473 ( .A1(n8162), .A2(n13329), .ZN(n8163) );
  MUX2_X1 U10474 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(P1_DATAO_REG_29__SCAN_IN), 
        .S(n10187), .Z(n8164) );
  INV_X1 U10475 ( .A(SI_29_), .ZN(n13215) );
  XNOR2_X1 U10476 ( .A(n8164), .B(n13215), .ZN(n8210) );
  NOR2_X1 U10477 ( .A1(n8164), .A2(SI_29_), .ZN(n8165) );
  AOI21_X2 U10478 ( .B1(n8211), .B2(n8210), .A(n8165), .ZN(n8188) );
  INV_X1 U10479 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n12627) );
  INV_X1 U10480 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n13866) );
  MUX2_X1 U10481 ( .A(n12627), .B(n13866), .S(n10187), .Z(n8166) );
  XNOR2_X1 U10482 ( .A(n8166), .B(SI_30_), .ZN(n8189) );
  NAND2_X1 U10483 ( .A1(n8188), .A2(n8189), .ZN(n8169) );
  INV_X1 U10484 ( .A(n8166), .ZN(n8167) );
  NAND2_X1 U10485 ( .A1(n8167), .A2(SI_30_), .ZN(n8168) );
  NAND2_X1 U10486 ( .A1(n8169), .A2(n8168), .ZN(n8172) );
  MUX2_X1 U10487 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n10187), .Z(n8170) );
  XNOR2_X1 U10488 ( .A(n8170), .B(SI_31_), .ZN(n8171) );
  NAND2_X1 U10489 ( .A1(n13861), .A2(n8212), .ZN(n8175) );
  NAND2_X1 U10490 ( .A1(n8173), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n8174) );
  MUX2_X1 U10491 ( .A(n14024), .B(n14118), .S(n8176), .Z(n8178) );
  NOR2_X1 U10492 ( .A1(n14118), .A2(n14024), .ZN(n8177) );
  OR2_X1 U10493 ( .A1(n8178), .A2(n8177), .ZN(n8259) );
  AND2_X1 U10494 ( .A1(n9915), .A2(n11493), .ZN(n8180) );
  NAND2_X1 U10495 ( .A1(n9264), .A2(n9502), .ZN(n10618) );
  OAI21_X1 U10496 ( .B1(n9666), .B2(n8180), .A(n10618), .ZN(n8261) );
  NAND2_X1 U10497 ( .A1(n11614), .A2(n8181), .ZN(n9454) );
  AND2_X1 U10498 ( .A1(n8261), .A2(n9454), .ZN(n8257) );
  NAND2_X1 U10499 ( .A1(n8259), .A2(n8257), .ZN(n8270) );
  INV_X1 U10500 ( .A(n8182), .ZN(n8186) );
  INV_X1 U10501 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n14441) );
  INV_X1 U10502 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n14125) );
  OR2_X1 U10503 ( .A1(n8205), .A2(n14125), .ZN(n8184) );
  NAND2_X1 U10504 ( .A1(n8137), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n8183) );
  OAI211_X1 U10505 ( .C1(n8185), .C2(n14441), .A(n8184), .B(n8183), .ZN(n14025) );
  OAI21_X1 U10506 ( .B1(n8186), .B2(n14024), .A(n14025), .ZN(n8187) );
  INV_X1 U10507 ( .A(n8187), .ZN(n8193) );
  INV_X1 U10508 ( .A(n8188), .ZN(n8190) );
  NAND2_X1 U10509 ( .A1(n12626), .A2(n8212), .ZN(n8192) );
  NAND2_X1 U10510 ( .A1(n8173), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n8191) );
  MUX2_X1 U10511 ( .A(n8193), .B(n14438), .S(n8215), .Z(n8223) );
  INV_X1 U10512 ( .A(n8223), .ZN(n8199) );
  NAND2_X1 U10513 ( .A1(n8215), .A2(n14024), .ZN(n8196) );
  INV_X1 U10514 ( .A(n14025), .ZN(n8194) );
  AOI21_X1 U10515 ( .B1(n8196), .B2(n8195), .A(n8194), .ZN(n8197) );
  AOI21_X1 U10516 ( .B1(n14438), .B2(n8176), .A(n8197), .ZN(n8222) );
  INV_X1 U10517 ( .A(n8222), .ZN(n8198) );
  AND2_X1 U10518 ( .A1(n8199), .A2(n8198), .ZN(n8266) );
  OR2_X1 U10519 ( .A1(n8270), .A2(n8266), .ZN(n8256) );
  INV_X1 U10520 ( .A(n8256), .ZN(n8217) );
  NAND2_X1 U10521 ( .A1(n8137), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n8209) );
  INV_X1 U10522 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n9560) );
  OR2_X1 U10523 ( .A1(n8201), .A2(n9560), .ZN(n8208) );
  INV_X1 U10524 ( .A(n8202), .ZN(n8203) );
  NAND2_X1 U10525 ( .A1(n8203), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n12551) );
  OR2_X1 U10526 ( .A1(n8119), .A2(n12551), .ZN(n8207) );
  INV_X1 U10527 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n8204) );
  OR2_X1 U10528 ( .A1(n8205), .A2(n8204), .ZN(n8206) );
  XNOR2_X1 U10529 ( .A(n8211), .B(n8210), .ZN(n13869) );
  NAND2_X1 U10530 ( .A1(n13869), .A2(n8212), .ZN(n8214) );
  NAND2_X1 U10531 ( .A1(n8173), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n8213) );
  INV_X1 U10532 ( .A(n12555), .ZN(n9565) );
  MUX2_X1 U10533 ( .A(n12074), .B(n9565), .S(n8215), .Z(n8225) );
  INV_X1 U10534 ( .A(n12074), .ZN(n14131) );
  MUX2_X1 U10535 ( .A(n14131), .B(n12555), .S(n8176), .Z(n8224) );
  NAND2_X1 U10536 ( .A1(n8225), .A2(n8224), .ZN(n8263) );
  XNOR2_X1 U10537 ( .A(n14118), .B(n8219), .ZN(n8258) );
  INV_X1 U10538 ( .A(n8258), .ZN(n8221) );
  INV_X1 U10539 ( .A(n8261), .ZN(n8220) );
  NAND2_X1 U10540 ( .A1(n8221), .A2(n8220), .ZN(n8268) );
  AND2_X1 U10541 ( .A1(n8223), .A2(n8222), .ZN(n8265) );
  OR2_X1 U10542 ( .A1(n8268), .A2(n8265), .ZN(n8264) );
  INV_X1 U10543 ( .A(n8264), .ZN(n8228) );
  INV_X1 U10544 ( .A(n8224), .ZN(n8227) );
  INV_X1 U10545 ( .A(n8225), .ZN(n8226) );
  NAND2_X1 U10546 ( .A1(n8227), .A2(n8226), .ZN(n8255) );
  NAND3_X1 U10547 ( .A1(n8229), .A2(n8228), .A3(n8255), .ZN(n8274) );
  XNOR2_X1 U10548 ( .A(n12555), .B(n12074), .ZN(n9543) );
  INV_X1 U10549 ( .A(n14146), .ZN(n13878) );
  INV_X1 U10550 ( .A(n14175), .ZN(n9465) );
  NAND2_X1 U10551 ( .A1(n14158), .A2(n9465), .ZN(n9541) );
  OR2_X1 U10552 ( .A1(n14158), .A2(n9465), .ZN(n8230) );
  NAND2_X1 U10553 ( .A1(n9541), .A2(n8230), .ZN(n14144) );
  INV_X1 U10554 ( .A(n14144), .ZN(n14150) );
  INV_X1 U10555 ( .A(n14147), .ZN(n8231) );
  XNOR2_X1 U10556 ( .A(n14366), .B(n8231), .ZN(n14171) );
  NAND2_X1 U10557 ( .A1(n14374), .A2(n14213), .ZN(n14170) );
  OR2_X1 U10558 ( .A1(n14374), .A2(n14213), .ZN(n8232) );
  NAND2_X1 U10559 ( .A1(n14170), .A2(n8232), .ZN(n14192) );
  XNOR2_X1 U10560 ( .A(n14377), .B(n14026), .ZN(n14205) );
  INV_X1 U10561 ( .A(n14027), .ZN(n14265) );
  XNOR2_X1 U10562 ( .A(n14271), .B(n14248), .ZN(n14266) );
  OR2_X1 U10563 ( .A1(n13949), .A2(n13984), .ZN(n9529) );
  NAND2_X1 U10564 ( .A1(n13949), .A2(n13984), .ZN(n8233) );
  NAND2_X1 U10565 ( .A1(n9529), .A2(n8233), .ZN(n12042) );
  XNOR2_X1 U10566 ( .A(n11736), .B(n11898), .ZN(n11599) );
  XNOR2_X1 U10567 ( .A(n11488), .B(n11824), .ZN(n11477) );
  INV_X1 U10568 ( .A(n14034), .ZN(n11352) );
  XNOR2_X1 U10569 ( .A(n11663), .B(n11418), .ZN(n11360) );
  XNOR2_X1 U10570 ( .A(n11767), .B(n11465), .ZN(n11161) );
  INV_X1 U10571 ( .A(n14037), .ZN(n9515) );
  XNOR2_X1 U10572 ( .A(n11471), .B(n9515), .ZN(n11231) );
  INV_X1 U10573 ( .A(n14039), .ZN(n10662) );
  XNOR2_X1 U10574 ( .A(n14002), .B(n10662), .ZN(n10645) );
  INV_X1 U10575 ( .A(n10645), .ZN(n8241) );
  NAND2_X1 U10576 ( .A1(n10900), .A2(n10837), .ZN(n9507) );
  NAND2_X1 U10577 ( .A1(n14839), .A2(n14041), .ZN(n8236) );
  NAND2_X1 U10578 ( .A1(n8237), .A2(n9505), .ZN(n10620) );
  INV_X1 U10579 ( .A(n10171), .ZN(n10178) );
  AND4_X1 U10580 ( .A1(n10611), .A2(n10178), .A3(n10509), .A4(n10822), .ZN(
        n8240) );
  INV_X1 U10581 ( .A(n14040), .ZN(n9508) );
  XNOR2_X1 U10582 ( .A(n10897), .B(n9508), .ZN(n10656) );
  INV_X1 U10583 ( .A(n10656), .ZN(n10660) );
  NAND4_X1 U10584 ( .A1(n8241), .A2(n10828), .A3(n8240), .A4(n10660), .ZN(
        n8242) );
  XNOR2_X1 U10585 ( .A(n11200), .B(n11241), .ZN(n11148) );
  OR4_X1 U10586 ( .A1(n11161), .A2(n11231), .A3(n8242), .A4(n11148), .ZN(n8243) );
  OR4_X1 U10587 ( .A1(n11477), .A2(n11413), .A3(n11360), .A4(n8243), .ZN(n8244) );
  NOR2_X1 U10588 ( .A1(n11599), .A2(n8244), .ZN(n8245) );
  NAND3_X1 U10589 ( .A1(n11771), .A2(n8245), .A3(n11649), .ZN(n8246) );
  NOR2_X1 U10590 ( .A1(n12042), .A2(n8246), .ZN(n8247) );
  XNOR2_X1 U10591 ( .A(n14425), .B(n14014), .ZN(n11838) );
  INV_X1 U10592 ( .A(n11838), .ZN(n11832) );
  XNOR2_X1 U10593 ( .A(n14404), .B(n14028), .ZN(n14280) );
  NAND3_X1 U10594 ( .A1(n14266), .A2(n8248), .A3(n14280), .ZN(n8249) );
  NOR2_X1 U10595 ( .A1(n14171), .A2(n8250), .ZN(n8251) );
  XNOR2_X1 U10596 ( .A(n8253), .B(n9502), .ZN(n8254) );
  NAND2_X1 U10597 ( .A1(n8258), .A2(n8257), .ZN(n8260) );
  MUX2_X1 U10598 ( .A(n8261), .B(n8260), .S(n8259), .Z(n8262) );
  OAI21_X1 U10599 ( .B1(n8264), .B2(n8263), .A(n8262), .ZN(n8272) );
  INV_X1 U10600 ( .A(n8265), .ZN(n8269) );
  INV_X1 U10601 ( .A(n8266), .ZN(n8267) );
  OAI22_X1 U10602 ( .A1(n8270), .A2(n8269), .B1(n8268), .B2(n8267), .ZN(n8271)
         );
  NAND2_X1 U10603 ( .A1(n8280), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8277) );
  INV_X1 U10604 ( .A(n9665), .ZN(n8278) );
  NAND2_X1 U10605 ( .A1(n6589), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8286) );
  MUX2_X1 U10606 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8286), .S(
        P1_IR_REG_25__SCAN_IN), .Z(n8288) );
  NOR2_X1 U10607 ( .A1(n12009), .A2(n11882), .ZN(n8289) );
  NAND2_X1 U10608 ( .A1(n11493), .A2(n12108), .ZN(n9449) );
  NAND2_X1 U10609 ( .A1(n9666), .A2(n9449), .ZN(n9460) );
  INV_X1 U10610 ( .A(n14059), .ZN(n9745) );
  INV_X1 U10611 ( .A(n8291), .ZN(n9747) );
  NAND3_X1 U10612 ( .A1(n10593), .A2(n9745), .A3(n14319), .ZN(n8292) );
  OAI211_X1 U10613 ( .C1(n14483), .C2(n11885), .A(n8292), .B(P1_B_REG_SCAN_IN), 
        .ZN(n8293) );
  NAND2_X1 U10614 ( .A1(n8294), .A2(n8293), .ZN(P1_U3242) );
  NOR2_X1 U10615 ( .A1(P3_IR_REG_7__SCAN_IN), .A2(P3_IR_REG_8__SCAN_IN), .ZN(
        n8295) );
  INV_X1 U10616 ( .A(P3_IR_REG_9__SCAN_IN), .ZN(n8301) );
  INV_X1 U10617 ( .A(P3_IR_REG_14__SCAN_IN), .ZN(n8300) );
  INV_X1 U10618 ( .A(P3_IR_REG_13__SCAN_IN), .ZN(n8299) );
  NAND2_X1 U10619 ( .A1(n8505), .A2(n8507), .ZN(n8501) );
  INV_X1 U10620 ( .A(n9808), .ZN(n8316) );
  NOR2_X1 U10621 ( .A1(P3_IR_REG_22__SCAN_IN), .A2(P3_IR_REG_21__SCAN_IN), 
        .ZN(n8309) );
  NOR2_X1 U10622 ( .A1(P3_IR_REG_24__SCAN_IN), .A2(P3_IR_REG_20__SCAN_IN), 
        .ZN(n8308) );
  NAND4_X1 U10623 ( .A1(n8309), .A2(n8308), .A3(n8317), .A4(n13121), .ZN(n8310) );
  NOR2_X1 U10624 ( .A1(n8313), .A2(n8453), .ZN(n8312) );
  MUX2_X1 U10625 ( .A(n8453), .B(n8312), .S(P3_IR_REG_26__SCAN_IN), .Z(n8314)
         );
  INV_X1 U10626 ( .A(n11878), .ZN(n8315) );
  INV_X1 U10627 ( .A(n11748), .ZN(n8319) );
  NAND2_X1 U10628 ( .A1(n8504), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8321) );
  MUX2_X1 U10629 ( .A(n8321), .B(P3_IR_REG_31__SCAN_IN), .S(n13121), .Z(n8323)
         );
  NAND2_X1 U10630 ( .A1(n8326), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8327) );
  NAND2_X1 U10631 ( .A1(n8324), .A2(n8453), .ZN(n8328) );
  MUX2_X1 U10632 ( .A(P3_REG2_REG_17__SCAN_IN), .B(P3_REG1_REG_17__SCAN_IN), 
        .S(n6489), .Z(n8452) );
  NOR2_X1 U10633 ( .A1(n8424), .A2(P3_IR_REG_9__SCAN_IN), .ZN(n8431) );
  NAND2_X1 U10634 ( .A1(n8431), .A2(n8330), .ZN(n8434) );
  NOR2_X1 U10635 ( .A1(n8339), .A2(P3_IR_REG_12__SCAN_IN), .ZN(n8337) );
  INV_X1 U10636 ( .A(P3_IR_REG_14__SCAN_IN), .ZN(n8331) );
  NAND2_X1 U10637 ( .A1(n8333), .A2(n8331), .ZN(n8446) );
  OAI21_X1 U10638 ( .B1(n8449), .B2(P3_IR_REG_16__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8332) );
  XNOR2_X1 U10639 ( .A(n8332), .B(P3_IR_REG_17__SCAN_IN), .ZN(n12802) );
  INV_X1 U10640 ( .A(n12802), .ZN(n10327) );
  NOR2_X1 U10641 ( .A1(n8333), .A2(n8453), .ZN(n8334) );
  MUX2_X1 U10642 ( .A(n8453), .B(n8334), .S(P3_IR_REG_14__SCAN_IN), .Z(n8336)
         );
  INV_X1 U10643 ( .A(n8446), .ZN(n8335) );
  MUX2_X1 U10644 ( .A(P3_REG2_REG_14__SCAN_IN), .B(P3_REG1_REG_14__SCAN_IN), 
        .S(n6490), .Z(n8445) );
  MUX2_X1 U10645 ( .A(P3_REG2_REG_13__SCAN_IN), .B(P3_REG1_REG_13__SCAN_IN), 
        .S(n6490), .Z(n8444) );
  OR2_X1 U10646 ( .A1(n8337), .A2(n8453), .ZN(n8338) );
  XNOR2_X1 U10647 ( .A(n8338), .B(P3_IR_REG_13__SCAN_IN), .ZN(n8540) );
  INV_X1 U10648 ( .A(n8540), .ZN(n12764) );
  MUX2_X1 U10649 ( .A(P3_REG2_REG_12__SCAN_IN), .B(P3_REG1_REG_12__SCAN_IN), 
        .S(n6489), .Z(n8443) );
  NAND2_X1 U10650 ( .A1(n8339), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8341) );
  INV_X1 U10651 ( .A(P3_IR_REG_12__SCAN_IN), .ZN(n8340) );
  MUX2_X1 U10652 ( .A(P3_REG2_REG_11__SCAN_IN), .B(P3_REG1_REG_11__SCAN_IN), 
        .S(n6490), .Z(n8442) );
  NAND2_X1 U10653 ( .A1(n8434), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8342) );
  XNOR2_X1 U10654 ( .A(n8342), .B(P3_IR_REG_11__SCAN_IN), .ZN(n8537) );
  INV_X1 U10655 ( .A(n8537), .ZN(n11529) );
  INV_X1 U10656 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n8344) );
  INV_X1 U10657 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n8343) );
  NAND2_X1 U10658 ( .A1(n8347), .A2(n8519), .ZN(n10422) );
  INV_X1 U10659 ( .A(n8347), .ZN(n8348) );
  INV_X1 U10660 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n15105) );
  NOR2_X1 U10661 ( .A1(n8350), .A2(n15105), .ZN(n15103) );
  NAND2_X1 U10662 ( .A1(n10423), .A2(n10422), .ZN(n8361) );
  INV_X1 U10663 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n8352) );
  INV_X1 U10664 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n8351) );
  MUX2_X1 U10665 ( .A(n8352), .B(n8351), .S(n6490), .Z(n8356) );
  INV_X1 U10666 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n8354) );
  INV_X1 U10667 ( .A(n8357), .ZN(n10450) );
  NAND2_X1 U10668 ( .A1(n8356), .A2(n10450), .ZN(n10430) );
  INV_X1 U10669 ( .A(n8356), .ZN(n8358) );
  NAND2_X1 U10670 ( .A1(n8358), .A2(n6496), .ZN(n8359) );
  NAND2_X1 U10671 ( .A1(n10430), .A2(n8359), .ZN(n10421) );
  INV_X1 U10672 ( .A(n10421), .ZN(n8360) );
  NAND2_X1 U10673 ( .A1(n8361), .A2(n8360), .ZN(n10431) );
  NAND2_X1 U10674 ( .A1(n10431), .A2(n10430), .ZN(n8370) );
  INV_X1 U10675 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n11013) );
  INV_X1 U10676 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n8362) );
  MUX2_X1 U10677 ( .A(n11013), .B(n8362), .S(n6490), .Z(n8366) );
  INV_X1 U10678 ( .A(P3_IR_REG_3__SCAN_IN), .ZN(n8365) );
  OR3_X1 U10679 ( .A1(P3_IR_REG_2__SCAN_IN), .A2(P3_IR_REG_1__SCAN_IN), .A3(
        P3_IR_REG_0__SCAN_IN), .ZN(n8363) );
  NAND2_X1 U10680 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(n8363), .ZN(n8364) );
  XNOR2_X1 U10681 ( .A(n8365), .B(n8364), .ZN(n9606) );
  INV_X1 U10682 ( .A(n9606), .ZN(n10549) );
  NAND2_X1 U10683 ( .A1(n8366), .A2(n10549), .ZN(n15117) );
  INV_X1 U10684 ( .A(n8366), .ZN(n8367) );
  NAND2_X1 U10685 ( .A1(n8367), .A2(n9606), .ZN(n8368) );
  NAND2_X1 U10686 ( .A1(n15117), .A2(n8368), .ZN(n10429) );
  INV_X1 U10687 ( .A(n10429), .ZN(n8369) );
  NAND2_X1 U10688 ( .A1(n8370), .A2(n8369), .ZN(n15118) );
  NAND2_X1 U10689 ( .A1(n15118), .A2(n15117), .ZN(n8380) );
  INV_X1 U10690 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n8371) );
  INV_X1 U10691 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n8471) );
  MUX2_X1 U10692 ( .A(n8371), .B(n8471), .S(n6489), .Z(n8376) );
  NAND2_X1 U10693 ( .A1(n8373), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8375) );
  INV_X1 U10694 ( .A(P3_IR_REG_4__SCAN_IN), .ZN(n8374) );
  XNOR2_X1 U10695 ( .A(n8375), .B(n8374), .ZN(n9597) );
  INV_X1 U10696 ( .A(n9597), .ZN(n15122) );
  NAND2_X1 U10697 ( .A1(n8376), .A2(n15122), .ZN(n15129) );
  INV_X1 U10698 ( .A(n8376), .ZN(n8377) );
  NAND2_X1 U10699 ( .A1(n8377), .A2(n9597), .ZN(n8378) );
  NAND2_X1 U10700 ( .A1(n15129), .A2(n8378), .ZN(n15116) );
  INV_X1 U10701 ( .A(n15116), .ZN(n8379) );
  NAND2_X1 U10702 ( .A1(n8380), .A2(n8379), .ZN(n15130) );
  NAND2_X1 U10703 ( .A1(n15130), .A2(n15129), .ZN(n8391) );
  INV_X1 U10704 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n8382) );
  INV_X1 U10705 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n8381) );
  MUX2_X1 U10706 ( .A(n8382), .B(n8381), .S(n6489), .Z(n8387) );
  NOR2_X1 U10707 ( .A1(n8373), .A2(P3_IR_REG_4__SCAN_IN), .ZN(n8385) );
  OR2_X1 U10708 ( .A1(n8385), .A2(n8453), .ZN(n8383) );
  MUX2_X1 U10709 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8383), .S(
        P3_IR_REG_5__SCAN_IN), .Z(n8386) );
  INV_X1 U10710 ( .A(P3_IR_REG_5__SCAN_IN), .ZN(n8384) );
  NAND2_X1 U10711 ( .A1(n8385), .A2(n8384), .ZN(n8393) );
  NAND2_X1 U10712 ( .A1(n8386), .A2(n8393), .ZN(n15138) );
  INV_X1 U10713 ( .A(n15138), .ZN(n10923) );
  NAND2_X1 U10714 ( .A1(n8387), .A2(n10923), .ZN(n10407) );
  INV_X1 U10715 ( .A(n8387), .ZN(n8388) );
  NAND2_X1 U10716 ( .A1(n8388), .A2(n15138), .ZN(n8389) );
  NAND2_X1 U10717 ( .A1(n10407), .A2(n8389), .ZN(n15128) );
  INV_X1 U10718 ( .A(n15128), .ZN(n8390) );
  NAND2_X1 U10719 ( .A1(n8391), .A2(n8390), .ZN(n15133) );
  NAND2_X1 U10720 ( .A1(n15133), .A2(n10407), .ZN(n8400) );
  INV_X1 U10721 ( .A(P3_REG2_REG_6__SCAN_IN), .ZN(n8527) );
  INV_X1 U10722 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n8474) );
  MUX2_X1 U10723 ( .A(n8527), .B(n8474), .S(n6489), .Z(n8396) );
  NAND2_X1 U10724 ( .A1(n8393), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8392) );
  MUX2_X1 U10725 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8392), .S(
        P3_IR_REG_6__SCAN_IN), .Z(n8395) );
  INV_X1 U10726 ( .A(n8393), .ZN(n8394) );
  NAND2_X1 U10727 ( .A1(n8394), .A2(n8406), .ZN(n8403) );
  NAND2_X1 U10728 ( .A1(n8396), .A2(n8528), .ZN(n15149) );
  INV_X1 U10729 ( .A(n8396), .ZN(n8397) );
  NAND2_X1 U10730 ( .A1(n8397), .A2(n11074), .ZN(n8398) );
  NAND2_X1 U10731 ( .A1(n15149), .A2(n8398), .ZN(n10406) );
  INV_X1 U10732 ( .A(n10406), .ZN(n8399) );
  NAND2_X1 U10733 ( .A1(n8400), .A2(n8399), .ZN(n15150) );
  INV_X1 U10734 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n8402) );
  INV_X1 U10735 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n8401) );
  MUX2_X1 U10736 ( .A(n8402), .B(n8401), .S(n6490), .Z(n8410) );
  NAND2_X1 U10737 ( .A1(n8403), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8404) );
  MUX2_X1 U10738 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8404), .S(
        P3_IR_REG_7__SCAN_IN), .Z(n8409) );
  INV_X1 U10739 ( .A(P3_IR_REG_7__SCAN_IN), .ZN(n8405) );
  NAND3_X1 U10740 ( .A1(n8407), .A2(n8406), .A3(n8405), .ZN(n8408) );
  OR2_X1 U10741 ( .A1(n8373), .A2(n8408), .ZN(n8414) );
  NAND2_X1 U10742 ( .A1(n8410), .A2(n15154), .ZN(n10529) );
  INV_X1 U10743 ( .A(n8410), .ZN(n8411) );
  NAND2_X1 U10744 ( .A1(n8411), .A2(n9618), .ZN(n8412) );
  NAND2_X1 U10745 ( .A1(n10529), .A2(n8412), .ZN(n15148) );
  AOI21_X1 U10746 ( .B1(n15150), .B2(n15149), .A(n15148), .ZN(n15152) );
  INV_X1 U10747 ( .A(n10529), .ZN(n8422) );
  INV_X1 U10748 ( .A(P3_REG2_REG_8__SCAN_IN), .ZN(n8413) );
  INV_X1 U10749 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n15276) );
  MUX2_X1 U10750 ( .A(n8413), .B(n15276), .S(n6489), .Z(n8418) );
  NAND2_X1 U10751 ( .A1(n8414), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8415) );
  MUX2_X1 U10752 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8415), .S(
        P3_IR_REG_8__SCAN_IN), .Z(n8416) );
  NAND2_X1 U10753 ( .A1(n8416), .A2(n8424), .ZN(n11206) );
  INV_X1 U10754 ( .A(n11206), .ZN(n8417) );
  NAND2_X1 U10755 ( .A1(n8418), .A2(n8417), .ZN(n10855) );
  INV_X1 U10756 ( .A(n8418), .ZN(n8419) );
  NAND2_X1 U10757 ( .A1(n8419), .A2(n11206), .ZN(n8420) );
  NAND2_X1 U10758 ( .A1(n10855), .A2(n8420), .ZN(n10530) );
  INV_X1 U10759 ( .A(n10530), .ZN(n8421) );
  INV_X1 U10760 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n11326) );
  INV_X1 U10761 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n8423) );
  MUX2_X1 U10762 ( .A(n11326), .B(n8423), .S(n6490), .Z(n8426) );
  NAND2_X1 U10763 ( .A1(n8424), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8425) );
  XNOR2_X1 U10764 ( .A(n8425), .B(P3_IR_REG_9__SCAN_IN), .ZN(n11306) );
  NAND2_X1 U10765 ( .A1(n8426), .A2(n11306), .ZN(n11452) );
  INV_X1 U10766 ( .A(n8426), .ZN(n8427) );
  INV_X1 U10767 ( .A(n11306), .ZN(n10860) );
  NAND2_X1 U10768 ( .A1(n8427), .A2(n10860), .ZN(n8428) );
  NAND2_X1 U10769 ( .A1(n11452), .A2(n8428), .ZN(n10854) );
  INV_X1 U10770 ( .A(n11452), .ZN(n8440) );
  INV_X1 U10771 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n8430) );
  INV_X1 U10772 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n8429) );
  MUX2_X1 U10773 ( .A(n8430), .B(n8429), .S(n6489), .Z(n8436) );
  NOR2_X1 U10774 ( .A1(n8431), .A2(n8453), .ZN(n8432) );
  MUX2_X1 U10775 ( .A(n8453), .B(n8432), .S(P3_IR_REG_10__SCAN_IN), .Z(n8433)
         );
  INV_X1 U10776 ( .A(n8433), .ZN(n8435) );
  NAND2_X1 U10777 ( .A1(n8435), .A2(n8434), .ZN(n11393) );
  INV_X1 U10778 ( .A(n11393), .ZN(n11458) );
  NAND2_X1 U10779 ( .A1(n8436), .A2(n11458), .ZN(n8441) );
  INV_X1 U10780 ( .A(n8436), .ZN(n8437) );
  NAND2_X1 U10781 ( .A1(n8437), .A2(n11393), .ZN(n8438) );
  NAND2_X1 U10782 ( .A1(n8441), .A2(n8438), .ZN(n11451) );
  INV_X1 U10783 ( .A(n11451), .ZN(n8439) );
  NAND2_X1 U10784 ( .A1(n11455), .A2(n8441), .ZN(n11430) );
  XNOR2_X1 U10785 ( .A(n8442), .B(n8537), .ZN(n11429) );
  NAND2_X1 U10786 ( .A1(n11430), .A2(n11429), .ZN(n11428) );
  OAI21_X1 U10787 ( .B1(n8442), .B2(n11529), .A(n11428), .ZN(n11513) );
  XNOR2_X1 U10788 ( .A(n8443), .B(n11516), .ZN(n11514) );
  XNOR2_X1 U10789 ( .A(n8444), .B(n8540), .ZN(n12760) );
  XNOR2_X1 U10790 ( .A(n12783), .B(P3_REG1_REG_14__SCAN_IN), .ZN(n12776) );
  XNOR2_X1 U10791 ( .A(n12783), .B(P3_REG2_REG_14__SCAN_IN), .ZN(n12774) );
  MUX2_X1 U10792 ( .A(n12776), .B(n12774), .S(n8552), .Z(n12779) );
  NAND2_X1 U10793 ( .A1(n8446), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8447) );
  XNOR2_X1 U10794 ( .A(n8447), .B(P3_IR_REG_15__SCAN_IN), .ZN(n14623) );
  MUX2_X1 U10795 ( .A(P3_REG2_REG_15__SCAN_IN), .B(P3_REG1_REG_15__SCAN_IN), 
        .S(n6489), .Z(n14630) );
  AOI21_X1 U10796 ( .B1(n8448), .B2(n14623), .A(n14628), .ZN(n14645) );
  INV_X1 U10797 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n8545) );
  INV_X1 U10798 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n8492) );
  MUX2_X1 U10799 ( .A(n8545), .B(n8492), .S(n6490), .Z(n8451) );
  NAND2_X1 U10800 ( .A1(n8449), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8450) );
  XNOR2_X1 U10801 ( .A(n8450), .B(P3_IR_REG_16__SCAN_IN), .ZN(n14646) );
  NOR2_X1 U10802 ( .A1(n8451), .A2(n14646), .ZN(n14641) );
  NAND2_X1 U10803 ( .A1(n8451), .A2(n14646), .ZN(n14642) );
  XOR2_X1 U10804 ( .A(n8452), .B(n12802), .Z(n12799) );
  OR2_X1 U10805 ( .A1(n8454), .A2(n8453), .ZN(n8455) );
  XNOR2_X1 U10806 ( .A(n8455), .B(P3_IR_REG_18__SCAN_IN), .ZN(n12820) );
  XNOR2_X1 U10807 ( .A(n8456), .B(n12820), .ZN(n12806) );
  MUX2_X1 U10808 ( .A(P3_REG2_REG_18__SCAN_IN), .B(P3_REG1_REG_18__SCAN_IN), 
        .S(n6490), .Z(n12807) );
  NAND2_X1 U10809 ( .A1(n8458), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8460) );
  XNOR2_X1 U10810 ( .A(n12345), .B(P3_REG2_REG_19__SCAN_IN), .ZN(n8551) );
  XNOR2_X1 U10811 ( .A(n12345), .B(P3_REG1_REG_19__SCAN_IN), .ZN(n8497) );
  MUX2_X1 U10812 ( .A(n8551), .B(n8497), .S(n6489), .Z(n8461) );
  XNOR2_X1 U10813 ( .A(n8462), .B(n8461), .ZN(n8517) );
  NAND2_X1 U10814 ( .A1(n9918), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8464) );
  INV_X1 U10815 ( .A(n14646), .ZN(n10153) );
  INV_X1 U10816 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n13182) );
  NOR3_X1 U10817 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), .A3(
        n13182), .ZN(n8467) );
  NOR2_X1 U10818 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(n13182), .ZN(n8466) );
  INV_X1 U10819 ( .A(n8467), .ZN(n8465) );
  NOR2_X1 U10820 ( .A1(n8343), .A2(n10160), .ZN(n10159) );
  NOR2_X1 U10821 ( .A1(n8467), .A2(n10159), .ZN(n10415) );
  AND2_X1 U10822 ( .A1(n6496), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n8468) );
  NOR2_X1 U10823 ( .A1(n10549), .A2(n8469), .ZN(n8470) );
  MUX2_X1 U10824 ( .A(n8471), .B(P3_REG1_REG_4__SCAN_IN), .S(n9597), .Z(n15113) );
  NOR2_X1 U10825 ( .A1(n10923), .A2(n8472), .ZN(n8473) );
  AOI22_X1 U10826 ( .A1(n8528), .A2(P3_REG1_REG_6__SCAN_IN), .B1(n8474), .B2(
        n11074), .ZN(n10401) );
  NOR2_X1 U10827 ( .A1(n8528), .A2(n8474), .ZN(n8475) );
  INV_X1 U10828 ( .A(n8476), .ZN(n8478) );
  NAND2_X1 U10829 ( .A1(P3_REG1_REG_8__SCAN_IN), .A2(n11206), .ZN(n8479) );
  OAI21_X1 U10830 ( .B1(P3_REG1_REG_8__SCAN_IN), .B2(n11206), .A(n8479), .ZN(
        n10533) );
  NOR2_X1 U10831 ( .A1(n8423), .A2(n10851), .ZN(n10850) );
  NOR2_X1 U10832 ( .A1(n11306), .A2(n8480), .ZN(n8481) );
  NAND2_X1 U10833 ( .A1(n11393), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n8483) );
  OR2_X1 U10834 ( .A1(n11393), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n8482) );
  NAND2_X1 U10835 ( .A1(n8483), .A2(n8482), .ZN(n11443) );
  NOR2_X1 U10836 ( .A1(n8537), .A2(n8484), .ZN(n8485) );
  INV_X1 U10837 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n14684) );
  NAND2_X1 U10838 ( .A1(P3_REG1_REG_12__SCAN_IN), .A2(n11516), .ZN(n8486) );
  OAI21_X1 U10839 ( .B1(P3_REG1_REG_12__SCAN_IN), .B2(n11516), .A(n8486), .ZN(
        n11511) );
  NOR2_X1 U10840 ( .A1(n8540), .A2(n8487), .ZN(n8488) );
  INV_X1 U10841 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n14673) );
  NOR2_X1 U10842 ( .A1(n12777), .A2(n12776), .ZN(n8489) );
  NOR2_X1 U10843 ( .A1(n14623), .A2(n8490), .ZN(n8491) );
  INV_X1 U10844 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n14627) );
  XNOR2_X1 U10845 ( .A(n14646), .B(n8492), .ZN(n14653) );
  INV_X1 U10846 ( .A(n12820), .ZN(n10468) );
  NAND2_X1 U10847 ( .A1(n10468), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n8496) );
  INV_X1 U10848 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n8494) );
  NAND2_X1 U10849 ( .A1(n12820), .A2(n8494), .ZN(n8495) );
  AND2_X1 U10850 ( .A1(n8496), .A2(n8495), .ZN(n12814) );
  NAND2_X1 U10851 ( .A1(n12817), .A2(n8496), .ZN(n8498) );
  INV_X1 U10852 ( .A(n13295), .ZN(n8500) );
  INV_X1 U10853 ( .A(n8509), .ZN(n8499) );
  NAND2_X1 U10854 ( .A1(n8500), .A2(n12549), .ZN(n8514) );
  NAND2_X1 U10855 ( .A1(n8501), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8502) );
  MUX2_X1 U10856 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8502), .S(
        P3_IR_REG_22__SCAN_IN), .Z(n8503) );
  INV_X1 U10857 ( .A(n8505), .ZN(n8506) );
  NAND2_X1 U10858 ( .A1(n8506), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8508) );
  NAND2_X1 U10859 ( .A1(n11001), .A2(n8509), .ZN(n8511) );
  AND2_X1 U10860 ( .A1(n8511), .A2(n11392), .ZN(n8512) );
  NAND2_X1 U10861 ( .A1(n8514), .A2(n8512), .ZN(n8554) );
  INV_X1 U10862 ( .A(n8512), .ZN(n8513) );
  NOR2_X1 U10863 ( .A1(n12167), .A2(P3_STATE_REG_SCAN_IN), .ZN(n12646) );
  MUX2_X1 U10864 ( .A(n12743), .B(n8554), .S(n6485), .Z(n15139) );
  NOR2_X1 U10865 ( .A1(n15139), .A2(n12345), .ZN(n8515) );
  AOI211_X1 U10866 ( .C1(P3_ADDR_REG_19__SCAN_IN), .C2(n15097), .A(n12646), 
        .B(n8515), .ZN(n8516) );
  INV_X1 U10867 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n15099) );
  NOR3_X1 U10868 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), .A3(
        n15099), .ZN(n8521) );
  INV_X1 U10869 ( .A(n8520), .ZN(n10158) );
  NOR2_X1 U10870 ( .A1(n10549), .A2(n8522), .ZN(n8523) );
  AOI22_X1 U10871 ( .A1(n15122), .A2(P3_REG2_REG_4__SCAN_IN), .B1(n8371), .B2(
        n9597), .ZN(n15111) );
  NOR2_X1 U10872 ( .A1(n10923), .A2(n8525), .ZN(n8526) );
  AOI22_X1 U10873 ( .A1(n8528), .A2(P3_REG2_REG_6__SCAN_IN), .B1(n8527), .B2(
        n11074), .ZN(n10398) );
  NAND2_X1 U10874 ( .A1(n8530), .A2(n9618), .ZN(n8529) );
  INV_X1 U10875 ( .A(n8529), .ZN(n8531) );
  OAI21_X1 U10876 ( .B1(n8530), .B2(n9618), .A(n8529), .ZN(n15147) );
  NOR2_X1 U10877 ( .A1(n8402), .A2(n15147), .ZN(n15146) );
  NAND2_X1 U10878 ( .A1(P3_REG2_REG_8__SCAN_IN), .A2(n11206), .ZN(n8532) );
  OAI21_X1 U10879 ( .B1(P3_REG2_REG_8__SCAN_IN), .B2(n11206), .A(n8532), .ZN(
        n10527) );
  NOR2_X1 U10880 ( .A1(n10528), .A2(n10527), .ZN(n10526) );
  XNOR2_X1 U10881 ( .A(n8533), .B(n11306), .ZN(n10849) );
  NOR2_X1 U10882 ( .A1(n11306), .A2(n8533), .ZN(n8534) );
  NOR2_X1 U10883 ( .A1(n10848), .A2(n8534), .ZN(n11448) );
  NAND2_X1 U10884 ( .A1(n11393), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n8536) );
  OR2_X1 U10885 ( .A1(n11393), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n8535) );
  NAND2_X1 U10886 ( .A1(n8536), .A2(n8535), .ZN(n11447) );
  NOR2_X1 U10887 ( .A1(n8537), .A2(n6611), .ZN(n8538) );
  INV_X1 U10888 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n11427) );
  NAND2_X1 U10889 ( .A1(P3_REG2_REG_12__SCAN_IN), .A2(n11516), .ZN(n8539) );
  OAI21_X1 U10890 ( .B1(P3_REG2_REG_12__SCAN_IN), .B2(n11516), .A(n8539), .ZN(
        n11509) );
  NOR2_X1 U10891 ( .A1(n11510), .A2(n11509), .ZN(n11508) );
  NOR2_X1 U10892 ( .A1(n8540), .A2(n8541), .ZN(n8542) );
  INV_X1 U10893 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n12758) );
  NOR2_X1 U10894 ( .A1(n14623), .A2(n8543), .ZN(n8544) );
  INV_X1 U10895 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n14622) );
  XNOR2_X1 U10896 ( .A(n8543), .B(n14623), .ZN(n14621) );
  AOI22_X1 U10897 ( .A1(P3_REG2_REG_16__SCAN_IN), .A2(n14646), .B1(n10153), 
        .B2(n8545), .ZN(n14639) );
  NOR2_X1 U10898 ( .A1(n14646), .A2(n8545), .ZN(n8546) );
  NAND2_X1 U10899 ( .A1(n10468), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n8549) );
  INV_X1 U10900 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n8547) );
  NAND2_X1 U10901 ( .A1(n12820), .A2(n8547), .ZN(n8548) );
  NAND2_X1 U10902 ( .A1(n8549), .A2(n8548), .ZN(n12808) );
  INV_X1 U10903 ( .A(n8549), .ZN(n8550) );
  INV_X1 U10904 ( .A(n6485), .ZN(n8553) );
  NAND2_X1 U10905 ( .A1(n8553), .A2(n8552), .ZN(n10232) );
  NOR2_X1 U10906 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), 
        .ZN(n8560) );
  NAND4_X1 U10907 ( .A1(n8560), .A2(n8559), .A3(n8558), .A4(n8557), .ZN(n8924)
         );
  NOR2_X1 U10908 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), 
        .ZN(n8562) );
  NOR2_X1 U10909 ( .A1(P2_IR_REG_24__SCAN_IN), .A2(P2_IR_REG_23__SCAN_IN), 
        .ZN(n8561) );
  NOR2_X1 U10910 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(P2_IR_REG_28__SCAN_IN), 
        .ZN(n8564) );
  NAND2_X1 U10911 ( .A1(n9174), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n8570) );
  NAND2_X1 U10912 ( .A1(n8575), .A2(n8574), .ZN(n8576) );
  NOR2_X1 U10913 ( .A1(n8924), .A2(n8576), .ZN(n8577) );
  NAND2_X1 U10914 ( .A1(n8782), .A2(n8577), .ZN(n8585) );
  INV_X1 U10915 ( .A(n8585), .ZN(n8579) );
  INV_X1 U10916 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n8578) );
  INV_X1 U10917 ( .A(n8583), .ZN(n8581) );
  INV_X1 U10918 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n8580) );
  NAND2_X1 U10919 ( .A1(n8581), .A2(n8580), .ZN(n8587) );
  NAND2_X1 U10920 ( .A1(n8585), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8586) );
  XNOR2_X2 U10921 ( .A(n8586), .B(P2_IR_REG_19__SCAN_IN), .ZN(n10368) );
  NAND2_X1 U10922 ( .A1(n8611), .A2(n14992), .ZN(n14988) );
  INV_X1 U10923 ( .A(n8587), .ZN(n8589) );
  INV_X1 U10924 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n8588) );
  NAND2_X1 U10925 ( .A1(n8589), .A2(n8588), .ZN(n9227) );
  NAND2_X1 U10926 ( .A1(n6484), .A2(SI_0_), .ZN(n8591) );
  XNOR2_X1 U10927 ( .A(n8591), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n13874) );
  INV_X1 U10928 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n8594) );
  NAND2_X1 U10929 ( .A1(P2_IR_REG_27__SCAN_IN), .A2(P2_IR_REG_26__SCAN_IN), 
        .ZN(n8592) );
  NAND2_X1 U10930 ( .A1(n8592), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8593) );
  OAI21_X1 U10931 ( .B1(n8594), .B2(P2_IR_REG_31__SCAN_IN), .A(n8593), .ZN(
        n8595) );
  INV_X1 U10932 ( .A(n8595), .ZN(n8596) );
  AOI21_X1 U10933 ( .B1(n8601), .B2(n8597), .A(n8596), .ZN(n8599) );
  INV_X1 U10934 ( .A(n9242), .ZN(n8601) );
  NAND2_X1 U10935 ( .A1(n8601), .A2(n8600), .ZN(n9244) );
  AND2_X1 U10936 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_28__SCAN_IN), 
        .ZN(n8602) );
  NAND2_X1 U10937 ( .A1(n9244), .A2(n8602), .ZN(n8609) );
  INV_X1 U10938 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n8605) );
  NAND2_X1 U10939 ( .A1(P2_IR_REG_27__SCAN_IN), .A2(P2_IR_REG_28__SCAN_IN), 
        .ZN(n8603) );
  NAND2_X1 U10940 ( .A1(n8603), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8604) );
  OAI21_X1 U10941 ( .B1(n8605), .B2(P2_IR_REG_31__SCAN_IN), .A(n8604), .ZN(
        n8606) );
  NAND2_X1 U10942 ( .A1(n8609), .A2(n8608), .ZN(n9250) );
  INV_X1 U10943 ( .A(n10369), .ZN(n11812) );
  NAND2_X1 U10944 ( .A1(n11812), .A2(n10368), .ZN(n8613) );
  INV_X1 U10945 ( .A(n9991), .ZN(n8612) );
  NAND2_X1 U10946 ( .A1(n8613), .A2(n8612), .ZN(n8614) );
  NAND2_X1 U10947 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), 
        .ZN(n8616) );
  MUX2_X1 U10948 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8616), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n8619) );
  INV_X1 U10949 ( .A(n8639), .ZN(n8618) );
  NAND2_X1 U10950 ( .A1(n8619), .A2(n8618), .ZN(n14857) );
  INV_X1 U10951 ( .A(n14857), .ZN(n8620) );
  NAND2_X2 U10952 ( .A1(n8638), .A2(n8621), .ZN(n8657) );
  INV_X1 U10953 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n9572) );
  NAND2_X1 U10954 ( .A1(n9174), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n8624) );
  NAND2_X1 U10955 ( .A1(n8664), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n8623) );
  NAND2_X1 U10956 ( .A1(n8683), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n8622) );
  NAND2_X1 U10957 ( .A1(n9998), .A2(n9230), .ZN(n8625) );
  NAND2_X1 U10958 ( .A1(n8626), .A2(n8625), .ZN(n8632) );
  NAND2_X1 U10959 ( .A1(n8631), .A2(n8632), .ZN(n8630) );
  NAND2_X1 U10960 ( .A1(n9230), .A2(n10987), .ZN(n8628) );
  NAND2_X1 U10961 ( .A1(n9998), .A2(n8663), .ZN(n8627) );
  NAND2_X1 U10962 ( .A1(n8628), .A2(n8627), .ZN(n8629) );
  NAND2_X1 U10963 ( .A1(n8630), .A2(n8629), .ZN(n8636) );
  INV_X1 U10964 ( .A(n8631), .ZN(n8634) );
  NAND2_X1 U10965 ( .A1(n8634), .A2(n8633), .ZN(n8635) );
  NAND2_X1 U10966 ( .A1(n8636), .A2(n8635), .ZN(n8656) );
  INV_X1 U10967 ( .A(n9628), .ZN(n8637) );
  INV_X1 U10968 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n9600) );
  INV_X1 U10969 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n8783) );
  NOR2_X1 U10970 ( .A1(n8639), .A2(n8783), .ZN(n8640) );
  MUX2_X1 U10971 ( .A(n8783), .B(n8640), .S(P2_IR_REG_2__SCAN_IN), .Z(n8641)
         );
  INV_X1 U10972 ( .A(n8641), .ZN(n8644) );
  INV_X1 U10973 ( .A(n8642), .ZN(n8643) );
  NAND2_X1 U10974 ( .A1(n8644), .A2(n8643), .ZN(n9723) );
  NOR2_X1 U10975 ( .A1(n7440), .A2(n8645), .ZN(n8646) );
  NAND2_X1 U10976 ( .A1(n9087), .A2(n10769), .ZN(n8653) );
  NAND2_X1 U10977 ( .A1(n9174), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n8650) );
  NAND2_X1 U10978 ( .A1(n8684), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n8649) );
  NAND2_X1 U10979 ( .A1(n8683), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n8648) );
  NAND2_X1 U10980 ( .A1(n13448), .A2(n9035), .ZN(n8652) );
  NAND2_X1 U10981 ( .A1(n8653), .A2(n8652), .ZN(n8655) );
  NAND2_X1 U10982 ( .A1(n9570), .A2(n6483), .ZN(n8662) );
  NOR2_X1 U10983 ( .A1(n8642), .A2(n8783), .ZN(n8658) );
  MUX2_X1 U10984 ( .A(n8783), .B(n8658), .S(P2_IR_REG_3__SCAN_IN), .Z(n8660)
         );
  AND2_X1 U10985 ( .A1(n8642), .A2(n8659), .ZN(n8679) );
  NOR2_X1 U10986 ( .A1(n8660), .A2(n8679), .ZN(n9760) );
  AOI22_X1 U10987 ( .A1(n8965), .A2(P1_DATAO_REG_3__SCAN_IN), .B1(n8964), .B2(
        n9760), .ZN(n8661) );
  INV_X1 U10988 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n8686) );
  NAND2_X1 U10989 ( .A1(n8664), .A2(n8686), .ZN(n8668) );
  NAND2_X1 U10990 ( .A1(n8683), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n8667) );
  NAND2_X1 U10991 ( .A1(n9174), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n8666) );
  NAND2_X1 U10992 ( .A1(n8684), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n8665) );
  NAND4_X1 U10993 ( .A1(n8668), .A2(n8667), .A3(n8666), .A4(n8665), .ZN(n13447) );
  AOI22_X1 U10994 ( .A1(n10375), .A2(n9181), .B1(n13447), .B2(n9087), .ZN(
        n8674) );
  INV_X1 U10995 ( .A(n8674), .ZN(n8669) );
  NAND2_X1 U10996 ( .A1(n8673), .A2(n8669), .ZN(n8672) );
  NAND2_X1 U10997 ( .A1(n10375), .A2(n9172), .ZN(n8670) );
  OAI21_X1 U10998 ( .B1(n10357), .B2(n9230), .A(n8670), .ZN(n8671) );
  NAND2_X1 U10999 ( .A1(n8672), .A2(n8671), .ZN(n8677) );
  INV_X1 U11000 ( .A(n8673), .ZN(n8675) );
  NAND2_X1 U11001 ( .A1(n8675), .A2(n8674), .ZN(n8676) );
  INV_X1 U11002 ( .A(n8679), .ZN(n8697) );
  NAND2_X1 U11003 ( .A1(n8697), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8680) );
  XNOR2_X1 U11004 ( .A(n8680), .B(P2_IR_REG_4__SCAN_IN), .ZN(n9699) );
  AOI22_X1 U11005 ( .A1(n8965), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n8964), .B2(
        n9699), .ZN(n8681) );
  NAND2_X1 U11006 ( .A1(n15049), .A2(n9087), .ZN(n8693) );
  NAND2_X1 U11007 ( .A1(n9173), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n8691) );
  NAND2_X1 U11008 ( .A1(n8684), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n8690) );
  INV_X1 U11009 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n8685) );
  NAND2_X1 U11010 ( .A1(n8686), .A2(n8685), .ZN(n8687) );
  NAND2_X1 U11011 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n8707) );
  AND2_X1 U11012 ( .A1(n8687), .A2(n8707), .ZN(n14978) );
  NAND2_X1 U11013 ( .A1(n8664), .A2(n14978), .ZN(n8689) );
  NAND2_X1 U11014 ( .A1(n9174), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n8688) );
  NAND4_X1 U11015 ( .A1(n8691), .A2(n8690), .A3(n8689), .A4(n8688), .ZN(n13446) );
  NAND2_X1 U11016 ( .A1(n13446), .A2(n9181), .ZN(n8692) );
  NAND2_X1 U11017 ( .A1(n8693), .A2(n8692), .ZN(n8695) );
  AOI22_X1 U11018 ( .A1(n15049), .A2(n9181), .B1(n13446), .B2(n9172), .ZN(
        n8694) );
  NAND2_X1 U11019 ( .A1(n9619), .A2(n6483), .ZN(n8704) );
  NAND2_X1 U11020 ( .A1(n8699), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8698) );
  MUX2_X1 U11021 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8698), .S(
        P2_IR_REG_5__SCAN_IN), .Z(n8702) );
  INV_X1 U11022 ( .A(n8699), .ZN(n8701) );
  INV_X1 U11023 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n8700) );
  NAND2_X1 U11024 ( .A1(n8701), .A2(n8700), .ZN(n8725) );
  NAND2_X1 U11025 ( .A1(n8702), .A2(n8725), .ZN(n9711) );
  INV_X1 U11026 ( .A(n9711), .ZN(n9731) );
  AOI22_X1 U11027 ( .A1(n8965), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n8964), .B2(
        n9731), .ZN(n8703) );
  NAND2_X1 U11028 ( .A1(n8704), .A2(n8703), .ZN(n15058) );
  NAND2_X1 U11029 ( .A1(n15058), .A2(n9181), .ZN(n8714) );
  NAND2_X1 U11030 ( .A1(n8684), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n8712) );
  NAND2_X1 U11031 ( .A1(n9173), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n8711) );
  INV_X1 U11032 ( .A(n8707), .ZN(n8705) );
  NAND2_X1 U11033 ( .A1(n8705), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n8744) );
  INV_X1 U11034 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n8706) );
  NAND2_X1 U11035 ( .A1(n8707), .A2(n8706), .ZN(n8708) );
  AND2_X1 U11036 ( .A1(n8744), .A2(n8708), .ZN(n10745) );
  NAND2_X1 U11037 ( .A1(n8664), .A2(n10745), .ZN(n8710) );
  NAND2_X1 U11038 ( .A1(n9174), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n8709) );
  NAND4_X1 U11039 ( .A1(n8712), .A2(n8711), .A3(n8710), .A4(n8709), .ZN(n13445) );
  NAND2_X1 U11040 ( .A1(n13445), .A2(n9172), .ZN(n8713) );
  NAND2_X1 U11041 ( .A1(n8714), .A2(n8713), .ZN(n8719) );
  INV_X1 U11042 ( .A(n13445), .ZN(n10363) );
  NAND2_X1 U11043 ( .A1(n15058), .A2(n9087), .ZN(n8715) );
  OAI21_X1 U11044 ( .B1(n10363), .B2(n9230), .A(n8715), .ZN(n8716) );
  NAND2_X1 U11045 ( .A1(n8717), .A2(n8716), .ZN(n8723) );
  INV_X1 U11046 ( .A(n8718), .ZN(n8721) );
  INV_X1 U11047 ( .A(n8719), .ZN(n8720) );
  NAND2_X1 U11048 ( .A1(n8721), .A2(n8720), .ZN(n8722) );
  OR2_X1 U11049 ( .A1(n9633), .A2(n8678), .ZN(n8728) );
  NAND2_X1 U11050 ( .A1(n8725), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8724) );
  MUX2_X1 U11051 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8724), .S(
        P2_IR_REG_6__SCAN_IN), .Z(n8726) );
  AOI22_X1 U11052 ( .A1(n8965), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n8964), .B2(
        n9847), .ZN(n8727) );
  NAND2_X1 U11053 ( .A1(n8728), .A2(n8727), .ZN(n10574) );
  NAND2_X1 U11054 ( .A1(n10574), .A2(n9172), .ZN(n8734) );
  NAND2_X1 U11055 ( .A1(n8684), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n8732) );
  NAND2_X1 U11056 ( .A1(n9173), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n8731) );
  XNOR2_X1 U11057 ( .A(n8744), .B(P2_REG3_REG_6__SCAN_IN), .ZN(n10881) );
  NAND2_X1 U11058 ( .A1(n8664), .A2(n10881), .ZN(n8730) );
  NAND2_X1 U11059 ( .A1(n9174), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n8729) );
  NAND4_X1 U11060 ( .A1(n8732), .A2(n8731), .A3(n8730), .A4(n8729), .ZN(n13444) );
  NAND2_X1 U11061 ( .A1(n13444), .A2(n9181), .ZN(n8733) );
  AOI22_X1 U11062 ( .A1(n10574), .A2(n9181), .B1(n13444), .B2(n9172), .ZN(
        n8735) );
  OR2_X1 U11063 ( .A1(n9639), .A2(n8678), .ZN(n8739) );
  NAND2_X1 U11064 ( .A1(n8761), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8737) );
  XNOR2_X1 U11065 ( .A(n8737), .B(P2_IR_REG_7__SCAN_IN), .ZN(n13456) );
  AOI22_X1 U11066 ( .A1(n8965), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n8964), .B2(
        n13456), .ZN(n8738) );
  NAND2_X1 U11067 ( .A1(n8739), .A2(n8738), .ZN(n10709) );
  NAND2_X1 U11068 ( .A1(n10709), .A2(n9181), .ZN(n8751) );
  NAND2_X1 U11069 ( .A1(n8684), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n8749) );
  INV_X2 U11070 ( .A(n8765), .ZN(n9173) );
  NAND2_X1 U11071 ( .A1(n9173), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n8748) );
  INV_X1 U11072 ( .A(n8744), .ZN(n8741) );
  AND2_X1 U11073 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_REG3_REG_7__SCAN_IN), 
        .ZN(n8740) );
  NAND2_X1 U11074 ( .A1(n8741), .A2(n8740), .ZN(n8768) );
  INV_X1 U11075 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n8743) );
  INV_X1 U11076 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n8742) );
  OAI21_X1 U11077 ( .B1(n8744), .B2(n8743), .A(n8742), .ZN(n8745) );
  AND2_X1 U11078 ( .A1(n8768), .A2(n8745), .ZN(n10587) );
  NAND2_X1 U11079 ( .A1(n8664), .A2(n10587), .ZN(n8747) );
  NAND2_X1 U11080 ( .A1(n9174), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n8746) );
  NAND4_X1 U11081 ( .A1(n8749), .A2(n8748), .A3(n8747), .A4(n8746), .ZN(n13443) );
  NAND2_X1 U11082 ( .A1(n13443), .A2(n9172), .ZN(n8750) );
  NAND2_X1 U11083 ( .A1(n8751), .A2(n8750), .ZN(n8756) );
  INV_X1 U11084 ( .A(n13443), .ZN(n10708) );
  NAND2_X1 U11085 ( .A1(n10709), .A2(n9172), .ZN(n8752) );
  OAI21_X1 U11086 ( .B1(n10708), .B2(n9230), .A(n8752), .ZN(n8753) );
  NAND2_X1 U11087 ( .A1(n8754), .A2(n8753), .ZN(n8760) );
  INV_X1 U11088 ( .A(n8755), .ZN(n8758) );
  INV_X1 U11089 ( .A(n8756), .ZN(n8757) );
  NAND2_X1 U11090 ( .A1(n8758), .A2(n8757), .ZN(n8759) );
  OR2_X1 U11091 ( .A1(n9647), .A2(n8678), .ZN(n8764) );
  OAI21_X1 U11092 ( .B1(n8761), .B2(P2_IR_REG_7__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8762) );
  XNOR2_X1 U11093 ( .A(n8762), .B(P2_IR_REG_8__SCAN_IN), .ZN(n13472) );
  AOI22_X1 U11094 ( .A1(n8965), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n13472), 
        .B2(n8964), .ZN(n8763) );
  NAND2_X1 U11095 ( .A1(n15068), .A2(n9172), .ZN(n8775) );
  NAND2_X1 U11096 ( .A1(n9173), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n8773) );
  NAND2_X1 U11097 ( .A1(n8684), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n8772) );
  INV_X1 U11098 ( .A(n8768), .ZN(n8766) );
  NAND2_X1 U11099 ( .A1(n8766), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n8791) );
  INV_X1 U11100 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n8767) );
  NAND2_X1 U11101 ( .A1(n8768), .A2(n8767), .ZN(n8769) );
  AND2_X1 U11102 ( .A1(n8791), .A2(n8769), .ZN(n10721) );
  NAND2_X1 U11103 ( .A1(n8664), .A2(n10721), .ZN(n8771) );
  NAND2_X1 U11104 ( .A1(n9174), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n8770) );
  NAND4_X1 U11105 ( .A1(n8773), .A2(n8772), .A3(n8771), .A4(n8770), .ZN(n13442) );
  NAND2_X1 U11106 ( .A1(n13442), .A2(n9181), .ZN(n8774) );
  NAND2_X1 U11107 ( .A1(n8775), .A2(n8774), .ZN(n8776) );
  NAND2_X1 U11108 ( .A1(n8777), .A2(n8776), .ZN(n8780) );
  AOI22_X1 U11109 ( .A1(n15068), .A2(n9181), .B1(n13442), .B2(n9172), .ZN(
        n8778) );
  NAND2_X1 U11110 ( .A1(n8780), .A2(n8779), .ZN(n8781) );
  OR2_X1 U11111 ( .A1(n9652), .A2(n8678), .ZN(n8789) );
  NOR2_X1 U11112 ( .A1(n8782), .A2(n8783), .ZN(n8784) );
  MUX2_X1 U11113 ( .A(n8783), .B(n8784), .S(P2_IR_REG_9__SCAN_IN), .Z(n8787)
         );
  INV_X1 U11114 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n8785) );
  NAND2_X1 U11115 ( .A1(n8782), .A2(n8785), .ZN(n8925) );
  INV_X1 U11116 ( .A(n8925), .ZN(n8786) );
  NOR2_X1 U11117 ( .A1(n8787), .A2(n8786), .ZN(n9902) );
  AOI22_X1 U11118 ( .A1(n8965), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n8964), .B2(
        n9902), .ZN(n8788) );
  NAND2_X1 U11119 ( .A1(n8789), .A2(n8788), .ZN(n10918) );
  NAND2_X1 U11120 ( .A1(n10918), .A2(n9181), .ZN(n8798) );
  NAND2_X1 U11121 ( .A1(n9173), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n8796) );
  NAND2_X1 U11122 ( .A1(n8684), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n8795) );
  NAND2_X1 U11123 ( .A1(n8791), .A2(n8790), .ZN(n8792) );
  AND2_X1 U11124 ( .A1(n8806), .A2(n8792), .ZN(n10912) );
  NAND2_X1 U11125 ( .A1(n8664), .A2(n10912), .ZN(n8794) );
  NAND2_X1 U11126 ( .A1(n9174), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n8793) );
  NAND4_X1 U11127 ( .A1(n8796), .A2(n8795), .A3(n8794), .A4(n8793), .ZN(n13441) );
  NAND2_X1 U11128 ( .A1(n13441), .A2(n9172), .ZN(n8797) );
  NAND2_X1 U11129 ( .A1(n8798), .A2(n8797), .ZN(n8800) );
  AOI22_X1 U11130 ( .A1(n10918), .A2(n9172), .B1(n9181), .B2(n13441), .ZN(
        n8799) );
  NAND2_X1 U11131 ( .A1(n8925), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8801) );
  XNOR2_X1 U11132 ( .A(n8801), .B(P2_IR_REG_10__SCAN_IN), .ZN(n10102) );
  AOI22_X1 U11133 ( .A1(n8965), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n8964), 
        .B2(n10102), .ZN(n8802) );
  NAND2_X1 U11134 ( .A1(n11059), .A2(n9087), .ZN(n8813) );
  NAND2_X1 U11135 ( .A1(n8684), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n8811) );
  NAND2_X1 U11136 ( .A1(n9173), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n8810) );
  INV_X1 U11137 ( .A(n8806), .ZN(n8804) );
  NAND2_X1 U11138 ( .A1(n8804), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n8840) );
  INV_X1 U11139 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n8805) );
  NAND2_X1 U11140 ( .A1(n8806), .A2(n8805), .ZN(n8807) );
  AND2_X1 U11141 ( .A1(n8840), .A2(n8807), .ZN(n11054) );
  NAND2_X1 U11142 ( .A1(n8664), .A2(n11054), .ZN(n8809) );
  NAND2_X1 U11143 ( .A1(n9174), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n8808) );
  NAND4_X1 U11144 ( .A1(n8811), .A2(n8810), .A3(n8809), .A4(n8808), .ZN(n13440) );
  NAND2_X1 U11145 ( .A1(n13440), .A2(n9181), .ZN(n8812) );
  NAND2_X1 U11146 ( .A1(n8813), .A2(n8812), .ZN(n8818) );
  NAND2_X1 U11147 ( .A1(n8817), .A2(n8818), .ZN(n8816) );
  INV_X1 U11148 ( .A(n13440), .ZN(n10955) );
  NAND2_X1 U11149 ( .A1(n11059), .A2(n9181), .ZN(n8814) );
  OAI21_X1 U11150 ( .B1(n10955), .B2(n9035), .A(n8814), .ZN(n8815) );
  NAND2_X1 U11151 ( .A1(n9932), .A2(n6483), .ZN(n8823) );
  NAND2_X1 U11152 ( .A1(n8832), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8821) );
  XNOR2_X1 U11153 ( .A(n8821), .B(P2_IR_REG_11__SCAN_IN), .ZN(n13494) );
  AOI22_X1 U11154 ( .A1(n8965), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n8964), 
        .B2(n13494), .ZN(n8822) );
  NAND2_X1 U11155 ( .A1(n11276), .A2(n9181), .ZN(n8829) );
  NAND2_X1 U11156 ( .A1(n8684), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n8827) );
  NAND2_X1 U11157 ( .A1(n9173), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n8826) );
  XNOR2_X1 U11158 ( .A(n8840), .B(P2_REG3_REG_11__SCAN_IN), .ZN(n11285) );
  NAND2_X1 U11159 ( .A1(n8664), .A2(n11285), .ZN(n8825) );
  NAND2_X1 U11160 ( .A1(n9174), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n8824) );
  NAND4_X1 U11161 ( .A1(n8827), .A2(n8826), .A3(n8825), .A4(n8824), .ZN(n13439) );
  NAND2_X1 U11162 ( .A1(n13439), .A2(n9087), .ZN(n8828) );
  NAND2_X1 U11163 ( .A1(n8829), .A2(n8828), .ZN(n8831) );
  AOI22_X1 U11164 ( .A1(n11276), .A2(n9172), .B1(n9181), .B2(n13439), .ZN(
        n8830) );
  NAND2_X1 U11165 ( .A1(n10167), .A2(n6483), .ZN(n8836) );
  NOR2_X1 U11166 ( .A1(n8832), .A2(P2_IR_REG_11__SCAN_IN), .ZN(n8856) );
  INV_X1 U11167 ( .A(n8856), .ZN(n8833) );
  NAND2_X1 U11168 ( .A1(n8833), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8834) );
  XNOR2_X1 U11169 ( .A(n8834), .B(P2_IR_REG_12__SCAN_IN), .ZN(n13497) );
  AOI22_X1 U11170 ( .A1(n8965), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n8964), 
        .B2(n13497), .ZN(n8835) );
  NAND2_X1 U11171 ( .A1(n14716), .A2(n9087), .ZN(n8847) );
  NAND2_X1 U11172 ( .A1(n8684), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n8845) );
  NAND2_X1 U11173 ( .A1(n9173), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n8844) );
  INV_X1 U11174 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n8838) );
  INV_X1 U11175 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n8837) );
  OAI21_X1 U11176 ( .B1(n8840), .B2(n8838), .A(n8837), .ZN(n8841) );
  NAND2_X1 U11177 ( .A1(P2_REG3_REG_11__SCAN_IN), .A2(P2_REG3_REG_12__SCAN_IN), 
        .ZN(n8839) );
  AND2_X1 U11178 ( .A1(n8841), .A2(n8864), .ZN(n14714) );
  NAND2_X1 U11179 ( .A1(n8664), .A2(n14714), .ZN(n8843) );
  NAND2_X1 U11180 ( .A1(n9174), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n8842) );
  NAND4_X1 U11181 ( .A1(n8845), .A2(n8844), .A3(n8843), .A4(n8842), .ZN(n13438) );
  NAND2_X1 U11182 ( .A1(n13438), .A2(n9181), .ZN(n8846) );
  NAND2_X1 U11183 ( .A1(n8847), .A2(n8846), .ZN(n8851) );
  INV_X1 U11184 ( .A(n13438), .ZN(n11252) );
  NAND2_X1 U11185 ( .A1(n14716), .A2(n9181), .ZN(n8848) );
  OAI21_X1 U11186 ( .B1(n11252), .B2(n9035), .A(n8848), .ZN(n8849) );
  INV_X1 U11187 ( .A(n8850), .ZN(n8853) );
  NAND2_X1 U11188 ( .A1(n8853), .A2(n8852), .ZN(n8854) );
  NAND2_X1 U11189 ( .A1(n10280), .A2(n6483), .ZN(n8861) );
  INV_X1 U11190 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n8855) );
  NAND2_X1 U11191 ( .A1(n8856), .A2(n8855), .ZN(n8858) );
  NAND2_X1 U11192 ( .A1(n8858), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8857) );
  MUX2_X1 U11193 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8857), .S(
        P2_IR_REG_13__SCAN_IN), .Z(n8859) );
  AND2_X1 U11194 ( .A1(n8859), .A2(n8894), .ZN(n14903) );
  AOI22_X1 U11195 ( .A1(n14903), .A2(n8964), .B1(n8965), .B2(
        P1_DATAO_REG_13__SCAN_IN), .ZN(n8860) );
  NAND2_X1 U11196 ( .A1(n11638), .A2(n9181), .ZN(n8871) );
  NAND2_X1 U11197 ( .A1(n9173), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n8869) );
  INV_X1 U11198 ( .A(n8864), .ZN(n8862) );
  NAND2_X1 U11199 ( .A1(n8862), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n8877) );
  INV_X1 U11200 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n8863) );
  NAND2_X1 U11201 ( .A1(n8864), .A2(n8863), .ZN(n8865) );
  AND2_X1 U11202 ( .A1(n8877), .A2(n8865), .ZN(n11627) );
  NAND2_X1 U11203 ( .A1(n8664), .A2(n11627), .ZN(n8868) );
  NAND2_X1 U11204 ( .A1(n9174), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n8867) );
  NAND2_X1 U11205 ( .A1(n8684), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n8866) );
  NAND4_X1 U11206 ( .A1(n8869), .A2(n8868), .A3(n8867), .A4(n8866), .ZN(n13437) );
  NAND2_X1 U11207 ( .A1(n13437), .A2(n9087), .ZN(n8870) );
  NAND2_X1 U11208 ( .A1(n8871), .A2(n8870), .ZN(n8873) );
  AOI22_X1 U11209 ( .A1(n11638), .A2(n9172), .B1(n9181), .B2(n13437), .ZN(
        n8872) );
  NAND2_X1 U11210 ( .A1(n10522), .A2(n6483), .ZN(n8876) );
  NAND2_X1 U11211 ( .A1(n8894), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8874) );
  XNOR2_X1 U11212 ( .A(n8874), .B(P2_IR_REG_14__SCAN_IN), .ZN(n14918) );
  AOI22_X1 U11213 ( .A1(n14918), .A2(n8964), .B1(n8965), .B2(
        P1_DATAO_REG_14__SCAN_IN), .ZN(n8875) );
  NAND2_X1 U11214 ( .A1(n14702), .A2(n9172), .ZN(n8884) );
  NAND2_X1 U11215 ( .A1(n8684), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n8882) );
  NAND2_X1 U11216 ( .A1(n8877), .A2(n11671), .ZN(n8878) );
  AND2_X1 U11217 ( .A1(n8897), .A2(n8878), .ZN(n14701) );
  NAND2_X1 U11218 ( .A1(n14701), .A2(n8664), .ZN(n8881) );
  NAND2_X1 U11219 ( .A1(n9173), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n8880) );
  NAND2_X1 U11220 ( .A1(n9174), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n8879) );
  NAND4_X1 U11221 ( .A1(n8882), .A2(n8881), .A3(n8880), .A4(n8879), .ZN(n13436) );
  NAND2_X1 U11222 ( .A1(n13436), .A2(n9181), .ZN(n8883) );
  NAND2_X1 U11223 ( .A1(n8884), .A2(n8883), .ZN(n8889) );
  NAND2_X1 U11224 ( .A1(n8888), .A2(n8889), .ZN(n8887) );
  INV_X1 U11225 ( .A(n13436), .ZN(n11559) );
  NAND2_X1 U11226 ( .A1(n14702), .A2(n9181), .ZN(n8885) );
  OAI21_X1 U11227 ( .B1(n11559), .B2(n9035), .A(n8885), .ZN(n8886) );
  NAND2_X1 U11228 ( .A1(n8887), .A2(n8886), .ZN(n8893) );
  INV_X1 U11229 ( .A(n8888), .ZN(n8891) );
  NAND2_X1 U11230 ( .A1(n8891), .A2(n8890), .ZN(n8892) );
  NAND2_X1 U11231 ( .A1(n10780), .A2(n6483), .ZN(n8896) );
  OAI21_X1 U11232 ( .B1(n8894), .B2(P2_IR_REG_14__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8911) );
  XNOR2_X1 U11233 ( .A(n8911), .B(P2_IR_REG_15__SCAN_IN), .ZN(n14923) );
  AOI22_X1 U11234 ( .A1(n14923), .A2(n8964), .B1(n8965), .B2(
        P1_DATAO_REG_15__SCAN_IN), .ZN(n8895) );
  NAND2_X1 U11235 ( .A1(n11802), .A2(n9181), .ZN(n8904) );
  NAND2_X1 U11236 ( .A1(n8897), .A2(n11727), .ZN(n8898) );
  NAND2_X1 U11237 ( .A1(n8917), .A2(n8898), .ZN(n11726) );
  NAND2_X1 U11238 ( .A1(n8684), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n8900) );
  NAND2_X1 U11239 ( .A1(n9173), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n8899) );
  AND2_X1 U11240 ( .A1(n8900), .A2(n8899), .ZN(n8902) );
  NAND2_X1 U11241 ( .A1(n9174), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n8901) );
  OAI211_X1 U11242 ( .C1(n11726), .C2(n9147), .A(n8902), .B(n8901), .ZN(n13435) );
  NAND2_X1 U11243 ( .A1(n13435), .A2(n9087), .ZN(n8903) );
  NAND2_X1 U11244 ( .A1(n8904), .A2(n8903), .ZN(n8907) );
  AOI22_X1 U11245 ( .A1(n11802), .A2(n9172), .B1(n9181), .B2(n13435), .ZN(
        n8905) );
  AOI21_X1 U11246 ( .B1(n8908), .B2(n8907), .A(n8905), .ZN(n8906) );
  INV_X1 U11247 ( .A(n8906), .ZN(n8909) );
  NAND2_X1 U11248 ( .A1(n10975), .A2(n6483), .ZN(n8915) );
  INV_X1 U11249 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n8910) );
  NAND2_X1 U11250 ( .A1(n8911), .A2(n8910), .ZN(n8912) );
  NAND2_X1 U11251 ( .A1(n8912), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8913) );
  XNOR2_X1 U11252 ( .A(n8913), .B(P2_IR_REG_16__SCAN_IN), .ZN(n14935) );
  AOI22_X1 U11253 ( .A1(n14935), .A2(n8964), .B1(P1_DATAO_REG_16__SCAN_IN), 
        .B2(n8965), .ZN(n8914) );
  NAND2_X1 U11254 ( .A1(n11964), .A2(n9172), .ZN(n8923) );
  INV_X1 U11255 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n8921) );
  INV_X1 U11256 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n11866) );
  NAND2_X1 U11257 ( .A1(n8917), .A2(n11866), .ZN(n8918) );
  NAND2_X1 U11258 ( .A1(n8930), .A2(n8918), .ZN(n11865) );
  OR2_X1 U11259 ( .A1(n11865), .A2(n9147), .ZN(n8920) );
  AOI22_X1 U11260 ( .A1(n8684), .A2(P2_REG1_REG_16__SCAN_IN), .B1(n9173), .B2(
        P2_REG2_REG_16__SCAN_IN), .ZN(n8919) );
  OAI211_X1 U11261 ( .C1(n9150), .C2(n8921), .A(n8920), .B(n8919), .ZN(n13434)
         );
  NAND2_X1 U11262 ( .A1(n13434), .A2(n9181), .ZN(n8922) );
  NAND2_X1 U11263 ( .A1(n8923), .A2(n8922), .ZN(n8941) );
  NAND2_X1 U11264 ( .A1(n11122), .A2(n6483), .ZN(n8928) );
  OR2_X1 U11265 ( .A1(n8925), .A2(n8924), .ZN(n8947) );
  NAND2_X1 U11266 ( .A1(n8947), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8926) );
  XNOR2_X1 U11267 ( .A(n8926), .B(P2_IR_REG_17__SCAN_IN), .ZN(n14943) );
  AOI22_X1 U11268 ( .A1(n8965), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n8964), 
        .B2(n14943), .ZN(n8927) );
  INV_X1 U11269 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n13505) );
  INV_X1 U11270 ( .A(n8930), .ZN(n8929) );
  INV_X1 U11271 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n12002) );
  NAND2_X1 U11272 ( .A1(n8930), .A2(n12002), .ZN(n8931) );
  NAND2_X1 U11273 ( .A1(n8951), .A2(n8931), .ZN(n12001) );
  OR2_X1 U11274 ( .A1(n12001), .A2(n9147), .ZN(n8933) );
  AOI22_X1 U11275 ( .A1(n9174), .A2(P2_REG0_REG_17__SCAN_IN), .B1(n9173), .B2(
        P2_REG2_REG_17__SCAN_IN), .ZN(n8932) );
  OAI211_X1 U11276 ( .C1(n6932), .C2(n13505), .A(n8933), .B(n8932), .ZN(n13567) );
  AOI22_X1 U11277 ( .A1(n13569), .A2(n9172), .B1(n8663), .B2(n13567), .ZN(
        n8936) );
  NAND2_X1 U11278 ( .A1(n13569), .A2(n9181), .ZN(n8935) );
  NAND2_X1 U11279 ( .A1(n13567), .A2(n9087), .ZN(n8934) );
  NAND2_X1 U11280 ( .A1(n8935), .A2(n8934), .ZN(n8944) );
  NAND2_X1 U11281 ( .A1(n8936), .A2(n8944), .ZN(n8937) );
  INV_X1 U11282 ( .A(n13434), .ZN(n11961) );
  NAND2_X1 U11283 ( .A1(n11964), .A2(n9181), .ZN(n8938) );
  OAI21_X1 U11284 ( .B1(n11961), .B2(n9035), .A(n8938), .ZN(n8939) );
  AOI21_X1 U11285 ( .B1(n8942), .B2(n8941), .A(n8940), .ZN(n8945) );
  NOR2_X1 U11286 ( .A1(n13569), .A2(n13567), .ZN(n8943) );
  NAND2_X1 U11287 ( .A1(n11377), .A2(n6483), .ZN(n8950) );
  OAI21_X1 U11288 ( .B1(n8947), .B2(P2_IR_REG_17__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8948) );
  XNOR2_X1 U11289 ( .A(n8948), .B(P2_IR_REG_18__SCAN_IN), .ZN(n14958) );
  AOI22_X1 U11290 ( .A1(n8965), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n8964), 
        .B2(n14958), .ZN(n8949) );
  NAND2_X1 U11291 ( .A1(n13745), .A2(n9172), .ZN(n8960) );
  INV_X1 U11292 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n13411) );
  NAND2_X1 U11293 ( .A1(n8951), .A2(n13411), .ZN(n8952) );
  AND2_X1 U11294 ( .A1(n8970), .A2(n8952), .ZN(n13748) );
  NAND2_X1 U11295 ( .A1(n13748), .A2(n8664), .ZN(n8958) );
  INV_X1 U11296 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8955) );
  NAND2_X1 U11297 ( .A1(n9173), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n8954) );
  NAND2_X1 U11298 ( .A1(n9174), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n8953) );
  OAI211_X1 U11299 ( .C1(n6932), .C2(n8955), .A(n8954), .B(n8953), .ZN(n8956)
         );
  INV_X1 U11300 ( .A(n8956), .ZN(n8957) );
  NAND2_X1 U11301 ( .A1(n8958), .A2(n8957), .ZN(n13566) );
  NAND2_X1 U11302 ( .A1(n13566), .A2(n9181), .ZN(n8959) );
  INV_X1 U11303 ( .A(n13566), .ZN(n13573) );
  NAND2_X1 U11304 ( .A1(n13745), .A2(n9181), .ZN(n8961) );
  OAI21_X1 U11305 ( .B1(n13573), .B2(n9181), .A(n8961), .ZN(n8962) );
  NAND2_X1 U11306 ( .A1(n8963), .A2(n6483), .ZN(n8967) );
  AOI22_X1 U11307 ( .A1(n8965), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n8964), 
        .B2(n10368), .ZN(n8966) );
  NAND2_X1 U11308 ( .A1(n13734), .A2(n9181), .ZN(n8979) );
  INV_X1 U11309 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n8969) );
  NAND2_X1 U11310 ( .A1(n8970), .A2(n8969), .ZN(n8971) );
  NAND2_X1 U11311 ( .A1(n8986), .A2(n8971), .ZN(n13730) );
  OR2_X1 U11312 ( .A1(n13730), .A2(n9147), .ZN(n8977) );
  INV_X1 U11313 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n8974) );
  NAND2_X1 U11314 ( .A1(n9174), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n8973) );
  NAND2_X1 U11315 ( .A1(n9173), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n8972) );
  OAI211_X1 U11316 ( .C1(n6932), .C2(n8974), .A(n8973), .B(n8972), .ZN(n8975)
         );
  INV_X1 U11317 ( .A(n8975), .ZN(n8976) );
  NAND2_X1 U11318 ( .A1(n13575), .A2(n9172), .ZN(n8978) );
  NAND2_X1 U11319 ( .A1(n8979), .A2(n8978), .ZN(n8981) );
  AOI22_X1 U11320 ( .A1(n13734), .A2(n9172), .B1(n9181), .B2(n13575), .ZN(
        n8980) );
  NOR2_X1 U11321 ( .A1(n8982), .A2(n8981), .ZN(n8983) );
  NAND2_X1 U11322 ( .A1(n11492), .A2(n6483), .ZN(n8985) );
  OR2_X1 U11323 ( .A1(n8657), .A2(n7139), .ZN(n8984) );
  NAND2_X1 U11324 ( .A1(n13822), .A2(n9172), .ZN(n8995) );
  INV_X1 U11325 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n13394) );
  NAND2_X1 U11326 ( .A1(n8986), .A2(n13394), .ZN(n8987) );
  AND2_X1 U11327 ( .A1(n9000), .A2(n8987), .ZN(n13719) );
  NAND2_X1 U11328 ( .A1(n13719), .A2(n8664), .ZN(n8993) );
  INV_X1 U11329 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n8990) );
  NAND2_X1 U11330 ( .A1(n9173), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n8989) );
  NAND2_X1 U11331 ( .A1(n8684), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n8988) );
  OAI211_X1 U11332 ( .C1(n8990), .C2(n9150), .A(n8989), .B(n8988), .ZN(n8991)
         );
  INV_X1 U11333 ( .A(n8991), .ZN(n8992) );
  NAND2_X1 U11334 ( .A1(n8993), .A2(n8992), .ZN(n13361) );
  NAND2_X1 U11335 ( .A1(n13361), .A2(n9035), .ZN(n8994) );
  AOI22_X1 U11336 ( .A1(n13822), .A2(n9181), .B1(n13361), .B2(n9172), .ZN(
        n8996) );
  NAND2_X1 U11337 ( .A1(n11613), .A2(n6483), .ZN(n8998) );
  OR2_X1 U11338 ( .A1(n8657), .A2(n11619), .ZN(n8997) );
  NAND2_X1 U11339 ( .A1(n13817), .A2(n9035), .ZN(n9008) );
  INV_X1 U11340 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n13362) );
  NAND2_X1 U11341 ( .A1(n9000), .A2(n13362), .ZN(n9001) );
  NAND2_X1 U11342 ( .A1(n9024), .A2(n9001), .ZN(n13704) );
  OR2_X1 U11343 ( .A1(n13704), .A2(n9147), .ZN(n9006) );
  INV_X1 U11344 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n13122) );
  NAND2_X1 U11345 ( .A1(n9174), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n9003) );
  NAND2_X1 U11346 ( .A1(n9173), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n9002) );
  OAI211_X1 U11347 ( .C1(n6932), .C2(n13122), .A(n9003), .B(n9002), .ZN(n9004)
         );
  INV_X1 U11348 ( .A(n9004), .ZN(n9005) );
  NAND2_X1 U11349 ( .A1(n9006), .A2(n9005), .ZN(n13433) );
  NAND2_X1 U11350 ( .A1(n13433), .A2(n9172), .ZN(n9007) );
  NAND2_X1 U11351 ( .A1(n9008), .A2(n9007), .ZN(n9013) );
  NAND2_X1 U11352 ( .A1(n9012), .A2(n9013), .ZN(n9011) );
  AOI22_X1 U11353 ( .A1(n13817), .A2(n9172), .B1(n9181), .B2(n13433), .ZN(
        n9009) );
  INV_X1 U11354 ( .A(n9009), .ZN(n9010) );
  NAND2_X1 U11355 ( .A1(n9011), .A2(n9010), .ZN(n9017) );
  NAND2_X1 U11356 ( .A1(n9015), .A2(n9014), .ZN(n9016) );
  INV_X1 U11357 ( .A(n9018), .ZN(n9020) );
  NAND2_X1 U11358 ( .A1(n9020), .A2(n9019), .ZN(n11809) );
  AND2_X1 U11359 ( .A1(n6483), .A2(n11810), .ZN(n9021) );
  NAND2_X1 U11360 ( .A1(n11809), .A2(n9021), .ZN(n9023) );
  OR2_X1 U11361 ( .A1(n8657), .A2(n11813), .ZN(n9022) );
  INV_X1 U11362 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n13403) );
  NAND2_X1 U11363 ( .A1(n9024), .A2(n13403), .ZN(n9025) );
  AND2_X1 U11364 ( .A1(n9044), .A2(n9025), .ZN(n13691) );
  NAND2_X1 U11365 ( .A1(n13691), .A2(n8664), .ZN(n9031) );
  INV_X1 U11366 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n9028) );
  NAND2_X1 U11367 ( .A1(n8684), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n9027) );
  NAND2_X1 U11368 ( .A1(n9173), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n9026) );
  OAI211_X1 U11369 ( .C1(n9028), .C2(n9150), .A(n9027), .B(n9026), .ZN(n9029)
         );
  INV_X1 U11370 ( .A(n9029), .ZN(n9030) );
  NAND2_X1 U11371 ( .A1(n9031), .A2(n9030), .ZN(n13545) );
  AND2_X1 U11372 ( .A1(n13545), .A2(n9181), .ZN(n9032) );
  AOI21_X1 U11373 ( .B1(n13811), .B2(n9172), .A(n9032), .ZN(n9038) );
  INV_X1 U11374 ( .A(n9038), .ZN(n9033) );
  INV_X1 U11375 ( .A(n13545), .ZN(n13579) );
  NAND2_X1 U11376 ( .A1(n13811), .A2(n9035), .ZN(n9034) );
  OAI21_X1 U11377 ( .B1(n13579), .B2(n9035), .A(n9034), .ZN(n9036) );
  INV_X1 U11378 ( .A(n9037), .ZN(n9039) );
  NAND2_X1 U11379 ( .A1(n9039), .A2(n9038), .ZN(n9040) );
  NAND2_X1 U11380 ( .A1(n11888), .A2(n6483), .ZN(n9042) );
  INV_X1 U11381 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n11892) );
  OR2_X1 U11382 ( .A1(n8657), .A2(n11892), .ZN(n9041) );
  NAND2_X1 U11383 ( .A1(n13806), .A2(n9181), .ZN(n9052) );
  NAND2_X1 U11384 ( .A1(n9044), .A2(n9043), .ZN(n9045) );
  NAND2_X1 U11385 ( .A1(n9058), .A2(n9045), .ZN(n13675) );
  INV_X1 U11386 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n9048) );
  NAND2_X1 U11387 ( .A1(n8684), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n9047) );
  NAND2_X1 U11388 ( .A1(n9173), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n9046) );
  OAI211_X1 U11389 ( .C1(n9048), .C2(n9150), .A(n9047), .B(n9046), .ZN(n9049)
         );
  INV_X1 U11390 ( .A(n9049), .ZN(n9050) );
  NAND2_X1 U11391 ( .A1(n13580), .A2(n9172), .ZN(n9051) );
  AOI22_X1 U11392 ( .A1(n13806), .A2(n9087), .B1(n9181), .B2(n13580), .ZN(
        n9053) );
  NAND2_X1 U11393 ( .A1(n11814), .A2(n6483), .ZN(n9055) );
  INV_X1 U11394 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n11816) );
  OR2_X1 U11395 ( .A1(n8657), .A2(n11816), .ZN(n9054) );
  NAND2_X1 U11396 ( .A1(n13795), .A2(n9172), .ZN(n9066) );
  INV_X1 U11397 ( .A(n9058), .ZN(n9056) );
  NAND2_X1 U11398 ( .A1(n9056), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n9079) );
  INV_X1 U11399 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n9057) );
  NAND2_X1 U11400 ( .A1(n9058), .A2(n9057), .ZN(n9059) );
  AND2_X1 U11401 ( .A1(n9079), .A2(n9059), .ZN(n13660) );
  NAND2_X1 U11402 ( .A1(n13660), .A2(n8664), .ZN(n9064) );
  INV_X1 U11403 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n13658) );
  NAND2_X1 U11404 ( .A1(n9174), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n9061) );
  NAND2_X1 U11405 ( .A1(n8684), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n9060) );
  OAI211_X1 U11406 ( .C1(n8765), .C2(n13658), .A(n9061), .B(n9060), .ZN(n9062)
         );
  INV_X1 U11407 ( .A(n9062), .ZN(n9063) );
  NAND2_X1 U11408 ( .A1(n9064), .A2(n9063), .ZN(n13550) );
  NAND2_X1 U11409 ( .A1(n13550), .A2(n9181), .ZN(n9065) );
  NAND2_X1 U11410 ( .A1(n9066), .A2(n9065), .ZN(n9071) );
  NAND2_X1 U11411 ( .A1(n9070), .A2(n9071), .ZN(n9069) );
  NAND2_X1 U11412 ( .A1(n13795), .A2(n9181), .ZN(n9067) );
  OAI21_X1 U11413 ( .B1(n13581), .B2(n9035), .A(n9067), .ZN(n9068) );
  NAND2_X1 U11414 ( .A1(n9069), .A2(n9068), .ZN(n9075) );
  INV_X1 U11415 ( .A(n9070), .ZN(n9073) );
  INV_X1 U11416 ( .A(n9071), .ZN(n9072) );
  NAND2_X1 U11417 ( .A1(n9073), .A2(n9072), .ZN(n9074) );
  NAND2_X1 U11418 ( .A1(n11879), .A2(n6483), .ZN(n9077) );
  OR2_X1 U11419 ( .A1(n8657), .A2(n11881), .ZN(n9076) );
  NAND2_X1 U11420 ( .A1(n13791), .A2(n8663), .ZN(n9089) );
  INV_X1 U11421 ( .A(n9079), .ZN(n9078) );
  NAND2_X1 U11422 ( .A1(n9078), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n9098) );
  INV_X1 U11423 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n13371) );
  NAND2_X1 U11424 ( .A1(n9079), .A2(n13371), .ZN(n9080) );
  NAND2_X1 U11425 ( .A1(n9098), .A2(n9080), .ZN(n13645) );
  INV_X1 U11426 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n9083) );
  NAND2_X1 U11427 ( .A1(n8684), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n9082) );
  NAND2_X1 U11428 ( .A1(n9173), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n9081) );
  OAI211_X1 U11429 ( .C1(n9083), .C2(n9150), .A(n9082), .B(n9081), .ZN(n9084)
         );
  INV_X1 U11430 ( .A(n9084), .ZN(n9085) );
  NAND2_X1 U11431 ( .A1(n13552), .A2(n9087), .ZN(n9088) );
  NAND2_X1 U11432 ( .A1(n9089), .A2(n9088), .ZN(n9091) );
  INV_X1 U11433 ( .A(n9091), .ZN(n9090) );
  AOI22_X1 U11434 ( .A1(n13791), .A2(n9087), .B1(n9181), .B2(n13552), .ZN(
        n9092) );
  INV_X1 U11435 ( .A(n9092), .ZN(n9093) );
  NAND2_X1 U11436 ( .A1(n12007), .A2(n6483), .ZN(n9096) );
  OR2_X1 U11437 ( .A1(n8657), .A2(n9094), .ZN(n9095) );
  NAND2_X1 U11438 ( .A1(n13635), .A2(n9172), .ZN(n9107) );
  INV_X1 U11439 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n9097) );
  NAND2_X1 U11440 ( .A1(n9098), .A2(n9097), .ZN(n9099) );
  NAND2_X1 U11441 ( .A1(n13632), .A2(n8664), .ZN(n9105) );
  INV_X1 U11442 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n9102) );
  NAND2_X1 U11443 ( .A1(n8684), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n9101) );
  NAND2_X1 U11444 ( .A1(n9173), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n9100) );
  OAI211_X1 U11445 ( .C1(n9102), .C2(n9150), .A(n9101), .B(n9100), .ZN(n9103)
         );
  INV_X1 U11446 ( .A(n9103), .ZN(n9104) );
  NAND2_X1 U11447 ( .A1(n13432), .A2(n9035), .ZN(n9106) );
  NAND2_X1 U11448 ( .A1(n9107), .A2(n9106), .ZN(n9109) );
  AOI22_X1 U11449 ( .A1(n13635), .A2(n9181), .B1(n13432), .B2(n9172), .ZN(
        n9108) );
  AOI21_X1 U11450 ( .B1(n9110), .B2(n9109), .A(n9108), .ZN(n9161) );
  NOR2_X1 U11451 ( .A1(n9110), .A2(n9109), .ZN(n9160) );
  NAND2_X1 U11452 ( .A1(n13861), .A2(n6483), .ZN(n9112) );
  INV_X1 U11453 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n13862) );
  OR2_X1 U11454 ( .A1(n8657), .A2(n13862), .ZN(n9111) );
  NAND2_X2 U11455 ( .A1(n9112), .A2(n9111), .ZN(n13528) );
  INV_X1 U11456 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n9115) );
  NAND2_X1 U11457 ( .A1(n9173), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n9114) );
  NAND2_X1 U11458 ( .A1(n8684), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n9113) );
  OAI211_X1 U11459 ( .C1(n9150), .C2(n9115), .A(n9114), .B(n9113), .ZN(n9774)
         );
  XNOR2_X1 U11460 ( .A(n13528), .B(n9774), .ZN(n9202) );
  NAND2_X1 U11461 ( .A1(n13869), .A2(n6483), .ZN(n9117) );
  OR2_X1 U11462 ( .A1(n8657), .A2(n13871), .ZN(n9116) );
  NAND2_X1 U11463 ( .A1(n9129), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n13562) );
  OR2_X1 U11464 ( .A1(n13562), .A2(n9147), .ZN(n9123) );
  INV_X1 U11465 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n9120) );
  NAND2_X1 U11466 ( .A1(n9173), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n9119) );
  NAND2_X1 U11467 ( .A1(n8684), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n9118) );
  OAI211_X1 U11468 ( .C1(n9120), .C2(n9150), .A(n9119), .B(n9118), .ZN(n9121)
         );
  INV_X1 U11469 ( .A(n9121), .ZN(n9122) );
  NAND2_X1 U11470 ( .A1(n9123), .A2(n9122), .ZN(n12615) );
  AND2_X1 U11471 ( .A1(n12615), .A2(n9172), .ZN(n9124) );
  AOI21_X1 U11472 ( .B1(n13763), .B2(n9035), .A(n9124), .ZN(n9185) );
  NAND2_X1 U11473 ( .A1(n13763), .A2(n9172), .ZN(n9126) );
  NAND2_X1 U11474 ( .A1(n12615), .A2(n9035), .ZN(n9125) );
  NAND2_X1 U11475 ( .A1(n9126), .A2(n9125), .ZN(n9184) );
  NAND2_X1 U11476 ( .A1(n9185), .A2(n9184), .ZN(n9190) );
  NAND2_X1 U11477 ( .A1(n12121), .A2(n6483), .ZN(n9128) );
  OR2_X1 U11478 ( .A1(n8657), .A2(n12278), .ZN(n9127) );
  NAND2_X2 U11479 ( .A1(n9128), .A2(n9127), .ZN(n13769) );
  INV_X1 U11480 ( .A(n9129), .ZN(n9146) );
  INV_X1 U11481 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n12618) );
  NAND2_X1 U11482 ( .A1(n9146), .A2(n12618), .ZN(n9130) );
  NAND2_X1 U11483 ( .A1(n13562), .A2(n9130), .ZN(n13609) );
  INV_X1 U11484 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n9133) );
  NAND2_X1 U11485 ( .A1(n8684), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n9132) );
  NAND2_X1 U11486 ( .A1(n9173), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n9131) );
  OAI211_X1 U11487 ( .C1(n9133), .C2(n9150), .A(n9132), .B(n9131), .ZN(n9134)
         );
  INV_X1 U11488 ( .A(n9134), .ZN(n9135) );
  AND2_X1 U11489 ( .A1(n13431), .A2(n9172), .ZN(n9137) );
  AOI21_X1 U11490 ( .B1(n13769), .B2(n9181), .A(n9137), .ZN(n9189) );
  NAND2_X1 U11491 ( .A1(n13769), .A2(n9172), .ZN(n9139) );
  NAND2_X1 U11492 ( .A1(n13431), .A2(n9181), .ZN(n9138) );
  NAND2_X1 U11493 ( .A1(n9139), .A2(n9138), .ZN(n9188) );
  NAND2_X1 U11494 ( .A1(n9189), .A2(n9188), .ZN(n9140) );
  AND2_X1 U11495 ( .A1(n9190), .A2(n9140), .ZN(n9141) );
  AND2_X1 U11496 ( .A1(n9202), .A2(n9141), .ZN(n9162) );
  NAND2_X1 U11497 ( .A1(n12047), .A2(n6483), .ZN(n9143) );
  OR2_X1 U11498 ( .A1(n8657), .A2(n12563), .ZN(n9142) );
  NAND2_X1 U11499 ( .A1(n9144), .A2(n13340), .ZN(n9145) );
  NAND2_X1 U11500 ( .A1(n9146), .A2(n9145), .ZN(n13621) );
  INV_X1 U11501 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n9151) );
  NAND2_X1 U11502 ( .A1(n8684), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n9149) );
  NAND2_X1 U11503 ( .A1(n9173), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n9148) );
  OAI211_X1 U11504 ( .C1(n9151), .C2(n9150), .A(n9149), .B(n9148), .ZN(n9152)
         );
  INV_X1 U11505 ( .A(n9152), .ZN(n9153) );
  AND2_X1 U11506 ( .A1(n13585), .A2(n9172), .ZN(n9155) );
  AOI21_X1 U11507 ( .B1(n13779), .B2(n9035), .A(n9155), .ZN(n9164) );
  NAND2_X1 U11508 ( .A1(n13779), .A2(n9172), .ZN(n9157) );
  NAND2_X1 U11509 ( .A1(n13585), .A2(n9181), .ZN(n9156) );
  NAND2_X1 U11510 ( .A1(n9157), .A2(n9156), .ZN(n9163) );
  NAND2_X1 U11511 ( .A1(n9164), .A2(n9163), .ZN(n9158) );
  AND2_X1 U11512 ( .A1(n9162), .A2(n9158), .ZN(n9159) );
  OAI21_X1 U11513 ( .B1(n9161), .B2(n9160), .A(n9159), .ZN(n9197) );
  INV_X1 U11514 ( .A(n9162), .ZN(n9165) );
  MUX2_X1 U11515 ( .A(n9774), .B(n9035), .S(n13528), .Z(n9167) );
  NAND2_X1 U11516 ( .A1(n9774), .A2(n9181), .ZN(n9166) );
  NAND2_X1 U11517 ( .A1(n9167), .A2(n9166), .ZN(n9187) );
  NAND2_X1 U11518 ( .A1(n12626), .A2(n6483), .ZN(n9170) );
  OR2_X1 U11519 ( .A1(n8657), .A2(n13866), .ZN(n9169) );
  NAND2_X1 U11520 ( .A1(n6713), .A2(n14992), .ZN(n9226) );
  NAND2_X1 U11521 ( .A1(n11523), .A2(n13516), .ZN(n9978) );
  AND2_X1 U11522 ( .A1(n11616), .A2(n9978), .ZN(n9171) );
  AND2_X1 U11523 ( .A1(n9226), .A2(n9171), .ZN(n9179) );
  NAND2_X1 U11524 ( .A1(n9172), .A2(n9774), .ZN(n9178) );
  NAND2_X1 U11525 ( .A1(n8684), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n9177) );
  NAND2_X1 U11526 ( .A1(n9173), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n9176) );
  NAND2_X1 U11527 ( .A1(n9174), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n9175) );
  AND3_X1 U11528 ( .A1(n9177), .A2(n9176), .A3(n9175), .ZN(n13589) );
  AOI21_X1 U11529 ( .B1(n9179), .B2(n9178), .A(n13589), .ZN(n9180) );
  AOI21_X1 U11530 ( .B1(n13521), .B2(n9181), .A(n9180), .ZN(n9199) );
  NAND2_X1 U11531 ( .A1(n13521), .A2(n9172), .ZN(n9183) );
  INV_X1 U11532 ( .A(n13589), .ZN(n13430) );
  NAND2_X1 U11533 ( .A1(n13430), .A2(n9181), .ZN(n9182) );
  NAND2_X1 U11534 ( .A1(n9183), .A2(n9182), .ZN(n9198) );
  OAI22_X1 U11535 ( .A1(n9199), .A2(n9198), .B1(n9185), .B2(n9184), .ZN(n9186)
         );
  NAND2_X1 U11536 ( .A1(n9187), .A2(n9186), .ZN(n9194) );
  INV_X1 U11537 ( .A(n9188), .ZN(n9192) );
  INV_X1 U11538 ( .A(n9189), .ZN(n9191) );
  NAND4_X1 U11539 ( .A1(n9202), .A2(n9192), .A3(n9191), .A4(n9190), .ZN(n9193)
         );
  NAND2_X1 U11540 ( .A1(n9194), .A2(n9193), .ZN(n9195) );
  NAND2_X1 U11541 ( .A1(n9197), .A2(n9196), .ZN(n9201) );
  NAND2_X1 U11542 ( .A1(n9199), .A2(n9198), .ZN(n9200) );
  NAND2_X1 U11543 ( .A1(n9201), .A2(n9200), .ZN(n9263) );
  INV_X1 U11544 ( .A(n9202), .ZN(n9222) );
  XOR2_X1 U11545 ( .A(n13430), .B(n13521), .Z(n9221) );
  INV_X1 U11546 ( .A(n12615), .ZN(n9203) );
  XNOR2_X1 U11547 ( .A(n13763), .B(n9203), .ZN(n13588) );
  NAND2_X1 U11548 ( .A1(n13769), .A2(n13431), .ZN(n13558) );
  OAI21_X1 U11549 ( .B1(n13769), .B2(n13431), .A(n13558), .ZN(n13587) );
  NAND2_X1 U11550 ( .A1(n13635), .A2(n13556), .ZN(n13584) );
  NAND2_X1 U11551 ( .A1(n13583), .A2(n13584), .ZN(n13629) );
  INV_X1 U11552 ( .A(n13433), .ZN(n13578) );
  XNOR2_X1 U11553 ( .A(n13817), .B(n13578), .ZN(n13706) );
  NAND2_X1 U11554 ( .A1(n13734), .A2(n13575), .ZN(n13538) );
  NAND2_X1 U11555 ( .A1(n13539), .A2(n13538), .ZN(n13727) );
  INV_X1 U11556 ( .A(n13435), .ZN(n11796) );
  XNOR2_X1 U11557 ( .A(n11802), .B(n11796), .ZN(n11560) );
  XNOR2_X1 U11558 ( .A(n14702), .B(n11559), .ZN(n11548) );
  INV_X1 U11559 ( .A(n13437), .ZN(n11556) );
  XNOR2_X1 U11560 ( .A(n11638), .B(n11556), .ZN(n11253) );
  XNOR2_X1 U11561 ( .A(n14716), .B(n11252), .ZN(n14717) );
  XNOR2_X1 U11562 ( .A(n11276), .B(n13439), .ZN(n11245) );
  INV_X1 U11563 ( .A(n13442), .ZN(n10729) );
  NAND2_X1 U11564 ( .A1(n15068), .A2(n10729), .ZN(n10726) );
  OR2_X1 U11565 ( .A1(n15068), .A2(n10729), .ZN(n9204) );
  NAND2_X1 U11566 ( .A1(n10726), .A2(n9204), .ZN(n10728) );
  XNOR2_X1 U11567 ( .A(n10709), .B(n10708), .ZN(n10705) );
  XNOR2_X1 U11568 ( .A(n10574), .B(n13444), .ZN(n10569) );
  INV_X1 U11569 ( .A(n9205), .ZN(n10076) );
  NAND2_X1 U11570 ( .A1(n10076), .A2(n14990), .ZN(n10075) );
  NAND2_X1 U11571 ( .A1(n9205), .A2(n6945), .ZN(n9206) );
  AND2_X1 U11572 ( .A1(n10075), .A2(n9206), .ZN(n15020) );
  NAND4_X1 U11573 ( .A1(n15020), .A2(n9207), .A3(n10349), .A4(n10343), .ZN(
        n9208) );
  NOR2_X1 U11574 ( .A1(n9208), .A2(n10356), .ZN(n9209) );
  XNOR2_X1 U11575 ( .A(n15058), .B(n13445), .ZN(n10751) );
  NAND4_X1 U11576 ( .A1(n10569), .A2(n9209), .A3(n14971), .A4(n10751), .ZN(
        n9210) );
  NOR3_X1 U11577 ( .A1(n10728), .A2(n10705), .A3(n9210), .ZN(n9211) );
  XNOR2_X1 U11578 ( .A(n10918), .B(n13441), .ZN(n10733) );
  NAND4_X1 U11579 ( .A1(n11245), .A2(n9211), .A3(n10953), .A4(n10733), .ZN(
        n9212) );
  OR4_X1 U11580 ( .A1(n11548), .A2(n11253), .A3(n14717), .A4(n9212), .ZN(n9213) );
  NOR2_X1 U11581 ( .A1(n11560), .A2(n9213), .ZN(n9214) );
  XNOR2_X1 U11582 ( .A(n13569), .B(n13567), .ZN(n11965) );
  XNOR2_X1 U11583 ( .A(n11964), .B(n13434), .ZN(n11959) );
  NAND4_X1 U11584 ( .A1(n13727), .A2(n9214), .A3(n11965), .A4(n11959), .ZN(
        n9216) );
  NAND2_X1 U11585 ( .A1(n13822), .A2(n13540), .ZN(n13576) );
  OR2_X1 U11586 ( .A1(n13822), .A2(n13540), .ZN(n9215) );
  NAND2_X1 U11587 ( .A1(n13576), .A2(n9215), .ZN(n13715) );
  XNOR2_X1 U11588 ( .A(n13745), .B(n13573), .ZN(n13742) );
  NOR4_X1 U11589 ( .A1(n13706), .A2(n9216), .A3(n13715), .A4(n13742), .ZN(
        n9217) );
  XOR2_X1 U11590 ( .A(n13581), .B(n13795), .Z(n13665) );
  NAND3_X1 U11591 ( .A1(n13687), .A2(n9217), .A3(n13665), .ZN(n9218) );
  INV_X1 U11592 ( .A(n13552), .ZN(n13582) );
  XNOR2_X1 U11593 ( .A(n13791), .B(n13582), .ZN(n13647) );
  NOR3_X1 U11594 ( .A1(n13629), .A2(n9218), .A3(n13647), .ZN(n9219) );
  NAND4_X1 U11595 ( .A1(n13587), .A2(n9219), .A3(n13617), .A4(n13669), .ZN(
        n9220) );
  XNOR2_X1 U11596 ( .A(n9223), .B(n10368), .ZN(n9224) );
  NOR2_X1 U11597 ( .A1(n9224), .A2(n11616), .ZN(n9257) );
  NAND2_X1 U11598 ( .A1(n11616), .A2(n9207), .ZN(n10370) );
  OR2_X1 U11599 ( .A1(n10370), .A2(n13516), .ZN(n9225) );
  AND2_X1 U11600 ( .A1(n9226), .A2(n9225), .ZN(n9255) );
  INV_X1 U11601 ( .A(n9255), .ZN(n9229) );
  INV_X1 U11602 ( .A(n9982), .ZN(n9671) );
  AND2_X1 U11603 ( .A1(n9671), .A2(P2_STATE_REG_SCAN_IN), .ZN(n11889) );
  OAI21_X1 U11604 ( .B1(n9257), .B2(n9229), .A(n11889), .ZN(n9262) );
  INV_X1 U11605 ( .A(n9774), .ZN(n13527) );
  OR3_X1 U11606 ( .A1(n13528), .A2(n13527), .A3(n9172), .ZN(n9232) );
  NAND3_X1 U11607 ( .A1(n13528), .A2(n13527), .A3(n9230), .ZN(n9231) );
  NOR2_X1 U11608 ( .A1(n11616), .A2(n11523), .ZN(n9233) );
  OAI22_X1 U11609 ( .A1(n10368), .A2(n9233), .B1(n6713), .B2(n9991), .ZN(n9234) );
  NAND2_X1 U11610 ( .A1(n11889), .A2(n9234), .ZN(n9235) );
  NOR2_X1 U11611 ( .A1(n7456), .A2(n9235), .ZN(n9236) );
  NAND2_X1 U11612 ( .A1(n9263), .A2(n9236), .ZN(n9261) );
  INV_X1 U11613 ( .A(P2_B_REG_SCAN_IN), .ZN(n13525) );
  NAND2_X1 U11614 ( .A1(n9238), .A2(n9237), .ZN(n9239) );
  NAND2_X1 U11615 ( .A1(n9242), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9243) );
  MUX2_X1 U11616 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9243), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n9245) );
  NAND2_X1 U11617 ( .A1(n9246), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9247) );
  MUX2_X1 U11618 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9247), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n9248) );
  NAND2_X1 U11619 ( .A1(n9969), .A2(n9966), .ZN(n9249) );
  INV_X1 U11620 ( .A(n15016), .ZN(n15013) );
  NAND2_X1 U11621 ( .A1(n6713), .A2(n11616), .ZN(n9987) );
  OR2_X1 U11622 ( .A1(n9987), .A2(n9251), .ZN(n13591) );
  NOR4_X1 U11623 ( .A1(n15013), .A2(n13526), .A3(n9978), .A4(n13591), .ZN(
        n9252) );
  AOI211_X1 U11624 ( .C1(n11889), .C2(n11812), .A(n13525), .B(n9252), .ZN(
        n9258) );
  NOR2_X1 U11625 ( .A1(n7456), .A2(n9258), .ZN(n9253) );
  INV_X1 U11626 ( .A(n9253), .ZN(n9259) );
  INV_X1 U11627 ( .A(n9258), .ZN(n9254) );
  AOI21_X1 U11628 ( .B1(n9255), .B2(n9254), .A(n9253), .ZN(n9256) );
  OAI222_X1 U11629 ( .A1(n9259), .A2(n10348), .B1(n11889), .B2(n9258), .C1(
        n9257), .C2(n9256), .ZN(n9260) );
  OAI211_X1 U11630 ( .C1(n9263), .C2(n9262), .A(n9261), .B(n9260), .ZN(
        P2_U3328) );
  INV_X4 U11631 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  NAND2_X1 U11632 ( .A1(n13949), .A2(n9275), .ZN(n9267) );
  NAND2_X1 U11633 ( .A1(n14320), .A2(n12057), .ZN(n9266) );
  NAND2_X1 U11634 ( .A1(n9267), .A2(n9266), .ZN(n9269) );
  NAND2_X1 U11635 ( .A1(n14483), .A2(n12108), .ZN(n9268) );
  INV_X2 U11636 ( .A(n9501), .ZN(n9295) );
  XNOR2_X1 U11637 ( .A(n9269), .B(n9295), .ZN(n9371) );
  AOI22_X1 U11638 ( .A1(n13949), .A2(n12061), .B1(n9278), .B2(n14320), .ZN(
        n9369) );
  INV_X1 U11639 ( .A(n9369), .ZN(n9370) );
  NAND2_X1 U11640 ( .A1(n14046), .A2(n12057), .ZN(n9272) );
  INV_X1 U11641 ( .A(n9265), .ZN(n9274) );
  NAND2_X1 U11642 ( .A1(n9274), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n9271) );
  AOI222_X1 U11643 ( .A1(n14046), .A2(n9278), .B1(n9274), .B2(
        P1_IR_REG_0__SCAN_IN), .C1(n9548), .C2(n12065), .ZN(n10134) );
  NAND2_X1 U11644 ( .A1(n10134), .A2(n10133), .ZN(n10132) );
  OAI21_X1 U11645 ( .B1(n9501), .B2(n10133), .A(n10132), .ZN(n10143) );
  AOI22_X1 U11646 ( .A1(n12065), .A2(n9913), .B1(n9275), .B2(n14345), .ZN(
        n9276) );
  XNOR2_X1 U11647 ( .A(n9276), .B(n9295), .ZN(n9281) );
  INV_X2 U11648 ( .A(n9278), .ZN(n9344) );
  OAI22_X1 U11649 ( .A1(n10177), .A2(n9344), .B1(n10184), .B2(n9287), .ZN(
        n9279) );
  XNOR2_X1 U11650 ( .A(n9281), .B(n9279), .ZN(n10144) );
  INV_X1 U11651 ( .A(n9279), .ZN(n9280) );
  OAI22_X1 U11652 ( .A1(n10510), .A2(n9344), .B1(n6691), .B2(n9287), .ZN(n9284) );
  XNOR2_X1 U11653 ( .A(n9284), .B(n9285), .ZN(n10139) );
  OAI21_X2 U11654 ( .B1(n10138), .B2(n10139), .A(n9286), .ZN(n10333) );
  AOI22_X1 U11655 ( .A1(n12066), .A2(n14042), .B1(n9275), .B2(n10605), .ZN(
        n9290) );
  XNOR2_X1 U11656 ( .A(n9290), .B(n9295), .ZN(n9291) );
  AOI22_X1 U11657 ( .A1(n9278), .A2(n14042), .B1(n12057), .B2(n10605), .ZN(
        n9292) );
  XNOR2_X1 U11658 ( .A(n9291), .B(n9292), .ZN(n10334) );
  INV_X1 U11659 ( .A(n9291), .ZN(n9294) );
  INV_X1 U11660 ( .A(n9292), .ZN(n9293) );
  AOI22_X1 U11661 ( .A1(n9278), .A2(n14041), .B1(n12065), .B2(n10837), .ZN(
        n9298) );
  XNOR2_X1 U11662 ( .A(n9297), .B(n9299), .ZN(n10692) );
  AOI22_X1 U11663 ( .A1(n12061), .A2(n14041), .B1(n9275), .B2(n10837), .ZN(
        n9296) );
  XOR2_X1 U11664 ( .A(n9295), .B(n9296), .Z(n10691) );
  INV_X1 U11665 ( .A(n9297), .ZN(n9300) );
  INV_X1 U11666 ( .A(n10897), .ZN(n10668) );
  OAI22_X1 U11667 ( .A1(n10668), .A2(n9287), .B1(n9508), .B2(n9344), .ZN(n9303) );
  AOI22_X1 U11668 ( .A1(n10897), .A2(n9275), .B1(n12065), .B2(n14040), .ZN(
        n9302) );
  XOR2_X1 U11669 ( .A(n9295), .B(n9302), .Z(n10895) );
  NAND2_X1 U11670 ( .A1(n14002), .A2(n9275), .ZN(n9305) );
  NAND2_X1 U11671 ( .A1(n14039), .A2(n12057), .ZN(n9304) );
  NAND2_X1 U11672 ( .A1(n9305), .A2(n9304), .ZN(n9306) );
  XNOR2_X1 U11673 ( .A(n9306), .B(n9295), .ZN(n9308) );
  AOI22_X1 U11674 ( .A1(n14002), .A2(n12061), .B1(n9278), .B2(n14039), .ZN(
        n9307) );
  XNOR2_X1 U11675 ( .A(n9308), .B(n9307), .ZN(n13993) );
  INV_X1 U11676 ( .A(n9307), .ZN(n9309) );
  AOI22_X1 U11677 ( .A1(n11200), .A2(n9275), .B1(n12065), .B2(n14038), .ZN(
        n9310) );
  XNOR2_X1 U11678 ( .A(n9310), .B(n9295), .ZN(n9312) );
  NOR2_X1 U11679 ( .A1(n11241), .A2(n9344), .ZN(n9311) );
  AOI21_X1 U11680 ( .B1(n11200), .B2(n12066), .A(n9311), .ZN(n9313) );
  XNOR2_X1 U11681 ( .A(n9312), .B(n9313), .ZN(n11193) );
  OR2_X1 U11682 ( .A1(n9313), .A2(n9312), .ZN(n9314) );
  NAND2_X1 U11683 ( .A1(n11471), .A2(n9275), .ZN(n9316) );
  NAND2_X1 U11684 ( .A1(n14037), .A2(n12061), .ZN(n9315) );
  NAND2_X1 U11685 ( .A1(n9316), .A2(n9315), .ZN(n9317) );
  XNOR2_X1 U11686 ( .A(n9317), .B(n9501), .ZN(n9320) );
  NOR2_X1 U11687 ( .A1(n9515), .A2(n9344), .ZN(n9318) );
  AOI21_X1 U11688 ( .B1(n11471), .B2(n12066), .A(n9318), .ZN(n9319) );
  NAND2_X1 U11689 ( .A1(n9320), .A2(n9319), .ZN(n9321) );
  OAI21_X1 U11690 ( .B1(n9320), .B2(n9319), .A(n9321), .ZN(n11463) );
  NOR2_X1 U11691 ( .A1(n11465), .A2(n9344), .ZN(n9322) );
  AOI21_X1 U11692 ( .B1(n11767), .B2(n12066), .A(n9322), .ZN(n9325) );
  AOI22_X1 U11693 ( .A1(n11767), .A2(n9275), .B1(n12066), .B2(n14036), .ZN(
        n9323) );
  XNOR2_X1 U11694 ( .A(n9323), .B(n9295), .ZN(n11762) );
  NAND2_X1 U11695 ( .A1(n11663), .A2(n9275), .ZN(n9327) );
  NAND2_X1 U11696 ( .A1(n14035), .A2(n12057), .ZN(n9326) );
  NAND2_X1 U11697 ( .A1(n9327), .A2(n9326), .ZN(n9328) );
  XNOR2_X1 U11698 ( .A(n9328), .B(n9501), .ZN(n9331) );
  NOR2_X1 U11699 ( .A1(n11418), .A2(n9344), .ZN(n9329) );
  AOI21_X1 U11700 ( .B1(n11663), .B2(n12066), .A(n9329), .ZN(n9330) );
  NOR2_X1 U11701 ( .A1(n9331), .A2(n9330), .ZN(n11656) );
  AOI22_X1 U11702 ( .A1(n11571), .A2(n12061), .B1(n9278), .B2(n14034), .ZN(
        n9334) );
  AOI22_X1 U11703 ( .A1(n11571), .A2(n9275), .B1(n12066), .B2(n14034), .ZN(
        n9332) );
  XNOR2_X1 U11704 ( .A(n9332), .B(n9295), .ZN(n9333) );
  XOR2_X1 U11705 ( .A(n9334), .B(n9333), .Z(n11822) );
  NOR2_X1 U11706 ( .A1(n11824), .A2(n9344), .ZN(n9336) );
  AOI21_X1 U11707 ( .B1(n11488), .B2(n12066), .A(n9336), .ZN(n9341) );
  NAND2_X1 U11708 ( .A1(n11488), .A2(n9275), .ZN(n9338) );
  NAND2_X1 U11709 ( .A1(n14033), .A2(n12061), .ZN(n9337) );
  NAND2_X1 U11710 ( .A1(n9338), .A2(n9337), .ZN(n9339) );
  XNOR2_X1 U11711 ( .A(n9339), .B(n9295), .ZN(n9340) );
  XOR2_X1 U11712 ( .A(n9341), .B(n9340), .Z(n11893) );
  INV_X1 U11713 ( .A(n9341), .ZN(n9342) );
  NOR2_X1 U11714 ( .A1(n11898), .A2(n9344), .ZN(n9345) );
  AOI21_X1 U11715 ( .B1(n11736), .B2(n12066), .A(n9345), .ZN(n9348) );
  AOI22_X1 U11716 ( .A1(n11736), .A2(n9275), .B1(n12066), .B2(n14032), .ZN(
        n9346) );
  XNOR2_X1 U11717 ( .A(n9346), .B(n9295), .ZN(n9347) );
  XOR2_X1 U11718 ( .A(n9348), .B(n9347), .Z(n12022) );
  INV_X1 U11719 ( .A(n9347), .ZN(n9350) );
  INV_X1 U11720 ( .A(n9348), .ZN(n9349) );
  NAND2_X1 U11721 ( .A1(n9350), .A2(n9349), .ZN(n9351) );
  AOI22_X1 U11722 ( .A1(n13892), .A2(n9275), .B1(n12066), .B2(n14031), .ZN(
        n9352) );
  XNOR2_X1 U11723 ( .A(n9352), .B(n9295), .ZN(n9354) );
  AOI22_X1 U11724 ( .A1(n13892), .A2(n12061), .B1(n9278), .B2(n14031), .ZN(
        n9355) );
  XNOR2_X1 U11725 ( .A(n9354), .B(n9355), .ZN(n13886) );
  INV_X1 U11726 ( .A(n13886), .ZN(n9353) );
  NAND2_X1 U11727 ( .A1(n9354), .A2(n9355), .ZN(n9356) );
  AOI22_X1 U11728 ( .A1(n14019), .A2(n9275), .B1(n12065), .B2(n14030), .ZN(
        n9357) );
  XNOR2_X1 U11729 ( .A(n9357), .B(n9295), .ZN(n9359) );
  INV_X1 U11730 ( .A(n9359), .ZN(n9358) );
  AOI22_X1 U11731 ( .A1(n14019), .A2(n12061), .B1(n9278), .B2(n14030), .ZN(
        n14009) );
  NAND2_X1 U11732 ( .A1(n14008), .A2(n14009), .ZN(n9361) );
  NAND2_X1 U11733 ( .A1(n9360), .A2(n9359), .ZN(n14007) );
  NAND2_X1 U11734 ( .A1(n14425), .A2(n9275), .ZN(n9363) );
  NAND2_X1 U11735 ( .A1(n12038), .A2(n12061), .ZN(n9362) );
  NAND2_X1 U11736 ( .A1(n9363), .A2(n9362), .ZN(n9364) );
  XNOR2_X1 U11737 ( .A(n9364), .B(n9295), .ZN(n9367) );
  AOI22_X1 U11738 ( .A1(n14425), .A2(n12061), .B1(n9278), .B2(n12038), .ZN(
        n9365) );
  XNOR2_X1 U11739 ( .A(n9367), .B(n9365), .ZN(n13932) );
  INV_X1 U11740 ( .A(n9365), .ZN(n9366) );
  XNOR2_X1 U11741 ( .A(n9371), .B(n9369), .ZN(n13943) );
  NAND2_X1 U11742 ( .A1(n14414), .A2(n9275), .ZN(n9373) );
  NAND2_X1 U11743 ( .A1(n14029), .A2(n12061), .ZN(n9372) );
  NAND2_X1 U11744 ( .A1(n9373), .A2(n9372), .ZN(n9374) );
  XNOR2_X1 U11745 ( .A(n9374), .B(n9295), .ZN(n9375) );
  AOI22_X1 U11746 ( .A1(n14414), .A2(n12061), .B1(n9278), .B2(n14029), .ZN(
        n9376) );
  XNOR2_X1 U11747 ( .A(n9375), .B(n9376), .ZN(n13982) );
  INV_X1 U11748 ( .A(n9375), .ZN(n9377) );
  NAND2_X1 U11749 ( .A1(n9377), .A2(n9376), .ZN(n9378) );
  AND2_X1 U11750 ( .A1(n14322), .A2(n9278), .ZN(n9379) );
  AOI21_X1 U11751 ( .B1(n14409), .B2(n12066), .A(n9379), .ZN(n9385) );
  NAND2_X1 U11752 ( .A1(n14409), .A2(n9275), .ZN(n9381) );
  NAND2_X1 U11753 ( .A1(n14322), .A2(n12061), .ZN(n9380) );
  NAND2_X1 U11754 ( .A1(n9381), .A2(n9380), .ZN(n9382) );
  XNOR2_X1 U11755 ( .A(n9382), .B(n9295), .ZN(n9387) );
  XOR2_X1 U11756 ( .A(n9385), .B(n9387), .Z(n13903) );
  AND2_X1 U11757 ( .A1(n14028), .A2(n9278), .ZN(n9383) );
  AOI21_X1 U11758 ( .B1(n14404), .B2(n12066), .A(n9383), .ZN(n9390) );
  AOI22_X1 U11759 ( .A1(n14404), .A2(n9275), .B1(n12066), .B2(n14028), .ZN(
        n9384) );
  XNOR2_X1 U11760 ( .A(n9384), .B(n9295), .ZN(n9389) );
  XOR2_X1 U11761 ( .A(n9390), .B(n9389), .Z(n13964) );
  INV_X1 U11762 ( .A(n13964), .ZN(n9388) );
  INV_X1 U11763 ( .A(n9385), .ZN(n9386) );
  NAND2_X1 U11764 ( .A1(n9387), .A2(n9386), .ZN(n13959) );
  OR2_X1 U11765 ( .A1(n9388), .A2(n13959), .ZN(n13961) );
  INV_X1 U11766 ( .A(n9389), .ZN(n9392) );
  INV_X1 U11767 ( .A(n9390), .ZN(n9391) );
  NAND2_X1 U11768 ( .A1(n9392), .A2(n9391), .ZN(n9393) );
  AND2_X1 U11769 ( .A1(n13961), .A2(n9393), .ZN(n9394) );
  NAND2_X1 U11770 ( .A1(n13962), .A2(n9394), .ZN(n13913) );
  AOI22_X1 U11771 ( .A1(n14271), .A2(n9275), .B1(n12065), .B2(n14248), .ZN(
        n9395) );
  XNOR2_X1 U11772 ( .A(n9395), .B(n9295), .ZN(n9398) );
  AOI22_X1 U11773 ( .A1(n14271), .A2(n12061), .B1(n9278), .B2(n14248), .ZN(
        n9397) );
  XNOR2_X1 U11774 ( .A(n9398), .B(n9397), .ZN(n13914) );
  INV_X1 U11775 ( .A(n13914), .ZN(n9396) );
  NAND2_X1 U11776 ( .A1(n9398), .A2(n9397), .ZN(n9399) );
  AOI22_X1 U11777 ( .A1(n14394), .A2(n9275), .B1(n12065), .B2(n14027), .ZN(
        n9400) );
  XNOR2_X1 U11778 ( .A(n9400), .B(n9295), .ZN(n9405) );
  INV_X1 U11779 ( .A(n14394), .ZN(n14259) );
  OR2_X1 U11780 ( .A1(n14259), .A2(n9287), .ZN(n9402) );
  NAND2_X1 U11781 ( .A1(n14027), .A2(n9278), .ZN(n9401) );
  NAND2_X1 U11782 ( .A1(n9402), .A2(n9401), .ZN(n9403) );
  XNOR2_X1 U11783 ( .A(n9405), .B(n9403), .ZN(n13973) );
  INV_X1 U11784 ( .A(n9403), .ZN(n9404) );
  NAND2_X1 U11785 ( .A1(n9405), .A2(n9404), .ZN(n9406) );
  NAND2_X1 U11786 ( .A1(n14385), .A2(n9275), .ZN(n9408) );
  NAND2_X1 U11787 ( .A1(n14249), .A2(n12057), .ZN(n9407) );
  NAND2_X1 U11788 ( .A1(n9408), .A2(n9407), .ZN(n9409) );
  XNOR2_X1 U11789 ( .A(n9409), .B(n9295), .ZN(n9410) );
  AOI22_X1 U11790 ( .A1(n14385), .A2(n12061), .B1(n9278), .B2(n14249), .ZN(
        n9411) );
  XNOR2_X1 U11791 ( .A(n9410), .B(n9411), .ZN(n13896) );
  INV_X1 U11792 ( .A(n9410), .ZN(n9412) );
  NAND2_X1 U11793 ( .A1(n9412), .A2(n9411), .ZN(n9413) );
  NAND2_X1 U11794 ( .A1(n14377), .A2(n9275), .ZN(n9416) );
  NAND2_X1 U11795 ( .A1(n14026), .A2(n12057), .ZN(n9415) );
  NAND2_X1 U11796 ( .A1(n9416), .A2(n9415), .ZN(n9417) );
  XNOR2_X1 U11797 ( .A(n9417), .B(n9295), .ZN(n9418) );
  AOI22_X1 U11798 ( .A1(n14377), .A2(n12061), .B1(n9278), .B2(n14026), .ZN(
        n9419) );
  XNOR2_X1 U11799 ( .A(n9418), .B(n9419), .ZN(n13953) );
  INV_X1 U11800 ( .A(n9418), .ZN(n9420) );
  NAND2_X1 U11801 ( .A1(n9420), .A2(n9419), .ZN(n13922) );
  NAND2_X1 U11802 ( .A1(n14374), .A2(n9275), .ZN(n9422) );
  NAND2_X1 U11803 ( .A1(n14174), .A2(n12057), .ZN(n9421) );
  NAND2_X1 U11804 ( .A1(n9422), .A2(n9421), .ZN(n9423) );
  XNOR2_X1 U11805 ( .A(n9423), .B(n9295), .ZN(n9427) );
  INV_X1 U11806 ( .A(n9427), .ZN(n9424) );
  AOI22_X1 U11807 ( .A1(n14374), .A2(n12061), .B1(n9278), .B2(n14174), .ZN(
        n9426) );
  NAND2_X1 U11808 ( .A1(n9424), .A2(n9426), .ZN(n9425) );
  AND2_X1 U11809 ( .A1(n13922), .A2(n9425), .ZN(n12051) );
  INV_X1 U11810 ( .A(n9425), .ZN(n9428) );
  XNOR2_X1 U11811 ( .A(n9427), .B(n9426), .ZN(n13925) );
  OR2_X1 U11812 ( .A1(n9428), .A2(n13925), .ZN(n12053) );
  NAND2_X1 U11813 ( .A1(n14366), .A2(n9275), .ZN(n9430) );
  NAND2_X1 U11814 ( .A1(n14147), .A2(n12057), .ZN(n9429) );
  NAND2_X1 U11815 ( .A1(n9430), .A2(n9429), .ZN(n9431) );
  XNOR2_X1 U11816 ( .A(n9431), .B(n9295), .ZN(n12048) );
  AOI22_X1 U11817 ( .A1(n14366), .A2(n12061), .B1(n9278), .B2(n14147), .ZN(
        n12049) );
  XNOR2_X1 U11818 ( .A(n12048), .B(n12049), .ZN(n12054) );
  INV_X1 U11819 ( .A(n12054), .ZN(n9432) );
  NAND2_X1 U11820 ( .A1(n11882), .A2(P1_B_REG_SCAN_IN), .ZN(n9433) );
  MUX2_X1 U11821 ( .A(n9433), .B(P1_B_REG_SCAN_IN), .S(n9447), .Z(n9435) );
  INV_X1 U11822 ( .A(n12009), .ZN(n9434) );
  OR2_X1 U11823 ( .A1(n9653), .A2(P1_D_REG_1__SCAN_IN), .ZN(n9436) );
  NAND2_X1 U11824 ( .A1(n12009), .A2(n11882), .ZN(n9657) );
  NOR4_X1 U11825 ( .A1(P1_D_REG_4__SCAN_IN), .A2(P1_D_REG_5__SCAN_IN), .A3(
        P1_D_REG_6__SCAN_IN), .A4(P1_D_REG_7__SCAN_IN), .ZN(n9445) );
  NOR4_X1 U11826 ( .A1(P1_D_REG_8__SCAN_IN), .A2(P1_D_REG_9__SCAN_IN), .A3(
        P1_D_REG_10__SCAN_IN), .A4(P1_D_REG_11__SCAN_IN), .ZN(n9444) );
  OR4_X1 U11827 ( .A1(P1_D_REG_31__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_2__SCAN_IN), .A4(P1_D_REG_3__SCAN_IN), .ZN(n9442) );
  NOR4_X1 U11828 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_17__SCAN_IN), .A3(
        P1_D_REG_18__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n9440) );
  NOR4_X1 U11829 ( .A1(P1_D_REG_12__SCAN_IN), .A2(P1_D_REG_15__SCAN_IN), .A3(
        P1_D_REG_13__SCAN_IN), .A4(P1_D_REG_14__SCAN_IN), .ZN(n9439) );
  NOR4_X1 U11830 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_27__SCAN_IN), .A4(P1_D_REG_28__SCAN_IN), .ZN(n9438) );
  NOR4_X1 U11831 ( .A1(P1_D_REG_21__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_23__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n9437) );
  NAND4_X1 U11832 ( .A1(n9440), .A2(n9439), .A3(n9438), .A4(n9437), .ZN(n9441)
         );
  NOR4_X1 U11833 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        n9442), .A4(n9441), .ZN(n9443) );
  AND3_X1 U11834 ( .A1(n9445), .A2(n9444), .A3(n9443), .ZN(n9555) );
  AND2_X1 U11835 ( .A1(n9555), .A2(P1_D_REG_0__SCAN_IN), .ZN(n9446) );
  OR2_X1 U11836 ( .A1(n9653), .A2(n9446), .ZN(n9448) );
  INV_X1 U11837 ( .A(n9447), .ZN(n11817) );
  NAND2_X1 U11838 ( .A1(n11817), .A2(n12009), .ZN(n9654) );
  AND2_X1 U11839 ( .A1(n9448), .A2(n9654), .ZN(n9562) );
  INV_X1 U11840 ( .A(n9666), .ZN(n9451) );
  AND2_X1 U11841 ( .A1(n11614), .A2(n9449), .ZN(n9450) );
  NAND2_X1 U11842 ( .A1(n9451), .A2(n14843), .ZN(n9452) );
  NOR2_X1 U11843 ( .A1(n9457), .A2(n9452), .ZN(n9453) );
  INV_X1 U11844 ( .A(n9454), .ZN(n9455) );
  NAND2_X1 U11845 ( .A1(n9455), .A2(n9915), .ZN(n10601) );
  NOR2_X1 U11846 ( .A1(n9457), .A2(n10601), .ZN(n9456) );
  NAND2_X1 U11847 ( .A1(n9463), .A2(n9456), .ZN(n9458) );
  INV_X1 U11848 ( .A(n9463), .ZN(n9459) );
  NAND2_X1 U11849 ( .A1(n9459), .A2(n9553), .ZN(n10135) );
  NAND3_X1 U11850 ( .A1(n10135), .A2(n9460), .A3(n9265), .ZN(n9461) );
  NAND2_X1 U11851 ( .A1(n9461), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9462) );
  NOR2_X1 U11852 ( .A1(n13989), .A2(n14178), .ZN(n9467) );
  NAND2_X1 U11853 ( .A1(n13999), .A2(n14321), .ZN(n14013) );
  AOI22_X1 U11854 ( .A1(n14011), .A2(n14174), .B1(P1_REG3_REG_26__SCAN_IN), 
        .B2(P1_U3086), .ZN(n9464) );
  OAI21_X1 U11855 ( .B1(n9465), .B2(n14013), .A(n9464), .ZN(n9466) );
  AOI211_X1 U11856 ( .C1(n14366), .C2(n14018), .A(n9467), .B(n9466), .ZN(n9468) );
  INV_X1 U11857 ( .A(n14374), .ZN(n14451) );
  NAND2_X1 U11858 ( .A1(n10177), .A2(n10184), .ZN(n9469) );
  NAND2_X1 U11859 ( .A1(n10510), .A2(n6691), .ZN(n9470) );
  NAND2_X1 U11860 ( .A1(n10621), .A2(n9470), .ZN(n10504) );
  NAND2_X1 U11861 ( .A1(n10504), .A2(n10503), .ZN(n10502) );
  NAND2_X1 U11862 ( .A1(n9471), .A2(n10518), .ZN(n9472) );
  NAND2_X1 U11863 ( .A1(n10502), .A2(n9472), .ZN(n10825) );
  NAND2_X1 U11864 ( .A1(n10900), .A2(n14839), .ZN(n9473) );
  NAND2_X1 U11865 ( .A1(n10823), .A2(n9473), .ZN(n10657) );
  NAND2_X1 U11866 ( .A1(n10657), .A2(n10656), .ZN(n10655) );
  OR2_X1 U11867 ( .A1(n14040), .A2(n10897), .ZN(n9474) );
  NAND2_X1 U11868 ( .A1(n10655), .A2(n9474), .ZN(n10643) );
  NAND2_X1 U11869 ( .A1(n10643), .A2(n10645), .ZN(n10642) );
  OR2_X1 U11870 ( .A1(n14002), .A2(n14039), .ZN(n9475) );
  NAND2_X1 U11871 ( .A1(n10642), .A2(n9475), .ZN(n11141) );
  OR2_X1 U11872 ( .A1(n11200), .A2(n14038), .ZN(n9476) );
  OR2_X1 U11873 ( .A1(n11471), .A2(n14037), .ZN(n9477) );
  NAND2_X1 U11874 ( .A1(n11361), .A2(n11360), .ZN(n11359) );
  OR2_X1 U11875 ( .A1(n11663), .A2(n14035), .ZN(n9478) );
  OR2_X1 U11876 ( .A1(n11571), .A2(n14034), .ZN(n9479) );
  OR2_X1 U11877 ( .A1(n11736), .A2(n14032), .ZN(n9480) );
  NAND2_X1 U11878 ( .A1(n13892), .A2(n14031), .ZN(n9482) );
  OR2_X1 U11879 ( .A1(n14019), .A2(n14030), .ZN(n9483) );
  OR2_X1 U11880 ( .A1(n14425), .A2(n12038), .ZN(n9484) );
  OR2_X1 U11881 ( .A1(n14414), .A2(n14029), .ZN(n9485) );
  NAND2_X1 U11882 ( .A1(n14414), .A2(n14029), .ZN(n9486) );
  INV_X1 U11883 ( .A(n14302), .ZN(n9488) );
  OR2_X1 U11884 ( .A1(n14409), .A2(n14322), .ZN(n9489) );
  INV_X1 U11885 ( .A(n14266), .ZN(n9490) );
  OR2_X1 U11886 ( .A1(n14271), .A2(n14248), .ZN(n9491) );
  NAND2_X1 U11887 ( .A1(n14253), .A2(n14252), .ZN(n14251) );
  OR2_X1 U11888 ( .A1(n14394), .A2(n14027), .ZN(n9492) );
  NAND2_X1 U11889 ( .A1(n14385), .A2(n14249), .ZN(n14204) );
  AND2_X1 U11890 ( .A1(n14210), .A2(n14204), .ZN(n9494) );
  OR2_X1 U11891 ( .A1(n14377), .A2(n14026), .ZN(n9495) );
  INV_X1 U11892 ( .A(n14158), .ZN(n9496) );
  NAND2_X1 U11893 ( .A1(n9496), .A2(n9465), .ZN(n9497) );
  XNOR2_X1 U11894 ( .A(n9498), .B(n9543), .ZN(n12560) );
  OAI21_X1 U11895 ( .B1(n9499), .B2(n9915), .A(n12108), .ZN(n9500) );
  AND2_X1 U11896 ( .A1(n11493), .A2(n9502), .ZN(n9503) );
  NAND2_X1 U11897 ( .A1(n9915), .A2(n9503), .ZN(n10515) );
  NAND2_X1 U11898 ( .A1(n9504), .A2(n8239), .ZN(n10610) );
  NAND2_X1 U11899 ( .A1(n10611), .A2(n10610), .ZN(n10609) );
  NAND2_X1 U11900 ( .A1(n10609), .A2(n9505), .ZN(n10508) );
  NAND2_X1 U11901 ( .A1(n10508), .A2(n10509), .ZN(n10506) );
  NAND2_X1 U11902 ( .A1(n10506), .A2(n9506), .ZN(n10827) );
  NAND2_X1 U11903 ( .A1(n10826), .A2(n9507), .ZN(n10661) );
  NAND2_X1 U11904 ( .A1(n10661), .A2(n10660), .ZN(n10659) );
  NAND2_X1 U11905 ( .A1(n10897), .A2(n9508), .ZN(n9509) );
  NAND2_X1 U11906 ( .A1(n10659), .A2(n9509), .ZN(n10646) );
  OR2_X1 U11907 ( .A1(n14002), .A2(n10662), .ZN(n9510) );
  NAND2_X1 U11908 ( .A1(n10646), .A2(n9510), .ZN(n9512) );
  NAND2_X1 U11909 ( .A1(n14002), .A2(n10662), .ZN(n9511) );
  NAND2_X1 U11910 ( .A1(n9512), .A2(n9511), .ZN(n11147) );
  AND2_X1 U11911 ( .A1(n11200), .A2(n11241), .ZN(n9514) );
  OR2_X1 U11912 ( .A1(n11200), .A2(n11241), .ZN(n9513) );
  INV_X1 U11913 ( .A(n11231), .ZN(n11239) );
  OR2_X1 U11914 ( .A1(n11471), .A2(n9515), .ZN(n9516) );
  NAND2_X1 U11915 ( .A1(n11767), .A2(n11465), .ZN(n9517) );
  NAND2_X1 U11916 ( .A1(n11159), .A2(n9517), .ZN(n11356) );
  OR2_X1 U11917 ( .A1(n11663), .A2(n11418), .ZN(n9520) );
  INV_X1 U11918 ( .A(n11413), .ZN(n11416) );
  INV_X1 U11919 ( .A(n11477), .ZN(n11480) );
  OR2_X1 U11920 ( .A1(n11488), .A2(n11824), .ZN(n9521) );
  NAND2_X1 U11921 ( .A1(n9522), .A2(n9521), .ZN(n11601) );
  INV_X1 U11922 ( .A(n11599), .ZN(n11602) );
  NAND2_X1 U11923 ( .A1(n11601), .A2(n11602), .ZN(n9524) );
  OR2_X1 U11924 ( .A1(n11736), .A2(n11898), .ZN(n9523) );
  NAND2_X1 U11925 ( .A1(n9524), .A2(n9523), .ZN(n11648) );
  NAND2_X1 U11926 ( .A1(n11648), .A2(n11649), .ZN(n9526) );
  AND2_X1 U11927 ( .A1(n14425), .A2(n14014), .ZN(n12034) );
  NAND2_X1 U11928 ( .A1(n11831), .A2(n9528), .ZN(n12036) );
  NAND2_X1 U11929 ( .A1(n12036), .A2(n9529), .ZN(n14318) );
  NAND2_X1 U11930 ( .A1(n14318), .A2(n14332), .ZN(n9531) );
  INV_X1 U11931 ( .A(n14029), .ZN(n13906) );
  OR2_X1 U11932 ( .A1(n14414), .A2(n13906), .ZN(n9530) );
  INV_X1 U11933 ( .A(n14280), .ZN(n14283) );
  INV_X1 U11934 ( .A(n14028), .ZN(n14264) );
  INV_X1 U11935 ( .A(n14248), .ZN(n14288) );
  NOR2_X1 U11936 ( .A1(n14271), .A2(n14288), .ZN(n9533) );
  INV_X1 U11937 ( .A(n14252), .ZN(n14246) );
  NAND2_X1 U11938 ( .A1(n14247), .A2(n14246), .ZN(n9535) );
  NAND2_X1 U11939 ( .A1(n14394), .A2(n14265), .ZN(n9534) );
  NAND2_X1 U11940 ( .A1(n9535), .A2(n9534), .ZN(n14228) );
  NAND2_X1 U11941 ( .A1(n14228), .A2(n14233), .ZN(n14230) );
  INV_X1 U11942 ( .A(n14249), .ZN(n9536) );
  NAND2_X1 U11943 ( .A1(n14385), .A2(n9536), .ZN(n9537) );
  NAND2_X1 U11944 ( .A1(n14230), .A2(n9537), .ZN(n14211) );
  INV_X1 U11945 ( .A(n14211), .ZN(n9538) );
  NAND2_X2 U11946 ( .A1(n9538), .A2(n14205), .ZN(n14215) );
  INV_X1 U11947 ( .A(n14026), .ZN(n9539) );
  OR2_X1 U11948 ( .A1(n14377), .A2(n9539), .ZN(n9540) );
  INV_X1 U11949 ( .A(n14366), .ZN(n14180) );
  NOR2_X1 U11950 ( .A1(n14180), .A2(n14147), .ZN(n14149) );
  NAND2_X1 U11951 ( .A1(n14130), .A2(n14135), .ZN(n14129) );
  NAND2_X1 U11952 ( .A1(n14129), .A2(n9542), .ZN(n9544) );
  XNOR2_X1 U11953 ( .A(n9544), .B(n6669), .ZN(n9547) );
  OR2_X1 U11954 ( .A1(n9915), .A2(n12108), .ZN(n9546) );
  NOR2_X1 U11955 ( .A1(n14345), .A2(n9548), .ZN(n10614) );
  NAND2_X1 U11956 ( .A1(n10614), .A2(n6691), .ZN(n10613) );
  OR2_X1 U11957 ( .A1(n10613), .A2(n10605), .ZN(n10831) );
  INV_X1 U11958 ( .A(n11471), .ZN(n14844) );
  AND2_X2 U11959 ( .A1(n11235), .A2(n14844), .ZN(n11233) );
  NAND2_X1 U11960 ( .A1(n12031), .A2(n11485), .ZN(n11642) );
  INV_X1 U11961 ( .A(n14138), .ZN(n14356) );
  AOI21_X1 U11962 ( .B1(n14136), .B2(n12555), .A(n14326), .ZN(n9550) );
  NAND2_X1 U11963 ( .A1(n9550), .A2(n12082), .ZN(n12558) );
  NAND2_X1 U11964 ( .A1(n9745), .A2(P1_B_REG_SCAN_IN), .ZN(n9551) );
  AND2_X1 U11965 ( .A1(n14321), .A2(n9551), .ZN(n12084) );
  NAND2_X1 U11966 ( .A1(n12084), .A2(n14025), .ZN(n12552) );
  OAI21_X1 U11967 ( .B1(n9653), .B2(P1_D_REG_0__SCAN_IN), .A(n9654), .ZN(n9557) );
  OR2_X1 U11968 ( .A1(n9653), .A2(n9555), .ZN(n9556) );
  NAND2_X1 U11969 ( .A1(n9557), .A2(n9556), .ZN(n10595) );
  INV_X1 U11970 ( .A(n10593), .ZN(n9558) );
  NOR2_X1 U11971 ( .A1(n10595), .A2(n9558), .ZN(n9559) );
  NAND2_X1 U11972 ( .A1(n14849), .A2(n14426), .ZN(n14468) );
  NAND2_X1 U11973 ( .A1(n9561), .A2(n7447), .ZN(P1_U3525) );
  AND2_X1 U11974 ( .A1(n9562), .A2(n10593), .ZN(n9563) );
  NAND2_X1 U11975 ( .A1(n9566), .A2(n7448), .ZN(P1_U3557) );
  INV_X1 U11976 ( .A(n9658), .ZN(n9569) );
  OR2_X2 U11977 ( .A1(n9569), .A2(n9265), .ZN(n14044) );
  INV_X2 U11978 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  OAI222_X1 U11979 ( .A1(P2_U3088), .A2(n9723), .B1(n13873), .B2(n9628), .C1(
        n9600), .C2(n13870), .ZN(P2_U3325) );
  OAI222_X1 U11980 ( .A1(P2_U3088), .A2(n14857), .B1(n13873), .B2(n9631), .C1(
        n9572), .C2(n13870), .ZN(P2_U3326) );
  INV_X1 U11981 ( .A(n9760), .ZN(n9771) );
  INV_X1 U11982 ( .A(n9570), .ZN(n9630) );
  INV_X1 U11983 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n9603) );
  OAI222_X1 U11984 ( .A1(P2_U3088), .A2(n9771), .B1(n13873), .B2(n9630), .C1(
        n9603), .C2(n13870), .ZN(P2_U3324) );
  INV_X2 U11985 ( .A(n13320), .ZN(n13333) );
  INV_X1 U11986 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n9571) );
  AND2_X1 U11987 ( .A1(n9571), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n9611) );
  NAND2_X1 U11988 ( .A1(n9592), .A2(n9611), .ZN(n9574) );
  NAND2_X1 U11989 ( .A1(n9572), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n9573) );
  NAND2_X1 U11990 ( .A1(n9574), .A2(n9573), .ZN(n9602) );
  INV_X1 U11991 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n9627) );
  NAND2_X1 U11992 ( .A1(n9627), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n9575) );
  NAND2_X1 U11993 ( .A1(n9602), .A2(n9575), .ZN(n9577) );
  NAND2_X1 U11994 ( .A1(n9600), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n9576) );
  AND2_X1 U11995 ( .A1(n9603), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n9578) );
  INV_X1 U11996 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n9629) );
  NAND2_X1 U11997 ( .A1(n9629), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n9579) );
  INV_X1 U11998 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n9626) );
  NAND2_X1 U11999 ( .A1(n9626), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n9580) );
  XNOR2_X1 U12000 ( .A(n9584), .B(n9583), .ZN(n10922) );
  INV_X2 U12001 ( .A(n12092), .ZN(n13335) );
  INV_X1 U12002 ( .A(SI_5_), .ZN(n10921) );
  OAI222_X1 U12003 ( .A1(n13333), .A2(n10922), .B1(n13335), .B2(n10921), .C1(
        n15138), .C2(P3_U3151), .ZN(P3_U3290) );
  INV_X1 U12004 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n9624) );
  NAND2_X1 U12005 ( .A1(n9624), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n9585) );
  NAND2_X1 U12006 ( .A1(n9632), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n9588) );
  INV_X1 U12007 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n9634) );
  NAND2_X1 U12008 ( .A1(n9634), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n9587) );
  NAND2_X1 U12009 ( .A1(n9588), .A2(n9587), .ZN(n9607) );
  XNOR2_X1 U12010 ( .A(n9637), .B(P2_DATAO_REG_7__SCAN_IN), .ZN(n9616) );
  XNOR2_X1 U12011 ( .A(n9646), .B(P2_DATAO_REG_8__SCAN_IN), .ZN(n9589) );
  XNOR2_X1 U12012 ( .A(n9621), .B(n9589), .ZN(n11205) );
  INV_X1 U12013 ( .A(n11205), .ZN(n9591) );
  INV_X1 U12014 ( .A(SI_8_), .ZN(n9590) );
  OAI222_X1 U12015 ( .A1(n13333), .A2(n9591), .B1(n13335), .B2(n9590), .C1(
        n11206), .C2(P3_U3151), .ZN(P3_U3287) );
  INV_X1 U12016 ( .A(SI_1_), .ZN(n9594) );
  XNOR2_X1 U12017 ( .A(n9592), .B(n9611), .ZN(n10284) );
  INV_X1 U12018 ( .A(n10284), .ZN(n9593) );
  XNOR2_X1 U12019 ( .A(n9596), .B(n9595), .ZN(n10797) );
  INV_X1 U12020 ( .A(SI_4_), .ZN(n10796) );
  OAI222_X1 U12021 ( .A1(n13333), .A2(n10797), .B1(n13335), .B2(n10796), .C1(
        n9597), .C2(P3_U3151), .ZN(P3_U3291) );
  INV_X1 U12022 ( .A(n9699), .ZN(n14869) );
  INV_X1 U12023 ( .A(n9598), .ZN(n9625) );
  INV_X1 U12024 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n9599) );
  OAI222_X1 U12025 ( .A1(P2_U3088), .A2(n14869), .B1(n13873), .B2(n9625), .C1(
        n9599), .C2(n13870), .ZN(P2_U3323) );
  XNOR2_X1 U12026 ( .A(n9600), .B(P2_DATAO_REG_2__SCAN_IN), .ZN(n9601) );
  XNOR2_X1 U12027 ( .A(n9602), .B(n9601), .ZN(n10448) );
  INV_X1 U12028 ( .A(SI_2_), .ZN(n10447) );
  OAI222_X1 U12029 ( .A1(n6496), .A2(P3_U3151), .B1(n13333), .B2(n10448), .C1(
        n10447), .C2(n13335), .ZN(P3_U3293) );
  XNOR2_X1 U12030 ( .A(n9603), .B(P2_DATAO_REG_3__SCAN_IN), .ZN(n9604) );
  XNOR2_X1 U12031 ( .A(n9605), .B(n9604), .ZN(n10548) );
  INV_X1 U12032 ( .A(SI_3_), .ZN(n10547) );
  OAI222_X1 U12033 ( .A1(n9606), .A2(P3_U3151), .B1(n13333), .B2(n10548), .C1(
        n10547), .C2(n13335), .ZN(P3_U3292) );
  XNOR2_X1 U12034 ( .A(n9608), .B(n9607), .ZN(n11071) );
  INV_X1 U12035 ( .A(n11071), .ZN(n9610) );
  INV_X1 U12036 ( .A(SI_6_), .ZN(n9609) );
  OAI222_X1 U12037 ( .A1(n11074), .A2(P3_U3151), .B1(n13333), .B2(n9610), .C1(
        n9609), .C2(n13335), .ZN(P3_U3289) );
  INV_X1 U12038 ( .A(n9611), .ZN(n9614) );
  NAND2_X1 U12039 ( .A1(n9612), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n9613) );
  NAND2_X1 U12040 ( .A1(n9614), .A2(n9613), .ZN(n10188) );
  INV_X1 U12041 ( .A(n10188), .ZN(n9615) );
  OAI222_X1 U12042 ( .A1(n15105), .A2(P3_U3151), .B1(n13333), .B2(n9615), .C1(
        n13279), .C2(n13335), .ZN(P3_U3295) );
  XNOR2_X1 U12043 ( .A(n9617), .B(n9616), .ZN(n11082) );
  INV_X1 U12044 ( .A(SI_7_), .ZN(n11083) );
  OAI222_X1 U12045 ( .A1(n9618), .A2(P3_U3151), .B1(n13333), .B2(n11082), .C1(
        n11083), .C2(n13335), .ZN(P3_U3288) );
  INV_X1 U12046 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n9620) );
  INV_X1 U12047 ( .A(n9619), .ZN(n9623) );
  OAI222_X1 U12048 ( .A1(n13870), .A2(n9620), .B1(n13873), .B2(n9623), .C1(
        P2_U3088), .C2(n9711), .ZN(P2_U3322) );
  XNOR2_X1 U12049 ( .A(n9651), .B(P2_DATAO_REG_9__SCAN_IN), .ZN(n9622) );
  XNOR2_X1 U12050 ( .A(n9636), .B(n9622), .ZN(n11304) );
  INV_X1 U12051 ( .A(SI_9_), .ZN(n11305) );
  OAI222_X1 U12052 ( .A1(n10860), .A2(P3_U3151), .B1(n13333), .B2(n11304), 
        .C1(n11305), .C2(n13335), .ZN(P3_U3286) );
  INV_X2 U12053 ( .A(n14473), .ZN(n14478) );
  AND2_X1 U12054 ( .A1(n8621), .A2(P1_U3086), .ZN(n11884) );
  INV_X2 U12055 ( .A(n11884), .ZN(n14480) );
  OAI222_X1 U12056 ( .A1(n14478), .A2(n9624), .B1(n14480), .B2(n9623), .C1(
        P1_U3086), .C2(n9884), .ZN(P1_U3350) );
  INV_X1 U12057 ( .A(n9799), .ZN(n14794) );
  OAI222_X1 U12058 ( .A1(n14478), .A2(n9626), .B1(n14480), .B2(n9625), .C1(
        n14794), .C2(P1_U3086), .ZN(P1_U3351) );
  INV_X1 U12059 ( .A(n14073), .ZN(n9788) );
  OAI222_X1 U12060 ( .A1(P1_U3086), .A2(n9788), .B1(n14480), .B2(n9628), .C1(
        n9627), .C2(n14478), .ZN(P1_U3353) );
  OAI222_X1 U12061 ( .A1(P1_U3086), .A2(n14090), .B1(n14480), .B2(n9630), .C1(
        n9629), .C2(n14478), .ZN(P1_U3352) );
  OAI222_X1 U12062 ( .A1(P1_U3086), .A2(n7526), .B1(n14480), .B2(n9631), .C1(
        n7499), .C2(n14478), .ZN(P1_U3354) );
  INV_X1 U12063 ( .A(n9847), .ZN(n9740) );
  OAI222_X1 U12064 ( .A1(P2_U3088), .A2(n9740), .B1(n13873), .B2(n9633), .C1(
        n9632), .C2(n13870), .ZN(P2_U3321) );
  INV_X1 U12065 ( .A(n9885), .ZN(n9950) );
  OAI222_X1 U12066 ( .A1(n14478), .A2(n9634), .B1(n14480), .B2(n9633), .C1(
        n9950), .C2(P1_U3086), .ZN(P1_U3349) );
  AND2_X1 U12067 ( .A1(n9651), .A2(P2_DATAO_REG_9__SCAN_IN), .ZN(n9635) );
  XNOR2_X1 U12068 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .ZN(n9640) );
  XNOR2_X1 U12069 ( .A(n9641), .B(n9640), .ZN(n11391) );
  OAI222_X1 U12070 ( .A1(n13333), .A2(n11391), .B1(n13335), .B2(n11394), .C1(
        n11393), .C2(P3_U3151), .ZN(P3_U3285) );
  INV_X1 U12071 ( .A(n13456), .ZN(n13449) );
  OAI222_X1 U12072 ( .A1(P2_U3088), .A2(n13449), .B1(n13873), .B2(n9639), .C1(
        n9637), .C2(n13870), .ZN(P2_U3320) );
  INV_X1 U12073 ( .A(n10011), .ZN(n10020) );
  OAI222_X1 U12074 ( .A1(n14478), .A2(n7136), .B1(n14480), .B2(n9639), .C1(
        n10020), .C2(P1_U3086), .ZN(P1_U3348) );
  NAND2_X1 U12075 ( .A1(n9778), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n9642) );
  NAND2_X1 U12076 ( .A1(n9936), .A2(P2_DATAO_REG_11__SCAN_IN), .ZN(n9662) );
  INV_X1 U12077 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n9933) );
  NAND2_X1 U12078 ( .A1(n9933), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n9644) );
  XNOR2_X1 U12079 ( .A(n9661), .B(n6642), .ZN(n11528) );
  OAI222_X1 U12080 ( .A1(n11529), .A2(P3_U3151), .B1(n13333), .B2(n11528), 
        .C1(n11530), .C2(n13335), .ZN(P3_U3284) );
  INV_X1 U12081 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n9645) );
  INV_X1 U12082 ( .A(n10023), .ZN(n10063) );
  OAI222_X1 U12083 ( .A1(n14478), .A2(n9645), .B1(n14480), .B2(n9647), .C1(
        n10063), .C2(P1_U3086), .ZN(P1_U3347) );
  INV_X1 U12084 ( .A(n13472), .ZN(n9648) );
  OAI222_X1 U12085 ( .A1(P2_U3088), .A2(n9648), .B1(n13873), .B2(n9647), .C1(
        n9646), .C2(n13870), .ZN(P2_U3319) );
  INV_X1 U12086 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n9650) );
  INV_X1 U12087 ( .A(n10042), .ZN(n9649) );
  OAI222_X1 U12088 ( .A1(n14478), .A2(n9650), .B1(n14480), .B2(n9652), .C1(
        n9649), .C2(P1_U3086), .ZN(P1_U3346) );
  INV_X1 U12089 ( .A(n9902), .ZN(n9871) );
  OAI222_X1 U12090 ( .A1(P2_U3088), .A2(n9871), .B1(n13873), .B2(n9652), .C1(
        n9651), .C2(n13870), .ZN(P2_U3318) );
  INV_X1 U12091 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n9656) );
  INV_X1 U12092 ( .A(n9654), .ZN(n9655) );
  AOI22_X1 U12093 ( .A1(n14831), .A2(n9656), .B1(n9658), .B2(n9655), .ZN(
        P1_U3445) );
  INV_X1 U12094 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n9660) );
  INV_X1 U12095 ( .A(n9657), .ZN(n9659) );
  AOI22_X1 U12096 ( .A1(n14831), .A2(n9660), .B1(n9659), .B2(n9658), .ZN(
        P1_U3446) );
  XNOR2_X1 U12097 ( .A(n6512), .B(n6641), .ZN(n11681) );
  INV_X1 U12098 ( .A(n11516), .ZN(n11682) );
  AOI222_X1 U12099 ( .A1(n11681), .A2(n13320), .B1(SI_12_), .B2(n12092), .C1(
        P3_STATE_REG_SCAN_IN), .C2(n11682), .ZN(n9663) );
  INV_X1 U12100 ( .A(n9663), .ZN(P3_U3283) );
  NAND2_X1 U12101 ( .A1(n9666), .A2(n9665), .ZN(n9668) );
  NAND2_X1 U12102 ( .A1(n9668), .A2(n9667), .ZN(n9742) );
  NAND2_X1 U12103 ( .A1(n9744), .A2(n9742), .ZN(n14815) );
  INV_X1 U12104 ( .A(n14815), .ZN(n14088) );
  NOR2_X1 U12105 ( .A1(n14088), .A2(P1_U4016), .ZN(P1_U3085) );
  OAI21_X1 U12106 ( .B1(n9671), .B2(n9987), .A(n9669), .ZN(n9670) );
  OAI21_X1 U12107 ( .B1(n9983), .B2(n9671), .A(n9670), .ZN(n9689) );
  NAND2_X1 U12108 ( .A1(n9689), .A2(n9251), .ZN(n14870) );
  OR2_X1 U12109 ( .A1(n9251), .A2(P2_U3088), .ZN(n12079) );
  INV_X1 U12110 ( .A(n13526), .ZN(n9672) );
  NOR2_X1 U12111 ( .A1(n12079), .A2(n9672), .ZN(n9673) );
  NAND2_X1 U12112 ( .A1(n9689), .A2(n9673), .ZN(n13511) );
  INV_X1 U12113 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n9674) );
  MUX2_X1 U12114 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n9674), .S(n9760), .Z(n9680)
         );
  INV_X1 U12115 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n9675) );
  MUX2_X1 U12116 ( .A(n9675), .B(P2_REG1_REG_2__SCAN_IN), .S(n9723), .Z(n9678)
         );
  INV_X1 U12117 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n9676) );
  MUX2_X1 U12118 ( .A(n9676), .B(P2_REG1_REG_1__SCAN_IN), .S(n14857), .Z(
        n14863) );
  AND2_X1 U12119 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n14864) );
  NAND2_X1 U12120 ( .A1(n14863), .A2(n14864), .ZN(n14862) );
  NAND2_X1 U12121 ( .A1(n8620), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n9712) );
  NAND2_X1 U12122 ( .A1(n14862), .A2(n9712), .ZN(n9677) );
  NAND2_X1 U12123 ( .A1(n9678), .A2(n9677), .ZN(n9762) );
  OR2_X1 U12124 ( .A1(n9723), .A2(n9675), .ZN(n9761) );
  NAND2_X1 U12125 ( .A1(n9762), .A2(n9761), .ZN(n9679) );
  NAND2_X1 U12126 ( .A1(n9680), .A2(n9679), .ZN(n9765) );
  NAND2_X1 U12127 ( .A1(n9760), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n9681) );
  NAND2_X1 U12128 ( .A1(n9765), .A2(n9681), .ZN(n14877) );
  INV_X1 U12129 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n15090) );
  MUX2_X1 U12130 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n15090), .S(n9699), .Z(
        n14876) );
  NAND2_X1 U12131 ( .A1(n14877), .A2(n14876), .ZN(n14875) );
  NAND2_X1 U12132 ( .A1(n9699), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n9686) );
  NAND2_X1 U12133 ( .A1(n14875), .A2(n9686), .ZN(n9684) );
  INV_X1 U12134 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n9682) );
  MUX2_X1 U12135 ( .A(n9682), .B(P2_REG1_REG_5__SCAN_IN), .S(n9711), .Z(n9683)
         );
  NAND2_X1 U12136 ( .A1(n9684), .A2(n9683), .ZN(n9725) );
  MUX2_X1 U12137 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n9682), .S(n9711), .Z(n9685)
         );
  NAND3_X1 U12138 ( .A1(n14875), .A2(n9686), .A3(n9685), .ZN(n9687) );
  AND3_X1 U12139 ( .A1(n14956), .A2(n9725), .A3(n9687), .ZN(n9709) );
  INV_X1 U12140 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n9707) );
  NOR2_X1 U12141 ( .A1(n12079), .A2(n13526), .ZN(n9688) );
  INV_X1 U12142 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n9690) );
  MUX2_X1 U12143 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n9690), .S(n9760), .Z(n9696)
         );
  NAND2_X1 U12144 ( .A1(n8620), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n9692) );
  INV_X1 U12145 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n10985) );
  NAND2_X1 U12146 ( .A1(n14857), .A2(n10985), .ZN(n9691) );
  AND2_X1 U12147 ( .A1(n9692), .A2(n9691), .ZN(n14861) );
  AND2_X1 U12148 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n14860) );
  NAND2_X1 U12149 ( .A1(n14861), .A2(n14860), .ZN(n14859) );
  NAND2_X1 U12150 ( .A1(n14859), .A2(n9692), .ZN(n9718) );
  XNOR2_X1 U12151 ( .A(n9723), .B(P2_REG2_REG_2__SCAN_IN), .ZN(n9717) );
  NAND2_X1 U12152 ( .A1(n9718), .A2(n9717), .ZN(n9695) );
  INV_X1 U12153 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n9693) );
  OR2_X1 U12154 ( .A1(n9723), .A2(n9693), .ZN(n9694) );
  NAND2_X1 U12155 ( .A1(n9695), .A2(n9694), .ZN(n9755) );
  NAND2_X1 U12156 ( .A1(n9696), .A2(n9755), .ZN(n9756) );
  NAND2_X1 U12157 ( .A1(n9760), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n9697) );
  NAND2_X1 U12158 ( .A1(n9756), .A2(n9697), .ZN(n14874) );
  INV_X1 U12159 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n9698) );
  MUX2_X1 U12160 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n9698), .S(n9699), .Z(n14873) );
  NAND2_X1 U12161 ( .A1(n14874), .A2(n14873), .ZN(n14872) );
  NAND2_X1 U12162 ( .A1(n9699), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n9704) );
  NAND2_X1 U12163 ( .A1(n14872), .A2(n9704), .ZN(n9702) );
  INV_X1 U12164 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n9700) );
  MUX2_X1 U12165 ( .A(n9700), .B(P2_REG2_REG_5__SCAN_IN), .S(n9711), .Z(n9701)
         );
  NAND2_X1 U12166 ( .A1(n9702), .A2(n9701), .ZN(n9736) );
  MUX2_X1 U12167 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n9700), .S(n9711), .Z(n9703)
         );
  NAND3_X1 U12168 ( .A1(n14872), .A2(n9704), .A3(n9703), .ZN(n9705) );
  NAND3_X1 U12169 ( .A1(n14961), .A2(n9736), .A3(n9705), .ZN(n9706) );
  OAI21_X1 U12170 ( .B1(n9707), .B2(n14901), .A(n9706), .ZN(n9708) );
  AND2_X1 U12171 ( .A1(P2_U3088), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n10276) );
  NOR3_X1 U12172 ( .A1(n9709), .A2(n9708), .A3(n10276), .ZN(n9710) );
  OAI21_X1 U12173 ( .B1(n9711), .B2(n14894), .A(n9710), .ZN(P2_U3219) );
  INV_X1 U12174 ( .A(n14901), .ZN(n14954) );
  MUX2_X1 U12175 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n9675), .S(n9723), .Z(n9713)
         );
  NAND3_X1 U12176 ( .A1(n9713), .A2(n14862), .A3(n9712), .ZN(n9714) );
  NAND2_X1 U12177 ( .A1(n9762), .A2(n9714), .ZN(n9716) );
  INV_X1 U12178 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n9715) );
  OAI22_X1 U12179 ( .A1(n13511), .A2(n9716), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9715), .ZN(n9721) );
  INV_X1 U12180 ( .A(n14961), .ZN(n10113) );
  XNOR2_X1 U12181 ( .A(n9718), .B(n9717), .ZN(n9719) );
  NOR2_X1 U12182 ( .A1(n10113), .A2(n9719), .ZN(n9720) );
  AOI211_X1 U12183 ( .C1(n14954), .C2(P2_ADDR_REG_2__SCAN_IN), .A(n9721), .B(
        n9720), .ZN(n9722) );
  OAI21_X1 U12184 ( .B1(n9723), .B2(n14894), .A(n9722), .ZN(P2_U3216) );
  NAND2_X1 U12185 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3088), .ZN(n10392) );
  NAND2_X1 U12186 ( .A1(n9731), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n9724) );
  NAND2_X1 U12187 ( .A1(n9725), .A2(n9724), .ZN(n9728) );
  INV_X1 U12188 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n9726) );
  MUX2_X1 U12189 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n9726), .S(n9847), .Z(n9727)
         );
  NAND2_X1 U12190 ( .A1(n9728), .A2(n9727), .ZN(n13454) );
  OAI211_X1 U12191 ( .C1(n9728), .C2(n9727), .A(n14956), .B(n13454), .ZN(n9729) );
  NAND2_X1 U12192 ( .A1(n10392), .A2(n9729), .ZN(n9730) );
  AOI21_X1 U12193 ( .B1(n14954), .B2(P2_ADDR_REG_6__SCAN_IN), .A(n9730), .ZN(
        n9739) );
  NAND2_X1 U12194 ( .A1(n9731), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n9735) );
  NAND2_X1 U12195 ( .A1(n9736), .A2(n9735), .ZN(n9733) );
  INV_X1 U12196 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n10887) );
  MUX2_X1 U12197 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n10887), .S(n9847), .Z(n9732) );
  NAND2_X1 U12198 ( .A1(n9733), .A2(n9732), .ZN(n13459) );
  MUX2_X1 U12199 ( .A(n10887), .B(P2_REG2_REG_6__SCAN_IN), .S(n9847), .Z(n9734) );
  NAND3_X1 U12200 ( .A1(n9736), .A2(n9735), .A3(n9734), .ZN(n9737) );
  NAND3_X1 U12201 ( .A1(n14961), .A2(n13459), .A3(n9737), .ZN(n9738) );
  OAI211_X1 U12202 ( .C1(n14894), .C2(n9740), .A(n9739), .B(n9738), .ZN(
        P2_U3220) );
  NAND2_X1 U12203 ( .A1(P1_U4016), .A2(n12038), .ZN(n9741) );
  OAI21_X1 U12204 ( .B1(P1_U4016), .B2(n7884), .A(n9741), .ZN(P1_U3576) );
  INV_X1 U12205 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n9754) );
  INV_X1 U12206 ( .A(n9742), .ZN(n9743) );
  AND2_X1 U12207 ( .A1(n9744), .A2(n9743), .ZN(n9794) );
  INV_X1 U12208 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n9748) );
  NAND3_X1 U12209 ( .A1(n14102), .A2(P1_IR_REG_0__SCAN_IN), .A3(n9748), .ZN(
        n9753) );
  NAND2_X1 U12210 ( .A1(n9745), .A2(n9795), .ZN(n9746) );
  NAND2_X1 U12211 ( .A1(n9747), .A2(n9746), .ZN(n14064) );
  AND2_X1 U12212 ( .A1(n14059), .A2(n9748), .ZN(n9749) );
  NOR2_X1 U12213 ( .A1(n14064), .A2(n9749), .ZN(n9750) );
  MUX2_X1 U12214 ( .A(n9750), .B(n14064), .S(P1_IR_REG_0__SCAN_IN), .Z(n9751)
         );
  AOI22_X1 U12215 ( .A1(n9794), .A2(n9751), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        P1_U3086), .ZN(n9752) );
  OAI211_X1 U12216 ( .C1(n14815), .C2(n9754), .A(n9753), .B(n9752), .ZN(
        P1_U3243) );
  INV_X1 U12217 ( .A(n9755), .ZN(n9759) );
  MUX2_X1 U12218 ( .A(n9690), .B(P2_REG2_REG_3__SCAN_IN), .S(n9760), .Z(n9758)
         );
  INV_X1 U12219 ( .A(n9756), .ZN(n9757) );
  AOI211_X1 U12220 ( .C1(n9759), .C2(n9758), .A(n9757), .B(n10113), .ZN(n9769)
         );
  AND2_X1 U12221 ( .A1(P2_U3088), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n10056) );
  INV_X1 U12222 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n9767) );
  MUX2_X1 U12223 ( .A(n9674), .B(P2_REG1_REG_3__SCAN_IN), .S(n9760), .Z(n9763)
         );
  NAND3_X1 U12224 ( .A1(n9763), .A2(n9762), .A3(n9761), .ZN(n9764) );
  NAND2_X1 U12225 ( .A1(n9765), .A2(n9764), .ZN(n9766) );
  OAI22_X1 U12226 ( .A1(n14901), .A2(n9767), .B1(n13511), .B2(n9766), .ZN(
        n9768) );
  NOR3_X1 U12227 ( .A1(n9769), .A2(n10056), .A3(n9768), .ZN(n9770) );
  OAI21_X1 U12228 ( .B1(n9771), .B2(n14894), .A(n9770), .ZN(P2_U3217) );
  XNOR2_X1 U12229 ( .A(n9873), .B(P1_DATAO_REG_13__SCAN_IN), .ZN(n11701) );
  OAI222_X1 U12230 ( .A1(n12764), .A2(P3_U3151), .B1(n13333), .B2(n11701), 
        .C1(n11702), .C2(n13335), .ZN(P3_U3282) );
  INV_X1 U12231 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n12318) );
  NAND2_X1 U12232 ( .A1(n6492), .A2(n9774), .ZN(n9775) );
  OAI21_X1 U12233 ( .B1(n6492), .B2(n12318), .A(n9775), .ZN(P2_U3562) );
  INV_X1 U12234 ( .A(n10102), .ZN(n9912) );
  INV_X1 U12235 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n9776) );
  OAI222_X1 U12236 ( .A1(P2_U3088), .A2(n9912), .B1(n13873), .B2(n9777), .C1(
        n9776), .C2(n13870), .ZN(P2_U3317) );
  INV_X1 U12237 ( .A(n10120), .ZN(n10115) );
  OAI222_X1 U12238 ( .A1(n14478), .A2(n9778), .B1(n14480), .B2(n9777), .C1(
        n10115), .C2(P1_U3086), .ZN(P1_U3345) );
  NAND2_X1 U12239 ( .A1(n13361), .A2(n6492), .ZN(n9779) );
  OAI21_X1 U12240 ( .B1(n7985), .B2(n6492), .A(n9779), .ZN(P2_U3551) );
  INV_X1 U12241 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n14995) );
  AOI22_X1 U12242 ( .A1(n14956), .A2(P2_REG1_REG_0__SCAN_IN), .B1(n14961), 
        .B2(P2_REG2_REG_0__SCAN_IN), .ZN(n9783) );
  INV_X1 U12243 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n15004) );
  NAND2_X1 U12244 ( .A1(n14961), .A2(n15004), .ZN(n9780) );
  OAI211_X1 U12245 ( .C1(P2_REG1_REG_0__SCAN_IN), .C2(n13511), .A(n14894), .B(
        n9780), .ZN(n9781) );
  INV_X1 U12246 ( .A(n9781), .ZN(n9782) );
  MUX2_X1 U12247 ( .A(n9783), .B(n9782), .S(P2_IR_REG_0__SCAN_IN), .Z(n9785)
         );
  NAND2_X1 U12248 ( .A1(n14954), .A2(P2_ADDR_REG_0__SCAN_IN), .ZN(n9784) );
  OAI211_X1 U12249 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n14995), .A(n9785), .B(
        n9784), .ZN(P2_U3214) );
  INV_X1 U12250 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n9786) );
  MUX2_X1 U12251 ( .A(n9786), .B(P1_REG1_REG_5__SCAN_IN), .S(n9884), .Z(n9792)
         );
  INV_X1 U12252 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n9787) );
  MUX2_X1 U12253 ( .A(n9787), .B(P1_REG1_REG_1__SCAN_IN), .S(n14052), .Z(
        n14050) );
  NAND2_X1 U12254 ( .A1(P1_REG1_REG_0__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n14049) );
  OR2_X1 U12255 ( .A1(n14050), .A2(n14049), .ZN(n14071) );
  NAND2_X1 U12256 ( .A1(n14052), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n14069) );
  INV_X1 U12257 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n14850) );
  MUX2_X1 U12258 ( .A(n14850), .B(P1_REG1_REG_2__SCAN_IN), .S(n14073), .Z(
        n14070) );
  AOI21_X1 U12259 ( .B1(n14071), .B2(n14069), .A(n14070), .ZN(n14068) );
  NOR2_X1 U12260 ( .A1(n9788), .A2(n14850), .ZN(n14089) );
  INV_X1 U12261 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n9789) );
  MUX2_X1 U12262 ( .A(n9789), .B(P1_REG1_REG_3__SCAN_IN), .S(n14090), .Z(n9790) );
  OAI21_X1 U12263 ( .B1(n14068), .B2(n14089), .A(n9790), .ZN(n14785) );
  NAND2_X1 U12264 ( .A1(n6752), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n14784) );
  INV_X1 U12265 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n14852) );
  MUX2_X1 U12266 ( .A(n14852), .B(P1_REG1_REG_4__SCAN_IN), .S(n9799), .Z(
        n14783) );
  AOI21_X1 U12267 ( .B1(n14785), .B2(n14784), .A(n14783), .ZN(n14787) );
  AOI21_X1 U12268 ( .B1(n9799), .B2(P1_REG1_REG_4__SCAN_IN), .A(n14787), .ZN(
        n9791) );
  NAND2_X1 U12269 ( .A1(n9791), .A2(n9792), .ZN(n9879) );
  OAI21_X1 U12270 ( .B1(n9792), .B2(n9791), .A(n9879), .ZN(n9804) );
  NOR2_X1 U12271 ( .A1(n8291), .A2(n14059), .ZN(n9793) );
  NAND2_X1 U12272 ( .A1(n9794), .A2(n9793), .ZN(n14807) );
  MUX2_X1 U12273 ( .A(n14341), .B(P1_REG2_REG_1__SCAN_IN), .S(n14052), .Z(
        n9796) );
  INV_X1 U12274 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n14065) );
  NOR3_X1 U12275 ( .A1(n9796), .A2(n14065), .A3(n9795), .ZN(n14078) );
  NOR2_X1 U12276 ( .A1(n7526), .A2(n14341), .ZN(n14074) );
  MUX2_X1 U12277 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n9797), .S(n14073), .Z(n9798) );
  OAI21_X1 U12278 ( .B1(n14078), .B2(n14074), .A(n9798), .ZN(n14085) );
  NAND2_X1 U12279 ( .A1(n14073), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n14084) );
  MUX2_X1 U12280 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n10600), .S(n14090), .Z(
        n14083) );
  AOI21_X1 U12281 ( .B1(n14085), .B2(n14084), .A(n14083), .ZN(n14791) );
  NOR2_X1 U12282 ( .A1(n14090), .A2(n10600), .ZN(n14790) );
  MUX2_X1 U12283 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n10830), .S(n9799), .Z(
        n14789) );
  OAI21_X1 U12284 ( .B1(n14791), .B2(n14790), .A(n14789), .ZN(n14788) );
  NAND2_X1 U12285 ( .A1(n9799), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n9801) );
  MUX2_X1 U12286 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n9883), .S(n9884), .Z(n9800)
         );
  AOI21_X1 U12287 ( .B1(n14788), .B2(n9801), .A(n9800), .ZN(n9888) );
  AND3_X1 U12288 ( .A1(n14788), .A2(n9801), .A3(n9800), .ZN(n9802) );
  NOR3_X1 U12289 ( .A1(n14807), .A2(n9888), .A3(n9802), .ZN(n9803) );
  AOI21_X1 U12290 ( .B1(n14102), .B2(n9804), .A(n9803), .ZN(n9807) );
  NAND2_X1 U12291 ( .A1(P1_U3086), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n10898) );
  INV_X1 U12292 ( .A(n10898), .ZN(n9805) );
  AOI21_X1 U12293 ( .B1(n14088), .B2(P1_ADDR_REG_5__SCAN_IN), .A(n9805), .ZN(
        n9806) );
  OAI211_X1 U12294 ( .C1(n9884), .C2(n14811), .A(n9807), .B(n9806), .ZN(
        P1_U3248) );
  XNOR2_X1 U12295 ( .A(n9808), .B(P3_B_REG_SCAN_IN), .ZN(n9809) );
  NOR2_X1 U12296 ( .A1(n10203), .A2(n10231), .ZN(n9812) );
  INV_X1 U12297 ( .A(P3_D_REG_2__SCAN_IN), .ZN(n9810) );
  NOR2_X1 U12298 ( .A1(n9829), .A2(n9810), .ZN(P3_U3263) );
  INV_X1 U12299 ( .A(P3_D_REG_4__SCAN_IN), .ZN(n9811) );
  NOR2_X1 U12300 ( .A1(n9829), .A2(n9811), .ZN(P3_U3261) );
  INV_X1 U12301 ( .A(P3_D_REG_7__SCAN_IN), .ZN(n9813) );
  NOR2_X1 U12302 ( .A1(n9829), .A2(n9813), .ZN(P3_U3258) );
  INV_X1 U12303 ( .A(P3_D_REG_8__SCAN_IN), .ZN(n9814) );
  NOR2_X1 U12304 ( .A1(n9829), .A2(n9814), .ZN(P3_U3257) );
  INV_X1 U12305 ( .A(P3_D_REG_9__SCAN_IN), .ZN(n9815) );
  NOR2_X1 U12306 ( .A1(n9829), .A2(n9815), .ZN(P3_U3256) );
  INV_X1 U12307 ( .A(P3_D_REG_6__SCAN_IN), .ZN(n9816) );
  NOR2_X1 U12308 ( .A1(n9829), .A2(n9816), .ZN(P3_U3259) );
  INV_X1 U12309 ( .A(P3_D_REG_11__SCAN_IN), .ZN(n13240) );
  NOR2_X1 U12310 ( .A1(n9829), .A2(n13240), .ZN(P3_U3254) );
  INV_X1 U12311 ( .A(P3_D_REG_12__SCAN_IN), .ZN(n9817) );
  NOR2_X1 U12312 ( .A1(n9829), .A2(n9817), .ZN(P3_U3253) );
  INV_X1 U12313 ( .A(P3_D_REG_13__SCAN_IN), .ZN(n9818) );
  NOR2_X1 U12314 ( .A1(n9829), .A2(n9818), .ZN(P3_U3252) );
  INV_X1 U12315 ( .A(P3_D_REG_5__SCAN_IN), .ZN(n9819) );
  NOR2_X1 U12316 ( .A1(n9812), .A2(n9819), .ZN(P3_U3260) );
  INV_X1 U12317 ( .A(P3_D_REG_15__SCAN_IN), .ZN(n9820) );
  NOR2_X1 U12318 ( .A1(n9829), .A2(n9820), .ZN(P3_U3250) );
  INV_X1 U12319 ( .A(P3_D_REG_16__SCAN_IN), .ZN(n9821) );
  NOR2_X1 U12320 ( .A1(n9829), .A2(n9821), .ZN(P3_U3249) );
  INV_X1 U12321 ( .A(P3_D_REG_17__SCAN_IN), .ZN(n9822) );
  NOR2_X1 U12322 ( .A1(n9829), .A2(n9822), .ZN(P3_U3248) );
  INV_X1 U12323 ( .A(P3_D_REG_18__SCAN_IN), .ZN(n9823) );
  NOR2_X1 U12324 ( .A1(n9829), .A2(n9823), .ZN(P3_U3247) );
  INV_X1 U12325 ( .A(P3_D_REG_10__SCAN_IN), .ZN(n9824) );
  NOR2_X1 U12326 ( .A1(n9829), .A2(n9824), .ZN(P3_U3255) );
  INV_X1 U12327 ( .A(P3_D_REG_19__SCAN_IN), .ZN(n9825) );
  NOR2_X1 U12328 ( .A1(n9829), .A2(n9825), .ZN(P3_U3246) );
  INV_X1 U12329 ( .A(P3_D_REG_3__SCAN_IN), .ZN(n9826) );
  NOR2_X1 U12330 ( .A1(n9812), .A2(n9826), .ZN(P3_U3262) );
  INV_X1 U12331 ( .A(P3_D_REG_20__SCAN_IN), .ZN(n9827) );
  NOR2_X1 U12332 ( .A1(n9812), .A2(n9827), .ZN(P3_U3245) );
  INV_X1 U12333 ( .A(P3_D_REG_14__SCAN_IN), .ZN(n9828) );
  NOR2_X1 U12334 ( .A1(n9829), .A2(n9828), .ZN(P3_U3251) );
  INV_X1 U12335 ( .A(P3_D_REG_22__SCAN_IN), .ZN(n9830) );
  NOR2_X1 U12336 ( .A1(n9812), .A2(n9830), .ZN(P3_U3243) );
  INV_X1 U12337 ( .A(P3_D_REG_23__SCAN_IN), .ZN(n9831) );
  NOR2_X1 U12338 ( .A1(n9812), .A2(n9831), .ZN(P3_U3242) );
  INV_X1 U12339 ( .A(P3_D_REG_24__SCAN_IN), .ZN(n9832) );
  NOR2_X1 U12340 ( .A1(n9812), .A2(n9832), .ZN(P3_U3241) );
  INV_X1 U12341 ( .A(P3_D_REG_25__SCAN_IN), .ZN(n9833) );
  NOR2_X1 U12342 ( .A1(n9812), .A2(n9833), .ZN(P3_U3240) );
  INV_X1 U12343 ( .A(P3_D_REG_26__SCAN_IN), .ZN(n13180) );
  NOR2_X1 U12344 ( .A1(n9812), .A2(n13180), .ZN(P3_U3239) );
  INV_X1 U12345 ( .A(P3_D_REG_21__SCAN_IN), .ZN(n9834) );
  NOR2_X1 U12346 ( .A1(n9812), .A2(n9834), .ZN(P3_U3244) );
  INV_X1 U12347 ( .A(P3_D_REG_27__SCAN_IN), .ZN(n9835) );
  NOR2_X1 U12348 ( .A1(n9812), .A2(n9835), .ZN(P3_U3238) );
  INV_X1 U12349 ( .A(P3_D_REG_28__SCAN_IN), .ZN(n9836) );
  NOR2_X1 U12350 ( .A1(n9812), .A2(n9836), .ZN(P3_U3237) );
  INV_X1 U12351 ( .A(P3_D_REG_29__SCAN_IN), .ZN(n9837) );
  NOR2_X1 U12352 ( .A1(n9829), .A2(n9837), .ZN(P3_U3236) );
  INV_X1 U12353 ( .A(P3_D_REG_30__SCAN_IN), .ZN(n9838) );
  NOR2_X1 U12354 ( .A1(n9829), .A2(n9838), .ZN(P3_U3235) );
  INV_X1 U12355 ( .A(P3_D_REG_31__SCAN_IN), .ZN(n9839) );
  NOR2_X1 U12356 ( .A1(n9829), .A2(n9839), .ZN(P3_U3234) );
  NOR2_X1 U12357 ( .A1(n13511), .A2(n9864), .ZN(n9856) );
  NAND2_X1 U12358 ( .A1(n9847), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n13453) );
  NAND2_X1 U12359 ( .A1(n13454), .A2(n13453), .ZN(n9842) );
  INV_X1 U12360 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n9840) );
  MUX2_X1 U12361 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n9840), .S(n13456), .Z(n9841) );
  NAND2_X1 U12362 ( .A1(n9842), .A2(n9841), .ZN(n13469) );
  NAND2_X1 U12363 ( .A1(n13456), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n13468) );
  NAND2_X1 U12364 ( .A1(n13469), .A2(n13468), .ZN(n9845) );
  INV_X1 U12365 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n9843) );
  MUX2_X1 U12366 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n9843), .S(n13472), .Z(n9844) );
  NAND2_X1 U12367 ( .A1(n9845), .A2(n9844), .ZN(n13471) );
  NAND2_X1 U12368 ( .A1(n13472), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n9846) );
  NAND2_X1 U12369 ( .A1(n13471), .A2(n9846), .ZN(n9866) );
  INV_X1 U12370 ( .A(n14894), .ZN(n14959) );
  NAND2_X1 U12371 ( .A1(n9847), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n13458) );
  NAND2_X1 U12372 ( .A1(n13459), .A2(n13458), .ZN(n9849) );
  INV_X1 U12373 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n10686) );
  MUX2_X1 U12374 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n10686), .S(n13456), .Z(
        n9848) );
  NAND2_X1 U12375 ( .A1(n9849), .A2(n9848), .ZN(n13475) );
  NAND2_X1 U12376 ( .A1(n13456), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n13474) );
  NAND2_X1 U12377 ( .A1(n13475), .A2(n13474), .ZN(n9851) );
  INV_X1 U12378 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n10719) );
  MUX2_X1 U12379 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n10719), .S(n13472), .Z(
        n9850) );
  NAND2_X1 U12380 ( .A1(n9851), .A2(n9850), .ZN(n13477) );
  NAND2_X1 U12381 ( .A1(n13472), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n9852) );
  NAND2_X1 U12382 ( .A1(n13477), .A2(n9852), .ZN(n9859) );
  INV_X1 U12383 ( .A(n9859), .ZN(n9854) );
  INV_X1 U12384 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n9853) );
  NOR3_X1 U12385 ( .A1(n9854), .A2(n10113), .A3(n9853), .ZN(n9855) );
  AOI211_X1 U12386 ( .C1(n9856), .C2(n9866), .A(n14959), .B(n9855), .ZN(n9872)
         );
  NAND2_X1 U12387 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3088), .ZN(n10914) );
  INV_X1 U12388 ( .A(n10914), .ZN(n9862) );
  MUX2_X1 U12389 ( .A(n9853), .B(P2_REG2_REG_9__SCAN_IN), .S(n9902), .Z(n9857)
         );
  OR2_X1 U12390 ( .A1(n9859), .A2(n9857), .ZN(n9897) );
  OR2_X1 U12391 ( .A1(n9902), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n9896) );
  INV_X1 U12392 ( .A(n9896), .ZN(n9858) );
  NAND2_X1 U12393 ( .A1(n9859), .A2(n9858), .ZN(n9860) );
  AOI21_X1 U12394 ( .B1(n9897), .B2(n9860), .A(n10113), .ZN(n9861) );
  AOI211_X1 U12395 ( .C1(n14954), .C2(P2_ADDR_REG_9__SCAN_IN), .A(n9862), .B(
        n9861), .ZN(n9870) );
  INV_X1 U12396 ( .A(n9866), .ZN(n9863) );
  NOR3_X1 U12397 ( .A1(n9863), .A2(n9902), .A3(P2_REG1_REG_9__SCAN_IN), .ZN(
        n9868) );
  INV_X1 U12398 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n9864) );
  MUX2_X1 U12399 ( .A(n9864), .B(P2_REG1_REG_9__SCAN_IN), .S(n9902), .Z(n9865)
         );
  OR2_X1 U12400 ( .A1(n9866), .A2(n9865), .ZN(n9904) );
  INV_X1 U12401 ( .A(n9904), .ZN(n9867) );
  OAI21_X1 U12402 ( .B1(n9868), .B2(n9867), .A(n14956), .ZN(n9869) );
  OAI211_X1 U12403 ( .C1(n9872), .C2(n9871), .A(n9870), .B(n9869), .ZN(
        P2_U3223) );
  NAND2_X1 U12404 ( .A1(n10283), .A2(n9874), .ZN(n9875) );
  NAND2_X1 U12405 ( .A1(n10524), .A2(P2_DATAO_REG_14__SCAN_IN), .ZN(n9937) );
  INV_X1 U12406 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n10523) );
  NAND2_X1 U12407 ( .A1(n10523), .A2(P1_DATAO_REG_14__SCAN_IN), .ZN(n9876) );
  NAND2_X1 U12408 ( .A1(n9937), .A2(n9876), .ZN(n9938) );
  XNOR2_X1 U12409 ( .A(n9939), .B(n9938), .ZN(n11940) );
  INV_X1 U12410 ( .A(n11940), .ZN(n9878) );
  OAI222_X1 U12411 ( .A1(n12783), .A2(P3_U3151), .B1(n13333), .B2(n9878), .C1(
        n9877), .C2(n13335), .ZN(P3_U3281) );
  OAI21_X1 U12412 ( .B1(n9880), .B2(P1_REG1_REG_5__SCAN_IN), .A(n9879), .ZN(
        n9882) );
  INV_X1 U12413 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n9942) );
  MUX2_X1 U12414 ( .A(n9942), .B(P1_REG1_REG_6__SCAN_IN), .S(n9885), .Z(n9881)
         );
  NOR2_X1 U12415 ( .A1(n9882), .A2(n9881), .ZN(n9948) );
  AOI211_X1 U12416 ( .C1(n9882), .C2(n9881), .A(n9948), .B(n14809), .ZN(n9892)
         );
  NOR2_X1 U12417 ( .A1(n9884), .A2(n9883), .ZN(n9887) );
  MUX2_X1 U12418 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n10942), .S(n9885), .Z(n9886) );
  OAI21_X1 U12419 ( .B1(n9888), .B2(n9887), .A(n9886), .ZN(n9949) );
  INV_X1 U12420 ( .A(n9949), .ZN(n9890) );
  NOR3_X1 U12421 ( .A1(n9888), .A2(n9887), .A3(n9886), .ZN(n9889) );
  NOR3_X1 U12422 ( .A1(n14807), .A2(n9890), .A3(n9889), .ZN(n9891) );
  NOR2_X1 U12423 ( .A1(n9892), .A2(n9891), .ZN(n9895) );
  INV_X1 U12424 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n9893) );
  NOR2_X1 U12425 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n9893), .ZN(n13997) );
  AOI21_X1 U12426 ( .B1(n14088), .B2(P1_ADDR_REG_6__SCAN_IN), .A(n13997), .ZN(
        n9894) );
  OAI211_X1 U12427 ( .C1(n9950), .C2(n14811), .A(n9895), .B(n9894), .ZN(
        P1_U3249) );
  NAND2_X1 U12428 ( .A1(n9897), .A2(n9896), .ZN(n9900) );
  INV_X1 U12429 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n9898) );
  MUX2_X1 U12430 ( .A(n9898), .B(P2_REG2_REG_10__SCAN_IN), .S(n10102), .Z(
        n9899) );
  AOI21_X1 U12431 ( .B1(n9900), .B2(n9899), .A(n10113), .ZN(n9901) );
  OR2_X1 U12432 ( .A1(n9900), .A2(n9899), .ZN(n10097) );
  NAND2_X1 U12433 ( .A1(n9901), .A2(n10097), .ZN(n9911) );
  NAND2_X1 U12434 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3088), .ZN(n11056)
         );
  INV_X1 U12435 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n10893) );
  MUX2_X1 U12436 ( .A(n10893), .B(P2_REG1_REG_10__SCAN_IN), .S(n10102), .Z(
        n9905) );
  OR2_X1 U12437 ( .A1(n9902), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n9903) );
  NAND2_X1 U12438 ( .A1(n9904), .A2(n9903), .ZN(n9906) );
  AOI21_X1 U12439 ( .B1(n9905), .B2(n9906), .A(n13511), .ZN(n9907) );
  OR2_X1 U12440 ( .A1(n9906), .A2(n9905), .ZN(n10108) );
  NAND2_X1 U12441 ( .A1(n9907), .A2(n10108), .ZN(n9908) );
  NAND2_X1 U12442 ( .A1(n11056), .A2(n9908), .ZN(n9909) );
  AOI21_X1 U12443 ( .B1(n14954), .B2(P2_ADDR_REG_10__SCAN_IN), .A(n9909), .ZN(
        n9910) );
  OAI211_X1 U12444 ( .C1(n14894), .C2(n9912), .A(n9911), .B(n9910), .ZN(
        P2_U3224) );
  INV_X1 U12445 ( .A(n10822), .ZN(n9914) );
  AOI22_X1 U12446 ( .A1(n9914), .A2(n14324), .B1(n14321), .B2(n14045), .ZN(
        n10818) );
  NAND3_X1 U12447 ( .A1(n9548), .A2(n11614), .A3(n9915), .ZN(n9916) );
  OAI211_X1 U12448 ( .C1(n14431), .C2(n10822), .A(n10818), .B(n9916), .ZN(
        n14433) );
  NAND2_X1 U12449 ( .A1(n14433), .A2(n14849), .ZN(n9917) );
  OAI21_X1 U12450 ( .B1(n14849), .B2(n7512), .A(n9917), .ZN(P1_U3459) );
  INV_X1 U12451 ( .A(P3_DATAO_REG_9__SCAN_IN), .ZN(n13276) );
  XNOR2_X2 U12452 ( .A(n9919), .B(P3_IR_REG_30__SCAN_IN), .ZN(n9922) );
  XNOR2_X2 U12453 ( .A(n9921), .B(P3_IR_REG_29__SCAN_IN), .ZN(n9926) );
  NAND2_X1 U12454 ( .A1(n12155), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n9930) );
  NAND2_X1 U12455 ( .A1(n10454), .A2(P3_REG0_REG_9__SCAN_IN), .ZN(n9929) );
  NOR2_X1 U12456 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_5__SCAN_IN), 
        .ZN(n9924) );
  INV_X1 U12457 ( .A(P3_REG3_REG_4__SCAN_IN), .ZN(n9923) );
  NAND2_X1 U12458 ( .A1(n9924), .A2(n9923), .ZN(n10929) );
  NOR2_X1 U12459 ( .A1(n11075), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n11093) );
  NAND2_X1 U12460 ( .A1(n11093), .A2(n11092), .ZN(n11095) );
  NAND2_X1 U12461 ( .A1(n11095), .A2(P3_REG3_REG_9__SCAN_IN), .ZN(n9925) );
  NAND2_X1 U12462 ( .A1(n11316), .A2(n9925), .ZN(n11505) );
  NAND2_X1 U12463 ( .A1(n10235), .A2(n11505), .ZN(n9928) );
  NAND2_X1 U12464 ( .A1(n6491), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n9927) );
  NAND4_X1 U12465 ( .A1(n9930), .A2(n9929), .A3(n9928), .A4(n9927), .ZN(n12411) );
  NAND2_X1 U12466 ( .A1(n12411), .A2(P3_U3897), .ZN(n9931) );
  OAI21_X1 U12467 ( .B1(P3_U3897), .B2(n13276), .A(n9931), .ZN(P3_U3500) );
  INV_X1 U12468 ( .A(n9932), .ZN(n9935) );
  INV_X1 U12469 ( .A(n14107), .ZN(n10116) );
  OAI222_X1 U12470 ( .A1(n14478), .A2(n9933), .B1(n14480), .B2(n9935), .C1(
        P1_U3086), .C2(n10116), .ZN(P1_U3344) );
  INV_X1 U12471 ( .A(n13494), .ZN(n9934) );
  OAI222_X1 U12472 ( .A1(n13870), .A2(n9936), .B1(n13873), .B2(n9935), .C1(
        P2_U3088), .C2(n9934), .ZN(P2_U3316) );
  XNOR2_X1 U12473 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .ZN(n9940) );
  XNOR2_X1 U12474 ( .A(n10150), .B(n9940), .ZN(n11976) );
  AOI222_X1 U12475 ( .A1(n11976), .A2(n13320), .B1(SI_15_), .B2(n12092), .C1(
        P3_STATE_REG_SCAN_IN), .C2(n14623), .ZN(n9941) );
  INV_X1 U12476 ( .A(n9941), .ZN(P3_U3280) );
  NOR2_X1 U12477 ( .A1(n9950), .A2(n9942), .ZN(n9946) );
  INV_X1 U12478 ( .A(n9946), .ZN(n9944) );
  INV_X1 U12479 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n10021) );
  MUX2_X1 U12480 ( .A(n10021), .B(P1_REG1_REG_7__SCAN_IN), .S(n10011), .Z(
        n9943) );
  NAND2_X1 U12481 ( .A1(n9944), .A2(n9943), .ZN(n9947) );
  MUX2_X1 U12482 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n10021), .S(n10011), .Z(
        n9945) );
  OAI21_X1 U12483 ( .B1(n9948), .B2(n9946), .A(n9945), .ZN(n10019) );
  OAI211_X1 U12484 ( .C1(n9948), .C2(n9947), .A(n10019), .B(n14102), .ZN(n9957) );
  NAND2_X1 U12485 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3086), .ZN(n11197) );
  OAI21_X1 U12486 ( .B1(n10942), .B2(n9950), .A(n9949), .ZN(n9953) );
  MUX2_X1 U12487 ( .A(n7658), .B(P1_REG2_REG_7__SCAN_IN), .S(n10011), .Z(n9951) );
  INV_X1 U12488 ( .A(n9951), .ZN(n9952) );
  NAND2_X1 U12489 ( .A1(n9953), .A2(n9952), .ZN(n10068) );
  OAI211_X1 U12490 ( .C1(n9953), .C2(n9952), .A(n14113), .B(n10068), .ZN(n9954) );
  NAND2_X1 U12491 ( .A1(n11197), .A2(n9954), .ZN(n9955) );
  AOI21_X1 U12492 ( .B1(n14088), .B2(P1_ADDR_REG_7__SCAN_IN), .A(n9955), .ZN(
        n9956) );
  OAI211_X1 U12493 ( .C1(n14811), .C2(n10020), .A(n9957), .B(n9956), .ZN(
        P1_U3250) );
  NOR4_X1 U12494 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_17__SCAN_IN), .A3(
        P2_D_REG_18__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n9961) );
  NOR4_X1 U12495 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_12__SCAN_IN), .A4(P2_D_REG_13__SCAN_IN), .ZN(n9960) );
  NOR4_X1 U12496 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n9959) );
  NOR4_X1 U12497 ( .A1(P2_D_REG_21__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .A3(
        P2_D_REG_23__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n9958) );
  NAND4_X1 U12498 ( .A1(n9961), .A2(n9960), .A3(n9959), .A4(n9958), .ZN(n9971)
         );
  NOR2_X1 U12499 ( .A1(P2_D_REG_19__SCAN_IN), .A2(P2_D_REG_16__SCAN_IN), .ZN(
        n9965) );
  NOR4_X1 U12500 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n9964) );
  NOR4_X1 U12501 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_8__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_10__SCAN_IN), .ZN(n9963) );
  NOR4_X1 U12502 ( .A1(P2_D_REG_3__SCAN_IN), .A2(P2_D_REG_4__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_6__SCAN_IN), .ZN(n9962) );
  NAND4_X1 U12503 ( .A1(n9965), .A2(n9964), .A3(n9963), .A4(n9962), .ZN(n9970)
         );
  INV_X1 U12504 ( .A(n9966), .ZN(n11880) );
  XNOR2_X1 U12505 ( .A(n11815), .B(P2_B_REG_SCAN_IN), .ZN(n9967) );
  NAND2_X1 U12506 ( .A1(n11880), .A2(n9967), .ZN(n9968) );
  NAND2_X1 U12507 ( .A1(n11815), .A2(n12011), .ZN(n9973) );
  INV_X1 U12508 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n15011) );
  NAND2_X1 U12509 ( .A1(n15006), .A2(n15011), .ZN(n9972) );
  NAND2_X1 U12510 ( .A1(n9973), .A2(n9972), .ZN(n15012) );
  INV_X1 U12511 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n15014) );
  NAND2_X1 U12512 ( .A1(n15006), .A2(n15014), .ZN(n9975) );
  NAND2_X1 U12513 ( .A1(n12011), .A2(n11880), .ZN(n9974) );
  NAND2_X1 U12514 ( .A1(n9975), .A2(n9974), .ZN(n15015) );
  NOR2_X1 U12515 ( .A1(n15012), .A2(n15015), .ZN(n9976) );
  NAND2_X1 U12516 ( .A1(n10677), .A2(n9976), .ZN(n9981) );
  NOR2_X1 U12517 ( .A1(n14989), .A2(n11523), .ZN(n10680) );
  NAND2_X1 U12518 ( .A1(n9989), .A2(n10680), .ZN(n9977) );
  INV_X1 U12519 ( .A(n9978), .ZN(n9986) );
  INV_X1 U12520 ( .A(n9998), .ZN(n10350) );
  INV_X1 U12521 ( .A(n9251), .ZN(n9979) );
  OR2_X1 U12522 ( .A1(n9987), .A2(n9979), .ZN(n13370) );
  OAI22_X1 U12523 ( .A1(n10350), .A2(n13591), .B1(n10357), .B2(n13370), .ZN(
        n10764) );
  INV_X1 U12524 ( .A(n10339), .ZN(n9980) );
  NAND2_X1 U12525 ( .A1(n9981), .A2(n9980), .ZN(n9985) );
  OR2_X1 U12526 ( .A1(n9987), .A2(n9986), .ZN(n10341) );
  AND3_X1 U12527 ( .A1(n9983), .A2(n9982), .A3(n10341), .ZN(n9984) );
  NAND2_X1 U12528 ( .A1(n9985), .A2(n9984), .ZN(n10053) );
  OR2_X1 U12529 ( .A1(n10053), .A2(P2_U3088), .ZN(n10074) );
  AOI22_X1 U12530 ( .A1(n13374), .A2(n10764), .B1(n10074), .B2(
        P2_REG3_REG_2__SCAN_IN), .ZN(n10010) );
  AND2_X1 U12531 ( .A1(n15077), .A2(n9987), .ZN(n9988) );
  NAND2_X1 U12532 ( .A1(n13448), .A2(n12605), .ZN(n9994) );
  NAND2_X1 U12533 ( .A1(n9993), .A2(n9994), .ZN(n10051) );
  INV_X1 U12534 ( .A(n9993), .ZN(n9996) );
  INV_X1 U12535 ( .A(n9994), .ZN(n9995) );
  NAND2_X1 U12536 ( .A1(n9996), .A2(n9995), .ZN(n9997) );
  INV_X1 U12537 ( .A(n10002), .ZN(n10000) );
  INV_X1 U12538 ( .A(n10001), .ZN(n9999) );
  NAND2_X1 U12539 ( .A1(n10000), .A2(n9999), .ZN(n10003) );
  MUX2_X1 U12540 ( .A(n12605), .B(n9992), .S(n6945), .Z(n10004) );
  NAND2_X1 U12541 ( .A1(n10004), .A2(n10075), .ZN(n10031) );
  NAND2_X1 U12542 ( .A1(n10030), .A2(n10005), .ZN(n10006) );
  NAND2_X1 U12543 ( .A1(n10006), .A2(n10007), .ZN(n10052) );
  OAI21_X1 U12544 ( .B1(n10007), .B2(n10006), .A(n10052), .ZN(n10008) );
  NAND2_X1 U12545 ( .A1(n13391), .A2(n10008), .ZN(n10009) );
  OAI211_X1 U12546 ( .C1(n6747), .C2(n13415), .A(n10010), .B(n10009), .ZN(
        P2_U3209) );
  NAND2_X1 U12547 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_U3086), .ZN(n11760) );
  OAI21_X1 U12548 ( .B1(n14815), .B2(n14485), .A(n11760), .ZN(n10018) );
  NAND2_X1 U12549 ( .A1(n10011), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n10067) );
  MUX2_X1 U12550 ( .A(n7686), .B(P1_REG2_REG_8__SCAN_IN), .S(n10023), .Z(
        n10066) );
  AOI21_X1 U12551 ( .B1(n10068), .B2(n10067), .A(n10066), .ZN(n10065) );
  NOR2_X1 U12552 ( .A1(n10063), .A2(n7686), .ZN(n10014) );
  MUX2_X1 U12553 ( .A(P1_REG2_REG_9__SCAN_IN), .B(n10012), .S(n10042), .Z(
        n10013) );
  OAI21_X1 U12554 ( .B1(n10065), .B2(n10014), .A(n10013), .ZN(n10045) );
  INV_X1 U12555 ( .A(n10045), .ZN(n10016) );
  NOR3_X1 U12556 ( .A1(n10065), .A2(n10014), .A3(n10013), .ZN(n10015) );
  NOR3_X1 U12557 ( .A1(n10016), .A2(n10015), .A3(n14807), .ZN(n10017) );
  AOI211_X1 U12558 ( .C1(n14108), .C2(n10042), .A(n10018), .B(n10017), .ZN(
        n10029) );
  OAI21_X1 U12559 ( .B1(n10021), .B2(n10020), .A(n10019), .ZN(n10061) );
  INV_X1 U12560 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n10022) );
  MUX2_X1 U12561 ( .A(n10022), .B(P1_REG1_REG_8__SCAN_IN), .S(n10023), .Z(
        n10062) );
  NOR2_X1 U12562 ( .A1(n10061), .A2(n10062), .ZN(n10060) );
  NOR2_X1 U12563 ( .A1(n10023), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n10024) );
  MUX2_X1 U12564 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n7709), .S(n10042), .Z(
        n10025) );
  OAI21_X1 U12565 ( .B1(n10060), .B2(n10024), .A(n10025), .ZN(n10038) );
  INV_X1 U12566 ( .A(n10038), .ZN(n10027) );
  NOR3_X1 U12567 ( .A1(n10060), .A2(n10025), .A3(n10024), .ZN(n10026) );
  OAI21_X1 U12568 ( .B1(n10027), .B2(n10026), .A(n14102), .ZN(n10028) );
  NAND2_X1 U12569 ( .A1(n10029), .A2(n10028), .ZN(P1_U3252) );
  OAI21_X1 U12570 ( .B1(n10032), .B2(n10031), .A(n10030), .ZN(n10033) );
  AOI22_X1 U12571 ( .A1(n13426), .A2(n10987), .B1(n13391), .B2(n10033), .ZN(
        n10037) );
  INV_X2 U12572 ( .A(n13370), .ZN(n13524) );
  NAND2_X1 U12573 ( .A1(n13524), .A2(n13448), .ZN(n10035) );
  NAND2_X1 U12574 ( .A1(n13420), .A2(n9205), .ZN(n10034) );
  NAND2_X1 U12575 ( .A1(n10035), .A2(n10034), .ZN(n10979) );
  AOI22_X1 U12576 ( .A1(n13374), .A2(n10979), .B1(n10074), .B2(
        P2_REG3_REG_1__SCAN_IN), .ZN(n10036) );
  NAND2_X1 U12577 ( .A1(n10037), .A2(n10036), .ZN(P2_U3194) );
  OAI21_X1 U12578 ( .B1(n10042), .B2(P1_REG1_REG_9__SCAN_IN), .A(n10038), .ZN(
        n10041) );
  INV_X1 U12579 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n10039) );
  MUX2_X1 U12580 ( .A(n10039), .B(P1_REG1_REG_10__SCAN_IN), .S(n10120), .Z(
        n10040) );
  NOR2_X1 U12581 ( .A1(n10041), .A2(n10040), .ZN(n10119) );
  AOI211_X1 U12582 ( .C1(n10041), .C2(n10040), .A(n14809), .B(n10119), .ZN(
        n10050) );
  NAND2_X1 U12583 ( .A1(n10042), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n10044) );
  MUX2_X1 U12584 ( .A(n11357), .B(P1_REG2_REG_10__SCAN_IN), .S(n10120), .Z(
        n10043) );
  AOI21_X1 U12585 ( .B1(n10045), .B2(n10044), .A(n10043), .ZN(n14111) );
  AND3_X1 U12586 ( .A1(n10045), .A2(n10044), .A3(n10043), .ZN(n10046) );
  NOR3_X1 U12587 ( .A1(n14111), .A2(n10046), .A3(n14807), .ZN(n10049) );
  NAND2_X1 U12588 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n11660)
         );
  NAND2_X1 U12589 ( .A1(n14088), .A2(P1_ADDR_REG_10__SCAN_IN), .ZN(n10047) );
  OAI211_X1 U12590 ( .C1(n14811), .C2(n10115), .A(n11660), .B(n10047), .ZN(
        n10048) );
  OR3_X1 U12591 ( .A1(n10050), .A2(n10049), .A3(n10048), .ZN(P1_U3253) );
  XNOR2_X1 U12592 ( .A(n10375), .B(n10389), .ZN(n10081) );
  NAND2_X1 U12593 ( .A1(n13447), .A2(n12605), .ZN(n10082) );
  XOR2_X1 U12594 ( .A(n10081), .B(n10082), .Z(n10084) );
  XNOR2_X1 U12595 ( .A(n10085), .B(n10084), .ZN(n10059) );
  NAND2_X1 U12596 ( .A1(n10053), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13372) );
  AOI22_X1 U12597 ( .A1(n13426), .A2(n10375), .B1(n8686), .B2(n13422), .ZN(
        n10058) );
  NAND2_X1 U12598 ( .A1(n13524), .A2(n13446), .ZN(n10055) );
  NAND2_X1 U12599 ( .A1(n13420), .A2(n13448), .ZN(n10054) );
  NAND2_X1 U12600 ( .A1(n10055), .A2(n10054), .ZN(n15039) );
  AOI21_X1 U12601 ( .B1(n13374), .B2(n15039), .A(n10056), .ZN(n10057) );
  OAI211_X1 U12602 ( .C1(n10059), .C2(n13428), .A(n10058), .B(n10057), .ZN(
        P2_U3190) );
  AOI21_X1 U12603 ( .B1(n10062), .B2(n10061), .A(n10060), .ZN(n10073) );
  AND2_X1 U12604 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n11467) );
  NOR2_X1 U12605 ( .A1(n14811), .A2(n10063), .ZN(n10064) );
  AOI211_X1 U12606 ( .C1(n14088), .C2(P1_ADDR_REG_8__SCAN_IN), .A(n11467), .B(
        n10064), .ZN(n10072) );
  INV_X1 U12607 ( .A(n10065), .ZN(n10070) );
  NAND3_X1 U12608 ( .A1(n10068), .A2(n10067), .A3(n10066), .ZN(n10069) );
  NAND3_X1 U12609 ( .A1(n10070), .A2(n14113), .A3(n10069), .ZN(n10071) );
  OAI211_X1 U12610 ( .C1(n10073), .C2(n14809), .A(n10072), .B(n10071), .ZN(
        P1_U3251) );
  NAND2_X1 U12611 ( .A1(n13524), .A2(n9998), .ZN(n14999) );
  AOI22_X1 U12612 ( .A1(n13426), .A2(n14990), .B1(P2_REG3_REG_0__SCAN_IN), 
        .B2(n10074), .ZN(n10080) );
  INV_X1 U12613 ( .A(n10075), .ZN(n10978) );
  NOR2_X1 U12614 ( .A1(n10076), .A2(n10086), .ZN(n10077) );
  MUX2_X1 U12615 ( .A(n10077), .B(n10086), .S(n14990), .Z(n10078) );
  OAI21_X1 U12616 ( .B1(n10978), .B2(n10078), .A(n13391), .ZN(n10079) );
  OAI211_X1 U12617 ( .C1(n14999), .C2(n13424), .A(n10080), .B(n10079), .ZN(
        P2_U3204) );
  INV_X1 U12618 ( .A(n10081), .ZN(n10083) );
  XNOR2_X1 U12619 ( .A(n15049), .B(n9992), .ZN(n10088) );
  NAND2_X1 U12620 ( .A1(n13446), .A2(n12610), .ZN(n10087) );
  NAND2_X1 U12621 ( .A1(n10088), .A2(n10087), .ZN(n10267) );
  OAI21_X1 U12622 ( .B1(n10088), .B2(n10087), .A(n10267), .ZN(n10089) );
  NOR2_X1 U12623 ( .A1(n10090), .A2(n10089), .ZN(n10269) );
  AOI21_X1 U12624 ( .B1(n10090), .B2(n10089), .A(n10269), .ZN(n10095) );
  NAND2_X1 U12625 ( .A1(n13524), .A2(n13445), .ZN(n10092) );
  NAND2_X1 U12626 ( .A1(n13420), .A2(n13447), .ZN(n10091) );
  NAND2_X1 U12627 ( .A1(n10092), .A2(n10091), .ZN(n14973) );
  AOI22_X1 U12628 ( .A1(n13374), .A2(n14973), .B1(P2_REG3_REG_4__SCAN_IN), 
        .B2(P2_U3088), .ZN(n10094) );
  AOI22_X1 U12629 ( .A1(n13426), .A2(n15049), .B1(n13422), .B2(n14978), .ZN(
        n10093) );
  OAI211_X1 U12630 ( .C1(n10095), .C2(n13428), .A(n10094), .B(n10093), .ZN(
        P2_U3202) );
  NAND2_X1 U12631 ( .A1(n10102), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n10096) );
  NAND2_X1 U12632 ( .A1(n10097), .A2(n10096), .ZN(n10101) );
  INV_X1 U12633 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n10098) );
  MUX2_X1 U12634 ( .A(n10098), .B(P2_REG2_REG_11__SCAN_IN), .S(n13494), .Z(
        n10100) );
  INV_X1 U12635 ( .A(n14888), .ZN(n10099) );
  AOI21_X1 U12636 ( .B1(n10101), .B2(n10100), .A(n10099), .ZN(n10114) );
  INV_X1 U12637 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n14766) );
  NAND2_X1 U12638 ( .A1(P2_REG3_REG_11__SCAN_IN), .A2(P2_U3088), .ZN(n11282)
         );
  OAI21_X1 U12639 ( .B1(n14901), .B2(n14766), .A(n11282), .ZN(n10111) );
  NAND2_X1 U12640 ( .A1(n10102), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n10107) );
  NAND2_X1 U12641 ( .A1(n10108), .A2(n10107), .ZN(n10105) );
  INV_X1 U12642 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n10103) );
  MUX2_X1 U12643 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n10103), .S(n13494), .Z(
        n10104) );
  NAND2_X1 U12644 ( .A1(n10105), .A2(n10104), .ZN(n13496) );
  MUX2_X1 U12645 ( .A(n10103), .B(P2_REG1_REG_11__SCAN_IN), .S(n13494), .Z(
        n10106) );
  NAND3_X1 U12646 ( .A1(n10108), .A2(n10107), .A3(n10106), .ZN(n10109) );
  AND3_X1 U12647 ( .A1(n13496), .A2(n14956), .A3(n10109), .ZN(n10110) );
  AOI211_X1 U12648 ( .C1(n14959), .C2(n13494), .A(n10111), .B(n10110), .ZN(
        n10112) );
  OAI21_X1 U12649 ( .B1(n10114), .B2(n10113), .A(n10112), .ZN(P2_U3225) );
  MUX2_X1 U12650 ( .A(n11484), .B(P1_REG2_REG_12__SCAN_IN), .S(n10126), .Z(
        n10118) );
  NOR2_X1 U12651 ( .A1(n10115), .A2(n11357), .ZN(n14110) );
  MUX2_X1 U12652 ( .A(P1_REG2_REG_11__SCAN_IN), .B(n11419), .S(n14107), .Z(
        n14109) );
  OAI21_X1 U12653 ( .B1(n14111), .B2(n14110), .A(n14109), .ZN(n14114) );
  OAI21_X1 U12654 ( .B1(n10116), .B2(n11419), .A(n14114), .ZN(n10117) );
  NOR2_X1 U12655 ( .A1(n10117), .A2(n10118), .ZN(n10258) );
  AOI21_X1 U12656 ( .B1(n10118), .B2(n10117), .A(n10258), .ZN(n10131) );
  AOI21_X1 U12657 ( .B1(n10120), .B2(P1_REG1_REG_10__SCAN_IN), .A(n10119), 
        .ZN(n14101) );
  NOR2_X1 U12658 ( .A1(n14107), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n10121) );
  AOI21_X1 U12659 ( .B1(n14107), .B2(P1_REG1_REG_11__SCAN_IN), .A(n10121), 
        .ZN(n14100) );
  NAND2_X1 U12660 ( .A1(n14101), .A2(n14100), .ZN(n14099) );
  INV_X1 U12661 ( .A(n10121), .ZN(n10124) );
  OR2_X1 U12662 ( .A1(n10126), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n10255) );
  NAND2_X1 U12663 ( .A1(n10126), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n10122) );
  NAND2_X1 U12664 ( .A1(n10255), .A2(n10122), .ZN(n10123) );
  AOI21_X1 U12665 ( .B1(n14099), .B2(n10124), .A(n10123), .ZN(n10257) );
  AND3_X1 U12666 ( .A1(n14099), .A2(n10124), .A3(n10123), .ZN(n10125) );
  OAI21_X1 U12667 ( .B1(n10257), .B2(n10125), .A(n14102), .ZN(n10130) );
  NOR2_X1 U12668 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n11897), .ZN(n10128) );
  INV_X1 U12669 ( .A(n10126), .ZN(n10259) );
  NOR2_X1 U12670 ( .A1(n14811), .A2(n10259), .ZN(n10127) );
  AOI211_X1 U12671 ( .C1(n14088), .C2(P1_ADDR_REG_12__SCAN_IN), .A(n10128), 
        .B(n10127), .ZN(n10129) );
  OAI211_X1 U12672 ( .C1(n10131), .C2(n14807), .A(n10130), .B(n10129), .ZN(
        P1_U3255) );
  OAI21_X1 U12673 ( .B1(n10134), .B2(n10133), .A(n10132), .ZN(n14060) );
  AOI22_X1 U12674 ( .A1(n14060), .A2(n13995), .B1(n9548), .B2(n14018), .ZN(
        n10137) );
  INV_X1 U12675 ( .A(n14013), .ZN(n13987) );
  NAND2_X1 U12676 ( .A1(n10135), .A2(n10593), .ZN(n10145) );
  AOI22_X1 U12677 ( .A1(n13987), .A2(n14045), .B1(P1_REG3_REG_0__SCAN_IN), 
        .B2(n10145), .ZN(n10136) );
  NAND2_X1 U12678 ( .A1(n10137), .A2(n10136), .ZN(P1_U3232) );
  XOR2_X1 U12679 ( .A(n10139), .B(n10138), .Z(n10142) );
  AOI22_X1 U12680 ( .A1(n10623), .A2(n14018), .B1(n10145), .B2(
        P1_REG3_REG_2__SCAN_IN), .ZN(n10141) );
  AOI22_X1 U12681 ( .A1(n13987), .A2(n14042), .B1(n14011), .B2(n14045), .ZN(
        n10140) );
  OAI211_X1 U12682 ( .C1(n10142), .C2(n14022), .A(n10141), .B(n10140), .ZN(
        P1_U3237) );
  XOR2_X1 U12683 ( .A(n10144), .B(n10143), .Z(n10148) );
  AOI22_X1 U12684 ( .A1(n14345), .A2(n14018), .B1(n10145), .B2(
        P1_REG3_REG_1__SCAN_IN), .ZN(n10147) );
  AOI22_X1 U12685 ( .A1(n13987), .A2(n14043), .B1(n14011), .B2(n14046), .ZN(
        n10146) );
  OAI211_X1 U12686 ( .C1(n10148), .C2(n14022), .A(n10147), .B(n10146), .ZN(
        P1_U3222) );
  NAND2_X1 U12687 ( .A1(n10781), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n10151) );
  AOI22_X1 U12688 ( .A1(P2_DATAO_REG_16__SCAN_IN), .A2(
        P1_DATAO_REG_16__SCAN_IN), .B1(n7884), .B2(n10976), .ZN(n10323) );
  XNOR2_X1 U12689 ( .A(n10324), .B(n7154), .ZN(n12130) );
  INV_X1 U12690 ( .A(n12130), .ZN(n10154) );
  OAI222_X1 U12691 ( .A1(n13333), .A2(n10154), .B1(n10153), .B2(P3_U3151), 
        .C1(n10152), .C2(n13335), .ZN(P3_U3279) );
  OAI21_X1 U12692 ( .B1(n15103), .B2(n10155), .A(n10423), .ZN(n10165) );
  INV_X1 U12693 ( .A(P3_ADDR_REG_1__SCAN_IN), .ZN(n10156) );
  INV_X1 U12694 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n10307) );
  OAI22_X1 U12695 ( .A1(n15168), .A2(n10156), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n10307), .ZN(n10164) );
  AOI21_X1 U12696 ( .B1(n8344), .B2(n10158), .A(n10157), .ZN(n10162) );
  AOI21_X1 U12697 ( .B1(n8343), .B2(n10160), .A(n10159), .ZN(n10161) );
  OAI22_X1 U12698 ( .A1(n10162), .A2(n15163), .B1(n15136), .B2(n10161), .ZN(
        n10163) );
  AOI211_X1 U12699 ( .C1(n15155), .C2(n10165), .A(n10164), .B(n10163), .ZN(
        n10166) );
  INV_X1 U12700 ( .A(n13497), .ZN(n14893) );
  INV_X1 U12701 ( .A(n10167), .ZN(n10168) );
  OAI222_X1 U12702 ( .A1(P2_U3088), .A2(n14893), .B1(n13873), .B2(n10168), 
        .C1(n13222), .C2(n13870), .ZN(P2_U3315) );
  OAI222_X1 U12703 ( .A1(n14478), .A2(n10169), .B1(n14480), .B2(n10168), .C1(
        n10259), .C2(P1_U3086), .ZN(P1_U3343) );
  OR2_X1 U12704 ( .A1(n10171), .A2(n10170), .ZN(n10173) );
  AND2_X1 U12705 ( .A1(n10173), .A2(n10172), .ZN(n10181) );
  INV_X1 U12706 ( .A(n10181), .ZN(n14347) );
  INV_X1 U12707 ( .A(n10614), .ZN(n10175) );
  NAND2_X1 U12708 ( .A1(n9548), .A2(n14345), .ZN(n10174) );
  NAND2_X1 U12709 ( .A1(n10175), .A2(n10174), .ZN(n14342) );
  AND2_X1 U12710 ( .A1(n14043), .A2(n14321), .ZN(n14338) );
  INV_X1 U12711 ( .A(n14338), .ZN(n10176) );
  OAI21_X1 U12712 ( .B1(n14342), .B2(n14326), .A(n10176), .ZN(n10183) );
  INV_X1 U12713 ( .A(n14319), .ZN(n14285) );
  INV_X1 U12714 ( .A(n14046), .ZN(n10182) );
  XNOR2_X1 U12715 ( .A(n14342), .B(n10177), .ZN(n10179) );
  MUX2_X1 U12716 ( .A(n10179), .B(n10178), .S(n14046), .Z(n10180) );
  OAI222_X1 U12717 ( .A1(n14285), .A2(n10182), .B1(n14155), .B2(n10181), .C1(
        n14282), .C2(n10180), .ZN(n14339) );
  AOI211_X1 U12718 ( .C1(n14381), .C2(n14347), .A(n10183), .B(n14339), .ZN(
        n10331) );
  OAI22_X1 U12719 ( .A1(n14468), .A2(n10184), .B1(n14849), .B2(n7518), .ZN(
        n10185) );
  INV_X1 U12720 ( .A(n10185), .ZN(n10186) );
  OAI21_X1 U12721 ( .B1(n10331), .B2(n6786), .A(n10186), .ZN(P1_U3462) );
  NAND2_X1 U12722 ( .A1(n12282), .A2(SI_0_), .ZN(n10190) );
  AND2_X2 U12723 ( .A1(n11392), .A2(n8621), .ZN(n10449) );
  NAND2_X1 U12724 ( .A1(n10449), .A2(n10188), .ZN(n10189) );
  OAI211_X1 U12725 ( .C1(n15105), .C2(n11392), .A(n10190), .B(n10189), .ZN(
        n10244) );
  INV_X1 U12726 ( .A(n10244), .ZN(n10500) );
  INV_X2 U12727 ( .A(n12328), .ZN(n12268) );
  NAND2_X1 U12728 ( .A1(n12268), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n10194) );
  NAND2_X1 U12729 ( .A1(n10235), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n10193) );
  NAND2_X1 U12730 ( .A1(n10454), .A2(P3_REG0_REG_0__SCAN_IN), .ZN(n10192) );
  NAND2_X1 U12731 ( .A1(n6495), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n10191) );
  NAND4_X2 U12732 ( .A1(n10194), .A2(n10193), .A3(n10192), .A4(n10191), .ZN(
        n15195) );
  NOR2_X2 U12733 ( .A1(n10500), .A2(n15195), .ZN(n12368) );
  NAND2_X1 U12734 ( .A1(n15195), .A2(n10500), .ZN(n12369) );
  INV_X1 U12735 ( .A(n12369), .ZN(n10195) );
  NOR2_X1 U12736 ( .A1(n12368), .A2(n10195), .ZN(n12511) );
  NAND2_X1 U12737 ( .A1(n10203), .A2(n10196), .ZN(n10198) );
  NAND2_X1 U12738 ( .A1(n11748), .A2(n11878), .ZN(n10197) );
  INV_X1 U12739 ( .A(P3_D_REG_0__SCAN_IN), .ZN(n10199) );
  NAND2_X1 U12740 ( .A1(n10200), .A2(n10199), .ZN(n10202) );
  NAND2_X1 U12741 ( .A1(n9808), .A2(n11878), .ZN(n10201) );
  INV_X1 U12742 ( .A(n10203), .ZN(n10215) );
  NOR2_X1 U12743 ( .A1(P3_D_REG_11__SCAN_IN), .A2(P3_D_REG_26__SCAN_IN), .ZN(
        n10207) );
  NOR4_X1 U12744 ( .A1(P3_D_REG_2__SCAN_IN), .A2(P3_D_REG_8__SCAN_IN), .A3(
        P3_D_REG_31__SCAN_IN), .A4(P3_D_REG_17__SCAN_IN), .ZN(n10206) );
  NOR4_X1 U12745 ( .A1(P3_D_REG_18__SCAN_IN), .A2(P3_D_REG_27__SCAN_IN), .A3(
        P3_D_REG_24__SCAN_IN), .A4(P3_D_REG_29__SCAN_IN), .ZN(n10205) );
  NOR4_X1 U12746 ( .A1(P3_D_REG_22__SCAN_IN), .A2(P3_D_REG_25__SCAN_IN), .A3(
        P3_D_REG_20__SCAN_IN), .A4(P3_D_REG_19__SCAN_IN), .ZN(n10204) );
  NAND4_X1 U12747 ( .A1(n10207), .A2(n10206), .A3(n10205), .A4(n10204), .ZN(
        n10213) );
  NOR4_X1 U12748 ( .A1(P3_D_REG_9__SCAN_IN), .A2(P3_D_REG_16__SCAN_IN), .A3(
        P3_D_REG_15__SCAN_IN), .A4(P3_D_REG_30__SCAN_IN), .ZN(n10211) );
  NOR4_X1 U12749 ( .A1(P3_D_REG_10__SCAN_IN), .A2(P3_D_REG_21__SCAN_IN), .A3(
        P3_D_REG_14__SCAN_IN), .A4(P3_D_REG_12__SCAN_IN), .ZN(n10210) );
  NOR4_X1 U12750 ( .A1(P3_D_REG_3__SCAN_IN), .A2(P3_D_REG_5__SCAN_IN), .A3(
        P3_D_REG_4__SCAN_IN), .A4(P3_D_REG_7__SCAN_IN), .ZN(n10209) );
  NOR4_X1 U12751 ( .A1(P3_D_REG_13__SCAN_IN), .A2(P3_D_REG_28__SCAN_IN), .A3(
        P3_D_REG_23__SCAN_IN), .A4(P3_D_REG_6__SCAN_IN), .ZN(n10208) );
  NAND4_X1 U12752 ( .A1(n10211), .A2(n10210), .A3(n10209), .A4(n10208), .ZN(
        n10212) );
  NOR2_X1 U12753 ( .A1(n10213), .A2(n10212), .ZN(n10214) );
  NAND3_X1 U12754 ( .A1(n10495), .A2(n10471), .A3(n10472), .ZN(n13294) );
  INV_X1 U12755 ( .A(n10482), .ZN(n10218) );
  NAND2_X1 U12756 ( .A1(n8311), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n10217) );
  INV_X1 U12757 ( .A(n10779), .ZN(n10481) );
  NAND2_X1 U12758 ( .A1(n10218), .A2(n12541), .ZN(n13292) );
  INV_X1 U12759 ( .A(n10471), .ZN(n13319) );
  NAND3_X1 U12760 ( .A1(n13319), .A2(n13317), .A3(n10472), .ZN(n13298) );
  NAND2_X1 U12761 ( .A1(n12367), .A2(n10779), .ZN(n10490) );
  INV_X1 U12762 ( .A(n10490), .ZN(n10219) );
  XNOR2_X1 U12763 ( .A(n13053), .B(n10219), .ZN(n10221) );
  NAND2_X1 U12764 ( .A1(n12367), .A2(n12345), .ZN(n10220) );
  NAND2_X1 U12765 ( .A1(n10221), .A2(n10220), .ZN(n13291) );
  NAND2_X1 U12766 ( .A1(n13291), .A2(n15261), .ZN(n10483) );
  OAI22_X1 U12767 ( .A1(n13294), .A2(n13292), .B1(n13298), .B2(n10483), .ZN(
        n10222) );
  INV_X1 U12768 ( .A(n13292), .ZN(n10223) );
  NAND2_X1 U12769 ( .A1(n13294), .A2(n10223), .ZN(n10226) );
  NAND2_X1 U12770 ( .A1(n13298), .A2(n13291), .ZN(n10224) );
  NAND2_X1 U12771 ( .A1(n10779), .A2(n12345), .ZN(n10476) );
  NAND2_X1 U12772 ( .A1(n11001), .A2(n10476), .ZN(n10488) );
  NAND4_X1 U12773 ( .A1(n10226), .A2(n10225), .A3(n10224), .A4(n10488), .ZN(
        n10227) );
  NAND2_X1 U12774 ( .A1(n10227), .A2(P3_STATE_REG_SCAN_IN), .ZN(n10230) );
  INV_X1 U12775 ( .A(n10476), .ZN(n12505) );
  AND2_X1 U12776 ( .A1(n13295), .A2(n12505), .ZN(n10233) );
  INV_X1 U12777 ( .A(n13297), .ZN(n10228) );
  NAND2_X1 U12778 ( .A1(n13294), .A2(n10228), .ZN(n10229) );
  NAND2_X1 U12779 ( .A1(n10230), .A2(n10229), .ZN(n10542) );
  OR2_X1 U12780 ( .A1(n10542), .A2(n10231), .ZN(n10461) );
  NAND2_X1 U12781 ( .A1(n10461), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n10246) );
  NAND2_X1 U12782 ( .A1(n10232), .A2(n11392), .ZN(n12545) );
  NAND2_X1 U12783 ( .A1(n10233), .A2(n13040), .ZN(n10234) );
  INV_X1 U12784 ( .A(n12328), .ZN(n12155) );
  NAND2_X1 U12785 ( .A1(n12155), .A2(P3_REG2_REG_1__SCAN_IN), .ZN(n10240) );
  NAND2_X1 U12786 ( .A1(n10235), .A2(P3_REG3_REG_1__SCAN_IN), .ZN(n10239) );
  INV_X1 U12787 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n10236) );
  AND4_X2 U12788 ( .A1(n10240), .A2(n10239), .A3(n10238), .A4(n10237), .ZN(
        n10444) );
  INV_X1 U12789 ( .A(n10242), .ZN(n10241) );
  OR2_X1 U12790 ( .A1(n13298), .A2(n10241), .ZN(n10243) );
  AOI22_X1 U12791 ( .A1(n12733), .A2(n10297), .B1(n12739), .B2(n10244), .ZN(
        n10245) );
  OAI211_X1 U12792 ( .C1(n12511), .C2(n12741), .A(n10246), .B(n10245), .ZN(
        P3_U3172) );
  INV_X1 U12793 ( .A(P3_DATAO_REG_23__SCAN_IN), .ZN(n13219) );
  NAND2_X1 U12794 ( .A1(n11534), .A2(n11533), .ZN(n11675) );
  NAND2_X1 U12795 ( .A1(n11945), .A2(n11944), .ZN(n11979) );
  NOR2_X1 U12796 ( .A1(n12207), .A2(n12637), .ZN(n10247) );
  OR2_X1 U12797 ( .A1(n12222), .A2(n10247), .ZN(n12958) );
  NAND2_X1 U12798 ( .A1(n12958), .A2(n10235), .ZN(n10253) );
  INV_X1 U12799 ( .A(P3_REG2_REG_23__SCAN_IN), .ZN(n10250) );
  NAND2_X1 U12800 ( .A1(n6491), .A2(P3_REG1_REG_23__SCAN_IN), .ZN(n10249) );
  NAND2_X1 U12801 ( .A1(n10454), .A2(P3_REG0_REG_23__SCAN_IN), .ZN(n10248) );
  OAI211_X1 U12802 ( .C1(n6487), .C2(n10250), .A(n10249), .B(n10248), .ZN(
        n10251) );
  INV_X1 U12803 ( .A(n10251), .ZN(n10252) );
  NAND2_X1 U12804 ( .A1(n12967), .A2(P3_U3897), .ZN(n10254) );
  OAI21_X1 U12805 ( .B1(P3_U3897), .B2(n13219), .A(n10254), .ZN(P3_U3514) );
  INV_X1 U12806 ( .A(n10255), .ZN(n10256) );
  NOR2_X1 U12807 ( .A1(n10257), .A2(n10256), .ZN(n10310) );
  XNOR2_X1 U12808 ( .A(n10316), .B(P1_REG1_REG_13__SCAN_IN), .ZN(n10309) );
  XNOR2_X1 U12809 ( .A(n10310), .B(n10309), .ZN(n10266) );
  NAND2_X1 U12810 ( .A1(P1_U3086), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n12024)
         );
  AOI21_X1 U12811 ( .B1(n11484), .B2(n10259), .A(n10258), .ZN(n10261) );
  INV_X1 U12812 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n11607) );
  MUX2_X1 U12813 ( .A(n11607), .B(P1_REG2_REG_13__SCAN_IN), .S(n10316), .Z(
        n10260) );
  NAND2_X1 U12814 ( .A1(n10261), .A2(n10260), .ZN(n10315) );
  OAI211_X1 U12815 ( .C1(n10261), .C2(n10260), .A(n14113), .B(n10315), .ZN(
        n10262) );
  NAND2_X1 U12816 ( .A1(n12024), .A2(n10262), .ZN(n10264) );
  NOR2_X1 U12817 ( .A1(n14811), .A2(n10316), .ZN(n10263) );
  AOI211_X1 U12818 ( .C1(n14088), .C2(P1_ADDR_REG_13__SCAN_IN), .A(n10264), 
        .B(n10263), .ZN(n10265) );
  OAI21_X1 U12819 ( .B1(n10266), .B2(n14809), .A(n10265), .ZN(P1_U3256) );
  INV_X1 U12820 ( .A(n10267), .ZN(n10268) );
  NOR2_X1 U12821 ( .A1(n10269), .A2(n10268), .ZN(n10273) );
  XNOR2_X1 U12822 ( .A(n15058), .B(n9992), .ZN(n10271) );
  NAND2_X1 U12823 ( .A1(n13445), .A2(n12605), .ZN(n10270) );
  NAND2_X1 U12824 ( .A1(n10271), .A2(n10270), .ZN(n10386) );
  OAI21_X1 U12825 ( .B1(n10271), .B2(n10270), .A(n10386), .ZN(n10272) );
  AOI21_X1 U12826 ( .B1(n10273), .B2(n10272), .A(n10388), .ZN(n10279) );
  NAND2_X1 U12827 ( .A1(n13524), .A2(n13444), .ZN(n10275) );
  NAND2_X1 U12828 ( .A1(n13420), .A2(n13446), .ZN(n10274) );
  NAND2_X1 U12829 ( .A1(n10275), .A2(n10274), .ZN(n15057) );
  AOI21_X1 U12830 ( .B1(n13374), .B2(n15057), .A(n10276), .ZN(n10278) );
  AOI22_X1 U12831 ( .A1(n13426), .A2(n15058), .B1(n13422), .B2(n10745), .ZN(
        n10277) );
  OAI211_X1 U12832 ( .C1(n10279), .C2(n13428), .A(n10278), .B(n10277), .ZN(
        P2_U3199) );
  INV_X1 U12833 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n10281) );
  INV_X1 U12834 ( .A(n10280), .ZN(n10282) );
  OAI222_X1 U12835 ( .A1(n13870), .A2(n10281), .B1(n13873), .B2(n10282), .C1(
        n13498), .C2(P2_U3088), .ZN(P2_U3314) );
  OAI222_X1 U12836 ( .A1(n14478), .A2(n10283), .B1(n14480), .B2(n10282), .C1(
        n10316), .C2(P1_U3086), .ZN(P1_U3342) );
  INV_X1 U12837 ( .A(n10461), .ZN(n10308) );
  NAND2_X1 U12838 ( .A1(n12282), .A2(SI_1_), .ZN(n10286) );
  NAND2_X1 U12839 ( .A1(n10449), .A2(n10284), .ZN(n10285) );
  INV_X1 U12840 ( .A(n15195), .ZN(n10293) );
  OR2_X1 U12841 ( .A1(n13297), .A2(n12545), .ZN(n10287) );
  NAND2_X1 U12842 ( .A1(n12155), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n10292) );
  NAND2_X1 U12843 ( .A1(n10235), .A2(P3_REG3_REG_2__SCAN_IN), .ZN(n10291) );
  NAND2_X1 U12844 ( .A1(n10454), .A2(P3_REG0_REG_2__SCAN_IN), .ZN(n10290) );
  NAND2_X1 U12845 ( .A1(n6495), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n10289) );
  OAI22_X1 U12846 ( .A1(n10293), .A2(n12736), .B1(n12723), .B2(n15198), .ZN(
        n10294) );
  AOI21_X1 U12847 ( .B1(n15190), .B2(n12739), .A(n10294), .ZN(n10306) );
  NAND2_X1 U12848 ( .A1(n12367), .A2(n12539), .ZN(n10295) );
  NAND2_X1 U12849 ( .A1(n10295), .A2(n10779), .ZN(n10296) );
  NAND2_X1 U12850 ( .A1(n10444), .A2(n15190), .ZN(n12374) );
  NAND2_X1 U12851 ( .A1(n10299), .A2(n10298), .ZN(n10303) );
  NAND2_X1 U12852 ( .A1(n15195), .A2(n10244), .ZN(n15191) );
  INV_X1 U12853 ( .A(n15191), .ZN(n10300) );
  NAND2_X1 U12854 ( .A1(n12368), .A2(n12375), .ZN(n10991) );
  OAI21_X1 U12855 ( .B1(n10300), .B2(n6486), .A(n10991), .ZN(n10301) );
  NAND2_X1 U12856 ( .A1(n10303), .A2(n10301), .ZN(n10446) );
  INV_X1 U12857 ( .A(n12368), .ZN(n15203) );
  NAND3_X1 U12858 ( .A1(n15203), .A2(n15202), .A3(n12151), .ZN(n10302) );
  OAI211_X1 U12859 ( .C1(n10303), .C2(n15191), .A(n10446), .B(n10302), .ZN(
        n10304) );
  NAND2_X1 U12860 ( .A1(n10304), .A2(n12709), .ZN(n10305) );
  OAI211_X1 U12861 ( .C1(n10308), .C2(n10307), .A(n10306), .B(n10305), .ZN(
        P3_U3162) );
  INV_X1 U12862 ( .A(n11172), .ZN(n11184) );
  AOI22_X1 U12863 ( .A1(n11172), .A2(n11183), .B1(P1_REG1_REG_14__SCAN_IN), 
        .B2(n11184), .ZN(n10314) );
  NAND2_X1 U12864 ( .A1(n10310), .A2(n10309), .ZN(n10311) );
  OAI21_X1 U12865 ( .B1(n10316), .B2(n10312), .A(n10311), .ZN(n10313) );
  NOR2_X1 U12866 ( .A1(n10314), .A2(n10313), .ZN(n11182) );
  AOI21_X1 U12867 ( .B1(n10314), .B2(n10313), .A(n11182), .ZN(n10322) );
  OAI21_X1 U12868 ( .B1(n11607), .B2(n10316), .A(n10315), .ZN(n10318) );
  XNOR2_X1 U12869 ( .A(n11184), .B(P1_REG2_REG_14__SCAN_IN), .ZN(n10317) );
  NAND2_X1 U12870 ( .A1(n10317), .A2(n10318), .ZN(n11173) );
  OAI211_X1 U12871 ( .C1(n10318), .C2(n10317), .A(n14113), .B(n11173), .ZN(
        n10321) );
  INV_X1 U12872 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n14512) );
  NAND2_X1 U12873 ( .A1(P1_U3086), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n13889)
         );
  OAI21_X1 U12874 ( .B1(n14815), .B2(n14512), .A(n13889), .ZN(n10319) );
  AOI21_X1 U12875 ( .B1(n14108), .B2(n11172), .A(n10319), .ZN(n10320) );
  OAI211_X1 U12876 ( .C1(n10322), .C2(n14809), .A(n10321), .B(n10320), .ZN(
        P1_U3257) );
  AOI22_X1 U12877 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(
        P2_DATAO_REG_17__SCAN_IN), .B1(n11123), .B2(n13208), .ZN(n10325) );
  INV_X1 U12878 ( .A(n10325), .ZN(n10326) );
  XNOR2_X1 U12879 ( .A(n10465), .B(n10326), .ZN(n12137) );
  INV_X1 U12880 ( .A(n12137), .ZN(n10329) );
  OAI222_X1 U12881 ( .A1(n13333), .A2(n10329), .B1(n13335), .B2(n10328), .C1(
        n10327), .C2(P3_U3151), .ZN(P3_U3278) );
  AOI22_X1 U12882 ( .A1(n14375), .A2(n14345), .B1(n14854), .B2(
        P1_REG1_REG_1__SCAN_IN), .ZN(n10330) );
  OAI21_X1 U12883 ( .B1(n10331), .B2(n14854), .A(n10330), .ZN(P1_U3529) );
  AOI211_X1 U12884 ( .C1(n10334), .C2(n10333), .A(n14022), .B(n10332), .ZN(
        n10338) );
  INV_X1 U12885 ( .A(n14011), .ZN(n13985) );
  MUX2_X1 U12886 ( .A(n13989), .B(P1_STATE_REG_SCAN_IN), .S(
        P1_REG3_REG_3__SCAN_IN), .Z(n10336) );
  AOI22_X1 U12887 ( .A1(n13987), .A2(n14041), .B1(n10605), .B2(n14018), .ZN(
        n10335) );
  OAI211_X1 U12888 ( .C1(n10510), .C2(n13985), .A(n10336), .B(n10335), .ZN(
        n10337) );
  OR2_X1 U12889 ( .A1(n10338), .A2(n10337), .ZN(P1_U3218) );
  INV_X1 U12890 ( .A(n15015), .ZN(n10673) );
  NOR2_X1 U12891 ( .A1(n10339), .A2(n10673), .ZN(n10340) );
  AND2_X1 U12892 ( .A1(n10677), .A2(n10340), .ZN(n10382) );
  NAND2_X1 U12893 ( .A1(n15016), .A2(n10341), .ZN(n10675) );
  AND2_X1 U12894 ( .A1(n9205), .A2(n14990), .ZN(n10981) );
  OAI22_X1 U12895 ( .A1(n10981), .A2(n10349), .B1(n10987), .B2(n9998), .ZN(
        n10766) );
  INV_X1 U12896 ( .A(n13448), .ZN(n10353) );
  NAND2_X1 U12897 ( .A1(n10353), .A2(n6747), .ZN(n10344) );
  NAND2_X1 U12898 ( .A1(n10345), .A2(n10344), .ZN(n10697) );
  INV_X1 U12899 ( .A(n15058), .ZN(n10748) );
  INV_X1 U12900 ( .A(n10574), .ZN(n10883) );
  INV_X1 U12901 ( .A(n13444), .ZN(n10366) );
  XNOR2_X1 U12902 ( .A(n10706), .B(n10705), .ZN(n10689) );
  NAND2_X1 U12903 ( .A1(n10978), .A2(n10349), .ZN(n10352) );
  NAND2_X1 U12904 ( .A1(n10350), .A2(n10987), .ZN(n10351) );
  NAND2_X1 U12905 ( .A1(n10352), .A2(n10351), .ZN(n10763) );
  NAND2_X1 U12906 ( .A1(n10763), .A2(n10343), .ZN(n10355) );
  NAND2_X1 U12907 ( .A1(n10353), .A2(n10769), .ZN(n10354) );
  INV_X1 U12908 ( .A(n10356), .ZN(n10702) );
  NAND2_X1 U12909 ( .A1(n10701), .A2(n10702), .ZN(n10359) );
  NAND2_X1 U12910 ( .A1(n10375), .A2(n10357), .ZN(n10358) );
  NAND2_X1 U12911 ( .A1(n10359), .A2(n10358), .ZN(n14972) );
  NAND2_X1 U12912 ( .A1(n14972), .A2(n14971), .ZN(n10362) );
  INV_X1 U12913 ( .A(n13446), .ZN(n10360) );
  NAND2_X1 U12914 ( .A1(n15049), .A2(n10360), .ZN(n10361) );
  NAND2_X1 U12915 ( .A1(n10362), .A2(n10361), .ZN(n10750) );
  NAND2_X1 U12916 ( .A1(n10750), .A2(n10751), .ZN(n10365) );
  NAND2_X1 U12917 ( .A1(n15058), .A2(n10363), .ZN(n10364) );
  NAND2_X1 U12918 ( .A1(n10365), .A2(n10364), .ZN(n10568) );
  NAND2_X1 U12919 ( .A1(n10574), .A2(n10366), .ZN(n10367) );
  XOR2_X1 U12920 ( .A(n10705), .B(n10711), .Z(n10374) );
  NAND2_X1 U12921 ( .A1(n6713), .A2(n10368), .ZN(n10371) );
  NAND2_X1 U12922 ( .A1(n13524), .A2(n13442), .ZN(n10373) );
  NAND2_X1 U12923 ( .A1(n13420), .A2(n13444), .ZN(n10372) );
  NAND2_X1 U12924 ( .A1(n10373), .A2(n10372), .ZN(n10586) );
  AOI21_X1 U12925 ( .B1(n10374), .B2(n15064), .A(n10586), .ZN(n10685) );
  INV_X1 U12926 ( .A(n10572), .ZN(n10377) );
  INV_X1 U12927 ( .A(n10709), .ZN(n10682) );
  NAND2_X1 U12928 ( .A1(n10682), .A2(n10572), .ZN(n10720) );
  INV_X1 U12929 ( .A(n10720), .ZN(n10376) );
  AOI211_X1 U12930 ( .C1(n10709), .C2(n10377), .A(n12610), .B(n10376), .ZN(
        n10684) );
  AOI21_X1 U12931 ( .B1(n15069), .B2(n10709), .A(n10684), .ZN(n10378) );
  OAI211_X1 U12932 ( .C1(n10689), .C2(n15061), .A(n10685), .B(n10378), .ZN(
        n10383) );
  NAND2_X1 U12933 ( .A1(n10383), .A2(n15096), .ZN(n10379) );
  OAI21_X1 U12934 ( .B1(n15096), .B2(n9840), .A(n10379), .ZN(P2_U3506) );
  INV_X1 U12935 ( .A(n15012), .ZN(n10380) );
  NOR2_X1 U12936 ( .A1(n10675), .A2(n10380), .ZN(n10381) );
  INV_X1 U12937 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n10385) );
  NAND2_X1 U12938 ( .A1(n10383), .A2(n15066), .ZN(n10384) );
  OAI21_X1 U12939 ( .B1(n15066), .B2(n10385), .A(n10384), .ZN(P2_U3451) );
  INV_X1 U12940 ( .A(n10386), .ZN(n10387) );
  XNOR2_X1 U12941 ( .A(n10574), .B(n12611), .ZN(n10582) );
  NAND2_X1 U12942 ( .A1(n13444), .A2(n12610), .ZN(n10581) );
  XNOR2_X1 U12943 ( .A(n10582), .B(n10581), .ZN(n10584) );
  XNOR2_X1 U12944 ( .A(n10585), .B(n10584), .ZN(n10396) );
  NAND2_X1 U12945 ( .A1(n13524), .A2(n13443), .ZN(n10391) );
  NAND2_X1 U12946 ( .A1(n13420), .A2(n13445), .ZN(n10390) );
  NAND2_X1 U12947 ( .A1(n10391), .A2(n10390), .ZN(n10570) );
  INV_X1 U12948 ( .A(n10392), .ZN(n10393) );
  AOI21_X1 U12949 ( .B1(n13374), .B2(n10570), .A(n10393), .ZN(n10395) );
  AOI22_X1 U12950 ( .A1(n13426), .A2(n10574), .B1(n13422), .B2(n10881), .ZN(
        n10394) );
  OAI211_X1 U12951 ( .C1(n10396), .C2(n13428), .A(n10395), .B(n10394), .ZN(
        P2_U3211) );
  AOI21_X1 U12952 ( .B1(n10399), .B2(n10398), .A(n10397), .ZN(n10412) );
  AOI21_X1 U12953 ( .B1(n6651), .B2(n10401), .A(n10400), .ZN(n10405) );
  INV_X1 U12954 ( .A(P3_REG3_REG_6__SCAN_IN), .ZN(n10402) );
  NOR2_X1 U12955 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10402), .ZN(n11118) );
  NOR2_X1 U12956 ( .A1(n15139), .A2(n11074), .ZN(n10403) );
  AOI211_X1 U12957 ( .C1(n15097), .C2(P3_ADDR_REG_6__SCAN_IN), .A(n11118), .B(
        n10403), .ZN(n10404) );
  OAI21_X1 U12958 ( .B1(n10405), .B2(n15136), .A(n10404), .ZN(n10410) );
  NAND3_X1 U12959 ( .A1(n15133), .A2(n10407), .A3(n10406), .ZN(n10408) );
  AOI21_X1 U12960 ( .B1(n15150), .B2(n10408), .A(n15131), .ZN(n10409) );
  NOR2_X1 U12961 ( .A1(n10410), .A2(n10409), .ZN(n10411) );
  OAI21_X1 U12962 ( .B1(n10412), .B2(n15163), .A(n10411), .ZN(P3_U3188) );
  AOI21_X1 U12963 ( .B1(n10415), .B2(n10414), .A(n10413), .ZN(n10417) );
  AOI22_X1 U12964 ( .A1(n15097), .A2(P3_ADDR_REG_2__SCAN_IN), .B1(
        P3_REG3_REG_2__SCAN_IN), .B2(P3_U3151), .ZN(n10416) );
  OAI21_X1 U12965 ( .B1(n10417), .B2(n15136), .A(n10416), .ZN(n10427) );
  AOI21_X1 U12966 ( .B1(n10419), .B2(n10418), .A(n6654), .ZN(n10420) );
  NOR2_X1 U12967 ( .A1(n15163), .A2(n10420), .ZN(n10426) );
  NAND3_X1 U12968 ( .A1(n10423), .A2(n10422), .A3(n10421), .ZN(n10424) );
  AOI21_X1 U12969 ( .B1(n10431), .B2(n10424), .A(n15131), .ZN(n10425) );
  NOR3_X1 U12970 ( .A1(n10427), .A2(n10426), .A3(n10425), .ZN(n10428) );
  OAI21_X1 U12971 ( .B1(n6496), .B2(n15139), .A(n10428), .ZN(P3_U3184) );
  NAND3_X1 U12972 ( .A1(n10431), .A2(n10430), .A3(n10429), .ZN(n10432) );
  AOI21_X1 U12973 ( .B1(n15118), .B2(n10432), .A(n15131), .ZN(n10442) );
  AOI21_X1 U12974 ( .B1(n11013), .B2(n10434), .A(n10433), .ZN(n10440) );
  INV_X1 U12975 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n11014) );
  NOR2_X1 U12976 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11014), .ZN(n10554) );
  AOI21_X1 U12977 ( .B1(n8362), .B2(n10436), .A(n10435), .ZN(n10437) );
  NOR2_X1 U12978 ( .A1(n15136), .A2(n10437), .ZN(n10438) );
  AOI211_X1 U12979 ( .C1(n15097), .C2(P3_ADDR_REG_3__SCAN_IN), .A(n10554), .B(
        n10438), .ZN(n10439) );
  OAI21_X1 U12980 ( .B1(n10440), .B2(n15163), .A(n10439), .ZN(n10441) );
  AOI211_X1 U12981 ( .C1(n15153), .C2(n10549), .A(n10442), .B(n10441), .ZN(
        n10443) );
  INV_X1 U12982 ( .A(n10443), .ZN(P3_U3185) );
  MUX2_X1 U12983 ( .A(n15176), .B(n12374), .S(n6486), .Z(n10445) );
  NAND2_X1 U12984 ( .A1(n12282), .A2(n10447), .ZN(n10453) );
  NAND2_X1 U12985 ( .A1(n10449), .A2(n10448), .ZN(n10452) );
  OR2_X1 U12986 ( .A1(n11392), .A2(n10450), .ZN(n10451) );
  XNOR2_X1 U12987 ( .A(n6486), .B(n10992), .ZN(n10557) );
  INV_X1 U12988 ( .A(n10993), .ZN(n12755) );
  XNOR2_X1 U12989 ( .A(n10557), .B(n12755), .ZN(n10555) );
  XOR2_X1 U12990 ( .A(n10556), .B(n10555), .Z(n10463) );
  INV_X1 U12991 ( .A(n10992), .ZN(n15184) );
  NAND2_X1 U12992 ( .A1(n12268), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n10458) );
  NAND2_X1 U12993 ( .A1(n10235), .A2(n11014), .ZN(n10457) );
  NAND2_X1 U12994 ( .A1(n10454), .A2(P3_REG0_REG_3__SCAN_IN), .ZN(n10456) );
  NAND2_X1 U12995 ( .A1(n6495), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n10455) );
  AND4_X2 U12996 ( .A1(n10458), .A2(n10457), .A3(n10456), .A4(n10455), .ZN(
        n15172) );
  INV_X1 U12997 ( .A(n15172), .ZN(n12754) );
  AOI22_X1 U12998 ( .A1(n12720), .A2(n10297), .B1(n12733), .B2(n12754), .ZN(
        n10459) );
  OAI21_X1 U12999 ( .B1(n12717), .B2(n15184), .A(n10459), .ZN(n10460) );
  AOI21_X1 U13000 ( .B1(P3_REG3_REG_2__SCAN_IN), .B2(n10461), .A(n10460), .ZN(
        n10462) );
  OAI21_X1 U13001 ( .B1(n10463), .B2(n12741), .A(n10462), .ZN(P3_U3177) );
  NAND2_X1 U13002 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(n11123), .ZN(n10464) );
  INV_X1 U13003 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n11380) );
  AOI22_X1 U13004 ( .A1(P2_DATAO_REG_18__SCAN_IN), .A2(n11380), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(n11378), .ZN(n10466) );
  INV_X1 U13005 ( .A(n10466), .ZN(n10467) );
  XNOR2_X1 U13006 ( .A(n10579), .B(n10467), .ZN(n12148) );
  INV_X1 U13007 ( .A(n12148), .ZN(n10470) );
  OAI222_X1 U13008 ( .A1(n13333), .A2(n10470), .B1(n13335), .B2(n10469), .C1(
        n10468), .C2(P3_U3151), .ZN(P3_U3277) );
  XNOR2_X1 U13009 ( .A(n10471), .B(n13317), .ZN(n10474) );
  INV_X1 U13010 ( .A(n10488), .ZN(n10475) );
  NOR2_X1 U13011 ( .A1(n13317), .A2(n10475), .ZN(n10478) );
  NAND2_X1 U13012 ( .A1(n10482), .A2(n10476), .ZN(n10491) );
  INV_X1 U13013 ( .A(n10491), .ZN(n10477) );
  INV_X1 U13014 ( .A(n13053), .ZN(n12546) );
  NAND2_X1 U13015 ( .A1(n10477), .A2(n12546), .ZN(n10999) );
  NAND2_X1 U13016 ( .A1(n10999), .A2(n12481), .ZN(n10489) );
  MUX2_X1 U13017 ( .A(n13317), .B(n10478), .S(n10489), .Z(n10479) );
  OR2_X1 U13018 ( .A1(n15261), .A2(n15206), .ZN(n10480) );
  INV_X1 U13019 ( .A(n12367), .ZN(n12363) );
  NAND2_X1 U13020 ( .A1(n12363), .A2(n10481), .ZN(n12347) );
  AOI21_X1 U13021 ( .B1(n15178), .B2(n10483), .A(n12511), .ZN(n10484) );
  AOI21_X1 U13022 ( .B1(n13040), .B2(n10297), .A(n10484), .ZN(n10499) );
  MUX2_X1 U13023 ( .A(n15099), .B(n10499), .S(n15211), .Z(n10487) );
  NAND2_X1 U13024 ( .A1(n15208), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n10486) );
  OAI211_X1 U13025 ( .C1(n10500), .C2(n13047), .A(n10487), .B(n10486), .ZN(
        P3_U3233) );
  AND2_X1 U13026 ( .A1(n10489), .A2(n10488), .ZN(n10494) );
  AOI22_X1 U13027 ( .A1(n10491), .A2(n12367), .B1(n13053), .B2(n10490), .ZN(
        n10492) );
  NAND2_X1 U13028 ( .A1(n10495), .A2(n10492), .ZN(n10493) );
  OAI21_X1 U13029 ( .B1(n10495), .B2(n10494), .A(n10493), .ZN(n10496) );
  INV_X1 U13030 ( .A(n10496), .ZN(n10497) );
  OAI21_X1 U13031 ( .B1(n10500), .B2(n15261), .A(n10499), .ZN(n13316) );
  NAND2_X1 U13032 ( .A1(n13316), .A2(n15281), .ZN(n10501) );
  OAI21_X1 U13033 ( .B1(n15281), .B2(n13182), .A(n10501), .ZN(P3_U3459) );
  OAI21_X1 U13034 ( .B1(n10504), .B2(n10503), .A(n10502), .ZN(n10505) );
  INV_X1 U13035 ( .A(n10505), .ZN(n10608) );
  OAI21_X1 U13036 ( .B1(n10509), .B2(n10508), .A(n10507), .ZN(n10513) );
  INV_X1 U13037 ( .A(n14321), .ZN(n14287) );
  OAI22_X1 U13038 ( .A1(n10510), .A2(n14285), .B1(n10900), .B2(n14287), .ZN(
        n10512) );
  NOR2_X1 U13039 ( .A1(n10608), .A2(n14155), .ZN(n10511) );
  AOI211_X1 U13040 ( .C1(n14324), .C2(n10513), .A(n10512), .B(n10511), .ZN(
        n10599) );
  AOI21_X1 U13041 ( .B1(n10613), .B2(n10605), .A(n14326), .ZN(n10514) );
  NAND2_X1 U13042 ( .A1(n10514), .A2(n10831), .ZN(n10603) );
  OAI211_X1 U13043 ( .C1(n10608), .C2(n10515), .A(n10599), .B(n10603), .ZN(
        n10520) );
  OAI22_X1 U13044 ( .A1(n14423), .A2(n10518), .B1(n14856), .B2(n9789), .ZN(
        n10516) );
  AOI21_X1 U13045 ( .B1(n10520), .B2(n14856), .A(n10516), .ZN(n10517) );
  INV_X1 U13046 ( .A(n10517), .ZN(P1_U3531) );
  OAI22_X1 U13047 ( .A1(n14468), .A2(n10518), .B1(n14849), .B2(n7546), .ZN(
        n10519) );
  AOI21_X1 U13048 ( .B1(n10520), .B2(n14849), .A(n10519), .ZN(n10521) );
  INV_X1 U13049 ( .A(n10521), .ZN(P1_U3468) );
  INV_X1 U13050 ( .A(n10522), .ZN(n10525) );
  OAI222_X1 U13051 ( .A1(n14478), .A2(n10523), .B1(n14480), .B2(n10525), .C1(
        n11184), .C2(P1_U3086), .ZN(P1_U3341) );
  INV_X1 U13052 ( .A(n14918), .ZN(n13499) );
  OAI222_X1 U13053 ( .A1(P2_U3088), .A2(n13499), .B1(n13873), .B2(n10525), 
        .C1(n10524), .C2(n13870), .ZN(P2_U3313) );
  AOI21_X1 U13054 ( .B1(n10528), .B2(n10527), .A(n10526), .ZN(n10540) );
  NAND2_X1 U13055 ( .A1(n10530), .A2(n10529), .ZN(n10531) );
  OAI21_X1 U13056 ( .B1(n15152), .B2(n10531), .A(n10856), .ZN(n10538) );
  AND2_X1 U13057 ( .A1(P3_U3151), .A2(P3_REG3_REG_8__SCAN_IN), .ZN(n11373) );
  AOI21_X1 U13058 ( .B1(n15097), .B2(P3_ADDR_REG_8__SCAN_IN), .A(n11373), .ZN(
        n10532) );
  OAI21_X1 U13059 ( .B1(n15139), .B2(n11206), .A(n10532), .ZN(n10537) );
  AOI21_X1 U13060 ( .B1(n10534), .B2(n10533), .A(n6645), .ZN(n10535) );
  NOR2_X1 U13061 ( .A1(n10535), .A2(n15136), .ZN(n10536) );
  AOI211_X1 U13062 ( .C1(n15155), .C2(n10538), .A(n10537), .B(n10536), .ZN(
        n10539) );
  OAI21_X1 U13063 ( .B1(n10540), .B2(n15163), .A(n10539), .ZN(P3_U3190) );
  INV_X1 U13064 ( .A(n12549), .ZN(n10541) );
  INV_X1 U13065 ( .A(n12732), .ZN(n11596) );
  NAND2_X1 U13066 ( .A1(n12268), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n10546) );
  NAND2_X1 U13067 ( .A1(n6495), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n10545) );
  XNOR2_X1 U13068 ( .A(P3_REG3_REG_4__SCAN_IN), .B(P3_REG3_REG_3__SCAN_IN), 
        .ZN(n10795) );
  NAND2_X1 U13069 ( .A1(n10235), .A2(n10795), .ZN(n10544) );
  NAND2_X1 U13070 ( .A1(n10454), .A2(P3_REG0_REG_4__SCAN_IN), .ZN(n10543) );
  NAND2_X1 U13071 ( .A1(n12282), .A2(n10547), .ZN(n10552) );
  NAND2_X1 U13072 ( .A1(n10449), .A2(n10548), .ZN(n10551) );
  OR2_X1 U13073 ( .A1(n11392), .A2(n10549), .ZN(n10550) );
  INV_X1 U13074 ( .A(n15223), .ZN(n10994) );
  OAI22_X1 U13075 ( .A1(n12717), .A2(n10994), .B1(n15198), .B2(n12736), .ZN(
        n10553) );
  AOI211_X1 U13076 ( .C1(n12733), .C2(n12753), .A(n10554), .B(n10553), .ZN(
        n10566) );
  NAND2_X1 U13077 ( .A1(n10556), .A2(n10555), .ZN(n10559) );
  NAND2_X1 U13078 ( .A1(n10557), .A2(n15198), .ZN(n10558) );
  XNOR2_X1 U13079 ( .A(n10560), .B(n15223), .ZN(n10801) );
  XNOR2_X1 U13080 ( .A(n10801), .B(n15172), .ZN(n10562) );
  AOI21_X1 U13081 ( .B1(n10561), .B2(n10562), .A(n12741), .ZN(n10564) );
  NAND2_X1 U13082 ( .A1(n10564), .A2(n10804), .ZN(n10565) );
  OAI211_X1 U13083 ( .C1(P3_REG3_REG_3__SCAN_IN), .C2(n11596), .A(n10566), .B(
        n10565), .ZN(P3_U3158) );
  INV_X1 U13084 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10577) );
  XNOR2_X1 U13085 ( .A(n10567), .B(n10569), .ZN(n10890) );
  XNOR2_X1 U13086 ( .A(n10568), .B(n10569), .ZN(n10571) );
  AOI21_X1 U13087 ( .B1(n10571), .B2(n15064), .A(n10570), .ZN(n10886) );
  INV_X1 U13088 ( .A(n10744), .ZN(n10573) );
  AOI211_X1 U13089 ( .C1(n10574), .C2(n10573), .A(n12605), .B(n10572), .ZN(
        n10885) );
  AOI21_X1 U13090 ( .B1(n15069), .B2(n10574), .A(n10885), .ZN(n10575) );
  OAI211_X1 U13091 ( .C1(n10890), .C2(n15061), .A(n10886), .B(n10575), .ZN(
        n13845) );
  NAND2_X1 U13092 ( .A1(n13845), .A2(n15066), .ZN(n10576) );
  OAI21_X1 U13093 ( .B1(n15066), .B2(n10577), .A(n10576), .ZN(P2_U3448) );
  NAND2_X1 U13094 ( .A1(P2_DATAO_REG_18__SCAN_IN), .A2(n11380), .ZN(n10578) );
  AOI22_X1 U13095 ( .A1(n10579), .A2(n10578), .B1(P1_DATAO_REG_18__SCAN_IN), 
        .B2(n11378), .ZN(n10775) );
  AOI22_X1 U13096 ( .A1(P2_DATAO_REG_19__SCAN_IN), .A2(n7142), .B1(
        P1_DATAO_REG_19__SCAN_IN), .B2(n11475), .ZN(n10774) );
  XNOR2_X1 U13097 ( .A(n10775), .B(n10774), .ZN(n12166) );
  INV_X1 U13098 ( .A(n12166), .ZN(n10580) );
  OAI222_X1 U13099 ( .A1(P3_U3151), .A2(n12345), .B1(n13335), .B2(n12163), 
        .C1(n13333), .C2(n10580), .ZN(P3_U3276) );
  INV_X1 U13100 ( .A(n10581), .ZN(n10583) );
  NAND2_X1 U13101 ( .A1(n13443), .A2(n12605), .ZN(n10629) );
  XNOR2_X1 U13102 ( .A(n10709), .B(n12611), .ZN(n10628) );
  XOR2_X1 U13103 ( .A(n10629), .B(n10628), .Z(n10630) );
  XOR2_X1 U13104 ( .A(n10631), .B(n10630), .Z(n10591) );
  AND2_X1 U13105 ( .A1(P2_U3088), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n13451) );
  AOI21_X1 U13106 ( .B1(n13374), .B2(n10586), .A(n13451), .ZN(n10589) );
  INV_X1 U13107 ( .A(n10587), .ZN(n10681) );
  OR2_X1 U13108 ( .A1(n13372), .A2(n10681), .ZN(n10588) );
  OAI211_X1 U13109 ( .C1(n13415), .C2(n10682), .A(n10589), .B(n10588), .ZN(
        n10590) );
  AOI21_X1 U13110 ( .B1(n10591), .B2(n13391), .A(n10590), .ZN(n10592) );
  INV_X1 U13111 ( .A(n10592), .ZN(P2_U3185) );
  AND2_X1 U13112 ( .A1(n10594), .A2(n10593), .ZN(n10597) );
  INV_X1 U13113 ( .A(n10595), .ZN(n10596) );
  INV_X1 U13114 ( .A(n10618), .ZN(n10598) );
  NAND2_X1 U13115 ( .A1(n14313), .A2(n10598), .ZN(n14165) );
  MUX2_X1 U13116 ( .A(n10600), .B(n10599), .S(n14313), .Z(n10607) );
  INV_X1 U13117 ( .A(n12553), .ZN(n10602) );
  OAI22_X1 U13118 ( .A1(n14243), .A2(n10603), .B1(P1_REG3_REG_3__SCAN_IN), 
        .B2(n14307), .ZN(n10604) );
  AOI21_X1 U13119 ( .B1(n14346), .B2(n10605), .A(n10604), .ZN(n10606) );
  OAI211_X1 U13120 ( .C1(n10608), .C2(n14165), .A(n10607), .B(n10606), .ZN(
        P1_U3290) );
  OAI21_X1 U13121 ( .B1(n10611), .B2(n10610), .A(n10609), .ZN(n10612) );
  AOI222_X1 U13122 ( .A1(n14324), .A2(n10612), .B1(n14042), .B2(n14321), .C1(
        n14045), .C2(n14319), .ZN(n14833) );
  INV_X1 U13123 ( .A(n14833), .ZN(n10617) );
  NOR2_X1 U13124 ( .A1(n14313), .A2(n9797), .ZN(n10616) );
  OAI211_X1 U13125 ( .C1(n10614), .C2(n6691), .A(n14427), .B(n10613), .ZN(
        n14832) );
  INV_X1 U13126 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n14066) );
  OAI22_X1 U13127 ( .A1(n14243), .A2(n14832), .B1(n14066), .B2(n14307), .ZN(
        n10615) );
  AOI211_X1 U13128 ( .C1(n10617), .C2(n14313), .A(n10616), .B(n10615), .ZN(
        n10625) );
  AND2_X1 U13129 ( .A1(n14155), .A2(n10618), .ZN(n10619) );
  OAI21_X1 U13130 ( .B1(n10622), .B2(n10620), .A(n10621), .ZN(n14836) );
  AOI22_X1 U13131 ( .A1(n14277), .A2(n14836), .B1(n14346), .B2(n10623), .ZN(
        n10624) );
  NAND2_X1 U13132 ( .A1(n10625), .A2(n10624), .ZN(P1_U3291) );
  NAND2_X1 U13133 ( .A1(P1_U4016), .A2(n14147), .ZN(n10626) );
  OAI21_X1 U13134 ( .B1(P1_U4016), .B2(n9094), .A(n10626), .ZN(P1_U3586) );
  INV_X1 U13135 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n14477) );
  NAND2_X1 U13136 ( .A1(n12615), .A2(n6492), .ZN(n10627) );
  OAI21_X1 U13137 ( .B1(n14477), .B2(n6492), .A(n10627), .ZN(P2_U3560) );
  XNOR2_X1 U13138 ( .A(n15068), .B(n9992), .ZN(n10633) );
  NAND2_X1 U13139 ( .A1(n13442), .A2(n12610), .ZN(n10632) );
  NAND2_X1 U13140 ( .A1(n10633), .A2(n10632), .ZN(n10905) );
  OAI21_X1 U13141 ( .B1(n10633), .B2(n10632), .A(n10905), .ZN(n10634) );
  AOI21_X1 U13142 ( .B1(n10635), .B2(n10634), .A(n10907), .ZN(n10641) );
  NAND2_X1 U13143 ( .A1(n13524), .A2(n13441), .ZN(n10637) );
  NAND2_X1 U13144 ( .A1(n13420), .A2(n13443), .ZN(n10636) );
  AND2_X1 U13145 ( .A1(n10637), .A2(n10636), .ZN(n10714) );
  NAND2_X1 U13146 ( .A1(n13422), .A2(n10721), .ZN(n10638) );
  NAND2_X1 U13147 ( .A1(P2_U3088), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n13464) );
  OAI211_X1 U13148 ( .C1(n13424), .C2(n10714), .A(n10638), .B(n13464), .ZN(
        n10639) );
  AOI21_X1 U13149 ( .B1(n15068), .B2(n13426), .A(n10639), .ZN(n10640) );
  OAI21_X1 U13150 ( .B1(n10641), .B2(n13428), .A(n10640), .ZN(P2_U3193) );
  OAI21_X1 U13151 ( .B1(n10643), .B2(n10645), .A(n10642), .ZN(n10939) );
  INV_X1 U13152 ( .A(n11142), .ZN(n10644) );
  AOI211_X1 U13153 ( .C1(n14002), .C2(n10658), .A(n14326), .B(n10644), .ZN(
        n10945) );
  XNOR2_X1 U13154 ( .A(n10646), .B(n10645), .ZN(n10650) );
  NAND2_X1 U13155 ( .A1(n14040), .A2(n14319), .ZN(n10648) );
  NAND2_X1 U13156 ( .A1(n14038), .A2(n14321), .ZN(n10647) );
  NAND2_X1 U13157 ( .A1(n10648), .A2(n10647), .ZN(n13998) );
  INV_X1 U13158 ( .A(n13998), .ZN(n10649) );
  OAI21_X1 U13159 ( .B1(n10650), .B2(n14282), .A(n10649), .ZN(n10940) );
  AOI211_X1 U13160 ( .C1(n14848), .C2(n10939), .A(n10945), .B(n10940), .ZN(
        n10654) );
  INV_X1 U13161 ( .A(n14002), .ZN(n10943) );
  OAI22_X1 U13162 ( .A1(n14468), .A2(n10943), .B1(n14849), .B2(n7626), .ZN(
        n10651) );
  INV_X1 U13163 ( .A(n10651), .ZN(n10652) );
  OAI21_X1 U13164 ( .B1(n10654), .B2(n6786), .A(n10652), .ZN(P1_U3477) );
  AOI22_X1 U13165 ( .A1(n14375), .A2(n14002), .B1(n14854), .B2(
        P1_REG1_REG_6__SCAN_IN), .ZN(n10653) );
  OAI21_X1 U13166 ( .B1(n10654), .B2(n14854), .A(n10653), .ZN(P1_U3534) );
  OAI21_X1 U13167 ( .B1(n10657), .B2(n10656), .A(n10655), .ZN(n10846) );
  OAI211_X1 U13168 ( .C1(n10832), .C2(n10668), .A(n14427), .B(n10658), .ZN(
        n10842) );
  INV_X1 U13169 ( .A(n10842), .ZN(n10667) );
  INV_X1 U13170 ( .A(n10846), .ZN(n10666) );
  OAI21_X1 U13171 ( .B1(n10661), .B2(n10660), .A(n10659), .ZN(n10664) );
  OAI22_X1 U13172 ( .A1(n10900), .A2(n14285), .B1(n10662), .B2(n14287), .ZN(
        n10663) );
  AOI21_X1 U13173 ( .B1(n10664), .B2(n14324), .A(n10663), .ZN(n10665) );
  OAI21_X1 U13174 ( .B1(n10666), .B2(n14155), .A(n10665), .ZN(n10843) );
  AOI211_X1 U13175 ( .C1(n14381), .C2(n10846), .A(n10667), .B(n10843), .ZN(
        n10672) );
  OAI22_X1 U13176 ( .A1(n14468), .A2(n10668), .B1(n14849), .B2(n7612), .ZN(
        n10669) );
  INV_X1 U13177 ( .A(n10669), .ZN(n10670) );
  OAI21_X1 U13178 ( .B1(n10672), .B2(n6786), .A(n10670), .ZN(P1_U3474) );
  AOI22_X1 U13179 ( .A1(n14375), .A2(n10897), .B1(n14854), .B2(
        P1_REG1_REG_5__SCAN_IN), .ZN(n10671) );
  OAI21_X1 U13180 ( .B1(n10672), .B2(n14854), .A(n10671), .ZN(P1_U3533) );
  NAND2_X1 U13181 ( .A1(n15012), .A2(n10673), .ZN(n10674) );
  NOR2_X1 U13182 ( .A1(n10675), .A2(n10674), .ZN(n10676) );
  NAND2_X1 U13183 ( .A1(n10677), .A2(n10676), .ZN(n10678) );
  NAND2_X1 U13184 ( .A1(n10347), .A2(n14988), .ZN(n10679) );
  OAI22_X1 U13185 ( .A1(n14968), .A2(n10682), .B1(n14996), .B2(n10681), .ZN(
        n10683) );
  AOI21_X1 U13186 ( .B1(n10684), .B2(n14722), .A(n10683), .ZN(n10688) );
  MUX2_X1 U13187 ( .A(n10686), .B(n10685), .S(n15002), .Z(n10687) );
  OAI211_X1 U13188 ( .C1(n10689), .C2(n13739), .A(n10688), .B(n10687), .ZN(
        P2_U3258) );
  OAI211_X1 U13189 ( .C1(n10692), .C2(n10691), .A(n10690), .B(n13995), .ZN(
        n10696) );
  AOI22_X1 U13190 ( .A1(n13987), .A2(n14040), .B1(n14011), .B2(n14042), .ZN(
        n10693) );
  NAND2_X1 U13191 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_U3086), .ZN(n14799) );
  OAI211_X1 U13192 ( .C1(n14839), .C2(n13980), .A(n10693), .B(n14799), .ZN(
        n10694) );
  INV_X1 U13193 ( .A(n10694), .ZN(n10695) );
  OAI211_X1 U13194 ( .C1(n13989), .C2(n10835), .A(n10696), .B(n10695), .ZN(
        P1_U3230) );
  XNOR2_X1 U13195 ( .A(n10697), .B(n10702), .ZN(n15043) );
  OR2_X1 U13196 ( .A1(n15042), .A2(n10768), .ZN(n10698) );
  AND3_X1 U13197 ( .A1(n10698), .A2(n14980), .A3(n10086), .ZN(n15038) );
  MUX2_X1 U13198 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n15039), .S(n15002), .Z(
        n10700) );
  OAI22_X1 U13199 ( .A1(n14968), .A2(n15042), .B1(P2_REG3_REG_3__SCAN_IN), 
        .B2(n14996), .ZN(n10699) );
  AOI211_X1 U13200 ( .C1(n15038), .C2(n14722), .A(n10700), .B(n10699), .ZN(
        n10704) );
  NAND2_X1 U13201 ( .A1(n15002), .A2(n15064), .ZN(n13755) );
  INV_X1 U13202 ( .A(n13755), .ZN(n13737) );
  XNOR2_X1 U13203 ( .A(n10702), .B(n10701), .ZN(n15046) );
  NAND2_X1 U13204 ( .A1(n13737), .A2(n15046), .ZN(n10703) );
  OAI211_X1 U13205 ( .C1(n15043), .C2(n13739), .A(n10704), .B(n10703), .ZN(
        P2_U3262) );
  XNOR2_X1 U13206 ( .A(n10732), .B(n10728), .ZN(n10718) );
  INV_X1 U13207 ( .A(n10718), .ZN(n15072) );
  INV_X1 U13208 ( .A(n14988), .ZN(n10707) );
  NAND2_X1 U13209 ( .A1(n15002), .A2(n10707), .ZN(n14984) );
  INV_X1 U13210 ( .A(n10347), .ZN(n10717) );
  AND2_X1 U13211 ( .A1(n10709), .A2(n10708), .ZN(n10710) );
  INV_X1 U13212 ( .A(n10727), .ZN(n10712) );
  AOI21_X1 U13213 ( .B1(n10728), .B2(n10713), .A(n10712), .ZN(n10715) );
  OAI21_X1 U13214 ( .B1(n10715), .B2(n14997), .A(n10714), .ZN(n10716) );
  AOI21_X1 U13215 ( .B1(n10718), .B2(n10717), .A(n10716), .ZN(n15071) );
  MUX2_X1 U13216 ( .A(n10719), .B(n15071), .S(n15002), .Z(n10725) );
  AOI211_X1 U13217 ( .C1(n15068), .C2(n10720), .A(n12610), .B(n6948), .ZN(
        n15067) );
  INV_X1 U13218 ( .A(n15068), .ZN(n10730) );
  INV_X1 U13219 ( .A(n10721), .ZN(n10722) );
  OAI22_X1 U13220 ( .A1(n10730), .A2(n14968), .B1(n14996), .B2(n10722), .ZN(
        n10723) );
  AOI21_X1 U13221 ( .B1(n15067), .B2(n14722), .A(n10723), .ZN(n10724) );
  OAI211_X1 U13222 ( .C1(n15072), .C2(n14984), .A(n10725), .B(n10724), .ZN(
        P2_U3257) );
  NAND2_X1 U13223 ( .A1(n10727), .A2(n10726), .ZN(n10869) );
  INV_X1 U13224 ( .A(n10733), .ZN(n10866) );
  XNOR2_X1 U13225 ( .A(n10869), .B(n10866), .ZN(n10758) );
  INV_X1 U13226 ( .A(n10728), .ZN(n10731) );
  XNOR2_X1 U13227 ( .A(n10867), .B(n10733), .ZN(n10754) );
  NAND2_X1 U13228 ( .A1(n10754), .A2(n14723), .ZN(n10742) );
  AOI21_X1 U13229 ( .B1(n10918), .B2(n10734), .A(n12605), .ZN(n10735) );
  AND2_X1 U13230 ( .A1(n10735), .A2(n10877), .ZN(n10755) );
  NAND2_X1 U13231 ( .A1(n13524), .A2(n13440), .ZN(n10737) );
  NAND2_X1 U13232 ( .A1(n13420), .A2(n13442), .ZN(n10736) );
  NAND2_X1 U13233 ( .A1(n10737), .A2(n10736), .ZN(n10913) );
  AOI22_X1 U13234 ( .A1(n15002), .A2(n10913), .B1(n10912), .B2(n14979), .ZN(
        n10739) );
  NAND2_X1 U13235 ( .A1(n15005), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n10738) );
  OAI211_X1 U13236 ( .C1(n6947), .C2(n14968), .A(n10739), .B(n10738), .ZN(
        n10740) );
  AOI21_X1 U13237 ( .B1(n14722), .B2(n10755), .A(n10740), .ZN(n10741) );
  OAI211_X1 U13238 ( .C1(n10758), .C2(n13755), .A(n10742), .B(n10741), .ZN(
        P2_U3256) );
  XNOR2_X1 U13239 ( .A(n10743), .B(n10751), .ZN(n15060) );
  AOI211_X1 U13240 ( .C1(n15058), .C2(n14981), .A(n12605), .B(n10744), .ZN(
        n15056) );
  AOI22_X1 U13241 ( .A1(n15002), .A2(n15057), .B1(n10745), .B2(n14979), .ZN(
        n10747) );
  OR2_X1 U13242 ( .A1(n15002), .A2(n9700), .ZN(n10746) );
  OAI211_X1 U13243 ( .C1(n14968), .C2(n10748), .A(n10747), .B(n10746), .ZN(
        n10749) );
  AOI21_X1 U13244 ( .B1(n15056), .B2(n14722), .A(n10749), .ZN(n10753) );
  XNOR2_X1 U13245 ( .A(n10750), .B(n10751), .ZN(n15063) );
  NAND2_X1 U13246 ( .A1(n15063), .A2(n13737), .ZN(n10752) );
  OAI211_X1 U13247 ( .C1(n15060), .C2(n13739), .A(n10753), .B(n10752), .ZN(
        P2_U3260) );
  NAND2_X1 U13248 ( .A1(n10754), .A2(n15035), .ZN(n10757) );
  AOI211_X1 U13249 ( .C1(n15069), .C2(n10918), .A(n10913), .B(n10755), .ZN(
        n10756) );
  OAI211_X1 U13250 ( .C1(n14997), .C2(n10758), .A(n10757), .B(n10756), .ZN(
        n10760) );
  NAND2_X1 U13251 ( .A1(n10760), .A2(n15096), .ZN(n10759) );
  OAI21_X1 U13252 ( .B1(n15096), .B2(n9864), .A(n10759), .ZN(P2_U3508) );
  INV_X1 U13253 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n10762) );
  NAND2_X1 U13254 ( .A1(n10760), .A2(n15066), .ZN(n10761) );
  OAI21_X1 U13255 ( .B1(n15066), .B2(n10762), .A(n10761), .ZN(P2_U3457) );
  XNOR2_X1 U13256 ( .A(n10343), .B(n10763), .ZN(n10765) );
  AOI21_X1 U13257 ( .B1(n10765), .B2(n15064), .A(n10764), .ZN(n15032) );
  XNOR2_X1 U13258 ( .A(n10767), .B(n10766), .ZN(n15036) );
  AOI22_X1 U13259 ( .A1(n15005), .A2(P2_REG2_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(n14979), .ZN(n10771) );
  AOI211_X1 U13260 ( .C1(n10769), .C2(n10983), .A(n12605), .B(n10768), .ZN(
        n15030) );
  NAND2_X1 U13261 ( .A1(n14722), .A2(n15030), .ZN(n10770) );
  OAI211_X1 U13262 ( .C1(n6747), .C2(n14968), .A(n10771), .B(n10770), .ZN(
        n10772) );
  AOI21_X1 U13263 ( .B1(n14723), .B2(n15036), .A(n10772), .ZN(n10773) );
  OAI21_X1 U13264 ( .B1(n15005), .B2(n15032), .A(n10773), .ZN(P2_U3263) );
  NAND2_X1 U13265 ( .A1(n10775), .A2(n10774), .ZN(n10776) );
  AOI22_X1 U13266 ( .A1(P2_DATAO_REG_20__SCAN_IN), .A2(n7139), .B1(
        P1_DATAO_REG_20__SCAN_IN), .B2(n7985), .ZN(n10962) );
  XNOR2_X1 U13267 ( .A(n10961), .B(n10962), .ZN(n12175) );
  INV_X1 U13268 ( .A(n12175), .ZN(n10778) );
  OAI222_X1 U13269 ( .A1(n10779), .A2(P3_U3151), .B1(n13333), .B2(n10778), 
        .C1(n10777), .C2(n13335), .ZN(P3_U3275) );
  INV_X1 U13270 ( .A(n10780), .ZN(n10782) );
  INV_X1 U13271 ( .A(n11186), .ZN(n14810) );
  OAI222_X1 U13272 ( .A1(n14478), .A2(n10781), .B1(n14480), .B2(n10782), .C1(
        P1_U3086), .C2(n14810), .ZN(P1_U3340) );
  INV_X1 U13273 ( .A(n14923), .ZN(n13501) );
  OAI222_X1 U13274 ( .A1(n13870), .A2(n10783), .B1(n13873), .B2(n10782), .C1(
        P2_U3088), .C2(n13501), .ZN(P2_U3312) );
  INV_X1 U13275 ( .A(P3_REG3_REG_24__SCAN_IN), .ZN(n12221) );
  INV_X1 U13276 ( .A(n12253), .ZN(n10785) );
  INV_X1 U13277 ( .A(P3_REG3_REG_26__SCAN_IN), .ZN(n10784) );
  NAND2_X1 U13278 ( .A1(n10785), .A2(n10784), .ZN(n12266) );
  INV_X1 U13279 ( .A(n12285), .ZN(n10787) );
  INV_X1 U13280 ( .A(P3_REG3_REG_28__SCAN_IN), .ZN(n10786) );
  NAND2_X1 U13281 ( .A1(n10787), .A2(n10786), .ZN(n12827) );
  INV_X1 U13282 ( .A(P3_REG0_REG_29__SCAN_IN), .ZN(n13206) );
  NAND2_X1 U13283 ( .A1(n12268), .A2(P3_REG2_REG_29__SCAN_IN), .ZN(n10790) );
  NAND2_X1 U13284 ( .A1(n6495), .A2(P3_REG1_REG_29__SCAN_IN), .ZN(n10789) );
  OAI211_X1 U13285 ( .C1(n10791), .C2(n13206), .A(n10790), .B(n10789), .ZN(
        n10792) );
  INV_X1 U13286 ( .A(n10792), .ZN(n10793) );
  NAND2_X1 U13287 ( .A1(n12743), .A2(P3_DATAO_REG_29__SCAN_IN), .ZN(n10794) );
  OAI21_X1 U13288 ( .B1(n12881), .B2(n12743), .A(n10794), .ZN(P3_U3520) );
  INV_X1 U13289 ( .A(n10795), .ZN(n11048) );
  NAND2_X1 U13290 ( .A1(n12282), .A2(n10796), .ZN(n10800) );
  NAND2_X1 U13291 ( .A1(n10449), .A2(n10797), .ZN(n10799) );
  OR2_X1 U13292 ( .A1(n11392), .A2(n15122), .ZN(n10798) );
  XNOR2_X1 U13293 ( .A(n6486), .B(n11021), .ZN(n10927) );
  XNOR2_X1 U13294 ( .A(n10927), .B(n12753), .ZN(n10806) );
  INV_X1 U13295 ( .A(n10801), .ZN(n10802) );
  NAND2_X1 U13296 ( .A1(n10802), .A2(n12754), .ZN(n10803) );
  OAI21_X1 U13297 ( .B1(n10806), .B2(n10805), .A(n11113), .ZN(n10807) );
  NAND2_X1 U13298 ( .A1(n10807), .A2(n12709), .ZN(n10816) );
  NAND2_X1 U13299 ( .A1(n12268), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n10812) );
  NAND2_X1 U13300 ( .A1(n6491), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n10811) );
  OAI21_X1 U13301 ( .B1(P3_REG3_REG_4__SCAN_IN), .B2(P3_REG3_REG_3__SCAN_IN), 
        .A(P3_REG3_REG_5__SCAN_IN), .ZN(n10808) );
  NAND2_X1 U13302 ( .A1(n10929), .A2(n10808), .ZN(n11035) );
  NAND2_X1 U13303 ( .A1(n10235), .A2(n11035), .ZN(n10810) );
  NAND2_X1 U13304 ( .A1(n10454), .A2(P3_REG0_REG_5__SCAN_IN), .ZN(n10809) );
  NAND2_X1 U13305 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(P3_U3151), .ZN(n15123) );
  INV_X1 U13306 ( .A(n15123), .ZN(n10814) );
  INV_X1 U13307 ( .A(n11021), .ZN(n15229) );
  OAI22_X1 U13308 ( .A1(n12717), .A2(n15229), .B1(n15172), .B2(n12736), .ZN(
        n10813) );
  AOI211_X1 U13309 ( .C1(n12733), .C2(n12752), .A(n10814), .B(n10813), .ZN(
        n10815) );
  OAI211_X1 U13310 ( .C1(n11048), .C2(n11596), .A(n10816), .B(n10815), .ZN(
        P3_U3170) );
  NOR2_X1 U13311 ( .A1(n14243), .A2(n14326), .ZN(n14344) );
  OAI21_X1 U13312 ( .B1(n14344), .B2(n14346), .A(n9548), .ZN(n10821) );
  INV_X1 U13313 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n10817) );
  OAI22_X1 U13314 ( .A1(n14830), .A2(n10818), .B1(n10817), .B2(n14307), .ZN(
        n10819) );
  AOI21_X1 U13315 ( .B1(P1_REG2_REG_0__SCAN_IN), .B2(n14830), .A(n10819), .ZN(
        n10820) );
  OAI211_X1 U13316 ( .C1(n14334), .C2(n10822), .A(n10821), .B(n10820), .ZN(
        P1_U3293) );
  OAI21_X1 U13317 ( .B1(n10825), .B2(n10824), .A(n10823), .ZN(n14841) );
  INV_X1 U13318 ( .A(n14841), .ZN(n10840) );
  OAI21_X1 U13319 ( .B1(n10828), .B2(n10827), .A(n10826), .ZN(n10829) );
  AOI222_X1 U13320 ( .A1(n14324), .A2(n10829), .B1(n14040), .B2(n14321), .C1(
        n14042), .C2(n14319), .ZN(n14838) );
  MUX2_X1 U13321 ( .A(n10830), .B(n14838), .S(n14313), .Z(n10839) );
  INV_X1 U13322 ( .A(n10831), .ZN(n10834) );
  INV_X1 U13323 ( .A(n10832), .ZN(n10833) );
  OAI211_X1 U13324 ( .C1(n14839), .C2(n10834), .A(n10833), .B(n14427), .ZN(
        n14837) );
  OAI22_X1 U13325 ( .A1(n14243), .A2(n14837), .B1(n10835), .B2(n14307), .ZN(
        n10836) );
  AOI21_X1 U13326 ( .B1(n14346), .B2(n10837), .A(n10836), .ZN(n10838) );
  OAI211_X1 U13327 ( .C1(n10840), .C2(n14334), .A(n10839), .B(n10838), .ZN(
        P1_U3289) );
  INV_X1 U13328 ( .A(n14165), .ZN(n14826) );
  INV_X1 U13329 ( .A(n14307), .ZN(n14819) );
  AOI22_X1 U13330 ( .A1(n14346), .A2(n10897), .B1(n14819), .B2(n10902), .ZN(
        n10841) );
  OAI21_X1 U13331 ( .B1(n14243), .B2(n10842), .A(n10841), .ZN(n10845) );
  MUX2_X1 U13332 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n10843), .S(n14313), .Z(
        n10844) );
  AOI211_X1 U13333 ( .C1(n14826), .C2(n10846), .A(n10845), .B(n10844), .ZN(
        n10847) );
  INV_X1 U13334 ( .A(n10847), .ZN(P1_U3288) );
  AOI21_X1 U13335 ( .B1(n11326), .B2(n10849), .A(n10848), .ZN(n10865) );
  AOI21_X1 U13336 ( .B1(n8423), .B2(n10851), .A(n10850), .ZN(n10852) );
  NOR2_X1 U13337 ( .A1(n10852), .A2(n15136), .ZN(n10863) );
  INV_X1 U13338 ( .A(n10853), .ZN(n11453) );
  NAND3_X1 U13339 ( .A1(n10856), .A2(n10855), .A3(n10854), .ZN(n10857) );
  AOI21_X1 U13340 ( .B1(n11453), .B2(n10857), .A(n15131), .ZN(n10862) );
  INV_X1 U13341 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n11501) );
  NOR2_X1 U13342 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11501), .ZN(n10858) );
  AOI21_X1 U13343 ( .B1(n15097), .B2(P3_ADDR_REG_9__SCAN_IN), .A(n10858), .ZN(
        n10859) );
  OAI21_X1 U13344 ( .B1(n15139), .B2(n10860), .A(n10859), .ZN(n10861) );
  NOR3_X1 U13345 ( .A1(n10863), .A2(n10862), .A3(n10861), .ZN(n10864) );
  OAI21_X1 U13346 ( .B1(n10865), .B2(n15163), .A(n10864), .ZN(P3_U3191) );
  INV_X1 U13347 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n10880) );
  XNOR2_X1 U13348 ( .A(n10949), .B(n10953), .ZN(n10969) );
  INV_X1 U13349 ( .A(n13441), .ZN(n10868) );
  NAND2_X1 U13350 ( .A1(n10869), .A2(n10868), .ZN(n10870) );
  XNOR2_X1 U13351 ( .A(n10954), .B(n10953), .ZN(n10875) );
  NAND2_X1 U13352 ( .A1(n13524), .A2(n13439), .ZN(n10873) );
  NAND2_X1 U13353 ( .A1(n13420), .A2(n13441), .ZN(n10872) );
  AND2_X1 U13354 ( .A1(n10873), .A2(n10872), .ZN(n11057) );
  INV_X1 U13355 ( .A(n11057), .ZN(n10874) );
  AOI21_X1 U13356 ( .B1(n10875), .B2(n15064), .A(n10874), .ZN(n10974) );
  INV_X1 U13357 ( .A(n10950), .ZN(n10876) );
  AOI211_X1 U13358 ( .C1(n11059), .C2(n10877), .A(n12610), .B(n10876), .ZN(
        n10972) );
  AOI21_X1 U13359 ( .B1(n15069), .B2(n11059), .A(n10972), .ZN(n10878) );
  OAI211_X1 U13360 ( .C1(n10969), .C2(n15061), .A(n10974), .B(n10878), .ZN(
        n10891) );
  NAND2_X1 U13361 ( .A1(n10891), .A2(n15066), .ZN(n10879) );
  OAI21_X1 U13362 ( .B1(n15066), .B2(n10880), .A(n10879), .ZN(P2_U3460) );
  INV_X1 U13363 ( .A(n10881), .ZN(n10882) );
  OAI22_X1 U13364 ( .A1(n14968), .A2(n10883), .B1(n14996), .B2(n10882), .ZN(
        n10884) );
  AOI21_X1 U13365 ( .B1(n10885), .B2(n14722), .A(n10884), .ZN(n10889) );
  MUX2_X1 U13366 ( .A(n10887), .B(n10886), .S(n15002), .Z(n10888) );
  OAI211_X1 U13367 ( .C1(n10890), .C2(n13739), .A(n10889), .B(n10888), .ZN(
        P2_U3259) );
  NAND2_X1 U13368 ( .A1(n10891), .A2(n15096), .ZN(n10892) );
  OAI21_X1 U13369 ( .B1(n15096), .B2(n10893), .A(n10892), .ZN(P2_U3509) );
  XNOR2_X1 U13370 ( .A(n10895), .B(n7106), .ZN(n10896) );
  XNOR2_X1 U13371 ( .A(n10894), .B(n10896), .ZN(n10904) );
  AOI22_X1 U13372 ( .A1(n13987), .A2(n14039), .B1(n10897), .B2(n14018), .ZN(
        n10899) );
  OAI211_X1 U13373 ( .C1(n10900), .C2(n13985), .A(n10899), .B(n10898), .ZN(
        n10901) );
  AOI21_X1 U13374 ( .B1(n10902), .B2(n14016), .A(n10901), .ZN(n10903) );
  OAI21_X1 U13375 ( .B1(n10904), .B2(n14022), .A(n10903), .ZN(P1_U3227) );
  INV_X1 U13376 ( .A(n10905), .ZN(n10906) );
  XNOR2_X1 U13377 ( .A(n10918), .B(n9992), .ZN(n10909) );
  NAND2_X1 U13378 ( .A1(n13441), .A2(n12610), .ZN(n10908) );
  NAND2_X1 U13379 ( .A1(n10909), .A2(n10908), .ZN(n11052) );
  OAI21_X1 U13380 ( .B1(n10909), .B2(n10908), .A(n11052), .ZN(n10910) );
  AOI21_X1 U13381 ( .B1(n10911), .B2(n10910), .A(n11053), .ZN(n10920) );
  INV_X1 U13382 ( .A(n10912), .ZN(n10916) );
  NAND2_X1 U13383 ( .A1(n13374), .A2(n10913), .ZN(n10915) );
  OAI211_X1 U13384 ( .C1(n13372), .C2(n10916), .A(n10915), .B(n10914), .ZN(
        n10917) );
  AOI21_X1 U13385 ( .B1(n10918), .B2(n13426), .A(n10917), .ZN(n10919) );
  OAI21_X1 U13386 ( .B1(n10920), .B2(n13428), .A(n10919), .ZN(P2_U3203) );
  NAND2_X1 U13387 ( .A1(n12282), .A2(n10921), .ZN(n10926) );
  NAND2_X1 U13388 ( .A1(n10449), .A2(n10922), .ZN(n10925) );
  OR2_X1 U13389 ( .A1(n11392), .A2(n10923), .ZN(n10924) );
  XNOR2_X1 U13390 ( .A(n6486), .B(n11020), .ZN(n11107) );
  XNOR2_X1 U13391 ( .A(n11107), .B(n12752), .ZN(n11110) );
  NAND2_X1 U13392 ( .A1(n10927), .A2(n11031), .ZN(n11108) );
  NAND2_X1 U13393 ( .A1(n11113), .A2(n11108), .ZN(n10928) );
  XOR2_X1 U13394 ( .A(n11110), .B(n10928), .Z(n10938) );
  NAND2_X1 U13395 ( .A1(n12268), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n10934) );
  NAND2_X1 U13396 ( .A1(n6491), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n10933) );
  NAND2_X1 U13397 ( .A1(n10929), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n10930) );
  NAND2_X1 U13398 ( .A1(n11075), .A2(n10930), .ZN(n11136) );
  NAND2_X1 U13399 ( .A1(n10235), .A2(n11136), .ZN(n10932) );
  NAND2_X1 U13400 ( .A1(n10454), .A2(P3_REG0_REG_6__SCAN_IN), .ZN(n10931) );
  AOI22_X1 U13401 ( .A1(n12720), .A2(n12753), .B1(n12739), .B2(n11020), .ZN(
        n10935) );
  NAND2_X1 U13402 ( .A1(P3_REG3_REG_5__SCAN_IN), .A2(P3_U3151), .ZN(n15143) );
  OAI211_X1 U13403 ( .C1(n11266), .C2(n12723), .A(n10935), .B(n15143), .ZN(
        n10936) );
  AOI21_X1 U13404 ( .B1(n11035), .B2(n12732), .A(n10936), .ZN(n10937) );
  OAI21_X1 U13405 ( .B1(n10938), .B2(n12741), .A(n10937), .ZN(P3_U3167) );
  INV_X1 U13406 ( .A(n10939), .ZN(n10948) );
  INV_X1 U13407 ( .A(n10940), .ZN(n10941) );
  MUX2_X1 U13408 ( .A(n10942), .B(n10941), .S(n14313), .Z(n10947) );
  OAI22_X1 U13409 ( .A1(n14823), .A2(n10943), .B1(n14000), .B2(n14307), .ZN(
        n10944) );
  AOI21_X1 U13410 ( .B1(n10945), .B2(n14817), .A(n10944), .ZN(n10946) );
  OAI211_X1 U13411 ( .C1(n10948), .C2(n14334), .A(n10947), .B(n10946), .ZN(
        P1_U3287) );
  INV_X1 U13412 ( .A(n11059), .ZN(n10968) );
  XOR2_X1 U13413 ( .A(n11245), .B(n11251), .Z(n15075) );
  AOI211_X1 U13414 ( .C1(n11276), .C2(n10950), .A(n12605), .B(n14720), .ZN(
        n15081) );
  INV_X1 U13415 ( .A(n11276), .ZN(n15078) );
  AOI22_X1 U13416 ( .A1(n15005), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n11285), 
        .B2(n14979), .ZN(n10951) );
  OAI21_X1 U13417 ( .B1(n15078), .B2(n14968), .A(n10951), .ZN(n10952) );
  AOI21_X1 U13418 ( .B1(n15081), .B2(n14722), .A(n10952), .ZN(n10960) );
  NAND2_X1 U13419 ( .A1(n10954), .A2(n10953), .ZN(n10957) );
  NAND2_X1 U13420 ( .A1(n11059), .A2(n10955), .ZN(n10956) );
  XOR2_X1 U13421 ( .A(n11246), .B(n11245), .Z(n10958) );
  AOI22_X1 U13422 ( .A1(n13420), .A2(n13440), .B1(n13524), .B2(n13438), .ZN(
        n11283) );
  OAI21_X1 U13423 ( .B1(n10958), .B2(n14997), .A(n11283), .ZN(n15079) );
  NAND2_X1 U13424 ( .A1(n15079), .A2(n15002), .ZN(n10959) );
  OAI211_X1 U13425 ( .C1(n15075), .C2(n13739), .A(n10960), .B(n10959), .ZN(
        P2_U3254) );
  INV_X1 U13426 ( .A(SI_21_), .ZN(n10966) );
  INV_X1 U13427 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n11615) );
  AOI22_X1 U13428 ( .A1(P2_DATAO_REG_21__SCAN_IN), .A2(
        P1_DATAO_REG_21__SCAN_IN), .B1(n11619), .B2(n11615), .ZN(n10963) );
  INV_X1 U13429 ( .A(n10963), .ZN(n10964) );
  XNOR2_X1 U13430 ( .A(n11062), .B(n10964), .ZN(n12190) );
  INV_X1 U13431 ( .A(n12190), .ZN(n10965) );
  OAI222_X1 U13432 ( .A1(P3_U3151), .A2(n12367), .B1(n13335), .B2(n10966), 
        .C1(n13333), .C2(n10965), .ZN(P3_U3274) );
  AOI22_X1 U13433 ( .A1(n15005), .A2(P2_REG2_REG_10__SCAN_IN), .B1(n11054), 
        .B2(n14979), .ZN(n10967) );
  OAI21_X1 U13434 ( .B1(n10968), .B2(n14968), .A(n10967), .ZN(n10971) );
  NOR2_X1 U13435 ( .A1(n10969), .A2(n13739), .ZN(n10970) );
  AOI211_X1 U13436 ( .C1(n10972), .C2(n14722), .A(n10971), .B(n10970), .ZN(
        n10973) );
  OAI21_X1 U13437 ( .B1(n15005), .B2(n10974), .A(n10973), .ZN(P2_U3255) );
  INV_X1 U13438 ( .A(n10975), .ZN(n10977) );
  OAI222_X1 U13439 ( .A1(n14478), .A2(n10976), .B1(n14480), .B2(n10977), .C1(
        n11289), .C2(P1_U3086), .ZN(P1_U3339) );
  INV_X1 U13440 ( .A(n14935), .ZN(n13504) );
  OAI222_X1 U13441 ( .A1(P2_U3088), .A2(n13504), .B1(n13870), .B2(n7884), .C1(
        n10977), .C2(n13873), .ZN(P2_U3311) );
  XNOR2_X1 U13442 ( .A(n10349), .B(n10978), .ZN(n10980) );
  AOI21_X1 U13443 ( .B1(n10980), .B2(n15064), .A(n10979), .ZN(n15025) );
  XNOR2_X1 U13444 ( .A(n10349), .B(n10981), .ZN(n15022) );
  NAND2_X1 U13445 ( .A1(n10987), .A2(n14990), .ZN(n10982) );
  NAND3_X1 U13446 ( .A1(n10983), .A2(n10086), .A3(n10982), .ZN(n15024) );
  INV_X1 U13447 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n10984) );
  OAI22_X1 U13448 ( .A1(n15002), .A2(n10985), .B1(n10984), .B2(n14996), .ZN(
        n10986) );
  AOI21_X1 U13449 ( .B1(n14715), .B2(n10987), .A(n10986), .ZN(n10988) );
  OAI21_X1 U13450 ( .B1(n14983), .B2(n15024), .A(n10988), .ZN(n10989) );
  AOI21_X1 U13451 ( .B1(n15022), .B2(n14723), .A(n10989), .ZN(n10990) );
  OAI21_X1 U13452 ( .B1(n15005), .B2(n15025), .A(n10990), .ZN(P2_U3264) );
  NAND2_X1 U13453 ( .A1(n10991), .A2(n12374), .ZN(n15171) );
  NAND2_X1 U13454 ( .A1(n12378), .A2(n12365), .ZN(n15174) );
  INV_X1 U13455 ( .A(n15174), .ZN(n15177) );
  NAND2_X1 U13456 ( .A1(n15172), .A2(n15223), .ZN(n12383) );
  NAND2_X1 U13457 ( .A1(n12754), .A2(n10994), .ZN(n12384) );
  AND2_X2 U13458 ( .A1(n12383), .A2(n12384), .ZN(n12512) );
  OR2_X1 U13459 ( .A1(n10995), .A2(n12512), .ZN(n10996) );
  NAND2_X1 U13460 ( .A1(n11018), .A2(n10996), .ZN(n15225) );
  INV_X1 U13461 ( .A(n15225), .ZN(n11017) );
  INV_X1 U13462 ( .A(n15206), .ZN(n10997) );
  OR2_X1 U13463 ( .A1(n10997), .A2(n12367), .ZN(n15186) );
  AND2_X1 U13464 ( .A1(n15261), .A2(n12505), .ZN(n10998) );
  NAND2_X1 U13465 ( .A1(n13291), .A2(n10998), .ZN(n11000) );
  NAND2_X1 U13466 ( .A1(n15225), .A2(n15204), .ZN(n11012) );
  INV_X1 U13467 ( .A(n12545), .ZN(n11002) );
  OAI22_X1 U13468 ( .A1(n15198), .A2(n15173), .B1(n11031), .B2(n15197), .ZN(
        n11003) );
  INV_X1 U13469 ( .A(n11003), .ZN(n11011) );
  NAND2_X1 U13470 ( .A1(n15198), .A2(n15184), .ZN(n11005) );
  AND2_X1 U13471 ( .A1(n15176), .A2(n11005), .ZN(n11004) );
  NAND2_X1 U13472 ( .A1(n15193), .A2(n11004), .ZN(n11008) );
  INV_X1 U13473 ( .A(n11005), .ZN(n11006) );
  OR2_X1 U13474 ( .A1(n11006), .A2(n15174), .ZN(n11007) );
  OR2_X1 U13475 ( .A1(n11027), .A2(n12512), .ZN(n11043) );
  NAND2_X1 U13476 ( .A1(n11027), .A2(n12512), .ZN(n11009) );
  NAND3_X1 U13477 ( .A1(n11043), .A2(n15200), .A3(n11009), .ZN(n11010) );
  AND3_X1 U13478 ( .A1(n11012), .A2(n11011), .A3(n11010), .ZN(n15227) );
  MUX2_X1 U13479 ( .A(n11013), .B(n15227), .S(n15211), .Z(n11016) );
  INV_X1 U13480 ( .A(n13047), .ZN(n12831) );
  AOI22_X1 U13481 ( .A1(n12831), .A2(n15223), .B1(n15208), .B2(n11014), .ZN(
        n11015) );
  OAI211_X1 U13482 ( .C1(n11017), .C2(n11224), .A(n11016), .B(n11015), .ZN(
        P3_U3230) );
  NAND2_X1 U13483 ( .A1(n11031), .A2(n11021), .ZN(n12387) );
  NAND2_X1 U13484 ( .A1(n12753), .A2(n15229), .ZN(n12388) );
  NAND2_X1 U13485 ( .A1(n12387), .A2(n12388), .ZN(n11040) );
  INV_X1 U13486 ( .A(n11040), .ZN(n12510) );
  NAND2_X1 U13487 ( .A1(n11041), .A2(n12510), .ZN(n11019) );
  NAND2_X1 U13488 ( .A1(n11128), .A2(n11020), .ZN(n12394) );
  INV_X1 U13489 ( .A(n11020), .ZN(n15234) );
  NAND2_X1 U13490 ( .A1(n12752), .A2(n15234), .ZN(n12392) );
  XOR2_X1 U13491 ( .A(n11088), .B(n12509), .Z(n15235) );
  NAND2_X1 U13492 ( .A1(n12753), .A2(n11021), .ZN(n11023) );
  INV_X1 U13493 ( .A(n11023), .ZN(n11022) );
  NOR2_X1 U13494 ( .A1(n11022), .A2(n11040), .ZN(n11025) );
  OR2_X1 U13495 ( .A1(n12512), .A2(n11025), .ZN(n11028) );
  NAND2_X1 U13496 ( .A1(n12754), .A2(n15223), .ZN(n11042) );
  AND2_X1 U13497 ( .A1(n11042), .A2(n11023), .ZN(n11024) );
  OR2_X1 U13498 ( .A1(n11025), .A2(n11024), .ZN(n11026) );
  INV_X1 U13499 ( .A(n11029), .ZN(n11030) );
  OAI21_X1 U13500 ( .B1(n11030), .B2(n7337), .A(n11070), .ZN(n11033) );
  OAI22_X1 U13501 ( .A1(n11031), .A2(n15173), .B1(n11266), .B2(n15197), .ZN(
        n11032) );
  AOI21_X1 U13502 ( .B1(n11033), .B2(n15200), .A(n11032), .ZN(n11034) );
  OAI21_X1 U13503 ( .B1(n15235), .B2(n13054), .A(n11034), .ZN(n15237) );
  NAND2_X1 U13504 ( .A1(n15237), .A2(n15211), .ZN(n11039) );
  INV_X1 U13505 ( .A(n11035), .ZN(n11036) );
  OAI22_X1 U13506 ( .A1(n13047), .A2(n15234), .B1(n11036), .B2(n11954), .ZN(
        n11037) );
  AOI21_X1 U13507 ( .B1(n15213), .B2(P3_REG2_REG_5__SCAN_IN), .A(n11037), .ZN(
        n11038) );
  OAI211_X1 U13508 ( .C1(n15235), .C2(n11224), .A(n11039), .B(n11038), .ZN(
        P3_U3228) );
  XNOR2_X1 U13509 ( .A(n11041), .B(n11040), .ZN(n15230) );
  NAND2_X1 U13510 ( .A1(n11043), .A2(n11042), .ZN(n11044) );
  XNOR2_X1 U13511 ( .A(n11044), .B(n12510), .ZN(n11046) );
  OAI22_X1 U13512 ( .A1(n11128), .A2(n15197), .B1(n15172), .B2(n15173), .ZN(
        n11045) );
  AOI21_X1 U13513 ( .B1(n11046), .B2(n15200), .A(n11045), .ZN(n11047) );
  OAI21_X1 U13514 ( .B1(n13054), .B2(n15230), .A(n11047), .ZN(n15232) );
  NAND2_X1 U13515 ( .A1(n15232), .A2(n15211), .ZN(n11051) );
  OAI22_X1 U13516 ( .A1(n13047), .A2(n15229), .B1(n11048), .B2(n11954), .ZN(
        n11049) );
  AOI21_X1 U13517 ( .B1(n15213), .B2(P3_REG2_REG_4__SCAN_IN), .A(n11049), .ZN(
        n11050) );
  OAI211_X1 U13518 ( .C1(n15230), .C2(n11224), .A(n11051), .B(n11050), .ZN(
        P3_U3229) );
  XNOR2_X1 U13519 ( .A(n11059), .B(n12611), .ZN(n11273) );
  NAND2_X1 U13520 ( .A1(n13440), .A2(n12610), .ZN(n11272) );
  XNOR2_X1 U13521 ( .A(n11273), .B(n11272), .ZN(n11275) );
  XNOR2_X1 U13522 ( .A(n6646), .B(n11275), .ZN(n11061) );
  NAND2_X1 U13523 ( .A1(n13422), .A2(n11054), .ZN(n11055) );
  OAI211_X1 U13524 ( .C1(n13424), .C2(n11057), .A(n11056), .B(n11055), .ZN(
        n11058) );
  AOI21_X1 U13525 ( .B1(n11059), .B2(n13426), .A(n11058), .ZN(n11060) );
  OAI21_X1 U13526 ( .B1(n11061), .B2(n13428), .A(n11060), .ZN(P2_U3189) );
  NAND2_X1 U13527 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(n11615), .ZN(n11063) );
  INV_X1 U13528 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n11064) );
  AOI22_X1 U13529 ( .A1(P2_DATAO_REG_22__SCAN_IN), .A2(n11813), .B1(
        P1_DATAO_REG_22__SCAN_IN), .B2(n11064), .ZN(n11225) );
  INV_X1 U13530 ( .A(n11225), .ZN(n11065) );
  XNOR2_X1 U13531 ( .A(n11226), .B(n11065), .ZN(n12203) );
  NOR2_X1 U13532 ( .A1(n13335), .A2(SI_22_), .ZN(n11066) );
  AOI21_X1 U13533 ( .B1(n13053), .B2(P3_STATE_REG_SCAN_IN), .A(n11066), .ZN(
        n11067) );
  OAI21_X1 U13534 ( .B1(n12203), .B2(n13333), .A(n11067), .ZN(n11068) );
  INV_X1 U13535 ( .A(n11068), .ZN(P3_U3273) );
  NAND2_X1 U13536 ( .A1(n11128), .A2(n15234), .ZN(n11069) );
  NAND2_X1 U13537 ( .A1(n10449), .A2(n11071), .ZN(n11073) );
  NAND2_X1 U13538 ( .A1(n12282), .A2(SI_6_), .ZN(n11072) );
  OAI211_X1 U13539 ( .C1(n11392), .C2(n11074), .A(n11073), .B(n11072), .ZN(
        n11137) );
  NAND2_X1 U13540 ( .A1(n11266), .A2(n11137), .ZN(n12396) );
  INV_X1 U13541 ( .A(n11137), .ZN(n15239) );
  NAND2_X1 U13542 ( .A1(n12751), .A2(n15239), .ZN(n12398) );
  NAND2_X1 U13543 ( .A1(n12751), .A2(n11137), .ZN(n11211) );
  NAND2_X1 U13544 ( .A1(n11215), .A2(n11211), .ZN(n11087) );
  NAND2_X1 U13545 ( .A1(n12268), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n11081) );
  NAND2_X1 U13546 ( .A1(n6491), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n11080) );
  INV_X1 U13547 ( .A(n11093), .ZN(n11077) );
  NAND2_X1 U13548 ( .A1(n11075), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n11076) );
  NAND2_X1 U13549 ( .A1(n11077), .A2(n11076), .ZN(n11261) );
  NAND2_X1 U13550 ( .A1(n10235), .A2(n11261), .ZN(n11079) );
  NAND2_X1 U13551 ( .A1(n10454), .A2(P3_REG0_REG_7__SCAN_IN), .ZN(n11078) );
  NAND2_X1 U13552 ( .A1(n12311), .A2(n11082), .ZN(n11086) );
  NAND2_X1 U13553 ( .A1(n12282), .A2(n11083), .ZN(n11085) );
  OR2_X1 U13554 ( .A1(n11392), .A2(n15154), .ZN(n11084) );
  NAND2_X1 U13555 ( .A1(n11371), .A2(n11210), .ZN(n12402) );
  NAND2_X1 U13556 ( .A1(n12750), .A2(n15244), .ZN(n12403) );
  NAND2_X1 U13557 ( .A1(n12402), .A2(n12403), .ZN(n12405) );
  XNOR2_X1 U13558 ( .A(n11087), .B(n12405), .ZN(n11102) );
  NAND2_X1 U13559 ( .A1(n11088), .A2(n12509), .ZN(n11089) );
  NAND2_X1 U13560 ( .A1(n11089), .A2(n12394), .ZN(n11125) );
  NAND2_X1 U13561 ( .A1(n11125), .A2(n12513), .ZN(n11127) );
  INV_X1 U13562 ( .A(n12405), .ZN(n12514) );
  NAND3_X1 U13563 ( .A1(n11127), .A2(n12405), .A3(n12396), .ZN(n11091) );
  NAND2_X1 U13564 ( .A1(n11204), .A2(n11091), .ZN(n15247) );
  NAND2_X1 U13565 ( .A1(n12268), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n11099) );
  NAND2_X1 U13566 ( .A1(n6491), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n11098) );
  OR2_X1 U13567 ( .A1(n11093), .A2(n11092), .ZN(n11094) );
  NAND2_X1 U13568 ( .A1(n11095), .A2(n11094), .ZN(n11220) );
  NAND2_X1 U13569 ( .A1(n10235), .A2(n11220), .ZN(n11097) );
  NAND2_X1 U13570 ( .A1(n10454), .A2(P3_REG0_REG_8__SCAN_IN), .ZN(n11096) );
  OAI22_X1 U13571 ( .A1(n11266), .A2(n15173), .B1(n11502), .B2(n15197), .ZN(
        n11100) );
  AOI21_X1 U13572 ( .B1(n15247), .B2(n15204), .A(n11100), .ZN(n11101) );
  OAI21_X1 U13573 ( .B1(n11102), .B2(n15178), .A(n11101), .ZN(n15245) );
  INV_X1 U13574 ( .A(n15245), .ZN(n11106) );
  AOI22_X1 U13575 ( .A1(n12831), .A2(n11210), .B1(n15208), .B2(n11261), .ZN(
        n11103) );
  OAI21_X1 U13576 ( .B1(n8402), .B2(n15211), .A(n11103), .ZN(n11104) );
  AOI21_X1 U13577 ( .B1(n15247), .B2(n15209), .A(n11104), .ZN(n11105) );
  OAI21_X1 U13578 ( .B1(n11106), .B2(n15213), .A(n11105), .ZN(P3_U3226) );
  INV_X1 U13579 ( .A(n11136), .ZN(n11121) );
  NAND2_X1 U13580 ( .A1(n11107), .A2(n11128), .ZN(n11109) );
  AND2_X1 U13581 ( .A1(n11108), .A2(n11109), .ZN(n11112) );
  INV_X1 U13582 ( .A(n11109), .ZN(n11111) );
  XNOR2_X1 U13583 ( .A(n12151), .B(n15239), .ZN(n11262) );
  XNOR2_X1 U13584 ( .A(n11262), .B(n12751), .ZN(n11114) );
  AOI21_X1 U13585 ( .B1(n11115), .B2(n11114), .A(n12741), .ZN(n11116) );
  NAND2_X1 U13586 ( .A1(n11116), .A2(n11264), .ZN(n11120) );
  OAI22_X1 U13587 ( .A1(n12717), .A2(n15239), .B1(n11128), .B2(n12736), .ZN(
        n11117) );
  AOI211_X1 U13588 ( .C1(n12733), .C2(n12750), .A(n11118), .B(n11117), .ZN(
        n11119) );
  OAI211_X1 U13589 ( .C1(n11121), .C2(n11596), .A(n11120), .B(n11119), .ZN(
        P3_U3179) );
  INV_X1 U13590 ( .A(n11122), .ZN(n11124) );
  INV_X1 U13591 ( .A(n11296), .ZN(n11578) );
  OAI222_X1 U13592 ( .A1(n14478), .A2(n11123), .B1(n14480), .B2(n11124), .C1(
        n11578), .C2(P1_U3086), .ZN(P1_U3338) );
  INV_X1 U13593 ( .A(n14943), .ZN(n13506) );
  OAI222_X1 U13594 ( .A1(n13870), .A2(n13208), .B1(n13873), .B2(n11124), .C1(
        n13506), .C2(P2_U3088), .ZN(P2_U3310) );
  OR2_X1 U13595 ( .A1(n11125), .A2(n12513), .ZN(n11126) );
  NAND2_X1 U13596 ( .A1(n11127), .A2(n11126), .ZN(n11130) );
  INV_X1 U13597 ( .A(n11130), .ZN(n15240) );
  OAI22_X1 U13598 ( .A1(n11128), .A2(n15173), .B1(n11371), .B2(n15197), .ZN(
        n11129) );
  AOI21_X1 U13599 ( .B1(n11130), .B2(n15204), .A(n11129), .ZN(n11134) );
  NAND2_X1 U13600 ( .A1(n11131), .A2(n12513), .ZN(n11132) );
  NAND3_X1 U13601 ( .A1(n11215), .A2(n15200), .A3(n11132), .ZN(n11133) );
  NAND2_X1 U13602 ( .A1(n11134), .A2(n11133), .ZN(n15241) );
  MUX2_X1 U13603 ( .A(n15241), .B(P3_REG2_REG_6__SCAN_IN), .S(n15213), .Z(
        n11135) );
  INV_X1 U13604 ( .A(n11135), .ZN(n11139) );
  AOI22_X1 U13605 ( .A1(n12831), .A2(n11137), .B1(n15208), .B2(n11136), .ZN(
        n11138) );
  OAI211_X1 U13606 ( .C1(n15240), .C2(n11224), .A(n11139), .B(n11138), .ZN(
        P3_U3227) );
  OAI21_X1 U13607 ( .B1(n11141), .B2(n11148), .A(n11140), .ZN(n14827) );
  NAND2_X1 U13608 ( .A1(n11142), .A2(n11200), .ZN(n11143) );
  NAND2_X1 U13609 ( .A1(n11143), .A2(n14427), .ZN(n11144) );
  NOR2_X1 U13610 ( .A1(n11235), .A2(n11144), .ZN(n14818) );
  INV_X1 U13611 ( .A(n14155), .ZN(n14209) );
  NAND2_X1 U13612 ( .A1(n14039), .A2(n14319), .ZN(n11146) );
  NAND2_X1 U13613 ( .A1(n14037), .A2(n14321), .ZN(n11145) );
  NAND2_X1 U13614 ( .A1(n11146), .A2(n11145), .ZN(n11196) );
  XNOR2_X1 U13615 ( .A(n11147), .B(n11148), .ZN(n11149) );
  NOR2_X1 U13616 ( .A1(n11149), .A2(n14282), .ZN(n11150) );
  AOI211_X1 U13617 ( .C1(n14209), .C2(n14827), .A(n11196), .B(n11150), .ZN(
        n14829) );
  INV_X1 U13618 ( .A(n14829), .ZN(n11151) );
  AOI211_X1 U13619 ( .C1(n14381), .C2(n14827), .A(n14818), .B(n11151), .ZN(
        n11155) );
  AOI22_X1 U13620 ( .A1(n14375), .A2(n11200), .B1(n14854), .B2(
        P1_REG1_REG_7__SCAN_IN), .ZN(n11152) );
  OAI21_X1 U13621 ( .B1(n11155), .B2(n14854), .A(n11152), .ZN(P1_U3535) );
  INV_X1 U13622 ( .A(n11200), .ZN(n14824) );
  OAI22_X1 U13623 ( .A1(n14468), .A2(n14824), .B1(n14849), .B2(n7657), .ZN(
        n11153) );
  INV_X1 U13624 ( .A(n11153), .ZN(n11154) );
  OAI21_X1 U13625 ( .B1(n11155), .B2(n6786), .A(n11154), .ZN(P1_U3480) );
  OAI21_X1 U13626 ( .B1(n11157), .B2(n11161), .A(n11156), .ZN(n11343) );
  INV_X1 U13627 ( .A(n11343), .ZN(n11171) );
  INV_X1 U13628 ( .A(n11159), .ZN(n11160) );
  AOI21_X1 U13629 ( .B1(n11161), .B2(n11158), .A(n11160), .ZN(n11164) );
  AOI22_X1 U13630 ( .A1(n14319), .A2(n14037), .B1(n14035), .B2(n14321), .ZN(
        n11163) );
  NAND2_X1 U13631 ( .A1(n11343), .A2(n14209), .ZN(n11162) );
  OAI211_X1 U13632 ( .C1(n11164), .C2(n14282), .A(n11163), .B(n11162), .ZN(
        n11341) );
  NAND2_X1 U13633 ( .A1(n11341), .A2(n14313), .ZN(n11170) );
  XNOR2_X1 U13634 ( .A(n11233), .B(n11345), .ZN(n11165) );
  NOR2_X1 U13635 ( .A1(n11165), .A2(n14326), .ZN(n11342) );
  INV_X1 U13636 ( .A(n11166), .ZN(n11757) );
  AOI22_X1 U13637 ( .A1(n14830), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n11757), 
        .B2(n14819), .ZN(n11167) );
  OAI21_X1 U13638 ( .B1(n14823), .B2(n11345), .A(n11167), .ZN(n11168) );
  AOI21_X1 U13639 ( .B1(n11342), .B2(n14817), .A(n11168), .ZN(n11169) );
  OAI211_X1 U13640 ( .C1(n11171), .C2(n14165), .A(n11170), .B(n11169), .ZN(
        P1_U3284) );
  NAND2_X1 U13641 ( .A1(n11172), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n11174) );
  NAND2_X1 U13642 ( .A1(n11174), .A2(n11173), .ZN(n11175) );
  NOR2_X1 U13643 ( .A1(n11186), .A2(n11175), .ZN(n11176) );
  XNOR2_X1 U13644 ( .A(n11186), .B(n11175), .ZN(n14805) );
  NOR2_X1 U13645 ( .A1(P1_REG2_REG_15__SCAN_IN), .A2(n14805), .ZN(n14804) );
  NOR2_X1 U13646 ( .A1(n11176), .A2(n14804), .ZN(n11181) );
  INV_X1 U13647 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n11178) );
  NAND2_X1 U13648 ( .A1(n11295), .A2(n11178), .ZN(n11177) );
  OAI21_X1 U13649 ( .B1(n11295), .B2(n11178), .A(n11177), .ZN(n11180) );
  NAND2_X1 U13650 ( .A1(n11289), .A2(n11178), .ZN(n11179) );
  OAI211_X1 U13651 ( .C1(n11289), .C2(n11178), .A(n11181), .B(n11179), .ZN(
        n11288) );
  OAI211_X1 U13652 ( .C1(n11181), .C2(n11180), .A(n11288), .B(n14113), .ZN(
        n11192) );
  NAND2_X1 U13653 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n13935)
         );
  XNOR2_X1 U13654 ( .A(n11289), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n11294) );
  AOI21_X1 U13655 ( .B1(n11184), .B2(n11183), .A(n11182), .ZN(n11185) );
  NOR2_X1 U13656 ( .A1(n11186), .A2(n11185), .ZN(n11187) );
  XNOR2_X1 U13657 ( .A(n11186), .B(n11185), .ZN(n14803) );
  NOR2_X1 U13658 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(n14803), .ZN(n14802) );
  NOR2_X1 U13659 ( .A1(n11187), .A2(n14802), .ZN(n11293) );
  XOR2_X1 U13660 ( .A(n11294), .B(n11293), .Z(n11188) );
  NAND2_X1 U13661 ( .A1(n14102), .A2(n11188), .ZN(n11189) );
  NAND2_X1 U13662 ( .A1(n13935), .A2(n11189), .ZN(n11190) );
  AOI21_X1 U13663 ( .B1(n14088), .B2(P1_ADDR_REG_16__SCAN_IN), .A(n11190), 
        .ZN(n11191) );
  OAI211_X1 U13664 ( .C1(n14811), .C2(n11289), .A(n11192), .B(n11191), .ZN(
        P1_U3259) );
  XNOR2_X1 U13665 ( .A(n11194), .B(n11193), .ZN(n11203) );
  INV_X1 U13666 ( .A(n11195), .ZN(n14820) );
  NAND2_X1 U13667 ( .A1(n13999), .A2(n11196), .ZN(n11198) );
  NAND2_X1 U13668 ( .A1(n11198), .A2(n11197), .ZN(n11199) );
  AOI21_X1 U13669 ( .B1(n14820), .B2(n14016), .A(n11199), .ZN(n11202) );
  NAND2_X1 U13670 ( .A1(n14018), .A2(n11200), .ZN(n11201) );
  OAI211_X1 U13671 ( .C1(n11203), .C2(n14022), .A(n11202), .B(n11201), .ZN(
        P1_U3213) );
  NAND2_X1 U13672 ( .A1(n12311), .A2(n11205), .ZN(n11209) );
  NAND2_X1 U13673 ( .A1(n12282), .A2(SI_8_), .ZN(n11208) );
  OR2_X1 U13674 ( .A1(n11392), .A2(n11206), .ZN(n11207) );
  NAND2_X1 U13675 ( .A1(n11502), .A2(n15249), .ZN(n11310) );
  INV_X1 U13676 ( .A(n15249), .ZN(n11315) );
  NAND2_X1 U13677 ( .A1(n12749), .A2(n11315), .ZN(n11312) );
  NAND2_X1 U13678 ( .A1(n11310), .A2(n11312), .ZN(n12518) );
  XNOR2_X1 U13679 ( .A(n11314), .B(n12518), .ZN(n11217) );
  INV_X1 U13680 ( .A(n11217), .ZN(n15250) );
  NAND2_X1 U13681 ( .A1(n12750), .A2(n11210), .ZN(n11212) );
  AND2_X1 U13682 ( .A1(n11211), .A2(n11212), .ZN(n11214) );
  INV_X1 U13683 ( .A(n11212), .ZN(n11213) );
  XOR2_X1 U13684 ( .A(n11311), .B(n12518), .Z(n11219) );
  OAI22_X1 U13685 ( .A1(n12412), .A2(n15197), .B1(n11371), .B2(n15173), .ZN(
        n11216) );
  AOI21_X1 U13686 ( .B1(n11217), .B2(n15204), .A(n11216), .ZN(n11218) );
  OAI21_X1 U13687 ( .B1(n11219), .B2(n15178), .A(n11218), .ZN(n15252) );
  NAND2_X1 U13688 ( .A1(n15252), .A2(n15211), .ZN(n11223) );
  INV_X1 U13689 ( .A(n11220), .ZN(n11376) );
  OAI22_X1 U13690 ( .A1(n13047), .A2(n15249), .B1(n11376), .B2(n11954), .ZN(
        n11221) );
  AOI21_X1 U13691 ( .B1(P3_REG2_REG_8__SCAN_IN), .B2(n15213), .A(n11221), .ZN(
        n11222) );
  OAI211_X1 U13692 ( .C1(n15250), .C2(n11224), .A(n11223), .B(n11222), .ZN(
        P3_U3225) );
  INV_X1 U13693 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n11887) );
  AOI22_X1 U13694 ( .A1(P2_DATAO_REG_23__SCAN_IN), .A2(
        P1_DATAO_REG_23__SCAN_IN), .B1(n11892), .B2(n11887), .ZN(n11740) );
  NAND2_X1 U13695 ( .A1(n11226), .A2(n11225), .ZN(n11227) );
  XNOR2_X1 U13696 ( .A(n11740), .B(n11739), .ZN(n12230) );
  NAND2_X1 U13697 ( .A1(n12230), .A2(n13320), .ZN(n11228) );
  OAI211_X1 U13698 ( .C1(n11229), .C2(n13335), .A(n11228), .B(n12549), .ZN(
        P3_U3272) );
  OAI21_X1 U13699 ( .B1(n11232), .B2(n11231), .A(n11230), .ZN(n14847) );
  INV_X1 U13700 ( .A(n11233), .ZN(n11234) );
  OAI211_X1 U13701 ( .C1(n14844), .C2(n11235), .A(n11234), .B(n14427), .ZN(
        n14842) );
  NOR2_X1 U13702 ( .A1(n14307), .A2(n11469), .ZN(n11236) );
  AOI21_X1 U13703 ( .B1(n14346), .B2(n11471), .A(n11236), .ZN(n11237) );
  OAI21_X1 U13704 ( .B1(n14842), .B2(n14243), .A(n11237), .ZN(n11243) );
  XNOR2_X1 U13705 ( .A(n11238), .B(n11239), .ZN(n11240) );
  OAI222_X1 U13706 ( .A1(n14287), .A2(n11465), .B1(n14285), .B2(n11241), .C1(
        n11240), .C2(n14282), .ZN(n14845) );
  MUX2_X1 U13707 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n14845), .S(n14313), .Z(
        n11242) );
  AOI211_X1 U13708 ( .C1(n14277), .C2(n14847), .A(n11243), .B(n11242), .ZN(
        n11244) );
  INV_X1 U13709 ( .A(n11244), .ZN(P1_U3285) );
  INV_X1 U13710 ( .A(n13439), .ZN(n11249) );
  NAND2_X1 U13711 ( .A1(n11276), .A2(n11249), .ZN(n11247) );
  XOR2_X1 U13712 ( .A(n11555), .B(n11253), .Z(n14740) );
  INV_X1 U13713 ( .A(n14716), .ZN(n14750) );
  NOR2_X1 U13714 ( .A1(n15078), .A2(n11249), .ZN(n11250) );
  XNOR2_X1 U13715 ( .A(n11547), .B(n11253), .ZN(n14746) );
  NAND2_X1 U13716 ( .A1(n14750), .A2(n14720), .ZN(n14719) );
  NAND2_X1 U13717 ( .A1(n11638), .A2(n14719), .ZN(n11254) );
  NAND3_X1 U13718 ( .A1(n14706), .A2(n10086), .A3(n11254), .ZN(n14742) );
  AOI22_X1 U13719 ( .A1(n13420), .A2(n13438), .B1(n13524), .B2(n13436), .ZN(
        n14741) );
  INV_X1 U13720 ( .A(n11627), .ZN(n11255) );
  OAI22_X1 U13721 ( .A1(n15005), .A2(n14741), .B1(n11255), .B2(n14996), .ZN(
        n11257) );
  INV_X1 U13722 ( .A(n11638), .ZN(n14743) );
  NOR2_X1 U13723 ( .A1(n14743), .A2(n14968), .ZN(n11256) );
  AOI211_X1 U13724 ( .C1(n15005), .C2(P2_REG2_REG_13__SCAN_IN), .A(n11257), 
        .B(n11256), .ZN(n11258) );
  OAI21_X1 U13725 ( .B1(n14983), .B2(n14742), .A(n11258), .ZN(n11259) );
  AOI21_X1 U13726 ( .B1(n14746), .B2(n14723), .A(n11259), .ZN(n11260) );
  OAI21_X1 U13727 ( .B1(n13755), .B2(n14740), .A(n11260), .ZN(P2_U3252) );
  INV_X1 U13728 ( .A(n11261), .ZN(n11271) );
  NAND2_X1 U13729 ( .A1(n11262), .A2(n12751), .ZN(n11263) );
  NAND2_X1 U13730 ( .A1(n11264), .A2(n11263), .ZN(n11265) );
  XNOR2_X1 U13731 ( .A(n12405), .B(n12292), .ZN(n11365) );
  OAI211_X1 U13732 ( .C1(n11265), .C2(n11365), .A(n11368), .B(n12709), .ZN(
        n11270) );
  NAND2_X1 U13733 ( .A1(P3_REG3_REG_7__SCAN_IN), .A2(P3_U3151), .ZN(n15166) );
  INV_X1 U13734 ( .A(n15166), .ZN(n11268) );
  OAI22_X1 U13735 ( .A1(n12717), .A2(n15244), .B1(n11266), .B2(n12736), .ZN(
        n11267) );
  AOI211_X1 U13736 ( .C1(n12733), .C2(n12749), .A(n11268), .B(n11267), .ZN(
        n11269) );
  OAI211_X1 U13737 ( .C1(n11271), .C2(n11596), .A(n11270), .B(n11269), .ZN(
        P3_U3153) );
  INV_X1 U13738 ( .A(n11272), .ZN(n11274) );
  AND2_X1 U13739 ( .A1(n13439), .A2(n12605), .ZN(n11278) );
  XNOR2_X1 U13740 ( .A(n11276), .B(n12611), .ZN(n11277) );
  NOR2_X1 U13741 ( .A1(n11277), .A2(n11278), .ZN(n11330) );
  AOI21_X1 U13742 ( .B1(n11278), .B2(n11277), .A(n11330), .ZN(n11279) );
  OAI21_X1 U13743 ( .B1(n11280), .B2(n11279), .A(n11332), .ZN(n11281) );
  NAND2_X1 U13744 ( .A1(n11281), .A2(n13391), .ZN(n11287) );
  OAI21_X1 U13745 ( .B1(n13424), .B2(n11283), .A(n11282), .ZN(n11284) );
  AOI21_X1 U13746 ( .B1(n11285), .B2(n13422), .A(n11284), .ZN(n11286) );
  OAI211_X1 U13747 ( .C1(n15078), .C2(n13415), .A(n11287), .B(n11286), .ZN(
        P2_U3208) );
  OAI21_X1 U13748 ( .B1(n11289), .B2(n11178), .A(n11288), .ZN(n11292) );
  NAND2_X1 U13749 ( .A1(n11296), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n11575) );
  INV_X1 U13750 ( .A(n11575), .ZN(n11290) );
  AOI21_X1 U13751 ( .B1(n7895), .B2(n11578), .A(n11290), .ZN(n11291) );
  NAND2_X1 U13752 ( .A1(n11291), .A2(n11292), .ZN(n11574) );
  OAI211_X1 U13753 ( .C1(n11292), .C2(n11291), .A(n14113), .B(n11574), .ZN(
        n11303) );
  NAND2_X1 U13754 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n13944)
         );
  AOI22_X1 U13755 ( .A1(P1_REG1_REG_16__SCAN_IN), .A2(n11295), .B1(n11294), 
        .B2(n11293), .ZN(n11298) );
  XNOR2_X1 U13756 ( .A(n11296), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n11297) );
  OR2_X1 U13757 ( .A1(n11298), .A2(n11297), .ZN(n11577) );
  NAND2_X1 U13758 ( .A1(n11298), .A2(n11297), .ZN(n11299) );
  NAND3_X1 U13759 ( .A1(n14102), .A2(n11577), .A3(n11299), .ZN(n11300) );
  NAND2_X1 U13760 ( .A1(n13944), .A2(n11300), .ZN(n11301) );
  AOI21_X1 U13761 ( .B1(n14088), .B2(P1_ADDR_REG_17__SCAN_IN), .A(n11301), 
        .ZN(n11302) );
  OAI211_X1 U13762 ( .C1(n14811), .C2(n11578), .A(n11303), .B(n11302), .ZN(
        P1_U3260) );
  NAND2_X1 U13763 ( .A1(n11304), .A2(n12311), .ZN(n11309) );
  NAND2_X1 U13764 ( .A1(n12282), .A2(n11305), .ZN(n11308) );
  OR2_X1 U13765 ( .A1(n11392), .A2(n11306), .ZN(n11307) );
  XNOR2_X1 U13766 ( .A(n12411), .B(n12413), .ZN(n12520) );
  NAND2_X1 U13767 ( .A1(n11311), .A2(n11310), .ZN(n11313) );
  NAND2_X1 U13768 ( .A1(n11313), .A2(n11312), .ZN(n11397) );
  XOR2_X1 U13769 ( .A(n6481), .B(n12520), .Z(n11324) );
  NAND2_X1 U13770 ( .A1(n12749), .A2(n15249), .ZN(n12408) );
  NAND2_X1 U13771 ( .A1(n11502), .A2(n11315), .ZN(n12407) );
  XNOR2_X1 U13772 ( .A(n11388), .B(n12520), .ZN(n15258) );
  NAND2_X1 U13773 ( .A1(n12155), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n11321) );
  NAND2_X1 U13774 ( .A1(n6491), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n11320) );
  AND2_X1 U13775 ( .A1(n11316), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n11317) );
  OR2_X1 U13776 ( .A1(n11317), .A2(n11399), .ZN(n11585) );
  NAND2_X1 U13777 ( .A1(n10235), .A2(n11585), .ZN(n11319) );
  NAND2_X1 U13778 ( .A1(n10454), .A2(P3_REG0_REG_10__SCAN_IN), .ZN(n11318) );
  OAI22_X1 U13779 ( .A1(n11502), .A2(n15173), .B1(n11542), .B2(n15197), .ZN(
        n11322) );
  AOI21_X1 U13780 ( .B1(n15258), .B2(n15204), .A(n11322), .ZN(n11323) );
  OAI21_X1 U13781 ( .B1(n11324), .B2(n15178), .A(n11323), .ZN(n15255) );
  INV_X1 U13782 ( .A(n15255), .ZN(n11329) );
  AOI22_X1 U13783 ( .A1(n12831), .A2(n12413), .B1(n15208), .B2(n11505), .ZN(
        n11325) );
  OAI21_X1 U13784 ( .B1(n11326), .B2(n15211), .A(n11325), .ZN(n11327) );
  AOI21_X1 U13785 ( .B1(n15258), .B2(n15209), .A(n11327), .ZN(n11328) );
  OAI21_X1 U13786 ( .B1(n11329), .B2(n15213), .A(n11328), .ZN(P3_U3224) );
  INV_X1 U13787 ( .A(n11330), .ZN(n11331) );
  XOR2_X1 U13788 ( .A(n12611), .B(n14716), .Z(n11632) );
  NAND2_X1 U13789 ( .A1(n13438), .A2(n12610), .ZN(n11631) );
  XNOR2_X1 U13790 ( .A(n11632), .B(n11631), .ZN(n11333) );
  XNOR2_X1 U13791 ( .A(n11633), .B(n11333), .ZN(n11340) );
  INV_X1 U13792 ( .A(n14714), .ZN(n11337) );
  NAND2_X1 U13793 ( .A1(n13524), .A2(n13437), .ZN(n11335) );
  NAND2_X1 U13794 ( .A1(n13420), .A2(n13439), .ZN(n11334) );
  NAND2_X1 U13795 ( .A1(n11335), .A2(n11334), .ZN(n14712) );
  AOI22_X1 U13796 ( .A1(n13374), .A2(n14712), .B1(P2_REG3_REG_12__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11336) );
  OAI21_X1 U13797 ( .B1(n11337), .B2(n13372), .A(n11336), .ZN(n11338) );
  AOI21_X1 U13798 ( .B1(n14716), .B2(n13426), .A(n11338), .ZN(n11339) );
  OAI21_X1 U13799 ( .B1(n11340), .B2(n13428), .A(n11339), .ZN(P2_U3196) );
  AOI211_X1 U13800 ( .C1(n14381), .C2(n11343), .A(n11342), .B(n11341), .ZN(
        n11349) );
  INV_X1 U13801 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n11344) );
  OAI22_X1 U13802 ( .A1(n11345), .A2(n14468), .B1(n14849), .B2(n11344), .ZN(
        n11346) );
  INV_X1 U13803 ( .A(n11346), .ZN(n11347) );
  OAI21_X1 U13804 ( .B1(n11349), .B2(n6786), .A(n11347), .ZN(P1_U3486) );
  AOI22_X1 U13805 ( .A1(n14375), .A2(n11767), .B1(n14854), .B2(
        P1_REG1_REG_9__SCAN_IN), .ZN(n11348) );
  OAI21_X1 U13806 ( .B1(n11349), .B2(n14854), .A(n11348), .ZN(P1_U3537) );
  AOI211_X1 U13807 ( .C1(n11663), .C2(n11351), .A(n14326), .B(n11350), .ZN(
        n11353) );
  OAI22_X1 U13808 ( .A1(n11352), .A2(n14287), .B1(n11465), .B2(n14285), .ZN(
        n11658) );
  OR2_X1 U13809 ( .A1(n11353), .A2(n11658), .ZN(n11382) );
  INV_X1 U13810 ( .A(n11354), .ZN(n11355) );
  AOI211_X1 U13811 ( .C1(n11360), .C2(n11356), .A(n14282), .B(n11355), .ZN(
        n11381) );
  AOI21_X1 U13812 ( .B1(n12108), .B2(n11382), .A(n11381), .ZN(n11364) );
  OAI22_X1 U13813 ( .A1(n14313), .A2(n11357), .B1(n11661), .B2(n14307), .ZN(
        n11358) );
  AOI21_X1 U13814 ( .B1(n11663), .B2(n14346), .A(n11358), .ZN(n11363) );
  OAI21_X1 U13815 ( .B1(n11361), .B2(n11360), .A(n11359), .ZN(n11383) );
  NAND2_X1 U13816 ( .A1(n11383), .A2(n14277), .ZN(n11362) );
  OAI211_X1 U13817 ( .C1(n11364), .C2(n14830), .A(n11363), .B(n11362), .ZN(
        P1_U3283) );
  INV_X1 U13818 ( .A(n11365), .ZN(n11366) );
  NAND2_X1 U13819 ( .A1(n11366), .A2(n12750), .ZN(n11367) );
  NAND2_X1 U13820 ( .A1(n11368), .A2(n11367), .ZN(n11370) );
  XNOR2_X1 U13821 ( .A(n12151), .B(n15249), .ZN(n11494) );
  XNOR2_X1 U13822 ( .A(n11494), .B(n11502), .ZN(n11369) );
  OAI211_X1 U13823 ( .C1(n11370), .C2(n11369), .A(n11496), .B(n12709), .ZN(
        n11375) );
  OAI22_X1 U13824 ( .A1(n12717), .A2(n15249), .B1(n11371), .B2(n12736), .ZN(
        n11372) );
  AOI211_X1 U13825 ( .C1(n12733), .C2(n12411), .A(n11373), .B(n11372), .ZN(
        n11374) );
  OAI211_X1 U13826 ( .C1(n11376), .C2(n11596), .A(n11375), .B(n11374), .ZN(
        P3_U3161) );
  INV_X1 U13827 ( .A(n11377), .ZN(n11379) );
  INV_X1 U13828 ( .A(n12100), .ZN(n11584) );
  OAI222_X1 U13829 ( .A1(n14478), .A2(n11378), .B1(n14480), .B2(n11379), .C1(
        P1_U3086), .C2(n11584), .ZN(P1_U3337) );
  INV_X1 U13830 ( .A(n14958), .ZN(n13507) );
  OAI222_X1 U13831 ( .A1(n13870), .A2(n11380), .B1(n13873), .B2(n11379), .C1(
        P2_U3088), .C2(n13507), .ZN(P2_U3309) );
  AOI211_X1 U13832 ( .C1(n14848), .C2(n11383), .A(n11382), .B(n11381), .ZN(
        n11387) );
  INV_X1 U13833 ( .A(n14468), .ZN(n11753) );
  NOR2_X1 U13834 ( .A1(n14849), .A2(n7737), .ZN(n11384) );
  AOI21_X1 U13835 ( .B1(n11663), .B2(n11753), .A(n11384), .ZN(n11385) );
  OAI21_X1 U13836 ( .B1(n11387), .B2(n6786), .A(n11385), .ZN(P1_U3489) );
  AOI22_X1 U13837 ( .A1(n11663), .A2(n14375), .B1(n14854), .B2(
        P1_REG1_REG_10__SCAN_IN), .ZN(n11386) );
  OAI21_X1 U13838 ( .B1(n11387), .B2(n14854), .A(n11386), .ZN(P1_U3538) );
  NAND2_X1 U13839 ( .A1(n11388), .A2(n12520), .ZN(n11390) );
  NAND2_X1 U13840 ( .A1(n12412), .A2(n12413), .ZN(n11389) );
  NAND2_X1 U13841 ( .A1(n11390), .A2(n11389), .ZN(n11526) );
  NAND2_X1 U13842 ( .A1(n11391), .A2(n12311), .ZN(n11396) );
  AOI22_X1 U13843 ( .A1(n12332), .A2(n11394), .B1(n12162), .B2(n11393), .ZN(
        n11395) );
  NAND2_X1 U13844 ( .A1(n11589), .A2(n11542), .ZN(n12418) );
  INV_X1 U13845 ( .A(n11589), .ZN(n15260) );
  NAND2_X1 U13846 ( .A1(n15260), .A2(n12748), .ZN(n12419) );
  NAND2_X1 U13847 ( .A1(n12418), .A2(n12419), .ZN(n11525) );
  XNOR2_X1 U13848 ( .A(n11526), .B(n11525), .ZN(n15263) );
  INV_X1 U13849 ( .A(n12413), .ZN(n15254) );
  OAI211_X1 U13850 ( .C1(n11398), .C2(n11525), .A(n11540), .B(n15200), .ZN(
        n11406) );
  NAND2_X1 U13851 ( .A1(n12268), .A2(P3_REG2_REG_11__SCAN_IN), .ZN(n11404) );
  NAND2_X1 U13852 ( .A1(n6491), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n11403) );
  NOR2_X1 U13853 ( .A1(n11399), .A2(n11431), .ZN(n11400) );
  OR2_X1 U13854 ( .A1(n11534), .A2(n11400), .ZN(n11792) );
  NAND2_X1 U13855 ( .A1(n10235), .A2(n11792), .ZN(n11402) );
  NAND2_X1 U13856 ( .A1(n10454), .A2(P3_REG0_REG_11__SCAN_IN), .ZN(n11401) );
  AOI22_X1 U13857 ( .A1(n12747), .A2(n13040), .B1(n15194), .B2(n12411), .ZN(
        n11405) );
  OAI211_X1 U13858 ( .C1(n13054), .C2(n15263), .A(n11406), .B(n11405), .ZN(
        n15265) );
  INV_X1 U13859 ( .A(n15265), .ZN(n11411) );
  INV_X1 U13860 ( .A(n15263), .ZN(n11409) );
  AOI22_X1 U13861 ( .A1(n12831), .A2(n11589), .B1(n15208), .B2(n11585), .ZN(
        n11407) );
  OAI21_X1 U13862 ( .B1(n8430), .B2(n15211), .A(n11407), .ZN(n11408) );
  AOI21_X1 U13863 ( .B1(n11409), .B2(n15209), .A(n11408), .ZN(n11410) );
  OAI21_X1 U13864 ( .B1(n11411), .B2(n15213), .A(n11410), .ZN(P3_U3223) );
  OAI21_X1 U13865 ( .B1(n11414), .B2(n11413), .A(n11412), .ZN(n11569) );
  INV_X1 U13866 ( .A(n11569), .ZN(n11424) );
  XNOR2_X1 U13867 ( .A(n11415), .B(n11416), .ZN(n11417) );
  OAI222_X1 U13868 ( .A1(n14287), .A2(n11824), .B1(n14285), .B2(n11418), .C1(
        n11417), .C2(n14282), .ZN(n11567) );
  NAND2_X1 U13869 ( .A1(n11567), .A2(n14313), .ZN(n11423) );
  AOI211_X1 U13870 ( .C1(n11571), .C2(n6894), .A(n14326), .B(n6640), .ZN(
        n11568) );
  INV_X1 U13871 ( .A(n11571), .ZN(n11830) );
  NOR2_X1 U13872 ( .A1(n11830), .A2(n14823), .ZN(n11421) );
  OAI22_X1 U13873 ( .A1(n14313), .A2(n11419), .B1(n11825), .B2(n14307), .ZN(
        n11420) );
  AOI211_X1 U13874 ( .C1(n11568), .C2(n14817), .A(n11421), .B(n11420), .ZN(
        n11422) );
  OAI211_X1 U13875 ( .C1(n11424), .C2(n14334), .A(n11423), .B(n11422), .ZN(
        P1_U3282) );
  AOI21_X1 U13876 ( .B1(n11427), .B2(n11426), .A(n11425), .ZN(n11440) );
  OAI21_X1 U13877 ( .B1(n11430), .B2(n11429), .A(n11428), .ZN(n11438) );
  NOR2_X1 U13878 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11431), .ZN(n11789) );
  AOI21_X1 U13879 ( .B1(n15097), .B2(P3_ADDR_REG_11__SCAN_IN), .A(n11789), 
        .ZN(n11432) );
  OAI21_X1 U13880 ( .B1(n15139), .B2(n11529), .A(n11432), .ZN(n11437) );
  AOI21_X1 U13881 ( .B1(n14684), .B2(n11434), .A(n11433), .ZN(n11435) );
  NOR2_X1 U13882 ( .A1(n11435), .A2(n15136), .ZN(n11436) );
  AOI211_X1 U13883 ( .C1(n15155), .C2(n11438), .A(n11437), .B(n11436), .ZN(
        n11439) );
  OAI21_X1 U13884 ( .B1(n11440), .B2(n15163), .A(n11439), .ZN(P3_U3193) );
  INV_X1 U13885 ( .A(n11441), .ZN(n11442) );
  AOI21_X1 U13886 ( .B1(n11444), .B2(n11443), .A(n11442), .ZN(n11460) );
  INV_X1 U13887 ( .A(n11445), .ZN(n11446) );
  AOI21_X1 U13888 ( .B1(n11448), .B2(n11447), .A(n11446), .ZN(n11450) );
  AND2_X1 U13889 ( .A1(P3_U3151), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n11593) );
  AOI21_X1 U13890 ( .B1(n15097), .B2(P3_ADDR_REG_10__SCAN_IN), .A(n11593), 
        .ZN(n11449) );
  OAI21_X1 U13891 ( .B1(n11450), .B2(n15163), .A(n11449), .ZN(n11457) );
  NAND3_X1 U13892 ( .A1(n11453), .A2(n11452), .A3(n11451), .ZN(n11454) );
  AOI21_X1 U13893 ( .B1(n11455), .B2(n11454), .A(n15131), .ZN(n11456) );
  AOI211_X1 U13894 ( .C1(n15153), .C2(n11458), .A(n11457), .B(n11456), .ZN(
        n11459) );
  OAI21_X1 U13895 ( .B1(n11460), .B2(n15136), .A(n11459), .ZN(P3_U3192) );
  INV_X1 U13896 ( .A(n11461), .ZN(n11462) );
  AOI21_X1 U13897 ( .B1(n11464), .B2(n11463), .A(n11462), .ZN(n11473) );
  NOR2_X1 U13898 ( .A1(n14013), .A2(n11465), .ZN(n11466) );
  AOI211_X1 U13899 ( .C1(n14011), .C2(n14038), .A(n11467), .B(n11466), .ZN(
        n11468) );
  OAI21_X1 U13900 ( .B1(n13989), .B2(n11469), .A(n11468), .ZN(n11470) );
  AOI21_X1 U13901 ( .B1(n11471), .B2(n14018), .A(n11470), .ZN(n11472) );
  OAI21_X1 U13902 ( .B1(n11473), .B2(n14022), .A(n11472), .ZN(P1_U3221) );
  INV_X1 U13903 ( .A(n8963), .ZN(n11474) );
  OAI222_X1 U13904 ( .A1(n13870), .A2(n7142), .B1(n13873), .B2(n11474), .C1(
        n13516), .C2(P2_U3088), .ZN(P2_U3308) );
  OAI222_X1 U13905 ( .A1(n14478), .A2(n11475), .B1(n14480), .B2(n11474), .C1(
        P1_U3086), .C2(n12108), .ZN(P1_U3336) );
  OAI21_X1 U13906 ( .B1(n11478), .B2(n11477), .A(n11476), .ZN(n11623) );
  INV_X1 U13907 ( .A(n11623), .ZN(n11491) );
  XNOR2_X1 U13908 ( .A(n11479), .B(n11480), .ZN(n11483) );
  NAND2_X1 U13909 ( .A1(n11623), .A2(n14209), .ZN(n11482) );
  AOI22_X1 U13910 ( .A1(n14321), .A2(n14032), .B1(n14034), .B2(n14319), .ZN(
        n11481) );
  OAI211_X1 U13911 ( .C1(n14282), .C2(n11483), .A(n11482), .B(n11481), .ZN(
        n11621) );
  NAND2_X1 U13912 ( .A1(n11621), .A2(n14313), .ZN(n11490) );
  OAI22_X1 U13913 ( .A1(n14313), .A2(n11484), .B1(n11899), .B2(n14307), .ZN(
        n11487) );
  INV_X1 U13914 ( .A(n11485), .ZN(n11606) );
  OAI211_X1 U13915 ( .C1(n6891), .C2(n6640), .A(n11606), .B(n14427), .ZN(
        n11620) );
  NOR2_X1 U13916 ( .A1(n11620), .A2(n14243), .ZN(n11486) );
  AOI211_X1 U13917 ( .C1(n14346), .C2(n11488), .A(n11487), .B(n11486), .ZN(
        n11489) );
  OAI211_X1 U13918 ( .C1(n11491), .C2(n14165), .A(n11490), .B(n11489), .ZN(
        P1_U3281) );
  INV_X1 U13919 ( .A(n11492), .ZN(n11522) );
  OAI222_X1 U13920 ( .A1(P1_U3086), .A2(n11493), .B1(n14478), .B2(n7985), .C1(
        n11522), .C2(n14480), .ZN(P1_U3335) );
  XNOR2_X1 U13921 ( .A(n12151), .B(n12413), .ZN(n11586) );
  XNOR2_X1 U13922 ( .A(n11586), .B(n12412), .ZN(n11500) );
  NAND2_X1 U13923 ( .A1(n11494), .A2(n12749), .ZN(n11495) );
  INV_X1 U13924 ( .A(n11500), .ZN(n11497) );
  INV_X1 U13925 ( .A(n11588), .ZN(n11498) );
  AOI21_X1 U13926 ( .B1(n11500), .B2(n11499), .A(n11498), .ZN(n11507) );
  OAI22_X1 U13927 ( .A1(n12723), .A2(n11542), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n11501), .ZN(n11504) );
  OAI22_X1 U13928 ( .A1(n12717), .A2(n15254), .B1(n11502), .B2(n12736), .ZN(
        n11503) );
  AOI211_X1 U13929 ( .C1(n11505), .C2(n12732), .A(n11504), .B(n11503), .ZN(
        n11506) );
  OAI21_X1 U13930 ( .B1(n11507), .B2(n12741), .A(n11506), .ZN(P3_U3171) );
  AOI21_X1 U13931 ( .B1(n11510), .B2(n11509), .A(n11508), .ZN(n11521) );
  XNOR2_X1 U13932 ( .A(n6636), .B(n11511), .ZN(n11519) );
  INV_X1 U13933 ( .A(n15136), .ZN(n15158) );
  AOI211_X1 U13934 ( .C1(n11514), .C2(n11513), .A(n15131), .B(n11512), .ZN(
        n11518) );
  AND2_X1 U13935 ( .A1(P3_U3151), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n11912) );
  AOI21_X1 U13936 ( .B1(n15097), .B2(P3_ADDR_REG_12__SCAN_IN), .A(n11912), 
        .ZN(n11515) );
  OAI21_X1 U13937 ( .B1(n15139), .B2(n11516), .A(n11515), .ZN(n11517) );
  AOI211_X1 U13938 ( .C1(n11519), .C2(n15158), .A(n11518), .B(n11517), .ZN(
        n11520) );
  OAI21_X1 U13939 ( .B1(n11521), .B2(n15163), .A(n11520), .ZN(P3_U3194) );
  OAI222_X1 U13940 ( .A1(n13870), .A2(n7139), .B1(P2_U3088), .B2(n11523), .C1(
        n13873), .C2(n11522), .ZN(P2_U3307) );
  NAND2_X1 U13941 ( .A1(n13054), .A2(n15186), .ZN(n11524) );
  NAND2_X1 U13942 ( .A1(n15211), .A2(n11524), .ZN(n12877) );
  INV_X1 U13943 ( .A(n11525), .ZN(n12519) );
  NAND2_X1 U13944 ( .A1(n11526), .A2(n12519), .ZN(n11527) );
  NAND2_X1 U13945 ( .A1(n11528), .A2(n12311), .ZN(n11532) );
  AOI22_X1 U13946 ( .A1(n12332), .A2(n11530), .B1(n12162), .B2(n11529), .ZN(
        n11531) );
  NAND2_X1 U13947 ( .A1(n11532), .A2(n11531), .ZN(n14679) );
  NAND2_X1 U13948 ( .A1(n14679), .A2(n12747), .ZN(n12424) );
  XNOR2_X1 U13949 ( .A(n11692), .B(n12522), .ZN(n14681) );
  NAND2_X1 U13950 ( .A1(n12155), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n11539) );
  NAND2_X1 U13951 ( .A1(n6491), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n11538) );
  OR2_X1 U13952 ( .A1(n11534), .A2(n11533), .ZN(n11535) );
  NAND2_X1 U13953 ( .A1(n11675), .A2(n11535), .ZN(n11911) );
  NAND2_X1 U13954 ( .A1(n10235), .A2(n11911), .ZN(n11537) );
  NAND2_X1 U13955 ( .A1(n10454), .A2(P3_REG0_REG_12__SCAN_IN), .ZN(n11536) );
  XNOR2_X1 U13956 ( .A(n11686), .B(n12522), .ZN(n11541) );
  OAI222_X1 U13957 ( .A1(n15197), .A2(n11926), .B1(n15173), .B2(n11542), .C1(
        n11541), .C2(n15178), .ZN(n14683) );
  NAND2_X1 U13958 ( .A1(n14683), .A2(n15211), .ZN(n11546) );
  INV_X1 U13959 ( .A(n11792), .ZN(n11543) );
  OAI22_X1 U13960 ( .A1(n13047), .A2(n14679), .B1(n11543), .B2(n11954), .ZN(
        n11544) );
  AOI21_X1 U13961 ( .B1(n15213), .B2(P3_REG2_REG_11__SCAN_IN), .A(n11544), 
        .ZN(n11545) );
  OAI211_X1 U13962 ( .C1(n12877), .C2(n14681), .A(n11546), .B(n11545), .ZN(
        P3_U3222) );
  NOR2_X1 U13963 ( .A1(n14704), .A2(n14705), .ZN(n14703) );
  NAND2_X1 U13964 ( .A1(n11550), .A2(n11560), .ZN(n11804) );
  OAI21_X1 U13965 ( .B1(n11550), .B2(n11560), .A(n11804), .ZN(n14731) );
  INV_X1 U13966 ( .A(n14731), .ZN(n11566) );
  INV_X1 U13967 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n11551) );
  OAI22_X1 U13968 ( .A1(n15002), .A2(n11551), .B1(n11726), .B2(n14996), .ZN(
        n11554) );
  INV_X1 U13969 ( .A(n11802), .ZN(n14728) );
  INV_X1 U13970 ( .A(n14707), .ZN(n11552) );
  OAI211_X1 U13971 ( .C1(n14728), .C2(n11552), .A(n10086), .B(n11797), .ZN(
        n14727) );
  NOR2_X1 U13972 ( .A1(n14727), .A2(n14983), .ZN(n11553) );
  AOI211_X1 U13973 ( .C1(n14715), .C2(n11802), .A(n11554), .B(n11553), .ZN(
        n11565) );
  NAND2_X1 U13974 ( .A1(n11638), .A2(n11556), .ZN(n11557) );
  XOR2_X1 U13975 ( .A(n11795), .B(n11560), .Z(n11561) );
  NOR2_X1 U13976 ( .A1(n11561), .A2(n14997), .ZN(n14730) );
  AND2_X1 U13977 ( .A1(n13420), .A2(n13436), .ZN(n11562) );
  AOI21_X1 U13978 ( .B1(n13434), .B2(n13524), .A(n11562), .ZN(n14726) );
  INV_X1 U13979 ( .A(n14726), .ZN(n11563) );
  OAI21_X1 U13980 ( .B1(n14730), .B2(n11563), .A(n15002), .ZN(n11564) );
  OAI211_X1 U13981 ( .C1(n11566), .C2(n13739), .A(n11565), .B(n11564), .ZN(
        P2_U3250) );
  AOI211_X1 U13982 ( .C1(n14848), .C2(n11569), .A(n11568), .B(n11567), .ZN(
        n11573) );
  AOI22_X1 U13983 ( .A1(n11571), .A2(n11753), .B1(P1_REG0_REG_11__SCAN_IN), 
        .B2(n6786), .ZN(n11570) );
  OAI21_X1 U13984 ( .B1(n11573), .B2(n6786), .A(n11570), .ZN(P1_U3492) );
  AOI22_X1 U13985 ( .A1(n11571), .A2(n14375), .B1(P1_REG1_REG_11__SCAN_IN), 
        .B2(n14854), .ZN(n11572) );
  OAI21_X1 U13986 ( .B1(n11573), .B2(n14854), .A(n11572), .ZN(P1_U3539) );
  NAND2_X1 U13987 ( .A1(n11575), .A2(n11574), .ZN(n12099) );
  XOR2_X1 U13988 ( .A(n12100), .B(n12099), .Z(n11576) );
  NAND2_X1 U13989 ( .A1(P1_REG2_REG_18__SCAN_IN), .A2(n11576), .ZN(n12101) );
  OAI211_X1 U13990 ( .C1(n11576), .C2(P1_REG2_REG_18__SCAN_IN), .A(n14113), 
        .B(n12101), .ZN(n11583) );
  NAND2_X1 U13991 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n13983)
         );
  INV_X1 U13992 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n14421) );
  OAI21_X1 U13993 ( .B1(n14421), .B2(n11578), .A(n11577), .ZN(n12095) );
  XNOR2_X1 U13994 ( .A(n12095), .B(n11584), .ZN(n11579) );
  NAND2_X1 U13995 ( .A1(P1_REG1_REG_18__SCAN_IN), .A2(n11579), .ZN(n12097) );
  OAI211_X1 U13996 ( .C1(P1_REG1_REG_18__SCAN_IN), .C2(n11579), .A(n14102), 
        .B(n12097), .ZN(n11580) );
  NAND2_X1 U13997 ( .A1(n13983), .A2(n11580), .ZN(n11581) );
  AOI21_X1 U13998 ( .B1(n14088), .B2(P1_ADDR_REG_18__SCAN_IN), .A(n11581), 
        .ZN(n11582) );
  OAI211_X1 U13999 ( .C1(n14811), .C2(n11584), .A(n11583), .B(n11582), .ZN(
        P1_U3261) );
  INV_X1 U14000 ( .A(n11585), .ZN(n11597) );
  NAND2_X1 U14001 ( .A1(n11586), .A2(n12412), .ZN(n11587) );
  XNOR2_X1 U14002 ( .A(n12151), .B(n11589), .ZN(n11781) );
  XNOR2_X1 U14003 ( .A(n11781), .B(n12748), .ZN(n11590) );
  OAI211_X1 U14004 ( .C1(n11591), .C2(n11590), .A(n6685), .B(n12709), .ZN(
        n11595) );
  OAI22_X1 U14005 ( .A1(n12717), .A2(n15260), .B1(n12412), .B2(n12736), .ZN(
        n11592) );
  AOI211_X1 U14006 ( .C1(n12733), .C2(n12747), .A(n11593), .B(n11592), .ZN(
        n11594) );
  OAI211_X1 U14007 ( .C1(n11597), .C2(n11596), .A(n11595), .B(n11594), .ZN(
        P3_U3157) );
  OAI21_X1 U14008 ( .B1(n11600), .B2(n11599), .A(n11598), .ZN(n11734) );
  INV_X1 U14009 ( .A(n11734), .ZN(n11612) );
  XNOR2_X1 U14010 ( .A(n11603), .B(n11602), .ZN(n11604) );
  OAI222_X1 U14011 ( .A1(n14287), .A2(n12025), .B1(n14285), .B2(n11824), .C1(
        n11604), .C2(n14282), .ZN(n11732) );
  NAND2_X1 U14012 ( .A1(n11732), .A2(n14313), .ZN(n11611) );
  INV_X1 U14013 ( .A(n11642), .ZN(n11605) );
  AOI211_X1 U14014 ( .C1(n11736), .C2(n11606), .A(n14326), .B(n11605), .ZN(
        n11733) );
  NOR2_X1 U14015 ( .A1(n12031), .A2(n14823), .ZN(n11609) );
  OAI22_X1 U14016 ( .A1(n14313), .A2(n11607), .B1(n12026), .B2(n14307), .ZN(
        n11608) );
  AOI211_X1 U14017 ( .C1(n11733), .C2(n14817), .A(n11609), .B(n11608), .ZN(
        n11610) );
  OAI211_X1 U14018 ( .C1(n11612), .C2(n14334), .A(n11611), .B(n11610), .ZN(
        P1_U3280) );
  INV_X1 U14019 ( .A(n11613), .ZN(n11618) );
  OAI222_X1 U14020 ( .A1(n14478), .A2(n11615), .B1(n14480), .B2(n11618), .C1(
        P1_U3086), .C2(n11614), .ZN(P1_U3334) );
  INV_X1 U14021 ( .A(n11616), .ZN(n11617) );
  OAI222_X1 U14022 ( .A1(n13870), .A2(n11619), .B1(n13873), .B2(n11618), .C1(
        n11617), .C2(P2_U3088), .ZN(P2_U3306) );
  OAI21_X1 U14023 ( .B1(n6891), .B2(n14843), .A(n11620), .ZN(n11622) );
  AOI211_X1 U14024 ( .C1(n14381), .C2(n11623), .A(n11622), .B(n11621), .ZN(
        n11626) );
  NAND2_X1 U14025 ( .A1(n6786), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n11624) );
  OAI21_X1 U14026 ( .B1(n11626), .B2(n6786), .A(n11624), .ZN(P1_U3495) );
  NAND2_X1 U14027 ( .A1(n14854), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n11625) );
  OAI21_X1 U14028 ( .B1(n11626), .B2(n14854), .A(n11625), .ZN(P1_U3540) );
  NAND2_X1 U14029 ( .A1(n13422), .A2(n11627), .ZN(n11628) );
  NAND2_X1 U14030 ( .A1(P2_U3088), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n14899)
         );
  OAI211_X1 U14031 ( .C1(n13424), .C2(n14741), .A(n11628), .B(n14899), .ZN(
        n11637) );
  XNOR2_X1 U14032 ( .A(n11638), .B(n12611), .ZN(n11630) );
  AND2_X1 U14033 ( .A1(n13437), .A2(n12605), .ZN(n11629) );
  NAND2_X1 U14034 ( .A1(n11630), .A2(n11629), .ZN(n11666) );
  OAI21_X1 U14035 ( .B1(n11630), .B2(n11629), .A(n11666), .ZN(n11635) );
  AOI211_X1 U14036 ( .C1(n11635), .C2(n11634), .A(n13428), .B(n11667), .ZN(
        n11636) );
  AOI211_X1 U14037 ( .C1(n11638), .C2(n13426), .A(n11637), .B(n11636), .ZN(
        n11639) );
  INV_X1 U14038 ( .A(n11639), .ZN(P2_U3206) );
  OAI21_X1 U14039 ( .B1(n11641), .B2(n9481), .A(n11640), .ZN(n11749) );
  AOI21_X1 U14040 ( .B1(n13892), .B2(n11642), .A(n14326), .ZN(n11643) );
  AND2_X1 U14041 ( .A1(n11643), .A2(n11773), .ZN(n11750) );
  NAND2_X1 U14042 ( .A1(n13892), .A2(n14346), .ZN(n11646) );
  NOR2_X1 U14043 ( .A1(n14307), .A2(n13890), .ZN(n11644) );
  AOI21_X1 U14044 ( .B1(n14830), .B2(P1_REG2_REG_14__SCAN_IN), .A(n11644), 
        .ZN(n11645) );
  NAND2_X1 U14045 ( .A1(n11646), .A2(n11645), .ZN(n11647) );
  AOI21_X1 U14046 ( .B1(n11750), .B2(n14817), .A(n11647), .ZN(n11655) );
  XNOR2_X1 U14047 ( .A(n11650), .B(n11649), .ZN(n11651) );
  NOR2_X1 U14048 ( .A1(n11651), .A2(n14282), .ZN(n11751) );
  NAND2_X1 U14049 ( .A1(n14032), .A2(n14319), .ZN(n11653) );
  NAND2_X1 U14050 ( .A1(n14030), .A2(n14321), .ZN(n11652) );
  NAND2_X1 U14051 ( .A1(n11653), .A2(n11652), .ZN(n13887) );
  OAI21_X1 U14052 ( .B1(n11751), .B2(n13887), .A(n14313), .ZN(n11654) );
  OAI211_X1 U14053 ( .C1(n11749), .C2(n14334), .A(n11655), .B(n11654), .ZN(
        P1_U3279) );
  NOR2_X1 U14054 ( .A1(n11656), .A2(n6643), .ZN(n11657) );
  XNOR2_X1 U14055 ( .A(n6647), .B(n11657), .ZN(n11665) );
  NAND2_X1 U14056 ( .A1(n13999), .A2(n11658), .ZN(n11659) );
  OAI211_X1 U14057 ( .C1(n13989), .C2(n11661), .A(n11660), .B(n11659), .ZN(
        n11662) );
  AOI21_X1 U14058 ( .B1(n11663), .B2(n14018), .A(n11662), .ZN(n11664) );
  OAI21_X1 U14059 ( .B1(n11665), .B2(n14022), .A(n11664), .ZN(P1_U3217) );
  XNOR2_X1 U14060 ( .A(n14702), .B(n12611), .ZN(n11720) );
  NAND2_X1 U14061 ( .A1(n13436), .A2(n12610), .ZN(n11721) );
  XNOR2_X1 U14062 ( .A(n11720), .B(n11721), .ZN(n11668) );
  OAI21_X1 U14063 ( .B1(n11669), .B2(n11668), .A(n6711), .ZN(n11670) );
  NAND2_X1 U14064 ( .A1(n11670), .A2(n13391), .ZN(n11674) );
  AOI22_X1 U14065 ( .A1(n13435), .A2(n13524), .B1(n13420), .B2(n13437), .ZN(
        n14698) );
  OAI22_X1 U14066 ( .A1(n13424), .A2(n14698), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n11671), .ZN(n11672) );
  AOI21_X1 U14067 ( .B1(n14701), .B2(n13422), .A(n11672), .ZN(n11673) );
  OAI211_X1 U14068 ( .C1(n14735), .C2(n13415), .A(n11674), .B(n11673), .ZN(
        P2_U3187) );
  NAND2_X1 U14069 ( .A1(n12268), .A2(P3_REG2_REG_13__SCAN_IN), .ZN(n11680) );
  NAND2_X1 U14070 ( .A1(n10454), .A2(P3_REG0_REG_13__SCAN_IN), .ZN(n11679) );
  NAND2_X1 U14071 ( .A1(n11675), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n11676) );
  NAND2_X1 U14072 ( .A1(n11706), .A2(n11676), .ZN(n11929) );
  NAND2_X1 U14073 ( .A1(n10235), .A2(n11929), .ZN(n11678) );
  NAND2_X1 U14074 ( .A1(n6491), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n11677) );
  NAND4_X1 U14075 ( .A1(n11680), .A2(n11679), .A3(n11678), .A4(n11677), .ZN(
        n12745) );
  NAND2_X1 U14076 ( .A1(n11681), .A2(n12311), .ZN(n11684) );
  AOI22_X1 U14077 ( .A1(n12332), .A2(SI_12_), .B1(n12162), .B2(n11682), .ZN(
        n11683) );
  NAND2_X1 U14078 ( .A1(n11684), .A2(n11683), .ZN(n11917) );
  OR2_X1 U14079 ( .A1(n11917), .A2(n11926), .ZN(n12429) );
  NAND2_X1 U14080 ( .A1(n11917), .A2(n11926), .ZN(n12428) );
  NAND2_X1 U14081 ( .A1(n14679), .A2(n11915), .ZN(n11685) );
  NAND2_X1 U14082 ( .A1(n11686), .A2(n11685), .ZN(n11688) );
  OR2_X1 U14083 ( .A1(n14679), .A2(n11915), .ZN(n11687) );
  OR2_X2 U14084 ( .A1(n11690), .A2(n12525), .ZN(n11700) );
  INV_X1 U14085 ( .A(n11700), .ZN(n11689) );
  AOI21_X1 U14086 ( .B1(n12525), .B2(n11690), .A(n11689), .ZN(n11691) );
  OAI222_X1 U14087 ( .A1(n15197), .A2(n12017), .B1(n15173), .B2(n11915), .C1(
        n15178), .C2(n11691), .ZN(n14675) );
  INV_X1 U14088 ( .A(n14675), .ZN(n11698) );
  NAND2_X1 U14089 ( .A1(n11692), .A2(n12421), .ZN(n11693) );
  OAI21_X1 U14090 ( .B1(n11694), .B2(n12525), .A(n11714), .ZN(n14677) );
  INV_X1 U14091 ( .A(n11917), .ZN(n14674) );
  AOI22_X1 U14092 ( .A1(n15213), .A2(P3_REG2_REG_12__SCAN_IN), .B1(n15208), 
        .B2(n11911), .ZN(n11695) );
  OAI21_X1 U14093 ( .B1(n14674), .B2(n13047), .A(n11695), .ZN(n11696) );
  AOI21_X1 U14094 ( .B1(n14677), .B2(n13050), .A(n11696), .ZN(n11697) );
  OAI21_X1 U14095 ( .B1(n11698), .B2(n15213), .A(n11697), .ZN(P3_U3221) );
  INV_X1 U14096 ( .A(n11926), .ZN(n12746) );
  OR2_X1 U14097 ( .A1(n11917), .A2(n12746), .ZN(n11699) );
  NAND2_X1 U14098 ( .A1(n11701), .A2(n12311), .ZN(n11704) );
  AOI22_X1 U14099 ( .A1(n12332), .A2(n11702), .B1(n12162), .B2(n12764), .ZN(
        n11703) );
  NAND2_X1 U14100 ( .A1(n11704), .A2(n11703), .ZN(n14669) );
  OR2_X1 U14101 ( .A1(n14669), .A2(n12745), .ZN(n12362) );
  NAND2_X1 U14102 ( .A1(n14669), .A2(n12745), .ZN(n12361) );
  NAND2_X1 U14103 ( .A1(n12362), .A2(n12361), .ZN(n11715) );
  OAI211_X1 U14104 ( .C1(n11705), .C2(n11715), .A(n11952), .B(n15200), .ZN(
        n11713) );
  NAND2_X1 U14105 ( .A1(n12155), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n11711) );
  NAND2_X1 U14106 ( .A1(n6491), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n11710) );
  AND2_X1 U14107 ( .A1(n11706), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n11707) );
  OR2_X1 U14108 ( .A1(n11707), .A2(n11945), .ZN(n12014) );
  NAND2_X1 U14109 ( .A1(n10235), .A2(n12014), .ZN(n11709) );
  NAND2_X1 U14110 ( .A1(n10454), .A2(P3_REG0_REG_14__SCAN_IN), .ZN(n11708) );
  AOI22_X1 U14111 ( .A1(n13040), .A2(n12744), .B1(n12746), .B2(n15194), .ZN(
        n11712) );
  NAND2_X1 U14112 ( .A1(n11713), .A2(n11712), .ZN(n14670) );
  INV_X1 U14113 ( .A(n14670), .ZN(n11719) );
  XNOR2_X1 U14114 ( .A(n11939), .B(n12526), .ZN(n14672) );
  AOI22_X1 U14115 ( .A1(n15213), .A2(P3_REG2_REG_13__SCAN_IN), .B1(n15208), 
        .B2(n11929), .ZN(n11716) );
  OAI21_X1 U14116 ( .B1(n14669), .B2(n13047), .A(n11716), .ZN(n11717) );
  AOI21_X1 U14117 ( .B1(n14672), .B2(n13050), .A(n11717), .ZN(n11718) );
  OAI21_X1 U14118 ( .B1(n11719), .B2(n15213), .A(n11718), .ZN(P3_U3220) );
  INV_X1 U14119 ( .A(n6711), .ZN(n11723) );
  INV_X1 U14120 ( .A(n11720), .ZN(n11722) );
  AND2_X1 U14121 ( .A1(n11722), .A2(n11721), .ZN(n11855) );
  NOR2_X1 U14122 ( .A1(n11723), .A2(n11855), .ZN(n11725) );
  XNOR2_X1 U14123 ( .A(n11802), .B(n9992), .ZN(n11857) );
  NAND2_X1 U14124 ( .A1(n13435), .A2(n12610), .ZN(n11856) );
  INV_X1 U14125 ( .A(n11856), .ZN(n11858) );
  XNOR2_X1 U14126 ( .A(n11857), .B(n11858), .ZN(n11724) );
  XNOR2_X1 U14127 ( .A(n11725), .B(n11724), .ZN(n11731) );
  NOR2_X1 U14128 ( .A1(n13372), .A2(n11726), .ZN(n11729) );
  OAI22_X1 U14129 ( .A1(n13424), .A2(n14726), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n11727), .ZN(n11728) );
  AOI211_X1 U14130 ( .C1(n11802), .C2(n13426), .A(n11729), .B(n11728), .ZN(
        n11730) );
  OAI21_X1 U14131 ( .B1(n11731), .B2(n13428), .A(n11730), .ZN(P2_U3213) );
  AOI211_X1 U14132 ( .C1(n14848), .C2(n11734), .A(n11733), .B(n11732), .ZN(
        n11738) );
  AOI22_X1 U14133 ( .A1(n11736), .A2(n11753), .B1(P1_REG0_REG_13__SCAN_IN), 
        .B2(n6786), .ZN(n11735) );
  OAI21_X1 U14134 ( .B1(n11738), .B2(n6786), .A(n11735), .ZN(P1_U3498) );
  AOI22_X1 U14135 ( .A1(n11736), .A2(n14375), .B1(P1_REG1_REG_13__SCAN_IN), 
        .B2(n14854), .ZN(n11737) );
  OAI21_X1 U14136 ( .B1(n11738), .B2(n14854), .A(n11737), .ZN(P1_U3541) );
  NAND2_X1 U14137 ( .A1(n11742), .A2(n11819), .ZN(n11744) );
  NAND2_X1 U14138 ( .A1(n11744), .A2(n11743), .ZN(n11872) );
  AOI22_X1 U14139 ( .A1(P2_DATAO_REG_25__SCAN_IN), .A2(n11881), .B1(
        P1_DATAO_REG_25__SCAN_IN), .B2(n6678), .ZN(n11873) );
  INV_X1 U14140 ( .A(n11873), .ZN(n11745) );
  XNOR2_X1 U14141 ( .A(n11872), .B(n11745), .ZN(n12238) );
  INV_X1 U14142 ( .A(n12238), .ZN(n11746) );
  OAI222_X1 U14143 ( .A1(n11748), .A2(P3_U3151), .B1(n13335), .B2(n11747), 
        .C1(n13333), .C2(n11746), .ZN(P3_U3270) );
  NOR2_X1 U14144 ( .A1(n11749), .A2(n14431), .ZN(n11752) );
  NOR4_X1 U14145 ( .A1(n11752), .A2(n11751), .A3(n11750), .A4(n13887), .ZN(
        n11756) );
  AOI22_X1 U14146 ( .A1(n13892), .A2(n11753), .B1(P1_REG0_REG_14__SCAN_IN), 
        .B2(n6786), .ZN(n11754) );
  OAI21_X1 U14147 ( .B1(n11756), .B2(n6786), .A(n11754), .ZN(P1_U3501) );
  AOI22_X1 U14148 ( .A1(n13892), .A2(n14375), .B1(P1_REG1_REG_14__SCAN_IN), 
        .B2(n14854), .ZN(n11755) );
  OAI21_X1 U14149 ( .B1(n11756), .B2(n14854), .A(n11755), .ZN(P1_U3542) );
  NAND2_X1 U14150 ( .A1(n13987), .A2(n14035), .ZN(n11761) );
  NAND2_X1 U14151 ( .A1(n14016), .A2(n11757), .ZN(n11759) );
  NAND2_X1 U14152 ( .A1(n14011), .A2(n14037), .ZN(n11758) );
  NAND4_X1 U14153 ( .A1(n11761), .A2(n11760), .A3(n11759), .A4(n11758), .ZN(
        n11766) );
  XNOR2_X1 U14154 ( .A(n11763), .B(n11762), .ZN(n11764) );
  NOR2_X1 U14155 ( .A1(n11764), .A2(n14022), .ZN(n11765) );
  AOI211_X1 U14156 ( .C1(n11767), .C2(n14018), .A(n11766), .B(n11765), .ZN(
        n11768) );
  INV_X1 U14157 ( .A(n11768), .ZN(P1_U3231) );
  XNOR2_X1 U14158 ( .A(n11769), .B(n11771), .ZN(n11770) );
  OAI222_X1 U14159 ( .A1(n14287), .A2(n14014), .B1(n14285), .B2(n12025), .C1(
        n14282), .C2(n11770), .ZN(n11933) );
  INV_X1 U14160 ( .A(n11933), .ZN(n11780) );
  XNOR2_X1 U14161 ( .A(n11772), .B(n11771), .ZN(n11935) );
  NAND2_X1 U14162 ( .A1(n14019), .A2(n11773), .ZN(n11774) );
  NAND2_X1 U14163 ( .A1(n11840), .A2(n11774), .ZN(n11932) );
  INV_X1 U14164 ( .A(n14344), .ZN(n11777) );
  AOI22_X1 U14165 ( .A1(n14830), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n14017), 
        .B2(n14819), .ZN(n11776) );
  NAND2_X1 U14166 ( .A1(n14019), .A2(n14346), .ZN(n11775) );
  OAI211_X1 U14167 ( .C1(n11932), .C2(n11777), .A(n11776), .B(n11775), .ZN(
        n11778) );
  AOI21_X1 U14168 ( .B1(n11935), .B2(n14277), .A(n11778), .ZN(n11779) );
  OAI21_X1 U14169 ( .B1(n11780), .B2(n14830), .A(n11779), .ZN(P1_U3278) );
  INV_X1 U14170 ( .A(n11781), .ZN(n11782) );
  NAND2_X1 U14171 ( .A1(n11782), .A2(n12748), .ZN(n11783) );
  XNOR2_X1 U14172 ( .A(n12292), .B(n14679), .ZN(n11785) );
  INV_X1 U14173 ( .A(n11785), .ZN(n11786) );
  NAND2_X1 U14174 ( .A1(n11904), .A2(n11905), .ZN(n11787) );
  XNOR2_X1 U14175 ( .A(n11787), .B(n11915), .ZN(n11794) );
  NOR2_X1 U14176 ( .A1(n12723), .A2(n11926), .ZN(n11788) );
  AOI211_X1 U14177 ( .C1(n12720), .C2(n12748), .A(n11789), .B(n11788), .ZN(
        n11790) );
  OAI21_X1 U14178 ( .B1(n12717), .B2(n14679), .A(n11790), .ZN(n11791) );
  AOI21_X1 U14179 ( .B1(n11792), .B2(n12732), .A(n11791), .ZN(n11793) );
  OAI21_X1 U14180 ( .B1(n11794), .B2(n12741), .A(n11793), .ZN(P3_U3176) );
  XOR2_X1 U14181 ( .A(n11960), .B(n11959), .Z(n11851) );
  AOI21_X1 U14182 ( .B1(n11964), .B2(n11797), .A(n12610), .ZN(n11798) );
  NAND2_X1 U14183 ( .A1(n11798), .A2(n11966), .ZN(n11847) );
  AOI22_X1 U14184 ( .A1(n13567), .A2(n13524), .B1(n13420), .B2(n13435), .ZN(
        n11867) );
  OAI22_X1 U14185 ( .A1(n15005), .A2(n11867), .B1(n11865), .B2(n14996), .ZN(
        n11800) );
  NOR2_X1 U14186 ( .A1(n6949), .A2(n14968), .ZN(n11799) );
  AOI211_X1 U14187 ( .C1(n15005), .C2(P2_REG2_REG_16__SCAN_IN), .A(n11800), 
        .B(n11799), .ZN(n11801) );
  OAI21_X1 U14188 ( .B1(n14983), .B2(n11847), .A(n11801), .ZN(n11807) );
  AND2_X1 U14189 ( .A1(n11805), .A2(n11959), .ZN(n11848) );
  NOR3_X1 U14190 ( .A1(n11963), .A2(n11848), .A3(n13739), .ZN(n11806) );
  AOI211_X1 U14191 ( .C1(n13737), .C2(n11851), .A(n11807), .B(n11806), .ZN(
        n11808) );
  INV_X1 U14192 ( .A(n11808), .ZN(P2_U3249) );
  NAND2_X1 U14193 ( .A1(n11810), .A2(n11809), .ZN(n11811) );
  OAI222_X1 U14194 ( .A1(n13870), .A2(n11813), .B1(P2_U3088), .B2(n11812), 
        .C1(n13873), .C2(n11811), .ZN(P2_U3305) );
  INV_X1 U14195 ( .A(n11814), .ZN(n11818) );
  OAI222_X1 U14196 ( .A1(n13870), .A2(n11816), .B1(n13873), .B2(n11818), .C1(
        P2_U3088), .C2(n11815), .ZN(P2_U3303) );
  OAI222_X1 U14197 ( .A1(n14478), .A2(n11819), .B1(n14480), .B2(n11818), .C1(
        P1_U3086), .C2(n11817), .ZN(P1_U3331) );
  OAI21_X1 U14198 ( .B1(n11822), .B2(n11821), .A(n11820), .ZN(n11823) );
  NAND2_X1 U14199 ( .A1(n11823), .A2(n13995), .ZN(n11829) );
  NAND2_X1 U14200 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n14104)
         );
  OAI21_X1 U14201 ( .B1(n14013), .B2(n11824), .A(n14104), .ZN(n11827) );
  NOR2_X1 U14202 ( .A1(n13989), .A2(n11825), .ZN(n11826) );
  AOI211_X1 U14203 ( .C1(n14011), .C2(n14035), .A(n11827), .B(n11826), .ZN(
        n11828) );
  OAI211_X1 U14204 ( .C1(n11830), .C2(n13980), .A(n11829), .B(n11828), .ZN(
        P1_U3236) );
  OAI21_X1 U14205 ( .B1(n11833), .B2(n11832), .A(n11831), .ZN(n11836) );
  AND2_X1 U14206 ( .A1(n14030), .A2(n14319), .ZN(n11834) );
  AOI21_X1 U14207 ( .B1(n14320), .B2(n14321), .A(n11834), .ZN(n13938) );
  INV_X1 U14208 ( .A(n13938), .ZN(n11835) );
  AOI21_X1 U14209 ( .B1(n11836), .B2(n14324), .A(n11835), .ZN(n14430) );
  OAI21_X1 U14210 ( .B1(n11839), .B2(n11838), .A(n11837), .ZN(n14424) );
  INV_X1 U14211 ( .A(n14425), .ZN(n11844) );
  NAND2_X1 U14212 ( .A1(n14425), .A2(n11840), .ZN(n11841) );
  AND2_X1 U14213 ( .A1(n12033), .A2(n11841), .ZN(n14428) );
  NAND2_X1 U14214 ( .A1(n14428), .A2(n14344), .ZN(n11843) );
  AOI22_X1 U14215 ( .A1(n14830), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n13934), 
        .B2(n14819), .ZN(n11842) );
  OAI211_X1 U14216 ( .C1(n11844), .C2(n14823), .A(n11843), .B(n11842), .ZN(
        n11845) );
  AOI21_X1 U14217 ( .B1(n14424), .B2(n14277), .A(n11845), .ZN(n11846) );
  OAI21_X1 U14218 ( .B1(n14430), .B2(n14830), .A(n11846), .ZN(P1_U3277) );
  OAI211_X1 U14219 ( .C1(n6949), .C2(n15077), .A(n11847), .B(n11867), .ZN(
        n11850) );
  NOR3_X1 U14220 ( .A1(n11963), .A2(n11848), .A3(n15061), .ZN(n11849) );
  AOI211_X1 U14221 ( .C1(n15064), .C2(n11851), .A(n11850), .B(n11849), .ZN(
        n11854) );
  NAND2_X1 U14222 ( .A1(n15094), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n11852) );
  OAI21_X1 U14223 ( .B1(n11854), .B2(n15094), .A(n11852), .ZN(P2_U3515) );
  INV_X1 U14224 ( .A(n15066), .ZN(n15083) );
  NAND2_X1 U14225 ( .A1(n15083), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n11853) );
  OAI21_X1 U14226 ( .B1(n11854), .B2(n15083), .A(n11853), .ZN(P2_U3478) );
  AOI21_X1 U14227 ( .B1(n11857), .B2(n11856), .A(n11855), .ZN(n11860) );
  INV_X1 U14228 ( .A(n11857), .ZN(n11859) );
  XNOR2_X1 U14229 ( .A(n11964), .B(n12611), .ZN(n11996) );
  NAND2_X1 U14230 ( .A1(n13434), .A2(n12610), .ZN(n11994) );
  XNOR2_X1 U14231 ( .A(n11996), .B(n11994), .ZN(n11862) );
  OAI21_X1 U14232 ( .B1(n11863), .B2(n11862), .A(n11997), .ZN(n11864) );
  NAND2_X1 U14233 ( .A1(n11864), .A2(n13391), .ZN(n11871) );
  INV_X1 U14234 ( .A(n11865), .ZN(n11869) );
  OAI22_X1 U14235 ( .A1(n13424), .A2(n11867), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n11866), .ZN(n11868) );
  AOI21_X1 U14236 ( .B1(n11869), .B2(n13422), .A(n11868), .ZN(n11870) );
  OAI211_X1 U14237 ( .C1(n6949), .C2(n13415), .A(n11871), .B(n11870), .ZN(
        P2_U3198) );
  NAND2_X1 U14238 ( .A1(n11873), .A2(n11872), .ZN(n11874) );
  AOI22_X1 U14239 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(n9094), .B1(
        P1_DATAO_REG_26__SCAN_IN), .B2(n12008), .ZN(n12086) );
  INV_X1 U14240 ( .A(n12086), .ZN(n11875) );
  XNOR2_X1 U14241 ( .A(n12085), .B(n11875), .ZN(n12250) );
  INV_X1 U14242 ( .A(n12250), .ZN(n11876) );
  OAI222_X1 U14243 ( .A1(n11878), .A2(P3_U3151), .B1(n13335), .B2(n11877), 
        .C1(n13333), .C2(n11876), .ZN(P3_U3269) );
  INV_X1 U14244 ( .A(n11879), .ZN(n11883) );
  OAI222_X1 U14245 ( .A1(n13870), .A2(n11881), .B1(n13873), .B2(n11883), .C1(
        P2_U3088), .C2(n11880), .ZN(P2_U3302) );
  OAI222_X1 U14246 ( .A1(n14478), .A2(n6678), .B1(n14480), .B2(n11883), .C1(
        P1_U3086), .C2(n11882), .ZN(P1_U3330) );
  NAND2_X1 U14247 ( .A1(n11888), .A2(n11884), .ZN(n11886) );
  OAI211_X1 U14248 ( .C1(n11887), .C2(n14478), .A(n11886), .B(n11885), .ZN(
        P1_U3332) );
  NAND2_X1 U14249 ( .A1(n11888), .A2(n12078), .ZN(n11891) );
  INV_X1 U14250 ( .A(n11889), .ZN(n11890) );
  OAI211_X1 U14251 ( .C1(n11892), .C2(n13870), .A(n11891), .B(n11890), .ZN(
        P2_U3304) );
  AOI21_X1 U14252 ( .B1(n11894), .B2(n11893), .A(n14022), .ZN(n11896) );
  NAND2_X1 U14253 ( .A1(n11896), .A2(n11895), .ZN(n11903) );
  OAI22_X1 U14254 ( .A1(n14013), .A2(n11898), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n11897), .ZN(n11901) );
  NOR2_X1 U14255 ( .A1(n13989), .A2(n11899), .ZN(n11900) );
  AOI211_X1 U14256 ( .C1(n14011), .C2(n14034), .A(n11901), .B(n11900), .ZN(
        n11902) );
  OAI211_X1 U14257 ( .C1(n6891), .C2(n13980), .A(n11903), .B(n11902), .ZN(
        P1_U3224) );
  XNOR2_X1 U14258 ( .A(n11917), .B(n12151), .ZN(n11920) );
  XNOR2_X1 U14259 ( .A(n11920), .B(n11926), .ZN(n11910) );
  INV_X1 U14260 ( .A(n11909), .ZN(n11907) );
  INV_X1 U14261 ( .A(n11910), .ZN(n11906) );
  NAND2_X1 U14262 ( .A1(n11907), .A2(n11906), .ZN(n11922) );
  INV_X1 U14263 ( .A(n11922), .ZN(n11908) );
  AOI21_X1 U14264 ( .B1(n11910), .B2(n11909), .A(n11908), .ZN(n11919) );
  NAND2_X1 U14265 ( .A1(n12732), .A2(n11911), .ZN(n11914) );
  AOI21_X1 U14266 ( .B1(n12733), .B2(n12745), .A(n11912), .ZN(n11913) );
  OAI211_X1 U14267 ( .C1(n11915), .C2(n12736), .A(n11914), .B(n11913), .ZN(
        n11916) );
  AOI21_X1 U14268 ( .B1(n11917), .B2(n12739), .A(n11916), .ZN(n11918) );
  OAI21_X1 U14269 ( .B1(n11919), .B2(n12741), .A(n11918), .ZN(P3_U3164) );
  NAND2_X1 U14270 ( .A1(n11920), .A2(n11926), .ZN(n11921) );
  XNOR2_X1 U14271 ( .A(n14669), .B(n12292), .ZN(n12012) );
  XNOR2_X1 U14272 ( .A(n12012), .B(n12017), .ZN(n11923) );
  XNOR2_X1 U14273 ( .A(n12013), .B(n11923), .ZN(n11931) );
  INV_X1 U14274 ( .A(P3_REG3_REG_13__SCAN_IN), .ZN(n11924) );
  NOR2_X1 U14275 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11924), .ZN(n12762) );
  AOI21_X1 U14276 ( .B1(n12733), .B2(n12744), .A(n12762), .ZN(n11925) );
  OAI21_X1 U14277 ( .B1(n11926), .B2(n12736), .A(n11925), .ZN(n11928) );
  NOR2_X1 U14278 ( .A1(n14669), .A2(n12717), .ZN(n11927) );
  AOI211_X1 U14279 ( .C1(n11929), .C2(n12732), .A(n11928), .B(n11927), .ZN(
        n11930) );
  OAI21_X1 U14280 ( .B1(n11931), .B2(n12741), .A(n11930), .ZN(P3_U3174) );
  OAI22_X1 U14281 ( .A1(n11932), .A2(n14326), .B1(n6904), .B2(n14843), .ZN(
        n11934) );
  AOI211_X1 U14282 ( .C1(n11935), .C2(n14848), .A(n11934), .B(n11933), .ZN(
        n11938) );
  NAND2_X1 U14283 ( .A1(n14854), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n11936) );
  OAI21_X1 U14284 ( .B1(n11938), .B2(n14854), .A(n11936), .ZN(P1_U3543) );
  NAND2_X1 U14285 ( .A1(n6786), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n11937) );
  OAI21_X1 U14286 ( .B1(n11938), .B2(n6786), .A(n11937), .ZN(P1_U3504) );
  NAND2_X1 U14287 ( .A1(n11940), .A2(n12311), .ZN(n11943) );
  INV_X1 U14288 ( .A(n12783), .ZN(n11941) );
  AOI22_X1 U14289 ( .A1(n12332), .A2(SI_14_), .B1(n12162), .B2(n11941), .ZN(
        n11942) );
  XNOR2_X1 U14290 ( .A(n14667), .B(n12737), .ZN(n11986) );
  XNOR2_X1 U14291 ( .A(n11987), .B(n11986), .ZN(n14664) );
  NAND2_X1 U14292 ( .A1(n12268), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n11950) );
  NAND2_X1 U14293 ( .A1(n6491), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n11949) );
  OR2_X1 U14294 ( .A1(n11945), .A2(n11944), .ZN(n11946) );
  NAND2_X1 U14295 ( .A1(n11979), .A2(n11946), .ZN(n12731) );
  NAND2_X1 U14296 ( .A1(n10235), .A2(n12731), .ZN(n11948) );
  NAND2_X1 U14297 ( .A1(n10454), .A2(P3_REG0_REG_15__SCAN_IN), .ZN(n11947) );
  OR2_X1 U14298 ( .A1(n14669), .A2(n12017), .ZN(n11951) );
  XNOR2_X1 U14299 ( .A(n11973), .B(n11986), .ZN(n11953) );
  OAI222_X1 U14300 ( .A1(n15197), .A2(n12727), .B1(n15173), .B2(n12017), .C1(
        n15178), .C2(n11953), .ZN(n14665) );
  NAND2_X1 U14301 ( .A1(n14665), .A2(n15211), .ZN(n11958) );
  INV_X1 U14302 ( .A(n12014), .ZN(n11955) );
  OAI22_X1 U14303 ( .A1(n15211), .A2(n6955), .B1(n11955), .B2(n11954), .ZN(
        n11956) );
  AOI21_X1 U14304 ( .B1(n14667), .B2(n12831), .A(n11956), .ZN(n11957) );
  OAI211_X1 U14305 ( .C1(n14664), .C2(n12877), .A(n11958), .B(n11957), .ZN(
        P3_U3219) );
  OR2_X1 U14306 ( .A1(n11964), .A2(n11961), .ZN(n11962) );
  XNOR2_X1 U14307 ( .A(n13572), .B(n11965), .ZN(n13844) );
  AOI21_X1 U14308 ( .B1(n6631), .B2(n11965), .A(n13536), .ZN(n13842) );
  AOI21_X1 U14309 ( .B1(n13569), .B2(n11966), .A(n12605), .ZN(n11967) );
  OR2_X1 U14310 ( .A1(n13569), .A2(n11966), .ZN(n13744) );
  NAND2_X1 U14311 ( .A1(n11967), .A2(n13744), .ZN(n13839) );
  AOI22_X1 U14312 ( .A1(n13566), .A2(n13524), .B1(n13420), .B2(n13434), .ZN(
        n13838) );
  OAI22_X1 U14313 ( .A1(n15005), .A2(n13838), .B1(n12001), .B2(n14996), .ZN(
        n11969) );
  INV_X1 U14314 ( .A(n13569), .ZN(n13840) );
  NOR2_X1 U14315 ( .A1(n13840), .A2(n14968), .ZN(n11968) );
  AOI211_X1 U14316 ( .C1(n15005), .C2(P2_REG2_REG_17__SCAN_IN), .A(n11969), 
        .B(n11968), .ZN(n11970) );
  OAI21_X1 U14317 ( .B1(n14983), .B2(n13839), .A(n11970), .ZN(n11971) );
  AOI21_X1 U14318 ( .B1(n13842), .B2(n14723), .A(n11971), .ZN(n11972) );
  OAI21_X1 U14319 ( .B1(n13755), .B2(n13844), .A(n11972), .ZN(P2_U3248) );
  NAND2_X1 U14320 ( .A1(n14667), .A2(n12744), .ZN(n11974) );
  NAND2_X1 U14321 ( .A1(n11975), .A2(n11974), .ZN(n12838) );
  NAND2_X1 U14322 ( .A1(n11976), .A2(n12311), .ZN(n11978) );
  AOI22_X1 U14323 ( .A1(n12332), .A2(SI_15_), .B1(n12162), .B2(n14623), .ZN(
        n11977) );
  NAND2_X1 U14324 ( .A1(n11978), .A2(n11977), .ZN(n13110) );
  OR2_X1 U14325 ( .A1(n13110), .A2(n12727), .ZN(n12359) );
  NAND2_X1 U14326 ( .A1(n13110), .A2(n12727), .ZN(n12445) );
  NAND2_X1 U14327 ( .A1(n12359), .A2(n12445), .ZN(n12837) );
  XNOR2_X1 U14328 ( .A(n12838), .B(n12441), .ZN(n11985) );
  NAND2_X1 U14329 ( .A1(n12268), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n11984) );
  NAND2_X1 U14330 ( .A1(n6495), .A2(P3_REG1_REG_16__SCAN_IN), .ZN(n11983) );
  NAND2_X1 U14331 ( .A1(n11979), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n11980) );
  NAND2_X1 U14332 ( .A1(n12140), .A2(n11980), .ZN(n13045) );
  NAND2_X1 U14333 ( .A1(n10235), .A2(n13045), .ZN(n11982) );
  NAND2_X1 U14334 ( .A1(n10454), .A2(P3_REG0_REG_16__SCAN_IN), .ZN(n11981) );
  NAND4_X1 U14335 ( .A1(n11984), .A2(n11983), .A3(n11982), .A4(n11981), .ZN(
        n13028) );
  AOI222_X1 U14336 ( .A1(n15200), .A2(n11985), .B1(n13028), .B2(n13040), .C1(
        n12744), .C2(n15194), .ZN(n13113) );
  INV_X1 U14337 ( .A(n11986), .ZN(n12528) );
  NAND2_X1 U14338 ( .A1(n11987), .A2(n12528), .ZN(n11989) );
  NAND2_X1 U14339 ( .A1(n14667), .A2(n12737), .ZN(n11988) );
  XNOR2_X1 U14340 ( .A(n12304), .B(n12441), .ZN(n13111) );
  INV_X1 U14341 ( .A(n13110), .ZN(n11991) );
  AOI22_X1 U14342 ( .A1(n15213), .A2(P3_REG2_REG_15__SCAN_IN), .B1(n15208), 
        .B2(n12731), .ZN(n11990) );
  OAI21_X1 U14343 ( .B1(n11991), .B2(n13047), .A(n11990), .ZN(n11992) );
  AOI21_X1 U14344 ( .B1(n13111), .B2(n13050), .A(n11992), .ZN(n11993) );
  OAI21_X1 U14345 ( .B1(n13113), .B2(n15213), .A(n11993), .ZN(P3_U3218) );
  XNOR2_X1 U14346 ( .A(n13569), .B(n12611), .ZN(n12566) );
  NAND2_X1 U14347 ( .A1(n13567), .A2(n12610), .ZN(n12564) );
  XNOR2_X1 U14348 ( .A(n12566), .B(n12564), .ZN(n11999) );
  INV_X1 U14349 ( .A(n11994), .ZN(n11995) );
  OAI21_X1 U14350 ( .B1(n11999), .B2(n11998), .A(n12568), .ZN(n12000) );
  NAND2_X1 U14351 ( .A1(n12000), .A2(n13391), .ZN(n12006) );
  INV_X1 U14352 ( .A(n12001), .ZN(n12004) );
  OAI22_X1 U14353 ( .A1(n13424), .A2(n13838), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12002), .ZN(n12003) );
  AOI21_X1 U14354 ( .B1(n12004), .B2(n13422), .A(n12003), .ZN(n12005) );
  OAI211_X1 U14355 ( .C1(n13840), .C2(n13415), .A(n12006), .B(n12005), .ZN(
        P2_U3200) );
  INV_X1 U14356 ( .A(n12007), .ZN(n12010) );
  OAI222_X1 U14357 ( .A1(P1_U3086), .A2(n12009), .B1(n14480), .B2(n12010), 
        .C1(n12008), .C2(n14478), .ZN(P1_U3329) );
  OAI222_X1 U14358 ( .A1(P2_U3088), .A2(n12011), .B1(n13870), .B2(n9094), .C1(
        n12010), .C2(n13873), .ZN(P2_U3301) );
  XNOR2_X1 U14359 ( .A(n14667), .B(n12151), .ZN(n12125) );
  XNOR2_X1 U14360 ( .A(n12125), .B(n12744), .ZN(n12123) );
  XNOR2_X1 U14361 ( .A(n12124), .B(n12123), .ZN(n12020) );
  NAND2_X1 U14362 ( .A1(n12732), .A2(n12014), .ZN(n12016) );
  AND2_X1 U14363 ( .A1(P3_U3151), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n12781) );
  AOI21_X1 U14364 ( .B1(n12733), .B2(n13039), .A(n12781), .ZN(n12015) );
  OAI211_X1 U14365 ( .C1(n12017), .C2(n12736), .A(n12016), .B(n12015), .ZN(
        n12018) );
  AOI21_X1 U14366 ( .B1(n14667), .B2(n12739), .A(n12018), .ZN(n12019) );
  OAI21_X1 U14367 ( .B1(n12020), .B2(n12741), .A(n12019), .ZN(P3_U3155) );
  OAI211_X1 U14368 ( .C1(n12023), .C2(n12022), .A(n12021), .B(n13995), .ZN(
        n12030) );
  OAI21_X1 U14369 ( .B1(n14013), .B2(n12025), .A(n12024), .ZN(n12028) );
  NOR2_X1 U14370 ( .A1(n13989), .A2(n12026), .ZN(n12027) );
  AOI211_X1 U14371 ( .C1(n14011), .C2(n14033), .A(n12028), .B(n12027), .ZN(
        n12029) );
  OAI211_X1 U14372 ( .C1(n12031), .C2(n13980), .A(n12030), .B(n12029), .ZN(
        P1_U3234) );
  INV_X1 U14373 ( .A(n14327), .ZN(n12032) );
  AOI211_X1 U14374 ( .C1(n13949), .C2(n12033), .A(n14326), .B(n12032), .ZN(
        n14418) );
  NOR2_X1 U14375 ( .A1(n14307), .A2(n13947), .ZN(n12041) );
  OAI21_X1 U14376 ( .B1(n12035), .B2(n12034), .A(n12042), .ZN(n12037) );
  NAND3_X1 U14377 ( .A1(n12037), .A2(n14324), .A3(n12036), .ZN(n12040) );
  AOI22_X1 U14378 ( .A1(n14029), .A2(n14321), .B1(n14319), .B2(n12038), .ZN(
        n12039) );
  NAND2_X1 U14379 ( .A1(n12040), .A2(n12039), .ZN(n14419) );
  AOI211_X1 U14380 ( .C1(n14418), .C2(n12108), .A(n12041), .B(n14419), .ZN(
        n12046) );
  AOI22_X1 U14381 ( .A1(n13949), .A2(n14346), .B1(n14830), .B2(
        P1_REG2_REG_17__SCAN_IN), .ZN(n12045) );
  XNOR2_X1 U14382 ( .A(n12043), .B(n12042), .ZN(n14420) );
  NAND2_X1 U14383 ( .A1(n14420), .A2(n14277), .ZN(n12044) );
  OAI211_X1 U14384 ( .C1(n12046), .C2(n14830), .A(n12045), .B(n12044), .ZN(
        P1_U3276) );
  INV_X1 U14385 ( .A(n12047), .ZN(n12562) );
  OAI222_X1 U14386 ( .A1(n14478), .A2(n12088), .B1(n14480), .B2(n12562), .C1(
        n14059), .C2(P1_U3086), .ZN(P1_U3328) );
  INV_X1 U14387 ( .A(n12048), .ZN(n12050) );
  NAND2_X1 U14388 ( .A1(n12050), .A2(n12049), .ZN(n12052) );
  INV_X1 U14389 ( .A(n12052), .ZN(n12056) );
  AND2_X1 U14390 ( .A1(n12054), .A2(n12053), .ZN(n12055) );
  NAND2_X1 U14391 ( .A1(n14158), .A2(n9275), .ZN(n12059) );
  NAND2_X1 U14392 ( .A1(n14175), .A2(n12057), .ZN(n12058) );
  NAND2_X1 U14393 ( .A1(n12059), .A2(n12058), .ZN(n12060) );
  XNOR2_X1 U14394 ( .A(n12060), .B(n9295), .ZN(n12062) );
  AOI22_X1 U14395 ( .A1(n14158), .A2(n12061), .B1(n9278), .B2(n14175), .ZN(
        n12063) );
  XNOR2_X1 U14396 ( .A(n12062), .B(n12063), .ZN(n13876) );
  INV_X1 U14397 ( .A(n12062), .ZN(n12064) );
  AOI22_X1 U14398 ( .A1(n14138), .A2(n9275), .B1(n12065), .B2(n14146), .ZN(
        n12069) );
  AOI22_X1 U14399 ( .A1(n14138), .A2(n12066), .B1(n9278), .B2(n14146), .ZN(
        n12067) );
  XNOR2_X1 U14400 ( .A(n12067), .B(n9295), .ZN(n12068) );
  XOR2_X1 U14401 ( .A(n12069), .B(n12068), .Z(n12070) );
  XNOR2_X1 U14402 ( .A(n12071), .B(n12070), .ZN(n12077) );
  AOI22_X1 U14403 ( .A1(n14011), .A2(n14175), .B1(P1_REG3_REG_28__SCAN_IN), 
        .B2(P1_U3086), .ZN(n12073) );
  NAND2_X1 U14404 ( .A1(n14016), .A2(n14137), .ZN(n12072) );
  OAI211_X1 U14405 ( .C1(n12074), .C2(n14013), .A(n12073), .B(n12072), .ZN(
        n12075) );
  AOI21_X1 U14406 ( .B1(n14138), .B2(n14018), .A(n12075), .ZN(n12076) );
  OAI21_X1 U14407 ( .B1(n12077), .B2(n14022), .A(n12076), .ZN(P1_U3220) );
  NAND2_X1 U14408 ( .A1(n12121), .A2(n12078), .ZN(n12080) );
  OAI211_X1 U14409 ( .C1(n13870), .C2(n12278), .A(n12080), .B(n12079), .ZN(
        P2_U3299) );
  NAND2_X1 U14410 ( .A1(n12082), .A2(n14438), .ZN(n12081) );
  NAND2_X1 U14411 ( .A1(n12081), .A2(n14427), .ZN(n12083) );
  INV_X1 U14412 ( .A(n14351), .ZN(n14120) );
  INV_X1 U14413 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n12277) );
  NOR2_X1 U14414 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(n12278), .ZN(n12090) );
  AOI22_X1 U14415 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(n12563), .B1(
        P1_DATAO_REG_27__SCAN_IN), .B2(n12088), .ZN(n12261) );
  OAI22_X1 U14416 ( .A1(n14477), .A2(P1_DATAO_REG_29__SCAN_IN), .B1(n13871), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n12115) );
  INV_X1 U14417 ( .A(n12316), .ZN(n12091) );
  AOI22_X1 U14418 ( .A1(P2_DATAO_REG_30__SCAN_IN), .A2(n13866), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n12627), .ZN(n12317) );
  AOI22_X1 U14419 ( .A1(n12333), .A2(n13320), .B1(n12092), .B2(SI_30_), .ZN(
        n12093) );
  OAI21_X1 U14420 ( .B1(n12094), .B2(P3_U3151), .A(n12093), .ZN(P3_U3265) );
  NAND2_X1 U14421 ( .A1(n12100), .A2(n12095), .ZN(n12096) );
  NAND2_X1 U14422 ( .A1(n12097), .A2(n12096), .ZN(n12098) );
  XOR2_X1 U14423 ( .A(n12098), .B(P1_REG1_REG_19__SCAN_IN), .Z(n12107) );
  INV_X1 U14424 ( .A(n12107), .ZN(n12105) );
  NAND2_X1 U14425 ( .A1(n12100), .A2(n12099), .ZN(n12102) );
  NAND2_X1 U14426 ( .A1(n12102), .A2(n12101), .ZN(n12103) );
  XOR2_X1 U14427 ( .A(P1_REG2_REG_19__SCAN_IN), .B(n12103), .Z(n12106) );
  OAI21_X1 U14428 ( .B1(n12106), .B2(n14807), .A(n14811), .ZN(n12104) );
  AOI21_X1 U14429 ( .B1(n12105), .B2(n14102), .A(n12104), .ZN(n12110) );
  AOI22_X1 U14430 ( .A1(n12107), .A2(n14102), .B1(n14113), .B2(n12106), .ZN(
        n12109) );
  MUX2_X1 U14431 ( .A(n12110), .B(n12109), .S(n12108), .Z(n12113) );
  NOR2_X1 U14432 ( .A1(n12111), .A2(P1_STATE_REG_SCAN_IN), .ZN(n13908) );
  INV_X1 U14433 ( .A(n13908), .ZN(n12112) );
  OAI211_X1 U14434 ( .C1(n12114), .C2(n14815), .A(n12113), .B(n12112), .ZN(
        P1_U3262) );
  INV_X1 U14435 ( .A(n12115), .ZN(n12116) );
  XNOR2_X1 U14436 ( .A(n12117), .B(n12116), .ZN(n12312) );
  INV_X1 U14437 ( .A(n12312), .ZN(n12120) );
  OAI222_X1 U14438 ( .A1(n13333), .A2(n12120), .B1(n12119), .B2(P3_U3151), 
        .C1(n13215), .C2(n13335), .ZN(P3_U3266) );
  INV_X1 U14439 ( .A(n12121), .ZN(n12122) );
  OAI222_X1 U14440 ( .A1(n14478), .A2(n12277), .B1(n14480), .B2(n12122), .C1(
        P1_U3086), .C2(n8291), .ZN(P1_U3327) );
  INV_X1 U14441 ( .A(n12125), .ZN(n12126) );
  XNOR2_X1 U14442 ( .A(n13110), .B(n12292), .ZN(n12728) );
  INV_X1 U14443 ( .A(n12728), .ZN(n12127) );
  NAND2_X1 U14444 ( .A1(n12127), .A2(n12727), .ZN(n12128) );
  NAND2_X1 U14445 ( .A1(n12130), .A2(n12311), .ZN(n12132) );
  AOI22_X1 U14446 ( .A1(n12332), .A2(SI_16_), .B1(n12162), .B2(n14646), .ZN(
        n12131) );
  XNOR2_X1 U14447 ( .A(n13106), .B(n12151), .ZN(n12134) );
  INV_X1 U14448 ( .A(n13028), .ZN(n12681) );
  XNOR2_X1 U14449 ( .A(n12134), .B(n12681), .ZN(n12669) );
  INV_X1 U14450 ( .A(n12669), .ZN(n12133) );
  INV_X1 U14451 ( .A(n12134), .ZN(n12135) );
  NAND2_X1 U14452 ( .A1(n12135), .A2(n13028), .ZN(n12136) );
  NAND2_X1 U14453 ( .A1(n12137), .A2(n12311), .ZN(n12139) );
  AOI22_X1 U14454 ( .A1(SI_17_), .A2(n12332), .B1(n12802), .B2(n12162), .ZN(
        n12138) );
  NAND2_X1 U14455 ( .A1(n12139), .A2(n12138), .ZN(n13102) );
  XNOR2_X1 U14456 ( .A(n13102), .B(n12292), .ZN(n12146) );
  NAND2_X1 U14457 ( .A1(n12268), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n12145) );
  NAND2_X1 U14458 ( .A1(n10454), .A2(P3_REG0_REG_17__SCAN_IN), .ZN(n12144) );
  NAND2_X1 U14459 ( .A1(n12140), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n12141) );
  NAND2_X1 U14460 ( .A1(n12152), .A2(n12141), .ZN(n13033) );
  NAND2_X1 U14461 ( .A1(n13033), .A2(n10235), .ZN(n12143) );
  NAND2_X1 U14462 ( .A1(n6491), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n12142) );
  XNOR2_X1 U14463 ( .A(n12146), .B(n13014), .ZN(n12678) );
  INV_X1 U14464 ( .A(n13014), .ZN(n13041) );
  NAND2_X1 U14465 ( .A1(n12146), .A2(n13041), .ZN(n12147) );
  NAND2_X1 U14466 ( .A1(n12677), .A2(n12147), .ZN(n12712) );
  NAND2_X1 U14467 ( .A1(n12148), .A2(n12311), .ZN(n12150) );
  AOI22_X1 U14468 ( .A1(n12332), .A2(SI_18_), .B1(n12162), .B2(n12820), .ZN(
        n12149) );
  NAND2_X1 U14469 ( .A1(n12150), .A2(n12149), .ZN(n13098) );
  XNOR2_X1 U14470 ( .A(n13098), .B(n12151), .ZN(n12159) );
  INV_X1 U14471 ( .A(n12168), .ZN(n12154) );
  NAND2_X1 U14472 ( .A1(n12152), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n12153) );
  NAND2_X1 U14473 ( .A1(n12154), .A2(n12153), .ZN(n13022) );
  NAND2_X1 U14474 ( .A1(n13022), .A2(n10235), .ZN(n12158) );
  AOI22_X1 U14475 ( .A1(n12268), .A2(P3_REG2_REG_18__SCAN_IN), .B1(n6495), 
        .B2(P3_REG1_REG_18__SCAN_IN), .ZN(n12157) );
  NAND2_X1 U14476 ( .A1(n10454), .A2(P3_REG0_REG_18__SCAN_IN), .ZN(n12156) );
  XNOR2_X1 U14477 ( .A(n12159), .B(n13029), .ZN(n12711) );
  NAND2_X1 U14478 ( .A1(n12712), .A2(n12711), .ZN(n12710) );
  INV_X1 U14479 ( .A(n12159), .ZN(n12160) );
  NAND2_X1 U14480 ( .A1(n12160), .A2(n13029), .ZN(n12161) );
  NAND2_X1 U14481 ( .A1(n12710), .A2(n12161), .ZN(n12645) );
  AOI22_X1 U14482 ( .A1(n12332), .A2(n12163), .B1(n12162), .B2(n12345), .ZN(
        n12164) );
  XNOR2_X1 U14483 ( .A(n13097), .B(n12151), .ZN(n12173) );
  NOR2_X1 U14484 ( .A1(n12168), .A2(n12167), .ZN(n12169) );
  OR2_X1 U14485 ( .A1(n12179), .A2(n12169), .ZN(n13006) );
  NAND2_X1 U14486 ( .A1(n13006), .A2(n10235), .ZN(n12172) );
  AOI22_X1 U14487 ( .A1(n12268), .A2(P3_REG2_REG_19__SCAN_IN), .B1(n6491), 
        .B2(P3_REG1_REG_19__SCAN_IN), .ZN(n12171) );
  NAND2_X1 U14488 ( .A1(n10454), .A2(P3_REG0_REG_19__SCAN_IN), .ZN(n12170) );
  XNOR2_X1 U14489 ( .A(n12173), .B(n13015), .ZN(n12644) );
  NAND2_X1 U14490 ( .A1(n12173), .A2(n12987), .ZN(n12174) );
  NAND2_X1 U14491 ( .A1(n12643), .A2(n12174), .ZN(n12698) );
  NAND2_X1 U14492 ( .A1(n12175), .A2(n12311), .ZN(n12177) );
  NAND2_X1 U14493 ( .A1(n12332), .A2(SI_20_), .ZN(n12176) );
  XNOR2_X1 U14494 ( .A(n13090), .B(n12151), .ZN(n12187) );
  OR2_X1 U14495 ( .A1(n12179), .A2(n12178), .ZN(n12180) );
  NAND2_X1 U14496 ( .A1(n12193), .A2(n12180), .ZN(n12994) );
  NAND2_X1 U14497 ( .A1(n12994), .A2(n10235), .ZN(n12186) );
  INV_X1 U14498 ( .A(P3_REG2_REG_20__SCAN_IN), .ZN(n12183) );
  NAND2_X1 U14499 ( .A1(n6491), .A2(P3_REG1_REG_20__SCAN_IN), .ZN(n12182) );
  NAND2_X1 U14500 ( .A1(n10454), .A2(P3_REG0_REG_20__SCAN_IN), .ZN(n12181) );
  OAI211_X1 U14501 ( .C1(n6487), .C2(n12183), .A(n12182), .B(n12181), .ZN(
        n12184) );
  INV_X1 U14502 ( .A(n12184), .ZN(n12185) );
  XNOR2_X1 U14503 ( .A(n12187), .B(n13000), .ZN(n12697) );
  INV_X1 U14504 ( .A(n12187), .ZN(n12188) );
  NAND2_X1 U14505 ( .A1(n12188), .A2(n13000), .ZN(n12189) );
  NAND2_X1 U14506 ( .A1(n12190), .A2(n12311), .ZN(n12192) );
  NAND2_X1 U14507 ( .A1(n12332), .A2(SI_21_), .ZN(n12191) );
  XNOR2_X1 U14508 ( .A(n13086), .B(n12151), .ZN(n12201) );
  NAND2_X1 U14509 ( .A1(n12193), .A2(P3_REG3_REG_21__SCAN_IN), .ZN(n12194) );
  NAND2_X1 U14510 ( .A1(n12206), .A2(n12194), .ZN(n12981) );
  NAND2_X1 U14511 ( .A1(n12981), .A2(n10235), .ZN(n12200) );
  INV_X1 U14512 ( .A(P3_REG2_REG_21__SCAN_IN), .ZN(n12197) );
  NAND2_X1 U14513 ( .A1(n6491), .A2(P3_REG1_REG_21__SCAN_IN), .ZN(n12196) );
  NAND2_X1 U14514 ( .A1(n10454), .A2(P3_REG0_REG_21__SCAN_IN), .ZN(n12195) );
  OAI211_X1 U14515 ( .C1(n6487), .C2(n12197), .A(n12196), .B(n12195), .ZN(
        n12198) );
  INV_X1 U14516 ( .A(n12198), .ZN(n12199) );
  XNOR2_X1 U14517 ( .A(n12201), .B(n12846), .ZN(n12655) );
  NAND2_X1 U14518 ( .A1(n12201), .A2(n12846), .ZN(n12202) );
  NAND2_X1 U14519 ( .A1(n12203), .A2(n12311), .ZN(n12205) );
  NAND2_X1 U14520 ( .A1(n12332), .A2(SI_22_), .ZN(n12204) );
  XNOR2_X1 U14521 ( .A(n13082), .B(n12292), .ZN(n12215) );
  XNOR2_X2 U14522 ( .A(n12217), .B(n12215), .ZN(n12703) );
  AND2_X1 U14523 ( .A1(n12206), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n12208) );
  OR2_X1 U14524 ( .A1(n12208), .A2(n12207), .ZN(n12971) );
  NAND2_X1 U14525 ( .A1(n12971), .A2(n10235), .ZN(n12214) );
  INV_X1 U14526 ( .A(P3_REG2_REG_22__SCAN_IN), .ZN(n12211) );
  NAND2_X1 U14527 ( .A1(n6495), .A2(P3_REG1_REG_22__SCAN_IN), .ZN(n12210) );
  NAND2_X1 U14528 ( .A1(n10454), .A2(P3_REG0_REG_22__SCAN_IN), .ZN(n12209) );
  OAI211_X1 U14529 ( .C1(n6487), .C2(n12211), .A(n12210), .B(n12209), .ZN(
        n12212) );
  INV_X1 U14530 ( .A(n12212), .ZN(n12213) );
  INV_X1 U14531 ( .A(n12215), .ZN(n12216) );
  AND2_X1 U14532 ( .A1(n12217), .A2(n12216), .ZN(n12218) );
  XOR2_X1 U14533 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n12219), .Z(n12623) );
  AND2_X1 U14534 ( .A1(n12332), .A2(SI_24_), .ZN(n12220) );
  XNOR2_X1 U14535 ( .A(n12946), .B(n12292), .ZN(n12688) );
  OR2_X1 U14536 ( .A1(n12222), .A2(n12221), .ZN(n12223) );
  NAND2_X1 U14537 ( .A1(n12241), .A2(n12223), .ZN(n12944) );
  NAND2_X1 U14538 ( .A1(n12944), .A2(n10235), .ZN(n12229) );
  INV_X1 U14539 ( .A(P3_REG2_REG_24__SCAN_IN), .ZN(n12226) );
  NAND2_X1 U14540 ( .A1(n6491), .A2(P3_REG1_REG_24__SCAN_IN), .ZN(n12225) );
  NAND2_X1 U14541 ( .A1(n10454), .A2(P3_REG0_REG_24__SCAN_IN), .ZN(n12224) );
  OAI211_X1 U14542 ( .C1(n6487), .C2(n12226), .A(n12225), .B(n12224), .ZN(
        n12227) );
  INV_X1 U14543 ( .A(n12227), .ZN(n12228) );
  NAND2_X1 U14544 ( .A1(n12230), .A2(n12311), .ZN(n12232) );
  NAND2_X1 U14545 ( .A1(n12332), .A2(SI_23_), .ZN(n12231) );
  XNOR2_X1 U14546 ( .A(n12960), .B(n12151), .ZN(n12686) );
  INV_X1 U14547 ( .A(n12686), .ZN(n12233) );
  OAI22_X1 U14548 ( .A1(n12688), .A2(n12922), .B1(n12937), .B2(n12233), .ZN(
        n12237) );
  OAI21_X1 U14549 ( .B1(n12686), .B2(n12967), .A(n12954), .ZN(n12235) );
  NOR2_X1 U14550 ( .A1(n12954), .A2(n12967), .ZN(n12234) );
  AOI22_X1 U14551 ( .A1(n12688), .A2(n12235), .B1(n12234), .B2(n12233), .ZN(
        n12236) );
  NAND2_X1 U14552 ( .A1(n12238), .A2(n12311), .ZN(n12240) );
  NAND2_X1 U14553 ( .A1(n12282), .A2(SI_25_), .ZN(n12239) );
  XNOR2_X1 U14554 ( .A(n13070), .B(n12151), .ZN(n12249) );
  NAND2_X1 U14555 ( .A1(n12241), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n12242) );
  NAND2_X1 U14556 ( .A1(n12253), .A2(n12242), .ZN(n12929) );
  NAND2_X1 U14557 ( .A1(n12929), .A2(n10235), .ZN(n12248) );
  INV_X1 U14558 ( .A(P3_REG2_REG_25__SCAN_IN), .ZN(n12245) );
  NAND2_X1 U14559 ( .A1(n6495), .A2(P3_REG1_REG_25__SCAN_IN), .ZN(n12244) );
  NAND2_X1 U14560 ( .A1(n10454), .A2(P3_REG0_REG_25__SCAN_IN), .ZN(n12243) );
  OAI211_X1 U14561 ( .C1(n6487), .C2(n12245), .A(n12244), .B(n12243), .ZN(
        n12246) );
  INV_X1 U14562 ( .A(n12246), .ZN(n12247) );
  XNOR2_X1 U14563 ( .A(n12249), .B(n12909), .ZN(n12663) );
  INV_X1 U14564 ( .A(n12909), .ZN(n12938) );
  NAND2_X1 U14565 ( .A1(n12250), .A2(n10449), .ZN(n12252) );
  NAND2_X1 U14566 ( .A1(n12332), .A2(SI_26_), .ZN(n12251) );
  XNOR2_X1 U14567 ( .A(n12918), .B(n12151), .ZN(n12260) );
  NAND2_X1 U14568 ( .A1(n12253), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n12254) );
  NAND2_X1 U14569 ( .A1(n12266), .A2(n12254), .ZN(n12916) );
  NAND2_X1 U14570 ( .A1(n12916), .A2(n10235), .ZN(n12259) );
  INV_X1 U14571 ( .A(P3_REG2_REG_26__SCAN_IN), .ZN(n12914) );
  NAND2_X1 U14572 ( .A1(n6491), .A2(P3_REG1_REG_26__SCAN_IN), .ZN(n12256) );
  NAND2_X1 U14573 ( .A1(n10454), .A2(P3_REG0_REG_26__SCAN_IN), .ZN(n12255) );
  OAI211_X1 U14574 ( .C1(n6487), .C2(n12914), .A(n12256), .B(n12255), .ZN(
        n12257) );
  INV_X1 U14575 ( .A(n12257), .ZN(n12258) );
  XNOR2_X1 U14576 ( .A(n12260), .B(n12858), .ZN(n12719) );
  INV_X1 U14577 ( .A(n12261), .ZN(n12262) );
  XNOR2_X1 U14578 ( .A(n12263), .B(n12262), .ZN(n13331) );
  NAND2_X1 U14579 ( .A1(n13331), .A2(n10449), .ZN(n12265) );
  NAND2_X1 U14580 ( .A1(n12282), .A2(SI_27_), .ZN(n12264) );
  XNOR2_X1 U14581 ( .A(n13062), .B(n12151), .ZN(n12276) );
  NAND2_X1 U14582 ( .A1(n12266), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n12267) );
  NAND2_X1 U14583 ( .A1(n12285), .A2(n12267), .ZN(n12903) );
  NAND2_X1 U14584 ( .A1(n12903), .A2(n10235), .ZN(n12274) );
  INV_X1 U14585 ( .A(P3_REG1_REG_27__SCAN_IN), .ZN(n12271) );
  NAND2_X1 U14586 ( .A1(n10454), .A2(P3_REG0_REG_27__SCAN_IN), .ZN(n12270) );
  NAND2_X1 U14587 ( .A1(n12268), .A2(P3_REG2_REG_27__SCAN_IN), .ZN(n12269) );
  OAI211_X1 U14588 ( .C1(n12290), .C2(n12271), .A(n12270), .B(n12269), .ZN(
        n12272) );
  INV_X1 U14589 ( .A(n12272), .ZN(n12273) );
  XNOR2_X1 U14590 ( .A(n12276), .B(n12880), .ZN(n12629) );
  INV_X1 U14591 ( .A(n12629), .ZN(n12275) );
  INV_X1 U14592 ( .A(n12276), .ZN(n12296) );
  AOI22_X1 U14593 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(n12278), .B1(
        P1_DATAO_REG_28__SCAN_IN), .B2(n12277), .ZN(n12279) );
  INV_X1 U14594 ( .A(n12279), .ZN(n12280) );
  XNOR2_X1 U14595 ( .A(n12281), .B(n12280), .ZN(n13328) );
  NAND2_X1 U14596 ( .A1(n13328), .A2(n10449), .ZN(n12284) );
  NAND2_X1 U14597 ( .A1(n12282), .A2(SI_28_), .ZN(n12283) );
  NAND2_X1 U14598 ( .A1(n12284), .A2(n12283), .ZN(n12836) );
  NAND2_X1 U14599 ( .A1(n12285), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n12286) );
  NAND2_X1 U14600 ( .A1(n12827), .A2(n12286), .ZN(n12888) );
  INV_X1 U14601 ( .A(P3_REG1_REG_28__SCAN_IN), .ZN(n12289) );
  NAND2_X1 U14602 ( .A1(n10454), .A2(P3_REG0_REG_28__SCAN_IN), .ZN(n12288) );
  NAND2_X1 U14603 ( .A1(n12268), .A2(P3_REG2_REG_28__SCAN_IN), .ZN(n12287) );
  OAI211_X1 U14604 ( .C1(n12290), .C2(n12289), .A(n12288), .B(n12287), .ZN(
        n12291) );
  OR2_X1 U14605 ( .A1(n12836), .A2(n12894), .ZN(n12495) );
  NAND2_X1 U14606 ( .A1(n12836), .A2(n12894), .ZN(n12497) );
  XNOR2_X1 U14607 ( .A(n12862), .B(n12292), .ZN(n12293) );
  INV_X1 U14608 ( .A(n12293), .ZN(n12297) );
  OAI211_X1 U14609 ( .C1(n12296), .C2(n12910), .A(n12297), .B(n12709), .ZN(
        n12302) );
  NAND3_X1 U14610 ( .A1(n12303), .A2(n12709), .A3(n12293), .ZN(n12301) );
  AOI22_X1 U14611 ( .A1(n12910), .A2(n12720), .B1(P3_REG3_REG_28__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12295) );
  NAND2_X1 U14612 ( .A1(n12888), .A2(n12732), .ZN(n12294) );
  OAI211_X1 U14613 ( .C1(n12881), .C2(n12723), .A(n12295), .B(n12294), .ZN(
        n12299) );
  NOR4_X1 U14614 ( .A1(n12297), .A2(n12296), .A3(n12910), .A4(n12741), .ZN(
        n12298) );
  AOI211_X1 U14615 ( .C1(n12739), .C2(n12836), .A(n12299), .B(n12298), .ZN(
        n12300) );
  OAI211_X1 U14616 ( .C1(n12303), .C2(n12302), .A(n12301), .B(n12300), .ZN(
        P3_U3160) );
  AND2_X1 U14617 ( .A1(n13066), .A2(n12923), .ZN(n12348) );
  XNOR2_X1 U14618 ( .A(n13106), .B(n13028), .ZN(n13043) );
  NAND2_X1 U14619 ( .A1(n13106), .A2(n12681), .ZN(n12446) );
  NAND2_X1 U14620 ( .A1(n12305), .A2(n12446), .ZN(n13032) );
  OR2_X1 U14621 ( .A1(n13102), .A2(n13014), .ZN(n12355) );
  NAND2_X1 U14622 ( .A1(n13102), .A2(n13014), .ZN(n12358) );
  OR2_X1 U14623 ( .A1(n13098), .A2(n12648), .ZN(n13002) );
  NAND2_X1 U14624 ( .A1(n13098), .A2(n12648), .ZN(n12451) );
  XNOR2_X1 U14625 ( .A(n13097), .B(n13015), .ZN(n13004) );
  AND2_X1 U14626 ( .A1(n13004), .A2(n13002), .ZN(n12306) );
  OR2_X1 U14627 ( .A1(n13097), .A2(n12987), .ZN(n12457) );
  NAND2_X1 U14628 ( .A1(n13090), .A2(n12658), .ZN(n12353) );
  NAND2_X1 U14629 ( .A1(n12354), .A2(n12353), .ZN(n12993) );
  NAND2_X1 U14630 ( .A1(n13086), .A2(n12846), .ZN(n12351) );
  OR2_X1 U14631 ( .A1(n13086), .A2(n12846), .ZN(n12352) );
  NAND2_X1 U14632 ( .A1(n12307), .A2(n12352), .ZN(n12970) );
  NAND2_X1 U14633 ( .A1(n13082), .A2(n12636), .ZN(n12464) );
  NAND2_X1 U14634 ( .A1(n12970), .A2(n12464), .ZN(n12308) );
  NAND2_X1 U14635 ( .A1(n12308), .A2(n12465), .ZN(n12951) );
  NAND2_X1 U14636 ( .A1(n12960), .A2(n12967), .ZN(n12934) );
  NAND2_X1 U14637 ( .A1(n13078), .A2(n12937), .ZN(n12309) );
  NAND2_X1 U14638 ( .A1(n12934), .A2(n12309), .ZN(n12852) );
  NAND2_X1 U14639 ( .A1(n12946), .A2(n12954), .ZN(n12471) );
  NAND2_X1 U14640 ( .A1(n13074), .A2(n12922), .ZN(n12473) );
  AND2_X1 U14641 ( .A1(n12939), .A2(n12934), .ZN(n12310) );
  NAND2_X1 U14642 ( .A1(n12953), .A2(n12310), .ZN(n12935) );
  NAND2_X1 U14643 ( .A1(n12935), .A2(n12473), .ZN(n12928) );
  XNOR2_X1 U14644 ( .A(n13070), .B(n12909), .ZN(n12927) );
  NAND2_X1 U14645 ( .A1(n13070), .A2(n12938), .ZN(n12480) );
  OR2_X1 U14646 ( .A1(n13062), .A2(n12880), .ZN(n12491) );
  NAND2_X1 U14647 ( .A1(n13062), .A2(n12880), .ZN(n12493) );
  NAND2_X1 U14648 ( .A1(n12887), .A2(n12886), .ZN(n12885) );
  NAND2_X1 U14649 ( .A1(n12312), .A2(n12311), .ZN(n12315) );
  OR2_X1 U14650 ( .A1(n12313), .A2(n13215), .ZN(n12314) );
  NAND2_X1 U14651 ( .A1(n12315), .A2(n12314), .ZN(n12872) );
  NAND2_X1 U14652 ( .A1(n12834), .A2(n12508), .ZN(n12340) );
  AOI22_X1 U14653 ( .A1(P1_DATAO_REG_31__SCAN_IN), .A2(n12318), .B1(
        P2_DATAO_REG_31__SCAN_IN), .B2(n13862), .ZN(n12319) );
  AND2_X1 U14654 ( .A1(n12332), .A2(SI_31_), .ZN(n12320) );
  INV_X1 U14655 ( .A(P3_REG2_REG_31__SCAN_IN), .ZN(n12323) );
  NAND2_X1 U14656 ( .A1(n6491), .A2(P3_REG1_REG_31__SCAN_IN), .ZN(n12322) );
  NAND2_X1 U14657 ( .A1(n10454), .A2(P3_REG0_REG_31__SCAN_IN), .ZN(n12321) );
  OAI211_X1 U14658 ( .C1(n6487), .C2(n12323), .A(n12322), .B(n12321), .ZN(
        n12324) );
  INV_X1 U14659 ( .A(n12324), .ZN(n12325) );
  NAND2_X1 U14660 ( .A1(n12331), .A2(n12325), .ZN(n12826) );
  NAND2_X1 U14661 ( .A1(n14658), .A2(n12826), .ZN(n12501) );
  INV_X1 U14662 ( .A(P3_REG2_REG_30__SCAN_IN), .ZN(n12833) );
  NAND2_X1 U14663 ( .A1(n6491), .A2(P3_REG1_REG_30__SCAN_IN), .ZN(n12327) );
  NAND2_X1 U14664 ( .A1(n10454), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n12326) );
  OAI211_X1 U14665 ( .C1(n6487), .C2(n12833), .A(n12327), .B(n12326), .ZN(
        n12329) );
  INV_X1 U14666 ( .A(n12329), .ZN(n12330) );
  NAND2_X1 U14667 ( .A1(n12331), .A2(n12330), .ZN(n12867) );
  OR2_X1 U14668 ( .A1(n12867), .A2(n14662), .ZN(n12334) );
  NAND2_X1 U14669 ( .A1(n12501), .A2(n12334), .ZN(n12506) );
  NAND2_X1 U14670 ( .A1(n12872), .A2(n12881), .ZN(n12507) );
  INV_X1 U14671 ( .A(n12507), .ZN(n12335) );
  NOR2_X1 U14672 ( .A1(n12506), .A2(n12335), .ZN(n12503) );
  INV_X1 U14673 ( .A(n14658), .ZN(n12342) );
  AND2_X1 U14674 ( .A1(n12867), .A2(n14662), .ZN(n12341) );
  NAND2_X1 U14675 ( .A1(n12500), .A2(n12342), .ZN(n12343) );
  NAND2_X1 U14676 ( .A1(n12344), .A2(n12343), .ZN(n12346) );
  INV_X1 U14677 ( .A(n12347), .ZN(n12544) );
  INV_X1 U14678 ( .A(n12348), .ZN(n12350) );
  MUX2_X1 U14679 ( .A(n12349), .B(n12350), .S(n12481), .Z(n12489) );
  MUX2_X1 U14680 ( .A(n12352), .B(n12351), .S(n11001), .Z(n12463) );
  MUX2_X1 U14681 ( .A(n12354), .B(n12353), .S(n12481), .Z(n12461) );
  XNOR2_X1 U14682 ( .A(n13086), .B(n12988), .ZN(n12980) );
  NAND2_X1 U14683 ( .A1(n13002), .A2(n12355), .ZN(n12356) );
  NAND2_X1 U14684 ( .A1(n12356), .A2(n12451), .ZN(n12357) );
  NAND2_X1 U14685 ( .A1(n13097), .A2(n12987), .ZN(n12456) );
  NAND3_X1 U14686 ( .A1(n12357), .A2(n11001), .A3(n12456), .ZN(n12453) );
  OAI21_X1 U14687 ( .B1(n13106), .B2(n12681), .A(n12359), .ZN(n12360) );
  NAND2_X1 U14688 ( .A1(n12360), .A2(n12481), .ZN(n12444) );
  MUX2_X1 U14689 ( .A(n12362), .B(n12361), .S(n11001), .Z(n12434) );
  NAND2_X1 U14690 ( .A1(n12369), .A2(n12363), .ZN(n12364) );
  NAND2_X1 U14691 ( .A1(n12374), .A2(n12364), .ZN(n12366) );
  NAND3_X1 U14692 ( .A1(n12384), .A2(n12365), .A3(n11001), .ZN(n12379) );
  NAND2_X1 U14693 ( .A1(n12366), .A2(n12379), .ZN(n12373) );
  NAND2_X1 U14694 ( .A1(n12368), .A2(n12367), .ZN(n12372) );
  NAND2_X1 U14695 ( .A1(n12375), .A2(n12369), .ZN(n12370) );
  NAND2_X1 U14696 ( .A1(n12370), .A2(n11001), .ZN(n12371) );
  NAND3_X1 U14697 ( .A1(n12373), .A2(n12372), .A3(n12371), .ZN(n12377) );
  MUX2_X1 U14698 ( .A(n12375), .B(n12374), .S(n11001), .Z(n12376) );
  NAND3_X1 U14699 ( .A1(n12377), .A2(n15177), .A3(n12376), .ZN(n12382) );
  NAND3_X1 U14700 ( .A1(n12383), .A2(n12378), .A3(n12481), .ZN(n12380) );
  NAND2_X1 U14701 ( .A1(n12380), .A2(n12379), .ZN(n12381) );
  NAND2_X1 U14702 ( .A1(n12382), .A2(n12381), .ZN(n12386) );
  MUX2_X1 U14703 ( .A(n12384), .B(n12383), .S(n11001), .Z(n12385) );
  NAND3_X1 U14704 ( .A1(n12386), .A2(n12510), .A3(n12385), .ZN(n12391) );
  MUX2_X1 U14705 ( .A(n12388), .B(n12387), .S(n12481), .Z(n12389) );
  AND2_X1 U14706 ( .A1(n12389), .A2(n12509), .ZN(n12390) );
  NAND2_X1 U14707 ( .A1(n12391), .A2(n12390), .ZN(n12395) );
  NAND3_X1 U14708 ( .A1(n12395), .A2(n12398), .A3(n12392), .ZN(n12393) );
  NAND2_X1 U14709 ( .A1(n12393), .A2(n12396), .ZN(n12401) );
  NAND2_X1 U14710 ( .A1(n12395), .A2(n12394), .ZN(n12399) );
  INV_X1 U14711 ( .A(n12396), .ZN(n12397) );
  AOI21_X1 U14712 ( .B1(n12399), .B2(n12398), .A(n12397), .ZN(n12400) );
  MUX2_X1 U14713 ( .A(n12401), .B(n12400), .S(n11001), .Z(n12406) );
  MUX2_X1 U14714 ( .A(n12403), .B(n12402), .S(n11001), .Z(n12404) );
  OAI211_X1 U14715 ( .C1(n12406), .C2(n12405), .A(n12404), .B(n12518), .ZN(
        n12410) );
  MUX2_X1 U14716 ( .A(n12408), .B(n12407), .S(n12481), .Z(n12409) );
  NAND3_X1 U14717 ( .A1(n12410), .A2(n12520), .A3(n12409), .ZN(n12417) );
  NAND2_X1 U14718 ( .A1(n12411), .A2(n12481), .ZN(n12415) );
  NAND2_X1 U14719 ( .A1(n12412), .A2(n11001), .ZN(n12414) );
  MUX2_X1 U14720 ( .A(n12415), .B(n12414), .S(n12413), .Z(n12416) );
  NAND2_X1 U14721 ( .A1(n12417), .A2(n12416), .ZN(n12423) );
  MUX2_X1 U14722 ( .A(n12419), .B(n12418), .S(n11001), .Z(n12420) );
  NAND2_X1 U14723 ( .A1(n12421), .A2(n12420), .ZN(n12422) );
  AOI21_X1 U14724 ( .B1(n12423), .B2(n12519), .A(n12422), .ZN(n12432) );
  NAND2_X1 U14725 ( .A1(n12429), .A2(n12424), .ZN(n12427) );
  NAND2_X1 U14726 ( .A1(n12428), .A2(n12425), .ZN(n12426) );
  MUX2_X1 U14727 ( .A(n12427), .B(n12426), .S(n12481), .Z(n12431) );
  MUX2_X1 U14728 ( .A(n12429), .B(n12428), .S(n11001), .Z(n12430) );
  OAI211_X1 U14729 ( .C1(n12432), .C2(n12431), .A(n12526), .B(n12430), .ZN(
        n12433) );
  NAND3_X1 U14730 ( .A1(n12528), .A2(n12434), .A3(n12433), .ZN(n12439) );
  NOR2_X1 U14731 ( .A1(n14667), .A2(n11001), .ZN(n12436) );
  AND2_X1 U14732 ( .A1(n14667), .A2(n11001), .ZN(n12435) );
  MUX2_X1 U14733 ( .A(n12436), .B(n12435), .S(n12737), .Z(n12437) );
  INV_X1 U14734 ( .A(n12437), .ZN(n12438) );
  NAND2_X1 U14735 ( .A1(n12439), .A2(n12438), .ZN(n12440) );
  NAND2_X1 U14736 ( .A1(n12441), .A2(n12440), .ZN(n12443) );
  INV_X1 U14737 ( .A(n12446), .ZN(n12442) );
  AOI21_X1 U14738 ( .B1(n12444), .B2(n12443), .A(n12442), .ZN(n12449) );
  AOI21_X1 U14739 ( .B1(n12446), .B2(n12445), .A(n12481), .ZN(n12448) );
  NAND2_X1 U14740 ( .A1(n13028), .A2(n11001), .ZN(n12447) );
  OAI22_X1 U14741 ( .A1(n12449), .A2(n12448), .B1(n13106), .B2(n12447), .ZN(
        n12450) );
  AOI22_X1 U14742 ( .A1(n12453), .A2(n7029), .B1(n13031), .B2(n12450), .ZN(
        n12455) );
  NAND3_X1 U14743 ( .A1(n12457), .A2(n12481), .A3(n12451), .ZN(n12452) );
  NAND2_X1 U14744 ( .A1(n12453), .A2(n12452), .ZN(n12454) );
  OAI21_X1 U14745 ( .B1(n12455), .B2(n13018), .A(n12454), .ZN(n12459) );
  MUX2_X1 U14746 ( .A(n12457), .B(n12456), .S(n12481), .Z(n12458) );
  NAND3_X1 U14747 ( .A1(n12459), .A2(n7027), .A3(n12458), .ZN(n12460) );
  NAND3_X1 U14748 ( .A1(n12461), .A2(n12980), .A3(n12460), .ZN(n12462) );
  AND2_X1 U14749 ( .A1(n12463), .A2(n12462), .ZN(n12467) );
  NAND2_X1 U14750 ( .A1(n12465), .A2(n12464), .ZN(n12969) );
  MUX2_X1 U14751 ( .A(n12465), .B(n12464), .S(n11001), .Z(n12466) );
  OAI21_X1 U14752 ( .B1(n12467), .B2(n12969), .A(n12466), .ZN(n12469) );
  NOR2_X1 U14753 ( .A1(n12967), .A2(n12481), .ZN(n12468) );
  AOI22_X1 U14754 ( .A1(n12469), .A2(n12950), .B1(n12468), .B2(n13078), .ZN(
        n12479) );
  INV_X1 U14755 ( .A(n12939), .ZN(n12478) );
  INV_X1 U14756 ( .A(n12934), .ZN(n12470) );
  NAND2_X1 U14757 ( .A1(n12473), .A2(n12470), .ZN(n12472) );
  NAND2_X1 U14758 ( .A1(n12472), .A2(n12471), .ZN(n12475) );
  INV_X1 U14759 ( .A(n12473), .ZN(n12474) );
  MUX2_X1 U14760 ( .A(n12475), .B(n12474), .S(n11001), .Z(n12476) );
  INV_X1 U14761 ( .A(n12476), .ZN(n12477) );
  OAI211_X1 U14762 ( .C1(n12479), .C2(n12478), .A(n12927), .B(n12477), .ZN(
        n12486) );
  NOR2_X1 U14763 ( .A1(n13070), .A2(n12938), .ZN(n12483) );
  INV_X1 U14764 ( .A(n12480), .ZN(n12482) );
  MUX2_X1 U14765 ( .A(n12483), .B(n12482), .S(n12481), .Z(n12484) );
  INV_X1 U14766 ( .A(n12484), .ZN(n12485) );
  NAND2_X1 U14767 ( .A1(n12486), .A2(n12485), .ZN(n12487) );
  NAND2_X1 U14768 ( .A1(n12913), .A2(n12487), .ZN(n12488) );
  NAND3_X1 U14769 ( .A1(n12489), .A2(n12897), .A3(n12488), .ZN(n12490) );
  OAI21_X1 U14770 ( .B1(n11001), .B2(n12491), .A(n12490), .ZN(n12492) );
  NAND2_X1 U14771 ( .A1(n12887), .A2(n12492), .ZN(n12499) );
  NAND2_X1 U14772 ( .A1(n12493), .A2(n11001), .ZN(n12494) );
  NAND2_X1 U14773 ( .A1(n12495), .A2(n12494), .ZN(n12496) );
  NAND3_X1 U14774 ( .A1(n12499), .A2(n12497), .A3(n12496), .ZN(n12498) );
  OAI211_X1 U14775 ( .C1(n12499), .C2(n11001), .A(n12498), .B(n12508), .ZN(
        n12502) );
  AOI22_X1 U14776 ( .A1(n12503), .A2(n12502), .B1(n12501), .B2(n12500), .ZN(
        n12504) );
  INV_X1 U14777 ( .A(n12506), .ZN(n12538) );
  INV_X1 U14778 ( .A(n12980), .ZN(n12532) );
  INV_X1 U14779 ( .A(n13004), .ZN(n12531) );
  NAND4_X1 U14780 ( .A1(n12511), .A2(n12510), .A3(n15177), .A4(n12509), .ZN(
        n12517) );
  INV_X1 U14781 ( .A(n15202), .ZN(n12515) );
  NAND4_X1 U14782 ( .A1(n12515), .A2(n12514), .A3(n12513), .A4(n12512), .ZN(
        n12516) );
  NOR2_X1 U14783 ( .A1(n12517), .A2(n12516), .ZN(n12521) );
  NAND4_X1 U14784 ( .A1(n12521), .A2(n12520), .A3(n12519), .A4(n12518), .ZN(
        n12523) );
  NOR2_X1 U14785 ( .A1(n12523), .A2(n12522), .ZN(n12524) );
  NAND3_X1 U14786 ( .A1(n12526), .A2(n12525), .A3(n12524), .ZN(n12527) );
  NOR2_X1 U14787 ( .A1(n12837), .A2(n12527), .ZN(n12529) );
  NAND4_X1 U14788 ( .A1(n13031), .A2(n12529), .A3(n13043), .A4(n12528), .ZN(
        n12530) );
  OR4_X1 U14789 ( .A1(n12532), .A2(n12531), .A3(n13018), .A4(n12530), .ZN(
        n12533) );
  NOR4_X1 U14790 ( .A1(n12852), .A2(n12993), .A3(n12969), .A4(n12533), .ZN(
        n12534) );
  NAND4_X1 U14791 ( .A1(n12927), .A2(n12913), .A3(n12939), .A4(n12534), .ZN(
        n12535) );
  NOR3_X1 U14792 ( .A1(n12862), .A2(n12859), .A3(n12535), .ZN(n12536) );
  NAND4_X1 U14793 ( .A1(n12538), .A2(n12863), .A3(n12537), .A4(n12536), .ZN(
        n12540) );
  XNOR2_X1 U14794 ( .A(n12540), .B(n12539), .ZN(n12542) );
  NOR3_X1 U14795 ( .A1(n13297), .A2(n6485), .A3(n12545), .ZN(n12548) );
  OAI21_X1 U14796 ( .B1(n12549), .B2(n12546), .A(P3_B_REG_SCAN_IN), .ZN(n12547) );
  OAI22_X1 U14797 ( .A1(n12553), .A2(n12552), .B1(n12551), .B2(n14307), .ZN(
        n12554) );
  AOI21_X1 U14798 ( .B1(P1_REG2_REG_29__SCAN_IN), .B2(n14830), .A(n12554), 
        .ZN(n12557) );
  NAND2_X1 U14799 ( .A1(n12555), .A2(n14346), .ZN(n12556) );
  OAI211_X1 U14800 ( .C1(n12558), .C2(n14243), .A(n12557), .B(n12556), .ZN(
        n12559) );
  AOI21_X1 U14801 ( .B1(n12560), .B2(n14277), .A(n12559), .ZN(n12561) );
  OAI21_X1 U14802 ( .B1(n12550), .B2(n14830), .A(n12561), .ZN(P1_U3356) );
  OAI222_X1 U14803 ( .A1(n13870), .A2(n12563), .B1(n13873), .B2(n12562), .C1(
        n13526), .C2(P2_U3088), .ZN(P2_U3300) );
  INV_X1 U14804 ( .A(n12564), .ZN(n12565) );
  XNOR2_X1 U14805 ( .A(n13745), .B(n12611), .ZN(n12570) );
  AND2_X1 U14806 ( .A1(n13566), .A2(n12605), .ZN(n12569) );
  NAND2_X1 U14807 ( .A1(n12570), .A2(n12569), .ZN(n12571) );
  OAI21_X1 U14808 ( .B1(n12570), .B2(n12569), .A(n12571), .ZN(n13408) );
  INV_X1 U14809 ( .A(n12571), .ZN(n12572) );
  XNOR2_X1 U14810 ( .A(n13734), .B(n12611), .ZN(n12575) );
  NAND2_X1 U14811 ( .A1(n13575), .A2(n12610), .ZN(n12573) );
  XNOR2_X1 U14812 ( .A(n12575), .B(n12573), .ZN(n13350) );
  INV_X1 U14813 ( .A(n12573), .ZN(n12574) );
  XNOR2_X1 U14814 ( .A(n13822), .B(n9992), .ZN(n12578) );
  NAND2_X1 U14815 ( .A1(n13361), .A2(n12610), .ZN(n12579) );
  AND2_X1 U14816 ( .A1(n12578), .A2(n12579), .ZN(n13388) );
  INV_X1 U14817 ( .A(n12578), .ZN(n12581) );
  INV_X1 U14818 ( .A(n12579), .ZN(n12580) );
  NAND2_X1 U14819 ( .A1(n12581), .A2(n12580), .ZN(n13387) );
  XNOR2_X1 U14820 ( .A(n13817), .B(n12611), .ZN(n12582) );
  NAND2_X1 U14821 ( .A1(n13433), .A2(n12610), .ZN(n12583) );
  XNOR2_X1 U14822 ( .A(n12582), .B(n12583), .ZN(n13360) );
  INV_X1 U14823 ( .A(n12582), .ZN(n12584) );
  XNOR2_X1 U14824 ( .A(n13811), .B(n12611), .ZN(n12588) );
  XNOR2_X1 U14825 ( .A(n12587), .B(n12588), .ZN(n13399) );
  INV_X1 U14826 ( .A(n13399), .ZN(n12586) );
  NAND2_X1 U14827 ( .A1(n13545), .A2(n12610), .ZN(n13398) );
  NAND2_X1 U14828 ( .A1(n12586), .A2(n12585), .ZN(n13400) );
  INV_X1 U14829 ( .A(n12587), .ZN(n12590) );
  INV_X1 U14830 ( .A(n12588), .ZN(n12589) );
  XNOR2_X1 U14831 ( .A(n13806), .B(n9992), .ZN(n12591) );
  NAND2_X1 U14832 ( .A1(n13580), .A2(n12610), .ZN(n13344) );
  XNOR2_X1 U14833 ( .A(n13795), .B(n12611), .ZN(n12594) );
  AND2_X1 U14834 ( .A1(n13550), .A2(n12605), .ZN(n12593) );
  NAND2_X1 U14835 ( .A1(n12594), .A2(n12593), .ZN(n12596) );
  OAI21_X1 U14836 ( .B1(n12594), .B2(n12593), .A(n12596), .ZN(n13380) );
  INV_X1 U14837 ( .A(n13380), .ZN(n12595) );
  XNOR2_X1 U14838 ( .A(n13791), .B(n9992), .ZN(n12598) );
  NAND2_X1 U14839 ( .A1(n13552), .A2(n12610), .ZN(n12597) );
  NOR2_X1 U14840 ( .A1(n12598), .A2(n12597), .ZN(n12599) );
  AOI21_X1 U14841 ( .B1(n12598), .B2(n12597), .A(n12599), .ZN(n13368) );
  INV_X1 U14842 ( .A(n12599), .ZN(n12600) );
  NAND2_X1 U14843 ( .A1(n13432), .A2(n12610), .ZN(n12602) );
  XNOR2_X1 U14844 ( .A(n13635), .B(n12611), .ZN(n12601) );
  XOR2_X1 U14845 ( .A(n12602), .B(n12601), .Z(n13419) );
  INV_X1 U14846 ( .A(n12601), .ZN(n12603) );
  NAND2_X1 U14847 ( .A1(n12603), .A2(n12602), .ZN(n12604) );
  XNOR2_X1 U14848 ( .A(n13779), .B(n12611), .ZN(n12607) );
  AND2_X1 U14849 ( .A1(n13585), .A2(n12605), .ZN(n12606) );
  NAND2_X1 U14850 ( .A1(n12607), .A2(n12606), .ZN(n12609) );
  OAI21_X1 U14851 ( .B1(n12607), .B2(n12606), .A(n12609), .ZN(n13336) );
  INV_X1 U14852 ( .A(n13336), .ZN(n12608) );
  NAND2_X1 U14853 ( .A1(n13431), .A2(n12610), .ZN(n12612) );
  XNOR2_X1 U14854 ( .A(n12612), .B(n12611), .ZN(n12613) );
  XNOR2_X1 U14855 ( .A(n13769), .B(n12613), .ZN(n12614) );
  NAND2_X1 U14856 ( .A1(n12615), .A2(n13524), .ZN(n12617) );
  NAND2_X1 U14857 ( .A1(n13585), .A2(n13420), .ZN(n12616) );
  NAND2_X1 U14858 ( .A1(n12617), .A2(n12616), .ZN(n13600) );
  OAI22_X1 U14859 ( .A1(n13609), .A2(n13372), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12618), .ZN(n12620) );
  INV_X1 U14860 ( .A(n13769), .ZN(n13607) );
  NOR2_X1 U14861 ( .A1(n13607), .A2(n13415), .ZN(n12619) );
  AOI211_X1 U14862 ( .C1(n13374), .C2(n13600), .A(n12620), .B(n12619), .ZN(
        n12621) );
  OAI21_X1 U14863 ( .B1(n12622), .B2(n13428), .A(n12621), .ZN(P2_U3192) );
  INV_X1 U14864 ( .A(SI_24_), .ZN(n12625) );
  INV_X1 U14865 ( .A(n12623), .ZN(n12624) );
  OAI222_X1 U14866 ( .A1(n9808), .A2(P3_U3151), .B1(n13335), .B2(n12625), .C1(
        n13333), .C2(n12624), .ZN(P3_U3271) );
  INV_X1 U14867 ( .A(n12626), .ZN(n13868) );
  OAI222_X1 U14868 ( .A1(n14480), .A2(n13868), .B1(P1_U3086), .B2(n12628), 
        .C1(n12627), .C2(n14478), .ZN(P1_U3325) );
  XNOR2_X1 U14869 ( .A(n12630), .B(n12629), .ZN(n12635) );
  AOI22_X1 U14870 ( .A1(n12858), .A2(n12720), .B1(P3_REG3_REG_27__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12632) );
  NAND2_X1 U14871 ( .A1(n12903), .A2(n12732), .ZN(n12631) );
  OAI211_X1 U14872 ( .C1(n12894), .C2(n12723), .A(n12632), .B(n12631), .ZN(
        n12633) );
  AOI21_X1 U14873 ( .B1(n13062), .B2(n12739), .A(n12633), .ZN(n12634) );
  OAI21_X1 U14874 ( .B1(n12635), .B2(n12741), .A(n12634), .ZN(P3_U3154) );
  XNOR2_X1 U14875 ( .A(n12685), .B(n12686), .ZN(n12687) );
  XNOR2_X1 U14876 ( .A(n12687), .B(n12937), .ZN(n12642) );
  NOR2_X1 U14877 ( .A1(n12636), .A2(n12736), .ZN(n12639) );
  OAI22_X1 U14878 ( .A1(n12922), .A2(n12723), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12637), .ZN(n12638) );
  AOI211_X1 U14879 ( .C1(n12958), .C2(n12732), .A(n12639), .B(n12638), .ZN(
        n12641) );
  NAND2_X1 U14880 ( .A1(n13078), .A2(n12739), .ZN(n12640) );
  OAI211_X1 U14881 ( .C1(n12642), .C2(n12741), .A(n12641), .B(n12640), .ZN(
        P3_U3156) );
  OAI211_X1 U14882 ( .C1(n12645), .C2(n12644), .A(n12643), .B(n12709), .ZN(
        n12651) );
  AOI21_X1 U14883 ( .B1(n12733), .B2(n13000), .A(n12646), .ZN(n12647) );
  OAI21_X1 U14884 ( .B1(n12648), .B2(n12736), .A(n12647), .ZN(n12649) );
  AOI21_X1 U14885 ( .B1(n13006), .B2(n12732), .A(n12649), .ZN(n12650) );
  OAI211_X1 U14886 ( .C1(n12717), .C2(n13097), .A(n12651), .B(n12650), .ZN(
        P3_U3159) );
  INV_X1 U14887 ( .A(n12652), .ZN(n12653) );
  AOI21_X1 U14888 ( .B1(n12655), .B2(n12654), .A(n12653), .ZN(n12661) );
  AOI22_X1 U14889 ( .A1(n12977), .A2(n12733), .B1(P3_REG3_REG_21__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12657) );
  NAND2_X1 U14890 ( .A1(n12732), .A2(n12981), .ZN(n12656) );
  OAI211_X1 U14891 ( .C1(n12658), .C2(n12736), .A(n12657), .B(n12656), .ZN(
        n12659) );
  AOI21_X1 U14892 ( .B1(n13086), .B2(n12739), .A(n12659), .ZN(n12660) );
  OAI21_X1 U14893 ( .B1(n12661), .B2(n12741), .A(n12660), .ZN(P3_U3163) );
  XOR2_X1 U14894 ( .A(n12663), .B(n12662), .Z(n12668) );
  AOI22_X1 U14895 ( .A1(n12954), .A2(n12720), .B1(P3_REG3_REG_25__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12665) );
  NAND2_X1 U14896 ( .A1(n12929), .A2(n12732), .ZN(n12664) );
  OAI211_X1 U14897 ( .C1(n12923), .C2(n12723), .A(n12665), .B(n12664), .ZN(
        n12666) );
  AOI21_X1 U14898 ( .B1(n13070), .B2(n12739), .A(n12666), .ZN(n12667) );
  OAI21_X1 U14899 ( .B1(n12668), .B2(n12741), .A(n12667), .ZN(P3_U3165) );
  INV_X1 U14900 ( .A(n13106), .ZN(n13048) );
  AOI21_X1 U14901 ( .B1(n12670), .B2(n12669), .A(n12741), .ZN(n12672) );
  NAND2_X1 U14902 ( .A1(n12672), .A2(n12671), .ZN(n12676) );
  NAND2_X1 U14903 ( .A1(n12733), .A2(n13041), .ZN(n12673) );
  NAND2_X1 U14904 ( .A1(P3_U3151), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n14647)
         );
  OAI211_X1 U14905 ( .C1(n12727), .C2(n12736), .A(n12673), .B(n14647), .ZN(
        n12674) );
  AOI21_X1 U14906 ( .B1(n12732), .B2(n13045), .A(n12674), .ZN(n12675) );
  OAI211_X1 U14907 ( .C1(n13048), .C2(n12717), .A(n12676), .B(n12675), .ZN(
        P3_U3166) );
  INV_X1 U14908 ( .A(n13102), .ZN(n13035) );
  OAI211_X1 U14909 ( .C1(n12679), .C2(n12678), .A(n12677), .B(n12709), .ZN(
        n12684) );
  NAND2_X1 U14910 ( .A1(n12733), .A2(n13029), .ZN(n12680) );
  NAND2_X1 U14911 ( .A1(P3_U3151), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n12794)
         );
  OAI211_X1 U14912 ( .C1(n12681), .C2(n12736), .A(n12680), .B(n12794), .ZN(
        n12682) );
  AOI21_X1 U14913 ( .B1(n12732), .B2(n13033), .A(n12682), .ZN(n12683) );
  OAI211_X1 U14914 ( .C1(n13035), .C2(n12717), .A(n12684), .B(n12683), .ZN(
        P3_U3168) );
  OAI22_X1 U14915 ( .A1(n12687), .A2(n12967), .B1(n12686), .B2(n12685), .ZN(
        n12690) );
  XNOR2_X1 U14916 ( .A(n12688), .B(n12922), .ZN(n12689) );
  XNOR2_X1 U14917 ( .A(n12690), .B(n12689), .ZN(n12695) );
  AOI22_X1 U14918 ( .A1(n12967), .A2(n12720), .B1(P3_REG3_REG_24__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12692) );
  NAND2_X1 U14919 ( .A1(n12732), .A2(n12944), .ZN(n12691) );
  OAI211_X1 U14920 ( .C1(n12938), .C2(n12723), .A(n12692), .B(n12691), .ZN(
        n12693) );
  AOI21_X1 U14921 ( .B1(n13074), .B2(n12739), .A(n12693), .ZN(n12694) );
  OAI21_X1 U14922 ( .B1(n12695), .B2(n12741), .A(n12694), .ZN(P3_U3169) );
  INV_X1 U14923 ( .A(n13090), .ZN(n12996) );
  OAI211_X1 U14924 ( .C1(n12698), .C2(n12697), .A(n12696), .B(n12709), .ZN(
        n12702) );
  AOI22_X1 U14925 ( .A1(n12733), .A2(n12988), .B1(P3_REG3_REG_20__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12699) );
  OAI21_X1 U14926 ( .B1(n13015), .B2(n12736), .A(n12699), .ZN(n12700) );
  AOI21_X1 U14927 ( .B1(n12994), .B2(n12732), .A(n12700), .ZN(n12701) );
  OAI211_X1 U14928 ( .C1(n12996), .C2(n12717), .A(n12702), .B(n12701), .ZN(
        P3_U3173) );
  XNOR2_X1 U14929 ( .A(n12703), .B(n12977), .ZN(n12708) );
  AOI22_X1 U14930 ( .A1(n12967), .A2(n12733), .B1(P3_REG3_REG_22__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12705) );
  NAND2_X1 U14931 ( .A1(n12732), .A2(n12971), .ZN(n12704) );
  OAI211_X1 U14932 ( .C1(n12846), .C2(n12736), .A(n12705), .B(n12704), .ZN(
        n12706) );
  AOI21_X1 U14933 ( .B1(n13082), .B2(n12739), .A(n12706), .ZN(n12707) );
  OAI21_X1 U14934 ( .B1(n12708), .B2(n12741), .A(n12707), .ZN(P3_U3175) );
  INV_X1 U14935 ( .A(n13098), .ZN(n13024) );
  OAI211_X1 U14936 ( .C1(n12712), .C2(n12711), .A(n12710), .B(n12709), .ZN(
        n12716) );
  NAND2_X1 U14937 ( .A1(n12733), .A2(n12987), .ZN(n12713) );
  NAND2_X1 U14938 ( .A1(P3_U3151), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n12813)
         );
  OAI211_X1 U14939 ( .C1(n13014), .C2(n12736), .A(n12713), .B(n12813), .ZN(
        n12714) );
  AOI21_X1 U14940 ( .B1(n12732), .B2(n13022), .A(n12714), .ZN(n12715) );
  OAI211_X1 U14941 ( .C1(n13024), .C2(n12717), .A(n12716), .B(n12715), .ZN(
        P3_U3178) );
  XOR2_X1 U14942 ( .A(n12719), .B(n12718), .Z(n12726) );
  AOI22_X1 U14943 ( .A1(n12909), .A2(n12720), .B1(P3_REG3_REG_26__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12722) );
  NAND2_X1 U14944 ( .A1(n12916), .A2(n12732), .ZN(n12721) );
  OAI211_X1 U14945 ( .C1(n12880), .C2(n12723), .A(n12722), .B(n12721), .ZN(
        n12724) );
  AOI21_X1 U14946 ( .B1(n13066), .B2(n12739), .A(n12724), .ZN(n12725) );
  OAI21_X1 U14947 ( .B1(n12726), .B2(n12741), .A(n12725), .ZN(P3_U3180) );
  XNOR2_X1 U14948 ( .A(n12728), .B(n12727), .ZN(n12729) );
  XNOR2_X1 U14949 ( .A(n12730), .B(n12729), .ZN(n12742) );
  NAND2_X1 U14950 ( .A1(n12732), .A2(n12731), .ZN(n12735) );
  AND2_X1 U14951 ( .A1(P3_U3151), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n14635) );
  AOI21_X1 U14952 ( .B1(n12733), .B2(n13028), .A(n14635), .ZN(n12734) );
  OAI211_X1 U14953 ( .C1(n12737), .C2(n12736), .A(n12735), .B(n12734), .ZN(
        n12738) );
  AOI21_X1 U14954 ( .B1(n13110), .B2(n12739), .A(n12738), .ZN(n12740) );
  OAI21_X1 U14955 ( .B1(n12742), .B2(n12741), .A(n12740), .ZN(P3_U3181) );
  MUX2_X1 U14956 ( .A(P3_DATAO_REG_31__SCAN_IN), .B(n12826), .S(P3_U3897), .Z(
        P3_U3522) );
  MUX2_X1 U14957 ( .A(P3_DATAO_REG_30__SCAN_IN), .B(n12867), .S(P3_U3897), .Z(
        P3_U3521) );
  INV_X1 U14958 ( .A(n12894), .ZN(n12868) );
  MUX2_X1 U14959 ( .A(P3_DATAO_REG_28__SCAN_IN), .B(n12868), .S(P3_U3897), .Z(
        P3_U3519) );
  MUX2_X1 U14960 ( .A(n12910), .B(P3_DATAO_REG_27__SCAN_IN), .S(n12743), .Z(
        P3_U3518) );
  MUX2_X1 U14961 ( .A(P3_DATAO_REG_26__SCAN_IN), .B(n12858), .S(P3_U3897), .Z(
        P3_U3517) );
  MUX2_X1 U14962 ( .A(n12909), .B(P3_DATAO_REG_25__SCAN_IN), .S(n12743), .Z(
        P3_U3516) );
  MUX2_X1 U14963 ( .A(n12954), .B(P3_DATAO_REG_24__SCAN_IN), .S(n12743), .Z(
        P3_U3515) );
  MUX2_X1 U14964 ( .A(n12977), .B(P3_DATAO_REG_22__SCAN_IN), .S(n12743), .Z(
        P3_U3513) );
  MUX2_X1 U14965 ( .A(P3_DATAO_REG_21__SCAN_IN), .B(n12988), .S(P3_U3897), .Z(
        P3_U3512) );
  MUX2_X1 U14966 ( .A(P3_DATAO_REG_20__SCAN_IN), .B(n13000), .S(P3_U3897), .Z(
        P3_U3511) );
  MUX2_X1 U14967 ( .A(P3_DATAO_REG_19__SCAN_IN), .B(n12987), .S(P3_U3897), .Z(
        P3_U3510) );
  MUX2_X1 U14968 ( .A(P3_DATAO_REG_18__SCAN_IN), .B(n13029), .S(P3_U3897), .Z(
        P3_U3509) );
  MUX2_X1 U14969 ( .A(P3_DATAO_REG_17__SCAN_IN), .B(n13041), .S(P3_U3897), .Z(
        P3_U3508) );
  MUX2_X1 U14970 ( .A(P3_DATAO_REG_16__SCAN_IN), .B(n13028), .S(P3_U3897), .Z(
        P3_U3507) );
  MUX2_X1 U14971 ( .A(P3_DATAO_REG_15__SCAN_IN), .B(n13039), .S(P3_U3897), .Z(
        P3_U3506) );
  MUX2_X1 U14972 ( .A(P3_DATAO_REG_14__SCAN_IN), .B(n12744), .S(P3_U3897), .Z(
        P3_U3505) );
  MUX2_X1 U14973 ( .A(P3_DATAO_REG_13__SCAN_IN), .B(n12745), .S(P3_U3897), .Z(
        P3_U3504) );
  MUX2_X1 U14974 ( .A(P3_DATAO_REG_12__SCAN_IN), .B(n12746), .S(P3_U3897), .Z(
        P3_U3503) );
  MUX2_X1 U14975 ( .A(P3_DATAO_REG_11__SCAN_IN), .B(n12747), .S(P3_U3897), .Z(
        P3_U3502) );
  MUX2_X1 U14976 ( .A(P3_DATAO_REG_10__SCAN_IN), .B(n12748), .S(P3_U3897), .Z(
        P3_U3501) );
  MUX2_X1 U14977 ( .A(P3_DATAO_REG_8__SCAN_IN), .B(n12749), .S(P3_U3897), .Z(
        P3_U3499) );
  MUX2_X1 U14978 ( .A(P3_DATAO_REG_7__SCAN_IN), .B(n12750), .S(P3_U3897), .Z(
        P3_U3498) );
  MUX2_X1 U14979 ( .A(P3_DATAO_REG_6__SCAN_IN), .B(n12751), .S(P3_U3897), .Z(
        P3_U3497) );
  MUX2_X1 U14980 ( .A(P3_DATAO_REG_5__SCAN_IN), .B(n12752), .S(P3_U3897), .Z(
        P3_U3496) );
  MUX2_X1 U14981 ( .A(P3_DATAO_REG_4__SCAN_IN), .B(n12753), .S(P3_U3897), .Z(
        P3_U3495) );
  MUX2_X1 U14982 ( .A(P3_DATAO_REG_3__SCAN_IN), .B(n12754), .S(P3_U3897), .Z(
        P3_U3494) );
  MUX2_X1 U14983 ( .A(P3_DATAO_REG_2__SCAN_IN), .B(n12755), .S(P3_U3897), .Z(
        P3_U3493) );
  MUX2_X1 U14984 ( .A(P3_DATAO_REG_1__SCAN_IN), .B(n10297), .S(P3_U3897), .Z(
        P3_U3492) );
  MUX2_X1 U14985 ( .A(P3_DATAO_REG_0__SCAN_IN), .B(n15195), .S(P3_U3897), .Z(
        P3_U3491) );
  AOI21_X1 U14986 ( .B1(n12758), .B2(n12757), .A(n12756), .ZN(n12772) );
  OAI21_X1 U14987 ( .B1(n12761), .B2(n12760), .A(n12759), .ZN(n12770) );
  AOI21_X1 U14988 ( .B1(n15097), .B2(P3_ADDR_REG_13__SCAN_IN), .A(n12762), 
        .ZN(n12763) );
  OAI21_X1 U14989 ( .B1(n15139), .B2(n12764), .A(n12763), .ZN(n12769) );
  AOI21_X1 U14990 ( .B1(n14673), .B2(n12766), .A(n12765), .ZN(n12767) );
  NOR2_X1 U14991 ( .A1(n12767), .A2(n15136), .ZN(n12768) );
  AOI211_X1 U14992 ( .C1(n15155), .C2(n12770), .A(n12769), .B(n12768), .ZN(
        n12771) );
  OAI21_X1 U14993 ( .B1(n12772), .B2(n15163), .A(n12771), .ZN(P3_U3195) );
  AOI21_X1 U14994 ( .B1(n12775), .B2(n12774), .A(n12773), .ZN(n12788) );
  XNOR2_X1 U14995 ( .A(n12777), .B(n12776), .ZN(n12786) );
  AOI211_X1 U14996 ( .C1(n12780), .C2(n12779), .A(n15131), .B(n12778), .ZN(
        n12785) );
  AOI21_X1 U14997 ( .B1(n15097), .B2(P3_ADDR_REG_14__SCAN_IN), .A(n12781), 
        .ZN(n12782) );
  OAI21_X1 U14998 ( .B1(n15139), .B2(n12783), .A(n12782), .ZN(n12784) );
  AOI211_X1 U14999 ( .C1(n12786), .C2(n15158), .A(n12785), .B(n12784), .ZN(
        n12787) );
  OAI21_X1 U15000 ( .B1(n12788), .B2(n15163), .A(n12787), .ZN(P3_U3196) );
  INV_X1 U15001 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n12791) );
  INV_X1 U15002 ( .A(n12810), .ZN(n12789) );
  AOI21_X1 U15003 ( .B1(n12791), .B2(n12790), .A(n12789), .ZN(n12804) );
  INV_X1 U15004 ( .A(P3_ADDR_REG_17__SCAN_IN), .ZN(n12796) );
  NOR2_X1 U15005 ( .A1(n12792), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n12793) );
  OAI21_X1 U15006 ( .B1(n12793), .B2(n12815), .A(n15158), .ZN(n12795) );
  OAI211_X1 U15007 ( .C1(n15168), .C2(n12796), .A(n12795), .B(n12794), .ZN(
        n12801) );
  AOI211_X1 U15008 ( .C1(n12799), .C2(n12798), .A(n15131), .B(n12797), .ZN(
        n12800) );
  AOI211_X1 U15009 ( .C1(n15153), .C2(n12802), .A(n12801), .B(n12800), .ZN(
        n12803) );
  OAI21_X1 U15010 ( .B1(n12804), .B2(n15163), .A(n12803), .ZN(P3_U3199) );
  AOI21_X1 U15011 ( .B1(n12807), .B2(n12806), .A(n12805), .ZN(n12823) );
  AND3_X1 U15012 ( .A1(n12810), .A2(n12809), .A3(n12808), .ZN(n12811) );
  OAI21_X1 U15013 ( .B1(n12812), .B2(n12811), .A(n8555), .ZN(n12822) );
  INV_X1 U15014 ( .A(P3_ADDR_REG_18__SCAN_IN), .ZN(n14614) );
  OAI21_X1 U15015 ( .B1(n15168), .B2(n14614), .A(n12813), .ZN(n12819) );
  OR3_X1 U15016 ( .A1(n12815), .A2(n6522), .A3(n12814), .ZN(n12816) );
  AOI21_X1 U15017 ( .B1(n12817), .B2(n12816), .A(n15136), .ZN(n12818) );
  AOI211_X1 U15018 ( .C1(n15153), .C2(n12820), .A(n12819), .B(n12818), .ZN(
        n12821) );
  OAI211_X1 U15019 ( .C1(n12823), .C2(n15131), .A(n12822), .B(n12821), .ZN(
        P3_U3200) );
  INV_X1 U15020 ( .A(P3_B_REG_SCAN_IN), .ZN(n12824) );
  NOR2_X1 U15021 ( .A1(n6485), .A2(n12824), .ZN(n12825) );
  NOR2_X1 U15022 ( .A1(n15197), .A2(n12825), .ZN(n12866) );
  NAND2_X1 U15023 ( .A1(n12826), .A2(n12866), .ZN(n14661) );
  INV_X1 U15024 ( .A(n12827), .ZN(n12828) );
  NAND2_X1 U15025 ( .A1(n12828), .A2(n15208), .ZN(n12871) );
  OAI21_X1 U15026 ( .B1(n15213), .B2(n14661), .A(n12871), .ZN(n12830) );
  AOI21_X1 U15027 ( .B1(n15213), .B2(P3_REG2_REG_31__SCAN_IN), .A(n12830), 
        .ZN(n12829) );
  OAI21_X1 U15028 ( .B1(n14658), .B2(n13047), .A(n12829), .ZN(P3_U3202) );
  AOI21_X1 U15029 ( .B1(n12831), .B2(n12337), .A(n12830), .ZN(n12832) );
  OAI21_X1 U15030 ( .B1(n12833), .B2(n15211), .A(n12832), .ZN(P3_U3203) );
  INV_X1 U15031 ( .A(n12863), .ZN(n12835) );
  INV_X1 U15032 ( .A(n12836), .ZN(n13061) );
  NAND2_X1 U15033 ( .A1(n12838), .A2(n12837), .ZN(n12840) );
  NAND2_X1 U15034 ( .A1(n13110), .A2(n13039), .ZN(n12839) );
  AND2_X1 U15035 ( .A1(n13106), .A2(n13028), .ZN(n12841) );
  OR2_X1 U15036 ( .A1(n13106), .A2(n13028), .ZN(n12842) );
  OR2_X1 U15037 ( .A1(n13098), .A2(n13029), .ZN(n12843) );
  AND2_X1 U15038 ( .A1(n13097), .A2(n13015), .ZN(n12844) );
  NAND2_X1 U15039 ( .A1(n13090), .A2(n13000), .ZN(n12845) );
  INV_X1 U15040 ( .A(n13086), .ZN(n12983) );
  NAND2_X1 U15041 ( .A1(n12983), .A2(n12846), .ZN(n12964) );
  OR2_X1 U15042 ( .A1(n13082), .A2(n12977), .ZN(n12847) );
  AND2_X1 U15043 ( .A1(n12964), .A2(n12847), .ZN(n12848) );
  NAND2_X1 U15044 ( .A1(n12965), .A2(n12848), .ZN(n12850) );
  NAND2_X1 U15045 ( .A1(n13082), .A2(n12977), .ZN(n12849) );
  NOR2_X1 U15046 ( .A1(n12960), .A2(n12937), .ZN(n12851) );
  NAND2_X1 U15047 ( .A1(n13074), .A2(n12954), .ZN(n12853) );
  NAND2_X1 U15048 ( .A1(n12940), .A2(n12853), .ZN(n12855) );
  NAND2_X1 U15049 ( .A1(n12946), .A2(n12922), .ZN(n12854) );
  NAND2_X1 U15050 ( .A1(n12855), .A2(n12854), .ZN(n12921) );
  OR2_X2 U15051 ( .A1(n12921), .A2(n12927), .ZN(n12925) );
  NAND2_X1 U15052 ( .A1(n13070), .A2(n12909), .ZN(n12856) );
  NAND2_X1 U15053 ( .A1(n12918), .A2(n12923), .ZN(n12857) );
  NAND2_X1 U15054 ( .A1(n13066), .A2(n12858), .ZN(n12895) );
  AND2_X1 U15055 ( .A1(n12859), .A2(n12895), .ZN(n12860) );
  INV_X1 U15056 ( .A(n13062), .ZN(n12905) );
  NAND2_X1 U15057 ( .A1(n12905), .A2(n12880), .ZN(n12861) );
  OAI21_X1 U15058 ( .B1(n12894), .B2(n13061), .A(n12883), .ZN(n12864) );
  XNOR2_X1 U15059 ( .A(n12864), .B(n12863), .ZN(n12865) );
  NAND2_X1 U15060 ( .A1(n12865), .A2(n15200), .ZN(n12870) );
  AOI22_X1 U15061 ( .A1(n12868), .A2(n15194), .B1(n12867), .B2(n12866), .ZN(
        n12869) );
  NAND2_X1 U15062 ( .A1(n12870), .A2(n12869), .ZN(n13052) );
  NAND2_X1 U15063 ( .A1(n13052), .A2(n15211), .ZN(n12876) );
  INV_X1 U15064 ( .A(n12871), .ZN(n12874) );
  INV_X1 U15065 ( .A(n12872), .ZN(n13055) );
  NOR2_X1 U15066 ( .A1(n13055), .A2(n13047), .ZN(n12873) );
  AOI211_X1 U15067 ( .C1(n15213), .C2(P3_REG2_REG_29__SCAN_IN), .A(n12874), 
        .B(n12873), .ZN(n12875) );
  OAI211_X1 U15068 ( .C1(n13056), .C2(n12877), .A(n12876), .B(n12875), .ZN(
        P3_U3204) );
  INV_X1 U15069 ( .A(n12878), .ZN(n12879) );
  AOI21_X1 U15070 ( .B1(n12879), .B2(n12887), .A(n15178), .ZN(n12884) );
  OAI22_X1 U15071 ( .A1(n12881), .A2(n15197), .B1(n12880), .B2(n15173), .ZN(
        n12882) );
  AOI21_X1 U15072 ( .B1(n12884), .B2(n12883), .A(n12882), .ZN(n13060) );
  OAI21_X1 U15073 ( .B1(n12887), .B2(n12886), .A(n12885), .ZN(n13058) );
  AOI22_X1 U15074 ( .A1(n12888), .A2(n15208), .B1(P3_REG2_REG_28__SCAN_IN), 
        .B2(n15213), .ZN(n12889) );
  OAI21_X1 U15075 ( .B1(n13061), .B2(n13047), .A(n12889), .ZN(n12890) );
  AOI21_X1 U15076 ( .B1(n13058), .B2(n13050), .A(n12890), .ZN(n12891) );
  OAI21_X1 U15077 ( .B1(n13060), .B2(n15213), .A(n12891), .ZN(P3_U3205) );
  OAI21_X1 U15078 ( .B1(n12897), .B2(n12893), .A(n12892), .ZN(n13063) );
  OAI22_X1 U15079 ( .A1(n12894), .A2(n15197), .B1(n12923), .B2(n15173), .ZN(
        n12902) );
  NAND2_X1 U15080 ( .A1(n12896), .A2(n12895), .ZN(n12898) );
  NAND2_X1 U15081 ( .A1(n12898), .A2(n12897), .ZN(n12899) );
  AOI21_X1 U15082 ( .B1(n12900), .B2(n12899), .A(n15178), .ZN(n12901) );
  AOI22_X1 U15083 ( .A1(n12903), .A2(n15208), .B1(P3_REG2_REG_27__SCAN_IN), 
        .B2(n15213), .ZN(n12904) );
  OAI21_X1 U15084 ( .B1(n12905), .B2(n13047), .A(n12904), .ZN(n12906) );
  AOI21_X1 U15085 ( .B1(n13063), .B2(n15209), .A(n12906), .ZN(n12907) );
  OAI21_X1 U15086 ( .B1(n13065), .B2(n15213), .A(n12907), .ZN(P3_U3206) );
  XNOR2_X1 U15087 ( .A(n12908), .B(n12913), .ZN(n12911) );
  AOI222_X1 U15088 ( .A1(n15200), .A2(n12911), .B1(n12910), .B2(n13040), .C1(
        n12909), .C2(n15194), .ZN(n13069) );
  XNOR2_X1 U15089 ( .A(n12913), .B(n12912), .ZN(n13067) );
  NOR2_X1 U15090 ( .A1(n15211), .A2(n12914), .ZN(n12915) );
  AOI21_X1 U15091 ( .B1(n12916), .B2(n15208), .A(n12915), .ZN(n12917) );
  OAI21_X1 U15092 ( .B1(n12918), .B2(n13047), .A(n12917), .ZN(n12919) );
  AOI21_X1 U15093 ( .B1(n13067), .B2(n13050), .A(n12919), .ZN(n12920) );
  OAI21_X1 U15094 ( .B1(n13069), .B2(n15213), .A(n12920), .ZN(P3_U3207) );
  AOI21_X1 U15095 ( .B1(n12921), .B2(n12927), .A(n15178), .ZN(n12926) );
  OAI22_X1 U15096 ( .A1(n12923), .A2(n15197), .B1(n12922), .B2(n15173), .ZN(
        n12924) );
  AOI21_X1 U15097 ( .B1(n12926), .B2(n12925), .A(n12924), .ZN(n13073) );
  XNOR2_X1 U15098 ( .A(n12928), .B(n12927), .ZN(n13071) );
  INV_X1 U15099 ( .A(n13070), .ZN(n12931) );
  AOI22_X1 U15100 ( .A1(n12929), .A2(n15208), .B1(P3_REG2_REG_25__SCAN_IN), 
        .B2(n15213), .ZN(n12930) );
  OAI21_X1 U15101 ( .B1(n12931), .B2(n13047), .A(n12930), .ZN(n12932) );
  AOI21_X1 U15102 ( .B1(n13071), .B2(n13050), .A(n12932), .ZN(n12933) );
  OAI21_X1 U15103 ( .B1(n13073), .B2(n15213), .A(n12933), .ZN(P3_U3208) );
  AND2_X1 U15104 ( .A1(n12953), .A2(n12934), .ZN(n12936) );
  OAI21_X1 U15105 ( .B1(n12936), .B2(n12939), .A(n12935), .ZN(n13075) );
  OAI22_X1 U15106 ( .A1(n12938), .A2(n15197), .B1(n12937), .B2(n15173), .ZN(
        n12943) );
  XNOR2_X1 U15107 ( .A(n6482), .B(n12939), .ZN(n12941) );
  NOR2_X1 U15108 ( .A1(n12941), .A2(n15178), .ZN(n12942) );
  AOI211_X1 U15109 ( .C1(n15204), .C2(n13075), .A(n12943), .B(n12942), .ZN(
        n13077) );
  AOI22_X1 U15110 ( .A1(n15208), .A2(n12944), .B1(n15213), .B2(
        P3_REG2_REG_24__SCAN_IN), .ZN(n12945) );
  OAI21_X1 U15111 ( .B1(n12946), .B2(n13047), .A(n12945), .ZN(n12947) );
  AOI21_X1 U15112 ( .B1(n13075), .B2(n15209), .A(n12947), .ZN(n12948) );
  OAI21_X1 U15113 ( .B1(n13077), .B2(n15213), .A(n12948), .ZN(P3_U3209) );
  XNOR2_X1 U15114 ( .A(n12949), .B(n12950), .ZN(n12957) );
  OR2_X1 U15115 ( .A1(n12951), .A2(n12950), .ZN(n12952) );
  NAND2_X1 U15116 ( .A1(n12953), .A2(n12952), .ZN(n13081) );
  AOI22_X1 U15117 ( .A1(n12954), .A2(n13040), .B1(n15194), .B2(n12977), .ZN(
        n12955) );
  OAI21_X1 U15118 ( .B1(n13081), .B2(n13054), .A(n12955), .ZN(n12956) );
  AOI21_X1 U15119 ( .B1(n12957), .B2(n15200), .A(n12956), .ZN(n13080) );
  INV_X1 U15120 ( .A(n13081), .ZN(n12962) );
  AOI22_X1 U15121 ( .A1(n15213), .A2(P3_REG2_REG_23__SCAN_IN), .B1(n12958), 
        .B2(n15208), .ZN(n12959) );
  OAI21_X1 U15122 ( .B1(n12960), .B2(n13047), .A(n12959), .ZN(n12961) );
  AOI21_X1 U15123 ( .B1(n12962), .B2(n15209), .A(n12961), .ZN(n12963) );
  OAI21_X1 U15124 ( .B1(n13080), .B2(n15213), .A(n12963), .ZN(P3_U3210) );
  NAND2_X1 U15125 ( .A1(n12965), .A2(n12964), .ZN(n12966) );
  XNOR2_X1 U15126 ( .A(n12966), .B(n12969), .ZN(n12968) );
  AOI222_X1 U15127 ( .A1(n15200), .A2(n12968), .B1(n12967), .B2(n13040), .C1(
        n12988), .C2(n15194), .ZN(n13085) );
  XNOR2_X1 U15128 ( .A(n12970), .B(n12969), .ZN(n13083) );
  INV_X1 U15129 ( .A(n13082), .ZN(n12973) );
  AOI22_X1 U15130 ( .A1(n15213), .A2(P3_REG2_REG_22__SCAN_IN), .B1(n15208), 
        .B2(n12971), .ZN(n12972) );
  OAI21_X1 U15131 ( .B1(n12973), .B2(n13047), .A(n12972), .ZN(n12974) );
  AOI21_X1 U15132 ( .B1(n13083), .B2(n13050), .A(n12974), .ZN(n12975) );
  OAI21_X1 U15133 ( .B1(n13085), .B2(n15213), .A(n12975), .ZN(P3_U3211) );
  XNOR2_X1 U15134 ( .A(n12976), .B(n12980), .ZN(n12978) );
  AOI222_X1 U15135 ( .A1(n15200), .A2(n12978), .B1(n12977), .B2(n13040), .C1(
        n13000), .C2(n15194), .ZN(n13089) );
  XOR2_X1 U15136 ( .A(n12980), .B(n12979), .Z(n13087) );
  AOI22_X1 U15137 ( .A1(n15213), .A2(P3_REG2_REG_21__SCAN_IN), .B1(n15208), 
        .B2(n12981), .ZN(n12982) );
  OAI21_X1 U15138 ( .B1(n12983), .B2(n13047), .A(n12982), .ZN(n12984) );
  AOI21_X1 U15139 ( .B1(n13087), .B2(n13050), .A(n12984), .ZN(n12985) );
  OAI21_X1 U15140 ( .B1(n13089), .B2(n15213), .A(n12985), .ZN(P3_U3212) );
  XNOR2_X1 U15141 ( .A(n12986), .B(n7027), .ZN(n12989) );
  AOI222_X1 U15142 ( .A1(n15200), .A2(n12989), .B1(n12988), .B2(n13040), .C1(
        n12987), .C2(n15194), .ZN(n13093) );
  INV_X1 U15143 ( .A(n12990), .ZN(n12991) );
  AOI21_X1 U15144 ( .B1(n12993), .B2(n12992), .A(n12991), .ZN(n13091) );
  AOI22_X1 U15145 ( .A1(n15213), .A2(P3_REG2_REG_20__SCAN_IN), .B1(n15208), 
        .B2(n12994), .ZN(n12995) );
  OAI21_X1 U15146 ( .B1(n12996), .B2(n13047), .A(n12995), .ZN(n12997) );
  AOI21_X1 U15147 ( .B1(n13091), .B2(n13050), .A(n12997), .ZN(n12998) );
  OAI21_X1 U15148 ( .B1(n13093), .B2(n15213), .A(n12998), .ZN(P3_U3213) );
  XOR2_X1 U15149 ( .A(n13004), .B(n12999), .Z(n13001) );
  AOI222_X1 U15150 ( .A1(n15200), .A2(n13001), .B1(n13000), .B2(n13040), .C1(
        n13029), .C2(n15194), .ZN(n13096) );
  AND2_X1 U15151 ( .A1(n13021), .A2(n13002), .ZN(n13005) );
  OAI21_X1 U15152 ( .B1(n13005), .B2(n13004), .A(n13003), .ZN(n13094) );
  AOI22_X1 U15153 ( .A1(n15213), .A2(P3_REG2_REG_19__SCAN_IN), .B1(n15208), 
        .B2(n13006), .ZN(n13007) );
  OAI21_X1 U15154 ( .B1(n13097), .B2(n13047), .A(n13007), .ZN(n13008) );
  AOI21_X1 U15155 ( .B1(n13094), .B2(n13050), .A(n13008), .ZN(n13009) );
  OAI21_X1 U15156 ( .B1(n13096), .B2(n15213), .A(n13009), .ZN(P3_U3214) );
  NAND2_X1 U15157 ( .A1(n13011), .A2(n13010), .ZN(n13012) );
  NAND2_X1 U15158 ( .A1(n13013), .A2(n13012), .ZN(n13017) );
  OAI22_X1 U15159 ( .A1(n13015), .A2(n15197), .B1(n13014), .B2(n15173), .ZN(
        n13016) );
  AOI21_X1 U15160 ( .B1(n13017), .B2(n15200), .A(n13016), .ZN(n13101) );
  NAND2_X1 U15161 ( .A1(n13019), .A2(n13018), .ZN(n13020) );
  AOI22_X1 U15162 ( .A1(n15213), .A2(P3_REG2_REG_18__SCAN_IN), .B1(n15208), 
        .B2(n13022), .ZN(n13023) );
  OAI21_X1 U15163 ( .B1(n13024), .B2(n13047), .A(n13023), .ZN(n13025) );
  AOI21_X1 U15164 ( .B1(n13099), .B2(n13050), .A(n13025), .ZN(n13026) );
  OAI21_X1 U15165 ( .B1(n13101), .B2(n15213), .A(n13026), .ZN(P3_U3215) );
  XOR2_X1 U15166 ( .A(n13027), .B(n13031), .Z(n13030) );
  AOI222_X1 U15167 ( .A1(n15200), .A2(n13030), .B1(n13029), .B2(n13040), .C1(
        n13028), .C2(n15194), .ZN(n13105) );
  XNOR2_X1 U15168 ( .A(n13032), .B(n13031), .ZN(n13103) );
  AOI22_X1 U15169 ( .A1(n15213), .A2(P3_REG2_REG_17__SCAN_IN), .B1(n15208), 
        .B2(n13033), .ZN(n13034) );
  OAI21_X1 U15170 ( .B1(n13035), .B2(n13047), .A(n13034), .ZN(n13036) );
  AOI21_X1 U15171 ( .B1(n13103), .B2(n13050), .A(n13036), .ZN(n13037) );
  OAI21_X1 U15172 ( .B1(n13105), .B2(n15213), .A(n13037), .ZN(P3_U3216) );
  XNOR2_X1 U15173 ( .A(n13038), .B(n13043), .ZN(n13042) );
  AOI222_X1 U15174 ( .A1(n15200), .A2(n13042), .B1(n13041), .B2(n13040), .C1(
        n13039), .C2(n15194), .ZN(n13109) );
  XNOR2_X1 U15175 ( .A(n13044), .B(n13043), .ZN(n13107) );
  AOI22_X1 U15176 ( .A1(n15213), .A2(P3_REG2_REG_16__SCAN_IN), .B1(n15208), 
        .B2(n13045), .ZN(n13046) );
  OAI21_X1 U15177 ( .B1(n13048), .B2(n13047), .A(n13046), .ZN(n13049) );
  AOI21_X1 U15178 ( .B1(n13107), .B2(n13050), .A(n13049), .ZN(n13051) );
  OAI21_X1 U15179 ( .B1(n13109), .B2(n15213), .A(n13051), .ZN(P3_U3217) );
  INV_X1 U15180 ( .A(n13052), .ZN(n13057) );
  NAND2_X1 U15181 ( .A1(n13053), .A2(n15206), .ZN(n15262) );
  MUX2_X1 U15182 ( .A(P3_REG1_REG_29__SCAN_IN), .B(n13301), .S(n15281), .Z(
        P3_U3488) );
  NAND2_X1 U15183 ( .A1(n13058), .A2(n15214), .ZN(n13059) );
  OAI211_X1 U15184 ( .C1(n13061), .C2(n15261), .A(n13060), .B(n13059), .ZN(
        n13302) );
  MUX2_X1 U15185 ( .A(P3_REG1_REG_28__SCAN_IN), .B(n13302), .S(n15281), .Z(
        P3_U3487) );
  INV_X1 U15186 ( .A(n15262), .ZN(n15257) );
  AOI22_X1 U15187 ( .A1(n13063), .A2(n15257), .B1(n15224), .B2(n13062), .ZN(
        n13064) );
  MUX2_X1 U15188 ( .A(P3_REG1_REG_27__SCAN_IN), .B(n13303), .S(n15281), .Z(
        P3_U3486) );
  AOI22_X1 U15189 ( .A1(n13067), .A2(n15214), .B1(n15224), .B2(n13066), .ZN(
        n13068) );
  NAND2_X1 U15190 ( .A1(n13069), .A2(n13068), .ZN(n13304) );
  MUX2_X1 U15191 ( .A(P3_REG1_REG_26__SCAN_IN), .B(n13304), .S(n15281), .Z(
        P3_U3485) );
  AOI22_X1 U15192 ( .A1(n13071), .A2(n15214), .B1(n15224), .B2(n13070), .ZN(
        n13072) );
  NAND2_X1 U15193 ( .A1(n13073), .A2(n13072), .ZN(n13305) );
  MUX2_X1 U15194 ( .A(P3_REG1_REG_25__SCAN_IN), .B(n13305), .S(n15281), .Z(
        P3_U3484) );
  AOI22_X1 U15195 ( .A1(n13075), .A2(n15257), .B1(n15224), .B2(n13074), .ZN(
        n13076) );
  NAND2_X1 U15196 ( .A1(n13077), .A2(n13076), .ZN(n13306) );
  MUX2_X1 U15197 ( .A(P3_REG1_REG_24__SCAN_IN), .B(n13306), .S(n15281), .Z(
        P3_U3483) );
  NAND2_X1 U15198 ( .A1(n13078), .A2(n15224), .ZN(n13079) );
  OAI211_X1 U15199 ( .C1(n13081), .C2(n15262), .A(n13080), .B(n13079), .ZN(
        n13307) );
  MUX2_X1 U15200 ( .A(P3_REG1_REG_23__SCAN_IN), .B(n13307), .S(n15281), .Z(
        P3_U3482) );
  AOI22_X1 U15201 ( .A1(n13083), .A2(n15214), .B1(n15224), .B2(n13082), .ZN(
        n13084) );
  NAND2_X1 U15202 ( .A1(n13085), .A2(n13084), .ZN(n13308) );
  MUX2_X1 U15203 ( .A(P3_REG1_REG_22__SCAN_IN), .B(n13308), .S(n15281), .Z(
        P3_U3481) );
  AOI22_X1 U15204 ( .A1(n13087), .A2(n15214), .B1(n15224), .B2(n13086), .ZN(
        n13088) );
  NAND2_X1 U15205 ( .A1(n13089), .A2(n13088), .ZN(n13309) );
  MUX2_X1 U15206 ( .A(P3_REG1_REG_21__SCAN_IN), .B(n13309), .S(n15281), .Z(
        P3_U3480) );
  AOI22_X1 U15207 ( .A1(n13091), .A2(n15214), .B1(n15224), .B2(n13090), .ZN(
        n13092) );
  NAND2_X1 U15208 ( .A1(n13093), .A2(n13092), .ZN(n13310) );
  MUX2_X1 U15209 ( .A(P3_REG1_REG_20__SCAN_IN), .B(n13310), .S(n15281), .Z(
        P3_U3479) );
  NAND2_X1 U15210 ( .A1(n13094), .A2(n15214), .ZN(n13095) );
  OAI211_X1 U15211 ( .C1(n13097), .C2(n15261), .A(n13096), .B(n13095), .ZN(
        n13311) );
  MUX2_X1 U15212 ( .A(P3_REG1_REG_19__SCAN_IN), .B(n13311), .S(n15281), .Z(
        P3_U3478) );
  AOI22_X1 U15213 ( .A1(n13099), .A2(n15214), .B1(n15224), .B2(n13098), .ZN(
        n13100) );
  NAND2_X1 U15214 ( .A1(n13101), .A2(n13100), .ZN(n13312) );
  MUX2_X1 U15215 ( .A(P3_REG1_REG_18__SCAN_IN), .B(n13312), .S(n15281), .Z(
        P3_U3477) );
  AOI22_X1 U15216 ( .A1(n13103), .A2(n15214), .B1(n15224), .B2(n13102), .ZN(
        n13104) );
  NAND2_X1 U15217 ( .A1(n13105), .A2(n13104), .ZN(n13313) );
  MUX2_X1 U15218 ( .A(P3_REG1_REG_17__SCAN_IN), .B(n13313), .S(n15281), .Z(
        P3_U3476) );
  AOI22_X1 U15219 ( .A1(n13107), .A2(n15214), .B1(n15224), .B2(n13106), .ZN(
        n13108) );
  NAND2_X1 U15220 ( .A1(n13109), .A2(n13108), .ZN(n13314) );
  MUX2_X1 U15221 ( .A(P3_REG1_REG_16__SCAN_IN), .B(n13314), .S(n15281), .Z(
        P3_U3475) );
  AOI22_X1 U15222 ( .A1(n13111), .A2(n15214), .B1(n15224), .B2(n13110), .ZN(
        n13112) );
  NAND2_X1 U15223 ( .A1(n13113), .A2(n13112), .ZN(n13315) );
  MUX2_X1 U15224 ( .A(P3_REG1_REG_15__SCAN_IN), .B(n13315), .S(n15281), .Z(
        n13290) );
  INV_X1 U15225 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n14739) );
  AOI22_X1 U15226 ( .A1(n14739), .A2(keyinput52), .B1(n6841), .B2(keyinput56), 
        .ZN(n13114) );
  OAI221_X1 U15227 ( .B1(n14739), .B2(keyinput52), .C1(n6841), .C2(keyinput56), 
        .A(n13114), .ZN(n13118) );
  INV_X1 U15228 ( .A(P2_D_REG_24__SCAN_IN), .ZN(n15007) );
  AOI22_X1 U15229 ( .A1(n15007), .A2(keyinput14), .B1(n13862), .B2(keyinput60), 
        .ZN(n13115) );
  OAI221_X1 U15230 ( .B1(n15007), .B2(keyinput14), .C1(n13862), .C2(keyinput60), .A(n13115), .ZN(n13117) );
  XNOR2_X1 U15231 ( .A(n14485), .B(keyinput6), .ZN(n13116) );
  NOR3_X1 U15232 ( .A1(n13118), .A2(n13117), .A3(n13116), .ZN(n13146) );
  INV_X1 U15233 ( .A(P1_D_REG_19__SCAN_IN), .ZN(n13209) );
  AOI22_X1 U15234 ( .A1(n13208), .A2(keyinput19), .B1(keyinput50), .B2(n13209), 
        .ZN(n13119) );
  OAI221_X1 U15235 ( .B1(n13208), .B2(keyinput19), .C1(n13209), .C2(keyinput50), .A(n13119), .ZN(n13127) );
  AOI22_X1 U15236 ( .A1(n13122), .A2(keyinput59), .B1(n13121), .B2(keyinput33), 
        .ZN(n13120) );
  OAI221_X1 U15237 ( .B1(n13122), .B2(keyinput59), .C1(n13121), .C2(keyinput33), .A(n13120), .ZN(n13126) );
  XNOR2_X1 U15238 ( .A(P3_IR_REG_7__SCAN_IN), .B(keyinput21), .ZN(n13124) );
  XNOR2_X1 U15239 ( .A(keyinput10), .B(P3_REG2_REG_22__SCAN_IN), .ZN(n13123)
         );
  NAND2_X1 U15240 ( .A1(n13124), .A2(n13123), .ZN(n13125) );
  NOR3_X1 U15241 ( .A1(n13127), .A2(n13126), .A3(n13125), .ZN(n13145) );
  INV_X1 U15242 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n14510) );
  AOI22_X1 U15243 ( .A1(n12245), .A2(keyinput36), .B1(keyinput18), .B2(n14510), 
        .ZN(n13128) );
  OAI221_X1 U15244 ( .B1(n12245), .B2(keyinput36), .C1(n14510), .C2(keyinput18), .A(n13128), .ZN(n13131) );
  AOI22_X1 U15245 ( .A1(n13179), .A2(keyinput62), .B1(keyinput13), .B2(n15169), 
        .ZN(n13129) );
  OAI221_X1 U15246 ( .B1(n13179), .B2(keyinput62), .C1(n15169), .C2(keyinput13), .A(n13129), .ZN(n13130) );
  NOR2_X1 U15247 ( .A1(n13131), .A2(n13130), .ZN(n13144) );
  INV_X1 U15248 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n14588) );
  AOI22_X1 U15249 ( .A1(n7479), .A2(keyinput41), .B1(keyinput12), .B2(n14588), 
        .ZN(n13132) );
  OAI221_X1 U15250 ( .B1(n7479), .B2(keyinput41), .C1(n14588), .C2(keyinput12), 
        .A(n13132), .ZN(n13142) );
  XNOR2_X1 U15251 ( .A(P2_REG2_REG_2__SCAN_IN), .B(keyinput2), .ZN(n13136) );
  XNOR2_X1 U15252 ( .A(P2_IR_REG_6__SCAN_IN), .B(keyinput7), .ZN(n13135) );
  XNOR2_X1 U15253 ( .A(P2_REG3_REG_17__SCAN_IN), .B(keyinput27), .ZN(n13134)
         );
  XNOR2_X1 U15254 ( .A(P3_IR_REG_10__SCAN_IN), .B(keyinput16), .ZN(n13133) );
  AND4_X1 U15255 ( .A1(n13136), .A2(n13135), .A3(n13134), .A4(n13133), .ZN(
        n13140) );
  XNOR2_X1 U15256 ( .A(keyinput20), .B(P3_REG0_REG_0__SCAN_IN), .ZN(n13139) );
  XNOR2_X1 U15257 ( .A(P1_IR_REG_16__SCAN_IN), .B(keyinput22), .ZN(n13138) );
  XNOR2_X1 U15258 ( .A(P1_IR_REG_7__SCAN_IN), .B(keyinput53), .ZN(n13137) );
  NAND4_X1 U15259 ( .A1(n13140), .A2(n13139), .A3(n13138), .A4(n13137), .ZN(
        n13141) );
  NOR2_X1 U15260 ( .A1(n13142), .A2(n13141), .ZN(n13143) );
  AND4_X1 U15261 ( .A1(n13146), .A2(n13145), .A3(n13144), .A4(n13143), .ZN(
        n13174) );
  AOI22_X1 U15262 ( .A1(P2_REG1_REG_4__SCAN_IN), .A2(keyinput34), .B1(
        P3_D_REG_11__SCAN_IN), .B2(keyinput8), .ZN(n13147) );
  OAI221_X1 U15263 ( .B1(P2_REG1_REG_4__SCAN_IN), .B2(keyinput34), .C1(
        P3_D_REG_11__SCAN_IN), .C2(keyinput8), .A(n13147), .ZN(n13154) );
  AOI22_X1 U15264 ( .A1(P1_WR_REG_SCAN_IN), .A2(keyinput32), .B1(
        P2_REG1_REG_30__SCAN_IN), .B2(keyinput5), .ZN(n13148) );
  OAI221_X1 U15265 ( .B1(P1_WR_REG_SCAN_IN), .B2(keyinput32), .C1(
        P2_REG1_REG_30__SCAN_IN), .C2(keyinput5), .A(n13148), .ZN(n13153) );
  AOI22_X1 U15266 ( .A1(P3_DATAO_REG_23__SCAN_IN), .A2(keyinput25), .B1(
        P1_REG3_REG_28__SCAN_IN), .B2(keyinput28), .ZN(n13149) );
  OAI221_X1 U15267 ( .B1(P3_DATAO_REG_23__SCAN_IN), .B2(keyinput25), .C1(
        P1_REG3_REG_28__SCAN_IN), .C2(keyinput28), .A(n13149), .ZN(n13152) );
  AOI22_X1 U15268 ( .A1(P3_REG1_REG_0__SCAN_IN), .A2(keyinput31), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(keyinput63), .ZN(n13150) );
  OAI221_X1 U15269 ( .B1(P3_REG1_REG_0__SCAN_IN), .B2(keyinput31), .C1(
        P2_DATAO_REG_7__SCAN_IN), .C2(keyinput63), .A(n13150), .ZN(n13151) );
  NOR4_X1 U15270 ( .A1(n13154), .A2(n13153), .A3(n13152), .A4(n13151), .ZN(
        n13173) );
  AOI22_X1 U15271 ( .A1(SI_10_), .A2(keyinput39), .B1(SI_29_), .B2(keyinput48), 
        .ZN(n13155) );
  OAI221_X1 U15272 ( .B1(SI_10_), .B2(keyinput39), .C1(SI_29_), .C2(keyinput48), .A(n13155), .ZN(n13162) );
  AOI22_X1 U15273 ( .A1(P3_REG2_REG_24__SCAN_IN), .A2(keyinput17), .B1(
        P3_REG0_REG_29__SCAN_IN), .B2(keyinput9), .ZN(n13156) );
  OAI221_X1 U15274 ( .B1(P3_REG2_REG_24__SCAN_IN), .B2(keyinput17), .C1(
        P3_REG0_REG_29__SCAN_IN), .C2(keyinput9), .A(n13156), .ZN(n13161) );
  AOI22_X1 U15275 ( .A1(P2_ADDR_REG_3__SCAN_IN), .A2(keyinput44), .B1(
        P1_DATAO_REG_7__SCAN_IN), .B2(keyinput42), .ZN(n13157) );
  OAI221_X1 U15276 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(keyinput44), .C1(
        P1_DATAO_REG_7__SCAN_IN), .C2(keyinput42), .A(n13157), .ZN(n13160) );
  AOI22_X1 U15277 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(keyinput35), .B1(
        P1_D_REG_31__SCAN_IN), .B2(keyinput51), .ZN(n13158) );
  OAI221_X1 U15278 ( .B1(P2_IR_REG_25__SCAN_IN), .B2(keyinput35), .C1(
        P1_D_REG_31__SCAN_IN), .C2(keyinput51), .A(n13158), .ZN(n13159) );
  NOR4_X1 U15279 ( .A1(n13162), .A2(n13161), .A3(n13160), .A4(n13159), .ZN(
        n13172) );
  AOI22_X1 U15280 ( .A1(P3_REG2_REG_15__SCAN_IN), .A2(keyinput43), .B1(
        P3_REG0_REG_18__SCAN_IN), .B2(keyinput40), .ZN(n13163) );
  OAI221_X1 U15281 ( .B1(P3_REG2_REG_15__SCAN_IN), .B2(keyinput43), .C1(
        P3_REG0_REG_18__SCAN_IN), .C2(keyinput40), .A(n13163), .ZN(n13170) );
  AOI22_X1 U15282 ( .A1(P1_REG1_REG_8__SCAN_IN), .A2(keyinput26), .B1(
        P3_REG2_REG_9__SCAN_IN), .B2(keyinput4), .ZN(n13164) );
  OAI221_X1 U15283 ( .B1(P1_REG1_REG_8__SCAN_IN), .B2(keyinput26), .C1(
        P3_REG2_REG_9__SCAN_IN), .C2(keyinput4), .A(n13164), .ZN(n13169) );
  AOI22_X1 U15284 ( .A1(P1_REG0_REG_26__SCAN_IN), .A2(keyinput61), .B1(
        P3_D_REG_26__SCAN_IN), .B2(keyinput37), .ZN(n13165) );
  OAI221_X1 U15285 ( .B1(P1_REG0_REG_26__SCAN_IN), .B2(keyinput61), .C1(
        P3_D_REG_26__SCAN_IN), .C2(keyinput37), .A(n13165), .ZN(n13168) );
  AOI22_X1 U15286 ( .A1(P2_DATAO_REG_8__SCAN_IN), .A2(keyinput30), .B1(
        P3_IR_REG_30__SCAN_IN), .B2(keyinput47), .ZN(n13166) );
  OAI221_X1 U15287 ( .B1(P2_DATAO_REG_8__SCAN_IN), .B2(keyinput30), .C1(
        P3_IR_REG_30__SCAN_IN), .C2(keyinput47), .A(n13166), .ZN(n13167) );
  NOR4_X1 U15288 ( .A1(n13170), .A2(n13169), .A3(n13168), .A4(n13167), .ZN(
        n13171) );
  AND4_X1 U15289 ( .A1(n13174), .A2(n13173), .A3(n13172), .A4(n13171), .ZN(
        n13288) );
  AOI22_X1 U15290 ( .A1(n9767), .A2(keyinput108), .B1(n15007), .B2(keyinput78), 
        .ZN(n13175) );
  OAI221_X1 U15291 ( .B1(n9767), .B2(keyinput108), .C1(n15007), .C2(keyinput78), .A(n13175), .ZN(n13186) );
  INV_X1 U15292 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n13177) );
  AOI22_X1 U15293 ( .A1(n13177), .A2(keyinput92), .B1(n14477), .B2(keyinput110), .ZN(n13176) );
  OAI221_X1 U15294 ( .B1(n13177), .B2(keyinput92), .C1(n14477), .C2(
        keyinput110), .A(n13176), .ZN(n13185) );
  AOI22_X1 U15295 ( .A1(n13180), .A2(keyinput101), .B1(keyinput126), .B2(
        n13179), .ZN(n13178) );
  OAI221_X1 U15296 ( .B1(n13180), .B2(keyinput101), .C1(n13179), .C2(
        keyinput126), .A(n13178), .ZN(n13184) );
  AOI22_X1 U15297 ( .A1(n14588), .A2(keyinput76), .B1(n13182), .B2(keyinput95), 
        .ZN(n13181) );
  OAI221_X1 U15298 ( .B1(n14588), .B2(keyinput76), .C1(n13182), .C2(keyinput95), .A(n13181), .ZN(n13183) );
  NOR4_X1 U15299 ( .A1(n13186), .A2(n13185), .A3(n13184), .A4(n13183), .ZN(
        n13266) );
  OAI22_X1 U15300 ( .A1(P2_DATAO_REG_0__SCAN_IN), .A2(keyinput121), .B1(
        keyinput64), .B2(P1_ADDR_REG_13__SCAN_IN), .ZN(n13187) );
  AOI221_X1 U15301 ( .B1(P2_DATAO_REG_0__SCAN_IN), .B2(keyinput121), .C1(
        P1_ADDR_REG_13__SCAN_IN), .C2(keyinput64), .A(n13187), .ZN(n13194) );
  OAI22_X1 U15302 ( .A1(P2_REG1_REG_14__SCAN_IN), .A2(keyinput116), .B1(
        keyinput75), .B2(P1_ADDR_REG_2__SCAN_IN), .ZN(n13188) );
  AOI221_X1 U15303 ( .B1(P2_REG1_REG_14__SCAN_IN), .B2(keyinput116), .C1(
        P1_ADDR_REG_2__SCAN_IN), .C2(keyinput75), .A(n13188), .ZN(n13193) );
  OAI22_X1 U15304 ( .A1(P3_REG0_REG_0__SCAN_IN), .A2(keyinput84), .B1(
        P2_IR_REG_6__SCAN_IN), .B2(keyinput71), .ZN(n13189) );
  AOI221_X1 U15305 ( .B1(P3_REG0_REG_0__SCAN_IN), .B2(keyinput84), .C1(
        keyinput71), .C2(P2_IR_REG_6__SCAN_IN), .A(n13189), .ZN(n13192) );
  OAI22_X1 U15306 ( .A1(P1_DATAO_REG_7__SCAN_IN), .A2(keyinput106), .B1(
        keyinput102), .B2(P3_REG2_REG_0__SCAN_IN), .ZN(n13190) );
  AOI221_X1 U15307 ( .B1(P1_DATAO_REG_7__SCAN_IN), .B2(keyinput106), .C1(
        P3_REG2_REG_0__SCAN_IN), .C2(keyinput102), .A(n13190), .ZN(n13191) );
  NAND4_X1 U15308 ( .A1(n13194), .A2(n13193), .A3(n13192), .A4(n13191), .ZN(
        n13204) );
  OAI22_X1 U15309 ( .A1(P2_REG1_REG_21__SCAN_IN), .A2(keyinput123), .B1(
        P1_ADDR_REG_9__SCAN_IN), .B2(keyinput70), .ZN(n13195) );
  AOI221_X1 U15310 ( .B1(P2_REG1_REG_21__SCAN_IN), .B2(keyinput123), .C1(
        keyinput70), .C2(P1_ADDR_REG_9__SCAN_IN), .A(n13195), .ZN(n13202) );
  OAI22_X1 U15311 ( .A1(P3_IR_REG_23__SCAN_IN), .A2(keyinput97), .B1(
        keyinput107), .B2(P3_REG2_REG_15__SCAN_IN), .ZN(n13196) );
  AOI221_X1 U15312 ( .B1(P3_IR_REG_23__SCAN_IN), .B2(keyinput97), .C1(
        P3_REG2_REG_15__SCAN_IN), .C2(keyinput107), .A(n13196), .ZN(n13201) );
  OAI22_X1 U15313 ( .A1(P1_REG0_REG_26__SCAN_IN), .A2(keyinput125), .B1(
        keyinput96), .B2(P1_WR_REG_SCAN_IN), .ZN(n13197) );
  AOI221_X1 U15314 ( .B1(P1_REG0_REG_26__SCAN_IN), .B2(keyinput125), .C1(
        P1_WR_REG_SCAN_IN), .C2(keyinput96), .A(n13197), .ZN(n13200) );
  OAI22_X1 U15315 ( .A1(P3_IR_REG_30__SCAN_IN), .A2(keyinput111), .B1(
        P2_REG1_REG_2__SCAN_IN), .B2(keyinput87), .ZN(n13198) );
  AOI221_X1 U15316 ( .B1(P3_IR_REG_30__SCAN_IN), .B2(keyinput111), .C1(
        keyinput87), .C2(P2_REG1_REG_2__SCAN_IN), .A(n13198), .ZN(n13199) );
  NAND4_X1 U15317 ( .A1(n13202), .A2(n13201), .A3(n13200), .A4(n13199), .ZN(
        n13203) );
  NOR2_X1 U15318 ( .A1(n13204), .A2(n13203), .ZN(n13231) );
  AOI22_X1 U15319 ( .A1(n15090), .A2(keyinput98), .B1(n13206), .B2(keyinput73), 
        .ZN(n13205) );
  OAI221_X1 U15320 ( .B1(n15090), .B2(keyinput98), .C1(n13206), .C2(keyinput73), .A(n13205), .ZN(n13212) );
  INV_X1 U15321 ( .A(SI_0_), .ZN(n13279) );
  AOI22_X1 U15322 ( .A1(n13279), .A2(keyinput118), .B1(n13208), .B2(keyinput83), .ZN(n13207) );
  OAI221_X1 U15323 ( .B1(n13279), .B2(keyinput118), .C1(n13208), .C2(
        keyinput83), .A(n13207), .ZN(n13211) );
  XNOR2_X1 U15324 ( .A(n13209), .B(keyinput114), .ZN(n13210) );
  NOR3_X1 U15325 ( .A1(n13212), .A2(n13211), .A3(n13210), .ZN(n13230) );
  AOI22_X1 U15326 ( .A1(n14503), .A2(keyinput109), .B1(n13658), .B2(
        keyinput122), .ZN(n13213) );
  OAI221_X1 U15327 ( .B1(n14503), .B2(keyinput109), .C1(n13658), .C2(
        keyinput122), .A(n13213), .ZN(n13217) );
  AOI22_X1 U15328 ( .A1(n13215), .A2(keyinput112), .B1(keyinput81), .B2(n12226), .ZN(n13214) );
  OAI221_X1 U15329 ( .B1(n13215), .B2(keyinput112), .C1(n12226), .C2(
        keyinput81), .A(n13214), .ZN(n13216) );
  NOR2_X1 U15330 ( .A1(n13217), .A2(n13216), .ZN(n13229) );
  AOI22_X1 U15331 ( .A1(n13219), .A2(keyinput89), .B1(n7479), .B2(keyinput105), 
        .ZN(n13218) );
  OAI221_X1 U15332 ( .B1(n13219), .B2(keyinput89), .C1(n7479), .C2(keyinput105), .A(n13218), .ZN(n13227) );
  INV_X1 U15333 ( .A(P3_REG0_REG_18__SCAN_IN), .ZN(n13221) );
  AOI22_X1 U15334 ( .A1(n13222), .A2(keyinput88), .B1(keyinput104), .B2(n13221), .ZN(n13220) );
  OAI221_X1 U15335 ( .B1(n13222), .B2(keyinput88), .C1(n13221), .C2(
        keyinput104), .A(n13220), .ZN(n13226) );
  XNOR2_X1 U15336 ( .A(keyinput67), .B(P2_REG3_REG_3__SCAN_IN), .ZN(n13224) );
  XNOR2_X1 U15337 ( .A(keyinput82), .B(P1_ADDR_REG_12__SCAN_IN), .ZN(n13223)
         );
  NAND2_X1 U15338 ( .A1(n13224), .A2(n13223), .ZN(n13225) );
  NOR3_X1 U15339 ( .A1(n13227), .A2(n13226), .A3(n13225), .ZN(n13228) );
  AND4_X1 U15340 ( .A1(n13231), .A2(n13230), .A3(n13229), .A4(n13228), .ZN(
        n13265) );
  OAI22_X1 U15341 ( .A1(P3_REG2_REG_22__SCAN_IN), .A2(keyinput74), .B1(
        keyinput119), .B2(P2_D_REG_19__SCAN_IN), .ZN(n13232) );
  AOI221_X1 U15342 ( .B1(P3_REG2_REG_22__SCAN_IN), .B2(keyinput74), .C1(
        P2_D_REG_19__SCAN_IN), .C2(keyinput119), .A(n13232), .ZN(n13239) );
  OAI22_X1 U15343 ( .A1(SI_10_), .A2(keyinput103), .B1(keyinput90), .B2(
        P1_REG1_REG_8__SCAN_IN), .ZN(n13233) );
  AOI221_X1 U15344 ( .B1(SI_10_), .B2(keyinput103), .C1(P1_REG1_REG_8__SCAN_IN), .C2(keyinput90), .A(n13233), .ZN(n13238) );
  OAI22_X1 U15345 ( .A1(P1_DATAO_REG_31__SCAN_IN), .A2(keyinput124), .B1(
        keyinput77), .B2(P3_ADDR_REG_7__SCAN_IN), .ZN(n13234) );
  AOI221_X1 U15346 ( .B1(P1_DATAO_REG_31__SCAN_IN), .B2(keyinput124), .C1(
        P3_ADDR_REG_7__SCAN_IN), .C2(keyinput77), .A(n13234), .ZN(n13237) );
  OAI22_X1 U15347 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(keyinput86), .B1(
        P2_REG3_REG_17__SCAN_IN), .B2(keyinput91), .ZN(n13235) );
  AOI221_X1 U15348 ( .B1(P1_IR_REG_16__SCAN_IN), .B2(keyinput86), .C1(
        keyinput91), .C2(P2_REG3_REG_17__SCAN_IN), .A(n13235), .ZN(n13236) );
  AND4_X1 U15349 ( .A1(n13239), .A2(n13238), .A3(n13237), .A4(n13236), .ZN(
        n13253) );
  XNOR2_X1 U15350 ( .A(n13240), .B(keyinput72), .ZN(n13251) );
  XNOR2_X1 U15351 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(keyinput127), .ZN(n13244)
         );
  XNOR2_X1 U15352 ( .A(P3_IR_REG_7__SCAN_IN), .B(keyinput85), .ZN(n13243) );
  XNOR2_X1 U15353 ( .A(P2_IR_REG_25__SCAN_IN), .B(keyinput99), .ZN(n13242) );
  XNOR2_X1 U15354 ( .A(P2_IR_REG_13__SCAN_IN), .B(keyinput79), .ZN(n13241) );
  NAND4_X1 U15355 ( .A1(n13244), .A2(n13243), .A3(n13242), .A4(n13241), .ZN(
        n13250) );
  XNOR2_X1 U15356 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(keyinput94), .ZN(n13248)
         );
  XNOR2_X1 U15357 ( .A(P3_IR_REG_10__SCAN_IN), .B(keyinput80), .ZN(n13247) );
  XNOR2_X1 U15358 ( .A(P1_IR_REG_7__SCAN_IN), .B(keyinput117), .ZN(n13246) );
  XNOR2_X1 U15359 ( .A(P2_REG2_REG_2__SCAN_IN), .B(keyinput66), .ZN(n13245) );
  NAND4_X1 U15360 ( .A1(n13248), .A2(n13247), .A3(n13246), .A4(n13245), .ZN(
        n13249) );
  NOR3_X1 U15361 ( .A1(n13251), .A2(n13250), .A3(n13249), .ZN(n13252) );
  NAND2_X1 U15362 ( .A1(n13253), .A2(n13252), .ZN(n13263) );
  OAI22_X1 U15363 ( .A1(P1_D_REG_31__SCAN_IN), .A2(keyinput115), .B1(
        keyinput113), .B2(P2_D_REG_16__SCAN_IN), .ZN(n13254) );
  AOI221_X1 U15364 ( .B1(P1_D_REG_31__SCAN_IN), .B2(keyinput115), .C1(
        P2_D_REG_16__SCAN_IN), .C2(keyinput113), .A(n13254), .ZN(n13261) );
  OAI22_X1 U15365 ( .A1(P3_D_REG_31__SCAN_IN), .A2(keyinput93), .B1(
        P2_REG1_REG_30__SCAN_IN), .B2(keyinput69), .ZN(n13255) );
  AOI221_X1 U15366 ( .B1(P3_D_REG_31__SCAN_IN), .B2(keyinput93), .C1(
        keyinput69), .C2(P2_REG1_REG_30__SCAN_IN), .A(n13255), .ZN(n13260) );
  OAI22_X1 U15367 ( .A1(n11326), .A2(keyinput68), .B1(n13276), .B2(keyinput65), 
        .ZN(n13256) );
  AOI221_X1 U15368 ( .B1(n11326), .B2(keyinput68), .C1(keyinput65), .C2(n13276), .A(n13256), .ZN(n13259) );
  OAI22_X1 U15369 ( .A1(n12245), .A2(keyinput100), .B1(keyinput120), .B2(
        P2_RD_REG_SCAN_IN), .ZN(n13257) );
  AOI221_X1 U15370 ( .B1(n12245), .B2(keyinput100), .C1(P2_RD_REG_SCAN_IN), 
        .C2(keyinput120), .A(n13257), .ZN(n13258) );
  NAND4_X1 U15371 ( .A1(n13261), .A2(n13260), .A3(n13259), .A4(n13258), .ZN(
        n13262) );
  NOR2_X1 U15372 ( .A1(n13263), .A2(n13262), .ZN(n13264) );
  NAND3_X1 U15373 ( .A1(n13266), .A2(n13265), .A3(n13264), .ZN(n13287) );
  AOI22_X1 U15374 ( .A1(P2_D_REG_19__SCAN_IN), .A2(keyinput55), .B1(
        P3_D_REG_31__SCAN_IN), .B2(keyinput29), .ZN(n13267) );
  OAI221_X1 U15375 ( .B1(P2_D_REG_19__SCAN_IN), .B2(keyinput55), .C1(
        P3_D_REG_31__SCAN_IN), .C2(keyinput29), .A(n13267), .ZN(n13274) );
  AOI22_X1 U15376 ( .A1(P2_DATAO_REG_0__SCAN_IN), .A2(keyinput57), .B1(
        P1_DATAO_REG_12__SCAN_IN), .B2(keyinput24), .ZN(n13268) );
  OAI221_X1 U15377 ( .B1(P2_DATAO_REG_0__SCAN_IN), .B2(keyinput57), .C1(
        P1_DATAO_REG_12__SCAN_IN), .C2(keyinput24), .A(n13268), .ZN(n13273) );
  AOI22_X1 U15378 ( .A1(P1_ADDR_REG_13__SCAN_IN), .A2(keyinput0), .B1(
        P2_IR_REG_13__SCAN_IN), .B2(keyinput15), .ZN(n13269) );
  OAI221_X1 U15379 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(keyinput0), .C1(
        P2_IR_REG_13__SCAN_IN), .C2(keyinput15), .A(n13269), .ZN(n13272) );
  AOI22_X1 U15380 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(keyinput3), .B1(n13658), 
        .B2(keyinput58), .ZN(n13270) );
  OAI221_X1 U15381 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(keyinput3), .C1(n13658), 
        .C2(keyinput58), .A(n13270), .ZN(n13271) );
  NOR4_X1 U15382 ( .A1(n13274), .A2(n13273), .A3(n13272), .A4(n13271), .ZN(
        n13286) );
  AOI22_X1 U15383 ( .A1(n14477), .A2(keyinput46), .B1(keyinput1), .B2(n13276), 
        .ZN(n13275) );
  OAI221_X1 U15384 ( .B1(n14477), .B2(keyinput46), .C1(n13276), .C2(keyinput1), 
        .A(n13275), .ZN(n13284) );
  INV_X1 U15385 ( .A(P2_D_REG_16__SCAN_IN), .ZN(n15008) );
  AOI22_X1 U15386 ( .A1(n15099), .A2(keyinput38), .B1(keyinput49), .B2(n15008), 
        .ZN(n13277) );
  OAI221_X1 U15387 ( .B1(n15099), .B2(keyinput38), .C1(n15008), .C2(keyinput49), .A(n13277), .ZN(n13283) );
  INV_X1 U15388 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n14532) );
  AOI22_X1 U15389 ( .A1(n13279), .A2(keyinput54), .B1(keyinput11), .B2(n14532), 
        .ZN(n13278) );
  OAI221_X1 U15390 ( .B1(n13279), .B2(keyinput54), .C1(n14532), .C2(keyinput11), .A(n13278), .ZN(n13282) );
  AOI22_X1 U15391 ( .A1(n14503), .A2(keyinput45), .B1(n9675), .B2(keyinput23), 
        .ZN(n13280) );
  OAI221_X1 U15392 ( .B1(n14503), .B2(keyinput45), .C1(n9675), .C2(keyinput23), 
        .A(n13280), .ZN(n13281) );
  NOR4_X1 U15393 ( .A1(n13284), .A2(n13283), .A3(n13282), .A4(n13281), .ZN(
        n13285) );
  NAND4_X1 U15394 ( .A1(n13288), .A2(n13287), .A3(n13286), .A4(n13285), .ZN(
        n13289) );
  XNOR2_X1 U15395 ( .A(n13290), .B(n13289), .ZN(P3_U3474) );
  INV_X1 U15396 ( .A(n13291), .ZN(n13293) );
  OAI22_X1 U15397 ( .A1(n13294), .A2(n13293), .B1(n13298), .B2(n13292), .ZN(
        n13296) );
  NAND2_X1 U15398 ( .A1(n13296), .A2(n13295), .ZN(n13300) );
  MUX2_X1 U15399 ( .A(n13301), .B(P3_REG0_REG_29__SCAN_IN), .S(n15268), .Z(
        P3_U3456) );
  MUX2_X1 U15400 ( .A(P3_REG0_REG_28__SCAN_IN), .B(n13302), .S(n15266), .Z(
        P3_U3455) );
  MUX2_X1 U15401 ( .A(P3_REG0_REG_27__SCAN_IN), .B(n13303), .S(n15266), .Z(
        P3_U3454) );
  MUX2_X1 U15402 ( .A(P3_REG0_REG_26__SCAN_IN), .B(n13304), .S(n15266), .Z(
        P3_U3453) );
  MUX2_X1 U15403 ( .A(P3_REG0_REG_25__SCAN_IN), .B(n13305), .S(n15266), .Z(
        P3_U3452) );
  MUX2_X1 U15404 ( .A(P3_REG0_REG_24__SCAN_IN), .B(n13306), .S(n15266), .Z(
        P3_U3451) );
  MUX2_X1 U15405 ( .A(P3_REG0_REG_23__SCAN_IN), .B(n13307), .S(n15266), .Z(
        P3_U3450) );
  MUX2_X1 U15406 ( .A(P3_REG0_REG_22__SCAN_IN), .B(n13308), .S(n15266), .Z(
        P3_U3449) );
  MUX2_X1 U15407 ( .A(P3_REG0_REG_21__SCAN_IN), .B(n13309), .S(n15266), .Z(
        P3_U3448) );
  MUX2_X1 U15408 ( .A(P3_REG0_REG_20__SCAN_IN), .B(n13310), .S(n15266), .Z(
        P3_U3447) );
  MUX2_X1 U15409 ( .A(P3_REG0_REG_19__SCAN_IN), .B(n13311), .S(n15266), .Z(
        P3_U3446) );
  MUX2_X1 U15410 ( .A(P3_REG0_REG_18__SCAN_IN), .B(n13312), .S(n15266), .Z(
        P3_U3444) );
  MUX2_X1 U15411 ( .A(P3_REG0_REG_17__SCAN_IN), .B(n13313), .S(n15266), .Z(
        P3_U3441) );
  MUX2_X1 U15412 ( .A(P3_REG0_REG_16__SCAN_IN), .B(n13314), .S(n15266), .Z(
        P3_U3438) );
  MUX2_X1 U15413 ( .A(P3_REG0_REG_15__SCAN_IN), .B(n13315), .S(n15266), .Z(
        P3_U3435) );
  MUX2_X1 U15414 ( .A(P3_REG0_REG_0__SCAN_IN), .B(n13316), .S(n15266), .Z(
        P3_U3390) );
  MUX2_X1 U15415 ( .A(P3_D_REG_1__SCAN_IN), .B(n13317), .S(n13318), .Z(
        P3_U3377) );
  MUX2_X1 U15416 ( .A(P3_D_REG_0__SCAN_IN), .B(n13319), .S(n13318), .Z(
        P3_U3376) );
  INV_X1 U15417 ( .A(SI_31_), .ZN(n13327) );
  NAND2_X1 U15418 ( .A1(n13321), .A2(n13320), .ZN(n13326) );
  INV_X1 U15419 ( .A(n13322), .ZN(n13324) );
  INV_X1 U15420 ( .A(P3_IR_REG_30__SCAN_IN), .ZN(n13323) );
  NAND4_X1 U15421 ( .A1(n13324), .A2(P3_STATE_REG_SCAN_IN), .A3(
        P3_IR_REG_31__SCAN_IN), .A4(n13323), .ZN(n13325) );
  OAI211_X1 U15422 ( .C1(n13327), .C2(n13335), .A(n13326), .B(n13325), .ZN(
        P3_U3264) );
  INV_X1 U15423 ( .A(n13328), .ZN(n13330) );
  OAI222_X1 U15424 ( .A1(n13333), .A2(n13330), .B1(n6485), .B2(P3_U3151), .C1(
        n13329), .C2(n13335), .ZN(P3_U3267) );
  INV_X1 U15425 ( .A(SI_27_), .ZN(n13334) );
  INV_X1 U15426 ( .A(n13331), .ZN(n13332) );
  OAI222_X1 U15427 ( .A1(P3_U3151), .A2(n6489), .B1(n13335), .B2(n13334), .C1(
        n13333), .C2(n13332), .ZN(P3_U3268) );
  AOI21_X1 U15428 ( .B1(n13337), .B2(n13336), .A(n13428), .ZN(n13339) );
  INV_X1 U15429 ( .A(n13431), .ZN(n13592) );
  OAI22_X1 U15430 ( .A1(n13592), .A2(n13370), .B1(n13556), .B2(n13591), .ZN(
        n13778) );
  OAI22_X1 U15431 ( .A1(n13621), .A2(n13372), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13340), .ZN(n13341) );
  AOI21_X1 U15432 ( .B1(n13778), .B2(n13374), .A(n13341), .ZN(n13342) );
  XOR2_X1 U15433 ( .A(n13344), .B(n13343), .Z(n13348) );
  OAI22_X1 U15434 ( .A1(n13581), .A2(n13370), .B1(n13579), .B2(n13591), .ZN(
        n13805) );
  AOI22_X1 U15435 ( .A1(n13805), .A2(n13374), .B1(P2_REG3_REG_23__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13345) );
  OAI21_X1 U15436 ( .B1(n13675), .B2(n13372), .A(n13345), .ZN(n13346) );
  AOI21_X1 U15437 ( .B1(n13806), .B2(n13426), .A(n13346), .ZN(n13347) );
  OAI21_X1 U15438 ( .B1(n13348), .B2(n13428), .A(n13347), .ZN(P2_U3188) );
  OAI21_X1 U15439 ( .B1(n13351), .B2(n13350), .A(n13349), .ZN(n13352) );
  NAND2_X1 U15440 ( .A1(n13352), .A2(n13391), .ZN(n13357) );
  INV_X1 U15441 ( .A(n13730), .ZN(n13355) );
  AND2_X1 U15442 ( .A1(n13566), .A2(n13420), .ZN(n13353) );
  AOI21_X1 U15443 ( .B1(n13361), .B2(n13524), .A(n13353), .ZN(n13825) );
  NAND2_X1 U15444 ( .A1(P2_U3088), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n13519)
         );
  OAI21_X1 U15445 ( .B1(n13424), .B2(n13825), .A(n13519), .ZN(n13354) );
  AOI21_X1 U15446 ( .B1(n13355), .B2(n13422), .A(n13354), .ZN(n13356) );
  OAI211_X1 U15447 ( .C1(n6703), .C2(n13415), .A(n13357), .B(n13356), .ZN(
        P2_U3191) );
  OAI211_X1 U15448 ( .C1(n13358), .C2(n13360), .A(n13359), .B(n13391), .ZN(
        n13366) );
  INV_X1 U15449 ( .A(n13704), .ZN(n13364) );
  AOI22_X1 U15450 ( .A1(n13545), .A2(n13524), .B1(n13420), .B2(n13361), .ZN(
        n13708) );
  OAI22_X1 U15451 ( .A1(n13708), .A2(n13424), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13362), .ZN(n13363) );
  AOI21_X1 U15452 ( .B1(n13364), .B2(n13422), .A(n13363), .ZN(n13365) );
  OAI211_X1 U15453 ( .C1(n13699), .C2(n13415), .A(n13366), .B(n13365), .ZN(
        P2_U3195) );
  INV_X1 U15454 ( .A(n13791), .ZN(n13640) );
  OAI211_X1 U15455 ( .C1(n13369), .C2(n13368), .A(n13367), .B(n13391), .ZN(
        n13376) );
  OAI22_X1 U15456 ( .A1(n13556), .A2(n13370), .B1(n13581), .B2(n13591), .ZN(
        n13649) );
  OAI22_X1 U15457 ( .A1(n13645), .A2(n13372), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13371), .ZN(n13373) );
  AOI21_X1 U15458 ( .B1(n13649), .B2(n13374), .A(n13373), .ZN(n13375) );
  OAI211_X1 U15459 ( .C1(n13640), .C2(n13415), .A(n13376), .B(n13375), .ZN(
        P2_U3197) );
  INV_X1 U15460 ( .A(n13378), .ZN(n13379) );
  AOI211_X1 U15461 ( .C1(n13380), .C2(n13377), .A(n13428), .B(n13379), .ZN(
        n13385) );
  AND2_X1 U15462 ( .A1(n13580), .A2(n13420), .ZN(n13381) );
  AOI21_X1 U15463 ( .B1(n13552), .B2(n13524), .A(n13381), .ZN(n13796) );
  NAND2_X1 U15464 ( .A1(n13795), .A2(n13426), .ZN(n13383) );
  AOI22_X1 U15465 ( .A1(n13660), .A2(n13422), .B1(P2_REG3_REG_24__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13382) );
  OAI211_X1 U15466 ( .C1(n13796), .C2(n13424), .A(n13383), .B(n13382), .ZN(
        n13384) );
  OR2_X1 U15467 ( .A1(n13385), .A2(n13384), .ZN(P2_U3201) );
  NOR2_X1 U15468 ( .A1(n13386), .A2(n7236), .ZN(n13390) );
  OAI22_X1 U15469 ( .A1(n13390), .A2(n13389), .B1(n13358), .B2(n13388), .ZN(
        n13392) );
  NAND2_X1 U15470 ( .A1(n13392), .A2(n13391), .ZN(n13397) );
  AND2_X1 U15471 ( .A1(n13575), .A2(n13420), .ZN(n13393) );
  AOI21_X1 U15472 ( .B1(n13433), .B2(n13524), .A(n13393), .ZN(n13716) );
  OAI22_X1 U15473 ( .A1(n13424), .A2(n13716), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13394), .ZN(n13395) );
  AOI21_X1 U15474 ( .B1(n13719), .B2(n13422), .A(n13395), .ZN(n13396) );
  OAI211_X1 U15475 ( .C1(n13722), .C2(n13415), .A(n13397), .B(n13396), .ZN(
        P2_U3205) );
  INV_X1 U15476 ( .A(n13811), .ZN(n13694) );
  AOI21_X1 U15477 ( .B1(n13399), .B2(n13398), .A(n13428), .ZN(n13401) );
  NAND2_X1 U15478 ( .A1(n13401), .A2(n13400), .ZN(n13406) );
  AND2_X1 U15479 ( .A1(n13433), .A2(n13420), .ZN(n13402) );
  AOI21_X1 U15480 ( .B1(n13580), .B2(n13524), .A(n13402), .ZN(n13685) );
  OAI22_X1 U15481 ( .A1(n13685), .A2(n13424), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13403), .ZN(n13404) );
  AOI21_X1 U15482 ( .B1(n13691), .B2(n13422), .A(n13404), .ZN(n13405) );
  OAI211_X1 U15483 ( .C1(n13694), .C2(n13415), .A(n13406), .B(n13405), .ZN(
        P2_U3207) );
  INV_X1 U15484 ( .A(n13745), .ZN(n13833) );
  AOI211_X1 U15485 ( .C1(n13409), .C2(n13408), .A(n13428), .B(n13407), .ZN(
        n13410) );
  INV_X1 U15486 ( .A(n13410), .ZN(n13414) );
  AOI22_X1 U15487 ( .A1(n13575), .A2(n13524), .B1(n13420), .B2(n13567), .ZN(
        n13831) );
  OAI22_X1 U15488 ( .A1(n13424), .A2(n13831), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13411), .ZN(n13412) );
  AOI21_X1 U15489 ( .B1(n13748), .B2(n13422), .A(n13412), .ZN(n13413) );
  OAI211_X1 U15490 ( .C1(n13833), .C2(n13415), .A(n13414), .B(n13413), .ZN(
        P2_U3210) );
  INV_X1 U15491 ( .A(n13417), .ZN(n13418) );
  AOI21_X1 U15492 ( .B1(n13419), .B2(n13416), .A(n13418), .ZN(n13429) );
  AND2_X1 U15493 ( .A1(n13552), .A2(n13420), .ZN(n13421) );
  AOI21_X1 U15494 ( .B1(n13585), .B2(n13524), .A(n13421), .ZN(n13783) );
  AOI22_X1 U15495 ( .A1(n13632), .A2(n13422), .B1(P2_REG3_REG_26__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13423) );
  OAI21_X1 U15496 ( .B1(n13783), .B2(n13424), .A(n13423), .ZN(n13425) );
  AOI21_X1 U15497 ( .B1(n13635), .B2(n13426), .A(n13425), .ZN(n13427) );
  OAI21_X1 U15498 ( .B1(n13429), .B2(n13428), .A(n13427), .ZN(P2_U3212) );
  MUX2_X1 U15499 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n13430), .S(n6492), .Z(
        P2_U3561) );
  MUX2_X1 U15500 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n13431), .S(n6492), .Z(
        P2_U3559) );
  MUX2_X1 U15501 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n13585), .S(n6492), .Z(
        P2_U3558) );
  MUX2_X1 U15502 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n13432), .S(n6492), .Z(
        P2_U3557) );
  MUX2_X1 U15503 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n13552), .S(n6492), .Z(
        P2_U3556) );
  MUX2_X1 U15504 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n13550), .S(n6492), .Z(
        P2_U3555) );
  MUX2_X1 U15505 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(n13580), .S(n6492), .Z(
        P2_U3554) );
  MUX2_X1 U15506 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n13545), .S(n6492), .Z(
        P2_U3553) );
  MUX2_X1 U15507 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n13433), .S(P2_U3947), .Z(
        P2_U3552) );
  MUX2_X1 U15508 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n13575), .S(P2_U3947), .Z(
        P2_U3550) );
  MUX2_X1 U15509 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n13566), .S(P2_U3947), .Z(
        P2_U3549) );
  MUX2_X1 U15510 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n13567), .S(n6492), .Z(
        P2_U3548) );
  MUX2_X1 U15511 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n13434), .S(n6492), .Z(
        P2_U3547) );
  MUX2_X1 U15512 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n13435), .S(n6492), .Z(
        P2_U3546) );
  MUX2_X1 U15513 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n13436), .S(n6492), .Z(
        P2_U3545) );
  MUX2_X1 U15514 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n13437), .S(n6492), .Z(
        P2_U3544) );
  MUX2_X1 U15515 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n13438), .S(n6492), .Z(
        P2_U3543) );
  MUX2_X1 U15516 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n13439), .S(n6492), .Z(
        P2_U3542) );
  MUX2_X1 U15517 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n13440), .S(n6492), .Z(
        P2_U3541) );
  MUX2_X1 U15518 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n13441), .S(n6492), .Z(
        P2_U3540) );
  MUX2_X1 U15519 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n13442), .S(n6492), .Z(
        P2_U3539) );
  MUX2_X1 U15520 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n13443), .S(n6492), .Z(
        P2_U3538) );
  MUX2_X1 U15521 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n13444), .S(n6492), .Z(
        P2_U3537) );
  MUX2_X1 U15522 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(n13445), .S(n6492), .Z(
        P2_U3536) );
  MUX2_X1 U15523 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n13446), .S(n6492), .Z(
        P2_U3535) );
  MUX2_X1 U15524 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(n13447), .S(n6492), .Z(
        P2_U3534) );
  MUX2_X1 U15525 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(n13448), .S(n6492), .Z(
        P2_U3533) );
  MUX2_X1 U15526 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n9998), .S(n6492), .Z(
        P2_U3532) );
  MUX2_X1 U15527 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n9205), .S(n6492), .Z(
        P2_U3531) );
  NOR2_X1 U15528 ( .A1(n14894), .A2(n13449), .ZN(n13450) );
  AOI211_X1 U15529 ( .C1(n14954), .C2(P2_ADDR_REG_7__SCAN_IN), .A(n13451), .B(
        n13450), .ZN(n13463) );
  MUX2_X1 U15530 ( .A(n9840), .B(P2_REG1_REG_7__SCAN_IN), .S(n13456), .Z(
        n13452) );
  NAND3_X1 U15531 ( .A1(n13454), .A2(n13453), .A3(n13452), .ZN(n13455) );
  NAND3_X1 U15532 ( .A1(n14956), .A2(n13469), .A3(n13455), .ZN(n13462) );
  MUX2_X1 U15533 ( .A(n10686), .B(P2_REG2_REG_7__SCAN_IN), .S(n13456), .Z(
        n13457) );
  NAND3_X1 U15534 ( .A1(n13459), .A2(n13458), .A3(n13457), .ZN(n13460) );
  NAND3_X1 U15535 ( .A1(n14961), .A2(n13475), .A3(n13460), .ZN(n13461) );
  NAND3_X1 U15536 ( .A1(n13463), .A2(n13462), .A3(n13461), .ZN(P2_U3221) );
  INV_X1 U15537 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n13465) );
  OAI21_X1 U15538 ( .B1(n14901), .B2(n13465), .A(n13464), .ZN(n13466) );
  AOI21_X1 U15539 ( .B1(n13472), .B2(n14959), .A(n13466), .ZN(n13480) );
  MUX2_X1 U15540 ( .A(n9843), .B(P2_REG1_REG_8__SCAN_IN), .S(n13472), .Z(
        n13467) );
  NAND3_X1 U15541 ( .A1(n13469), .A2(n13468), .A3(n13467), .ZN(n13470) );
  NAND3_X1 U15542 ( .A1(n14956), .A2(n13471), .A3(n13470), .ZN(n13479) );
  MUX2_X1 U15543 ( .A(n10719), .B(P2_REG2_REG_8__SCAN_IN), .S(n13472), .Z(
        n13473) );
  NAND3_X1 U15544 ( .A1(n13475), .A2(n13474), .A3(n13473), .ZN(n13476) );
  NAND3_X1 U15545 ( .A1(n14961), .A2(n13477), .A3(n13476), .ZN(n13478) );
  NAND3_X1 U15546 ( .A1(n13480), .A2(n13479), .A3(n13478), .ZN(P2_U3222) );
  NAND2_X1 U15547 ( .A1(P2_REG2_REG_17__SCAN_IN), .A2(n14943), .ZN(n13490) );
  INV_X1 U15548 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n13482) );
  INV_X1 U15549 ( .A(n13490), .ZN(n13481) );
  AOI21_X1 U15550 ( .B1(n13482), .B2(n13506), .A(n13481), .ZN(n14948) );
  INV_X1 U15551 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n13489) );
  XOR2_X1 U15552 ( .A(P2_REG2_REG_16__SCAN_IN), .B(n14935), .Z(n14933) );
  INV_X1 U15553 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n13484) );
  INV_X1 U15554 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n13483) );
  OR2_X1 U15555 ( .A1(n13494), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n14886) );
  MUX2_X1 U15556 ( .A(n13483), .B(P2_REG2_REG_12__SCAN_IN), .S(n13497), .Z(
        n14887) );
  AOI21_X1 U15557 ( .B1(n14888), .B2(n14886), .A(n14887), .ZN(n14890) );
  AOI21_X1 U15558 ( .B1(n13483), .B2(n14893), .A(n14890), .ZN(n14906) );
  MUX2_X1 U15559 ( .A(P2_REG2_REG_13__SCAN_IN), .B(n13484), .S(n14903), .Z(
        n14905) );
  NAND2_X1 U15560 ( .A1(n14906), .A2(n14905), .ZN(n14904) );
  OAI21_X1 U15561 ( .B1(n13484), .B2(n13498), .A(n14904), .ZN(n13485) );
  NAND2_X1 U15562 ( .A1(n14918), .A2(n13485), .ZN(n13486) );
  XNOR2_X1 U15563 ( .A(n13485), .B(n13499), .ZN(n14914) );
  NAND2_X1 U15564 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n14914), .ZN(n14913) );
  NAND2_X1 U15565 ( .A1(n13486), .A2(n14913), .ZN(n13487) );
  NAND2_X1 U15566 ( .A1(n14923), .A2(n13487), .ZN(n13488) );
  XOR2_X1 U15567 ( .A(n14923), .B(n13487), .Z(n14925) );
  NAND2_X1 U15568 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n14925), .ZN(n14924) );
  NAND2_X1 U15569 ( .A1(n13488), .A2(n14924), .ZN(n14934) );
  NAND2_X1 U15570 ( .A1(n14933), .A2(n14934), .ZN(n14932) );
  OAI21_X1 U15571 ( .B1(n13504), .B2(n13489), .A(n14932), .ZN(n14949) );
  NAND2_X1 U15572 ( .A1(n14948), .A2(n14949), .ZN(n14947) );
  NAND2_X1 U15573 ( .A1(n13490), .A2(n14947), .ZN(n13491) );
  NOR2_X1 U15574 ( .A1(n14958), .A2(n13491), .ZN(n13492) );
  XNOR2_X1 U15575 ( .A(n13491), .B(n14958), .ZN(n14960) );
  NOR2_X1 U15576 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n14960), .ZN(n14962) );
  NOR2_X1 U15577 ( .A1(n13492), .A2(n14962), .ZN(n13493) );
  XNOR2_X1 U15578 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n13493), .ZN(n13513) );
  XNOR2_X1 U15579 ( .A(n13506), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n14945) );
  INV_X1 U15580 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n13503) );
  XOR2_X1 U15581 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n14935), .Z(n14937) );
  INV_X1 U15582 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n14747) );
  INV_X1 U15583 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n14754) );
  NAND2_X1 U15584 ( .A1(n13494), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n13495) );
  AND2_X1 U15585 ( .A1(n13496), .A2(n13495), .ZN(n14883) );
  MUX2_X1 U15586 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n14754), .S(n13497), .Z(
        n14882) );
  AND2_X1 U15587 ( .A1(n14883), .A2(n14882), .ZN(n14885) );
  AOI21_X1 U15588 ( .B1(n14754), .B2(n14893), .A(n14885), .ZN(n14909) );
  MUX2_X1 U15589 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n14747), .S(n14903), .Z(
        n14908) );
  NAND2_X1 U15590 ( .A1(n14909), .A2(n14908), .ZN(n14907) );
  OAI21_X1 U15591 ( .B1(n14747), .B2(n13498), .A(n14907), .ZN(n14917) );
  MUX2_X1 U15592 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n14739), .S(n14918), .Z(
        n14916) );
  NAND2_X1 U15593 ( .A1(n14917), .A2(n14916), .ZN(n14915) );
  OAI21_X1 U15594 ( .B1(n13499), .B2(n14739), .A(n14915), .ZN(n13500) );
  NAND2_X1 U15595 ( .A1(n14923), .A2(n13500), .ZN(n13502) );
  XNOR2_X1 U15596 ( .A(n13501), .B(n13500), .ZN(n14927) );
  NAND2_X1 U15597 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n14927), .ZN(n14926) );
  NAND2_X1 U15598 ( .A1(n13502), .A2(n14926), .ZN(n14938) );
  NAND2_X1 U15599 ( .A1(n14937), .A2(n14938), .ZN(n14936) );
  OAI21_X1 U15600 ( .B1(n13504), .B2(n13503), .A(n14936), .ZN(n14946) );
  NAND2_X1 U15601 ( .A1(n14945), .A2(n14946), .ZN(n14944) );
  OAI21_X1 U15602 ( .B1(n13506), .B2(n13505), .A(n14944), .ZN(n13508) );
  XNOR2_X1 U15603 ( .A(n13507), .B(n13508), .ZN(n14957) );
  NAND2_X1 U15604 ( .A1(P2_REG1_REG_18__SCAN_IN), .A2(n14957), .ZN(n14955) );
  NAND2_X1 U15605 ( .A1(n14958), .A2(n13508), .ZN(n13509) );
  NAND2_X1 U15606 ( .A1(n14955), .A2(n13509), .ZN(n13510) );
  XOR2_X1 U15607 ( .A(n13510), .B(P2_REG1_REG_19__SCAN_IN), .Z(n13515) );
  OAI21_X1 U15608 ( .B1(n13515), .B2(n13511), .A(n14894), .ZN(n13512) );
  AOI21_X1 U15609 ( .B1(n13513), .B2(n14961), .A(n13512), .ZN(n13518) );
  INV_X1 U15610 ( .A(n13513), .ZN(n13514) );
  AOI22_X1 U15611 ( .A1(n13515), .A2(n14956), .B1(n14961), .B2(n13514), .ZN(
        n13517) );
  MUX2_X1 U15612 ( .A(n13518), .B(n13517), .S(n13516), .Z(n13520) );
  OAI211_X1 U15613 ( .C1(n7496), .C2(n14901), .A(n13520), .B(n13519), .ZN(
        P2_U3233) );
  NAND2_X1 U15614 ( .A1(n13561), .A2(n13759), .ZN(n13531) );
  OAI21_X1 U15615 ( .B1(n13526), .B2(n13525), .A(n13524), .ZN(n13590) );
  NOR2_X1 U15616 ( .A1(n15005), .A2(n13757), .ZN(n13533) );
  NOR2_X1 U15617 ( .A1(n13522), .A2(n14968), .ZN(n13529) );
  AOI211_X1 U15618 ( .C1(P2_REG2_REG_31__SCAN_IN), .C2(n15005), .A(n13533), 
        .B(n13529), .ZN(n13530) );
  OAI21_X1 U15619 ( .B1(n14983), .B2(n13756), .A(n13530), .ZN(P2_U3234) );
  OAI211_X1 U15620 ( .C1(n13561), .C2(n13759), .A(n10086), .B(n13531), .ZN(
        n13758) );
  NOR2_X1 U15621 ( .A1(n13759), .A2(n14968), .ZN(n13532) );
  AOI211_X1 U15622 ( .C1(n15005), .C2(P2_REG2_REG_30__SCAN_IN), .A(n13533), 
        .B(n13532), .ZN(n13534) );
  OAI21_X1 U15623 ( .B1(n14983), .B2(n13758), .A(n13534), .ZN(P2_U3235) );
  NAND2_X1 U15624 ( .A1(n13712), .A2(n6559), .ZN(n13542) );
  NAND2_X1 U15625 ( .A1(n13722), .A2(n13540), .ZN(n13541) );
  NAND2_X1 U15626 ( .A1(n13699), .A2(n13578), .ZN(n13543) );
  NAND2_X1 U15627 ( .A1(n13811), .A2(n13545), .ZN(n13546) );
  INV_X1 U15628 ( .A(n13806), .ZN(n13679) );
  INV_X1 U15629 ( .A(n13580), .ZN(n13547) );
  NAND2_X1 U15630 ( .A1(n13679), .A2(n13547), .ZN(n13548) );
  NAND2_X1 U15631 ( .A1(n13795), .A2(n13550), .ZN(n13551) );
  INV_X1 U15632 ( .A(n13628), .ZN(n13555) );
  INV_X1 U15633 ( .A(n13635), .ZN(n13785) );
  NOR2_X1 U15634 ( .A1(n13785), .A2(n13556), .ZN(n13553) );
  INV_X1 U15635 ( .A(n13553), .ZN(n13554) );
  NAND2_X1 U15636 ( .A1(n13785), .A2(n13556), .ZN(n13557) );
  INV_X1 U15637 ( .A(n13587), .ZN(n13604) );
  NAND2_X1 U15638 ( .A1(n13603), .A2(n13558), .ZN(n13560) );
  INV_X1 U15639 ( .A(n13588), .ZN(n13559) );
  XNOR2_X1 U15640 ( .A(n13560), .B(n13559), .ZN(n13760) );
  INV_X1 U15641 ( .A(n13760), .ZN(n13597) );
  AOI211_X1 U15642 ( .C1(n13763), .C2(n13606), .A(n12610), .B(n13561), .ZN(
        n13762) );
  INV_X1 U15643 ( .A(n13562), .ZN(n13563) );
  AOI22_X1 U15644 ( .A1(n13563), .A2(n14979), .B1(P2_REG2_REG_29__SCAN_IN), 
        .B2(n15005), .ZN(n13564) );
  OAI21_X1 U15645 ( .B1(n13764), .B2(n14968), .A(n13564), .ZN(n13565) );
  AOI21_X1 U15646 ( .B1(n13762), .B2(n14722), .A(n13565), .ZN(n13596) );
  NAND2_X1 U15647 ( .A1(n13833), .A2(n13566), .ZN(n13574) );
  INV_X1 U15648 ( .A(n13567), .ZN(n13568) );
  NAND2_X1 U15649 ( .A1(n13569), .A2(n13568), .ZN(n13571) );
  NOR2_X1 U15650 ( .A1(n13569), .A2(n13568), .ZN(n13570) );
  INV_X1 U15651 ( .A(n13576), .ZN(n13577) );
  INV_X1 U15652 ( .A(n13669), .ZN(n13672) );
  NAND2_X1 U15653 ( .A1(n13795), .A2(n13581), .ZN(n13646) );
  INV_X1 U15654 ( .A(n13585), .ZN(n13586) );
  NAND2_X1 U15655 ( .A1(n13598), .A2(n13587), .ZN(n13601) );
  OAI22_X1 U15656 ( .A1(n13592), .A2(n13591), .B1(n13590), .B2(n13589), .ZN(
        n13593) );
  INV_X1 U15657 ( .A(n13593), .ZN(n13594) );
  NAND2_X1 U15658 ( .A1(n13761), .A2(n15002), .ZN(n13595) );
  OAI211_X1 U15659 ( .C1(n13597), .C2(n13739), .A(n13596), .B(n13595), .ZN(
        P2_U3236) );
  INV_X1 U15660 ( .A(n13598), .ZN(n13599) );
  AOI21_X1 U15661 ( .B1(n13599), .B2(n13604), .A(n14997), .ZN(n13602) );
  INV_X1 U15662 ( .A(n13768), .ZN(n13613) );
  OAI211_X1 U15663 ( .C1(n13620), .C2(n13607), .A(n10086), .B(n13606), .ZN(
        n13771) );
  INV_X1 U15664 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n13608) );
  OAI22_X1 U15665 ( .A1(n13609), .A2(n14996), .B1(n13608), .B2(n15002), .ZN(
        n13610) );
  AOI21_X1 U15666 ( .B1(n13769), .B2(n14715), .A(n13610), .ZN(n13611) );
  OAI21_X1 U15667 ( .B1(n13771), .B2(n14983), .A(n13611), .ZN(n13612) );
  AOI21_X1 U15668 ( .B1(n13613), .B2(n14723), .A(n13612), .ZN(n13614) );
  OAI21_X1 U15669 ( .B1(n15005), .B2(n13773), .A(n13614), .ZN(P2_U3237) );
  XOR2_X1 U15670 ( .A(n13615), .B(n13617), .Z(n13782) );
  NAND2_X1 U15671 ( .A1(n13616), .A2(n13617), .ZN(n13775) );
  NAND3_X1 U15672 ( .A1(n13776), .A2(n13775), .A3(n14723), .ZN(n13627) );
  NAND2_X1 U15673 ( .A1(n13630), .A2(n13779), .ZN(n13618) );
  NAND2_X1 U15674 ( .A1(n13618), .A2(n10086), .ZN(n13619) );
  NOR2_X1 U15675 ( .A1(n13620), .A2(n13619), .ZN(n13777) );
  INV_X1 U15676 ( .A(n13621), .ZN(n13622) );
  AOI22_X1 U15677 ( .A1(n13622), .A2(n14979), .B1(P2_REG2_REG_27__SCAN_IN), 
        .B2(n15005), .ZN(n13624) );
  NAND2_X1 U15678 ( .A1(n13778), .A2(n15002), .ZN(n13623) );
  OAI211_X1 U15679 ( .C1(n6944), .C2(n14968), .A(n13624), .B(n13623), .ZN(
        n13625) );
  AOI21_X1 U15680 ( .B1(n13777), .B2(n14722), .A(n13625), .ZN(n13626) );
  OAI211_X1 U15681 ( .C1(n13782), .C2(n13755), .A(n13627), .B(n13626), .ZN(
        P2_U3238) );
  XNOR2_X1 U15682 ( .A(n13628), .B(n13629), .ZN(n13789) );
  XNOR2_X1 U15683 ( .A(n6535), .B(n13629), .ZN(n13787) );
  AOI21_X1 U15684 ( .B1(n13642), .B2(n13635), .A(n12610), .ZN(n13631) );
  NAND2_X1 U15685 ( .A1(n13631), .A2(n13630), .ZN(n13784) );
  AOI22_X1 U15686 ( .A1(n13632), .A2(n14979), .B1(P2_REG2_REG_26__SCAN_IN), 
        .B2(n15005), .ZN(n13633) );
  OAI21_X1 U15687 ( .B1(n13783), .B2(n15005), .A(n13633), .ZN(n13634) );
  AOI21_X1 U15688 ( .B1(n13635), .B2(n14715), .A(n13634), .ZN(n13636) );
  OAI21_X1 U15689 ( .B1(n13784), .B2(n14983), .A(n13636), .ZN(n13637) );
  AOI21_X1 U15690 ( .B1(n13787), .B2(n13737), .A(n13637), .ZN(n13638) );
  OAI21_X1 U15691 ( .B1(n13789), .B2(n13739), .A(n13638), .ZN(P2_U3239) );
  XNOR2_X1 U15692 ( .A(n13639), .B(n13647), .ZN(n13794) );
  OR2_X1 U15693 ( .A1(n13657), .A2(n13640), .ZN(n13641) );
  AND3_X1 U15694 ( .A1(n13642), .A2(n10086), .A3(n13641), .ZN(n13790) );
  NAND2_X1 U15695 ( .A1(n13791), .A2(n14715), .ZN(n13644) );
  NAND2_X1 U15696 ( .A1(n15005), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n13643) );
  OAI211_X1 U15697 ( .C1(n14996), .C2(n13645), .A(n13644), .B(n13643), .ZN(
        n13652) );
  NAND3_X1 U15698 ( .A1(n13664), .A2(n13647), .A3(n13646), .ZN(n13648) );
  AOI21_X1 U15699 ( .B1(n6564), .B2(n13648), .A(n14997), .ZN(n13650) );
  NOR2_X1 U15700 ( .A1(n13650), .A2(n13649), .ZN(n13793) );
  NOR2_X1 U15701 ( .A1(n13793), .A2(n15005), .ZN(n13651) );
  AOI211_X1 U15702 ( .C1(n13790), .C2(n14722), .A(n13652), .B(n13651), .ZN(
        n13653) );
  OAI21_X1 U15703 ( .B1(n13794), .B2(n13739), .A(n13653), .ZN(P2_U3240) );
  OAI21_X1 U15704 ( .B1(n6517), .B2(n13549), .A(n13654), .ZN(n13802) );
  NAND2_X1 U15705 ( .A1(n13673), .A2(n13795), .ZN(n13655) );
  NAND2_X1 U15706 ( .A1(n13655), .A2(n10086), .ZN(n13656) );
  NOR2_X1 U15707 ( .A1(n13657), .A2(n13656), .ZN(n13799) );
  NAND2_X1 U15708 ( .A1(n13795), .A2(n14715), .ZN(n13662) );
  NOR2_X1 U15709 ( .A1(n15002), .A2(n13658), .ZN(n13659) );
  AOI21_X1 U15710 ( .B1(n13660), .B2(n14979), .A(n13659), .ZN(n13661) );
  OAI211_X1 U15711 ( .C1(n15005), .C2(n13796), .A(n13662), .B(n13661), .ZN(
        n13663) );
  AOI21_X1 U15712 ( .B1(n13799), .B2(n14722), .A(n13663), .ZN(n13668) );
  OAI21_X1 U15713 ( .B1(n13666), .B2(n13665), .A(n13664), .ZN(n13800) );
  NAND2_X1 U15714 ( .A1(n13800), .A2(n13737), .ZN(n13667) );
  OAI211_X1 U15715 ( .C1(n13802), .C2(n13739), .A(n13668), .B(n13667), .ZN(
        P2_U3241) );
  XNOR2_X1 U15716 ( .A(n13670), .B(n13669), .ZN(n13809) );
  OAI21_X1 U15717 ( .B1(n6562), .B2(n13672), .A(n13671), .ZN(n13803) );
  NAND2_X1 U15718 ( .A1(n13803), .A2(n14723), .ZN(n13682) );
  INV_X1 U15719 ( .A(n13673), .ZN(n13674) );
  AOI211_X1 U15720 ( .C1(n13806), .C2(n13689), .A(n12610), .B(n13674), .ZN(
        n13804) );
  INV_X1 U15721 ( .A(n13675), .ZN(n13676) );
  AOI22_X1 U15722 ( .A1(n13676), .A2(n14979), .B1(n15005), .B2(
        P2_REG2_REG_23__SCAN_IN), .ZN(n13678) );
  NAND2_X1 U15723 ( .A1(n13805), .A2(n15002), .ZN(n13677) );
  OAI211_X1 U15724 ( .C1(n13679), .C2(n14968), .A(n13678), .B(n13677), .ZN(
        n13680) );
  AOI21_X1 U15725 ( .B1(n13804), .B2(n14722), .A(n13680), .ZN(n13681) );
  OAI211_X1 U15726 ( .C1(n13809), .C2(n13755), .A(n13682), .B(n13681), .ZN(
        P2_U3242) );
  OAI211_X1 U15727 ( .C1(n13684), .C2(n13687), .A(n13683), .B(n15064), .ZN(
        n13686) );
  OAI21_X1 U15728 ( .B1(n6561), .B2(n7402), .A(n13688), .ZN(n13814) );
  INV_X1 U15729 ( .A(n13814), .ZN(n13696) );
  AOI21_X1 U15730 ( .B1(n13811), .B2(n13701), .A(n12610), .ZN(n13690) );
  AND2_X1 U15731 ( .A1(n13690), .A2(n13689), .ZN(n13810) );
  NAND2_X1 U15732 ( .A1(n13810), .A2(n14722), .ZN(n13693) );
  AOI22_X1 U15733 ( .A1(n15005), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n13691), 
        .B2(n14979), .ZN(n13692) );
  OAI211_X1 U15734 ( .C1(n13694), .C2(n14968), .A(n13693), .B(n13692), .ZN(
        n13695) );
  AOI21_X1 U15735 ( .B1(n13696), .B2(n14723), .A(n13695), .ZN(n13697) );
  OAI21_X1 U15736 ( .B1(n15005), .B2(n13813), .A(n13697), .ZN(P2_U3243) );
  XOR2_X1 U15737 ( .A(n13698), .B(n13706), .Z(n13819) );
  OR2_X1 U15738 ( .A1(n13718), .A2(n13699), .ZN(n13700) );
  AND3_X1 U15739 ( .A1(n13701), .A2(n10086), .A3(n13700), .ZN(n13816) );
  NAND2_X1 U15740 ( .A1(n13817), .A2(n14715), .ZN(n13703) );
  NAND2_X1 U15741 ( .A1(n15005), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n13702) );
  OAI211_X1 U15742 ( .C1(n14996), .C2(n13704), .A(n13703), .B(n13702), .ZN(
        n13705) );
  AOI21_X1 U15743 ( .B1(n13816), .B2(n14722), .A(n13705), .ZN(n13711) );
  AOI21_X1 U15744 ( .B1(n13707), .B2(n13706), .A(n6581), .ZN(n13709) );
  OAI21_X1 U15745 ( .B1(n13709), .B2(n14997), .A(n13708), .ZN(n13815) );
  NAND2_X1 U15746 ( .A1(n13815), .A2(n15002), .ZN(n13710) );
  OAI211_X1 U15747 ( .C1(n13819), .C2(n13739), .A(n13711), .B(n13710), .ZN(
        P2_U3244) );
  XOR2_X1 U15748 ( .A(n13712), .B(n13715), .Z(n13824) );
  AOI21_X1 U15749 ( .B1(n13715), .B2(n13714), .A(n13713), .ZN(n13717) );
  OAI21_X1 U15750 ( .B1(n13717), .B2(n14997), .A(n13716), .ZN(n13820) );
  AOI211_X1 U15751 ( .C1(n13822), .C2(n13729), .A(n12610), .B(n13718), .ZN(
        n13821) );
  NAND2_X1 U15752 ( .A1(n13821), .A2(n14722), .ZN(n13721) );
  AOI22_X1 U15753 ( .A1(n15005), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n13719), 
        .B2(n14979), .ZN(n13720) );
  OAI211_X1 U15754 ( .C1(n13722), .C2(n14968), .A(n13721), .B(n13720), .ZN(
        n13723) );
  AOI21_X1 U15755 ( .B1(n13820), .B2(n15002), .A(n13723), .ZN(n13724) );
  OAI21_X1 U15756 ( .B1(n13824), .B2(n13739), .A(n13724), .ZN(P2_U3245) );
  XNOR2_X1 U15757 ( .A(n13725), .B(n13727), .ZN(n13830) );
  XOR2_X1 U15758 ( .A(n13727), .B(n13726), .Z(n13828) );
  NAND2_X1 U15759 ( .A1(n13734), .A2(n13746), .ZN(n13728) );
  NAND3_X1 U15760 ( .A1(n13729), .A2(n10086), .A3(n13728), .ZN(n13826) );
  OR2_X1 U15761 ( .A1(n14996), .A2(n13730), .ZN(n13732) );
  NAND2_X1 U15762 ( .A1(n15005), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n13731) );
  OAI211_X1 U15763 ( .C1(n13825), .C2(n15005), .A(n13732), .B(n13731), .ZN(
        n13733) );
  AOI21_X1 U15764 ( .B1(n13734), .B2(n14715), .A(n13733), .ZN(n13735) );
  OAI21_X1 U15765 ( .B1(n13826), .B2(n14983), .A(n13735), .ZN(n13736) );
  AOI21_X1 U15766 ( .B1(n13828), .B2(n13737), .A(n13736), .ZN(n13738) );
  OAI21_X1 U15767 ( .B1(n13830), .B2(n13739), .A(n13738), .ZN(P2_U3246) );
  XNOR2_X1 U15768 ( .A(n13740), .B(n13742), .ZN(n13837) );
  OAI21_X1 U15769 ( .B1(n13743), .B2(n13742), .A(n13741), .ZN(n13835) );
  AOI21_X1 U15770 ( .B1(n13745), .B2(n13744), .A(n12610), .ZN(n13747) );
  NAND2_X1 U15771 ( .A1(n13747), .A2(n13746), .ZN(n13832) );
  INV_X1 U15772 ( .A(n13748), .ZN(n13749) );
  OAI22_X1 U15773 ( .A1(n15005), .A2(n13831), .B1(n13749), .B2(n14996), .ZN(
        n13751) );
  NOR2_X1 U15774 ( .A1(n13833), .A2(n14968), .ZN(n13750) );
  AOI211_X1 U15775 ( .C1(n15005), .C2(P2_REG2_REG_18__SCAN_IN), .A(n13751), 
        .B(n13750), .ZN(n13752) );
  OAI21_X1 U15776 ( .B1(n14983), .B2(n13832), .A(n13752), .ZN(n13753) );
  AOI21_X1 U15777 ( .B1(n13835), .B2(n14723), .A(n13753), .ZN(n13754) );
  OAI21_X1 U15778 ( .B1(n13755), .B2(n13837), .A(n13754), .ZN(P2_U3247) );
  OAI211_X1 U15779 ( .C1(n13522), .C2(n15077), .A(n13756), .B(n13757), .ZN(
        n13846) );
  MUX2_X1 U15780 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n13846), .S(n15096), .Z(
        P2_U3530) );
  OAI211_X1 U15781 ( .C1(n13759), .C2(n15077), .A(n13758), .B(n13757), .ZN(
        n13847) );
  MUX2_X1 U15782 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n13847), .S(n15096), .Z(
        P2_U3529) );
  NAND2_X1 U15783 ( .A1(n13760), .A2(n15035), .ZN(n13767) );
  INV_X1 U15784 ( .A(n13762), .ZN(n13765) );
  INV_X1 U15785 ( .A(n13763), .ZN(n13764) );
  NAND2_X1 U15786 ( .A1(n13767), .A2(n7446), .ZN(n13848) );
  MUX2_X1 U15787 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n13848), .S(n15096), .Z(
        P2_U3528) );
  NAND2_X1 U15788 ( .A1(n13769), .A2(n15069), .ZN(n13770) );
  NAND3_X1 U15789 ( .A1(n13776), .A2(n13775), .A3(n15035), .ZN(n13781) );
  AOI211_X1 U15790 ( .C1(n15069), .C2(n13779), .A(n13778), .B(n13777), .ZN(
        n13780) );
  OAI211_X1 U15791 ( .C1(n14997), .C2(n13782), .A(n13781), .B(n13780), .ZN(
        n13850) );
  MUX2_X1 U15792 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n13850), .S(n15096), .Z(
        P2_U3526) );
  OAI211_X1 U15793 ( .C1(n13785), .C2(n15077), .A(n13784), .B(n13783), .ZN(
        n13786) );
  AOI21_X1 U15794 ( .B1(n13787), .B2(n15064), .A(n13786), .ZN(n13788) );
  MUX2_X1 U15795 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n13851), .S(n15096), .Z(
        P2_U3525) );
  AOI21_X1 U15796 ( .B1(n15069), .B2(n13791), .A(n13790), .ZN(n13792) );
  OAI211_X1 U15797 ( .C1(n13794), .C2(n15061), .A(n13793), .B(n13792), .ZN(
        n13852) );
  MUX2_X1 U15798 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n13852), .S(n15096), .Z(
        P2_U3524) );
  INV_X1 U15799 ( .A(n13795), .ZN(n13797) );
  OAI21_X1 U15800 ( .B1(n13797), .B2(n15077), .A(n13796), .ZN(n13798) );
  AOI211_X1 U15801 ( .C1(n13800), .C2(n15064), .A(n13799), .B(n13798), .ZN(
        n13801) );
  OAI21_X1 U15802 ( .B1(n13802), .B2(n15061), .A(n13801), .ZN(n13853) );
  MUX2_X1 U15803 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n13853), .S(n15096), .Z(
        P2_U3523) );
  NAND2_X1 U15804 ( .A1(n13803), .A2(n15035), .ZN(n13808) );
  AOI211_X1 U15805 ( .C1(n15069), .C2(n13806), .A(n13805), .B(n13804), .ZN(
        n13807) );
  OAI211_X1 U15806 ( .C1(n14997), .C2(n13809), .A(n13808), .B(n13807), .ZN(
        n13854) );
  MUX2_X1 U15807 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n13854), .S(n15096), .Z(
        P2_U3522) );
  AOI21_X1 U15808 ( .B1(n15069), .B2(n13811), .A(n13810), .ZN(n13812) );
  OAI211_X1 U15809 ( .C1(n13814), .C2(n15061), .A(n13813), .B(n13812), .ZN(
        n13855) );
  MUX2_X1 U15810 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n13855), .S(n15096), .Z(
        P2_U3521) );
  AOI211_X1 U15811 ( .C1(n15069), .C2(n13817), .A(n13816), .B(n13815), .ZN(
        n13818) );
  OAI21_X1 U15812 ( .B1(n13819), .B2(n15061), .A(n13818), .ZN(n13856) );
  MUX2_X1 U15813 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n13856), .S(n15096), .Z(
        P2_U3520) );
  AOI211_X1 U15814 ( .C1(n15069), .C2(n13822), .A(n13821), .B(n13820), .ZN(
        n13823) );
  OAI21_X1 U15815 ( .B1(n13824), .B2(n15061), .A(n13823), .ZN(n13857) );
  MUX2_X1 U15816 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n13857), .S(n15096), .Z(
        P2_U3519) );
  OAI211_X1 U15817 ( .C1(n6703), .C2(n15077), .A(n13826), .B(n13825), .ZN(
        n13827) );
  AOI21_X1 U15818 ( .B1(n13828), .B2(n15064), .A(n13827), .ZN(n13829) );
  OAI21_X1 U15819 ( .B1(n13830), .B2(n15061), .A(n13829), .ZN(n13858) );
  MUX2_X1 U15820 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n13858), .S(n15096), .Z(
        P2_U3518) );
  OAI211_X1 U15821 ( .C1(n13833), .C2(n15077), .A(n13832), .B(n13831), .ZN(
        n13834) );
  AOI21_X1 U15822 ( .B1(n13835), .B2(n15035), .A(n13834), .ZN(n13836) );
  OAI21_X1 U15823 ( .B1(n14997), .B2(n13837), .A(n13836), .ZN(n13859) );
  MUX2_X1 U15824 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n13859), .S(n15096), .Z(
        P2_U3517) );
  OAI211_X1 U15825 ( .C1(n13840), .C2(n15077), .A(n13839), .B(n13838), .ZN(
        n13841) );
  AOI21_X1 U15826 ( .B1(n13842), .B2(n15035), .A(n13841), .ZN(n13843) );
  OAI21_X1 U15827 ( .B1(n14997), .B2(n13844), .A(n13843), .ZN(n13860) );
  MUX2_X1 U15828 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n13860), .S(n15096), .Z(
        P2_U3516) );
  MUX2_X1 U15829 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n13845), .S(n15096), .Z(
        P2_U3505) );
  MUX2_X1 U15830 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n13846), .S(n15066), .Z(
        P2_U3498) );
  MUX2_X1 U15831 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n13847), .S(n15066), .Z(
        P2_U3497) );
  MUX2_X1 U15832 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n13848), .S(n15066), .Z(
        P2_U3496) );
  MUX2_X1 U15833 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n13849), .S(n15066), .Z(
        P2_U3495) );
  MUX2_X1 U15834 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n13850), .S(n15066), .Z(
        P2_U3494) );
  MUX2_X1 U15835 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n13852), .S(n15066), .Z(
        P2_U3492) );
  MUX2_X1 U15836 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n13853), .S(n15066), .Z(
        P2_U3491) );
  MUX2_X1 U15837 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n13854), .S(n15066), .Z(
        P2_U3490) );
  MUX2_X1 U15838 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n13855), .S(n15066), .Z(
        P2_U3489) );
  MUX2_X1 U15839 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n13856), .S(n15066), .Z(
        P2_U3488) );
  MUX2_X1 U15840 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n13857), .S(n15066), .Z(
        P2_U3487) );
  MUX2_X1 U15841 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n13858), .S(n15066), .Z(
        P2_U3486) );
  MUX2_X1 U15842 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n13859), .S(n15066), .Z(
        P2_U3484) );
  MUX2_X1 U15843 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n13860), .S(n15066), .Z(
        P2_U3481) );
  INV_X1 U15844 ( .A(n13861), .ZN(n14475) );
  NAND3_X1 U15845 ( .A1(n8565), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_STATE_REG_SCAN_IN), .ZN(n13863) );
  OAI22_X1 U15846 ( .A1(n8567), .A2(n13863), .B1(n13862), .B2(n13870), .ZN(
        n13864) );
  INV_X1 U15847 ( .A(n13864), .ZN(n13865) );
  OAI21_X1 U15848 ( .B1(n14475), .B2(n13873), .A(n13865), .ZN(P2_U3296) );
  INV_X1 U15849 ( .A(n13869), .ZN(n14479) );
  OAI222_X1 U15850 ( .A1(n13873), .A2(n14479), .B1(P2_U3088), .B2(n13872), 
        .C1(n13871), .C2(n13870), .ZN(P2_U3298) );
  MUX2_X1 U15851 ( .A(n13874), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3327) );
  XOR2_X1 U15852 ( .A(n13876), .B(n13875), .Z(n13882) );
  NOR2_X1 U15853 ( .A1(n13989), .A2(n14159), .ZN(n13880) );
  AOI22_X1 U15854 ( .A1(n14011), .A2(n14147), .B1(P1_REG3_REG_27__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13877) );
  OAI21_X1 U15855 ( .B1(n13878), .B2(n14013), .A(n13877), .ZN(n13879) );
  AOI211_X1 U15856 ( .C1(n14158), .C2(n14018), .A(n13880), .B(n13879), .ZN(
        n13881) );
  OAI21_X1 U15857 ( .B1(n13882), .B2(n14022), .A(n13881), .ZN(P1_U3214) );
  INV_X1 U15858 ( .A(n13883), .ZN(n13884) );
  AOI21_X1 U15859 ( .B1(n13886), .B2(n13885), .A(n13884), .ZN(n13894) );
  NAND2_X1 U15860 ( .A1(n13999), .A2(n13887), .ZN(n13888) );
  OAI211_X1 U15861 ( .C1(n13989), .C2(n13890), .A(n13889), .B(n13888), .ZN(
        n13891) );
  AOI21_X1 U15862 ( .B1(n13892), .B2(n14018), .A(n13891), .ZN(n13893) );
  OAI21_X1 U15863 ( .B1(n13894), .B2(n14022), .A(n13893), .ZN(P1_U3215) );
  XOR2_X1 U15864 ( .A(n13896), .B(n13895), .Z(n13902) );
  NAND2_X1 U15865 ( .A1(n14027), .A2(n14319), .ZN(n13898) );
  NAND2_X1 U15866 ( .A1(n14026), .A2(n14321), .ZN(n13897) );
  NAND2_X1 U15867 ( .A1(n13898), .A2(n13897), .ZN(n14231) );
  AOI22_X1 U15868 ( .A1(n14231), .A2(n13999), .B1(P1_REG3_REG_23__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13899) );
  OAI21_X1 U15869 ( .B1(n13989), .B2(n14239), .A(n13899), .ZN(n13900) );
  AOI21_X1 U15870 ( .B1(n14385), .B2(n14018), .A(n13900), .ZN(n13901) );
  OAI21_X1 U15871 ( .B1(n13902), .B2(n14022), .A(n13901), .ZN(P1_U3216) );
  AOI21_X1 U15872 ( .B1(n13904), .B2(n13903), .A(n14022), .ZN(n13905) );
  OR2_X1 U15873 ( .A1(n13904), .A2(n13903), .ZN(n13960) );
  NAND2_X1 U15874 ( .A1(n13905), .A2(n13960), .ZN(n13910) );
  OAI22_X1 U15875 ( .A1(n14264), .A2(n14287), .B1(n13906), .B2(n14285), .ZN(
        n14305) );
  NOR2_X1 U15876 ( .A1(n13989), .A2(n14308), .ZN(n13907) );
  AOI211_X1 U15877 ( .C1(n13999), .C2(n14305), .A(n13908), .B(n13907), .ZN(
        n13909) );
  OAI211_X1 U15878 ( .C1(n9549), .C2(n13980), .A(n13910), .B(n13909), .ZN(
        P1_U3219) );
  INV_X1 U15879 ( .A(n13911), .ZN(n13912) );
  AOI21_X1 U15880 ( .B1(n13914), .B2(n13913), .A(n13912), .ZN(n13921) );
  NOR2_X1 U15881 ( .A1(n13915), .A2(P1_STATE_REG_SCAN_IN), .ZN(n13916) );
  AOI21_X1 U15882 ( .B1(n14027), .B2(n13987), .A(n13916), .ZN(n13918) );
  NAND2_X1 U15883 ( .A1(n14011), .A2(n14028), .ZN(n13917) );
  OAI211_X1 U15884 ( .C1(n13989), .C2(n14272), .A(n13918), .B(n13917), .ZN(
        n13919) );
  AOI21_X1 U15885 ( .B1(n14271), .B2(n14018), .A(n13919), .ZN(n13920) );
  OAI21_X1 U15886 ( .B1(n13921), .B2(n14022), .A(n13920), .ZN(P1_U3223) );
  NAND2_X1 U15887 ( .A1(n13923), .A2(n13922), .ZN(n13924) );
  XOR2_X1 U15888 ( .A(n13925), .B(n13924), .Z(n13931) );
  NAND2_X1 U15889 ( .A1(n14026), .A2(n14319), .ZN(n13927) );
  NAND2_X1 U15890 ( .A1(n14147), .A2(n14321), .ZN(n13926) );
  NAND2_X1 U15891 ( .A1(n13927), .A2(n13926), .ZN(n14189) );
  AOI22_X1 U15892 ( .A1(n13999), .A2(n14189), .B1(P1_REG3_REG_25__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13928) );
  OAI21_X1 U15893 ( .B1(n13989), .B2(n14198), .A(n13928), .ZN(n13929) );
  AOI21_X1 U15894 ( .B1(n14374), .B2(n14018), .A(n13929), .ZN(n13930) );
  OAI21_X1 U15895 ( .B1(n13931), .B2(n14022), .A(n13930), .ZN(P1_U3225) );
  XOR2_X1 U15896 ( .A(n13933), .B(n13932), .Z(n13941) );
  INV_X1 U15897 ( .A(n13999), .ZN(n13937) );
  NAND2_X1 U15898 ( .A1(n14016), .A2(n13934), .ZN(n13936) );
  OAI211_X1 U15899 ( .C1(n13938), .C2(n13937), .A(n13936), .B(n13935), .ZN(
        n13939) );
  AOI21_X1 U15900 ( .B1(n14425), .B2(n14018), .A(n13939), .ZN(n13940) );
  OAI21_X1 U15901 ( .B1(n13941), .B2(n14022), .A(n13940), .ZN(P1_U3226) );
  XOR2_X1 U15902 ( .A(n13943), .B(n13942), .Z(n13951) );
  OAI21_X1 U15903 ( .B1(n13985), .B2(n14014), .A(n13944), .ZN(n13945) );
  AOI21_X1 U15904 ( .B1(n13987), .B2(n14029), .A(n13945), .ZN(n13946) );
  OAI21_X1 U15905 ( .B1(n13989), .B2(n13947), .A(n13946), .ZN(n13948) );
  AOI21_X1 U15906 ( .B1(n13949), .B2(n14018), .A(n13948), .ZN(n13950) );
  OAI21_X1 U15907 ( .B1(n13951), .B2(n14022), .A(n13950), .ZN(P1_U3228) );
  XOR2_X1 U15908 ( .A(n13953), .B(n13952), .Z(n13958) );
  NOR2_X1 U15909 ( .A1(n13989), .A2(n14222), .ZN(n13956) );
  AOI22_X1 U15910 ( .A1(n14249), .A2(n14011), .B1(P1_REG3_REG_24__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13954) );
  OAI21_X1 U15911 ( .B1(n14213), .B2(n14013), .A(n13954), .ZN(n13955) );
  AOI211_X1 U15912 ( .C1(n14377), .C2(n14018), .A(n13956), .B(n13955), .ZN(
        n13957) );
  OAI21_X1 U15913 ( .B1(n13958), .B2(n14022), .A(n13957), .ZN(P1_U3229) );
  INV_X1 U15914 ( .A(n14404), .ZN(n14296) );
  NAND2_X1 U15915 ( .A1(n13960), .A2(n13959), .ZN(n13965) );
  AND2_X1 U15916 ( .A1(n13962), .A2(n13961), .ZN(n13963) );
  OAI211_X1 U15917 ( .C1(n13965), .C2(n13964), .A(n13963), .B(n13995), .ZN(
        n13970) );
  OAI22_X1 U15918 ( .A1(n14288), .A2(n14013), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13966), .ZN(n13968) );
  NOR2_X1 U15919 ( .A1(n13989), .A2(n14292), .ZN(n13967) );
  AOI211_X1 U15920 ( .C1(n14011), .C2(n14322), .A(n13968), .B(n13967), .ZN(
        n13969) );
  OAI211_X1 U15921 ( .C1(n14296), .C2(n13980), .A(n13970), .B(n13969), .ZN(
        P1_U3233) );
  OAI21_X1 U15922 ( .B1(n13973), .B2(n13972), .A(n13971), .ZN(n13974) );
  NAND2_X1 U15923 ( .A1(n13974), .A2(n13995), .ZN(n13979) );
  INV_X1 U15924 ( .A(n13975), .ZN(n14256) );
  AOI22_X1 U15925 ( .A1(n14249), .A2(n13987), .B1(P1_REG3_REG_22__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13976) );
  OAI21_X1 U15926 ( .B1(n14288), .B2(n13985), .A(n13976), .ZN(n13977) );
  AOI21_X1 U15927 ( .B1(n14256), .B2(n14016), .A(n13977), .ZN(n13978) );
  OAI211_X1 U15928 ( .C1(n13980), .C2(n14259), .A(n13979), .B(n13978), .ZN(
        P1_U3235) );
  XOR2_X1 U15929 ( .A(n13982), .B(n13981), .Z(n13992) );
  OAI21_X1 U15930 ( .B1(n13985), .B2(n13984), .A(n13983), .ZN(n13986) );
  AOI21_X1 U15931 ( .B1(n13987), .B2(n14322), .A(n13986), .ZN(n13988) );
  OAI21_X1 U15932 ( .B1(n13989), .B2(n14328), .A(n13988), .ZN(n13990) );
  AOI21_X1 U15933 ( .B1(n14414), .B2(n14018), .A(n13990), .ZN(n13991) );
  OAI21_X1 U15934 ( .B1(n13992), .B2(n14022), .A(n13991), .ZN(P1_U3238) );
  XOR2_X1 U15935 ( .A(n13994), .B(n13993), .Z(n13996) );
  NAND2_X1 U15936 ( .A1(n13996), .A2(n13995), .ZN(n14006) );
  AOI21_X1 U15937 ( .B1(n13999), .B2(n13998), .A(n13997), .ZN(n14005) );
  INV_X1 U15938 ( .A(n14000), .ZN(n14001) );
  NAND2_X1 U15939 ( .A1(n14016), .A2(n14001), .ZN(n14004) );
  NAND2_X1 U15940 ( .A1(n14018), .A2(n14002), .ZN(n14003) );
  NAND4_X1 U15941 ( .A1(n14006), .A2(n14005), .A3(n14004), .A4(n14003), .ZN(
        P1_U3239) );
  NAND2_X1 U15942 ( .A1(n14008), .A2(n14007), .ZN(n14010) );
  XNOR2_X1 U15943 ( .A(n14010), .B(n14009), .ZN(n14023) );
  NAND2_X1 U15944 ( .A1(n14011), .A2(n14031), .ZN(n14012) );
  NAND2_X1 U15945 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n14813)
         );
  OAI211_X1 U15946 ( .C1(n14014), .C2(n14013), .A(n14012), .B(n14813), .ZN(
        n14015) );
  AOI21_X1 U15947 ( .B1(n14017), .B2(n14016), .A(n14015), .ZN(n14021) );
  NAND2_X1 U15948 ( .A1(n14019), .A2(n14018), .ZN(n14020) );
  OAI211_X1 U15949 ( .C1(n14023), .C2(n14022), .A(n14021), .B(n14020), .ZN(
        P1_U3241) );
  MUX2_X1 U15950 ( .A(n14024), .B(P1_DATAO_REG_31__SCAN_IN), .S(n14044), .Z(
        P1_U3591) );
  MUX2_X1 U15951 ( .A(n14025), .B(P1_DATAO_REG_30__SCAN_IN), .S(n14044), .Z(
        P1_U3590) );
  MUX2_X1 U15952 ( .A(n14131), .B(P1_DATAO_REG_29__SCAN_IN), .S(n14044), .Z(
        P1_U3589) );
  MUX2_X1 U15953 ( .A(n14146), .B(P1_DATAO_REG_28__SCAN_IN), .S(n14044), .Z(
        P1_U3588) );
  MUX2_X1 U15954 ( .A(n14175), .B(P1_DATAO_REG_27__SCAN_IN), .S(n14044), .Z(
        P1_U3587) );
  MUX2_X1 U15955 ( .A(n14174), .B(P1_DATAO_REG_25__SCAN_IN), .S(n14044), .Z(
        P1_U3585) );
  MUX2_X1 U15956 ( .A(n14026), .B(P1_DATAO_REG_24__SCAN_IN), .S(n14044), .Z(
        P1_U3584) );
  MUX2_X1 U15957 ( .A(n14249), .B(P1_DATAO_REG_23__SCAN_IN), .S(n14044), .Z(
        P1_U3583) );
  MUX2_X1 U15958 ( .A(n14027), .B(P1_DATAO_REG_22__SCAN_IN), .S(n14044), .Z(
        P1_U3582) );
  MUX2_X1 U15959 ( .A(n14248), .B(P1_DATAO_REG_21__SCAN_IN), .S(n14044), .Z(
        P1_U3581) );
  MUX2_X1 U15960 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n14028), .S(P1_U4016), .Z(
        P1_U3580) );
  MUX2_X1 U15961 ( .A(n14322), .B(P1_DATAO_REG_19__SCAN_IN), .S(n14044), .Z(
        P1_U3579) );
  MUX2_X1 U15962 ( .A(n14029), .B(P1_DATAO_REG_18__SCAN_IN), .S(n14044), .Z(
        P1_U3578) );
  MUX2_X1 U15963 ( .A(n14320), .B(P1_DATAO_REG_17__SCAN_IN), .S(n14044), .Z(
        P1_U3577) );
  MUX2_X1 U15964 ( .A(n14030), .B(P1_DATAO_REG_15__SCAN_IN), .S(n14044), .Z(
        P1_U3575) );
  MUX2_X1 U15965 ( .A(n14031), .B(P1_DATAO_REG_14__SCAN_IN), .S(n14044), .Z(
        P1_U3574) );
  MUX2_X1 U15966 ( .A(n14032), .B(P1_DATAO_REG_13__SCAN_IN), .S(n14044), .Z(
        P1_U3573) );
  MUX2_X1 U15967 ( .A(n14033), .B(P1_DATAO_REG_12__SCAN_IN), .S(n14044), .Z(
        P1_U3572) );
  MUX2_X1 U15968 ( .A(n14034), .B(P1_DATAO_REG_11__SCAN_IN), .S(n14044), .Z(
        P1_U3571) );
  MUX2_X1 U15969 ( .A(n14035), .B(P1_DATAO_REG_10__SCAN_IN), .S(n14044), .Z(
        P1_U3570) );
  MUX2_X1 U15970 ( .A(n14036), .B(P1_DATAO_REG_9__SCAN_IN), .S(n14044), .Z(
        P1_U3569) );
  MUX2_X1 U15971 ( .A(n14037), .B(P1_DATAO_REG_8__SCAN_IN), .S(n14044), .Z(
        P1_U3568) );
  MUX2_X1 U15972 ( .A(n14038), .B(P1_DATAO_REG_7__SCAN_IN), .S(n14044), .Z(
        P1_U3567) );
  MUX2_X1 U15973 ( .A(n14039), .B(P1_DATAO_REG_6__SCAN_IN), .S(n14044), .Z(
        P1_U3566) );
  MUX2_X1 U15974 ( .A(n14040), .B(P1_DATAO_REG_5__SCAN_IN), .S(n14044), .Z(
        P1_U3565) );
  MUX2_X1 U15975 ( .A(n14041), .B(P1_DATAO_REG_4__SCAN_IN), .S(n14044), .Z(
        P1_U3564) );
  MUX2_X1 U15976 ( .A(n14042), .B(P1_DATAO_REG_3__SCAN_IN), .S(n14044), .Z(
        P1_U3563) );
  MUX2_X1 U15977 ( .A(n14043), .B(P1_DATAO_REG_2__SCAN_IN), .S(n14044), .Z(
        P1_U3562) );
  MUX2_X1 U15978 ( .A(n14045), .B(P1_DATAO_REG_1__SCAN_IN), .S(n14044), .Z(
        P1_U3561) );
  MUX2_X1 U15979 ( .A(n14046), .B(P1_DATAO_REG_0__SCAN_IN), .S(n14044), .Z(
        P1_U3560) );
  INV_X1 U15980 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n14047) );
  OAI22_X1 U15981 ( .A1(n14815), .A2(n14487), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14047), .ZN(n14048) );
  AOI21_X1 U15982 ( .B1(n14108), .B2(n14052), .A(n14048), .ZN(n14058) );
  NAND2_X1 U15983 ( .A1(n14050), .A2(n14049), .ZN(n14051) );
  NAND3_X1 U15984 ( .A1(n14102), .A2(n14071), .A3(n14051), .ZN(n14057) );
  NAND2_X1 U15985 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n14061) );
  INV_X1 U15986 ( .A(n14061), .ZN(n14055) );
  MUX2_X1 U15987 ( .A(P1_REG2_REG_1__SCAN_IN), .B(n14341), .S(n14052), .Z(
        n14054) );
  INV_X1 U15988 ( .A(n14078), .ZN(n14053) );
  OAI211_X1 U15989 ( .C1(n14055), .C2(n14054), .A(n14113), .B(n14053), .ZN(
        n14056) );
  NAND3_X1 U15990 ( .A1(n14058), .A2(n14057), .A3(n14056), .ZN(P1_U3244) );
  MUX2_X1 U15991 ( .A(n14061), .B(n14060), .S(n14059), .Z(n14062) );
  NOR2_X1 U15992 ( .A1(n14062), .A2(n8291), .ZN(n14063) );
  AOI211_X1 U15993 ( .C1(n14065), .C2(n14064), .A(n14044), .B(n14063), .ZN(
        n14798) );
  INV_X1 U15994 ( .A(n14798), .ZN(n14082) );
  OAI22_X1 U15995 ( .A1(n14815), .A2(n14532), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14066), .ZN(n14067) );
  AOI21_X1 U15996 ( .B1(n14108), .B2(n14073), .A(n14067), .ZN(n14081) );
  INV_X1 U15997 ( .A(n14068), .ZN(n14093) );
  NAND3_X1 U15998 ( .A1(n14071), .A2(n14070), .A3(n14069), .ZN(n14072) );
  NAND3_X1 U15999 ( .A1(n14102), .A2(n14093), .A3(n14072), .ZN(n14080) );
  MUX2_X1 U16000 ( .A(n9797), .B(P1_REG2_REG_2__SCAN_IN), .S(n14073), .Z(
        n14076) );
  INV_X1 U16001 ( .A(n14074), .ZN(n14075) );
  NAND2_X1 U16002 ( .A1(n14076), .A2(n14075), .ZN(n14077) );
  OAI211_X1 U16003 ( .C1(n14078), .C2(n14077), .A(n14113), .B(n14085), .ZN(
        n14079) );
  NAND4_X1 U16004 ( .A1(n14082), .A2(n14081), .A3(n14080), .A4(n14079), .ZN(
        P1_U3245) );
  INV_X1 U16005 ( .A(n14791), .ZN(n14087) );
  NAND3_X1 U16006 ( .A1(n14085), .A2(n14084), .A3(n14083), .ZN(n14086) );
  NAND3_X1 U16007 ( .A1(n14113), .A2(n14087), .A3(n14086), .ZN(n14098) );
  NAND2_X1 U16008 ( .A1(n14108), .A2(n6752), .ZN(n14097) );
  AOI22_X1 U16009 ( .A1(n14088), .A2(P1_ADDR_REG_3__SCAN_IN), .B1(
        P1_REG3_REG_3__SCAN_IN), .B2(P1_U3086), .ZN(n14096) );
  INV_X1 U16010 ( .A(n14089), .ZN(n14092) );
  MUX2_X1 U16011 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n9789), .S(n14090), .Z(
        n14091) );
  NAND3_X1 U16012 ( .A1(n14093), .A2(n14092), .A3(n14091), .ZN(n14094) );
  NAND3_X1 U16013 ( .A1(n14102), .A2(n14785), .A3(n14094), .ZN(n14095) );
  NAND4_X1 U16014 ( .A1(n14098), .A2(n14097), .A3(n14096), .A4(n14095), .ZN(
        P1_U3246) );
  OAI21_X1 U16015 ( .B1(n14101), .B2(n14100), .A(n14099), .ZN(n14103) );
  NAND2_X1 U16016 ( .A1(n14103), .A2(n14102), .ZN(n14117) );
  INV_X1 U16017 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n14105) );
  OAI21_X1 U16018 ( .B1(n14815), .B2(n14105), .A(n14104), .ZN(n14106) );
  AOI21_X1 U16019 ( .B1(n14108), .B2(n14107), .A(n14106), .ZN(n14116) );
  OR3_X1 U16020 ( .A1(n14111), .A2(n14110), .A3(n14109), .ZN(n14112) );
  NAND3_X1 U16021 ( .A1(n14114), .A2(n14113), .A3(n14112), .ZN(n14115) );
  NAND3_X1 U16022 ( .A1(n14117), .A2(n14116), .A3(n14115), .ZN(P1_U3254) );
  XNOR2_X1 U16023 ( .A(n14119), .B(n14118), .ZN(n14352) );
  NAND2_X1 U16024 ( .A1(n14352), .A2(n14344), .ZN(n14122) );
  NOR2_X1 U16025 ( .A1(n14830), .A2(n14120), .ZN(n14123) );
  AOI21_X1 U16026 ( .B1(n14830), .B2(P1_REG2_REG_31__SCAN_IN), .A(n14123), 
        .ZN(n14121) );
  OAI211_X1 U16027 ( .C1(n14437), .C2(n14823), .A(n14122), .B(n14121), .ZN(
        P1_U3263) );
  INV_X1 U16028 ( .A(n14123), .ZN(n14124) );
  OAI21_X1 U16029 ( .B1(n14313), .B2(n14125), .A(n14124), .ZN(n14126) );
  AOI21_X1 U16030 ( .B1(n14438), .B2(n14346), .A(n14126), .ZN(n14127) );
  OAI21_X1 U16031 ( .B1(n14128), .B2(n14243), .A(n14127), .ZN(P1_U3264) );
  OAI21_X1 U16032 ( .B1(n14135), .B2(n14130), .A(n14129), .ZN(n14132) );
  AOI21_X1 U16033 ( .B1(n14135), .B2(n14134), .A(n14133), .ZN(n14358) );
  OAI211_X1 U16034 ( .C1(n14156), .C2(n14356), .A(n14427), .B(n14136), .ZN(
        n14355) );
  AOI22_X1 U16035 ( .A1(n14830), .A2(P1_REG2_REG_28__SCAN_IN), .B1(n14137), 
        .B2(n14819), .ZN(n14140) );
  NAND2_X1 U16036 ( .A1(n14138), .A2(n14346), .ZN(n14139) );
  OAI211_X1 U16037 ( .C1(n14355), .C2(n14243), .A(n14140), .B(n14139), .ZN(
        n14141) );
  AOI21_X1 U16038 ( .B1(n14358), .B2(n14277), .A(n14141), .ZN(n14142) );
  OAI21_X1 U16039 ( .B1(n14359), .B2(n14830), .A(n14142), .ZN(P1_U3265) );
  OAI21_X1 U16040 ( .B1(n14145), .B2(n14144), .A(n14143), .ZN(n14363) );
  INV_X1 U16041 ( .A(n14363), .ZN(n14166) );
  AOI22_X1 U16042 ( .A1(n14319), .A2(n14147), .B1(n14146), .B2(n14321), .ZN(
        n14154) );
  INV_X1 U16043 ( .A(n14148), .ZN(n14152) );
  NOR3_X1 U16044 ( .A1(n14168), .A2(n14150), .A3(n14149), .ZN(n14151) );
  OAI21_X1 U16045 ( .B1(n14152), .B2(n14151), .A(n14324), .ZN(n14153) );
  NAND2_X1 U16046 ( .A1(n14361), .A2(n14313), .ZN(n14164) );
  INV_X1 U16047 ( .A(n14181), .ZN(n14157) );
  AOI211_X1 U16048 ( .C1(n14158), .C2(n14157), .A(n14326), .B(n14156), .ZN(
        n14362) );
  NOR2_X1 U16049 ( .A1(n9496), .A2(n14823), .ZN(n14162) );
  OAI22_X1 U16050 ( .A1(n14313), .A2(n14160), .B1(n14159), .B2(n14307), .ZN(
        n14161) );
  AOI211_X1 U16051 ( .C1(n14362), .C2(n14817), .A(n14162), .B(n14161), .ZN(
        n14163) );
  OAI211_X1 U16052 ( .C1(n14166), .C2(n14165), .A(n14164), .B(n14163), .ZN(
        P1_U3266) );
  XNOR2_X1 U16053 ( .A(n14167), .B(n14171), .ZN(n14369) );
  INV_X1 U16054 ( .A(n14168), .ZN(n14173) );
  NAND3_X1 U16055 ( .A1(n14169), .A2(n14171), .A3(n14170), .ZN(n14172) );
  NAND2_X1 U16056 ( .A1(n14173), .A2(n14172), .ZN(n14176) );
  AOI222_X1 U16057 ( .A1(n14324), .A2(n14176), .B1(n14175), .B2(n14321), .C1(
        n14174), .C2(n14319), .ZN(n14368) );
  NAND2_X1 U16058 ( .A1(n14830), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n14177) );
  OAI21_X1 U16059 ( .B1(n14307), .B2(n14178), .A(n14177), .ZN(n14179) );
  AOI21_X1 U16060 ( .B1(n14366), .B2(n14346), .A(n14179), .ZN(n14184) );
  OAI21_X1 U16061 ( .B1(n14194), .B2(n14180), .A(n14427), .ZN(n14182) );
  NOR2_X1 U16062 ( .A1(n14182), .A2(n14181), .ZN(n14365) );
  NAND2_X1 U16063 ( .A1(n14365), .A2(n14817), .ZN(n14183) );
  OAI211_X1 U16064 ( .C1(n14368), .C2(n14830), .A(n14184), .B(n14183), .ZN(
        n14185) );
  INV_X1 U16065 ( .A(n14185), .ZN(n14186) );
  OAI21_X1 U16066 ( .B1(n14369), .B2(n14334), .A(n14186), .ZN(P1_U3267) );
  NAND2_X1 U16067 ( .A1(n14187), .A2(n14192), .ZN(n14188) );
  NAND2_X1 U16068 ( .A1(n14169), .A2(n14188), .ZN(n14190) );
  AOI21_X1 U16069 ( .B1(n14190), .B2(n14324), .A(n14189), .ZN(n14371) );
  OAI21_X1 U16070 ( .B1(n14193), .B2(n14192), .A(n14191), .ZN(n14372) );
  INV_X1 U16071 ( .A(n14372), .ZN(n14202) );
  INV_X1 U16072 ( .A(n14194), .ZN(n14196) );
  AOI21_X1 U16073 ( .B1(n14220), .B2(n14374), .A(n14326), .ZN(n14195) );
  NAND2_X1 U16074 ( .A1(n14196), .A2(n14195), .ZN(n14370) );
  NAND2_X1 U16075 ( .A1(n14830), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n14197) );
  OAI21_X1 U16076 ( .B1(n14307), .B2(n14198), .A(n14197), .ZN(n14199) );
  AOI21_X1 U16077 ( .B1(n14374), .B2(n14346), .A(n14199), .ZN(n14200) );
  OAI21_X1 U16078 ( .B1(n14370), .B2(n14243), .A(n14200), .ZN(n14201) );
  AOI21_X1 U16079 ( .B1(n14202), .B2(n14277), .A(n14201), .ZN(n14203) );
  OAI21_X1 U16080 ( .B1(n14830), .B2(n14371), .A(n14203), .ZN(P1_U3268) );
  NAND2_X1 U16081 ( .A1(n14236), .A2(n14204), .ZN(n14206) );
  NAND2_X1 U16082 ( .A1(n14206), .A2(n14205), .ZN(n14207) );
  NAND2_X1 U16083 ( .A1(n14208), .A2(n14207), .ZN(n14382) );
  NAND2_X1 U16084 ( .A1(n14382), .A2(n14209), .ZN(n14218) );
  AOI21_X1 U16085 ( .B1(n14211), .B2(n14210), .A(n14282), .ZN(n14216) );
  NAND2_X1 U16086 ( .A1(n14249), .A2(n14319), .ZN(n14212) );
  OAI21_X1 U16087 ( .B1(n14213), .B2(n14287), .A(n14212), .ZN(n14214) );
  AOI21_X1 U16088 ( .B1(n14216), .B2(n14215), .A(n14214), .ZN(n14217) );
  INV_X1 U16089 ( .A(n14219), .ZN(n14237) );
  AOI21_X1 U16090 ( .B1(n14237), .B2(n14377), .A(n14326), .ZN(n14221) );
  NAND2_X1 U16091 ( .A1(n14221), .A2(n14220), .ZN(n14378) );
  OAI22_X1 U16092 ( .A1(n14313), .A2(n14223), .B1(n14222), .B2(n14307), .ZN(
        n14224) );
  AOI21_X1 U16093 ( .B1(n14377), .B2(n14346), .A(n14224), .ZN(n14225) );
  OAI21_X1 U16094 ( .B1(n14378), .B2(n14243), .A(n14225), .ZN(n14226) );
  AOI21_X1 U16095 ( .B1(n14382), .B2(n14826), .A(n14226), .ZN(n14227) );
  OAI21_X1 U16096 ( .B1(n14384), .B2(n14830), .A(n14227), .ZN(P1_U3269) );
  OR2_X1 U16097 ( .A1(n14228), .A2(n14233), .ZN(n14229) );
  NAND2_X1 U16098 ( .A1(n14230), .A2(n14229), .ZN(n14232) );
  AOI21_X1 U16099 ( .B1(n14232), .B2(n14324), .A(n14231), .ZN(n14389) );
  NAND2_X1 U16100 ( .A1(n14234), .A2(n14233), .ZN(n14235) );
  AND2_X1 U16101 ( .A1(n14236), .A2(n14235), .ZN(n14386) );
  AOI21_X1 U16102 ( .B1(n14385), .B2(n14254), .A(n14326), .ZN(n14238) );
  NAND2_X1 U16103 ( .A1(n14238), .A2(n14237), .ZN(n14387) );
  INV_X1 U16104 ( .A(n14239), .ZN(n14240) );
  AOI22_X1 U16105 ( .A1(n14240), .A2(n14819), .B1(P1_REG2_REG_23__SCAN_IN), 
        .B2(n14830), .ZN(n14242) );
  NAND2_X1 U16106 ( .A1(n14385), .A2(n14346), .ZN(n14241) );
  OAI211_X1 U16107 ( .C1(n14387), .C2(n14243), .A(n14242), .B(n14241), .ZN(
        n14244) );
  AOI21_X1 U16108 ( .B1(n14386), .B2(n14277), .A(n14244), .ZN(n14245) );
  OAI21_X1 U16109 ( .B1(n14389), .B2(n14830), .A(n14245), .ZN(P1_U3270) );
  XNOR2_X1 U16110 ( .A(n14247), .B(n14246), .ZN(n14250) );
  AOI222_X1 U16111 ( .A1(n14324), .A2(n14250), .B1(n14249), .B2(n14321), .C1(
        n14248), .C2(n14319), .ZN(n14396) );
  OAI21_X1 U16112 ( .B1(n14253), .B2(n14252), .A(n14251), .ZN(n14392) );
  INV_X1 U16113 ( .A(n14254), .ZN(n14255) );
  AOI211_X1 U16114 ( .C1(n14394), .C2(n14268), .A(n14326), .B(n14255), .ZN(
        n14393) );
  NAND2_X1 U16115 ( .A1(n14393), .A2(n14817), .ZN(n14258) );
  AOI22_X1 U16116 ( .A1(n14256), .A2(n14819), .B1(n14830), .B2(
        P1_REG2_REG_22__SCAN_IN), .ZN(n14257) );
  OAI211_X1 U16117 ( .C1(n14823), .C2(n14259), .A(n14258), .B(n14257), .ZN(
        n14260) );
  AOI21_X1 U16118 ( .B1(n14277), .B2(n14392), .A(n14260), .ZN(n14261) );
  OAI21_X1 U16119 ( .B1(n14830), .B2(n14396), .A(n14261), .ZN(P1_U3271) );
  XNOR2_X1 U16120 ( .A(n14262), .B(n14266), .ZN(n14263) );
  OAI222_X1 U16121 ( .A1(n14287), .A2(n14265), .B1(n14285), .B2(n14264), .C1(
        n14263), .C2(n14282), .ZN(n14398) );
  INV_X1 U16122 ( .A(n14398), .ZN(n14279) );
  XNOR2_X1 U16123 ( .A(n14267), .B(n14266), .ZN(n14400) );
  INV_X1 U16124 ( .A(n14294), .ZN(n14270) );
  INV_X1 U16125 ( .A(n14268), .ZN(n14269) );
  AOI211_X1 U16126 ( .C1(n14271), .C2(n14270), .A(n14326), .B(n14269), .ZN(
        n14399) );
  NAND2_X1 U16127 ( .A1(n14399), .A2(n14817), .ZN(n14275) );
  INV_X1 U16128 ( .A(n14272), .ZN(n14273) );
  AOI22_X1 U16129 ( .A1(n14830), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n14273), 
        .B2(n14819), .ZN(n14274) );
  OAI211_X1 U16130 ( .C1(n14461), .C2(n14823), .A(n14275), .B(n14274), .ZN(
        n14276) );
  AOI21_X1 U16131 ( .B1(n14277), .B2(n14400), .A(n14276), .ZN(n14278) );
  OAI21_X1 U16132 ( .B1(n14830), .B2(n14279), .A(n14278), .ZN(P1_U3272) );
  XNOR2_X1 U16133 ( .A(n14281), .B(n14280), .ZN(n14407) );
  AOI21_X1 U16134 ( .B1(n14284), .B2(n14283), .A(n14282), .ZN(n14291) );
  OAI22_X1 U16135 ( .A1(n14288), .A2(n14287), .B1(n14286), .B2(n14285), .ZN(
        n14289) );
  AOI21_X1 U16136 ( .B1(n14291), .B2(n14290), .A(n14289), .ZN(n14405) );
  OAI21_X1 U16137 ( .B1(n14292), .B2(n14307), .A(n14405), .ZN(n14293) );
  NAND2_X1 U16138 ( .A1(n14293), .A2(n14313), .ZN(n14299) );
  AOI211_X1 U16139 ( .C1(n14404), .C2(n14311), .A(n14326), .B(n14294), .ZN(
        n14403) );
  INV_X1 U16140 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n14295) );
  OAI22_X1 U16141 ( .A1(n14296), .A2(n14823), .B1(n14295), .B2(n14313), .ZN(
        n14297) );
  AOI21_X1 U16142 ( .B1(n14403), .B2(n14817), .A(n14297), .ZN(n14298) );
  OAI211_X1 U16143 ( .C1(n14407), .C2(n14334), .A(n14299), .B(n14298), .ZN(
        P1_U3273) );
  INV_X1 U16144 ( .A(n14300), .ZN(n14301) );
  AOI21_X1 U16145 ( .B1(n14303), .B2(n14302), .A(n14301), .ZN(n14412) );
  XNOR2_X1 U16146 ( .A(n6686), .B(n7045), .ZN(n14306) );
  AOI21_X1 U16147 ( .B1(n14306), .B2(n14324), .A(n14305), .ZN(n14410) );
  OAI21_X1 U16148 ( .B1(n14308), .B2(n14307), .A(n14410), .ZN(n14309) );
  NAND2_X1 U16149 ( .A1(n14309), .A2(n14313), .ZN(n14317) );
  INV_X1 U16150 ( .A(n14311), .ZN(n14312) );
  AOI211_X1 U16151 ( .C1(n14409), .C2(n14325), .A(n14326), .B(n14312), .ZN(
        n14408) );
  INV_X1 U16152 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n14314) );
  OAI22_X1 U16153 ( .A1(n9549), .A2(n14823), .B1(n14314), .B2(n14313), .ZN(
        n14315) );
  AOI21_X1 U16154 ( .B1(n14408), .B2(n14817), .A(n14315), .ZN(n14316) );
  OAI211_X1 U16155 ( .C1(n14412), .C2(n14334), .A(n14317), .B(n14316), .ZN(
        P1_U3274) );
  XOR2_X1 U16156 ( .A(n14318), .B(n14332), .Z(n14323) );
  AOI222_X1 U16157 ( .A1(n14324), .A2(n14323), .B1(n14322), .B2(n14321), .C1(
        n14320), .C2(n14319), .ZN(n14416) );
  AOI211_X1 U16158 ( .C1(n14414), .C2(n14327), .A(n14326), .B(n14310), .ZN(
        n14413) );
  INV_X1 U16159 ( .A(n14414), .ZN(n14331) );
  INV_X1 U16160 ( .A(n14328), .ZN(n14329) );
  AOI22_X1 U16161 ( .A1(n14830), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n14329), 
        .B2(n14819), .ZN(n14330) );
  OAI21_X1 U16162 ( .B1(n14331), .B2(n14823), .A(n14330), .ZN(n14336) );
  XOR2_X1 U16163 ( .A(n14333), .B(n14332), .Z(n14417) );
  NOR2_X1 U16164 ( .A1(n14417), .A2(n14334), .ZN(n14335) );
  AOI211_X1 U16165 ( .C1(n14413), .C2(n14817), .A(n14336), .B(n14335), .ZN(
        n14337) );
  OAI21_X1 U16166 ( .B1(n14830), .B2(n14416), .A(n14337), .ZN(P1_U3275) );
  NOR2_X1 U16167 ( .A1(n14339), .A2(n14338), .ZN(n14340) );
  MUX2_X1 U16168 ( .A(n14341), .B(n14340), .S(n14313), .Z(n14350) );
  INV_X1 U16169 ( .A(n14342), .ZN(n14343) );
  AOI22_X1 U16170 ( .A1(n14344), .A2(n14343), .B1(P1_REG3_REG_1__SCAN_IN), 
        .B2(n14819), .ZN(n14349) );
  AOI22_X1 U16171 ( .A1(n14826), .A2(n14347), .B1(n14346), .B2(n14345), .ZN(
        n14348) );
  NAND3_X1 U16172 ( .A1(n14350), .A2(n14349), .A3(n14348), .ZN(P1_U3292) );
  INV_X1 U16173 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n14353) );
  AOI21_X1 U16174 ( .B1(n14352), .B2(n14427), .A(n14351), .ZN(n14434) );
  MUX2_X1 U16175 ( .A(n14353), .B(n14434), .S(n14856), .Z(n14354) );
  OAI21_X1 U16176 ( .B1(n14437), .B2(n14423), .A(n14354), .ZN(P1_U3559) );
  OAI21_X1 U16177 ( .B1(n14356), .B2(n14843), .A(n14355), .ZN(n14357) );
  AOI21_X1 U16178 ( .B1(n14358), .B2(n14848), .A(n14357), .ZN(n14360) );
  MUX2_X1 U16179 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n14444), .S(n14856), .Z(
        P1_U3556) );
  INV_X1 U16180 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n14364) );
  AOI21_X1 U16181 ( .B1(n14426), .B2(n14366), .A(n14365), .ZN(n14367) );
  OAI211_X1 U16182 ( .C1(n14431), .C2(n14369), .A(n14368), .B(n14367), .ZN(
        n14447) );
  MUX2_X1 U16183 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n14447), .S(n14856), .Z(
        P1_U3554) );
  OAI211_X1 U16184 ( .C1(n14372), .C2(n14431), .A(n14371), .B(n14370), .ZN(
        n14448) );
  MUX2_X1 U16185 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n14448), .S(n14856), .Z(
        n14373) );
  AOI21_X1 U16186 ( .B1(n14375), .B2(n14374), .A(n14373), .ZN(n14376) );
  INV_X1 U16187 ( .A(n14376), .ZN(P1_U3553) );
  INV_X1 U16188 ( .A(n14377), .ZN(n14379) );
  OAI21_X1 U16189 ( .B1(n14379), .B2(n14843), .A(n14378), .ZN(n14380) );
  AOI21_X1 U16190 ( .B1(n14382), .B2(n14381), .A(n14380), .ZN(n14383) );
  NAND2_X1 U16191 ( .A1(n14384), .A2(n14383), .ZN(n14452) );
  MUX2_X1 U16192 ( .A(n14452), .B(P1_REG1_REG_24__SCAN_IN), .S(n14854), .Z(
        P1_U3552) );
  INV_X1 U16193 ( .A(n14385), .ZN(n14456) );
  NAND2_X1 U16194 ( .A1(n14386), .A2(n14848), .ZN(n14388) );
  AND3_X1 U16195 ( .A1(n14389), .A2(n14388), .A3(n14387), .ZN(n14453) );
  MUX2_X1 U16196 ( .A(n14390), .B(n14453), .S(n14856), .Z(n14391) );
  OAI21_X1 U16197 ( .B1(n14456), .B2(n14423), .A(n14391), .ZN(P1_U3551) );
  INV_X1 U16198 ( .A(n14392), .ZN(n14397) );
  AOI21_X1 U16199 ( .B1(n14426), .B2(n14394), .A(n14393), .ZN(n14395) );
  OAI211_X1 U16200 ( .C1(n14431), .C2(n14397), .A(n14396), .B(n14395), .ZN(
        n14457) );
  MUX2_X1 U16201 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n14457), .S(n14856), .Z(
        P1_U3550) );
  AOI211_X1 U16202 ( .C1(n14848), .C2(n14400), .A(n14399), .B(n14398), .ZN(
        n14458) );
  MUX2_X1 U16203 ( .A(n14401), .B(n14458), .S(n14856), .Z(n14402) );
  OAI21_X1 U16204 ( .B1(n14461), .B2(n14423), .A(n14402), .ZN(P1_U3549) );
  AOI21_X1 U16205 ( .B1(n14426), .B2(n14404), .A(n14403), .ZN(n14406) );
  OAI211_X1 U16206 ( .C1(n14431), .C2(n14407), .A(n14406), .B(n14405), .ZN(
        n14462) );
  MUX2_X1 U16207 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n14462), .S(n14856), .Z(
        P1_U3548) );
  AOI21_X1 U16208 ( .B1(n14426), .B2(n14409), .A(n14408), .ZN(n14411) );
  OAI211_X1 U16209 ( .C1(n14412), .C2(n14431), .A(n14411), .B(n14410), .ZN(
        n14463) );
  MUX2_X1 U16210 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n14463), .S(n14856), .Z(
        P1_U3547) );
  AOI21_X1 U16211 ( .B1(n14426), .B2(n14414), .A(n14413), .ZN(n14415) );
  OAI211_X1 U16212 ( .C1(n14431), .C2(n14417), .A(n14416), .B(n14415), .ZN(
        n14464) );
  MUX2_X1 U16213 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n14464), .S(n14856), .Z(
        P1_U3546) );
  AOI211_X1 U16214 ( .C1(n14848), .C2(n14420), .A(n14419), .B(n14418), .ZN(
        n14465) );
  MUX2_X1 U16215 ( .A(n14421), .B(n14465), .S(n14856), .Z(n14422) );
  OAI21_X1 U16216 ( .B1(n14469), .B2(n14423), .A(n14422), .ZN(P1_U3545) );
  INV_X1 U16217 ( .A(n14424), .ZN(n14432) );
  AOI22_X1 U16218 ( .A1(n14428), .A2(n14427), .B1(n14426), .B2(n14425), .ZN(
        n14429) );
  OAI211_X1 U16219 ( .C1(n14432), .C2(n14431), .A(n14430), .B(n14429), .ZN(
        n14470) );
  MUX2_X1 U16220 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n14470), .S(n14856), .Z(
        P1_U3544) );
  MUX2_X1 U16221 ( .A(P1_REG1_REG_0__SCAN_IN), .B(n14433), .S(n14856), .Z(
        P1_U3528) );
  MUX2_X1 U16222 ( .A(n14435), .B(n14434), .S(n14849), .Z(n14436) );
  OAI21_X1 U16223 ( .B1(n14437), .B2(n14468), .A(n14436), .ZN(P1_U3527) );
  INV_X1 U16224 ( .A(n14438), .ZN(n14443) );
  INV_X1 U16225 ( .A(n14439), .ZN(n14440) );
  MUX2_X1 U16226 ( .A(n14441), .B(n14440), .S(n14849), .Z(n14442) );
  OAI21_X1 U16227 ( .B1(n14443), .B2(n14468), .A(n14442), .ZN(P1_U3526) );
  MUX2_X1 U16228 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n14444), .S(n14849), .Z(
        P1_U3524) );
  MUX2_X1 U16229 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n14447), .S(n14849), .Z(
        P1_U3522) );
  MUX2_X1 U16230 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n14448), .S(n14849), .Z(
        n14449) );
  INV_X1 U16231 ( .A(n14449), .ZN(n14450) );
  OAI21_X1 U16232 ( .B1(n14451), .B2(n14468), .A(n14450), .ZN(P1_U3521) );
  MUX2_X1 U16233 ( .A(n14452), .B(P1_REG0_REG_24__SCAN_IN), .S(n6786), .Z(
        P1_U3520) );
  INV_X1 U16234 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n14454) );
  MUX2_X1 U16235 ( .A(n14454), .B(n14453), .S(n14849), .Z(n14455) );
  OAI21_X1 U16236 ( .B1(n14456), .B2(n14468), .A(n14455), .ZN(P1_U3519) );
  MUX2_X1 U16237 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n14457), .S(n14849), .Z(
        P1_U3518) );
  INV_X1 U16238 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n14459) );
  MUX2_X1 U16239 ( .A(n14459), .B(n14458), .S(n14849), .Z(n14460) );
  OAI21_X1 U16240 ( .B1(n14461), .B2(n14468), .A(n14460), .ZN(P1_U3517) );
  MUX2_X1 U16241 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n14462), .S(n14849), .Z(
        P1_U3516) );
  MUX2_X1 U16242 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n14463), .S(n14849), .Z(
        P1_U3515) );
  MUX2_X1 U16243 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n14464), .S(n14849), .Z(
        P1_U3513) );
  INV_X1 U16244 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n14466) );
  MUX2_X1 U16245 ( .A(n14466), .B(n14465), .S(n14849), .Z(n14467) );
  OAI21_X1 U16246 ( .B1(n14469), .B2(n14468), .A(n14467), .ZN(P1_U3510) );
  MUX2_X1 U16247 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n14470), .S(n14849), .Z(
        P1_U3507) );
  NOR4_X1 U16248 ( .A1(n14471), .A2(P1_IR_REG_30__SCAN_IN), .A3(n7672), .A4(
        P1_U3086), .ZN(n14472) );
  AOI21_X1 U16249 ( .B1(n14473), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n14472), 
        .ZN(n14474) );
  OAI21_X1 U16250 ( .B1(n14475), .B2(n14480), .A(n14474), .ZN(P1_U3324) );
  OAI222_X1 U16251 ( .A1(n14480), .A2(n14479), .B1(n14478), .B2(n14477), .C1(
        n14476), .C2(P1_U3086), .ZN(P1_U3326) );
  MUX2_X1 U16252 ( .A(n14483), .B(n14482), .S(P1_U3086), .Z(P1_U3333) );
  MUX2_X1 U16253 ( .A(n14484), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  INV_X1 U16254 ( .A(P3_ADDR_REG_16__SCAN_IN), .ZN(n14649) );
  XOR2_X1 U16255 ( .A(P1_ADDR_REG_16__SCAN_IN), .B(n14649), .Z(n14515) );
  INV_X1 U16256 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n14816) );
  INV_X1 U16257 ( .A(P3_ADDR_REG_14__SCAN_IN), .ZN(n14516) );
  NOR2_X1 U16258 ( .A1(P1_ADDR_REG_14__SCAN_IN), .A2(n14516), .ZN(n14513) );
  INV_X1 U16259 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n14571) );
  AND2_X1 U16260 ( .A1(n14571), .A2(P1_ADDR_REG_13__SCAN_IN), .ZN(n14511) );
  INV_X1 U16261 ( .A(P3_ADDR_REG_12__SCAN_IN), .ZN(n14520) );
  NOR2_X1 U16262 ( .A1(P1_ADDR_REG_12__SCAN_IN), .A2(n14520), .ZN(n14519) );
  INV_X1 U16263 ( .A(P3_ADDR_REG_11__SCAN_IN), .ZN(n14509) );
  INV_X1 U16264 ( .A(P3_ADDR_REG_10__SCAN_IN), .ZN(n14507) );
  NAND2_X1 U16265 ( .A1(P3_ADDR_REG_9__SCAN_IN), .A2(n14485), .ZN(n14505) );
  INV_X1 U16266 ( .A(P3_ADDR_REG_9__SCAN_IN), .ZN(n14486) );
  AOI22_X1 U16267 ( .A1(P1_ADDR_REG_9__SCAN_IN), .A2(n14486), .B1(
        P3_ADDR_REG_9__SCAN_IN), .B2(n14485), .ZN(n14563) );
  NOR2_X1 U16268 ( .A1(n14490), .A2(n15125), .ZN(n14492) );
  NOR2_X1 U16269 ( .A1(n14493), .A2(n15145), .ZN(n14495) );
  NOR2_X1 U16270 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n14548), .ZN(n14494) );
  INV_X1 U16271 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n14552) );
  NOR2_X1 U16272 ( .A1(P3_ADDR_REG_6__SCAN_IN), .A2(n14552), .ZN(n14497) );
  NOR2_X1 U16273 ( .A1(P3_ADDR_REG_7__SCAN_IN), .A2(n14498), .ZN(n14500) );
  XOR2_X1 U16274 ( .A(n15169), .B(n14498), .Z(n14556) );
  NOR2_X1 U16275 ( .A1(n14556), .A2(n14557), .ZN(n14499) );
  NAND2_X1 U16276 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n14503), .ZN(n14501) );
  OAI21_X1 U16277 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(n14503), .A(n14501), .ZN(
        n14527) );
  NOR2_X1 U16278 ( .A1(n14528), .A2(n14527), .ZN(n14502) );
  NAND2_X1 U16279 ( .A1(n14505), .A2(n14504), .ZN(n14526) );
  XNOR2_X1 U16280 ( .A(n14507), .B(P1_ADDR_REG_10__SCAN_IN), .ZN(n14525) );
  NOR2_X1 U16281 ( .A1(n14526), .A2(n14525), .ZN(n14506) );
  XNOR2_X1 U16282 ( .A(n14509), .B(P1_ADDR_REG_11__SCAN_IN), .ZN(n14523) );
  OAI22_X1 U16283 ( .A1(n14513), .A2(n14518), .B1(P3_ADDR_REG_14__SCAN_IN), 
        .B2(n14512), .ZN(n14578) );
  INV_X1 U16284 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n14624) );
  XNOR2_X1 U16285 ( .A(P1_ADDR_REG_15__SCAN_IN), .B(n14624), .ZN(n14577) );
  NOR2_X1 U16286 ( .A1(n14578), .A2(n14577), .ZN(n14514) );
  XOR2_X1 U16287 ( .A(n14515), .B(n14584), .Z(n14582) );
  INV_X1 U16288 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n14580) );
  XNOR2_X1 U16289 ( .A(n14516), .B(P1_ADDR_REG_14__SCAN_IN), .ZN(n14517) );
  XOR2_X1 U16290 ( .A(n14518), .B(n14517), .Z(n14574) );
  INV_X1 U16291 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n14898) );
  AOI21_X1 U16292 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(n14520), .A(n14519), 
        .ZN(n14522) );
  XNOR2_X1 U16293 ( .A(n14522), .B(n14521), .ZN(n14769) );
  XOR2_X1 U16294 ( .A(n14524), .B(n14523), .Z(n14764) );
  XOR2_X1 U16295 ( .A(n14526), .B(n14525), .Z(n14601) );
  XOR2_X1 U16296 ( .A(n14528), .B(n14527), .Z(n14562) );
  INV_X1 U16297 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n14801) );
  NAND2_X1 U16298 ( .A1(P2_ADDR_REG_4__SCAN_IN), .A2(n14530), .ZN(n14547) );
  XNOR2_X1 U16299 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(n14531), .ZN(n15290) );
  XOR2_X1 U16300 ( .A(n14532), .B(P3_ADDR_REG_2__SCAN_IN), .Z(n14534) );
  XOR2_X1 U16301 ( .A(n14534), .B(n14533), .Z(n14542) );
  NAND2_X1 U16302 ( .A1(P2_ADDR_REG_1__SCAN_IN), .A2(n14538), .ZN(n14540) );
  AOI21_X1 U16303 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(n15109), .A(n14537), .ZN(
        n15286) );
  INV_X1 U16304 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n15285) );
  NOR2_X1 U16305 ( .A1(n15286), .A2(n15285), .ZN(n15294) );
  NAND2_X1 U16306 ( .A1(n15294), .A2(n15293), .ZN(n14539) );
  NAND2_X1 U16307 ( .A1(n14542), .A2(n14541), .ZN(n14544) );
  NAND2_X1 U16308 ( .A1(n14595), .A2(P2_ADDR_REG_2__SCAN_IN), .ZN(n14543) );
  NAND2_X1 U16309 ( .A1(n14544), .A2(n14543), .ZN(n15291) );
  NOR2_X1 U16310 ( .A1(n15290), .A2(n15291), .ZN(n14545) );
  NAND2_X1 U16311 ( .A1(n15290), .A2(n15291), .ZN(n15289) );
  NAND2_X1 U16312 ( .A1(n14547), .A2(n14546), .ZN(n14550) );
  XNOR2_X1 U16313 ( .A(n14549), .B(n14550), .ZN(n15284) );
  NAND2_X1 U16314 ( .A1(n14551), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n14555) );
  XNOR2_X1 U16315 ( .A(n14552), .B(P3_ADDR_REG_6__SCAN_IN), .ZN(n14553) );
  XNOR2_X1 U16316 ( .A(n14554), .B(n14553), .ZN(n14596) );
  XOR2_X1 U16317 ( .A(n14557), .B(n14556), .Z(n15288) );
  NAND2_X1 U16318 ( .A1(n15287), .A2(n15288), .ZN(n14560) );
  NAND2_X1 U16319 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n14558), .ZN(n14559) );
  XNOR2_X1 U16320 ( .A(n14564), .B(n14563), .ZN(n14566) );
  NAND2_X1 U16321 ( .A1(n14565), .A2(n14566), .ZN(n14567) );
  NOR2_X1 U16322 ( .A1(n14601), .A2(n14602), .ZN(n14568) );
  INV_X1 U16323 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n14603) );
  NAND2_X1 U16324 ( .A1(n14601), .A2(n14602), .ZN(n14600) );
  NOR2_X1 U16325 ( .A1(n14764), .A2(n14765), .ZN(n14569) );
  NAND2_X1 U16326 ( .A1(n14764), .A2(n14765), .ZN(n14763) );
  XNOR2_X1 U16327 ( .A(P1_ADDR_REG_13__SCAN_IN), .B(n14571), .ZN(n14572) );
  XNOR2_X1 U16328 ( .A(n14573), .B(n14572), .ZN(n14773) );
  INV_X1 U16329 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n14900) );
  NOR2_X1 U16330 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(n14775), .ZN(n14576) );
  XNOR2_X1 U16331 ( .A(n14578), .B(n14577), .ZN(n14779) );
  NAND2_X1 U16332 ( .A1(n14780), .A2(n14779), .ZN(n14579) );
  OR2_X1 U16333 ( .A1(n14649), .A2(P1_ADDR_REG_16__SCAN_IN), .ZN(n14583) );
  AOI22_X1 U16334 ( .A1(P1_ADDR_REG_16__SCAN_IN), .A2(n14649), .B1(n14584), 
        .B2(n14583), .ZN(n14589) );
  XOR2_X1 U16335 ( .A(n14588), .B(n14589), .Z(n14590) );
  XNOR2_X1 U16336 ( .A(P3_ADDR_REG_17__SCAN_IN), .B(n14590), .ZN(n14585) );
  NOR2_X1 U16337 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n14614), .ZN(n14587) );
  AOI21_X1 U16338 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n14614), .A(n14587), 
        .ZN(n14612) );
  NAND2_X1 U16339 ( .A1(n14589), .A2(n14588), .ZN(n14592) );
  NAND2_X1 U16340 ( .A1(P3_ADDR_REG_17__SCAN_IN), .A2(n14590), .ZN(n14591) );
  NAND2_X1 U16341 ( .A1(n14592), .A2(n14591), .ZN(n14611) );
  XNOR2_X1 U16342 ( .A(n14612), .B(n14611), .ZN(n14607) );
  XNOR2_X1 U16343 ( .A(P2_ADDR_REG_18__SCAN_IN), .B(n14606), .ZN(SUB_1596_U62)
         );
  AOI21_X1 U16344 ( .B1(P1_WR_REG_SCAN_IN), .B2(P2_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n14593) );
  OAI21_X1 U16345 ( .B1(P1_WR_REG_SCAN_IN), .B2(P2_WR_REG_SCAN_IN), .A(n14593), 
        .ZN(U28) );
  AOI21_X1 U16346 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(
        P3_RD_REG_SCAN_IN), .ZN(n14594) );
  OAI21_X1 U16347 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(n14594), 
        .ZN(U29) );
  XOR2_X1 U16348 ( .A(n14595), .B(P2_ADDR_REG_2__SCAN_IN), .Z(SUB_1596_U61) );
  XOR2_X1 U16349 ( .A(n14597), .B(n14596), .Z(SUB_1596_U57) );
  XNOR2_X1 U16350 ( .A(n14598), .B(P2_ADDR_REG_8__SCAN_IN), .ZN(SUB_1596_U55)
         );
  XOR2_X1 U16351 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n14599), .Z(SUB_1596_U54) );
  OAI21_X1 U16352 ( .B1(n14602), .B2(n14601), .A(n14600), .ZN(n14604) );
  XOR2_X1 U16353 ( .A(n14604), .B(n14603), .Z(SUB_1596_U70) );
  XNOR2_X1 U16354 ( .A(P2_ADDR_REG_17__SCAN_IN), .B(n14605), .ZN(SUB_1596_U63)
         );
  NOR2_X1 U16355 ( .A1(n14608), .A2(n14607), .ZN(n14609) );
  NOR2_X2 U16356 ( .A1(n14610), .A2(n14609), .ZN(n14619) );
  NAND2_X1 U16357 ( .A1(n14612), .A2(n14611), .ZN(n14613) );
  OAI21_X1 U16358 ( .B1(n14614), .B2(P1_ADDR_REG_18__SCAN_IN), .A(n14613), 
        .ZN(n14617) );
  XNOR2_X1 U16359 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(P1_ADDR_REG_19__SCAN_IN), 
        .ZN(n14615) );
  XNOR2_X1 U16360 ( .A(n14615), .B(P3_ADDR_REG_19__SCAN_IN), .ZN(n14616) );
  XNOR2_X1 U16361 ( .A(n14617), .B(n14616), .ZN(n14618) );
  XNOR2_X1 U16362 ( .A(n14619), .B(n14618), .ZN(SUB_1596_U4) );
  AOI21_X1 U16363 ( .B1(n14622), .B2(n14621), .A(n14620), .ZN(n14637) );
  OAI22_X1 U16364 ( .A1(n15139), .A2(n6725), .B1(n15168), .B2(n14624), .ZN(
        n14634) );
  AOI21_X1 U16365 ( .B1(n14627), .B2(n14626), .A(n14625), .ZN(n14632) );
  AOI21_X1 U16366 ( .B1(n14630), .B2(n14629), .A(n14628), .ZN(n14631) );
  OAI22_X1 U16367 ( .A1(n14632), .A2(n15136), .B1(n14631), .B2(n15131), .ZN(
        n14633) );
  NOR3_X1 U16368 ( .A1(n14635), .A2(n14634), .A3(n14633), .ZN(n14636) );
  OAI21_X1 U16369 ( .B1(n14637), .B2(n15163), .A(n14636), .ZN(P3_U3197) );
  AOI21_X1 U16370 ( .B1(n14640), .B2(n14639), .A(n14638), .ZN(n14657) );
  INV_X1 U16371 ( .A(n14641), .ZN(n14643) );
  NAND2_X1 U16372 ( .A1(n14643), .A2(n14642), .ZN(n14644) );
  XNOR2_X1 U16373 ( .A(n14645), .B(n14644), .ZN(n14651) );
  NAND2_X1 U16374 ( .A1(n15153), .A2(n14646), .ZN(n14648) );
  OAI211_X1 U16375 ( .C1(n14649), .C2(n15168), .A(n14648), .B(n14647), .ZN(
        n14650) );
  AOI21_X1 U16376 ( .B1(n14651), .B2(n15155), .A(n14650), .ZN(n14656) );
  AOI21_X1 U16377 ( .B1(n6545), .B2(n14653), .A(n14652), .ZN(n14654) );
  OR2_X1 U16378 ( .A1(n14654), .A2(n15136), .ZN(n14655) );
  OAI211_X1 U16379 ( .C1(n14657), .C2(n15163), .A(n14656), .B(n14655), .ZN(
        P3_U3198) );
  OR2_X1 U16380 ( .A1(n14658), .A2(n15261), .ZN(n14659) );
  INV_X1 U16381 ( .A(P3_REG1_REG_31__SCAN_IN), .ZN(n14660) );
  AOI22_X1 U16382 ( .A1(n15281), .A2(n14685), .B1(n14660), .B2(n15279), .ZN(
        P3_U3490) );
  OAI21_X1 U16383 ( .B1(n14662), .B2(n15261), .A(n14661), .ZN(n14687) );
  OAI22_X1 U16384 ( .A1(n15279), .A2(n14687), .B1(P3_REG1_REG_30__SCAN_IN), 
        .B2(n15281), .ZN(n14663) );
  INV_X1 U16385 ( .A(n14663), .ZN(P3_U3489) );
  NOR2_X1 U16386 ( .A1(n14664), .A2(n14680), .ZN(n14666) );
  AOI211_X1 U16387 ( .C1(n15224), .C2(n14667), .A(n14666), .B(n14665), .ZN(
        n14689) );
  INV_X1 U16388 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n14668) );
  AOI22_X1 U16389 ( .A1(n15281), .A2(n14689), .B1(n14668), .B2(n15279), .ZN(
        P3_U3473) );
  NOR2_X1 U16390 ( .A1(n14669), .A2(n15261), .ZN(n14671) );
  AOI211_X1 U16391 ( .C1(n14672), .C2(n15214), .A(n14671), .B(n14670), .ZN(
        n14691) );
  AOI22_X1 U16392 ( .A1(n15281), .A2(n14691), .B1(n14673), .B2(n15279), .ZN(
        P3_U3472) );
  NOR2_X1 U16393 ( .A1(n14674), .A2(n15261), .ZN(n14676) );
  AOI211_X1 U16394 ( .C1(n15214), .C2(n14677), .A(n14676), .B(n14675), .ZN(
        n14693) );
  INV_X1 U16395 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n14678) );
  AOI22_X1 U16396 ( .A1(n15281), .A2(n14693), .B1(n14678), .B2(n15279), .ZN(
        P3_U3471) );
  OAI22_X1 U16397 ( .A1(n14681), .A2(n14680), .B1(n15261), .B2(n14679), .ZN(
        n14682) );
  NOR2_X1 U16398 ( .A1(n14683), .A2(n14682), .ZN(n14695) );
  AOI22_X1 U16399 ( .A1(n15281), .A2(n14695), .B1(n14684), .B2(n15279), .ZN(
        P3_U3470) );
  INV_X1 U16400 ( .A(P3_REG0_REG_31__SCAN_IN), .ZN(n14686) );
  AOI22_X1 U16401 ( .A1(n15268), .A2(n14686), .B1(n14685), .B2(n15266), .ZN(
        P3_U3458) );
  OAI22_X1 U16402 ( .A1(n15266), .A2(P3_REG0_REG_30__SCAN_IN), .B1(n14687), 
        .B2(n15268), .ZN(n14688) );
  INV_X1 U16403 ( .A(n14688), .ZN(P3_U3457) );
  INV_X1 U16404 ( .A(P3_REG0_REG_14__SCAN_IN), .ZN(n14690) );
  AOI22_X1 U16405 ( .A1(n15268), .A2(n14690), .B1(n14689), .B2(n15266), .ZN(
        P3_U3432) );
  INV_X1 U16406 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n14692) );
  AOI22_X1 U16407 ( .A1(n15268), .A2(n14692), .B1(n14691), .B2(n15266), .ZN(
        P3_U3429) );
  INV_X1 U16408 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n14694) );
  AOI22_X1 U16409 ( .A1(n15268), .A2(n14694), .B1(n14693), .B2(n15266), .ZN(
        P3_U3426) );
  INV_X1 U16410 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n14696) );
  AOI22_X1 U16411 ( .A1(n15268), .A2(n14696), .B1(n14695), .B2(n15266), .ZN(
        P3_U3423) );
  XNOR2_X1 U16412 ( .A(n14697), .B(n14705), .ZN(n14700) );
  INV_X1 U16413 ( .A(n14698), .ZN(n14699) );
  AOI21_X1 U16414 ( .B1(n14700), .B2(n15064), .A(n14699), .ZN(n14733) );
  AOI222_X1 U16415 ( .A1(n14702), .A2(n14715), .B1(n14701), .B2(n14979), .C1(
        P2_REG2_REG_14__SCAN_IN), .C2(n15005), .ZN(n14710) );
  AOI21_X1 U16416 ( .B1(n14705), .B2(n14704), .A(n14703), .ZN(n14738) );
  OAI211_X1 U16417 ( .C1(n14735), .C2(n6951), .A(n10086), .B(n14707), .ZN(
        n14734) );
  INV_X1 U16418 ( .A(n14734), .ZN(n14708) );
  AOI22_X1 U16419 ( .A1(n14738), .A2(n14723), .B1(n14722), .B2(n14708), .ZN(
        n14709) );
  OAI211_X1 U16420 ( .C1(n15005), .C2(n14733), .A(n14710), .B(n14709), .ZN(
        P2_U3251) );
  XOR2_X1 U16421 ( .A(n14711), .B(n14717), .Z(n14713) );
  AOI21_X1 U16422 ( .B1(n14713), .B2(n15064), .A(n14712), .ZN(n14748) );
  AOI222_X1 U16423 ( .A1(n14716), .A2(n14715), .B1(n14714), .B2(n14979), .C1(
        P2_REG2_REG_12__SCAN_IN), .C2(n15005), .ZN(n14725) );
  XNOR2_X1 U16424 ( .A(n14718), .B(n14717), .ZN(n14753) );
  OAI211_X1 U16425 ( .C1(n14750), .C2(n14720), .A(n10086), .B(n14719), .ZN(
        n14749) );
  INV_X1 U16426 ( .A(n14749), .ZN(n14721) );
  AOI22_X1 U16427 ( .A1(n14753), .A2(n14723), .B1(n14722), .B2(n14721), .ZN(
        n14724) );
  OAI211_X1 U16428 ( .C1(n15005), .C2(n14748), .A(n14725), .B(n14724), .ZN(
        P2_U3253) );
  OAI211_X1 U16429 ( .C1(n14728), .C2(n15077), .A(n14727), .B(n14726), .ZN(
        n14729) );
  AOI211_X1 U16430 ( .C1(n14731), .C2(n15035), .A(n14730), .B(n14729), .ZN(
        n14756) );
  INV_X1 U16431 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n14732) );
  AOI22_X1 U16432 ( .A1(n15096), .A2(n14756), .B1(n14732), .B2(n15094), .ZN(
        P2_U3514) );
  INV_X1 U16433 ( .A(n14733), .ZN(n14737) );
  OAI21_X1 U16434 ( .B1(n14735), .B2(n15077), .A(n14734), .ZN(n14736) );
  AOI211_X1 U16435 ( .C1(n14738), .C2(n15035), .A(n14737), .B(n14736), .ZN(
        n14758) );
  AOI22_X1 U16436 ( .A1(n15096), .A2(n14758), .B1(n14739), .B2(n15094), .ZN(
        P2_U3513) );
  NOR2_X1 U16437 ( .A1(n14740), .A2(n14997), .ZN(n14745) );
  OAI211_X1 U16438 ( .C1(n14743), .C2(n15077), .A(n14742), .B(n14741), .ZN(
        n14744) );
  AOI211_X1 U16439 ( .C1(n14746), .C2(n15035), .A(n14745), .B(n14744), .ZN(
        n14760) );
  AOI22_X1 U16440 ( .A1(n15096), .A2(n14760), .B1(n14747), .B2(n15094), .ZN(
        P2_U3512) );
  INV_X1 U16441 ( .A(n14748), .ZN(n14752) );
  OAI21_X1 U16442 ( .B1(n14750), .B2(n15077), .A(n14749), .ZN(n14751) );
  AOI211_X1 U16443 ( .C1(n14753), .C2(n15035), .A(n14752), .B(n14751), .ZN(
        n14762) );
  AOI22_X1 U16444 ( .A1(n15096), .A2(n14762), .B1(n14754), .B2(n15094), .ZN(
        P2_U3511) );
  INV_X1 U16445 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n14755) );
  AOI22_X1 U16446 ( .A1(n15066), .A2(n14756), .B1(n14755), .B2(n15083), .ZN(
        P2_U3475) );
  INV_X1 U16447 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n14757) );
  AOI22_X1 U16448 ( .A1(n15066), .A2(n14758), .B1(n14757), .B2(n15083), .ZN(
        P2_U3472) );
  INV_X1 U16449 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n14759) );
  AOI22_X1 U16450 ( .A1(n15066), .A2(n14760), .B1(n14759), .B2(n15083), .ZN(
        P2_U3469) );
  INV_X1 U16451 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n14761) );
  AOI22_X1 U16452 ( .A1(n15066), .A2(n14762), .B1(n14761), .B2(n15083), .ZN(
        P2_U3466) );
  OAI21_X1 U16453 ( .B1(n14765), .B2(n14764), .A(n14763), .ZN(n14767) );
  XOR2_X1 U16454 ( .A(n14767), .B(n14766), .Z(SUB_1596_U69) );
  AOI21_X1 U16455 ( .B1(n14770), .B2(n14769), .A(n14768), .ZN(n14771) );
  XOR2_X1 U16456 ( .A(n14771), .B(P2_ADDR_REG_12__SCAN_IN), .Z(SUB_1596_U68)
         );
  OAI21_X1 U16457 ( .B1(n14773), .B2(n6638), .A(n14772), .ZN(n14774) );
  XOR2_X1 U16458 ( .A(n14774), .B(n14900), .Z(SUB_1596_U67) );
  NOR2_X1 U16459 ( .A1(n14776), .A2(n14775), .ZN(n14777) );
  XOR2_X1 U16460 ( .A(P2_ADDR_REG_14__SCAN_IN), .B(n14777), .Z(SUB_1596_U66)
         );
  AOI21_X1 U16461 ( .B1(n14780), .B2(n14779), .A(n14778), .ZN(n14781) );
  XOR2_X1 U16462 ( .A(n14781), .B(P2_ADDR_REG_15__SCAN_IN), .Z(SUB_1596_U65)
         );
  XNOR2_X1 U16463 ( .A(P2_ADDR_REG_16__SCAN_IN), .B(n6480), .ZN(SUB_1596_U64)
         );
  AND3_X1 U16464 ( .A1(n14785), .A2(n14784), .A3(n14783), .ZN(n14786) );
  NOR3_X1 U16465 ( .A1(n14809), .A2(n14787), .A3(n14786), .ZN(n14797) );
  INV_X1 U16466 ( .A(n14788), .ZN(n14793) );
  NOR3_X1 U16467 ( .A1(n14791), .A2(n14790), .A3(n14789), .ZN(n14792) );
  NOR3_X1 U16468 ( .A1(n14807), .A2(n14793), .A3(n14792), .ZN(n14796) );
  NOR2_X1 U16469 ( .A1(n14811), .A2(n14794), .ZN(n14795) );
  NOR4_X1 U16470 ( .A1(n14798), .A2(n14797), .A3(n14796), .A4(n14795), .ZN(
        n14800) );
  OAI211_X1 U16471 ( .C1(n14815), .C2(n14801), .A(n14800), .B(n14799), .ZN(
        P1_U3247) );
  AOI21_X1 U16472 ( .B1(P1_REG1_REG_15__SCAN_IN), .B2(n14803), .A(n14802), 
        .ZN(n14808) );
  AOI21_X1 U16473 ( .B1(P1_REG2_REG_15__SCAN_IN), .B2(n14805), .A(n14804), 
        .ZN(n14806) );
  OAI222_X1 U16474 ( .A1(n14811), .A2(n14810), .B1(n14809), .B2(n14808), .C1(
        n14807), .C2(n14806), .ZN(n14812) );
  INV_X1 U16475 ( .A(n14812), .ZN(n14814) );
  OAI211_X1 U16476 ( .C1(n14816), .C2(n14815), .A(n14814), .B(n14813), .ZN(
        P1_U3258) );
  NAND2_X1 U16477 ( .A1(n14818), .A2(n14817), .ZN(n14822) );
  AOI22_X1 U16478 ( .A1(n14830), .A2(P1_REG2_REG_7__SCAN_IN), .B1(n14820), 
        .B2(n14819), .ZN(n14821) );
  OAI211_X1 U16479 ( .C1(n14824), .C2(n14823), .A(n14822), .B(n14821), .ZN(
        n14825) );
  AOI21_X1 U16480 ( .B1(n14827), .B2(n14826), .A(n14825), .ZN(n14828) );
  OAI21_X1 U16481 ( .B1(n14830), .B2(n14829), .A(n14828), .ZN(P1_U3286) );
  AND2_X1 U16482 ( .A1(n14831), .A2(P1_D_REG_31__SCAN_IN), .ZN(P1_U3294) );
  AND2_X1 U16483 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n14831), .ZN(P1_U3295) );
  AND2_X1 U16484 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n14831), .ZN(P1_U3296) );
  AND2_X1 U16485 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n14831), .ZN(P1_U3297) );
  AND2_X1 U16486 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n14831), .ZN(P1_U3298) );
  AND2_X1 U16487 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n14831), .ZN(P1_U3299) );
  AND2_X1 U16488 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n14831), .ZN(P1_U3300) );
  AND2_X1 U16489 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n14831), .ZN(P1_U3301) );
  AND2_X1 U16490 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n14831), .ZN(P1_U3302) );
  AND2_X1 U16491 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n14831), .ZN(P1_U3303) );
  AND2_X1 U16492 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n14831), .ZN(P1_U3304) );
  AND2_X1 U16493 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n14831), .ZN(P1_U3305) );
  AND2_X1 U16494 ( .A1(n14831), .A2(P1_D_REG_19__SCAN_IN), .ZN(P1_U3306) );
  AND2_X1 U16495 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n14831), .ZN(P1_U3307) );
  AND2_X1 U16496 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n14831), .ZN(P1_U3308) );
  AND2_X1 U16497 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n14831), .ZN(P1_U3309) );
  AND2_X1 U16498 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n14831), .ZN(P1_U3310) );
  AND2_X1 U16499 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n14831), .ZN(P1_U3311) );
  AND2_X1 U16500 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n14831), .ZN(P1_U3312) );
  AND2_X1 U16501 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n14831), .ZN(P1_U3313) );
  AND2_X1 U16502 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n14831), .ZN(P1_U3314) );
  AND2_X1 U16503 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n14831), .ZN(P1_U3315) );
  AND2_X1 U16504 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n14831), .ZN(P1_U3316) );
  AND2_X1 U16505 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n14831), .ZN(P1_U3317) );
  AND2_X1 U16506 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n14831), .ZN(P1_U3318) );
  AND2_X1 U16507 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n14831), .ZN(P1_U3319) );
  AND2_X1 U16508 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n14831), .ZN(P1_U3320) );
  AND2_X1 U16509 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n14831), .ZN(P1_U3321) );
  AND2_X1 U16510 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n14831), .ZN(P1_U3322) );
  AND2_X1 U16511 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n14831), .ZN(P1_U3323) );
  OAI211_X1 U16512 ( .C1(n6691), .C2(n14843), .A(n14833), .B(n14832), .ZN(
        n14835) );
  AOI21_X1 U16513 ( .B1(n14848), .B2(n14836), .A(n14835), .ZN(n14851) );
  AOI22_X1 U16514 ( .A1(n14849), .A2(n14851), .B1(n7479), .B2(n6786), .ZN(
        P1_U3465) );
  OAI211_X1 U16515 ( .C1(n14839), .C2(n14843), .A(n14838), .B(n14837), .ZN(
        n14840) );
  AOI21_X1 U16516 ( .B1(n14848), .B2(n14841), .A(n14840), .ZN(n14853) );
  AOI22_X1 U16517 ( .A1(n14849), .A2(n14853), .B1(n7571), .B2(n6786), .ZN(
        P1_U3471) );
  OAI21_X1 U16518 ( .B1(n14844), .B2(n14843), .A(n14842), .ZN(n14846) );
  AOI211_X1 U16519 ( .C1(n14848), .C2(n14847), .A(n14846), .B(n14845), .ZN(
        n14855) );
  AOI22_X1 U16520 ( .A1(n14849), .A2(n14855), .B1(n7685), .B2(n6786), .ZN(
        P1_U3483) );
  AOI22_X1 U16521 ( .A1(n14856), .A2(n14851), .B1(n14850), .B2(n14854), .ZN(
        P1_U3530) );
  AOI22_X1 U16522 ( .A1(n14856), .A2(n14853), .B1(n14852), .B2(n14854), .ZN(
        P1_U3532) );
  AOI22_X1 U16523 ( .A1(n14856), .A2(n14855), .B1(n10022), .B2(n14854), .ZN(
        P1_U3536) );
  NOR2_X1 U16524 ( .A1(n14954), .A2(P2_U3947), .ZN(P2_U3087) );
  OAI21_X1 U16525 ( .B1(n14870), .B2(n14857), .A(P2_STATE_REG_SCAN_IN), .ZN(
        n14858) );
  OAI21_X1 U16526 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(P2_STATE_REG_SCAN_IN), 
        .A(n14858), .ZN(n14868) );
  OAI211_X1 U16527 ( .C1(n14861), .C2(n14860), .A(n14961), .B(n14859), .ZN(
        n14867) );
  NAND2_X1 U16528 ( .A1(P2_ADDR_REG_1__SCAN_IN), .A2(n14954), .ZN(n14866) );
  OAI211_X1 U16529 ( .C1(n14864), .C2(n14863), .A(n14956), .B(n14862), .ZN(
        n14865) );
  NAND4_X1 U16530 ( .A1(n14868), .A2(n14867), .A3(n14866), .A4(n14865), .ZN(
        P2_U3215) );
  OAI21_X1 U16531 ( .B1(n14870), .B2(n14869), .A(P2_STATE_REG_SCAN_IN), .ZN(
        n14871) );
  OAI21_X1 U16532 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(P2_STATE_REG_SCAN_IN), 
        .A(n14871), .ZN(n14881) );
  OAI211_X1 U16533 ( .C1(n14874), .C2(n14873), .A(n14961), .B(n14872), .ZN(
        n14880) );
  OAI211_X1 U16534 ( .C1(n14877), .C2(n14876), .A(n14956), .B(n14875), .ZN(
        n14879) );
  NAND2_X1 U16535 ( .A1(P2_ADDR_REG_4__SCAN_IN), .A2(n14954), .ZN(n14878) );
  NAND4_X1 U16536 ( .A1(n14881), .A2(n14880), .A3(n14879), .A4(n14878), .ZN(
        P2_U3218) );
  NOR2_X1 U16537 ( .A1(n14883), .A2(n14882), .ZN(n14884) );
  OAI21_X1 U16538 ( .B1(n14885), .B2(n14884), .A(n14956), .ZN(n14892) );
  AND3_X1 U16539 ( .A1(n14888), .A2(n14887), .A3(n14886), .ZN(n14889) );
  OAI21_X1 U16540 ( .B1(n14890), .B2(n14889), .A(n14961), .ZN(n14891) );
  OAI211_X1 U16541 ( .C1(n14894), .C2(n14893), .A(n14892), .B(n14891), .ZN(
        n14895) );
  INV_X1 U16542 ( .A(n14895), .ZN(n14897) );
  NAND2_X1 U16543 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3088), .ZN(n14896)
         );
  OAI211_X1 U16544 ( .C1(n14898), .C2(n14901), .A(n14897), .B(n14896), .ZN(
        P2_U3226) );
  OAI21_X1 U16545 ( .B1(n14901), .B2(n14900), .A(n14899), .ZN(n14902) );
  AOI21_X1 U16546 ( .B1(n14903), .B2(n14959), .A(n14902), .ZN(n14912) );
  OAI211_X1 U16547 ( .C1(n14906), .C2(n14905), .A(n14904), .B(n14961), .ZN(
        n14911) );
  OAI211_X1 U16548 ( .C1(n14909), .C2(n14908), .A(n14907), .B(n14956), .ZN(
        n14910) );
  NAND3_X1 U16549 ( .A1(n14912), .A2(n14911), .A3(n14910), .ZN(P2_U3227) );
  AOI22_X1 U16550 ( .A1(n14954), .A2(P2_ADDR_REG_14__SCAN_IN), .B1(
        P2_REG3_REG_14__SCAN_IN), .B2(P2_U3088), .ZN(n14922) );
  OAI211_X1 U16551 ( .C1(n14914), .C2(P2_REG2_REG_14__SCAN_IN), .A(n14961), 
        .B(n14913), .ZN(n14921) );
  OAI211_X1 U16552 ( .C1(n14917), .C2(n14916), .A(n14915), .B(n14956), .ZN(
        n14920) );
  NAND2_X1 U16553 ( .A1(n14959), .A2(n14918), .ZN(n14919) );
  NAND4_X1 U16554 ( .A1(n14922), .A2(n14921), .A3(n14920), .A4(n14919), .ZN(
        P2_U3228) );
  AOI22_X1 U16555 ( .A1(n14954), .A2(P2_ADDR_REG_15__SCAN_IN), .B1(
        P2_REG3_REG_15__SCAN_IN), .B2(P2_U3088), .ZN(n14931) );
  NAND2_X1 U16556 ( .A1(n14959), .A2(n14923), .ZN(n14930) );
  OAI211_X1 U16557 ( .C1(n14925), .C2(P2_REG2_REG_15__SCAN_IN), .A(n14961), 
        .B(n14924), .ZN(n14929) );
  OAI211_X1 U16558 ( .C1(P2_REG1_REG_15__SCAN_IN), .C2(n14927), .A(n14956), 
        .B(n14926), .ZN(n14928) );
  NAND4_X1 U16559 ( .A1(n14931), .A2(n14930), .A3(n14929), .A4(n14928), .ZN(
        P2_U3229) );
  AOI22_X1 U16560 ( .A1(n14954), .A2(P2_ADDR_REG_16__SCAN_IN), .B1(
        P2_REG3_REG_16__SCAN_IN), .B2(P2_U3088), .ZN(n14942) );
  OAI211_X1 U16561 ( .C1(n14934), .C2(n14933), .A(n14961), .B(n14932), .ZN(
        n14941) );
  NAND2_X1 U16562 ( .A1(n14959), .A2(n14935), .ZN(n14940) );
  OAI211_X1 U16563 ( .C1(n14938), .C2(n14937), .A(n14956), .B(n14936), .ZN(
        n14939) );
  NAND4_X1 U16564 ( .A1(n14942), .A2(n14941), .A3(n14940), .A4(n14939), .ZN(
        P2_U3230) );
  AOI22_X1 U16565 ( .A1(n14954), .A2(P2_ADDR_REG_17__SCAN_IN), .B1(
        P2_REG3_REG_17__SCAN_IN), .B2(P2_U3088), .ZN(n14953) );
  NAND2_X1 U16566 ( .A1(n14959), .A2(n14943), .ZN(n14952) );
  OAI211_X1 U16567 ( .C1(n14946), .C2(n14945), .A(n14944), .B(n14956), .ZN(
        n14951) );
  OAI211_X1 U16568 ( .C1(n14949), .C2(n14948), .A(n14947), .B(n14961), .ZN(
        n14950) );
  NAND4_X1 U16569 ( .A1(n14953), .A2(n14952), .A3(n14951), .A4(n14950), .ZN(
        P2_U3231) );
  AOI22_X1 U16570 ( .A1(n14954), .A2(P2_ADDR_REG_18__SCAN_IN), .B1(
        P2_REG3_REG_18__SCAN_IN), .B2(P2_U3088), .ZN(n14967) );
  OAI211_X1 U16571 ( .C1(P2_REG1_REG_18__SCAN_IN), .C2(n14957), .A(n14956), 
        .B(n14955), .ZN(n14966) );
  NAND2_X1 U16572 ( .A1(n14959), .A2(n14958), .ZN(n14965) );
  AND2_X1 U16573 ( .A1(n14960), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n14963) );
  OAI21_X1 U16574 ( .B1(n14963), .B2(n14962), .A(n14961), .ZN(n14964) );
  NAND4_X1 U16575 ( .A1(n14967), .A2(n14966), .A3(n14965), .A4(n14964), .ZN(
        P2_U3232) );
  NOR2_X1 U16576 ( .A1(n14968), .A2(n6701), .ZN(n14977) );
  INV_X1 U16577 ( .A(n14971), .ZN(n14969) );
  XNOR2_X1 U16578 ( .A(n14970), .B(n14969), .ZN(n15048) );
  XNOR2_X1 U16579 ( .A(n14972), .B(n14971), .ZN(n14974) );
  AOI21_X1 U16580 ( .B1(n14974), .B2(n15064), .A(n14973), .ZN(n15053) );
  OAI21_X1 U16581 ( .B1(n15048), .B2(n10347), .A(n15053), .ZN(n14975) );
  MUX2_X1 U16582 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n14975), .S(n15002), .Z(
        n14976) );
  AOI211_X1 U16583 ( .C1(n14979), .C2(n14978), .A(n14977), .B(n14976), .ZN(
        n14987) );
  AOI21_X1 U16584 ( .B1(n14980), .B2(n15049), .A(n12605), .ZN(n14982) );
  NAND2_X1 U16585 ( .A1(n14982), .A2(n14981), .ZN(n15051) );
  OAI22_X1 U16586 ( .A1(n14984), .A2(n15048), .B1(n14983), .B2(n15051), .ZN(
        n14985) );
  INV_X1 U16587 ( .A(n14985), .ZN(n14986) );
  NAND2_X1 U16588 ( .A1(n14987), .A2(n14986), .ZN(P2_U3261) );
  OR2_X1 U16589 ( .A1(n15020), .A2(n14988), .ZN(n14994) );
  INV_X1 U16590 ( .A(n14989), .ZN(n14991) );
  NAND2_X1 U16591 ( .A1(n14991), .A2(n14990), .ZN(n15018) );
  OR2_X1 U16592 ( .A1(n15018), .A2(n14992), .ZN(n14993) );
  OAI211_X1 U16593 ( .C1(n14996), .C2(n14995), .A(n14994), .B(n14993), .ZN(
        n15001) );
  AND2_X1 U16594 ( .A1(n10347), .A2(n14997), .ZN(n14998) );
  OR2_X1 U16595 ( .A1(n15020), .A2(n14998), .ZN(n15000) );
  NAND2_X1 U16596 ( .A1(n15000), .A2(n14999), .ZN(n15017) );
  NOR2_X1 U16597 ( .A1(n15001), .A2(n15017), .ZN(n15003) );
  AOI22_X1 U16598 ( .A1(n15005), .A2(n15004), .B1(n15003), .B2(n15002), .ZN(
        P2_U3265) );
  AND2_X1 U16599 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n15010), .ZN(P2_U3266) );
  AND2_X1 U16600 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n15010), .ZN(P2_U3267) );
  AND2_X1 U16601 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n15010), .ZN(P2_U3268) );
  AND2_X1 U16602 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n15010), .ZN(P2_U3269) );
  AND2_X1 U16603 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n15010), .ZN(P2_U3270) );
  AND2_X1 U16604 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n15010), .ZN(P2_U3271) );
  AND2_X1 U16605 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n15010), .ZN(P2_U3272) );
  NOR2_X1 U16606 ( .A1(n15009), .A2(n15007), .ZN(P2_U3273) );
  AND2_X1 U16607 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n15010), .ZN(P2_U3274) );
  AND2_X1 U16608 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n15010), .ZN(P2_U3275) );
  AND2_X1 U16609 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n15010), .ZN(P2_U3276) );
  AND2_X1 U16610 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n15010), .ZN(P2_U3277) );
  AND2_X1 U16611 ( .A1(n15010), .A2(P2_D_REG_19__SCAN_IN), .ZN(P2_U3278) );
  AND2_X1 U16612 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n15010), .ZN(P2_U3279) );
  AND2_X1 U16613 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n15010), .ZN(P2_U3280) );
  NOR2_X1 U16614 ( .A1(n15009), .A2(n15008), .ZN(P2_U3281) );
  AND2_X1 U16615 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n15010), .ZN(P2_U3282) );
  AND2_X1 U16616 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n15010), .ZN(P2_U3283) );
  AND2_X1 U16617 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n15010), .ZN(P2_U3284) );
  AND2_X1 U16618 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n15010), .ZN(P2_U3285) );
  AND2_X1 U16619 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n15010), .ZN(P2_U3286) );
  AND2_X1 U16620 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n15010), .ZN(P2_U3287) );
  AND2_X1 U16621 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n15010), .ZN(P2_U3288) );
  AND2_X1 U16622 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n15010), .ZN(P2_U3289) );
  AND2_X1 U16623 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n15010), .ZN(P2_U3290) );
  AND2_X1 U16624 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n15010), .ZN(P2_U3291) );
  AND2_X1 U16625 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n15010), .ZN(P2_U3292) );
  AND2_X1 U16626 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n15010), .ZN(P2_U3293) );
  AND2_X1 U16627 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n15010), .ZN(P2_U3294) );
  AND2_X1 U16628 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n15010), .ZN(P2_U3295) );
  AOI22_X1 U16629 ( .A1(n15016), .A2(n15012), .B1(n15011), .B2(n15013), .ZN(
        P2_U3416) );
  AOI22_X1 U16630 ( .A1(n15016), .A2(n15015), .B1(n15014), .B2(n15013), .ZN(
        P2_U3417) );
  INV_X1 U16631 ( .A(n15017), .ZN(n15019) );
  OAI211_X1 U16632 ( .C1(n15020), .C2(n15076), .A(n15019), .B(n15018), .ZN(
        n15085) );
  OAI22_X1 U16633 ( .A1(n15083), .A2(n15085), .B1(P2_REG0_REG_0__SCAN_IN), 
        .B2(n15066), .ZN(n15021) );
  INV_X1 U16634 ( .A(n15021), .ZN(P2_U3430) );
  INV_X1 U16635 ( .A(n15022), .ZN(n15023) );
  AOI21_X1 U16636 ( .B1(n10347), .B2(n15076), .A(n15023), .ZN(n15028) );
  OAI211_X1 U16637 ( .C1(n15026), .C2(n15077), .A(n15025), .B(n15024), .ZN(
        n15027) );
  NOR2_X1 U16638 ( .A1(n15028), .A2(n15027), .ZN(n15087) );
  INV_X1 U16639 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n15029) );
  AOI22_X1 U16640 ( .A1(n15066), .A2(n15087), .B1(n15029), .B2(n15083), .ZN(
        P2_U3433) );
  INV_X1 U16641 ( .A(n15030), .ZN(n15031) );
  OAI21_X1 U16642 ( .B1(n6747), .B2(n15077), .A(n15031), .ZN(n15034) );
  INV_X1 U16643 ( .A(n15032), .ZN(n15033) );
  AOI211_X1 U16644 ( .C1(n15036), .C2(n15035), .A(n15034), .B(n15033), .ZN(
        n15088) );
  INV_X1 U16645 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n15037) );
  AOI22_X1 U16646 ( .A1(n15066), .A2(n15088), .B1(n15037), .B2(n15083), .ZN(
        P2_U3436) );
  INV_X1 U16647 ( .A(n15038), .ZN(n15041) );
  INV_X1 U16648 ( .A(n15039), .ZN(n15040) );
  OAI211_X1 U16649 ( .C1(n15042), .C2(n15077), .A(n15041), .B(n15040), .ZN(
        n15045) );
  AOI21_X1 U16650 ( .B1(n10347), .B2(n15076), .A(n15043), .ZN(n15044) );
  AOI211_X1 U16651 ( .C1(n15064), .C2(n15046), .A(n15045), .B(n15044), .ZN(
        n15089) );
  INV_X1 U16652 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n15047) );
  AOI22_X1 U16653 ( .A1(n15066), .A2(n15089), .B1(n15047), .B2(n15083), .ZN(
        P2_U3439) );
  OR2_X1 U16654 ( .A1(n15048), .A2(n15061), .ZN(n15054) );
  NAND2_X1 U16655 ( .A1(n15049), .A2(n15069), .ZN(n15050) );
  AND2_X1 U16656 ( .A1(n15051), .A2(n15050), .ZN(n15052) );
  INV_X1 U16657 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n15055) );
  AOI22_X1 U16658 ( .A1(n15066), .A2(n15091), .B1(n15055), .B2(n15083), .ZN(
        P2_U3442) );
  AOI211_X1 U16659 ( .C1(n15069), .C2(n15058), .A(n15057), .B(n15056), .ZN(
        n15059) );
  OAI21_X1 U16660 ( .B1(n15061), .B2(n15060), .A(n15059), .ZN(n15062) );
  AOI21_X1 U16661 ( .B1(n15064), .B2(n15063), .A(n15062), .ZN(n15092) );
  INV_X1 U16662 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n15065) );
  AOI22_X1 U16663 ( .A1(n15066), .A2(n15092), .B1(n15065), .B2(n15083), .ZN(
        P2_U3445) );
  AOI21_X1 U16664 ( .B1(n15069), .B2(n15068), .A(n15067), .ZN(n15070) );
  OAI211_X1 U16665 ( .C1(n15072), .C2(n15076), .A(n15071), .B(n15070), .ZN(
        n15073) );
  INV_X1 U16666 ( .A(n15073), .ZN(n15093) );
  INV_X1 U16667 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n15074) );
  AOI22_X1 U16668 ( .A1(n15066), .A2(n15093), .B1(n15074), .B2(n15083), .ZN(
        P2_U3454) );
  AOI21_X1 U16669 ( .B1(n10347), .B2(n15076), .A(n15075), .ZN(n15082) );
  NOR2_X1 U16670 ( .A1(n15078), .A2(n15077), .ZN(n15080) );
  NOR4_X1 U16671 ( .A1(n15082), .A2(n15081), .A3(n15080), .A4(n15079), .ZN(
        n15095) );
  INV_X1 U16672 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n15084) );
  AOI22_X1 U16673 ( .A1(n15066), .A2(n15095), .B1(n15084), .B2(n15083), .ZN(
        P2_U3463) );
  OAI22_X1 U16674 ( .A1(n15094), .A2(n15085), .B1(P2_REG1_REG_0__SCAN_IN), 
        .B2(n15096), .ZN(n15086) );
  INV_X1 U16675 ( .A(n15086), .ZN(P2_U3499) );
  AOI22_X1 U16676 ( .A1(n15096), .A2(n15087), .B1(n9676), .B2(n15094), .ZN(
        P2_U3500) );
  AOI22_X1 U16677 ( .A1(n15096), .A2(n15088), .B1(n9675), .B2(n15094), .ZN(
        P2_U3501) );
  AOI22_X1 U16678 ( .A1(n15096), .A2(n15089), .B1(n9674), .B2(n15094), .ZN(
        P2_U3502) );
  AOI22_X1 U16679 ( .A1(n15096), .A2(n15091), .B1(n15090), .B2(n15094), .ZN(
        P2_U3503) );
  AOI22_X1 U16680 ( .A1(n15096), .A2(n15092), .B1(n9682), .B2(n15094), .ZN(
        P2_U3504) );
  AOI22_X1 U16681 ( .A1(n15096), .A2(n15093), .B1(n9843), .B2(n15094), .ZN(
        P2_U3507) );
  AOI22_X1 U16682 ( .A1(n15096), .A2(n15095), .B1(n10103), .B2(n15094), .ZN(
        P2_U3510) );
  NOR2_X1 U16683 ( .A1(P3_U3897), .A2(n15097), .ZN(P3_U3150) );
  MUX2_X1 U16684 ( .A(n15099), .B(n13182), .S(n6490), .Z(n15100) );
  NOR2_X1 U16685 ( .A1(n15100), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n15102) );
  NAND3_X1 U16686 ( .A1(n15163), .A2(n15136), .A3(n15131), .ZN(n15101) );
  OAI21_X1 U16687 ( .B1(n15103), .B2(n15102), .A(n15101), .ZN(n15108) );
  INV_X1 U16688 ( .A(P3_REG3_REG_0__SCAN_IN), .ZN(n15104) );
  OAI22_X1 U16689 ( .A1(n15139), .A2(n15105), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n15104), .ZN(n15106) );
  INV_X1 U16690 ( .A(n15106), .ZN(n15107) );
  OAI211_X1 U16691 ( .C1(n15109), .C2(n15168), .A(n15108), .B(n15107), .ZN(
        P3_U3182) );
  AOI21_X1 U16692 ( .B1(n6649), .B2(n15111), .A(n15110), .ZN(n15115) );
  AOI21_X1 U16693 ( .B1(n6650), .B2(n15113), .A(n15112), .ZN(n15114) );
  OAI22_X1 U16694 ( .A1(n15115), .A2(n15163), .B1(n15136), .B2(n15114), .ZN(
        n15121) );
  NAND3_X1 U16695 ( .A1(n15118), .A2(n15117), .A3(n15116), .ZN(n15119) );
  AOI21_X1 U16696 ( .B1(n15130), .B2(n15119), .A(n15131), .ZN(n15120) );
  AOI211_X1 U16697 ( .C1(n15153), .C2(n15122), .A(n15121), .B(n15120), .ZN(
        n15124) );
  OAI211_X1 U16698 ( .C1(n15125), .C2(n15168), .A(n15124), .B(n15123), .ZN(
        P3_U3186) );
  AOI21_X1 U16699 ( .B1(n8382), .B2(n15126), .A(n6652), .ZN(n15127) );
  NOR2_X1 U16700 ( .A1(n15127), .A2(n15163), .ZN(n15142) );
  NAND3_X1 U16701 ( .A1(n15130), .A2(n15129), .A3(n15128), .ZN(n15132) );
  AOI21_X1 U16702 ( .B1(n15133), .B2(n15132), .A(n15131), .ZN(n15141) );
  AOI21_X1 U16703 ( .B1(n15135), .B2(n8381), .A(n15134), .ZN(n15137) );
  OAI22_X1 U16704 ( .A1(n15139), .A2(n15138), .B1(n15137), .B2(n15136), .ZN(
        n15140) );
  NOR3_X1 U16705 ( .A1(n15142), .A2(n15141), .A3(n15140), .ZN(n15144) );
  OAI211_X1 U16706 ( .C1(n15145), .C2(n15168), .A(n15144), .B(n15143), .ZN(
        P3_U3187) );
  AOI21_X1 U16707 ( .B1(n15147), .B2(n8402), .A(n15146), .ZN(n15164) );
  AND3_X1 U16708 ( .A1(n15150), .A2(n15149), .A3(n15148), .ZN(n15151) );
  OR2_X1 U16709 ( .A1(n15152), .A2(n15151), .ZN(n15156) );
  AOI22_X1 U16710 ( .A1(n15156), .A2(n15155), .B1(n15154), .B2(n15153), .ZN(
        n15162) );
  AND2_X1 U16711 ( .A1(n15157), .A2(n8401), .ZN(n15159) );
  OAI21_X1 U16712 ( .B1(n15160), .B2(n15159), .A(n15158), .ZN(n15161) );
  OAI211_X1 U16713 ( .C1(n15164), .C2(n15163), .A(n15162), .B(n15161), .ZN(
        n15165) );
  INV_X1 U16714 ( .A(n15165), .ZN(n15167) );
  OAI211_X1 U16715 ( .C1(n15169), .C2(n15168), .A(n15167), .B(n15166), .ZN(
        P3_U3189) );
  OAI21_X1 U16716 ( .B1(n15171), .B2(n15177), .A(n15170), .ZN(n15221) );
  OAI22_X1 U16717 ( .A1(n10444), .A2(n15173), .B1(n15172), .B2(n15197), .ZN(
        n15182) );
  NAND2_X1 U16718 ( .A1(n15193), .A2(n15176), .ZN(n15175) );
  NAND2_X1 U16719 ( .A1(n15175), .A2(n15174), .ZN(n15180) );
  NAND3_X1 U16720 ( .A1(n15193), .A2(n15177), .A3(n15176), .ZN(n15179) );
  AOI21_X1 U16721 ( .B1(n15180), .B2(n15179), .A(n15178), .ZN(n15181) );
  AOI211_X1 U16722 ( .C1(n15204), .C2(n15221), .A(n15182), .B(n15181), .ZN(
        n15183) );
  INV_X1 U16723 ( .A(n15183), .ZN(n15219) );
  INV_X1 U16724 ( .A(n15221), .ZN(n15187) );
  NOR2_X1 U16725 ( .A1(n15184), .A2(n15261), .ZN(n15220) );
  INV_X1 U16726 ( .A(n15220), .ZN(n15185) );
  OAI22_X1 U16727 ( .A1(n15187), .A2(n15186), .B1(n15206), .B2(n15185), .ZN(
        n15188) );
  AOI211_X1 U16728 ( .C1(n15208), .C2(P3_REG3_REG_2__SCAN_IN), .A(n15219), .B(
        n15188), .ZN(n15189) );
  AOI22_X1 U16729 ( .A1(n15213), .A2(n8352), .B1(n15189), .B2(n15211), .ZN(
        P3_U3231) );
  NAND2_X1 U16730 ( .A1(n15190), .A2(n15224), .ZN(n15216) );
  OR2_X1 U16731 ( .A1(n15202), .A2(n15191), .ZN(n15192) );
  NAND2_X1 U16732 ( .A1(n15193), .A2(n15192), .ZN(n15201) );
  NAND2_X1 U16733 ( .A1(n15195), .A2(n15194), .ZN(n15196) );
  OAI21_X1 U16734 ( .B1(n15198), .B2(n15197), .A(n15196), .ZN(n15199) );
  AOI21_X1 U16735 ( .B1(n15201), .B2(n15200), .A(n15199), .ZN(n15218) );
  XNOR2_X1 U16736 ( .A(n15203), .B(n15202), .ZN(n15215) );
  NAND2_X1 U16737 ( .A1(n15215), .A2(n15204), .ZN(n15205) );
  OAI211_X1 U16738 ( .C1(n15206), .C2(n15216), .A(n15218), .B(n15205), .ZN(
        n15207) );
  INV_X1 U16739 ( .A(n15207), .ZN(n15212) );
  AOI22_X1 U16740 ( .A1(n15209), .A2(n15215), .B1(P3_REG3_REG_1__SCAN_IN), 
        .B2(n15208), .ZN(n15210) );
  OAI221_X1 U16741 ( .B1(n15213), .B2(n15212), .C1(n15211), .C2(n8344), .A(
        n15210), .ZN(P3_U3232) );
  NAND2_X1 U16742 ( .A1(n15215), .A2(n15214), .ZN(n15217) );
  AND3_X1 U16743 ( .A1(n15218), .A2(n15217), .A3(n15216), .ZN(n15269) );
  AOI22_X1 U16744 ( .A1(n15268), .A2(n10236), .B1(n15269), .B2(n15266), .ZN(
        P3_U3393) );
  INV_X1 U16745 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n15222) );
  AOI211_X1 U16746 ( .C1(n15257), .C2(n15221), .A(n15220), .B(n15219), .ZN(
        n15270) );
  AOI22_X1 U16747 ( .A1(n15268), .A2(n15222), .B1(n15270), .B2(n15266), .ZN(
        P3_U3396) );
  INV_X1 U16748 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n15228) );
  AOI22_X1 U16749 ( .A1(n15225), .A2(n15257), .B1(n15224), .B2(n15223), .ZN(
        n15226) );
  AND2_X1 U16750 ( .A1(n15227), .A2(n15226), .ZN(n15271) );
  AOI22_X1 U16751 ( .A1(n15268), .A2(n15228), .B1(n15271), .B2(n15266), .ZN(
        P3_U3399) );
  INV_X1 U16752 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n15233) );
  OAI22_X1 U16753 ( .A1(n15230), .A2(n15262), .B1(n15261), .B2(n15229), .ZN(
        n15231) );
  NOR2_X1 U16754 ( .A1(n15232), .A2(n15231), .ZN(n15272) );
  AOI22_X1 U16755 ( .A1(n15268), .A2(n15233), .B1(n15272), .B2(n15266), .ZN(
        P3_U3402) );
  INV_X1 U16756 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n15238) );
  OAI22_X1 U16757 ( .A1(n15235), .A2(n15262), .B1(n15261), .B2(n15234), .ZN(
        n15236) );
  NOR2_X1 U16758 ( .A1(n15237), .A2(n15236), .ZN(n15273) );
  AOI22_X1 U16759 ( .A1(n15268), .A2(n15238), .B1(n15273), .B2(n15266), .ZN(
        P3_U3405) );
  INV_X1 U16760 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n15243) );
  OAI22_X1 U16761 ( .A1(n15240), .A2(n15262), .B1(n15239), .B2(n15261), .ZN(
        n15242) );
  NOR2_X1 U16762 ( .A1(n15242), .A2(n15241), .ZN(n15274) );
  AOI22_X1 U16763 ( .A1(n15268), .A2(n15243), .B1(n15274), .B2(n15266), .ZN(
        P3_U3408) );
  INV_X1 U16764 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n15248) );
  NOR2_X1 U16765 ( .A1(n15244), .A2(n15261), .ZN(n15246) );
  AOI211_X1 U16766 ( .C1(n15257), .C2(n15247), .A(n15246), .B(n15245), .ZN(
        n15275) );
  AOI22_X1 U16767 ( .A1(n15268), .A2(n15248), .B1(n15275), .B2(n15266), .ZN(
        P3_U3411) );
  INV_X1 U16768 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n15253) );
  OAI22_X1 U16769 ( .A1(n15250), .A2(n15262), .B1(n15249), .B2(n15261), .ZN(
        n15251) );
  NOR2_X1 U16770 ( .A1(n15252), .A2(n15251), .ZN(n15277) );
  AOI22_X1 U16771 ( .A1(n15268), .A2(n15253), .B1(n15277), .B2(n15266), .ZN(
        P3_U3414) );
  INV_X1 U16772 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n15259) );
  NOR2_X1 U16773 ( .A1(n15254), .A2(n15261), .ZN(n15256) );
  AOI211_X1 U16774 ( .C1(n15258), .C2(n15257), .A(n15256), .B(n15255), .ZN(
        n15278) );
  AOI22_X1 U16775 ( .A1(n15268), .A2(n15259), .B1(n15278), .B2(n15266), .ZN(
        P3_U3417) );
  INV_X1 U16776 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n15267) );
  OAI22_X1 U16777 ( .A1(n15263), .A2(n15262), .B1(n15261), .B2(n15260), .ZN(
        n15264) );
  NOR2_X1 U16778 ( .A1(n15265), .A2(n15264), .ZN(n15280) );
  AOI22_X1 U16779 ( .A1(n15268), .A2(n15267), .B1(n15280), .B2(n15266), .ZN(
        P3_U3420) );
  AOI22_X1 U16780 ( .A1(n15281), .A2(n15269), .B1(n8343), .B2(n15279), .ZN(
        P3_U3460) );
  AOI22_X1 U16781 ( .A1(n15281), .A2(n15270), .B1(n8351), .B2(n15279), .ZN(
        P3_U3461) );
  AOI22_X1 U16782 ( .A1(n15281), .A2(n15271), .B1(n8362), .B2(n15279), .ZN(
        P3_U3462) );
  AOI22_X1 U16783 ( .A1(n15281), .A2(n15272), .B1(n8471), .B2(n15279), .ZN(
        P3_U3463) );
  AOI22_X1 U16784 ( .A1(n15281), .A2(n15273), .B1(n8381), .B2(n15279), .ZN(
        P3_U3464) );
  AOI22_X1 U16785 ( .A1(n15281), .A2(n15274), .B1(n8474), .B2(n15279), .ZN(
        P3_U3465) );
  AOI22_X1 U16786 ( .A1(n15281), .A2(n15275), .B1(n8401), .B2(n15279), .ZN(
        P3_U3466) );
  AOI22_X1 U16787 ( .A1(n15281), .A2(n15277), .B1(n15276), .B2(n15279), .ZN(
        P3_U3467) );
  AOI22_X1 U16788 ( .A1(n15281), .A2(n15278), .B1(n8423), .B2(n15279), .ZN(
        P3_U3468) );
  AOI22_X1 U16789 ( .A1(n15281), .A2(n15280), .B1(n8429), .B2(n15279), .ZN(
        P3_U3469) );
  XOR2_X1 U16790 ( .A(n15283), .B(n15282), .Z(SUB_1596_U59) );
  XNOR2_X1 U16791 ( .A(n15284), .B(P2_ADDR_REG_5__SCAN_IN), .ZN(SUB_1596_U58)
         );
  AOI21_X1 U16792 ( .B1(n15286), .B2(n15285), .A(n15294), .ZN(SUB_1596_U53) );
  XOR2_X1 U16793 ( .A(n15287), .B(n15288), .Z(SUB_1596_U56) );
  OAI21_X1 U16794 ( .B1(n15291), .B2(n15290), .A(n15289), .ZN(n15292) );
  XOR2_X1 U16795 ( .A(n15292), .B(n9767), .Z(SUB_1596_U60) );
  XOR2_X1 U16796 ( .A(n15294), .B(n15293), .Z(SUB_1596_U5) );
  NAND3_X1 U7521 ( .A1(n7473), .A2(n6720), .A3(n7059), .ZN(n7486) );
  NAND2_X2 U9791 ( .A1(n7481), .A2(n14476), .ZN(n8205) );
  OR2_X1 U7302 ( .A1(n7623), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n7550) );
  CLKBUF_X3 U7304 ( .A(n9168), .Z(n6483) );
  CLKBUF_X1 U7463 ( .A(n8201), .Z(n8185) );
  CLKBUF_X1 U7264 ( .A(n8638), .Z(n9669) );
  CLKBUF_X1 U7296 ( .A(n7477), .Z(n7475) );
  NAND2_X1 U7346 ( .A1(n8876), .A2(n8875), .ZN(n14702) );
  CLKBUF_X1 U7474 ( .A(n8611), .Z(n11616) );
  CLKBUF_X1 U7517 ( .A(n8510), .Z(n6485) );
  INV_X1 U7568 ( .A(n7481), .ZN(n12628) );
  CLKBUF_X1 U8617 ( .A(n14782), .Z(n6480) );
endmodule

