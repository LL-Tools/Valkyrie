

module b17_C_2inp_gates_syn ( P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, 
        DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, 
        DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, 
        DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, 
        DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, 
        DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, 
        READY1, READY2, P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN, 
        P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN, 
        P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN, 
        P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN, 
        P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN, 
        P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN, 
        P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN, 
        P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN, 
        P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN, 
        P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN, 
        P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN, 
        P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN, 
        P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN, 
        P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN, 
        P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN, 
        P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN, 
        P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN, 
        P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, 
        P1_REIP_REG_6__SCAN_IN, P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, 
        P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, 
        P1_REIP_REG_0__SCAN_IN, P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, 
        P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, 
        P1_EBX_REG_26__SCAN_IN, P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, 
        P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, 
        P1_EBX_REG_20__SCAN_IN, P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, 
        P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, 
        P1_EBX_REG_14__SCAN_IN, P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, 
        P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, 
        P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, 
        P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, 
        P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, 
        P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, 
        P1_EAX_REG_28__SCAN_IN, P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, 
        P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, 
        P1_EAX_REG_22__SCAN_IN, P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, 
        P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, 
        P1_EAX_REG_16__SCAN_IN, P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, 
        P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, 
        P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, 
        P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, 
        P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, 
        P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, U355, 
        U356, U357, U358, U359, U360, U361, U362, U363, U364, U366, U367, U368, 
        U369, U370, U371, U372, U373, U374, U375, U347, U348, U349, U350, U351, 
        U352, U353, U354, U365, U376, U247, U246, U245, U244, U243, U242, U241, 
        U240, U239, U238, U237, U236, U235, U234, U233, U232, U231, U230, U229, 
        U228, U227, U226, U225, U224, U223, U222, U221, U220, U219, U218, U217, 
        U216, U251, U252, U253, U254, U255, U256, U257, U258, U259, U260, U261, 
        U262, U263, U264, U265, U266, U267, U268, U269, U270, U271, U272, U273, 
        U274, U275, U276, U277, U278, U279, U280, U281, U282, U212, U215, U213, 
        U214, P3_U3274, P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, 
        P3_U3059, P3_U3058, P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, 
        P3_U3052, P3_U3051, P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, 
        P3_U3045, P3_U3044, P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, 
        P3_U3038, P3_U3037, P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, 
        P3_U3031, P3_U3030, P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, 
        P3_U3026, P3_U3025, P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, 
        P3_U3019, P3_U3018, P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, 
        P3_U3012, P3_U3011, P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, 
        P3_U3005, P3_U3004, P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, 
        P3_U3282, P3_U2998, P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, 
        P3_U2992, P3_U2991, P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, 
        P3_U2985, P3_U2984, P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, 
        P3_U2978, P3_U2977, P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, 
        P3_U2971, P3_U2970, P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, 
        P3_U2964, P3_U2963, P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, 
        P3_U2957, P3_U2956, P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, 
        P3_U2950, P3_U2949, P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, 
        P3_U2943, P3_U2942, P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, 
        P3_U2936, P3_U2935, P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, 
        P3_U2929, P3_U2928, P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, 
        P3_U2922, P3_U2921, P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, 
        P3_U2915, P3_U2914, P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, 
        P3_U2908, P3_U2907, P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, 
        P3_U2901, P3_U2900, P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, 
        P3_U2894, P3_U2893, P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, 
        P3_U2887, P3_U2886, P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, 
        P3_U2880, P3_U2879, P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, 
        P3_U2873, P3_U2872, P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, 
        P3_U3285, P3_U3288, P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, 
        P3_U2864, P3_U2863, P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, 
        P3_U2857, P3_U2856, P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, 
        P3_U2850, P3_U2849, P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, 
        P3_U2843, P3_U2842, P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, 
        P3_U2836, P3_U2835, P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, 
        P3_U2829, P3_U2828, P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, 
        P3_U2822, P3_U2821, P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, 
        P3_U2815, P3_U2814, P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, 
        P3_U2808, P3_U2807, P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, 
        P3_U2801, P3_U2800, P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, 
        P3_U2794, P3_U2793, P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, 
        P3_U2787, P3_U2786, P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, 
        P3_U2780, P3_U2779, P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, 
        P3_U2773, P3_U2772, P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, 
        P3_U2766, P3_U2765, P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, 
        P3_U2759, P3_U2758, P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, 
        P3_U2752, P3_U2751, P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, 
        P3_U2745, P3_U2744, P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, 
        P3_U2738, P3_U2737, P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, 
        P3_U2731, P3_U2730, P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, 
        P3_U2724, P3_U2723, P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, 
        P3_U2717, P3_U2716, P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, 
        P3_U2710, P3_U2709, P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, 
        P3_U2703, P3_U2702, P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, 
        P3_U2696, P3_U2695, P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, 
        P3_U2689, P3_U2688, P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, 
        P3_U2682, P3_U2681, P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, 
        P3_U2675, P3_U2674, P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, 
        P3_U2668, P3_U2667, P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, 
        P3_U2661, P3_U2660, P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, 
        P3_U2654, P3_U2653, P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, 
        P3_U2647, P3_U2646, P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, 
        P3_U2640, P3_U2639, P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, 
        P3_U3295, P3_U2636, P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, 
        P3_U3298, P3_U3299, P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, 
        P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, 
        P2_U3179, P2_U3593, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, 
        P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, 
        P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, 
        P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, 
        P2_U3152, P2_U3151, P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, 
        P2_U3145, P2_U3144, P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, 
        P2_U3138, P2_U3137, P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, 
        P2_U3131, P2_U3130, P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, 
        P2_U3124, P2_U3123, P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, 
        P2_U3117, P2_U3116, P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, 
        P2_U3110, P2_U3109, P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, 
        P2_U3103, P2_U3102, P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, 
        P2_U3096, P2_U3095, P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, 
        P2_U3089, P2_U3088, P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, 
        P2_U3082, P2_U3081, P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, 
        P2_U3075, P2_U3074, P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, 
        P2_U3068, P2_U3067, P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, 
        P2_U3061, P2_U3060, P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, 
        P2_U3054, P2_U3053, P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, 
        P2_U3595, P2_U3596, P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, 
        P2_U3603, P2_U3604, P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, 
        P2_U3042, P2_U3041, P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, 
        P2_U3035, P2_U3034, P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, 
        P2_U3028, P2_U3027, P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, 
        P2_U3021, P2_U3020, P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, 
        P2_U3014, P2_U3013, P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, 
        P2_U3007, P2_U3006, P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, 
        P2_U3000, P2_U2999, P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, 
        P2_U2993, P2_U2992, P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, 
        P2_U2986, P2_U2985, P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, 
        P2_U2979, P2_U2978, P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, 
        P2_U2972, P2_U2971, P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, 
        P2_U2965, P2_U2964, P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, 
        P2_U2958, P2_U2957, P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, 
        P2_U2951, P2_U2950, P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, 
        P2_U2944, P2_U2943, P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, 
        P2_U2937, P2_U2936, P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, 
        P2_U2930, P2_U2929, P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, 
        P2_U2923, P2_U2922, P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, 
        P2_U2916, P2_U2915, P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, 
        P2_U2909, P2_U2908, P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, 
        P2_U2902, P2_U2901, P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, 
        P2_U2895, P2_U2894, P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, 
        P2_U2888, P2_U2887, P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, 
        P2_U2881, P2_U2880, P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, 
        P2_U2874, P2_U2873, P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, 
        P2_U2867, P2_U2866, P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, 
        P2_U2860, P2_U2859, P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, 
        P2_U2853, P2_U2852, P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, 
        P2_U2846, P2_U2845, P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, 
        P2_U2839, P2_U2838, P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, 
        P2_U2832, P2_U2831, P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, 
        P2_U2825, P2_U2824, P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, 
        P2_U2819, P2_U3609, P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, 
        P2_U2815, P2_U3612, P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, 
        P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, 
        P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, 
        P1_U3212, P1_U3211, P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, 
        P1_U3205, P1_U3204, P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, 
        P1_U3198, P1_U3197, P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, 
        P1_U3193, P1_U3192, P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, 
        P1_U3186, P1_U3185, P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, 
        P1_U3179, P1_U3178, P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, 
        P1_U3172, P1_U3171, P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, 
        P1_U3165, P1_U3164, P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, 
        P1_U3159, P1_U3158, P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, 
        P1_U3152, P1_U3151, P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, 
        P1_U3145, P1_U3144, P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, 
        P1_U3138, P1_U3137, P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, 
        P1_U3131, P1_U3130, P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, 
        P1_U3124, P1_U3123, P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, 
        P1_U3117, P1_U3116, P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, 
        P1_U3110, P1_U3109, P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, 
        P1_U3103, P1_U3102, P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, 
        P1_U3096, P1_U3095, P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, 
        P1_U3089, P1_U3088, P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, 
        P1_U3082, P1_U3081, P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, 
        P1_U3075, P1_U3074, P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, 
        P1_U3068, P1_U3067, P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, 
        P1_U3061, P1_U3060, P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, 
        P1_U3054, P1_U3053, P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, 
        P1_U3047, P1_U3046, P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, 
        P1_U3040, P1_U3039, P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, 
        P1_U3033, P1_U3468, P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, 
        P1_U3475, P1_U3476, P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, 
        P1_U3028, P1_U3027, P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, 
        P1_U3021, P1_U3020, P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, 
        P1_U3014, P1_U3013, P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, 
        P1_U3007, P1_U3006, P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, 
        P1_U3000, P1_U2999, P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, 
        P1_U2993, P1_U2992, P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, 
        P1_U2986, P1_U2985, P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, 
        P1_U2979, P1_U2978, P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, 
        P1_U2972, P1_U2971, P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, 
        P1_U2965, P1_U2964, P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, 
        P1_U2958, P1_U2957, P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, 
        P1_U2951, P1_U2950, P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, 
        P1_U2944, P1_U2943, P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, 
        P1_U2937, P1_U2936, P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, 
        P1_U2930, P1_U2929, P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, 
        P1_U2923, P1_U2922, P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, 
        P1_U2916, P1_U2915, P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, 
        P1_U2909, P1_U2908, P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, 
        P1_U2902, P1_U2901, P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, 
        P1_U2895, P1_U2894, P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, 
        P1_U2888, P1_U2887, P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, 
        P1_U2881, P1_U2880, P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, 
        P1_U2874, P1_U2873, P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, 
        P1_U2867, P1_U2866, P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, 
        P1_U2860, P1_U2859, P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, 
        P1_U2853, P1_U2852, P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, 
        P1_U2846, P1_U2845, P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, 
        P1_U2839, P1_U2838, P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, 
        P1_U2832, P1_U2831, P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, 
        P1_U2825, P1_U2824, P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, 
        P1_U2818, P1_U2817, P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, 
        P1_U2811, P1_U2810, P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, 
        P1_U3483, P1_U2806, P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, 
        P1_U2803, P1_U2802, P1_U3487, P1_U2801, keyinput127, keyinput126, 
        keyinput125, keyinput124, keyinput123, keyinput122, keyinput121, 
        keyinput120, keyinput119, keyinput118, keyinput117, keyinput116, 
        keyinput115, keyinput114, keyinput113, keyinput112, keyinput111, 
        keyinput110, keyinput109, keyinput108, keyinput107, keyinput106, 
        keyinput105, keyinput104, keyinput103, keyinput102, keyinput101, 
        keyinput100, keyinput99, keyinput98, keyinput97, keyinput96, 
        keyinput95, keyinput94, keyinput93, keyinput92, keyinput91, keyinput90, 
        keyinput89, keyinput88, keyinput87, keyinput86, keyinput85, keyinput84, 
        keyinput83, keyinput82, keyinput81, keyinput80, keyinput79, keyinput78, 
        keyinput77, keyinput76, keyinput75, keyinput74, keyinput73, keyinput72, 
        keyinput71, keyinput70, keyinput69, keyinput68, keyinput67, keyinput66, 
        keyinput65, keyinput64, keyinput63, keyinput62, keyinput61, keyinput60, 
        keyinput59, keyinput58, keyinput57, keyinput56, keyinput55, keyinput54, 
        keyinput53, keyinput52, keyinput51, keyinput50, keyinput49, keyinput48, 
        keyinput47, keyinput46, keyinput45, keyinput44, keyinput43, keyinput42, 
        keyinput41, keyinput40, keyinput39, keyinput38, keyinput37, keyinput36, 
        keyinput35, keyinput34, keyinput33, keyinput32, keyinput31, keyinput30, 
        keyinput29, keyinput28, keyinput27, keyinput26, keyinput25, keyinput24, 
        keyinput23, keyinput22, keyinput21, keyinput20, keyinput19, keyinput18, 
        keyinput17, keyinput16, keyinput15, keyinput14, keyinput13, keyinput12, 
        keyinput11, keyinput10, keyinput9, keyinput8, keyinput7, keyinput6, 
        keyinput5, keyinput4, keyinput3, keyinput2, keyinput1, keyinput0 );
  input P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_,
         DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_,
         DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_,
         DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_,
         DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_,
         DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2,
         P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN, keyinput127, keyinput126, keyinput125,
         keyinput124, keyinput123, keyinput122, keyinput121, keyinput120,
         keyinput119, keyinput118, keyinput117, keyinput116, keyinput115,
         keyinput114, keyinput113, keyinput112, keyinput111, keyinput110,
         keyinput109, keyinput108, keyinput107, keyinput106, keyinput105,
         keyinput104, keyinput103, keyinput102, keyinput101, keyinput100,
         keyinput99, keyinput98, keyinput97, keyinput96, keyinput95,
         keyinput94, keyinput93, keyinput92, keyinput91, keyinput90,
         keyinput89, keyinput88, keyinput87, keyinput86, keyinput85,
         keyinput84, keyinput83, keyinput82, keyinput81, keyinput80,
         keyinput79, keyinput78, keyinput77, keyinput76, keyinput75,
         keyinput74, keyinput73, keyinput72, keyinput71, keyinput70,
         keyinput69, keyinput68, keyinput67, keyinput66, keyinput65,
         keyinput64, keyinput63, keyinput62, keyinput61, keyinput60,
         keyinput59, keyinput58, keyinput57, keyinput56, keyinput55,
         keyinput54, keyinput53, keyinput52, keyinput51, keyinput50,
         keyinput49, keyinput48, keyinput47, keyinput46, keyinput45,
         keyinput44, keyinput43, keyinput42, keyinput41, keyinput40,
         keyinput39, keyinput38, keyinput37, keyinput36, keyinput35,
         keyinput34, keyinput33, keyinput32, keyinput31, keyinput30,
         keyinput29, keyinput28, keyinput27, keyinput26, keyinput25,
         keyinput24, keyinput23, keyinput22, keyinput21, keyinput20,
         keyinput19, keyinput18, keyinput17, keyinput16, keyinput15,
         keyinput14, keyinput13, keyinput12, keyinput11, keyinput10, keyinput9,
         keyinput8, keyinput7, keyinput6, keyinput5, keyinput4, keyinput3,
         keyinput2, keyinput1, keyinput0;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9747, n9748, n9749, n9750, n9751, n9752, n9753,
         n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763,
         n9764, n9765, n9766, n9769, n9770, n9771, n9772, n9773, n9774, n9775,
         n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785,
         n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795,
         n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805,
         n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815,
         n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825,
         n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835,
         n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845,
         n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855,
         n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865,
         n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875,
         n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885,
         n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895,
         n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905,
         n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915,
         n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925,
         n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935,
         n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945,
         n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955,
         n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965,
         n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975,
         n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985,
         n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995,
         n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004,
         n10005, n10006, n10007, n10008, n10009, n10010, n10011, n10012,
         n10013, n10014, n10015, n10016, n10017, n10018, n10019, n10020,
         n10021, n10022, n10023, n10024, n10025, n10026, n10027, n10028,
         n10029, n10030, n10031, n10032, n10033, n10034, n10035, n10036,
         n10037, n10038, n10039, n10040, n10041, n10042, n10043, n10044,
         n10045, n10046, n10047, n10048, n10049, n10050, n10051, n10052,
         n10053, n10054, n10055, n10056, n10057, n10058, n10059, n10060,
         n10061, n10062, n10063, n10064, n10065, n10066, n10067, n10068,
         n10069, n10070, n10071, n10072, n10073, n10074, n10075, n10076,
         n10077, n10078, n10079, n10080, n10081, n10082, n10083, n10084,
         n10085, n10086, n10087, n10088, n10089, n10090, n10091, n10092,
         n10093, n10094, n10095, n10096, n10097, n10098, n10099, n10100,
         n10101, n10102, n10103, n10104, n10105, n10106, n10107, n10108,
         n10109, n10110, n10111, n10112, n10113, n10114, n10115, n10116,
         n10117, n10118, n10119, n10120, n10121, n10122, n10123, n10124,
         n10125, n10126, n10127, n10128, n10129, n10130, n10131, n10132,
         n10133, n10134, n10135, n10136, n10137, n10138, n10139, n10140,
         n10141, n10142, n10143, n10144, n10145, n10146, n10147, n10148,
         n10149, n10150, n10151, n10152, n10153, n10154, n10155, n10156,
         n10157, n10158, n10159, n10160, n10161, n10162, n10163, n10164,
         n10165, n10166, n10167, n10168, n10169, n10170, n10171, n10172,
         n10173, n10174, n10175, n10176, n10177, n10178, n10179, n10180,
         n10181, n10182, n10183, n10184, n10185, n10186, n10187, n10188,
         n10189, n10190, n10191, n10192, n10193, n10194, n10195, n10196,
         n10197, n10198, n10199, n10200, n10201, n10202, n10203, n10204,
         n10205, n10206, n10207, n10208, n10209, n10210, n10211, n10212,
         n10213, n10214, n10215, n10216, n10217, n10218, n10219, n10220,
         n10221, n10222, n10223, n10224, n10225, n10226, n10227, n10228,
         n10229, n10230, n10231, n10232, n10233, n10234, n10235, n10236,
         n10237, n10238, n10239, n10240, n10241, n10242, n10243, n10244,
         n10245, n10246, n10247, n10248, n10249, n10250, n10251, n10252,
         n10253, n10254, n10255, n10256, n10257, n10258, n10259, n10260,
         n10261, n10262, n10263, n10264, n10265, n10266, n10267, n10268,
         n10269, n10270, n10271, n10272, n10273, n10274, n10275, n10276,
         n10277, n10278, n10279, n10280, n10281, n10282, n10283, n10284,
         n10285, n10286, n10287, n10288, n10289, n10290, n10291, n10292,
         n10293, n10294, n10296, n10297, n10298, n10299, n10300, n10301,
         n10302, n10303, n10304, n10305, n10306, n10307, n10308, n10309,
         n10310, n10311, n10312, n10313, n10314, n10315, n10316, n10317,
         n10318, n10319, n10320, n10321, n10322, n10323, n10324, n10325,
         n10326, n10327, n10328, n10329, n10330, n10331, n10332, n10333,
         n10334, n10335, n10336, n10337, n10338, n10339, n10340, n10341,
         n10342, n10343, n10344, n10345, n10346, n10347, n10348, n10349,
         n10350, n10351, n10352, n10353, n10354, n10355, n10356, n10357,
         n10358, n10359, n10360, n10361, n10362, n10363, n10364, n10365,
         n10366, n10367, n10368, n10369, n10370, n10371, n10372, n10373,
         n10374, n10375, n10376, n10377, n10378, n10379, n10380, n10381,
         n10382, n10383, n10384, n10385, n10386, n10387, n10388, n10389,
         n10390, n10391, n10392, n10393, n10394, n10395, n10396, n10397,
         n10398, n10399, n10400, n10401, n10402, n10403, n10404, n10405,
         n10406, n10407, n10408, n10409, n10410, n10411, n10412, n10413,
         n10414, n10415, n10416, n10417, n10418, n10419, n10420, n10421,
         n10422, n10423, n10424, n10425, n10426, n10427, n10428, n10429,
         n10430, n10431, n10432, n10433, n10434, n10435, n10436, n10437,
         n10438, n10439, n10440, n10441, n10442, n10443, n10444, n10445,
         n10446, n10447, n10448, n10449, n10450, n10451, n10452, n10453,
         n10454, n10455, n10456, n10457, n10458, n10459, n10460, n10461,
         n10462, n10463, n10464, n10465, n10466, n10467, n10468, n10469,
         n10470, n10471, n10472, n10473, n10474, n10475, n10476, n10477,
         n10478, n10479, n10480, n10481, n10482, n10483, n10484, n10485,
         n10486, n10487, n10488, n10489, n10490, n10491, n10492, n10493,
         n10494, n10495, n10496, n10497, n10498, n10499, n10500, n10501,
         n10502, n10503, n10504, n10505, n10506, n10507, n10508, n10509,
         n10510, n10511, n10512, n10513, n10514, n10515, n10516, n10517,
         n10518, n10519, n10520, n10521, n10522, n10523, n10524, n10525,
         n10526, n10527, n10528, n10529, n10530, n10531, n10532, n10533,
         n10534, n10535, n10536, n10537, n10538, n10539, n10540, n10541,
         n10542, n10543, n10544, n10545, n10546, n10547, n10548, n10549,
         n10550, n10551, n10552, n10553, n10554, n10555, n10556, n10557,
         n10558, n10559, n10560, n10561, n10562, n10563, n10564, n10565,
         n10566, n10567, n10568, n10569, n10570, n10571, n10572, n10573,
         n10574, n10575, n10576, n10577, n10578, n10579, n10580, n10581,
         n10582, n10583, n10584, n10585, n10586, n10587, n10588, n10589,
         n10590, n10591, n10592, n10593, n10594, n10595, n10596, n10597,
         n10598, n10599, n10600, n10601, n10602, n10603, n10604, n10605,
         n10606, n10607, n10608, n10609, n10610, n10611, n10612, n10613,
         n10614, n10615, n10616, n10617, n10618, n10619, n10620, n10621,
         n10622, n10623, n10624, n10625, n10626, n10627, n10628, n10629,
         n10630, n10631, n10632, n10633, n10634, n10635, n10636, n10637,
         n10638, n10639, n10640, n10641, n10642, n10643, n10644, n10645,
         n10646, n10647, n10648, n10649, n10650, n10651, n10652, n10653,
         n10654, n10655, n10656, n10657, n10658, n10659, n10660, n10661,
         n10662, n10663, n10664, n10665, n10666, n10667, n10668, n10669,
         n10670, n10671, n10672, n10673, n10674, n10675, n10676, n10677,
         n10678, n10679, n10680, n10681, n10682, n10683, n10684, n10685,
         n10686, n10687, n10688, n10689, n10690, n10691, n10692, n10693,
         n10694, n10695, n10696, n10697, n10698, n10699, n10700, n10701,
         n10702, n10703, n10704, n10705, n10706, n10707, n10708, n10709,
         n10710, n10711, n10712, n10713, n10714, n10715, n10716, n10717,
         n10718, n10719, n10720, n10721, n10722, n10723, n10724, n10725,
         n10726, n10727, n10728, n10729, n10730, n10731, n10732, n10733,
         n10734, n10735, n10736, n10737, n10738, n10739, n10740, n10741,
         n10742, n10743, n10744, n10745, n10746, n10747, n10748, n10749,
         n10750, n10751, n10752, n10753, n10754, n10755, n10756, n10757,
         n10758, n10759, n10760, n10761, n10762, n10763, n10764, n10765,
         n10766, n10767, n10768, n10769, n10770, n10771, n10772, n10773,
         n10774, n10775, n10776, n10777, n10778, n10779, n10780, n10781,
         n10782, n10783, n10784, n10785, n10786, n10787, n10788, n10789,
         n10790, n10791, n10792, n10793, n10794, n10795, n10796, n10797,
         n10798, n10799, n10800, n10801, n10802, n10803, n10804, n10805,
         n10806, n10807, n10808, n10809, n10810, n10811, n10812, n10813,
         n10814, n10815, n10816, n10817, n10818, n10819, n10820, n10821,
         n10822, n10823, n10824, n10825, n10826, n10827, n10828, n10829,
         n10830, n10831, n10832, n10833, n10834, n10835, n10836, n10837,
         n10838, n10839, n10840, n10841, n10842, n10843, n10844, n10845,
         n10846, n10847, n10848, n10849, n10850, n10851, n10852, n10853,
         n10854, n10855, n10856, n10857, n10858, n10859, n10860, n10861,
         n10862, n10863, n10864, n10865, n10866, n10867, n10868, n10869,
         n10870, n10871, n10872, n10873, n10874, n10875, n10876, n10877,
         n10878, n10879, n10880, n10881, n10882, n10883, n10884, n10885,
         n10886, n10887, n10888, n10889, n10890, n10891, n10892, n10893,
         n10894, n10895, n10896, n10897, n10898, n10899, n10900, n10901,
         n10902, n10903, n10904, n10905, n10906, n10907, n10908, n10909,
         n10910, n10911, n10912, n10913, n10914, n10915, n10916, n10917,
         n10918, n10919, n10920, n10921, n10922, n10923, n10924, n10925,
         n10926, n10927, n10928, n10929, n10930, n10931, n10932, n10933,
         n10934, n10935, n10936, n10937, n10938, n10939, n10940, n10941,
         n10942, n10943, n10944, n10945, n10946, n10947, n10948, n10949,
         n10950, n10951, n10952, n10953, n10954, n10955, n10956, n10957,
         n10958, n10959, n10960, n10961, n10962, n10963, n10964, n10965,
         n10966, n10967, n10968, n10969, n10970, n10971, n10972, n10973,
         n10974, n10975, n10976, n10977, n10978, n10979, n10980, n10981,
         n10982, n10983, n10984, n10985, n10986, n10987, n10988, n10989,
         n10990, n10991, n10992, n10993, n10994, n10995, n10996, n10997,
         n10998, n10999, n11000, n11001, n11002, n11003, n11004, n11005,
         n11006, n11007, n11008, n11009, n11010, n11011, n11012, n11013,
         n11014, n11015, n11016, n11017, n11018, n11019, n11020, n11021,
         n11022, n11023, n11024, n11025, n11026, n11027, n11028, n11029,
         n11030, n11031, n11032, n11033, n11034, n11035, n11036, n11037,
         n11038, n11039, n11040, n11041, n11042, n11043, n11044, n11045,
         n11046, n11047, n11048, n11049, n11050, n11051, n11052, n11053,
         n11054, n11055, n11056, n11057, n11058, n11059, n11060, n11061,
         n11062, n11063, n11064, n11065, n11066, n11067, n11068, n11069,
         n11070, n11071, n11072, n11073, n11074, n11075, n11076, n11077,
         n11078, n11079, n11080, n11081, n11082, n11083, n11084, n11085,
         n11086, n11087, n11088, n11089, n11090, n11091, n11092, n11093,
         n11094, n11095, n11096, n11097, n11098, n11099, n11100, n11101,
         n11102, n11103, n11104, n11105, n11106, n11107, n11108, n11109,
         n11110, n11111, n11112, n11113, n11114, n11115, n11116, n11117,
         n11118, n11119, n11120, n11121, n11122, n11123, n11124, n11125,
         n11126, n11127, n11128, n11129, n11130, n11131, n11132, n11133,
         n11134, n11135, n11136, n11137, n11138, n11139, n11140, n11141,
         n11142, n11143, n11144, n11145, n11146, n11147, n11148, n11149,
         n11150, n11151, n11152, n11153, n11154, n11155, n11156, n11157,
         n11158, n11159, n11160, n11161, n11162, n11163, n11164, n11165,
         n11166, n11167, n11168, n11169, n11170, n11171, n11172, n11173,
         n11174, n11175, n11176, n11177, n11178, n11179, n11180, n11181,
         n11182, n11183, n11184, n11185, n11186, n11187, n11188, n11189,
         n11190, n11191, n11192, n11193, n11194, n11195, n11196, n11197,
         n11198, n11199, n11200, n11201, n11202, n11203, n11204, n11205,
         n11206, n11207, n11208, n11209, n11210, n11211, n11212, n11213,
         n11214, n11215, n11216, n11217, n11218, n11219, n11220, n11221,
         n11222, n11223, n11224, n11225, n11226, n11227, n11228, n11229,
         n11230, n11231, n11232, n11233, n11234, n11235, n11236, n11237,
         n11238, n11239, n11240, n11241, n11242, n11243, n11244, n11245,
         n11246, n11247, n11248, n11249, n11250, n11251, n11252, n11253,
         n11254, n11255, n11256, n11257, n11258, n11259, n11260, n11261,
         n11262, n11263, n11264, n11265, n11266, n11267, n11268, n11269,
         n11270, n11271, n11272, n11273, n11274, n11275, n11276, n11277,
         n11278, n11279, n11280, n11281, n11282, n11283, n11284, n11285,
         n11286, n11287, n11288, n11289, n11290, n11291, n11292, n11293,
         n11294, n11295, n11296, n11297, n11298, n11299, n11300, n11301,
         n11302, n11303, n11304, n11305, n11306, n11307, n11308, n11309,
         n11310, n11311, n11312, n11313, n11314, n11315, n11316, n11317,
         n11318, n11319, n11320, n11321, n11322, n11323, n11324, n11325,
         n11326, n11327, n11328, n11329, n11330, n11331, n11332, n11333,
         n11334, n11335, n11336, n11337, n11338, n11339, n11340, n11341,
         n11342, n11343, n11344, n11345, n11346, n11347, n11348, n11349,
         n11350, n11351, n11352, n11353, n11354, n11355, n11356, n11357,
         n11358, n11359, n11360, n11361, n11362, n11363, n11364, n11365,
         n11366, n11367, n11368, n11369, n11370, n11371, n11372, n11373,
         n11374, n11375, n11376, n11377, n11378, n11379, n11380, n11381,
         n11382, n11383, n11384, n11385, n11386, n11387, n11388, n11389,
         n11390, n11391, n11392, n11393, n11394, n11395, n11396, n11397,
         n11398, n11399, n11400, n11401, n11402, n11403, n11404, n11405,
         n11406, n11407, n11408, n11409, n11410, n11411, n11412, n11413,
         n11414, n11415, n11416, n11417, n11418, n11419, n11420, n11421,
         n11422, n11423, n11424, n11425, n11426, n11427, n11428, n11429,
         n11430, n11431, n11432, n11433, n11434, n11435, n11436, n11437,
         n11438, n11439, n11440, n11441, n11442, n11443, n11444, n11445,
         n11446, n11447, n11448, n11449, n11450, n11451, n11452, n11453,
         n11454, n11455, n11456, n11457, n11458, n11459, n11460, n11461,
         n11462, n11463, n11464, n11465, n11466, n11467, n11468, n11469,
         n11470, n11471, n11472, n11473, n11474, n11475, n11476, n11477,
         n11478, n11479, n11480, n11481, n11482, n11483, n11484, n11485,
         n11486, n11487, n11488, n11489, n11490, n11491, n11492, n11493,
         n11494, n11495, n11496, n11497, n11498, n11499, n11500, n11501,
         n11502, n11503, n11504, n11505, n11506, n11507, n11508, n11509,
         n11510, n11511, n11512, n11513, n11514, n11515, n11516, n11517,
         n11518, n11519, n11520, n11521, n11522, n11523, n11524, n11525,
         n11526, n11527, n11528, n11529, n11530, n11531, n11532, n11533,
         n11534, n11535, n11536, n11537, n11538, n11539, n11540, n11541,
         n11542, n11543, n11544, n11545, n11546, n11547, n11548, n11549,
         n11550, n11551, n11552, n11553, n11554, n11555, n11556, n11557,
         n11558, n11559, n11560, n11561, n11562, n11563, n11564, n11565,
         n11566, n11567, n11568, n11569, n11570, n11571, n11572, n11573,
         n11574, n11575, n11576, n11577, n11578, n11579, n11580, n11581,
         n11582, n11583, n11584, n11585, n11586, n11587, n11588, n11589,
         n11590, n11591, n11592, n11593, n11594, n11595, n11596, n11597,
         n11598, n11599, n11600, n11601, n11602, n11603, n11604, n11605,
         n11606, n11607, n11608, n11609, n11610, n11611, n11612, n11613,
         n11614, n11615, n11616, n11617, n11618, n11619, n11620, n11621,
         n11622, n11623, n11624, n11625, n11626, n11627, n11628, n11629,
         n11630, n11631, n11632, n11633, n11634, n11635, n11636, n11637,
         n11638, n11639, n11640, n11641, n11642, n11643, n11644, n11645,
         n11646, n11647, n11648, n11649, n11650, n11651, n11652, n11653,
         n11654, n11655, n11656, n11657, n11658, n11659, n11660, n11661,
         n11662, n11663, n11664, n11665, n11666, n11667, n11668, n11669,
         n11670, n11671, n11672, n11673, n11674, n11675, n11676, n11677,
         n11678, n11679, n11680, n11681, n11682, n11683, n11684, n11685,
         n11686, n11687, n11688, n11689, n11690, n11691, n11692, n11693,
         n11694, n11695, n11696, n11697, n11698, n11699, n11700, n11701,
         n11702, n11703, n11704, n11705, n11706, n11707, n11708, n11709,
         n11710, n11711, n11712, n11713, n11714, n11715, n11716, n11717,
         n11718, n11719, n11720, n11721, n11722, n11723, n11724, n11725,
         n11726, n11727, n11728, n11729, n11730, n11731, n11732, n11733,
         n11734, n11735, n11736, n11737, n11738, n11739, n11740, n11741,
         n11742, n11743, n11744, n11745, n11746, n11747, n11748, n11749,
         n11750, n11751, n11752, n11753, n11754, n11755, n11756, n11757,
         n11758, n11759, n11760, n11761, n11762, n11763, n11764, n11765,
         n11766, n11767, n11768, n11769, n11770, n11771, n11772, n11773,
         n11774, n11775, n11776, n11777, n11778, n11779, n11780, n11781,
         n11782, n11783, n11784, n11785, n11786, n11787, n11788, n11789,
         n11790, n11791, n11792, n11793, n11794, n11795, n11796, n11797,
         n11798, n11799, n11800, n11801, n11802, n11803, n11804, n11805,
         n11806, n11807, n11808, n11809, n11810, n11811, n11812, n11813,
         n11814, n11815, n11816, n11817, n11818, n11819, n11820, n11821,
         n11822, n11823, n11824, n11825, n11826, n11827, n11828, n11829,
         n11830, n11831, n11832, n11833, n11834, n11835, n11836, n11837,
         n11838, n11839, n11840, n11841, n11842, n11843, n11844, n11845,
         n11846, n11847, n11848, n11849, n11850, n11851, n11852, n11853,
         n11854, n11855, n11856, n11857, n11858, n11859, n11860, n11861,
         n11862, n11863, n11864, n11865, n11866, n11867, n11868, n11869,
         n11870, n11871, n11872, n11873, n11874, n11875, n11876, n11877,
         n11878, n11879, n11880, n11881, n11882, n11883, n11884, n11885,
         n11886, n11887, n11888, n11889, n11890, n11891, n11892, n11893,
         n11894, n11895, n11896, n11897, n11898, n11899, n11900, n11901,
         n11902, n11903, n11904, n11905, n11906, n11907, n11908, n11909,
         n11910, n11911, n11912, n11913, n11914, n11915, n11916, n11917,
         n11918, n11919, n11920, n11921, n11922, n11923, n11924, n11925,
         n11926, n11927, n11928, n11929, n11930, n11931, n11932, n11933,
         n11934, n11935, n11936, n11937, n11938, n11939, n11940, n11941,
         n11942, n11943, n11944, n11945, n11946, n11947, n11948, n11949,
         n11950, n11951, n11952, n11953, n11954, n11955, n11956, n11957,
         n11958, n11959, n11960, n11961, n11962, n11963, n11964, n11965,
         n11966, n11967, n11968, n11969, n11970, n11971, n11972, n11973,
         n11974, n11975, n11976, n11977, n11978, n11979, n11980, n11981,
         n11982, n11983, n11984, n11985, n11986, n11987, n11988, n11989,
         n11990, n11991, n11992, n11993, n11994, n11995, n11996, n11997,
         n11998, n11999, n12000, n12001, n12002, n12003, n12004, n12005,
         n12006, n12007, n12008, n12009, n12010, n12011, n12012, n12013,
         n12014, n12015, n12016, n12017, n12018, n12019, n12020, n12021,
         n12022, n12023, n12024, n12025, n12026, n12027, n12028, n12029,
         n12030, n12031, n12032, n12033, n12034, n12035, n12036, n12037,
         n12038, n12039, n12040, n12041, n12042, n12043, n12044, n12045,
         n12046, n12047, n12048, n12049, n12050, n12051, n12052, n12053,
         n12054, n12055, n12056, n12057, n12058, n12059, n12060, n12061,
         n12062, n12063, n12064, n12065, n12066, n12067, n12068, n12069,
         n12070, n12071, n12072, n12073, n12074, n12075, n12076, n12077,
         n12078, n12079, n12080, n12081, n12082, n12083, n12084, n12085,
         n12086, n12087, n12088, n12089, n12090, n12091, n12092, n12093,
         n12094, n12095, n12096, n12097, n12098, n12099, n12100, n12101,
         n12102, n12103, n12104, n12105, n12106, n12107, n12108, n12109,
         n12110, n12111, n12112, n12113, n12114, n12115, n12116, n12117,
         n12118, n12119, n12120, n12121, n12122, n12123, n12124, n12125,
         n12126, n12127, n12128, n12129, n12130, n12131, n12132, n12133,
         n12134, n12135, n12136, n12137, n12138, n12139, n12140, n12141,
         n12142, n12143, n12144, n12145, n12146, n12147, n12148, n12149,
         n12150, n12151, n12152, n12153, n12154, n12155, n12156, n12157,
         n12158, n12159, n12160, n12161, n12162, n12163, n12164, n12165,
         n12166, n12167, n12168, n12169, n12170, n12171, n12172, n12173,
         n12174, n12175, n12176, n12177, n12178, n12179, n12180, n12181,
         n12182, n12183, n12184, n12185, n12186, n12187, n12188, n12189,
         n12190, n12191, n12192, n12193, n12194, n12195, n12196, n12197,
         n12198, n12199, n12200, n12201, n12202, n12203, n12204, n12205,
         n12206, n12207, n12208, n12209, n12210, n12211, n12212, n12213,
         n12214, n12215, n12216, n12217, n12218, n12219, n12220, n12221,
         n12222, n12223, n12224, n12225, n12226, n12227, n12228, n12229,
         n12230, n12231, n12232, n12233, n12234, n12235, n12236, n12237,
         n12238, n12239, n12240, n12241, n12242, n12243, n12244, n12245,
         n12246, n12247, n12248, n12249, n12250, n12251, n12252, n12253,
         n12254, n12255, n12256, n12257, n12258, n12259, n12260, n12261,
         n12262, n12263, n12264, n12265, n12266, n12267, n12268, n12269,
         n12270, n12271, n12272, n12273, n12274, n12275, n12276, n12277,
         n12278, n12279, n12280, n12281, n12282, n12283, n12284, n12285,
         n12286, n12287, n12288, n12289, n12290, n12291, n12292, n12293,
         n12294, n12295, n12296, n12297, n12298, n12299, n12300, n12301,
         n12302, n12303, n12304, n12305, n12306, n12307, n12308, n12309,
         n12310, n12311, n12312, n12313, n12314, n12315, n12316, n12317,
         n12318, n12319, n12320, n12321, n12322, n12323, n12324, n12325,
         n12326, n12327, n12328, n12329, n12330, n12331, n12332, n12333,
         n12334, n12335, n12336, n12337, n12338, n12339, n12340, n12341,
         n12342, n12343, n12344, n12345, n12346, n12347, n12348, n12349,
         n12350, n12351, n12352, n12353, n12354, n12355, n12356, n12357,
         n12358, n12359, n12360, n12361, n12362, n12363, n12364, n12365,
         n12366, n12367, n12368, n12369, n12370, n12371, n12372, n12373,
         n12374, n12375, n12376, n12377, n12378, n12379, n12380, n12381,
         n12382, n12383, n12384, n12385, n12386, n12387, n12388, n12389,
         n12390, n12391, n12392, n12393, n12394, n12395, n12396, n12397,
         n12398, n12399, n12400, n12401, n12402, n12403, n12404, n12405,
         n12406, n12407, n12408, n12409, n12410, n12411, n12412, n12413,
         n12414, n12415, n12416, n12417, n12418, n12419, n12420, n12421,
         n12422, n12423, n12424, n12425, n12426, n12427, n12428, n12429,
         n12430, n12431, n12432, n12433, n12434, n12435, n12436, n12437,
         n12438, n12439, n12440, n12441, n12442, n12443, n12444, n12445,
         n12446, n12447, n12448, n12449, n12450, n12451, n12452, n12453,
         n12454, n12455, n12456, n12457, n12458, n12459, n12460, n12461,
         n12462, n12463, n12464, n12465, n12466, n12467, n12468, n12469,
         n12470, n12471, n12472, n12473, n12474, n12475, n12476, n12477,
         n12478, n12479, n12480, n12481, n12482, n12483, n12484, n12485,
         n12486, n12487, n12488, n12489, n12490, n12491, n12492, n12493,
         n12494, n12495, n12496, n12497, n12498, n12499, n12500, n12501,
         n12502, n12503, n12504, n12505, n12506, n12507, n12508, n12509,
         n12510, n12511, n12512, n12513, n12514, n12515, n12516, n12517,
         n12518, n12519, n12520, n12521, n12522, n12523, n12524, n12525,
         n12526, n12527, n12528, n12529, n12530, n12531, n12532, n12533,
         n12534, n12535, n12536, n12537, n12538, n12539, n12540, n12541,
         n12542, n12543, n12544, n12545, n12546, n12547, n12548, n12549,
         n12550, n12551, n12552, n12553, n12554, n12555, n12556, n12557,
         n12558, n12559, n12561, n12562, n12563, n12564, n12565, n12566,
         n12567, n12568, n12569, n12570, n12571, n12572, n12573, n12574,
         n12575, n12576, n12577, n12578, n12579, n12580, n12581, n12582,
         n12583, n12584, n12585, n12586, n12587, n12588, n12589, n12590,
         n12591, n12592, n12593, n12594, n12595, n12596, n12597, n12598,
         n12599, n12600, n12601, n12602, n12603, n12604, n12605, n12606,
         n12607, n12608, n12609, n12610, n12611, n12612, n12613, n12614,
         n12615, n12616, n12617, n12618, n12619, n12620, n12621, n12622,
         n12623, n12624, n12625, n12626, n12627, n12628, n12629, n12630,
         n12631, n12632, n12633, n12634, n12635, n12636, n12637, n12638,
         n12639, n12640, n12641, n12642, n12643, n12644, n12645, n12646,
         n12647, n12648, n12649, n12650, n12651, n12652, n12653, n12654,
         n12655, n12656, n12657, n12658, n12659, n12660, n12661, n12662,
         n12663, n12664, n12665, n12666, n12667, n12668, n12669, n12670,
         n12671, n12672, n12673, n12674, n12675, n12676, n12677, n12678,
         n12679, n12680, n12681, n12682, n12683, n12684, n12685, n12686,
         n12687, n12688, n12689, n12690, n12691, n12692, n12693, n12694,
         n12695, n12696, n12697, n12698, n12699, n12700, n12701, n12702,
         n12703, n12704, n12705, n12706, n12707, n12708, n12709, n12710,
         n12711, n12712, n12713, n12714, n12715, n12716, n12717, n12718,
         n12719, n12720, n12721, n12722, n12723, n12724, n12725, n12726,
         n12727, n12728, n12729, n12730, n12731, n12732, n12733, n12734,
         n12735, n12736, n12737, n12738, n12739, n12740, n12741, n12742,
         n12743, n12744, n12745, n12746, n12747, n12748, n12749, n12750,
         n12751, n12752, n12753, n12754, n12755, n12756, n12757, n12758,
         n12759, n12760, n12761, n12762, n12763, n12764, n12765, n12766,
         n12767, n12768, n12769, n12770, n12771, n12772, n12773, n12774,
         n12775, n12776, n12777, n12778, n12779, n12780, n12781, n12782,
         n12783, n12784, n12785, n12786, n12787, n12788, n12789, n12790,
         n12791, n12792, n12793, n12794, n12795, n12796, n12797, n12798,
         n12799, n12800, n12801, n12802, n12803, n12804, n12805, n12806,
         n12807, n12808, n12809, n12810, n12811, n12812, n12813, n12814,
         n12815, n12816, n12817, n12818, n12819, n12820, n12821, n12822,
         n12823, n12824, n12825, n12826, n12827, n12828, n12829, n12830,
         n12831, n12832, n12833, n12834, n12835, n12836, n12837, n12838,
         n12839, n12840, n12841, n12842, n12843, n12844, n12845, n12846,
         n12847, n12848, n12849, n12850, n12851, n12852, n12853, n12854,
         n12855, n12856, n12857, n12858, n12859, n12860, n12861, n12862,
         n12863, n12864, n12865, n12866, n12867, n12868, n12869, n12870,
         n12871, n12872, n12873, n12874, n12875, n12876, n12877, n12878,
         n12879, n12880, n12881, n12882, n12883, n12884, n12885, n12886,
         n12887, n12888, n12889, n12890, n12891, n12892, n12893, n12894,
         n12895, n12896, n12897, n12898, n12899, n12900, n12901, n12902,
         n12903, n12904, n12905, n12906, n12907, n12908, n12909, n12910,
         n12911, n12912, n12913, n12914, n12915, n12916, n12917, n12918,
         n12919, n12920, n12921, n12922, n12923, n12924, n12925, n12926,
         n12927, n12928, n12929, n12930, n12931, n12932, n12933, n12934,
         n12935, n12936, n12937, n12938, n12939, n12940, n12941, n12942,
         n12943, n12944, n12945, n12946, n12947, n12948, n12949, n12950,
         n12951, n12952, n12953, n12954, n12955, n12956, n12957, n12958,
         n12959, n12960, n12961, n12962, n12963, n12964, n12965, n12966,
         n12967, n12968, n12969, n12970, n12971, n12972, n12973, n12974,
         n12975, n12976, n12977, n12978, n12979, n12980, n12981, n12982,
         n12983, n12984, n12985, n12986, n12987, n12988, n12989, n12990,
         n12991, n12992, n12993, n12994, n12995, n12996, n12997, n12998,
         n12999, n13000, n13001, n13002, n13003, n13004, n13005, n13006,
         n13007, n13008, n13009, n13010, n13011, n13012, n13013, n13014,
         n13015, n13016, n13017, n13018, n13019, n13020, n13021, n13022,
         n13023, n13024, n13025, n13026, n13027, n13028, n13029, n13030,
         n13031, n13032, n13033, n13034, n13035, n13036, n13037, n13038,
         n13039, n13040, n13041, n13042, n13043, n13044, n13045, n13046,
         n13047, n13048, n13049, n13050, n13051, n13052, n13053, n13054,
         n13055, n13056, n13057, n13058, n13059, n13060, n13061, n13062,
         n13063, n13064, n13065, n13066, n13067, n13068, n13069, n13070,
         n13071, n13072, n13073, n13074, n13075, n13076, n13077, n13078,
         n13079, n13080, n13081, n13082, n13083, n13084, n13085, n13086,
         n13087, n13088, n13089, n13090, n13091, n13092, n13093, n13094,
         n13095, n13096, n13097, n13098, n13099, n13100, n13101, n13102,
         n13103, n13104, n13105, n13106, n13107, n13108, n13109, n13110,
         n13111, n13112, n13113, n13114, n13115, n13116, n13117, n13118,
         n13119, n13120, n13121, n13122, n13123, n13124, n13125, n13126,
         n13127, n13128, n13129, n13130, n13131, n13132, n13133, n13134,
         n13135, n13136, n13137, n13138, n13139, n13140, n13141, n13142,
         n13143, n13144, n13145, n13146, n13147, n13148, n13149, n13150,
         n13151, n13152, n13153, n13154, n13155, n13156, n13157, n13158,
         n13159, n13160, n13161, n13162, n13163, n13164, n13165, n13166,
         n13167, n13168, n13169, n13170, n13171, n13172, n13173, n13174,
         n13175, n13176, n13177, n13178, n13179, n13180, n13181, n13182,
         n13183, n13184, n13185, n13186, n13187, n13188, n13189, n13190,
         n13191, n13192, n13193, n13194, n13195, n13196, n13197, n13198,
         n13199, n13200, n13201, n13202, n13203, n13204, n13205, n13206,
         n13207, n13208, n13209, n13210, n13211, n13212, n13213, n13214,
         n13215, n13216, n13217, n13218, n13219, n13220, n13221, n13222,
         n13223, n13224, n13225, n13226, n13227, n13228, n13229, n13230,
         n13231, n13232, n13233, n13234, n13235, n13236, n13237, n13238,
         n13239, n13240, n13241, n13242, n13243, n13244, n13245, n13246,
         n13247, n13248, n13249, n13250, n13251, n13252, n13253, n13254,
         n13255, n13256, n13257, n13258, n13259, n13260, n13261, n13262,
         n13263, n13264, n13265, n13266, n13267, n13268, n13269, n13270,
         n13271, n13272, n13273, n13274, n13275, n13276, n13277, n13278,
         n13279, n13280, n13281, n13282, n13283, n13284, n13285, n13286,
         n13287, n13288, n13289, n13290, n13291, n13292, n13293, n13294,
         n13295, n13296, n13297, n13298, n13299, n13300, n13301, n13302,
         n13303, n13304, n13305, n13306, n13307, n13308, n13309, n13310,
         n13311, n13312, n13313, n13314, n13315, n13316, n13317, n13318,
         n13319, n13320, n13321, n13322, n13323, n13324, n13325, n13326,
         n13327, n13328, n13329, n13330, n13331, n13332, n13333, n13334,
         n13335, n13336, n13337, n13338, n13339, n13340, n13341, n13342,
         n13343, n13344, n13345, n13346, n13347, n13348, n13349, n13350,
         n13351, n13352, n13353, n13354, n13355, n13356, n13357, n13358,
         n13359, n13360, n13361, n13362, n13363, n13364, n13365, n13366,
         n13367, n13368, n13369, n13370, n13371, n13372, n13373, n13374,
         n13375, n13376, n13377, n13378, n13379, n13380, n13381, n13382,
         n13383, n13384, n13385, n13386, n13387, n13388, n13389, n13390,
         n13391, n13392, n13393, n13394, n13395, n13396, n13397, n13398,
         n13399, n13400, n13401, n13402, n13403, n13404, n13405, n13406,
         n13407, n13408, n13409, n13410, n13411, n13412, n13413, n13414,
         n13415, n13416, n13417, n13418, n13419, n13420, n13421, n13422,
         n13423, n13424, n13425, n13426, n13427, n13428, n13429, n13430,
         n13431, n13432, n13433, n13434, n13435, n13436, n13437, n13438,
         n13439, n13440, n13441, n13442, n13443, n13444, n13445, n13446,
         n13447, n13448, n13449, n13450, n13451, n13452, n13453, n13454,
         n13455, n13456, n13457, n13458, n13459, n13460, n13461, n13462,
         n13463, n13464, n13465, n13466, n13467, n13468, n13469, n13470,
         n13471, n13472, n13473, n13474, n13475, n13476, n13477, n13478,
         n13479, n13480, n13481, n13482, n13483, n13484, n13485, n13486,
         n13487, n13488, n13489, n13490, n13491, n13492, n13493, n13494,
         n13495, n13496, n13497, n13498, n13499, n13500, n13501, n13502,
         n13503, n13504, n13505, n13506, n13507, n13508, n13509, n13510,
         n13511, n13512, n13513, n13514, n13515, n13516, n13517, n13518,
         n13519, n13520, n13521, n13522, n13523, n13524, n13525, n13526,
         n13527, n13528, n13529, n13530, n13531, n13532, n13533, n13534,
         n13535, n13536, n13537, n13538, n13539, n13540, n13541, n13542,
         n13543, n13544, n13545, n13546, n13547, n13548, n13549, n13550,
         n13551, n13552, n13553, n13554, n13555, n13556, n13557, n13558,
         n13559, n13560, n13561, n13562, n13563, n13564, n13565, n13566,
         n13567, n13568, n13569, n13570, n13571, n13572, n13573, n13574,
         n13575, n13576, n13577, n13578, n13579, n13580, n13581, n13582,
         n13583, n13584, n13585, n13586, n13587, n13588, n13589, n13590,
         n13591, n13592, n13593, n13594, n13595, n13596, n13597, n13598,
         n13599, n13600, n13601, n13602, n13603, n13604, n13605, n13606,
         n13607, n13608, n13609, n13610, n13611, n13612, n13613, n13614,
         n13615, n13616, n13617, n13618, n13619, n13620, n13621, n13622,
         n13623, n13624, n13625, n13626, n13627, n13628, n13629, n13630,
         n13631, n13632, n13633, n13634, n13635, n13636, n13637, n13638,
         n13639, n13640, n13641, n13642, n13643, n13644, n13645, n13646,
         n13647, n13648, n13649, n13650, n13651, n13652, n13653, n13654,
         n13655, n13656, n13657, n13658, n13659, n13660, n13661, n13662,
         n13663, n13664, n13665, n13666, n13667, n13668, n13669, n13670,
         n13671, n13672, n13673, n13674, n13675, n13676, n13677, n13678,
         n13679, n13680, n13681, n13682, n13683, n13684, n13685, n13686,
         n13687, n13688, n13689, n13690, n13691, n13692, n13693, n13694,
         n13695, n13696, n13697, n13698, n13699, n13700, n13701, n13702,
         n13703, n13704, n13705, n13706, n13707, n13708, n13709, n13710,
         n13711, n13712, n13713, n13714, n13715, n13716, n13717, n13718,
         n13719, n13720, n13721, n13722, n13723, n13724, n13725, n13726,
         n13727, n13728, n13729, n13730, n13731, n13732, n13733, n13734,
         n13735, n13736, n13737, n13738, n13739, n13740, n13741, n13742,
         n13743, n13744, n13745, n13746, n13747, n13748, n13749, n13750,
         n13751, n13752, n13753, n13754, n13755, n13756, n13757, n13758,
         n13759, n13760, n13761, n13762, n13763, n13764, n13765, n13766,
         n13767, n13768, n13769, n13770, n13771, n13772, n13773, n13774,
         n13775, n13776, n13777, n13778, n13779, n13780, n13781, n13782,
         n13783, n13784, n13785, n13786, n13787, n13788, n13789, n13790,
         n13791, n13792, n13793, n13794, n13795, n13796, n13797, n13798,
         n13799, n13800, n13801, n13802, n13803, n13804, n13805, n13806,
         n13807, n13808, n13809, n13810, n13811, n13812, n13813, n13814,
         n13815, n13816, n13817, n13818, n13819, n13820, n13821, n13822,
         n13823, n13824, n13825, n13826, n13827, n13828, n13829, n13830,
         n13831, n13832, n13833, n13834, n13835, n13836, n13837, n13838,
         n13839, n13840, n13841, n13842, n13843, n13844, n13845, n13846,
         n13847, n13848, n13849, n13850, n13851, n13852, n13853, n13854,
         n13855, n13856, n13857, n13858, n13859, n13860, n13861, n13862,
         n13863, n13864, n13865, n13866, n13867, n13868, n13869, n13870,
         n13871, n13872, n13873, n13874, n13875, n13876, n13877, n13878,
         n13879, n13880, n13881, n13882, n13883, n13884, n13885, n13886,
         n13887, n13888, n13889, n13890, n13891, n13892, n13893, n13894,
         n13895, n13896, n13897, n13898, n13899, n13900, n13901, n13902,
         n13903, n13904, n13905, n13906, n13907, n13908, n13909, n13910,
         n13911, n13912, n13913, n13914, n13915, n13916, n13917, n13918,
         n13919, n13920, n13921, n13922, n13923, n13924, n13925, n13926,
         n13927, n13928, n13929, n13930, n13931, n13932, n13933, n13934,
         n13935, n13936, n13937, n13938, n13939, n13940, n13941, n13942,
         n13943, n13944, n13945, n13946, n13947, n13948, n13949, n13950,
         n13951, n13952, n13953, n13954, n13955, n13956, n13957, n13958,
         n13959, n13960, n13961, n13962, n13963, n13964, n13965, n13966,
         n13967, n13968, n13969, n13970, n13971, n13972, n13973, n13974,
         n13975, n13976, n13977, n13978, n13979, n13980, n13981, n13982,
         n13983, n13984, n13985, n13986, n13987, n13988, n13989, n13990,
         n13991, n13992, n13993, n13994, n13995, n13996, n13997, n13998,
         n13999, n14000, n14001, n14002, n14003, n14004, n14005, n14006,
         n14007, n14008, n14009, n14010, n14011, n14012, n14013, n14014,
         n14015, n14016, n14017, n14018, n14019, n14020, n14021, n14022,
         n14023, n14024, n14025, n14026, n14027, n14028, n14029, n14030,
         n14031, n14032, n14033, n14034, n14035, n14036, n14037, n14038,
         n14039, n14040, n14041, n14042, n14043, n14044, n14045, n14046,
         n14047, n14048, n14049, n14050, n14051, n14052, n14053, n14054,
         n14055, n14056, n14057, n14058, n14059, n14060, n14061, n14062,
         n14063, n14064, n14065, n14066, n14067, n14068, n14069, n14070,
         n14071, n14072, n14073, n14074, n14075, n14076, n14077, n14078,
         n14079, n14080, n14081, n14082, n14083, n14084, n14085, n14086,
         n14087, n14088, n14089, n14090, n14091, n14092, n14093, n14094,
         n14095, n14096, n14097, n14098, n14099, n14100, n14101, n14102,
         n14103, n14104, n14105, n14106, n14107, n14108, n14109, n14110,
         n14111, n14112, n14113, n14114, n14115, n14116, n14117, n14118,
         n14119, n14120, n14121, n14122, n14123, n14124, n14125, n14126,
         n14127, n14128, n14129, n14130, n14131, n14132, n14133, n14134,
         n14135, n14136, n14137, n14138, n14139, n14140, n14141, n14142,
         n14143, n14144, n14145, n14146, n14147, n14148, n14149, n14150,
         n14151, n14152, n14153, n14154, n14155, n14156, n14157, n14158,
         n14159, n14160, n14161, n14162, n14163, n14164, n14165, n14166,
         n14167, n14168, n14169, n14170, n14171, n14172, n14173, n14174,
         n14175, n14176, n14177, n14178, n14179, n14180, n14181, n14182,
         n14183, n14184, n14185, n14186, n14187, n14188, n14189, n14190,
         n14191, n14192, n14193, n14194, n14195, n14196, n14197, n14198,
         n14199, n14200, n14201, n14202, n14203, n14204, n14205, n14206,
         n14207, n14208, n14209, n14210, n14211, n14212, n14213, n14214,
         n14215, n14216, n14217, n14218, n14219, n14220, n14221, n14222,
         n14223, n14224, n14225, n14226, n14227, n14228, n14229, n14230,
         n14231, n14232, n14233, n14234, n14235, n14236, n14237, n14238,
         n14239, n14240, n14241, n14242, n14243, n14244, n14245, n14246,
         n14247, n14248, n14249, n14250, n14251, n14252, n14253, n14254,
         n14255, n14256, n14257, n14258, n14259, n14260, n14261, n14262,
         n14263, n14264, n14265, n14266, n14267, n14268, n14269, n14270,
         n14271, n14272, n14273, n14274, n14275, n14276, n14277, n14278,
         n14279, n14280, n14281, n14282, n14283, n14284, n14285, n14286,
         n14287, n14288, n14289, n14290, n14291, n14292, n14293, n14294,
         n14295, n14296, n14297, n14298, n14299, n14300, n14301, n14302,
         n14303, n14304, n14305, n14306, n14307, n14308, n14309, n14310,
         n14311, n14312, n14313, n14314, n14315, n14316, n14317, n14318,
         n14319, n14320, n14321, n14322, n14323, n14324, n14325, n14326,
         n14327, n14328, n14329, n14330, n14331, n14332, n14333, n14334,
         n14335, n14336, n14337, n14338, n14339, n14340, n14341, n14342,
         n14343, n14344, n14345, n14346, n14347, n14348, n14349, n14350,
         n14351, n14352, n14353, n14354, n14355, n14356, n14357, n14358,
         n14359, n14360, n14361, n14362, n14363, n14364, n14365, n14366,
         n14367, n14368, n14369, n14370, n14371, n14372, n14373, n14374,
         n14375, n14376, n14377, n14378, n14379, n14380, n14381, n14382,
         n14383, n14384, n14385, n14386, n14387, n14388, n14389, n14390,
         n14391, n14392, n14393, n14394, n14395, n14396, n14397, n14398,
         n14399, n14400, n14401, n14402, n14403, n14404, n14405, n14406,
         n14407, n14408, n14409, n14410, n14411, n14412, n14413, n14414,
         n14415, n14416, n14417, n14418, n14419, n14420, n14421, n14422,
         n14423, n14424, n14425, n14426, n14427, n14428, n14429, n14430,
         n14431, n14432, n14433, n14434, n14435, n14436, n14437, n14438,
         n14439, n14440, n14441, n14442, n14443, n14444, n14445, n14446,
         n14447, n14448, n14449, n14450, n14451, n14452, n14453, n14454,
         n14455, n14456, n14457, n14458, n14459, n14460, n14461, n14462,
         n14463, n14464, n14465, n14466, n14467, n14468, n14469, n14470,
         n14471, n14472, n14473, n14474, n14475, n14476, n14477, n14478,
         n14479, n14480, n14481, n14482, n14483, n14484, n14485, n14486,
         n14487, n14488, n14489, n14490, n14491, n14492, n14493, n14494,
         n14495, n14496, n14497, n14498, n14499, n14500, n14501, n14502,
         n14503, n14504, n14505, n14506, n14507, n14508, n14509, n14510,
         n14511, n14512, n14513, n14514, n14515, n14516, n14517, n14518,
         n14519, n14520, n14521, n14522, n14523, n14524, n14525, n14526,
         n14527, n14528, n14529, n14530, n14531, n14532, n14533, n14534,
         n14535, n14536, n14537, n14538, n14539, n14540, n14541, n14542,
         n14543, n14544, n14545, n14546, n14547, n14548, n14549, n14550,
         n14551, n14552, n14553, n14554, n14555, n14556, n14557, n14558,
         n14559, n14560, n14561, n14562, n14563, n14564, n14565, n14566,
         n14567, n14568, n14569, n14570, n14571, n14572, n14573, n14574,
         n14575, n14576, n14577, n14578, n14579, n14580, n14581, n14582,
         n14583, n14584, n14585, n14586, n14587, n14588, n14589, n14590,
         n14591, n14592, n14593, n14594, n14595, n14596, n14597, n14598,
         n14599, n14600, n14601, n14602, n14603, n14604, n14605, n14606,
         n14607, n14608, n14609, n14610, n14611, n14612, n14613, n14614,
         n14615, n14616, n14617, n14618, n14619, n14620, n14621, n14622,
         n14623, n14624, n14625, n14626, n14627, n14628, n14629, n14630,
         n14631, n14632, n14633, n14634, n14635, n14636, n14637, n14638,
         n14639, n14640, n14641, n14642, n14643, n14644, n14645, n14646,
         n14647, n14648, n14649, n14650, n14651, n14652, n14653, n14654,
         n14655, n14656, n14657, n14658, n14659, n14660, n14661, n14662,
         n14663, n14664, n14665, n14666, n14667, n14668, n14669, n14670,
         n14671, n14672, n14673, n14674, n14675, n14676, n14677, n14678,
         n14679, n14680, n14681, n14682, n14683, n14684, n14685, n14686,
         n14687, n14688, n14689, n14690, n14691, n14692, n14693, n14694,
         n14695, n14696, n14697, n14698, n14699, n14700, n14701, n14702,
         n14703, n14704, n14705, n14706, n14707, n14708, n14709, n14710,
         n14711, n14712, n14713, n14714, n14715, n14716, n14717, n14718,
         n14719, n14720, n14721, n14722, n14723, n14724, n14725, n14726,
         n14727, n14728, n14729, n14730, n14731, n14732, n14733, n14734,
         n14735, n14736, n14737, n14738, n14739, n14740, n14741, n14742,
         n14743, n14744, n14745, n14746, n14747, n14748, n14749, n14750,
         n14751, n14752, n14753, n14754, n14755, n14756, n14757, n14758,
         n14759, n14760, n14761, n14762, n14763, n14764, n14765, n14766,
         n14767, n14768, n14769, n14770, n14771, n14772, n14773, n14774,
         n14775, n14776, n14777, n14778, n14779, n14780, n14781, n14782,
         n14783, n14784, n14785, n14786, n14787, n14788, n14789, n14790,
         n14791, n14792, n14793, n14794, n14795, n14796, n14797, n14798,
         n14799, n14800, n14801, n14802, n14803, n14804, n14805, n14806,
         n14807, n14808, n14809, n14810, n14811, n14812, n14813, n14814,
         n14815, n14816, n14817, n14818, n14819, n14820, n14821, n14822,
         n14823, n14824, n14825, n14826, n14827, n14828, n14829, n14830,
         n14831, n14832, n14833, n14834, n14835, n14836, n14837, n14838,
         n14839, n14840, n14841, n14842, n14843, n14844, n14845, n14846,
         n14847, n14848, n14849, n14850, n14851, n14852, n14853, n14854,
         n14855, n14856, n14857, n14858, n14859, n14860, n14861, n14862,
         n14863, n14864, n14865, n14866, n14867, n14868, n14869, n14870,
         n14871, n14872, n14873, n14874, n14875, n14876, n14877, n14878,
         n14879, n14880, n14881, n14882, n14883, n14884, n14885, n14886,
         n14887, n14888, n14889, n14890, n14891, n14892, n14893, n14894,
         n14895, n14896, n14897, n14898, n14899, n14900, n14901, n14902,
         n14903, n14904, n14905, n14906, n14907, n14908, n14909, n14910,
         n14911, n14912, n14913, n14914, n14915, n14916, n14917, n14918,
         n14919, n14920, n14921, n14922, n14923, n14924, n14925, n14926,
         n14927, n14928, n14929, n14930, n14931, n14932, n14933, n14934,
         n14935, n14936, n14937, n14938, n14939, n14940, n14941, n14942,
         n14943, n14944, n14945, n14946, n14947, n14948, n14949, n14950,
         n14951, n14952, n14953, n14954, n14955, n14956, n14957, n14958,
         n14959, n14960, n14961, n14962, n14963, n14964, n14965, n14966,
         n14967, n14968, n14969, n14970, n14971, n14972, n14973, n14974,
         n14975, n14976, n14977, n14978, n14979, n14980, n14981, n14982,
         n14983, n14984, n14985, n14986, n14987, n14988, n14989, n14990,
         n14991, n14992, n14993, n14994, n14995, n14996, n14997, n14998,
         n14999, n15000, n15001, n15002, n15003, n15004, n15005, n15006,
         n15007, n15008, n15009, n15010, n15011, n15012, n15013, n15014,
         n15015, n15016, n15017, n15018, n15019, n15020, n15021, n15022,
         n15023, n15024, n15025, n15026, n15027, n15028, n15029, n15030,
         n15031, n15032, n15033, n15034, n15035, n15036, n15037, n15038,
         n15039, n15040, n15041, n15042, n15043, n15044, n15045, n15046,
         n15047, n15048, n15049, n15050, n15051, n15052, n15053, n15054,
         n15055, n15056, n15057, n15058, n15059, n15060, n15061, n15062,
         n15063, n15064, n15065, n15066, n15067, n15068, n15069, n15070,
         n15071, n15072, n15073, n15074, n15075, n15076, n15077, n15078,
         n15079, n15080, n15081, n15082, n15083, n15084, n15085, n15086,
         n15087, n15088, n15089, n15090, n15091, n15092, n15093, n15094,
         n15095, n15096, n15097, n15098, n15099, n15100, n15101, n15102,
         n15103, n15104, n15105, n15106, n15107, n15108, n15109, n15110,
         n15111, n15112, n15113, n15114, n15115, n15116, n15117, n15118,
         n15119, n15120, n15121, n15122, n15123, n15124, n15125, n15126,
         n15127, n15128, n15129, n15130, n15131, n15132, n15133, n15134,
         n15135, n15136, n15137, n15138, n15139, n15140, n15141, n15142,
         n15143, n15144, n15145, n15146, n15147, n15148, n15149, n15150,
         n15151, n15152, n15153, n15154, n15155, n15156, n15157, n15158,
         n15159, n15160, n15161, n15162, n15163, n15164, n15165, n15166,
         n15167, n15168, n15169, n15170, n15171, n15172, n15173, n15174,
         n15175, n15176, n15177, n15178, n15179, n15180, n15181, n15182,
         n15183, n15184, n15185, n15186, n15187, n15188, n15189, n15190,
         n15191, n15192, n15193, n15194, n15195, n15196, n15197, n15198,
         n15199, n15200, n15201, n15202, n15203, n15204, n15205, n15206,
         n15207, n15208, n15209, n15210, n15211, n15212, n15213, n15214,
         n15215, n15216, n15217, n15218, n15219, n15220, n15221, n15222,
         n15223, n15224, n15225, n15226, n15227, n15228, n15229, n15230,
         n15231, n15232, n15233, n15234, n15235, n15236, n15237, n15238,
         n15239, n15240, n15241, n15242, n15243, n15244, n15245, n15246,
         n15247, n15248, n15249, n15250, n15251, n15252, n15253, n15254,
         n15255, n15256, n15257, n15258, n15259, n15260, n15261, n15262,
         n15263, n15264, n15265, n15266, n15267, n15268, n15269, n15270,
         n15271, n15272, n15273, n15274, n15275, n15276, n15277, n15278,
         n15279, n15280, n15281, n15282, n15283, n15284, n15285, n15286,
         n15287, n15288, n15289, n15290, n15291, n15292, n15293, n15294,
         n15295, n15296, n15297, n15298, n15299, n15300, n15301, n15302,
         n15303, n15304, n15305, n15306, n15307, n15308, n15309, n15310,
         n15311, n15312, n15313, n15314, n15315, n15316, n15317, n15318,
         n15319, n15320, n15321, n15322, n15323, n15324, n15325, n15326,
         n15327, n15328, n15329, n15330, n15331, n15332, n15333, n15334,
         n15335, n15336, n15337, n15338, n15339, n15340, n15341, n15342,
         n15343, n15344, n15345, n15346, n15347, n15348, n15349, n15350,
         n15351, n15352, n15353, n15354, n15355, n15356, n15357, n15358,
         n15359, n15360, n15361, n15362, n15363, n15364, n15365, n15366,
         n15367, n15368, n15369, n15370, n15371, n15372, n15373, n15374,
         n15375, n15376, n15377, n15378, n15379, n15380, n15381, n15382,
         n15383, n15384, n15385, n15386, n15387, n15388, n15389, n15390,
         n15391, n15392, n15393, n15394, n15395, n15396, n15397, n15398,
         n15399, n15400, n15401, n15402, n15403, n15404, n15405, n15406,
         n15407, n15408, n15409, n15410, n15411, n15412, n15413, n15414,
         n15415, n15416, n15417, n15418, n15419, n15420, n15421, n15422,
         n15423, n15424, n15425, n15426, n15427, n15428, n15429, n15430,
         n15431, n15432, n15433, n15434, n15435, n15436, n15437, n15438,
         n15439, n15440, n15441, n15442, n15443, n15444, n15445, n15446,
         n15447, n15448, n15449, n15450, n15451, n15452, n15453, n15454,
         n15455, n15456, n15457, n15458, n15459, n15460, n15461, n15462,
         n15463, n15464, n15465, n15466, n15467, n15468, n15469, n15470,
         n15471, n15472, n15473, n15474, n15475, n15476, n15477, n15478,
         n15479, n15480, n15481, n15482, n15483, n15484, n15485, n15486,
         n15487, n15488, n15489, n15490, n15491, n15492, n15493, n15494,
         n15495, n15496, n15497, n15498, n15499, n15500, n15501, n15502,
         n15503, n15504, n15505, n15506, n15507, n15508, n15509, n15510,
         n15511, n15512, n15513, n15514, n15515, n15516, n15517, n15518,
         n15519, n15520, n15521, n15522, n15523, n15524, n15525, n15526,
         n15527, n15528, n15529, n15530, n15531, n15532, n15533, n15534,
         n15535, n15536, n15537, n15538, n15539, n15540, n15541, n15542,
         n15543, n15544, n15545, n15546, n15547, n15548, n15549, n15550,
         n15551, n15552, n15553, n15554, n15555, n15556, n15557, n15558,
         n15559, n15560, n15561, n15562, n15563, n15564, n15565, n15566,
         n15567, n15568, n15569, n15570, n15571, n15572, n15573, n15574,
         n15575, n15576, n15577, n15578, n15579, n15580, n15581, n15582,
         n15583, n15584, n15585, n15586, n15587, n15588, n15589, n15590,
         n15591, n15592, n15593, n15594, n15595, n15596, n15597, n15598,
         n15599, n15600, n15601, n15602, n15603, n15604, n15605, n15606,
         n15607, n15608, n15609, n15610, n15611, n15612, n15613, n15614,
         n15615, n15616, n15617, n15618, n15619, n15620, n15621, n15622,
         n15623, n15624, n15625, n15626, n15627, n15628, n15629, n15630,
         n15631, n15632, n15633, n15634, n15635, n15636, n15637, n15638,
         n15639, n15640, n15641, n15642, n15643, n15644, n15645, n15646,
         n15647, n15648, n15649, n15650, n15651, n15652, n15653, n15654,
         n15655, n15656, n15657, n15658, n15659, n15660, n15661, n15662,
         n15663, n15664, n15665, n15666, n15667, n15668, n15669, n15670,
         n15671, n15672, n15673, n15674, n15675, n15676, n15677, n15678,
         n15679, n15680, n15681, n15682, n15683, n15684, n15685, n15686,
         n15687, n15688, n15689, n15690, n15691, n15692, n15693, n15694,
         n15695, n15696, n15697, n15698, n15699, n15700, n15701, n15702,
         n15703, n15704, n15705, n15706, n15707, n15708, n15709, n15710,
         n15711, n15712, n15713, n15714, n15715, n15716, n15717, n15718,
         n15719, n15720, n15721, n15722, n15723, n15724, n15725, n15726,
         n15727, n15728, n15729, n15730, n15731, n15732, n15733, n15734,
         n15735, n15736, n15737, n15738, n15739, n15740, n15741, n15742,
         n15743, n15744, n15745, n15746, n15747, n15748, n15749, n15750,
         n15751, n15752, n15753, n15754, n15755, n15756, n15757, n15758,
         n15759, n15760, n15761, n15762, n15763, n15764, n15765, n15766,
         n15767, n15768, n15769, n15770, n15771, n15772, n15773, n15774,
         n15775, n15776, n15777, n15778, n15779, n15780, n15781, n15782,
         n15783, n15784, n15785, n15786, n15787, n15788, n15789, n15790,
         n15791, n15792, n15793, n15794, n15795, n15796, n15797, n15798,
         n15799, n15800, n15801, n15802, n15803, n15804, n15805, n15806,
         n15807, n15808, n15809, n15810, n15811, n15812, n15813, n15814,
         n15815, n15816, n15817, n15818, n15819, n15820, n15821, n15822,
         n15823, n15824, n15825, n15826, n15827, n15828, n15829, n15830,
         n15831, n15832, n15833, n15834, n15835, n15836, n15837, n15838,
         n15839, n15840, n15841, n15842, n15843, n15844, n15845, n15846,
         n15847, n15848, n15849, n15850, n15851, n15852, n15853, n15854,
         n15855, n15856, n15857, n15858, n15859, n15860, n15861, n15862,
         n15863, n15864, n15865, n15866, n15867, n15868, n15869, n15870,
         n15871, n15872, n15873, n15874, n15875, n15876, n15877, n15878,
         n15879, n15880, n15881, n15882, n15883, n15884, n15885, n15886,
         n15887, n15888, n15889, n15890, n15891, n15892, n15893, n15894,
         n15895, n15896, n15897, n15898, n15899, n15900, n15901, n15902,
         n15903, n15904, n15905, n15906, n15907, n15908, n15909, n15910,
         n15911, n15912, n15913, n15914, n15915, n15916, n15917, n15918,
         n15919, n15920, n15921, n15922, n15923, n15924, n15925, n15926,
         n15927, n15928, n15929, n15930, n15931, n15932, n15933, n15934,
         n15935, n15936, n15937, n15938, n15939, n15940, n15941, n15942,
         n15943, n15944, n15945, n15946, n15947, n15948, n15949, n15950,
         n15951, n15952, n15953, n15954, n15955, n15956, n15957, n15958,
         n15959, n15960, n15961, n15962, n15963, n15964, n15965, n15966,
         n15967, n15968, n15969, n15970, n15971, n15972, n15973, n15974,
         n15975, n15976, n15977, n15978, n15979, n15980, n15981, n15982,
         n15983, n15984, n15985, n15986, n15987, n15988, n15989, n15990,
         n15991, n15992, n15993, n15994, n15995, n15996, n15997, n15998,
         n15999, n16000, n16001, n16002, n16003, n16004, n16005, n16006,
         n16007, n16008, n16009, n16010, n16011, n16012, n16013, n16014,
         n16015, n16016, n16017, n16018, n16019, n16020, n16021, n16022,
         n16023, n16024, n16025, n16026, n16027, n16028, n16029, n16030,
         n16031, n16032, n16033, n16034, n16035, n16036, n16037, n16038,
         n16039, n16040, n16041, n16042, n16043, n16044, n16045, n16046,
         n16047, n16048, n16049, n16050, n16051, n16052, n16053, n16054,
         n16055, n16056, n16057, n16058, n16059, n16060, n16061, n16062,
         n16063, n16064, n16065, n16066, n16067, n16068, n16069, n16070,
         n16071, n16072, n16073, n16074, n16075, n16076, n16077, n16078,
         n16079, n16080, n16081, n16082, n16083, n16084, n16085, n16086,
         n16087, n16088, n16089, n16090, n16091, n16092, n16093, n16094,
         n16095, n16096, n16097, n16098, n16099, n16100, n16101, n16102,
         n16103, n16104, n16105, n16106, n16107, n16108, n16109, n16110,
         n16111, n16112, n16113, n16114, n16115, n16116, n16117, n16118,
         n16119, n16120, n16121, n16122, n16123, n16124, n16125, n16126,
         n16127, n16128, n16129, n16130, n16131, n16132, n16133, n16134,
         n16135, n16136, n16137, n16138, n16139, n16140, n16141, n16142,
         n16143, n16144, n16145, n16146, n16147, n16148, n16149, n16150,
         n16151, n16152, n16153, n16154, n16155, n16156, n16157, n16158,
         n16159, n16160, n16161, n16162, n16163, n16164, n16165, n16166,
         n16167, n16168, n16169, n16170, n16171, n16172, n16173, n16174,
         n16175, n16176, n16177, n16178, n16179, n16180, n16181, n16182,
         n16183, n16184, n16185, n16186, n16187, n16188, n16189, n16190,
         n16191, n16192, n16193, n16194, n16195, n16196, n16197, n16198,
         n16199, n16200, n16201, n16202, n16203, n16204, n16205, n16206,
         n16207, n16208, n16209, n16210, n16211, n16212, n16213, n16214,
         n16215, n16216, n16217, n16218, n16219, n16220, n16221, n16222,
         n16223, n16224, n16225, n16226, n16227, n16228, n16229, n16230,
         n16231, n16232, n16233, n16234, n16235, n16236, n16237, n16238,
         n16239, n16240, n16241, n16242, n16243, n16244, n16245, n16246,
         n16247, n16248, n16249, n16250, n16251, n16252, n16253, n16254,
         n16255, n16256, n16257, n16258, n16259, n16260, n16261, n16262,
         n16263, n16264, n16265, n16266, n16267, n16268, n16269, n16270,
         n16271, n16272, n16273, n16274, n16275, n16276, n16277, n16278,
         n16279, n16280, n16281, n16282, n16283, n16284, n16285, n16286,
         n16287, n16288, n16289, n16290, n16291, n16292, n16293, n16294,
         n16295, n16296, n16297, n16298, n16299, n16300, n16301, n16302,
         n16303, n16304, n16305, n16306, n16307, n16308, n16309, n16310,
         n16311, n16312, n16313, n16314, n16315, n16316, n16317, n16318,
         n16319, n16320, n16321, n16322, n16323, n16324, n16325, n16326,
         n16327, n16328, n16329, n16330, n16331, n16332, n16333, n16334,
         n16335, n16336, n16337, n16338, n16339, n16340, n16341, n16342,
         n16343, n16344, n16345, n16346, n16347, n16348, n16349, n16350,
         n16351, n16352, n16353, n16354, n16355, n16356, n16357, n16358,
         n16359, n16360, n16361, n16362, n16363, n16364, n16365, n16366,
         n16367, n16368, n16369, n16370, n16371, n16372, n16373, n16374,
         n16375, n16376, n16377, n16378, n16379, n16380, n16381, n16382,
         n16383, n16384, n16385, n16386, n16387, n16388, n16389, n16390,
         n16391, n16392, n16393, n16394, n16395, n16396, n16397, n16398,
         n16399, n16400, n16401, n16402, n16403, n16404, n16405, n16406,
         n16407, n16408, n16409, n16410, n16411, n16412, n16413, n16414,
         n16415, n16416, n16417, n16418, n16419, n16420, n16421, n16422,
         n16423, n16424, n16425, n16426, n16427, n16428, n16429, n16430,
         n16431, n16432, n16433, n16434, n16435, n16436, n16437, n16438,
         n16439, n16440, n16441, n16442, n16443, n16444, n16445, n16446,
         n16447, n16448, n16449, n16450, n16451, n16452, n16453, n16454,
         n16455, n16456, n16457, n16458, n16459, n16460, n16461, n16462,
         n16463, n16464, n16465, n16466, n16467, n16468, n16469, n16470,
         n16471, n16472, n16473, n16474, n16475, n16476, n16477, n16478,
         n16479, n16480, n16481, n16482, n16483, n16484, n16485, n16486,
         n16487, n16488, n16489, n16490, n16491, n16492, n16493, n16494,
         n16495, n16496, n16497, n16498, n16499, n16500, n16501, n16502,
         n16503, n16504, n16505, n16506, n16507, n16508, n16509, n16510,
         n16511, n16512, n16513, n16514, n16515, n16516, n16517, n16518,
         n16519, n16520, n16521, n16522, n16523, n16524, n16525, n16526,
         n16527, n16528, n16529, n16530, n16531, n16532, n16533, n16534,
         n16535, n16536, n16537, n16538, n16539, n16540, n16541, n16542,
         n16543, n16544, n16545, n16546, n16547, n16548, n16549, n16550,
         n16551, n16552, n16553, n16554, n16555, n16556, n16557, n16558,
         n16559, n16560, n16561, n16562, n16563, n16564, n16565, n16566,
         n16567, n16568, n16569, n16570, n16571, n16572, n16573, n16574,
         n16575, n16576, n16577, n16578, n16579, n16580, n16581, n16582,
         n16583, n16584, n16585, n16586, n16587, n16588, n16589, n16590,
         n16591, n16592, n16593, n16594, n16595, n16596, n16597, n16598,
         n16599, n16600, n16601, n16602, n16603, n16604, n16605, n16606,
         n16607, n16608, n16609, n16610, n16611, n16612, n16613, n16614,
         n16615, n16616, n16617, n16618, n16619, n16620, n16621, n16622,
         n16623, n16624, n16625, n16626, n16627, n16628, n16629, n16630,
         n16631, n16632, n16633, n16634, n16635, n16636, n16637, n16638,
         n16639, n16640, n16641, n16642, n16643, n16644, n16645, n16646,
         n16647, n16648, n16649, n16650, n16651, n16652, n16653, n16654,
         n16655, n16656, n16657, n16658, n16659, n16660, n16661, n16662,
         n16663, n16664, n16665, n16666, n16667, n16668, n16669, n16670,
         n16671, n16672, n16673, n16674, n16675, n16676, n16677, n16678,
         n16679, n16680, n16681, n16682, n16683, n16684, n16685, n16686,
         n16687, n16688, n16689, n16690, n16691, n16692, n16693, n16694,
         n16695, n16696, n16697, n16698, n16699, n16700, n16701, n16702,
         n16703, n16704, n16705, n16706, n16707, n16708, n16709, n16710,
         n16711, n16712, n16713, n16714, n16715, n16716, n16717, n16718,
         n16719, n16720, n16721, n16722, n16723, n16724, n16725, n16726,
         n16727, n16728, n16729, n16730, n16731, n16732, n16733, n16734,
         n16735, n16736, n16737, n16738, n16739, n16740, n16741, n16742,
         n16743, n16744, n16745, n16746, n16747, n16748, n16749, n16750,
         n16751, n16752, n16753, n16754, n16755, n16756, n16757, n16758,
         n16759, n16760, n16761, n16762, n16763, n16764, n16765, n16766,
         n16767, n16768, n16769, n16770, n16771, n16772, n16773, n16774,
         n16775, n16776, n16777, n16778, n16779, n16780, n16781, n16782,
         n16783, n16784, n16785, n16786, n16787, n16788, n16789, n16790,
         n16791, n16792, n16793, n16794, n16795, n16796, n16797, n16798,
         n16799, n16800, n16801, n16802, n16803, n16804, n16805, n16806,
         n16807, n16808, n16809, n16810, n16811, n16812, n16813, n16814,
         n16815, n16816, n16817, n16818, n16819, n16820, n16821, n16822,
         n16823, n16824, n16825, n16826, n16827, n16828, n16829, n16830,
         n16831, n16832, n16833, n16834, n16835, n16836, n16837, n16838,
         n16839, n16840, n16841, n16842, n16843, n16844, n16845, n16846,
         n16847, n16848, n16849, n16850, n16851, n16852, n16853, n16854,
         n16855, n16856, n16857, n16858, n16859, n16860, n16861, n16862,
         n16863, n16864, n16865, n16866, n16867, n16868, n16869, n16870,
         n16871, n16872, n16873, n16874, n16875, n16876, n16877, n16878,
         n16879, n16880, n16881, n16882, n16883, n16884, n16885, n16886,
         n16887, n16888, n16889, n16890, n16891, n16892, n16893, n16894,
         n16895, n16896, n16897, n16898, n16899, n16900, n16901, n16902,
         n16903, n16904, n16905, n16906, n16907, n16908, n16909, n16910,
         n16911, n16912, n16913, n16914, n16915, n16916, n16917, n16918,
         n16919, n16920, n16921, n16922, n16923, n16924, n16925, n16926,
         n16927, n16928, n16929, n16930, n16931, n16932, n16933, n16934,
         n16935, n16936, n16937, n16938, n16939, n16940, n16941, n16942,
         n16943, n16944, n16945, n16946, n16947, n16948, n16949, n16950,
         n16951, n16952, n16953, n16954, n16955, n16956, n16957, n16958,
         n16959, n16960, n16961, n16962, n16963, n16964, n16965, n16966,
         n16967, n16968, n16969, n16970, n16971, n16972, n16973, n16974,
         n16975, n16976, n16977, n16978, n16979, n16980, n16981, n16982,
         n16983, n16984, n16985, n16986, n16987, n16988, n16989, n16990,
         n16991, n16992, n16993, n16994, n16995, n16996, n16997, n16998,
         n16999, n17000, n17001, n17002, n17003, n17004, n17005, n17006,
         n17007, n17008, n17009, n17010, n17011, n17012, n17013, n17014,
         n17015, n17016, n17017, n17018, n17019, n17020, n17021, n17022,
         n17023, n17024, n17025, n17026, n17027, n17028, n17029, n17030,
         n17031, n17032, n17033, n17034, n17035, n17036, n17037, n17038,
         n17039, n17040, n17041, n17042, n17043, n17044, n17045, n17046,
         n17047, n17048, n17049, n17050, n17051, n17052, n17053, n17054,
         n17055, n17056, n17057, n17058, n17059, n17060, n17061, n17062,
         n17063, n17064, n17065, n17066, n17067, n17068, n17069, n17070,
         n17071, n17072, n17073, n17074, n17075, n17076, n17077, n17078,
         n17079, n17080, n17081, n17082, n17083, n17084, n17085, n17086,
         n17087, n17088, n17089, n17090, n17091, n17092, n17093, n17094,
         n17095, n17096, n17097, n17098, n17099, n17100, n17101, n17102,
         n17103, n17104, n17105, n17106, n17107, n17108, n17109, n17110,
         n17111, n17112, n17113, n17114, n17115, n17116, n17117, n17118,
         n17119, n17120, n17121, n17122, n17123, n17124, n17125, n17126,
         n17127, n17128, n17129, n17130, n17131, n17132, n17133, n17134,
         n17135, n17136, n17137, n17138, n17139, n17140, n17141, n17142,
         n17143, n17144, n17145, n17146, n17147, n17148, n17149, n17150,
         n17151, n17152, n17153, n17154, n17155, n17156, n17157, n17158,
         n17159, n17160, n17161, n17162, n17163, n17164, n17165, n17166,
         n17167, n17168, n17169, n17170, n17171, n17172, n17173, n17174,
         n17175, n17176, n17177, n17178, n17179, n17180, n17181, n17182,
         n17183, n17184, n17185, n17186, n17187, n17188, n17189, n17190,
         n17191, n17192, n17193, n17194, n17195, n17196, n17197, n17198,
         n17199, n17200, n17201, n17202, n17203, n17204, n17205, n17206,
         n17207, n17208, n17209, n17210, n17211, n17212, n17213, n17214,
         n17215, n17216, n17217, n17218, n17219, n17220, n17221, n17222,
         n17223, n17224, n17225, n17226, n17227, n17228, n17229, n17230,
         n17231, n17232, n17233, n17234, n17235, n17236, n17237, n17238,
         n17239, n17240, n17241, n17242, n17243, n17244, n17245, n17246,
         n17247, n17248, n17249, n17250, n17251, n17252, n17253, n17254,
         n17255, n17256, n17257, n17258, n17259, n17260, n17261, n17262,
         n17263, n17264, n17265, n17266, n17267, n17268, n17269, n17270,
         n17271, n17272, n17273, n17274, n17275, n17276, n17277, n17278,
         n17279, n17280, n17281, n17282, n17283, n17284, n17285, n17286,
         n17287, n17288, n17289, n17290, n17291, n17292, n17293, n17294,
         n17295, n17296, n17297, n17298, n17299, n17300, n17301, n17302,
         n17303, n17304, n17305, n17306, n17307, n17308, n17309, n17310,
         n17311, n17312, n17313, n17314, n17315, n17316, n17317, n17318,
         n17319, n17320, n17321, n17322, n17323, n17324, n17325, n17326,
         n17327, n17328, n17329, n17330, n17331, n17332, n17333, n17334,
         n17335, n17336, n17337, n17338, n17339, n17340, n17341, n17342,
         n17343, n17344, n17345, n17346, n17347, n17348, n17349, n17350,
         n17351, n17352, n17353, n17354, n17355, n17356, n17357, n17358,
         n17359, n17360, n17361, n17362, n17363, n17364, n17365, n17366,
         n17367, n17368, n17369, n17370, n17371, n17372, n17373, n17374,
         n17375, n17376, n17377, n17378, n17379, n17380, n17381, n17382,
         n17383, n17384, n17385, n17386, n17387, n17388, n17389, n17390,
         n17391, n17392, n17393, n17394, n17395, n17396, n17397, n17398,
         n17399, n17400, n17401, n17402, n17403, n17404, n17405, n17406,
         n17407, n17408, n17409, n17410, n17411, n17412, n17413, n17414,
         n17415, n17416, n17417, n17418, n17419, n17420, n17421, n17422,
         n17423, n17424, n17425, n17426, n17427, n17428, n17429, n17430,
         n17431, n17432, n17433, n17434, n17435, n17436, n17437, n17438,
         n17439, n17440, n17441, n17442, n17443, n17444, n17445, n17446,
         n17447, n17448, n17449, n17450, n17451, n17452, n17453, n17454,
         n17455, n17456, n17457, n17458, n17459, n17460, n17461, n17462,
         n17463, n17464, n17465, n17466, n17467, n17468, n17469, n17470,
         n17471, n17472, n17473, n17474, n17475, n17476, n17477, n17478,
         n17479, n17480, n17481, n17482, n17483, n17484, n17485, n17486,
         n17487, n17488, n17489, n17490, n17491, n17492, n17493, n17494,
         n17495, n17496, n17497, n17498, n17499, n17500, n17501, n17502,
         n17503, n17504, n17505, n17506, n17507, n17508, n17509, n17510,
         n17511, n17512, n17513, n17514, n17515, n17516, n17517, n17518,
         n17519, n17520, n17521, n17522, n17523, n17524, n17525, n17526,
         n17527, n17528, n17529, n17530, n17531, n17532, n17533, n17534,
         n17535, n17536, n17537, n17538, n17539, n17540, n17541, n17542,
         n17543, n17544, n17545, n17546, n17547, n17548, n17549, n17550,
         n17551, n17552, n17553, n17554, n17555, n17556, n17557, n17558,
         n17559, n17560, n17561, n17562, n17563, n17564, n17565, n17566,
         n17567, n17568, n17569, n17570, n17571, n17572, n17573, n17574,
         n17575, n17576, n17577, n17578, n17579, n17580, n17581, n17582,
         n17583, n17584, n17585, n17586, n17587, n17588, n17589, n17590,
         n17591, n17592, n17593, n17594, n17595, n17596, n17597, n17598,
         n17599, n17600, n17601, n17602, n17603, n17604, n17605, n17606,
         n17607, n17608, n17609, n17610, n17611, n17612, n17613, n17614,
         n17615, n17616, n17617, n17618, n17619, n17620, n17621, n17622,
         n17623, n17624, n17625, n17626, n17627, n17628, n17629, n17630,
         n17631, n17632, n17633, n17634, n17635, n17636, n17637, n17638,
         n17639, n17640, n17641, n17642, n17643, n17644, n17645, n17646,
         n17647, n17648, n17649, n17650, n17651, n17652, n17653, n17654,
         n17655, n17656, n17657, n17658, n17659, n17660, n17661, n17662,
         n17663, n17664, n17665, n17666, n17667, n17668, n17669, n17670,
         n17671, n17672, n17673, n17674, n17675, n17676, n17677, n17678,
         n17679, n17680, n17681, n17682, n17683, n17684, n17685, n17686,
         n17687, n17688, n17689, n17690, n17691, n17692, n17693, n17694,
         n17695, n17696, n17697, n17698, n17699, n17700, n17701, n17702,
         n17703, n17704, n17705, n17706, n17707, n17708, n17709, n17710,
         n17711, n17712, n17713, n17714, n17715, n17716, n17717, n17718,
         n17719, n17720, n17721, n17722, n17723, n17724, n17725, n17726,
         n17727, n17728, n17729, n17730, n17731, n17732, n17733, n17734,
         n17735, n17736, n17737, n17738, n17739, n17740, n17741, n17742,
         n17743, n17744, n17745, n17746, n17747, n17748, n17749, n17750,
         n17751, n17752, n17753, n17754, n17755, n17756, n17757, n17758,
         n17759, n17760, n17761, n17762, n17763, n17764, n17765, n17766,
         n17767, n17768, n17769, n17770, n17771, n17772, n17773, n17774,
         n17775, n17776, n17777, n17778, n17779, n17780, n17781, n17782,
         n17783, n17784, n17785, n17786, n17787, n17788, n17789, n17790,
         n17791, n17792, n17793, n17794, n17795, n17796, n17797, n17798,
         n17799, n17800, n17801, n17802, n17803, n17804, n17805, n17806,
         n17807, n17808, n17809, n17810, n17811, n17812, n17813, n17814,
         n17815, n17816, n17817, n17818, n17819, n17820, n17821, n17822,
         n17823, n17824, n17825, n17826, n17827, n17828, n17829, n17830,
         n17831, n17832, n17833, n17834, n17835, n17836, n17837, n17838,
         n17839, n17840, n17841, n17842, n17843, n17844, n17845, n17846,
         n17847, n17848, n17849, n17850, n17851, n17852, n17853, n17854,
         n17855, n17856, n17857, n17858, n17859, n17860, n17861, n17862,
         n17863, n17864, n17865, n17866, n17867, n17868, n17869, n17870,
         n17871, n17872, n17873, n17874, n17875, n17876, n17877, n17878,
         n17879, n17880, n17881, n17882, n17883, n17884, n17885, n17886,
         n17887, n17888, n17889, n17890, n17891, n17892, n17893, n17894,
         n17895, n17896, n17897, n17898, n17899, n17900, n17901, n17902,
         n17903, n17904, n17905, n17906, n17907, n17908, n17909, n17910,
         n17911, n17912, n17913, n17914, n17915, n17916, n17917, n17918,
         n17919, n17920, n17921, n17922, n17923, n17924, n17925, n17926,
         n17927, n17928, n17929, n17930, n17931, n17932, n17933, n17934,
         n17935, n17936, n17937, n17938, n17939, n17940, n17941, n17942,
         n17943, n17944, n17945, n17946, n17947, n17948, n17949, n17950,
         n17951, n17952, n17953, n17954, n17955, n17956, n17957, n17958,
         n17959, n17960, n17961, n17962, n17963, n17964, n17965, n17966,
         n17967, n17968, n17969, n17970, n17971, n17972, n17973, n17974,
         n17975, n17976, n17977, n17978, n17979, n17980, n17981, n17982,
         n17983, n17984, n17985, n17986, n17987, n17988, n17989, n17990,
         n17991, n17992, n17993, n17994, n17995, n17996, n17997, n17998,
         n17999, n18000, n18001, n18002, n18003, n18004, n18005, n18006,
         n18007, n18008, n18009, n18010, n18011, n18012, n18013, n18014,
         n18015, n18016, n18017, n18018, n18019, n18020, n18021, n18022,
         n18023, n18024, n18025, n18026, n18027, n18028, n18029, n18030,
         n18031, n18032, n18033, n18034, n18035, n18036, n18037, n18038,
         n18039, n18040, n18041, n18042, n18043, n18044, n18045, n18046,
         n18047, n18048, n18049, n18050, n18051, n18052, n18053, n18054,
         n18055, n18056, n18057, n18058, n18059, n18060, n18061, n18062,
         n18063, n18064, n18065, n18066, n18067, n18068, n18069, n18070,
         n18071, n18072, n18073, n18074, n18075, n18076, n18077, n18078,
         n18079, n18080, n18081, n18082, n18083, n18084, n18085, n18086,
         n18087, n18088, n18089, n18090, n18091, n18092, n18093, n18094,
         n18095, n18096, n18097, n18098, n18099, n18100, n18101, n18102,
         n18103, n18104, n18105, n18106, n18107, n18108, n18109, n18110,
         n18111, n18112, n18113, n18114, n18115, n18116, n18117, n18118,
         n18119, n18120, n18121, n18122, n18123, n18124, n18125, n18126,
         n18127, n18128, n18129, n18130, n18131, n18132, n18133, n18134,
         n18135, n18136, n18137, n18138, n18139, n18140, n18141, n18142,
         n18143, n18144, n18145, n18146, n18147, n18148, n18149, n18150,
         n18151, n18152, n18153, n18154, n18155, n18156, n18157, n18158,
         n18159, n18160, n18161, n18162, n18163, n18164, n18165, n18166,
         n18167, n18168, n18169, n18170, n18171, n18172, n18173, n18174,
         n18175, n18176, n18177, n18178, n18179, n18180, n18181, n18182,
         n18183, n18184, n18185, n18186, n18187, n18188, n18189, n18190,
         n18191, n18192, n18193, n18194, n18195, n18196, n18197, n18198,
         n18199, n18200, n18201, n18202, n18203, n18204, n18205, n18206,
         n18207, n18208, n18209, n18210, n18211, n18212, n18213, n18214,
         n18215, n18216, n18217, n18218, n18219, n18220, n18221, n18222,
         n18223, n18224, n18225, n18226, n18227, n18228, n18229, n18230,
         n18231, n18232, n18233, n18234, n18235, n18236, n18237, n18238,
         n18239, n18240, n18241, n18242, n18243, n18244, n18245, n18246,
         n18247, n18248, n18249, n18250, n18251, n18252, n18253, n18254,
         n18255, n18256, n18257, n18258, n18259, n18260, n18261, n18262,
         n18263, n18264, n18265, n18266, n18268, n18269, n18270, n18271,
         n18272, n18273, n18274, n18275, n18276, n18277, n18278, n18279,
         n18280, n18281, n18282, n18283, n18284, n18285, n18286, n18287,
         n18288, n18289, n18290, n18291, n18292, n18293, n18294, n18295,
         n18296, n18297, n18298, n18299, n18300, n18301, n18302, n18303,
         n18304, n18305, n18306, n18307, n18308, n18309, n18310, n18311,
         n18312, n18313, n18314, n18315, n18316, n18317, n18318, n18319,
         n18320, n18321, n18322, n18323, n18324, n18325, n18326, n18327,
         n18328, n18329, n18330, n18331, n18332, n18333, n18334, n18335,
         n18336, n18337, n18338, n18339, n18340, n18341, n18342, n18343,
         n18344, n18345, n18346, n18347, n18348, n18349, n18350, n18351,
         n18352, n18353, n18354, n18355, n18356, n18357, n18358, n18359,
         n18360, n18361, n18362, n18363, n18364, n18365, n18366, n18367,
         n18368, n18369, n18370, n18371, n18372, n18373, n18374, n18375,
         n18376, n18377, n18378, n18379, n18380, n18381, n18382, n18383,
         n18384, n18385, n18386, n18387, n18388, n18389, n18390, n18391,
         n18392, n18393, n18394, n18395, n18396, n18397, n18398, n18399,
         n18400, n18401, n18402, n18403, n18404, n18405, n18406, n18407,
         n18408, n18409, n18410, n18411, n18412, n18413, n18414, n18415,
         n18416, n18417, n18418, n18419, n18420, n18421, n18422, n18423,
         n18424, n18425, n18426, n18427, n18428, n18429, n18430, n18431,
         n18432, n18433, n18434, n18435, n18436, n18437, n18438, n18439,
         n18440, n18441, n18442, n18443, n18444, n18445, n18446, n18447,
         n18448, n18449, n18450, n18451, n18452, n18453, n18454, n18455,
         n18456, n18457, n18458, n18459, n18460, n18461, n18462, n18463,
         n18464, n18465, n18466, n18467, n18468, n18469, n18470, n18471,
         n18472, n18473, n18474, n18475, n18476, n18477, n18478, n18479,
         n18480, n18481, n18482, n18483, n18484, n18485, n18486, n18487,
         n18488, n18489, n18490, n18491, n18492, n18493, n18494, n18495,
         n18496, n18497, n18498, n18499, n18500, n18501, n18502, n18503,
         n18504, n18505, n18506, n18507, n18508, n18509, n18510, n18511,
         n18512, n18513, n18514, n18515, n18516, n18517, n18518, n18519,
         n18520, n18521, n18522, n18523, n18524, n18525, n18526, n18527,
         n18528, n18529, n18530, n18531, n18532, n18533, n18534, n18535,
         n18536, n18537, n18538, n18539, n18540, n18541, n18542, n18543,
         n18544, n18545, n18546, n18547, n18548, n18549, n18550, n18551,
         n18552, n18553, n18554, n18555, n18556, n18557, n18558, n18559,
         n18560, n18561, n18562, n18563, n18564, n18565, n18566, n18567,
         n18568, n18569, n18570, n18571, n18572, n18573, n18574, n18575,
         n18576, n18577, n18578, n18579, n18580, n18581, n18582, n18583,
         n18584, n18585, n18586, n18587, n18588, n18589, n18590, n18591,
         n18592, n18593, n18594, n18595, n18596, n18597, n18598, n18599,
         n18600, n18601, n18602, n18603, n18604, n18605, n18606, n18607,
         n18608, n18609, n18610, n18611, n18612, n18613, n18614, n18615,
         n18616, n18617, n18618, n18619, n18620, n18621, n18622, n18623,
         n18624, n18625, n18626, n18627, n18628, n18629, n18630, n18631,
         n18632, n18633, n18634, n18635, n18636, n18637, n18638, n18639,
         n18640, n18641, n18642, n18643, n18644, n18645, n18646, n18647,
         n18648, n18649, n18650, n18651, n18652, n18653, n18654, n18655,
         n18656, n18657, n18658, n18659, n18660, n18661, n18662, n18663,
         n18664, n18665, n18666, n18667, n18668, n18669, n18670, n18671,
         n18672, n18673, n18674, n18675, n18676, n18677, n18678, n18679,
         n18680, n18681, n18682, n18683, n18684, n18685, n18686, n18687,
         n18688, n18689, n18690, n18691, n18692, n18693, n18694, n18695,
         n18696, n18697, n18698, n18699, n18700, n18701, n18702, n18703,
         n18704, n18705, n18706, n18707, n18708, n18709, n18710, n18711,
         n18712, n18713, n18714, n18715, n18716, n18717, n18718, n18719,
         n18720, n18721, n18722, n18723, n18724, n18725, n18726, n18727,
         n18728, n18729, n18730, n18731, n18732, n18733, n18734, n18735,
         n18736, n18737, n18738, n18739, n18740, n18741, n18742, n18743,
         n18744, n18745, n18746, n18747, n18748, n18749, n18750, n18751,
         n18752, n18753, n18754, n18755, n18756, n18757, n18758, n18759,
         n18760, n18761, n18762, n18763, n18764, n18765, n18766, n18767,
         n18768, n18769, n18770, n18771, n18772, n18773, n18774, n18775,
         n18776, n18777, n18778, n18779, n18780, n18781, n18782, n18783,
         n18784, n18785, n18786, n18787, n18788, n18789, n18790, n18791,
         n18792, n18793, n18794, n18795, n18796, n18797, n18798, n18799,
         n18800, n18801, n18802, n18803, n18804, n18805, n18806, n18807,
         n18808, n18809, n18810, n18811, n18812, n18813, n18814, n18815,
         n18816, n18817, n18818, n18819, n18820, n18821, n18822, n18823,
         n18824, n18825, n18826, n18827, n18828, n18829, n18830, n18831,
         n18832, n18833, n18834, n18835, n18836, n18837, n18838, n18839,
         n18840, n18841, n18842, n18843, n18844, n18845, n18846, n18847,
         n18848, n18849, n18850, n18851, n18852, n18853, n18854, n18855,
         n18856, n18857, n18858, n18859, n18860, n18861, n18862, n18863,
         n18864, n18865, n18866, n18867, n18868, n18869, n18870, n18871,
         n18872, n18873, n18874, n18875, n18876, n18877, n18878, n18879,
         n18880, n18881, n18882, n18883, n18884, n18885, n18886, n18887,
         n18888, n18889, n18890, n18891, n18892, n18893, n18894, n18895,
         n18896, n18897, n18898, n18899, n18900, n18901, n18902, n18903,
         n18904, n18905, n18906, n18907, n18908, n18909, n18910, n18911,
         n18912, n18913, n18914, n18915, n18916, n18917, n18918, n18919,
         n18920, n18921, n18922, n18923, n18924, n18925, n18926, n18927,
         n18928, n18929, n18930, n18931, n18932, n18933, n18934, n18935,
         n18936, n18937, n18938, n18939, n18940, n18941, n18942, n18943,
         n18944, n18945, n18946, n18947, n18948, n18949, n18950, n18951,
         n18952, n18953, n18954, n18955, n18956, n18957, n18958, n18959,
         n18960, n18961, n18962, n18963, n18964, n18965, n18966, n18967,
         n18968, n18969, n18970, n18971, n18972, n18973, n18974, n18975,
         n18976, n18977, n18978, n18979, n18980, n18981, n18982, n18983,
         n18984, n18985, n18986, n18987, n18988, n18989, n18990, n18991,
         n18992, n18993, n18994, n18995, n18996, n18997, n18998, n18999,
         n19000, n19001, n19002, n19003, n19004, n19005, n19006, n19007,
         n19008, n19009, n19010, n19011, n19012, n19013, n19014, n19015,
         n19016, n19017, n19018, n19019, n19020, n19021, n19022, n19023,
         n19024, n19025, n19026, n19027, n19028, n19029, n19030, n19031,
         n19032, n19033, n19034, n19035, n19036, n19037, n19038, n19039,
         n19040, n19041, n19042, n19043, n19044, n19045, n19046, n19047,
         n19048, n19049, n19050, n19051, n19052, n19053, n19054, n19055,
         n19056, n19057, n19058, n19059, n19060, n19061, n19062, n19063,
         n19064, n19065, n19066, n19067, n19068, n19069, n19070, n19071,
         n19072, n19073, n19074, n19075, n19076, n19077, n19078, n19079,
         n19080, n19081, n19082, n19083, n19084, n19085, n19086, n19087,
         n19088, n19089, n19090, n19091, n19092, n19093, n19094, n19095,
         n19096, n19097, n19098, n19099, n19100, n19101, n19102, n19103,
         n19104, n19105, n19106, n19107, n19108, n19109, n19110, n19111,
         n19112, n19113, n19114, n19115, n19116, n19117, n19118, n19119,
         n19120, n19121, n19122, n19123, n19124, n19125, n19126, n19127,
         n19128, n19129, n19130, n19131, n19132, n19133, n19134, n19135,
         n19136, n19137, n19138, n19139, n19140, n19141, n19142, n19143,
         n19144, n19145, n19146, n19147, n19148, n19149, n19150, n19151,
         n19152, n19153, n19154, n19155, n19156, n19157, n19158, n19159,
         n19160, n19161, n19162, n19163, n19164, n19165, n19166, n19167,
         n19168, n19169, n19170, n19171, n19172, n19173, n19174, n19175,
         n19176, n19177, n19178, n19179, n19180, n19181, n19182, n19183,
         n19184, n19185, n19186, n19187, n19188, n19189, n19190, n19191,
         n19192, n19193, n19194, n19195, n19196, n19197, n19198, n19199,
         n19200, n19201, n19202, n19203, n19204, n19205, n19206, n19207,
         n19208, n19209, n19210, n19211, n19212, n19213, n19214, n19215,
         n19216, n19217, n19218, n19219, n19220, n19221, n19222, n19223,
         n19224, n19225, n19226, n19227, n19228, n19229, n19230, n19231,
         n19232, n19233, n19234, n19235, n19236, n19237, n19238, n19239,
         n19240, n19241, n19242, n19243, n19244, n19245, n19246, n19247,
         n19248, n19249, n19250, n19251, n19252, n19253, n19254, n19255,
         n19256, n19257, n19258, n19259, n19260, n19261, n19262, n19263,
         n19264, n19265, n19266, n19267, n19268, n19269, n19270, n19271,
         n19272, n19273, n19274, n19275, n19276, n19277, n19278, n19279,
         n19280, n19281, n19282, n19283, n19284, n19285, n19286, n19287,
         n19288, n19289, n19290, n19291, n19292, n19293, n19294, n19295,
         n19296, n19297, n19298, n19299, n19300, n19301, n19302, n19303,
         n19304, n19305, n19306, n19307, n19308, n19309, n19310, n19311,
         n19312, n19313, n19314, n19315, n19316, n19317, n19318, n19319,
         n19320, n19321, n19322, n19323, n19324, n19325, n19326, n19327,
         n19328, n19329, n19330, n19331, n19332, n19333, n19334, n19335,
         n19336, n19337, n19338, n19339, n19340, n19341, n19342, n19343,
         n19344, n19345, n19346, n19347, n19348, n19349, n19350, n19351,
         n19352, n19353, n19354, n19355, n19356, n19357, n19358, n19359,
         n19360, n19361, n19362, n19363, n19364, n19365, n19366, n19367,
         n19368, n19369, n19370, n19371, n19372, n19373, n19374, n19375,
         n19376, n19377, n19378, n19379, n19380, n19381, n19382, n19383,
         n19384, n19385, n19386, n19387, n19388, n19389, n19390, n19391,
         n19392, n19393, n19394, n19395, n19396, n19397, n19398, n19399,
         n19400, n19401, n19402, n19403, n19404, n19405, n19406, n19407,
         n19408, n19409, n19410, n19411, n19412, n19413, n19414, n19415,
         n19416, n19417, n19418, n19419, n19420, n19421, n19422, n19423,
         n19424, n19425, n19426, n19427, n19428, n19429, n19430, n19431,
         n19432, n19433, n19434, n19435, n19436, n19437, n19438, n19439,
         n19440, n19441, n19442, n19443, n19444, n19445, n19446, n19447,
         n19448, n19449, n19450, n19451, n19452, n19453, n19454, n19455,
         n19456, n19457, n19458, n19459, n19460, n19461, n19462, n19463,
         n19464, n19465, n19466, n19467, n19468, n19469, n19470, n19471,
         n19472, n19473, n19474, n19475, n19476, n19477, n19478, n19479,
         n19480, n19481, n19482, n19483, n19484, n19485, n19486, n19487,
         n19488, n19489, n19490, n19491, n19492, n19493, n19494, n19495,
         n19496, n19497, n19498, n19499, n19500, n19501, n19502, n19503,
         n19504, n19505, n19506, n19507, n19508, n19509, n19510, n19511,
         n19512, n19513, n19514, n19515, n19516, n19517, n19518, n19519,
         n19520, n19521, n19522, n19523, n19524, n19525, n19526, n19527,
         n19528, n19529, n19530, n19531, n19532, n19533, n19534, n19535,
         n19536, n19537, n19538, n19539, n19540, n19541, n19542, n19543,
         n19544, n19545, n19546, n19547, n19548, n19549, n19550, n19551,
         n19552, n19553, n19554, n19555, n19556, n19557, n19558, n19559,
         n19560, n19561, n19562, n19563, n19564, n19565, n19566, n19567,
         n19568, n19569, n19570, n19571, n19572, n19573, n19574, n19575,
         n19576, n19577, n19578, n19579, n19580, n19581, n19582, n19583,
         n19584, n19585, n19586, n19587, n19588, n19589, n19590, n19591,
         n19592, n19593, n19594, n19595, n19596, n19597, n19598, n19599,
         n19600, n19601, n19602, n19603, n19604, n19605, n19606, n19607,
         n19608, n19609, n19610, n19611, n19612, n19613, n19614, n19615,
         n19616, n19617, n19618, n19619, n19620, n19621, n19622, n19623,
         n19624, n19625, n19626, n19627, n19628, n19629, n19630, n19631,
         n19632, n19633, n19634, n19635, n19636, n19637, n19638, n19639,
         n19640, n19641, n19642, n19643, n19644, n19645, n19646, n19647,
         n19648, n19649, n19650, n19651, n19652, n19653, n19654, n19655,
         n19656, n19657, n19658, n19659, n19660, n19661, n19662, n19663,
         n19664, n19665, n19666, n19667, n19668, n19669, n19670, n19671,
         n19672, n19673, n19674, n19675, n19676, n19677, n19678, n19679,
         n19680, n19681, n19682, n19683, n19684, n19685, n19686, n19687,
         n19688, n19689, n19690, n19691, n19692, n19693, n19694, n19695,
         n19696, n19697, n19698, n19699, n19700, n19701, n19702, n19703,
         n19704, n19705, n19706, n19707, n19708, n19709, n19710, n19711,
         n19712, n19713, n19714, n19715, n19716, n19717, n19718, n19719,
         n19720, n19721, n19722, n19723, n19724, n19725, n19726, n19727,
         n19728, n19729, n19730, n19731, n19732, n19733, n19734, n19735,
         n19736, n19737, n19738, n19739, n19740, n19741, n19742, n19743,
         n19744, n19745, n19746, n19747, n19748, n19749, n19750, n19751,
         n19752, n19753, n19754, n19755, n19756, n19757, n19758, n19759,
         n19760, n19761, n19762, n19763, n19764, n19765, n19766, n19767,
         n19768, n19769, n19770, n19771, n19772, n19773, n19774, n19775,
         n19776, n19777, n19778, n19779, n19780, n19781, n19782, n19783,
         n19784, n19785, n19786, n19787, n19788, n19789, n19790, n19791,
         n19792, n19793, n19794, n19795, n19796, n19797, n19798, n19799,
         n19800, n19801, n19802, n19803, n19804, n19805, n19806, n19807,
         n19808, n19809, n19810, n19811, n19812, n19813, n19814, n19815,
         n19816, n19817, n19818, n19819, n19820, n19821, n19822, n19823,
         n19824, n19825, n19826, n19827, n19828, n19829, n19830, n19831,
         n19832, n19833, n19834, n19835, n19836, n19837, n19838, n19839,
         n19840, n19841, n19842, n19843, n19844, n19845, n19846, n19847,
         n19848, n19849, n19850, n19851, n19852, n19853, n19854, n19855,
         n19856, n19857, n19858, n19859, n19860, n19861, n19862, n19863,
         n19864, n19865, n19866, n19867, n19868, n19869, n19870, n19871,
         n19872, n19873, n19874, n19875, n19876, n19877, n19878, n19879,
         n19880, n19881, n19882, n19883, n19884, n19885, n19886, n19887,
         n19888, n19889, n19890, n19891, n19892, n19893, n19894, n19895,
         n19896, n19897, n19898, n19899, n19900, n19901, n19902, n19903,
         n19904, n19905, n19906, n19907, n19908, n19909, n19910, n19911,
         n19912, n19913, n19914, n19915, n19916, n19917, n19918, n19919,
         n19920, n19921, n19922, n19923, n19924, n19925, n19926, n19927,
         n19928, n19929, n19930, n19931, n19932, n19933, n19934, n19935,
         n19936, n19937, n19938, n19939, n19940, n19941, n19942, n19943,
         n19944, n19945, n19946, n19947, n19948, n19949, n19950, n19951,
         n19952, n19953, n19954, n19955, n19956, n19957, n19958, n19959,
         n19960, n19961, n19962, n19963, n19964, n19965, n19966, n19967,
         n19968, n19969, n19970, n19971, n19972, n19973, n19974, n19975,
         n19976, n19977, n19978, n19979, n19980, n19981, n19982, n19983,
         n19984, n19985, n19986, n19987, n19988, n19989, n19990, n19991,
         n19992, n19993, n19994, n19995, n19996, n19997, n19998, n19999,
         n20000, n20001, n20002, n20003, n20004, n20005, n20006, n20007,
         n20008, n20009, n20010, n20011, n20012, n20013, n20014, n20015,
         n20016, n20017, n20018, n20019, n20020, n20021, n20022, n20023,
         n20024, n20025, n20026, n20027, n20028, n20029, n20030, n20031,
         n20032, n20033, n20034, n20035, n20036, n20037, n20038, n20039,
         n20040, n20041, n20042, n20043, n20044, n20045, n20046, n20047,
         n20048, n20049, n20050, n20051, n20052, n20053, n20054, n20055,
         n20056, n20057, n20058, n20059, n20060, n20061, n20062, n20063,
         n20064, n20065, n20066, n20067, n20068, n20069, n20070, n20071,
         n20072, n20073, n20074, n20075, n20076, n20077, n20078, n20079,
         n20080, n20081, n20082, n20083, n20084, n20085, n20086, n20087,
         n20088, n20089, n20090, n20091, n20092, n20093, n20094, n20095,
         n20096, n20097, n20098, n20099, n20100, n20101, n20102, n20103,
         n20105, n20106, n20107, n20108, n20109, n20110, n20111, n20112,
         n20113, n20114, n20115, n20116, n20117, n20118, n20119, n20120,
         n20121, n20122, n20123, n20124, n20125, n20126, n20127, n20128,
         n20129, n20130, n20131, n20132, n20133, n20134, n20135, n20136,
         n20137, n20138, n20139, n20140, n20141, n20142, n20143, n20144,
         n20145, n20146, n20147, n20148, n20149, n20150, n20151, n20152,
         n20153, n20154, n20155, n20156, n20157, n20158, n20159, n20160,
         n20161, n20162, n20163, n20164, n20165, n20166, n20167, n20168,
         n20169, n20170, n20171, n20172, n20173, n20174, n20175, n20176,
         n20177, n20178, n20179, n20180, n20181, n20182, n20183, n20184,
         n20185, n20186, n20187, n20188, n20189, n20190, n20191, n20192,
         n20193, n20194, n20195, n20196, n20197, n20198, n20199, n20200,
         n20201, n20202, n20203, n20204, n20205, n20206, n20207, n20208,
         n20209, n20210, n20211, n20212, n20213, n20214, n20215, n20216,
         n20217, n20218, n20219, n20220, n20221, n20222, n20223, n20224,
         n20225, n20226, n20227, n20228, n20229, n20230, n20231, n20232,
         n20233, n20234, n20235, n20236, n20237, n20238, n20239, n20240,
         n20241, n20242, n20243, n20244, n20245, n20246, n20247, n20248,
         n20249, n20250, n20251, n20252, n20253, n20254, n20255, n20256,
         n20257, n20258, n20259, n20260, n20261, n20262, n20263, n20264,
         n20265, n20266, n20267, n20268, n20269, n20270, n20271, n20272,
         n20273, n20274, n20275, n20276, n20277, n20278, n20279, n20280,
         n20281, n20282, n20283, n20284, n20285, n20286, n20287, n20288,
         n20289, n20290, n20291, n20292, n20293, n20294, n20295, n20296,
         n20297, n20298, n20299, n20300, n20301, n20302, n20303, n20304,
         n20305, n20306, n20307, n20308, n20309, n20310, n20311, n20312,
         n20313, n20314, n20315, n20316, n20317, n20318, n20319, n20320,
         n20321, n20322, n20323, n20324, n20325, n20326, n20327, n20328,
         n20329, n20330, n20331, n20332, n20333, n20334, n20335, n20336,
         n20337, n20338, n20339, n20340, n20341, n20342, n20343, n20344,
         n20345, n20346, n20347, n20348, n20349, n20350, n20351, n20352,
         n20353, n20354, n20355, n20356, n20357, n20358, n20359, n20360,
         n20361, n20362, n20363, n20364, n20365, n20366, n20367, n20368,
         n20369, n20370, n20371, n20372, n20373, n20374, n20375, n20376,
         n20377, n20378, n20379, n20380, n20381, n20382, n20383, n20384,
         n20385, n20386, n20387, n20388, n20389, n20390, n20391, n20392,
         n20393, n20394, n20395, n20396, n20397, n20398, n20399, n20400,
         n20401, n20402, n20403, n20404, n20405, n20406, n20407, n20408,
         n20409, n20410, n20411, n20412, n20413, n20414, n20415, n20416,
         n20417, n20418, n20419, n20420, n20421, n20422, n20423, n20424,
         n20425, n20426, n20427, n20428, n20429, n20430, n20431, n20432,
         n20433, n20434, n20435, n20436, n20437, n20438, n20439, n20440,
         n20441, n20442, n20443, n20444, n20445, n20446, n20447, n20448,
         n20449, n20450, n20451, n20452, n20453, n20454, n20455, n20456,
         n20457, n20458, n20459, n20460, n20461, n20462, n20463, n20464,
         n20465, n20466, n20467, n20468, n20469, n20470, n20471, n20472,
         n20473, n20474, n20475, n20476, n20477, n20478, n20479, n20480,
         n20481, n20482, n20483, n20484, n20485, n20486, n20487, n20488,
         n20489, n20490, n20491, n20492, n20493, n20494, n20495, n20496,
         n20497, n20498, n20499, n20500, n20501, n20502, n20503, n20504,
         n20505, n20506, n20507, n20508, n20509, n20510, n20511, n20512,
         n20513, n20514, n20515, n20516, n20517, n20518, n20519, n20520,
         n20521, n20522, n20523, n20524, n20525, n20526, n20527, n20528,
         n20529, n20530, n20531, n20532, n20533, n20534, n20535, n20536,
         n20537, n20538, n20539, n20540, n20541, n20542, n20543, n20544,
         n20545, n20546, n20547, n20548, n20549, n20550, n20551, n20552,
         n20553, n20554, n20555, n20556, n20557, n20558, n20559, n20560,
         n20561, n20562, n20563, n20564, n20565, n20566, n20567, n20568,
         n20569, n20570, n20571, n20572, n20573, n20574, n20575, n20576,
         n20577, n20578, n20579, n20580, n20581, n20582, n20583, n20584,
         n20585, n20586, n20587, n20588, n20589, n20591, n20592, n20593,
         n20594, n20595, n20596, n20597, n20598, n20599, n20600, n20601,
         n20602, n20603, n20604, n20605, n20606, n20607, n20608, n20609,
         n20610, n20611, n20612, n20613, n20614, n20615, n20616, n20617,
         n20618, n20619, n20620, n20621, n20622, n20623, n20624, n20625,
         n20626, n20627, n20628, n20629, n20630, n20631, n20632, n20633,
         n20634, n20635, n20636, n20637, n20638, n20639, n20640, n20641,
         n20642, n20643, n20644, n20645, n20646, n20647, n20648, n20649,
         n20650, n20651, n20652, n20653, n20654, n20655, n20656, n20657,
         n20658, n20659, n20660, n20661, n20662, n20663, n20664, n20665,
         n20666, n20667, n20668, n20669, n20670, n20671, n20672, n20673,
         n20674, n20675, n20676, n20677, n20678, n20679, n20680, n20681,
         n20682, n20683, n20684, n20685, n20686, n20687, n20688, n20689,
         n20690, n20691, n20692, n20693, n20694, n20695, n20696, n20697,
         n20698, n20699, n20700, n20701, n20702, n20703, n20704, n20705,
         n20706, n20707, n20708, n20709, n20710, n20711, n20712, n20713,
         n20714, n20715, n20716, n20717, n20718, n20719, n20720, n20721,
         n20722, n20723, n20724, n20725, n20726, n20727, n20728, n20729,
         n20730, n20731, n20732, n20733, n20734, n20735, n20736, n20737,
         n20738, n20739, n20740, n20741, n20742, n20743, n20744, n20745,
         n20746, n20747, n20748, n20749, n20750, n20751, n20752, n20753,
         n20754, n20755, n20756, n20757, n20758, n20759, n20760, n20761,
         n20762, n20763, n20764, n20765, n20766, n20767, n20768, n20769,
         n20770, n20771, n20772, n20773, n20774, n20775, n20776, n20777,
         n20778, n20779, n20780, n20781, n20782, n20783, n20784, n20785,
         n20786, n20787, n20788, n20789, n20790, n20791, n20792, n20793,
         n20794, n20795, n20796, n20797, n20798, n20799, n20800, n20801,
         n20802, n20803, n20804, n20805, n20806, n20807, n20808, n20809,
         n20810, n20811, n20812, n20813, n20814, n20815, n20816, n20817,
         n20818, n20819, n20820, n20821, n20822, n20823, n20824, n20825,
         n20826, n20827, n20828, n20829, n20830, n20831, n20832, n20833,
         n20834, n20835, n20836, n20837, n20838, n20839, n20840, n20841,
         n20842, n20843, n20844, n20845, n20846, n20847, n20848, n20849,
         n20850, n20851, n20852, n20853, n20854, n20855, n20856, n20857,
         n20858, n20859, n20860, n20861, n20862, n20863, n20864, n20865,
         n20866, n20867, n20868, n20869, n20870, n20871, n20872, n20873,
         n20874, n20875, n20876, n20877, n20878, n20879, n20880, n20881,
         n20882, n20883, n20884, n20885, n20886, n20887, n20888, n20889,
         n20890, n20891, n20892, n20893, n20894, n20895, n20896, n20897,
         n20898, n20899, n20900, n20901, n20902, n20903, n20904, n20905,
         n20906, n20907, n20908, n20909, n20910, n20911, n20912, n20913,
         n20914, n20915, n20916, n20917, n20918, n20919, n20920, n20921,
         n20922, n20923, n20924, n20925, n20926, n20927, n20928, n20929,
         n20930, n20931, n20932, n20933, n20934, n20935, n20936, n20937,
         n20938, n20939, n20940, n20941, n20942, n20943, n20944, n20945,
         n20946, n20947, n20948, n20949, n20950, n20951, n20952, n20953,
         n20954, n20955, n20956, n20957, n20958, n20959, n20960, n20961,
         n20962, n20963, n20964, n20965, n20966, n20967, n20968, n20969,
         n20970, n20971, n20972, n20973, n20974, n20975, n20976, n20977,
         n20978, n20979, n20980, n20981, n20982, n20983, n20984, n20985,
         n20986, n20987, n20988, n20989, n20990, n20991, n20992, n20993,
         n20994, n20995, n20996, n20997, n20998, n20999, n21000, n21001,
         n21002, n21003, n21004, n21005, n21006, n21007, n21008, n21009,
         n21010, n21011, n21012, n21013, n21014, n21015, n21016, n21017,
         n21018, n21019, n21020, n21021, n21022, n21023, n21024, n21025,
         n21026, n21027, n21028, n21029, n21030, n21031, n21032, n21033,
         n21034, n21035, n21036, n21037, n21038, n21039, n21040, n21041,
         n21042, n21043, n21044, n21045, n21046, n21047, n21048, n21049,
         n21050, n21051, n21052, n21053, n21054, n21055, n21056, n21057,
         n21058, n21059, n21060, n21061, n21062, n21063, n21064, n21065,
         n21066, n21067, n21068, n21069, n21070, n21071, n21072, n21073,
         n21074, n21075, n21076, n21077, n21078, n21079, n21080, n21081,
         n21082, n21083, n21084, n21085, n21086, n21087, n21088, n21089,
         n21090, n21091, n21092, n21093, n21094, n21095, n21096, n21097,
         n21098, n21099, n21100, n21101, n21102, n21103, n21104, n21105,
         n21106, n21107, n21108, n21109, n21110, n21111, n21112, n21113,
         n21114, n21115, n21116, n21117, n21118, n21119, n21120, n21121,
         n21122, n21123, n21124, n21125, n21126, n21127, n21128, n21129,
         n21130, n21131, n21132, n21133, n21134, n21135, n21136, n21137,
         n21138, n21139, n21140, n21141, n21142, n21143, n21144, n21145,
         n21146, n21147, n21148, n21149, n21150, n21151, n21152, n21153,
         n21154, n21155, n21156, n21157, n21158, n21159, n21160, n21161,
         n21162, n21163, n21164, n21165, n21166, n21167, n21168, n21169,
         n21170, n21171, n21172, n21173, n21174, n21175, n21176, n21177,
         n21178, n21179, n21180, n21181, n21182, n21183, n21184, n21185,
         n21186, n21187, n21188, n21189, n21190, n21191, n21192, n21193,
         n21194, n21195, n21196, n21197, n21198, n21199, n21200, n21201,
         n21202, n21203, n21204, n21205, n21206, n21207, n21208, n21209,
         n21210, n21211, n21212, n21213, n21214, n21215, n21216, n21217,
         n21218, n21219, n21220, n21221, n21222, n21223, n21224, n21225,
         n21226, n21227, n21228, n21229, n21230, n21231, n21232, n21233,
         n21234, n21235, n21236, n21237, n21238, n21239, n21240, n21241,
         n21242, n21243, n21244, n21245, n21246, n21247, n21248, n21249,
         n21250, n21251, n21252, n21253, n21254, n21255, n21256, n21257,
         n21258, n21259, n21260, n21261, n21262, n21263, n21264, n21265,
         n21266, n21267, n21268, n21269, n21270, n21271, n21272, n21273,
         n21274, n21275, n21276, n21277, n21278, n21279, n21280, n21281,
         n21282, n21283, n21284, n21285, n21286, n21287, n21288, n21289,
         n21290, n21291, n21292, n21293, n21294, n21295, n21296, n21297;

  NOR2_X1 U11154 ( .A1(n19040), .A2(n9752), .ZN(n12760) );
  CLKBUF_X1 U11155 ( .A(n10469), .Z(n9759) );
  OR2_X1 U11156 ( .A1(n10418), .A2(n10421), .ZN(n10616) );
  OR2_X1 U11157 ( .A1(n10418), .A2(n10436), .ZN(n10620) );
  OR2_X1 U11158 ( .A1(n10418), .A2(n10425), .ZN(n20367) );
  OR3_X2 U11159 ( .A1(n13412), .A2(n15873), .A3(n10436), .ZN(n20300) );
  INV_X1 U11160 ( .A(n18053), .ZN(n19061) );
  NOR2_X1 U11161 ( .A1(n18676), .A2(n18682), .ZN(n18675) );
  CLKBUF_X1 U11162 ( .A(n12866), .Z(n12867) );
  INV_X1 U11163 ( .A(n14919), .ZN(n14957) );
  CLKBUF_X2 U11164 ( .A(n12684), .Z(n18002) );
  AND2_X1 U11165 ( .A1(n14989), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10507) );
  AND2_X1 U11166 ( .A1(n14932), .A2(n10461), .ZN(n10499) );
  AND2_X1 U11167 ( .A1(n14932), .A2(n13748), .ZN(n14885) );
  AND2_X1 U11168 ( .A1(n10317), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14910) );
  CLKBUF_X2 U11169 ( .A(n14927), .Z(n9761) );
  NAND2_X1 U11170 ( .A1(n11736), .A2(n11996), .ZN(n13743) );
  CLKBUF_X2 U11171 ( .A(n11162), .Z(n9715) );
  CLKBUF_X2 U11172 ( .A(n12588), .Z(n12539) );
  INV_X1 U11173 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n19656) );
  OR2_X1 U11174 ( .A1(n20755), .A2(n20750), .ZN(n11692) );
  NAND2_X2 U11175 ( .A1(n11127), .A2(n10226), .ZN(n13392) );
  INV_X1 U11176 ( .A(n13350), .ZN(n10336) );
  AND2_X1 U11177 ( .A1(n13305), .A2(n13599), .ZN(n11162) );
  AND2_X2 U11178 ( .A1(n10448), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n9739) );
  INV_X1 U11179 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13749) );
  AND2_X2 U11180 ( .A1(n13762), .A2(n14882), .ZN(n10317) );
  INV_X1 U11183 ( .A(n10894), .ZN(n10900) );
  OR2_X1 U11184 ( .A1(n16044), .A2(n16050), .ZN(n10827) );
  BUF_X1 U11185 ( .A(n10336), .Z(n13436) );
  BUF_X1 U11186 ( .A(n11238), .Z(n9749) );
  NAND2_X1 U11187 ( .A1(n9757), .A2(n10291), .ZN(n14473) );
  AND2_X1 U11188 ( .A1(n10440), .A2(n10441), .ZN(n9887) );
  INV_X1 U11190 ( .A(n14917), .ZN(n14956) );
  CLKBUF_X3 U11191 ( .A(n11752), .Z(n9713) );
  OR2_X1 U11192 ( .A1(n11768), .A2(n11771), .ZN(n13327) );
  NAND2_X1 U11193 ( .A1(n10412), .A2(n10215), .ZN(n20514) );
  NAND2_X1 U11195 ( .A1(n12663), .A2(n19674), .ZN(n17610) );
  AND2_X1 U11196 ( .A1(n12192), .A2(n13624), .ZN(n13625) );
  NAND2_X1 U11197 ( .A1(n9736), .A2(n11192), .ZN(n13649) );
  OR2_X1 U11198 ( .A1(n10822), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n10825) );
  NOR2_X1 U11200 ( .A1(n15932), .A2(n15933), .ZN(n11981) );
  NAND2_X1 U11201 ( .A1(n11976), .A2(n11975), .ZN(n15932) );
  INV_X1 U11202 ( .A(n20755), .ZN(n10469) );
  BUF_X1 U11203 ( .A(n10608), .Z(n9763) );
  OR2_X1 U11204 ( .A1(n17610), .A2(n12675), .ZN(n17827) );
  OR2_X1 U11205 ( .A1(n19506), .A2(n12675), .ZN(n17983) );
  INV_X1 U11206 ( .A(n16622), .ZN(n20850) );
  AND2_X1 U11207 ( .A1(n16963), .A2(n16962), .ZN(n17028) );
  INV_X1 U11208 ( .A(n12755), .ZN(n19056) );
  INV_X2 U11209 ( .A(n12838), .ZN(n17971) );
  OR2_X1 U11210 ( .A1(n18167), .A2(n9862), .ZN(n18137) );
  NAND2_X1 U11211 ( .A1(n12923), .A2(n17103), .ZN(n12931) );
  INV_X1 U11212 ( .A(n20808), .ZN(n16617) );
  INV_X1 U11213 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n20333) );
  INV_X4 U11215 ( .A(n10201), .ZN(n17864) );
  NAND2_X2 U11216 ( .A1(n14754), .A2(n10809), .ZN(n14757) );
  AND2_X1 U11217 ( .A1(n11050), .A2(n15828), .ZN(n11322) );
  AND2_X4 U11218 ( .A1(n13746), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10315) );
  NOR2_X2 U11220 ( .A1(n10897), .A2(n10896), .ZN(n10906) );
  NAND2_X2 U11221 ( .A1(n9930), .A2(n9928), .ZN(n11314) );
  OAI21_X2 U11222 ( .B1(n11685), .B2(n11686), .A(n11687), .ZN(n10848) );
  NOR2_X2 U11223 ( .A1(n18664), .A2(n18663), .ZN(n18662) );
  AOI21_X2 U11224 ( .B1(n16523), .B2(n10221), .A(n19546), .ZN(n18049) );
  OR3_X1 U11225 ( .A1(n10435), .A2(n13420), .A3(n10436), .ZN(n10659) );
  OR2_X1 U11226 ( .A1(n10435), .A2(n19923), .ZN(n10433) );
  NOR2_X2 U11228 ( .A1(n15855), .A2(n15854), .ZN(n15856) );
  NOR2_X2 U11229 ( .A1(n10714), .A2(n9946), .ZN(n10727) );
  XNOR2_X2 U11230 ( .A(n11361), .B(n11341), .ZN(n13729) );
  NAND2_X2 U11231 ( .A1(n11340), .A2(n11339), .ZN(n11361) );
  XNOR2_X2 U11233 ( .A(n10702), .B(n14394), .ZN(n14381) );
  NOR4_X2 U11234 ( .A1(n18698), .A2(n18715), .A3(n18697), .A4(n18696), .ZN(
        n18708) );
  XNOR2_X2 U11235 ( .A(n10653), .B(n10926), .ZN(n14259) );
  NAND2_X2 U11236 ( .A1(n10652), .A2(n19903), .ZN(n10653) );
  AND2_X4 U11237 ( .A1(n9761), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14951) );
  AND2_X1 U11238 ( .A1(n11463), .A2(n16645), .ZN(n16648) );
  OR2_X1 U11239 ( .A1(n16119), .A2(n16185), .ZN(n16187) );
  NAND2_X1 U11240 ( .A1(n12446), .A2(n10175), .ZN(n15180) );
  OR2_X1 U11241 ( .A1(n18473), .A2(n18509), .ZN(n18433) );
  CLKBUF_X2 U11242 ( .A(n18560), .Z(n9716) );
  OR2_X1 U11243 ( .A1(n10420), .A2(n10436), .ZN(n20549) );
  INV_X1 U11244 ( .A(n10420), .ZN(n10412) );
  INV_X1 U11245 ( .A(n15888), .ZN(n13259) );
  CLKBUF_X2 U11246 ( .A(n14197), .Z(n9719) );
  AOI21_X1 U11247 ( .B1(n10392), .B2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A(
        n10381), .ZN(n10386) );
  OAI21_X1 U11248 ( .B1(n12770), .B2(n16452), .A(n19477), .ZN(n19505) );
  NOR2_X1 U11249 ( .A1(n18272), .A2(n12757), .ZN(n19477) );
  INV_X1 U11250 ( .A(n10925), .ZN(n11019) );
  AND2_X1 U11251 ( .A1(n11197), .A2(n9950), .ZN(n9949) );
  INV_X1 U11252 ( .A(n11500), .ZN(n11510) );
  NAND2_X1 U11254 ( .A1(n18053), .A2(n12755), .ZN(n12946) );
  NAND3_X1 U11255 ( .A1(n12827), .A2(n12826), .A3(n10204), .ZN(n18683) );
  NAND2_X1 U11256 ( .A1(n10273), .A2(n10272), .ZN(n20098) );
  INV_X4 U11257 ( .A(n12705), .ZN(n12899) );
  INV_X4 U11258 ( .A(n17913), .ZN(n17970) );
  INV_X4 U11259 ( .A(n17975), .ZN(n12840) );
  BUF_X2 U11260 ( .A(n11158), .Z(n9762) );
  BUF_X2 U11261 ( .A(n11385), .Z(n12603) );
  CLKBUF_X2 U11262 ( .A(n11223), .Z(n12604) );
  INV_X1 U11263 ( .A(n12833), .ZN(n17946) );
  BUF_X2 U11265 ( .A(n11153), .Z(n12413) );
  NOR2_X1 U11266 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n20699) );
  INV_X1 U11267 ( .A(n12831), .ZN(n12726) );
  NOR2_X1 U11268 ( .A1(n12675), .A2(n12674), .ZN(n12833) );
  INV_X4 U11269 ( .A(n17966), .ZN(n17948) );
  INV_X4 U11270 ( .A(n12829), .ZN(n9714) );
  INV_X2 U11271 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11043) );
  INV_X2 U11272 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11262) );
  NOR2_X1 U11273 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n14932) );
  INV_X2 U11274 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10230) );
  OR2_X1 U11275 ( .A1(n15619), .A2(n16792), .ZN(n9994) );
  XNOR2_X1 U11276 ( .A(n11467), .B(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14760) );
  AND2_X1 U11277 ( .A1(n12029), .A2(n9789), .ZN(n10072) );
  AOI21_X1 U11278 ( .B1(n12053), .B2(n17010), .A(n9966), .ZN(n11042) );
  OAI22_X1 U11279 ( .A1(n16646), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .B1(
        n16648), .B2(n11464), .ZN(n15620) );
  AND2_X1 U11280 ( .A1(n10153), .A2(n10152), .ZN(n16104) );
  XNOR2_X1 U11281 ( .A(n14800), .B(n13034), .ZN(n14801) );
  XNOR2_X1 U11282 ( .A(n9967), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n12053) );
  OR2_X1 U11283 ( .A1(n9801), .A2(n16656), .ZN(n16755) );
  NAND2_X1 U11284 ( .A1(n16033), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n9967) );
  NOR2_X1 U11285 ( .A1(n16034), .A2(n16206), .ZN(n16033) );
  NAND2_X1 U11286 ( .A1(n9792), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n16034) );
  OR2_X1 U11287 ( .A1(n16053), .A2(n10192), .ZN(n16045) );
  XNOR2_X1 U11288 ( .A(n12634), .B(n12633), .ZN(n15148) );
  AOI21_X1 U11289 ( .B1(n17094), .B2(n17095), .A(n9900), .ZN(n17148) );
  AOI211_X1 U11290 ( .C1(n17131), .C2(n18596), .A(n17130), .B(n17129), .ZN(
        n17135) );
  AOI21_X1 U11291 ( .B1(n18335), .B2(n18334), .A(n18333), .ZN(n18340) );
  NAND2_X1 U11292 ( .A1(n14757), .A2(n10812), .ZN(n16060) );
  OR2_X1 U11293 ( .A1(n15906), .A2(n15905), .ZN(n10055) );
  AOI21_X1 U11294 ( .B1(n16351), .B2(n16349), .A(n16090), .ZN(n16944) );
  AND2_X1 U11295 ( .A1(n16400), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n16987) );
  AND2_X1 U11296 ( .A1(n12534), .A2(n9825), .ZN(n14734) );
  AOI21_X1 U11297 ( .B1(n12941), .B2(n12940), .A(n17160), .ZN(n12942) );
  OR2_X1 U11298 ( .A1(n10223), .A2(n15582), .ZN(n16591) );
  OR2_X1 U11299 ( .A1(n15520), .A2(n15430), .ZN(n15518) );
  NOR2_X1 U11300 ( .A1(n16508), .A2(n10210), .ZN(n17090) );
  NOR2_X1 U11301 ( .A1(n15914), .A2(n15913), .ZN(n15912) );
  NOR2_X1 U11302 ( .A1(n17159), .A2(n12931), .ZN(n17151) );
  NAND2_X1 U11303 ( .A1(n9908), .A2(n10095), .ZN(n16508) );
  OR2_X1 U11304 ( .A1(n10178), .A2(n15530), .ZN(n15520) );
  AND2_X1 U11305 ( .A1(n9957), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n9931) );
  NAND2_X1 U11306 ( .A1(n18352), .A2(n10094), .ZN(n17159) );
  NAND2_X1 U11307 ( .A1(n9921), .A2(n9919), .ZN(n14645) );
  NAND2_X1 U11308 ( .A1(n16848), .A2(n16849), .ZN(n16847) );
  AND2_X1 U11309 ( .A1(n12939), .A2(n9782), .ZN(n10094) );
  NAND2_X1 U11310 ( .A1(n9909), .A2(n12936), .ZN(n18352) );
  OR2_X1 U11311 ( .A1(n10115), .A2(n16673), .ZN(n9957) );
  NAND2_X1 U11312 ( .A1(n9774), .A2(n10905), .ZN(n10185) );
  AOI21_X1 U11313 ( .B1(n10118), .B2(n10116), .A(n9849), .ZN(n10115) );
  AND2_X1 U11314 ( .A1(n11981), .A2(n11980), .ZN(n12041) );
  NOR2_X1 U11315 ( .A1(n14808), .A2(n14809), .ZN(n15894) );
  OR2_X1 U11316 ( .A1(n14560), .A2(n14561), .ZN(n14563) );
  AND2_X1 U11317 ( .A1(n10904), .A2(n14394), .ZN(n10905) );
  NAND2_X1 U11318 ( .A1(n15920), .A2(n9786), .ZN(n16914) );
  XNOR2_X1 U11319 ( .A(n14820), .B(n14819), .ZN(n15467) );
  XNOR2_X1 U11320 ( .A(n10130), .B(n14816), .ZN(n15160) );
  NOR2_X1 U11321 ( .A1(n19014), .A2(n18769), .ZN(n18817) );
  NOR2_X1 U11322 ( .A1(n15746), .A2(n11450), .ZN(n9959) );
  INV_X1 U11323 ( .A(n12133), .ZN(n10130) );
  INV_X1 U11324 ( .A(n14799), .ZN(n13034) );
  AOI21_X1 U11325 ( .B1(n9924), .B2(n13833), .A(n9793), .ZN(n9923) );
  OR2_X1 U11326 ( .A1(n16198), .A2(n10936), .ZN(n9774) );
  NAND2_X1 U11327 ( .A1(n10891), .A2(n10890), .ZN(n14263) );
  NOR2_X1 U11328 ( .A1(n12130), .A2(n13064), .ZN(n13063) );
  OR2_X1 U11329 ( .A1(n15997), .A2(n15929), .ZN(n15927) );
  AND2_X1 U11330 ( .A1(n18418), .A2(n18433), .ZN(n18465) );
  AOI21_X1 U11331 ( .B1(n9922), .B2(n16728), .A(n9920), .ZN(n9919) );
  AND2_X1 U11332 ( .A1(n15747), .A2(n11456), .ZN(n11457) );
  AND2_X1 U11333 ( .A1(n9818), .A2(n16729), .ZN(n9922) );
  OR2_X1 U11334 ( .A1(n18735), .A2(n12933), .ZN(n10099) );
  NOR2_X1 U11335 ( .A1(n15664), .A2(n16687), .ZN(n15747) );
  NAND2_X1 U11336 ( .A1(n10893), .A2(n10926), .ZN(n14260) );
  NOR2_X1 U11337 ( .A1(n18474), .A2(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n18473) );
  OR2_X1 U11338 ( .A1(n15776), .A2(n15779), .ZN(n15664) );
  NAND2_X1 U11339 ( .A1(n12993), .A2(n18592), .ZN(n18512) );
  NOR2_X1 U11340 ( .A1(n14128), .A2(n16137), .ZN(n14435) );
  INV_X1 U11341 ( .A(n15988), .ZN(n10075) );
  NAND2_X1 U11342 ( .A1(n18757), .A2(n18800), .ZN(n18418) );
  INV_X1 U11343 ( .A(n11455), .ZN(n16687) );
  INV_X1 U11344 ( .A(n19963), .ZN(n13637) );
  OR2_X1 U11345 ( .A1(n11408), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n16737) );
  AND2_X1 U11346 ( .A1(n16581), .A2(n10138), .ZN(n15496) );
  AND2_X1 U11347 ( .A1(n18088), .A2(P3_EAX_REG_24__SCAN_IN), .ZN(n18083) );
  NAND2_X1 U11348 ( .A1(n13696), .A2(n13443), .ZN(n19963) );
  AND2_X1 U11349 ( .A1(n16692), .A2(n11448), .ZN(n16689) );
  AND2_X1 U11350 ( .A1(n15759), .A2(n11447), .ZN(n11455) );
  OAI211_X1 U11351 ( .C1(n12208), .C2(n12300), .A(n12207), .B(n12206), .ZN(
        n13818) );
  NAND2_X1 U11352 ( .A1(n11426), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n14352) );
  INV_X1 U11353 ( .A(n18833), .ZN(n18757) );
  OAI21_X1 U11354 ( .B1(n18510), .B2(n18836), .A(n12931), .ZN(n18479) );
  NOR2_X1 U11355 ( .A1(n10825), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n9936) );
  NAND2_X1 U11356 ( .A1(n17112), .A2(n18816), .ZN(n18833) );
  NAND2_X1 U11357 ( .A1(n11378), .A2(n9971), .ZN(n12208) );
  OR2_X1 U11358 ( .A1(n16673), .A2(n11425), .ZN(n11426) );
  NAND2_X1 U11359 ( .A1(n11316), .A2(n11315), .ZN(n11338) );
  AND2_X1 U11360 ( .A1(n13698), .A2(n13697), .ZN(n13696) );
  OAI21_X1 U11361 ( .B1(n15813), .B2(n12300), .A(n12191), .ZN(n13624) );
  AND2_X1 U11362 ( .A1(n11411), .A2(n11494), .ZN(n11444) );
  NAND2_X1 U11363 ( .A1(n9973), .A2(n9972), .ZN(n9971) );
  OR2_X1 U11364 ( .A1(n11400), .A2(n11399), .ZN(n12209) );
  XNOR2_X1 U11365 ( .A(n11411), .B(n11410), .ZN(n12143) );
  NOR2_X1 U11366 ( .A1(n12988), .A2(n18946), .ZN(n12989) );
  OR2_X1 U11367 ( .A1(n11336), .A2(n11364), .ZN(n15813) );
  NAND2_X1 U11368 ( .A1(n10804), .A2(n10824), .ZN(n10802) );
  OR2_X1 U11369 ( .A1(n10782), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n10804) );
  NOR2_X1 U11370 ( .A1(n18603), .A2(n18946), .ZN(n18602) );
  NAND2_X1 U11371 ( .A1(n10412), .A2(n10422), .ZN(n13810) );
  AOI211_X1 U11372 ( .C1(n9763), .C2(n20333), .A(n20291), .B(n20699), .ZN(
        n13962) );
  NAND2_X1 U11373 ( .A1(n10419), .A2(n10215), .ZN(n20404) );
  OAI22_X1 U11374 ( .A1(n14157), .A2(n20549), .B1(n10616), .B2(n14991), .ZN(
        n10482) );
  NOR2_X2 U11375 ( .A1(n19660), .A2(n18677), .ZN(n18547) );
  NOR2_X1 U11376 ( .A1(n10770), .A2(n10750), .ZN(n10781) );
  NAND2_X1 U11377 ( .A1(n10427), .A2(n10426), .ZN(n20129) );
  CLKBUF_X1 U11378 ( .A(n14705), .Z(n15598) );
  CLKBUF_X1 U11379 ( .A(n14707), .Z(n15596) );
  NAND2_X1 U11380 ( .A1(n12175), .A2(n12178), .ZN(n15812) );
  NAND2_X1 U11381 ( .A1(n10754), .A2(n10741), .ZN(n10770) );
  AND2_X1 U11382 ( .A1(n10736), .A2(n9944), .ZN(n10754) );
  NOR2_X1 U11383 ( .A1(n14233), .A2(n14095), .ZN(n21165) );
  NOR2_X1 U11384 ( .A1(n13888), .A2(n14095), .ZN(n21128) );
  NOR2_X1 U11385 ( .A1(n13980), .A2(n14095), .ZN(n21158) );
  NOR2_X1 U11386 ( .A1(n13881), .A2(n14095), .ZN(n21134) );
  NOR2_X1 U11387 ( .A1(n13863), .A2(n14095), .ZN(n21114) );
  NOR2_X1 U11388 ( .A1(n13871), .A2(n14095), .ZN(n21140) );
  NOR2_X1 U11389 ( .A1(n13972), .A2(n14095), .ZN(n21146) );
  NOR2_X1 U11390 ( .A1(n13876), .A2(n14095), .ZN(n21152) );
  NOR2_X2 U11391 ( .A1(n20921), .A2(n13951), .ZN(n13652) );
  NOR2_X1 U11392 ( .A1(n18628), .A2(n18629), .ZN(n18627) );
  AND2_X1 U11393 ( .A1(n17942), .A2(P3_EBX_REG_11__SCAN_IN), .ZN(n17910) );
  INV_X2 U11394 ( .A(n13695), .ZN(n9717) );
  NAND2_X2 U11395 ( .A1(n15603), .A2(n13394), .ZN(n15610) );
  AND2_X1 U11396 ( .A1(n10730), .A2(n10731), .ZN(n10736) );
  AND2_X1 U11397 ( .A1(n14265), .A2(n11787), .ZN(n13401) );
  OR2_X1 U11398 ( .A1(n11250), .A2(n11249), .ZN(n11260) );
  OR2_X1 U11399 ( .A1(n11275), .A2(n11274), .ZN(n11276) );
  XNOR2_X1 U11400 ( .A(n10093), .B(n10092), .ZN(n18628) );
  OAI21_X1 U11401 ( .B1(n9905), .B2(n18644), .A(n9903), .ZN(n10093) );
  NOR2_X1 U11402 ( .A1(n19715), .A2(n12785), .ZN(n17621) );
  NAND2_X1 U11403 ( .A1(n13527), .A2(n16486), .ZN(n20773) );
  NOR2_X2 U11404 ( .A1(n20092), .A2(n20551), .ZN(n20093) );
  NOR2_X2 U11405 ( .A1(n9759), .A2(n20120), .ZN(n20087) );
  NOR2_X2 U11406 ( .A1(n14301), .A2(n20551), .ZN(n13591) );
  NOR2_X2 U11407 ( .A1(n20088), .A2(n20551), .ZN(n20089) );
  NOR2_X1 U11408 ( .A1(n18948), .A2(n18995), .ZN(n19006) );
  OAI21_X1 U11409 ( .B1(n19493), .B2(n19505), .A(n19492), .ZN(n19515) );
  XNOR2_X1 U11410 ( .A(n10917), .B(n10916), .ZN(n10919) );
  XNOR2_X1 U11411 ( .A(n10386), .B(n10385), .ZN(n10397) );
  XNOR2_X1 U11412 ( .A(n11036), .B(n11038), .ZN(n12056) );
  AND2_X1 U11413 ( .A1(n10375), .A2(n10374), .ZN(n10399) );
  OR2_X1 U11414 ( .A1(n18652), .A2(n18976), .ZN(n9905) );
  OR2_X1 U11415 ( .A1(n9730), .A2(n12861), .ZN(n12863) );
  AOI21_X1 U11416 ( .B1(n10392), .B2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n10372), .ZN(n10398) );
  NAND2_X1 U11417 ( .A1(n10700), .A2(n10699), .ZN(n10707) );
  INV_X2 U11418 ( .A(n18315), .ZN(n18310) );
  AND2_X1 U11419 ( .A1(n16455), .A2(n16454), .ZN(n16522) );
  AOI21_X1 U11420 ( .B1(n10392), .B2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        n10395), .ZN(n10916) );
  AND2_X1 U11421 ( .A1(n10650), .A2(n10649), .ZN(n10700) );
  AND2_X1 U11422 ( .A1(n11206), .A2(n11205), .ZN(n11252) );
  AOI21_X1 U11423 ( .B1(n11188), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n11187), 
        .ZN(n11189) );
  AND2_X1 U11424 ( .A1(n10350), .A2(n10362), .ZN(n10360) );
  NOR2_X1 U11425 ( .A1(n10645), .A2(n10646), .ZN(n10650) );
  NAND2_X1 U11426 ( .A1(n10049), .A2(n13743), .ZN(n10048) );
  AND2_X1 U11427 ( .A1(n9879), .A2(n9878), .ZN(n10362) );
  AOI21_X1 U11428 ( .B1(n11204), .B2(n11203), .A(n11202), .ZN(n11205) );
  NAND2_X1 U11429 ( .A1(n12848), .A2(n12864), .ZN(n12849) );
  OR2_X1 U11430 ( .A1(n11760), .A2(n11761), .ZN(n11766) );
  NOR2_X1 U11431 ( .A1(n12767), .A2(n19044), .ZN(n17263) );
  NAND2_X1 U11432 ( .A1(n9881), .A2(n9880), .ZN(n10361) );
  AND2_X1 U11433 ( .A1(n11563), .A2(n11184), .ZN(n11206) );
  INV_X1 U11434 ( .A(n12864), .ZN(n12974) );
  NAND2_X1 U11435 ( .A1(n9895), .A2(n9891), .ZN(n12864) );
  INV_X2 U11436 ( .A(n10925), .ZN(n11026) );
  NAND2_X1 U11437 ( .A1(n13796), .A2(n10354), .ZN(n10931) );
  NAND2_X1 U11438 ( .A1(n9943), .A2(n9942), .ZN(n10579) );
  NAND2_X1 U11439 ( .A1(n19040), .A2(n9751), .ZN(n16521) );
  NOR2_X1 U11440 ( .A1(n10925), .A2(n10352), .ZN(n10358) );
  NAND2_X1 U11441 ( .A1(n11751), .A2(n11750), .ZN(n13372) );
  AND2_X1 U11442 ( .A1(n11759), .A2(n11758), .ZN(n13263) );
  INV_X1 U11443 ( .A(n12847), .ZN(n9895) );
  AND2_X1 U11444 ( .A1(n13051), .A2(n11194), .ZN(n13299) );
  NAND3_X1 U11445 ( .A1(n9951), .A2(n9949), .A3(n9948), .ZN(n11182) );
  CLKBUF_X1 U11446 ( .A(n10861), .Z(n13737) );
  AND2_X1 U11447 ( .A1(n11992), .A2(n9882), .ZN(n10343) );
  INV_X1 U11448 ( .A(n19700), .ZN(n9751) );
  INV_X1 U11449 ( .A(n10363), .ZN(n10354) );
  INV_X2 U11450 ( .A(n12128), .ZN(n12132) );
  AND3_X1 U11451 ( .A1(n9804), .A2(n12811), .A3(n9896), .ZN(n12847) );
  AND2_X1 U11452 ( .A1(n13369), .A2(n10469), .ZN(n11992) );
  OAI211_X1 U11453 ( .C1(n17913), .C2(n18014), .A(n12725), .B(n12724), .ZN(
        n18143) );
  AND2_X2 U11454 ( .A1(n14299), .A2(n11782), .ZN(n12037) );
  INV_X1 U11455 ( .A(n18191), .ZN(n9891) );
  AND2_X1 U11456 ( .A1(n10536), .A2(n10535), .ZN(n11762) );
  NAND2_X1 U11457 ( .A1(n11178), .A2(n13880), .ZN(n11198) );
  NOR2_X1 U11458 ( .A1(n11567), .A2(n11097), .ZN(n11132) );
  INV_X1 U11459 ( .A(n11195), .ZN(n12128) );
  NAND2_X1 U11460 ( .A1(n13880), .A2(n11554), .ZN(n11567) );
  AND2_X1 U11461 ( .A1(n9800), .A2(n9892), .ZN(n18191) );
  AOI211_X1 U11462 ( .C1(n12840), .C2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A(
        n12723), .B(n12722), .ZN(n12724) );
  AND2_X1 U11463 ( .A1(n10561), .A2(n13368), .ZN(n14299) );
  NAND4_X2 U11464 ( .A1(n11994), .A2(n13436), .A3(n10561), .A4(n20121), .ZN(
        n9882) );
  OAI211_X1 U11465 ( .C1(n17946), .C2(n17789), .A(n12704), .B(n12703), .ZN(
        n12755) );
  INV_X1 U11467 ( .A(n20098), .ZN(n11990) );
  NAND2_X1 U11468 ( .A1(n20750), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n20754) );
  NAND2_X1 U11469 ( .A1(n11068), .A2(n10202), .ZN(n11554) );
  NAND3_X2 U11470 ( .A1(n11174), .A2(n11173), .A3(n11172), .ZN(n11177) );
  OR2_X1 U11471 ( .A1(n11216), .A2(n11215), .ZN(n11423) );
  INV_X2 U11472 ( .A(n10306), .ZN(n10838) );
  OR2_X1 U11473 ( .A1(n11229), .A2(n11228), .ZN(n11309) );
  INV_X1 U11474 ( .A(n11192), .ZN(n13936) );
  AND4_X1 U11475 ( .A1(n11111), .A2(n11110), .A3(n11109), .A4(n11108), .ZN(
        n11127) );
  AND3_X1 U11476 ( .A1(n12825), .A2(n12824), .A3(n12823), .ZN(n10204) );
  AND3_X1 U11477 ( .A1(n11126), .A2(n11125), .A3(n11124), .ZN(n10226) );
  AND2_X1 U11478 ( .A1(n11161), .A2(n11160), .ZN(n11174) );
  NAND2_X2 U11479 ( .A1(n10225), .A2(n9787), .ZN(n14704) );
  NAND4_X2 U11480 ( .A1(n11096), .A2(n11095), .A3(n11094), .A4(n11093), .ZN(
        n11677) );
  OR3_X1 U11481 ( .A1(n12837), .A2(n12845), .A3(n9894), .ZN(n9893) );
  INV_X1 U11482 ( .A(n11994), .ZN(n10335) );
  AND4_X1 U11483 ( .A1(n11144), .A2(n11143), .A3(n11142), .A4(n11141), .ZN(
        n11150) );
  NAND2_X1 U11484 ( .A1(n10248), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10249) );
  AND4_X1 U11485 ( .A1(n11088), .A2(n11087), .A3(n11086), .A4(n11085), .ZN(
        n11094) );
  AND4_X1 U11486 ( .A1(n11136), .A2(n11135), .A3(n11134), .A4(n11133), .ZN(
        n11152) );
  AND4_X1 U11487 ( .A1(n11092), .A2(n11091), .A3(n11090), .A4(n11089), .ZN(
        n11093) );
  NAND2_X1 U11488 ( .A1(n10271), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10272) );
  AND4_X1 U11489 ( .A1(n11072), .A2(n11071), .A3(n11070), .A4(n11069), .ZN(
        n10225) );
  AND4_X1 U11490 ( .A1(n11157), .A2(n11156), .A3(n11155), .A4(n11154), .ZN(
        n11161) );
  AND4_X1 U11491 ( .A1(n11148), .A2(n11147), .A3(n11146), .A4(n11145), .ZN(
        n11149) );
  NAND2_X1 U11492 ( .A1(n10259), .A2(n10208), .ZN(n10260) );
  NAND2_X1 U11493 ( .A1(n9962), .A2(n9960), .ZN(n11994) );
  AND4_X1 U11494 ( .A1(n11073), .A2(n11075), .A3(n11074), .A4(n11076), .ZN(
        n9787) );
  AND4_X1 U11495 ( .A1(n11102), .A2(n11101), .A3(n11100), .A4(n11099), .ZN(
        n11107) );
  AND4_X1 U11496 ( .A1(n11115), .A2(n11114), .A3(n11113), .A4(n11112), .ZN(
        n11126) );
  AND4_X1 U11497 ( .A1(n11119), .A2(n11118), .A3(n11117), .A4(n11116), .ZN(
        n11125) );
  AND4_X1 U11498 ( .A1(n11080), .A2(n11079), .A3(n11078), .A4(n11077), .ZN(
        n11096) );
  AND4_X1 U11499 ( .A1(n11048), .A2(n11047), .A3(n11046), .A4(n11045), .ZN(
        n11057) );
  AND4_X1 U11500 ( .A1(n11106), .A2(n11105), .A3(n11104), .A4(n11103), .ZN(
        n10227) );
  INV_X2 U11501 ( .A(U214), .ZN(n17216) );
  INV_X2 U11502 ( .A(n17946), .ZN(n17967) );
  INV_X1 U11503 ( .A(n12882), .ZN(n12705) );
  AND3_X1 U11504 ( .A1(n10256), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        n10255), .ZN(n10259) );
  AND2_X2 U11505 ( .A1(n15129), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10631) );
  AND4_X1 U11506 ( .A1(n10270), .A2(n10269), .A3(n10268), .A4(n10267), .ZN(
        n10271) );
  NAND4_X1 U11507 ( .A1(n9961), .A2(n10235), .A3(n10236), .A4(n10238), .ZN(
        n9960) );
  AND4_X1 U11508 ( .A1(n11084), .A2(n11083), .A3(n11082), .A4(n11081), .ZN(
        n11095) );
  AND4_X1 U11509 ( .A1(n11123), .A2(n11122), .A3(n11121), .A4(n11120), .ZN(
        n11124) );
  AND4_X1 U11510 ( .A1(n11140), .A2(n11139), .A3(n11138), .A4(n11137), .ZN(
        n11151) );
  AND4_X1 U11511 ( .A1(n9978), .A2(n9977), .A3(n9976), .A4(n9975), .ZN(n11160)
         );
  NAND2_X2 U11512 ( .A1(n19710), .A2(n19578), .ZN(n19636) );
  INV_X2 U11513 ( .A(n17253), .ZN(U215) );
  NAND2_X2 U11514 ( .A1(n19710), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n19640) );
  CLKBUF_X3 U11515 ( .A(n11322), .Z(n9756) );
  INV_X2 U11516 ( .A(n13597), .ZN(n11098) );
  CLKBUF_X2 U11517 ( .A(n11322), .Z(n9755) );
  CLKBUF_X2 U11518 ( .A(n11238), .Z(n9750) );
  INV_X1 U11519 ( .A(n17983), .ZN(n17992) );
  BUF_X2 U11520 ( .A(n12612), .Z(n9745) );
  NAND2_X2 U11521 ( .A1(n12666), .A2(n19656), .ZN(n17975) );
  AND2_X1 U11522 ( .A1(n10290), .A2(n10291), .ZN(n9866) );
  NAND2_X1 U11523 ( .A1(n12662), .A2(n12661), .ZN(n12838) );
  INV_X2 U11524 ( .A(n12684), .ZN(n17958) );
  AND2_X1 U11525 ( .A1(n10286), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9868) );
  AND3_X1 U11526 ( .A1(n10280), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        n10279), .ZN(n10283) );
  AND2_X1 U11527 ( .A1(n10262), .A2(n10291), .ZN(n10266) );
  OR2_X2 U11528 ( .A1(n12636), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n16823) );
  OR3_X2 U11529 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(n12674), .ZN(n12829) );
  INV_X2 U11530 ( .A(n17258), .ZN(n17260) );
  BUF_X2 U11531 ( .A(n10315), .Z(n13745) );
  AND2_X1 U11532 ( .A1(n10316), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n10309) );
  AND2_X2 U11533 ( .A1(n10448), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10444) );
  NAND2_X2 U11534 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n19497), .ZN(
        n17995) );
  AND2_X2 U11535 ( .A1(n11051), .A2(n11052), .ZN(n11385) );
  AND2_X2 U11536 ( .A1(n10460), .A2(n14932), .ZN(n10498) );
  BUF_X2 U11537 ( .A(n11163), .Z(n9737) );
  AND3_X1 U11538 ( .A1(n10216), .A2(n11460), .A3(n11641), .ZN(n9723) );
  AND2_X2 U11539 ( .A1(n15828), .A2(n11044), .ZN(n11238) );
  AND2_X1 U11540 ( .A1(n14745), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11049) );
  AND2_X1 U11541 ( .A1(n11262), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11051) );
  AND2_X2 U11542 ( .A1(n13316), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13599) );
  AND2_X2 U11543 ( .A1(n11262), .A2(n10100), .ZN(n15828) );
  OR3_X2 U11544 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(n19506), .ZN(n17966) );
  AND2_X4 U11545 ( .A1(n13305), .A2(n11052), .ZN(n11163) );
  NAND2_X1 U11546 ( .A1(n19666), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12675) );
  NAND3_X1 U11547 ( .A1(n19674), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n12676) );
  NOR2_X2 U11548 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11044) );
  AND2_X1 U11549 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13748) );
  INV_X2 U11550 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13316) );
  NOR2_X1 U11551 ( .A1(n17103), .A2(n18687), .ZN(n18560) );
  INV_X1 U11552 ( .A(n11738), .ZN(n9721) );
  AND2_X1 U11553 ( .A1(n12098), .A2(n11712), .ZN(n9725) );
  INV_X1 U11554 ( .A(n9725), .ZN(n11738) );
  NAND2_X1 U11555 ( .A1(n9915), .A2(n9913), .ZN(n9722) );
  NAND2_X1 U11556 ( .A1(n11461), .A2(n9723), .ZN(n11462) );
  CLKBUF_X1 U11557 ( .A(n11197), .Z(n9724) );
  NAND2_X1 U11558 ( .A1(n9915), .A2(n9913), .ZN(n13060) );
  OAI22_X1 U11559 ( .A1(n13401), .A2(n13400), .B1(n11790), .B2(n11953), .ZN(
        n13399) );
  NOR2_X2 U11560 ( .A1(n13701), .A2(n13702), .ZN(n13703) );
  AOI211_X2 U11561 ( .C1(n16216), .C2(n17052), .A(n16215), .B(n16214), .ZN(
        n16217) );
  NOR2_X4 U11562 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13762) );
  NOR2_X1 U11563 ( .A1(n18627), .A2(n9729), .ZN(n9726) );
  NOR2_X1 U11564 ( .A1(n9726), .A2(n9727), .ZN(n9907) );
  AND2_X1 U11565 ( .A1(n9728), .A2(n18613), .ZN(n9727) );
  INV_X1 U11566 ( .A(n12911), .ZN(n9728) );
  OR2_X1 U11567 ( .A1(n12897), .A2(n12911), .ZN(n9729) );
  NOR2_X1 U11568 ( .A1(n18662), .A2(n12850), .ZN(n9730) );
  INV_X1 U11569 ( .A(n9909), .ZN(n9731) );
  AND2_X1 U11570 ( .A1(n10402), .A2(n10407), .ZN(n19923) );
  AOI22_X1 U11571 ( .A1(n18674), .A2(n18512), .B1(n18560), .B2(n17112), .ZN(
        n18586) );
  AND2_X1 U11572 ( .A1(n13350), .A2(n10306), .ZN(n13374) );
  XNOR2_X2 U11574 ( .A(n10656), .B(n10657), .ZN(n10892) );
  CLKBUF_X1 U11575 ( .A(n16727), .Z(n9732) );
  CLKBUF_X1 U11576 ( .A(n13553), .Z(n9733) );
  NAND2_X1 U11577 ( .A1(n13294), .A2(n11276), .ZN(n9734) );
  XNOR2_X1 U11578 ( .A(n11338), .B(n11317), .ZN(n13553) );
  NAND2_X1 U11579 ( .A1(n13294), .A2(n11276), .ZN(n13298) );
  NOR2_X1 U11580 ( .A1(n11291), .A2(n11290), .ZN(n11294) );
  NOR2_X1 U11581 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n12676), .ZN(
        n9735) );
  INV_X1 U11582 ( .A(n11177), .ZN(n9736) );
  INV_X2 U11583 ( .A(n11177), .ZN(n13951) );
  NOR3_X2 U11584 ( .A1(n9751), .A2(n12755), .A3(n12995), .ZN(n18272) );
  NOR2_X1 U11585 ( .A1(n11182), .A2(n10207), .ZN(n11488) );
  XNOR2_X1 U11586 ( .A(n10878), .B(n11777), .ZN(n20034) );
  OR2_X1 U11587 ( .A1(n13393), .A2(n11185), .ZN(n15821) );
  OAI21_X2 U11588 ( .B1(n10894), .B2(n10826), .A(n19889), .ZN(n10702) );
  NAND2_X2 U11589 ( .A1(n10909), .A2(n10697), .ZN(n10894) );
  NAND2_X1 U11590 ( .A1(n13392), .A2(n13049), .ZN(n11179) );
  AND2_X1 U11591 ( .A1(n11050), .A2(n11049), .ZN(n9738) );
  AND2_X2 U11592 ( .A1(n11050), .A2(n11049), .ZN(n12395) );
  NOR2_X4 U11594 ( .A1(n13420), .A2(n10184), .ZN(n20162) );
  NAND2_X2 U11595 ( .A1(n11189), .A2(n11257), .ZN(n11268) );
  NAND2_X2 U11596 ( .A1(n11050), .A2(n13305), .ZN(n13597) );
  AND2_X4 U11597 ( .A1(n11044), .A2(n13305), .ZN(n9741) );
  NAND2_X1 U11598 ( .A1(n10412), .A2(n10415), .ZN(n20476) );
  AND2_X1 U11599 ( .A1(n13305), .A2(n13599), .ZN(n9742) );
  AND2_X1 U11600 ( .A1(n13305), .A2(n13599), .ZN(n9743) );
  AND2_X1 U11601 ( .A1(n11049), .A2(n11052), .ZN(n9744) );
  AND2_X2 U11602 ( .A1(n11049), .A2(n11052), .ZN(n12588) );
  BUF_X4 U11603 ( .A(n12612), .Z(n9764) );
  INV_X4 U11604 ( .A(n12797), .ZN(n17972) );
  AND2_X2 U11606 ( .A1(n13762), .A2(n14882), .ZN(n9747) );
  NAND2_X2 U11607 ( .A1(n9953), .A2(n11259), .ZN(n12176) );
  NAND2_X2 U11608 ( .A1(n9917), .A2(n20978), .ZN(n9953) );
  OAI211_X2 U11609 ( .C1(n10920), .C2(n14877), .A(n10360), .B(n10359), .ZN(
        n10404) );
  NAND2_X2 U11610 ( .A1(n9952), .A2(n11190), .ZN(n11254) );
  OAI21_X2 U11611 ( .B1(n14771), .B2(n10826), .A(n14785), .ZN(n14774) );
  NAND2_X2 U11612 ( .A1(n10539), .A2(n10878), .ZN(n14771) );
  OAI21_X4 U11613 ( .B1(n12176), .B2(n11412), .A(n11306), .ZN(n11313) );
  AND2_X2 U11614 ( .A1(n13746), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n9753) );
  AND2_X1 U11615 ( .A1(n20755), .A2(n20333), .ZN(n11752) );
  INV_X2 U11616 ( .A(n14929), .ZN(n9757) );
  INV_X2 U11617 ( .A(n14929), .ZN(n9758) );
  NAND3_X4 U11618 ( .A1(n14882), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14929) );
  OR2_X1 U11619 ( .A1(n13861), .A2(n10228), .ZN(n20978) );
  NAND2_X1 U11620 ( .A1(n10228), .A2(n13861), .ZN(n11267) );
  XNOR2_X1 U11621 ( .A(n9926), .B(n11257), .ZN(n13861) );
  XNOR2_X2 U11622 ( .A(n11313), .B(n13476), .ZN(n13449) );
  AND2_X2 U11623 ( .A1(n11050), .A2(n11049), .ZN(n9760) );
  NAND2_X2 U11624 ( .A1(n11335), .A2(n11296), .ZN(n13856) );
  OAI21_X2 U11625 ( .B1(n16060), .B2(n16063), .A(n16061), .ZN(n16041) );
  NAND2_X1 U11626 ( .A1(n11275), .A2(n11274), .ZN(n13294) );
  AOI22_X1 U11627 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n12057), .B1(n12056), 
        .B2(n20749), .ZN(n9765) );
  INV_X1 U11628 ( .A(n14197), .ZN(n9766) );
  AOI22_X1 U11631 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n12057), .B1(n12056), 
        .B2(n20749), .ZN(n14197) );
  AND2_X2 U11632 ( .A1(n10573), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10460) );
  OR2_X1 U11633 ( .A1(n10364), .A2(n10363), .ZN(n9877) );
  AND2_X1 U11634 ( .A1(n16673), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11427) );
  NOR2_X1 U11635 ( .A1(n13314), .A2(n20767), .ZN(n13527) );
  NAND2_X1 U11636 ( .A1(n13393), .A2(n11554), .ZN(n11197) );
  NAND3_X1 U11637 ( .A1(n11677), .A2(n11192), .A3(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n11520) );
  NAND2_X1 U11638 ( .A1(n14771), .A2(n9812), .ZN(n9872) );
  AND2_X1 U11639 ( .A1(n13592), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10344) );
  NAND2_X1 U11640 ( .A1(n11735), .A2(n13119), .ZN(n9878) );
  NAND2_X1 U11641 ( .A1(n12882), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n12805) );
  NAND2_X1 U11642 ( .A1(n9735), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n12804) );
  NOR2_X1 U11643 ( .A1(n18182), .A2(n12894), .ZN(n12909) );
  OAI211_X1 U11644 ( .C1(n16524), .C2(n12945), .A(n12762), .B(n9858), .ZN(
        n12763) );
  NAND2_X1 U11645 ( .A1(n11429), .A2(n11277), .ZN(n11500) );
  INV_X1 U11646 ( .A(n11520), .ZN(n11529) );
  NOR2_X1 U11647 ( .A1(n9936), .A2(n10815), .ZN(n10845) );
  OR2_X1 U11648 ( .A1(n16130), .A2(n16307), .ZN(n16120) );
  OR2_X1 U11649 ( .A1(n16185), .A2(n12004), .ZN(n16130) );
  NAND2_X1 U11650 ( .A1(n10908), .A2(n10907), .ZN(n16148) );
  INV_X1 U11651 ( .A(n10909), .ZN(n10908) );
  INV_X1 U11652 ( .A(n10929), .ZN(n11027) );
  NAND2_X1 U11653 ( .A1(n10396), .A2(n10397), .ZN(n10001) );
  NAND2_X1 U11654 ( .A1(n13412), .A2(n13419), .ZN(n13418) );
  OR2_X1 U11655 ( .A1(n14878), .A2(n13360), .ZN(n13427) );
  NAND2_X1 U11656 ( .A1(n11709), .A2(n11708), .ZN(n13132) );
  INV_X1 U11657 ( .A(n9904), .ZN(n9903) );
  NAND2_X1 U11658 ( .A1(n14692), .A2(n19484), .ZN(n16455) );
  AND4_X1 U11659 ( .A1(n11167), .A2(n11166), .A3(n11165), .A4(n11164), .ZN(
        n11173) );
  AND2_X1 U11660 ( .A1(n10176), .A2(n12514), .ZN(n10175) );
  AND2_X1 U11661 ( .A1(n10116), .A2(n16645), .ZN(n10114) );
  NAND2_X1 U11662 ( .A1(n11462), .A2(n16673), .ZN(n15637) );
  NAND2_X1 U11663 ( .A1(n11543), .A2(n11542), .ZN(n11679) );
  AOI21_X1 U11664 ( .B1(n15899), .B2(n10050), .A(n9834), .ZN(n10052) );
  INV_X1 U11665 ( .A(n10053), .ZN(n10050) );
  OR2_X1 U11666 ( .A1(n10190), .A2(n9965), .ZN(n9963) );
  OR2_X1 U11667 ( .A1(n10191), .A2(n10829), .ZN(n10190) );
  OAI21_X1 U11668 ( .B1(n16157), .B2(n16096), .A(n9807), .ZN(n10151) );
  AND2_X1 U11669 ( .A1(n10148), .A2(n9820), .ZN(n10147) );
  OR2_X1 U11670 ( .A1(n16179), .A2(n10708), .ZN(n10160) );
  NAND2_X1 U11671 ( .A1(n10906), .A2(n14384), .ZN(n10187) );
  OAI21_X1 U11672 ( .B1(n14691), .B2(n9863), .A(n14694), .ZN(n16523) );
  AND2_X1 U11673 ( .A1(n18272), .A2(n17101), .ZN(n9863) );
  INV_X1 U11674 ( .A(n19040), .ZN(n17101) );
  INV_X1 U11675 ( .A(n12931), .ZN(n18509) );
  OAI211_X1 U11676 ( .C1(n17720), .C2(n17958), .A(n12922), .B(n12921), .ZN(
        n17103) );
  NAND2_X1 U11677 ( .A1(n13255), .A2(n13651), .ZN(n21285) );
  CLKBUF_X1 U11678 ( .A(n19965), .Z(n19969) );
  NOR2_X1 U11679 ( .A1(n11507), .A2(n9985), .ZN(n11512) );
  AND2_X1 U11680 ( .A1(n11529), .A2(n11513), .ZN(n9985) );
  OAI21_X1 U11681 ( .B1(n11506), .B2(n11524), .A(n11505), .ZN(n11511) );
  NAND2_X1 U11682 ( .A1(n11512), .A2(n11511), .ZN(n9984) );
  NAND2_X1 U11683 ( .A1(n11526), .A2(n11513), .ZN(n9983) );
  AND2_X1 U11684 ( .A1(n11500), .A2(n11496), .ZN(n11516) );
  NAND2_X1 U11685 ( .A1(n12395), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n9977) );
  BUF_X1 U11686 ( .A(n11390), .Z(n12605) );
  NAND2_X1 U11687 ( .A1(n11364), .A2(n11363), .ZN(n9973) );
  NAND2_X1 U11688 ( .A1(n9797), .A2(n11307), .ZN(n10111) );
  NAND2_X1 U11689 ( .A1(n13936), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11429) );
  NAND2_X1 U11690 ( .A1(n13880), .A2(n11175), .ZN(n9951) );
  NAND2_X1 U11691 ( .A1(n11185), .A2(n11179), .ZN(n9948) );
  NAND2_X1 U11692 ( .A1(n10274), .A2(n11990), .ZN(n10346) );
  AND3_X1 U11693 ( .A1(n11994), .A2(n13368), .A3(n10325), .ZN(n10274) );
  NOR2_X1 U11694 ( .A1(n10707), .A2(n10705), .ZN(n10712) );
  NAND2_X1 U11695 ( .A1(n14785), .A2(n9871), .ZN(n9870) );
  AND2_X1 U11696 ( .A1(n10826), .A2(n17065), .ZN(n9871) );
  NAND2_X1 U11697 ( .A1(n11988), .A2(n11990), .ZN(n9881) );
  NOR2_X2 U11698 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10461) );
  INV_X1 U11699 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10229) );
  NAND2_X1 U11700 ( .A1(n12956), .A2(n12758), .ZN(n12766) );
  INV_X1 U11701 ( .A(n18175), .ZN(n12967) );
  AOI21_X1 U11702 ( .B1(n9895), .B2(n18683), .A(n9891), .ZN(n12973) );
  NAND2_X1 U11703 ( .A1(n20845), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13937) );
  NOR2_X1 U11704 ( .A1(n11198), .A2(n14704), .ZN(n13051) );
  NOR2_X1 U11705 ( .A1(n14764), .A2(n15182), .ZN(n10183) );
  OR2_X1 U11706 ( .A1(n15512), .A2(n15510), .ZN(n12426) );
  NAND2_X1 U11707 ( .A1(n13996), .A2(n13990), .ZN(n10173) );
  NOR2_X1 U11708 ( .A1(n10135), .A2(n11675), .ZN(n10134) );
  INV_X1 U11709 ( .A(n10136), .ZN(n10135) );
  NAND2_X1 U11710 ( .A1(n11364), .A2(n9816), .ZN(n11411) );
  NAND2_X1 U11711 ( .A1(n10133), .A2(n11596), .ZN(n10132) );
  INV_X1 U11712 ( .A(n13559), .ZN(n10133) );
  OR2_X1 U11713 ( .A1(n11332), .A2(n11331), .ZN(n11355) );
  NAND2_X1 U11714 ( .A1(n12128), .A2(n13275), .ZN(n11589) );
  INV_X1 U11715 ( .A(n13457), .ZN(n11596) );
  NAND2_X1 U11716 ( .A1(n11182), .A2(n13936), .ZN(n11563) );
  NOR2_X1 U11717 ( .A1(n10111), .A2(n10107), .ZN(n10101) );
  INV_X1 U11718 ( .A(n10111), .ZN(n10105) );
  AND2_X1 U11719 ( .A1(n11230), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10104) );
  NAND2_X1 U11720 ( .A1(n9927), .A2(n11256), .ZN(n9926) );
  NAND2_X1 U11721 ( .A1(n11268), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n9927) );
  AOI21_X1 U11722 ( .B1(n10107), .B2(n11307), .A(n10164), .ZN(n10163) );
  NAND2_X1 U11723 ( .A1(n11230), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10166) );
  AND2_X1 U11724 ( .A1(n11267), .A2(n9954), .ZN(n9917) );
  NAND2_X1 U11725 ( .A1(n10727), .A2(n19958), .ZN(n10733) );
  NAND2_X1 U11726 ( .A1(n10824), .A2(n10733), .ZN(n10730) );
  NAND2_X1 U11727 ( .A1(n10712), .A2(n10704), .ZN(n10714) );
  NOR2_X1 U11728 ( .A1(n10578), .A2(n10579), .ZN(n10572) );
  NAND2_X1 U11729 ( .A1(n10571), .A2(n10572), .ZN(n10646) );
  AND2_X1 U11730 ( .A1(n14480), .A2(n13636), .ZN(n10062) );
  NOR2_X1 U11731 ( .A1(n14436), .A2(n16107), .ZN(n10015) );
  INV_X1 U11732 ( .A(n10931), .ZN(n10929) );
  INV_X1 U11733 ( .A(n9890), .ZN(n13027) );
  OR2_X1 U11734 ( .A1(n10832), .A2(n9850), .ZN(n9934) );
  INV_X1 U11735 ( .A(n13028), .ZN(n9935) );
  NAND2_X2 U11736 ( .A1(n10351), .A2(n10354), .ZN(n10925) );
  NOR2_X1 U11737 ( .A1(n16158), .A2(n16096), .ZN(n10150) );
  AND2_X1 U11738 ( .A1(n14303), .A2(n14372), .ZN(n10066) );
  INV_X1 U11739 ( .A(n13575), .ZN(n10063) );
  NAND2_X1 U11740 ( .A1(n10065), .A2(n13473), .ZN(n10064) );
  INV_X1 U11741 ( .A(n13403), .ZN(n10065) );
  INV_X1 U11742 ( .A(n10703), .ZN(n9886) );
  NOR2_X1 U11743 ( .A1(n10158), .A2(n16991), .ZN(n10157) );
  INV_X1 U11744 ( .A(n10159), .ZN(n10158) );
  OAI21_X1 U11745 ( .B1(n16991), .B2(n10156), .A(n10224), .ZN(n10155) );
  NAND2_X1 U11746 ( .A1(n10159), .A2(n10708), .ZN(n10156) );
  AND2_X1 U11747 ( .A1(n10711), .A2(n16403), .ZN(n10159) );
  OR2_X1 U11748 ( .A1(n13368), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n10213) );
  INV_X1 U11749 ( .A(n12037), .ZN(n11972) );
  NOR2_X1 U11750 ( .A1(n13468), .A2(n10006), .ZN(n10005) );
  INV_X1 U11751 ( .A(n13504), .ZN(n10006) );
  INV_X1 U11752 ( .A(n10696), .ZN(n9970) );
  AND3_X1 U11753 ( .A1(n10324), .A2(n10323), .A3(n20333), .ZN(n11782) );
  MUX2_X1 U11754 ( .A(n10328), .B(n13374), .S(n11990), .Z(n10330) );
  AND2_X1 U11755 ( .A1(n9875), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n9874) );
  NAND2_X1 U11756 ( .A1(n10306), .A2(n11782), .ZN(n11953) );
  INV_X1 U11757 ( .A(n18412), .ZN(n10038) );
  INV_X1 U11758 ( .A(n12674), .ZN(n12677) );
  NOR2_X1 U11759 ( .A1(n19656), .A2(n12676), .ZN(n12684) );
  INV_X1 U11760 ( .A(n12665), .ZN(n12666) );
  OR2_X1 U11761 ( .A1(n12769), .A2(n19493), .ZN(n16452) );
  NOR2_X1 U11762 ( .A1(n18602), .A2(n12926), .ZN(n12927) );
  INV_X1 U11763 ( .A(n9907), .ZN(n12925) );
  XOR2_X1 U11764 ( .A(n12894), .B(n12980), .Z(n12881) );
  NAND2_X1 U11765 ( .A1(n19044), .A2(n19048), .ZN(n19493) );
  AND2_X1 U11766 ( .A1(n12839), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n9860) );
  AND2_X1 U11767 ( .A1(n9779), .A2(n9840), .ZN(n10138) );
  NOR2_X1 U11768 ( .A1(n12577), .A2(n13024), .ZN(n12578) );
  NAND2_X1 U11769 ( .A1(n12534), .A2(n9810), .ZN(n13014) );
  NAND2_X1 U11770 ( .A1(n12534), .A2(n12533), .ZN(n14763) );
  NAND2_X1 U11771 ( .A1(n9847), .A2(n9980), .ZN(n9979) );
  NAND2_X1 U11772 ( .A1(n12117), .A2(n12116), .ZN(n9916) );
  OR2_X1 U11773 ( .A1(n16673), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11428) );
  INV_X1 U11774 ( .A(n13824), .ZN(n11607) );
  INV_X1 U11775 ( .A(n13823), .ZN(n11608) );
  NAND2_X1 U11776 ( .A1(n9996), .A2(n9995), .ZN(n15788) );
  INV_X1 U11777 ( .A(n20932), .ZN(n9996) );
  INV_X1 U11778 ( .A(n20934), .ZN(n9995) );
  NAND2_X1 U11779 ( .A1(n11312), .A2(n11311), .ZN(n13474) );
  NAND4_X1 U11780 ( .A1(n11260), .A2(n11251), .A3(n11259), .A4(n9953), .ZN(
        n12175) );
  NOR2_X1 U11781 ( .A1(n9990), .A2(n9817), .ZN(n13314) );
  NOR2_X1 U11782 ( .A1(n11533), .A2(n9991), .ZN(n9990) );
  NAND2_X1 U11783 ( .A1(n11534), .A2(n9992), .ZN(n9991) );
  NOR2_X1 U11784 ( .A1(n15812), .A2(n12170), .ZN(n21006) );
  OR2_X1 U11785 ( .A1(n15812), .A2(n14398), .ZN(n14587) );
  AND2_X1 U11786 ( .A1(n16839), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n11537) );
  NAND2_X2 U11787 ( .A1(n20755), .A2(n20750), .ZN(n11730) );
  AND2_X1 U11788 ( .A1(n11987), .A2(n11986), .ZN(n13754) );
  NAND2_X1 U11789 ( .A1(n10830), .A2(n13029), .ZN(n13033) );
  AND2_X1 U11790 ( .A1(n10000), .A2(n9799), .ZN(n14857) );
  OR2_X1 U11791 ( .A1(n15890), .A2(n15900), .ZN(n10053) );
  NOR2_X1 U11792 ( .A1(n15075), .A2(n15076), .ZN(n15899) );
  AOI21_X1 U11793 ( .B1(n16914), .B2(n16912), .A(n15005), .ZN(n15028) );
  NAND2_X1 U11794 ( .A1(n14903), .A2(n15998), .ZN(n15997) );
  NAND2_X1 U11795 ( .A1(n12084), .A2(n10078), .ZN(n11036) );
  AND2_X1 U11796 ( .A1(n9781), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10078) );
  NAND2_X1 U11797 ( .A1(n15856), .A2(n10019), .ZN(n14808) );
  NOR2_X1 U11798 ( .A1(n10020), .A2(n13037), .ZN(n10019) );
  INV_X1 U11799 ( .A(n10021), .ZN(n10020) );
  INV_X1 U11800 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n14786) );
  AND2_X1 U11801 ( .A1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n16121), .ZN(
        n10913) );
  NOR2_X1 U11802 ( .A1(n16120), .A2(n16297), .ZN(n10914) );
  AND2_X1 U11803 ( .A1(n19757), .A2(n10792), .ZN(n16118) );
  AOI21_X1 U11804 ( .B1(n16944), .B2(n16941), .A(n16091), .ZN(n16170) );
  NAND2_X1 U11805 ( .A1(n9784), .A2(n14285), .ZN(n14284) );
  NAND2_X1 U11806 ( .A1(n14382), .A2(n14381), .ZN(n9885) );
  NAND2_X1 U11807 ( .A1(n10901), .A2(n10900), .ZN(n10902) );
  NAND2_X1 U11808 ( .A1(n9889), .A2(n9888), .ZN(n10539) );
  AND2_X1 U11809 ( .A1(n13427), .A2(n13361), .ZN(n13362) );
  INV_X1 U11810 ( .A(n11692), .ZN(n13142) );
  AND2_X1 U11811 ( .A1(n20098), .A2(n11994), .ZN(n10308) );
  NAND2_X1 U11812 ( .A1(n10161), .A2(n15888), .ZN(n10184) );
  OR2_X1 U11813 ( .A1(n20706), .A2(n20718), .ZN(n20473) );
  NAND2_X1 U11814 ( .A1(n13582), .A2(n13581), .ZN(n20512) );
  NAND2_X1 U11815 ( .A1(n17082), .A2(n20749), .ZN(n13582) );
  INV_X1 U11816 ( .A(n20750), .ZN(n13592) );
  OR2_X1 U11817 ( .A1(n20706), .A2(n20074), .ZN(n20308) );
  INV_X1 U11818 ( .A(n20512), .ZN(n20551) );
  NAND2_X1 U11819 ( .A1(n17576), .A2(n18370), .ZN(n10026) );
  OR2_X1 U11820 ( .A1(n17344), .A2(n10027), .ZN(n10025) );
  NAND2_X1 U11821 ( .A1(n18370), .A2(n10028), .ZN(n10027) );
  NAND2_X1 U11822 ( .A1(n17576), .A2(n10038), .ZN(n10035) );
  OR2_X1 U11823 ( .A1(n17370), .A2(n10036), .ZN(n10034) );
  NAND2_X1 U11824 ( .A1(n10038), .A2(n10037), .ZN(n10036) );
  INV_X1 U11825 ( .A(n18425), .ZN(n10037) );
  NAND2_X1 U11826 ( .A1(n12658), .A2(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12660) );
  AND2_X1 U11827 ( .A1(n9735), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n9894)
         );
  NOR2_X1 U11828 ( .A1(n17913), .A2(n19081), .ZN(n12834) );
  NAND2_X1 U11829 ( .A1(n17970), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n12823) );
  NOR2_X1 U11830 ( .A1(n9770), .A2(n18368), .ZN(n18355) );
  NAND2_X1 U11831 ( .A1(n10032), .A2(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n10031) );
  INV_X1 U11832 ( .A(n18447), .ZN(n10032) );
  AND3_X1 U11833 ( .A1(n17507), .A2(n10212), .A3(n10043), .ZN(n18468) );
  AND2_X1 U11834 ( .A1(n10045), .A2(n10044), .ZN(n10043) );
  INV_X1 U11835 ( .A(n18484), .ZN(n10044) );
  INV_X1 U11836 ( .A(n18374), .ZN(n18384) );
  INV_X1 U11837 ( .A(n10093), .ZN(n12896) );
  NOR2_X1 U11838 ( .A1(n18873), .A2(n19515), .ZN(n18931) );
  INV_X1 U11839 ( .A(n19044), .ZN(n12947) );
  NOR2_X1 U11840 ( .A1(n12681), .A2(n12680), .ZN(n12682) );
  NOR2_X1 U11841 ( .A1(n10129), .A2(n9813), .ZN(n10128) );
  INV_X1 U11842 ( .A(n15159), .ZN(n10129) );
  AND2_X1 U11843 ( .A1(n20845), .A2(n13933), .ZN(n20808) );
  XNOR2_X1 U11844 ( .A(n14734), .B(n13048), .ZN(n15612) );
  AOI21_X1 U11845 ( .B1(n16722), .B2(n14723), .A(n13025), .ZN(n13026) );
  AND2_X1 U11846 ( .A1(n14815), .A2(n13065), .ZN(n15469) );
  XNOR2_X1 U11847 ( .A(n13023), .B(n15692), .ZN(n15699) );
  NAND2_X1 U11848 ( .A1(n15620), .A2(n13021), .ZN(n11467) );
  NOR2_X1 U11849 ( .A1(n15733), .A2(n15788), .ZN(n15738) );
  NAND2_X1 U11850 ( .A1(n11679), .A2(n11552), .ZN(n16792) );
  NAND2_X1 U11851 ( .A1(n11679), .A2(n11678), .ZN(n20925) );
  INV_X1 U11852 ( .A(n16792), .ZN(n20927) );
  INV_X1 U11853 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n16839) );
  INV_X1 U11854 ( .A(n16847), .ZN(n10077) );
  CLKBUF_X1 U11855 ( .A(n19910), .Z(n19897) );
  XNOR2_X1 U11856 ( .A(n9999), .B(n11031), .ZN(n12092) );
  XOR2_X1 U11857 ( .A(n11731), .B(n15892), .Z(n16845) );
  AOI21_X1 U11858 ( .B1(n13354), .B2(n13744), .A(n17088), .ZN(n19965) );
  OR2_X1 U11859 ( .A1(n12092), .A2(n16202), .ZN(n9998) );
  NAND2_X1 U11860 ( .A1(n13114), .A2(n11032), .ZN(n20055) );
  AND2_X1 U11861 ( .A1(n20055), .A2(n20713), .ZN(n20051) );
  AND2_X1 U11862 ( .A1(n20055), .A2(n13252), .ZN(n17008) );
  OR2_X1 U11863 ( .A1(n9792), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14805) );
  NAND2_X1 U11864 ( .A1(n16869), .A2(n17074), .ZN(n10071) );
  NOR3_X1 U11865 ( .A1(n10070), .A2(n14844), .A3(n10069), .ZN(n10068) );
  INV_X1 U11866 ( .A(n16207), .ZN(n10069) );
  NOR2_X1 U11867 ( .A1(n16208), .A2(n10828), .ZN(n10070) );
  OR2_X1 U11868 ( .A1(n9792), .A2(n13035), .ZN(n14798) );
  INV_X1 U11869 ( .A(n20068), .ZN(n17052) );
  INV_X1 U11870 ( .A(n20062), .ZN(n17074) );
  INV_X1 U11871 ( .A(n17048), .ZN(n20057) );
  OR2_X1 U11872 ( .A1(n14878), .A2(n13352), .ZN(n20727) );
  INV_X1 U11873 ( .A(n13512), .ZN(n13513) );
  INV_X1 U11874 ( .A(n20245), .ZN(n20223) );
  NOR2_X1 U11875 ( .A1(n17401), .A2(n18462), .ZN(n17400) );
  NOR2_X1 U11876 ( .A1(n17962), .A2(n17986), .ZN(n17942) );
  NAND2_X1 U11877 ( .A1(P3_EBX_REG_9__SCAN_IN), .A2(n17987), .ZN(n17986) );
  OR2_X1 U11878 ( .A1(n16456), .A2(n19546), .ZN(n9857) );
  OR2_X1 U11879 ( .A1(n18198), .A2(P3_EAX_REG_30__SCAN_IN), .ZN(n9861) );
  NAND2_X1 U11880 ( .A1(n18062), .A2(n18190), .ZN(n18060) );
  NOR2_X1 U11881 ( .A1(n18073), .A2(n18211), .ZN(n18068) );
  NAND2_X1 U11882 ( .A1(n18068), .A2(P3_EAX_REG_29__SCAN_IN), .ZN(n18062) );
  INV_X1 U11883 ( .A(n18098), .ZN(n18130) );
  INV_X1 U11884 ( .A(n18104), .ZN(n18131) );
  NAND2_X1 U11885 ( .A1(n10218), .A2(n9844), .ZN(n9862) );
  INV_X1 U11886 ( .A(n18114), .ZN(n18190) );
  NAND2_X1 U11887 ( .A1(n18049), .A2(P3_EAX_REG_1__SCAN_IN), .ZN(n18199) );
  INV_X1 U11888 ( .A(n18192), .ZN(n18196) );
  INV_X1 U11889 ( .A(n9901), .ZN(n9900) );
  NAND2_X1 U11890 ( .A1(n19012), .A2(n17103), .ZN(n18877) );
  NAND2_X1 U11891 ( .A1(n19040), .A2(n18931), .ZN(n19483) );
  INV_X1 U11892 ( .A(n18995), .ZN(n19014) );
  NOR2_X1 U11893 ( .A1(n17149), .A2(n19014), .ZN(n19012) );
  OAI21_X1 U11894 ( .B1(n12760), .B2(n12947), .A(n12946), .ZN(n9858) );
  AOI21_X1 U11895 ( .B1(n12839), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A(
        n9856), .ZN(n9855) );
  OAI22_X1 U11896 ( .A1(n17975), .A2(n17918), .B1(n17995), .B2(n17915), .ZN(
        n9856) );
  NAND2_X1 U11897 ( .A1(n17864), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n9854) );
  NAND2_X1 U11898 ( .A1(n9745), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n11141) );
  OR2_X1 U11899 ( .A1(n11351), .A2(n11350), .ZN(n11379) );
  NAND2_X1 U11900 ( .A1(n11490), .A2(n15821), .ZN(n11193) );
  AND2_X1 U11901 ( .A1(n11193), .A2(n11198), .ZN(n11186) );
  OR2_X1 U11902 ( .A1(n11244), .A2(n11243), .ZN(n11303) );
  OAI22_X1 U11903 ( .A1(n9982), .A2(n11519), .B1(n11518), .B2(n11517), .ZN(
        n11522) );
  AOI22_X1 U11904 ( .A1(n9984), .A2(n9983), .B1(n11514), .B2(n11515), .ZN(
        n9982) );
  NAND2_X1 U11905 ( .A1(n10333), .A2(n10332), .ZN(n11711) );
  NOR2_X1 U11906 ( .A1(n9945), .A2(n9777), .ZN(n9944) );
  CLKBUF_X1 U11907 ( .A(n14929), .Z(n14930) );
  NOR2_X1 U11908 ( .A1(n9969), .A2(n11777), .ZN(n9968) );
  INV_X1 U11909 ( .A(n10470), .ZN(n9969) );
  AND2_X1 U11910 ( .A1(n10644), .A2(n10643), .ZN(n10657) );
  OAI22_X1 U11911 ( .A1(n10472), .A2(n13810), .B1(n20367), .B2(n14164), .ZN(
        n10473) );
  NAND2_X1 U11912 ( .A1(n13119), .A2(n20755), .ZN(n10363) );
  NAND2_X1 U11913 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n14933) );
  NAND2_X1 U11914 ( .A1(n11711), .A2(n13368), .ZN(n11988) );
  AND2_X1 U11915 ( .A1(n10237), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9961) );
  NAND2_X1 U11916 ( .A1(n10336), .A2(n10306), .ZN(n10337) );
  AND2_X1 U11917 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n10449), .ZN(
        n10447) );
  AND2_X1 U11918 ( .A1(n20732), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10865) );
  AND2_X1 U11919 ( .A1(n12950), .A2(n12948), .ZN(n12771) );
  NOR2_X1 U11920 ( .A1(n10137), .A2(n15183), .ZN(n10136) );
  INV_X1 U11921 ( .A(n15479), .ZN(n10137) );
  NAND2_X1 U11922 ( .A1(n12606), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n11145) );
  NAND2_X1 U11923 ( .A1(n11385), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n9975) );
  NAND2_X1 U11924 ( .A1(n11159), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n9978) );
  AND2_X1 U11925 ( .A1(n15484), .A2(n10177), .ZN(n10176) );
  NOR2_X1 U11926 ( .A1(n15491), .A2(n15500), .ZN(n10177) );
  OR2_X1 U11927 ( .A1(n12406), .A2(n15519), .ZN(n15510) );
  OR2_X1 U11928 ( .A1(n12390), .A2(n15435), .ZN(n12371) );
  AND2_X1 U11929 ( .A1(n12285), .A2(n10181), .ZN(n10180) );
  INV_X1 U11930 ( .A(n15440), .ZN(n10181) );
  INV_X1 U11931 ( .A(n11377), .ZN(n9972) );
  NAND2_X1 U11932 ( .A1(n10113), .A2(n9931), .ZN(n11463) );
  INV_X1 U11933 ( .A(n15515), .ZN(n10139) );
  NAND2_X1 U11934 ( .A1(n9959), .A2(n15659), .ZN(n10118) );
  NAND2_X1 U11935 ( .A1(n10117), .A2(n15659), .ZN(n10116) );
  NAND2_X1 U11936 ( .A1(n10144), .A2(n10143), .ZN(n10142) );
  INV_X1 U11937 ( .A(n14292), .ZN(n10144) );
  NAND2_X1 U11938 ( .A1(n13275), .A2(n12132), .ZN(n11673) );
  NAND2_X1 U11939 ( .A1(n11585), .A2(n10125), .ZN(n11588) );
  AND2_X1 U11940 ( .A1(n11177), .A2(n9821), .ZN(n10123) );
  NAND2_X1 U11941 ( .A1(n13314), .A2(n9989), .ZN(n11535) );
  AND2_X1 U11942 ( .A1(n12320), .A2(n11177), .ZN(n9989) );
  AND2_X2 U11943 ( .A1(n11043), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11050) );
  AND2_X1 U11944 ( .A1(n11529), .A2(n11494), .ZN(n11524) );
  NAND2_X1 U11945 ( .A1(n9954), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n9992) );
  AND2_X1 U11946 ( .A1(n11475), .A2(n11476), .ZN(n11495) );
  NOR2_X1 U11947 ( .A1(n11063), .A2(n11062), .ZN(n11068) );
  OAI21_X1 U11948 ( .B1(n21291), .B2(n16835), .A(n16498), .ZN(n13858) );
  NAND2_X1 U11949 ( .A1(n14055), .A2(n9954), .ZN(n11334) );
  INV_X1 U11950 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n21009) );
  NOR2_X1 U11951 ( .A1(n13033), .A2(n10837), .ZN(n10840) );
  AND2_X1 U11952 ( .A1(n10736), .A2(n10763), .ZN(n10762) );
  NAND2_X1 U11953 ( .A1(n10838), .A2(P2_EBX_REG_2__SCAN_IN), .ZN(n9942) );
  NAND2_X1 U11954 ( .A1(n10850), .A2(n10306), .ZN(n9943) );
  NAND2_X1 U11955 ( .A1(n10391), .A2(n10390), .ZN(n10917) );
  NAND2_X1 U11956 ( .A1(n15054), .A2(n15053), .ZN(n15078) );
  AOI21_X1 U11957 ( .B1(n15028), .B2(n10060), .A(n10059), .ZN(n15052) );
  AND2_X1 U11958 ( .A1(n15027), .A2(n15917), .ZN(n10059) );
  OR2_X1 U11959 ( .A1(n15027), .A2(n15917), .ZN(n10060) );
  NOR2_X1 U11960 ( .A1(n10518), .A2(n10517), .ZN(n11756) );
  NOR2_X1 U11961 ( .A1(n12089), .A2(n10080), .ZN(n10079) );
  NOR2_X1 U11962 ( .A1(n10023), .A2(n10022), .ZN(n10021) );
  INV_X1 U11963 ( .A(n15910), .ZN(n10022) );
  INV_X1 U11964 ( .A(n15846), .ZN(n10023) );
  NAND2_X1 U11965 ( .A1(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n10086) );
  NOR2_X1 U11966 ( .A1(n16971), .A2(n10083), .ZN(n10082) );
  INV_X1 U11967 ( .A(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n10083) );
  NOR2_X1 U11968 ( .A1(n17014), .A2(n10091), .ZN(n10090) );
  INV_X1 U11969 ( .A(n12061), .ZN(n10089) );
  NAND2_X1 U11970 ( .A1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n12060) );
  AND2_X1 U11971 ( .A1(n15837), .A2(n15960), .ZN(n10073) );
  NAND2_X1 U11972 ( .A1(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n10191) );
  NAND2_X1 U11973 ( .A1(n12006), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n9965) );
  OR2_X1 U11974 ( .A1(n15865), .A2(n11790), .ZN(n10818) );
  NAND2_X1 U11975 ( .A1(n9807), .A2(n16096), .ZN(n10148) );
  AND2_X1 U11976 ( .A1(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n10219), .ZN(
        n16121) );
  NOR2_X1 U11977 ( .A1(n10012), .A2(n10011), .ZN(n10010) );
  INV_X1 U11978 ( .A(n13715), .ZN(n10011) );
  INV_X1 U11979 ( .A(n10966), .ZN(n10012) );
  NAND2_X1 U11980 ( .A1(n14263), .A2(n14260), .ZN(n10899) );
  NAND2_X1 U11981 ( .A1(n9872), .A2(n9869), .ZN(n9873) );
  AND2_X1 U11982 ( .A1(n14772), .A2(n9870), .ZN(n9869) );
  NAND2_X1 U11983 ( .A1(n10384), .A2(n10383), .ZN(n10385) );
  OAI211_X1 U11984 ( .C1(n10931), .C2(n10380), .A(n10379), .B(n10378), .ZN(
        n10381) );
  NOR2_X1 U11985 ( .A1(n10506), .A2(n10505), .ZN(n11748) );
  INV_X1 U11986 ( .A(n14933), .ZN(n10449) );
  NAND2_X1 U11987 ( .A1(n13426), .A2(n13425), .ZN(n13431) );
  INV_X1 U11988 ( .A(n10447), .ZN(n10870) );
  NOR2_X1 U11989 ( .A1(n13420), .A2(n10425), .ZN(n10426) );
  NAND2_X1 U11990 ( .A1(n13412), .A2(n15873), .ZN(n10418) );
  AOI22_X1 U11991 ( .A1(n10315), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n10316), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10275) );
  NAND2_X1 U11992 ( .A1(n20711), .A2(n20512), .ZN(n13587) );
  CLKBUF_X1 U11993 ( .A(n12797), .Z(n17643) );
  NAND2_X1 U11994 ( .A1(n12663), .A2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12674) );
  INV_X1 U11995 ( .A(n12810), .ZN(n9898) );
  AOI21_X1 U11996 ( .B1(n17864), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A(
        n12803), .ZN(n12809) );
  NOR2_X1 U11997 ( .A1(n17958), .A2(n12802), .ZN(n12803) );
  AND2_X1 U11998 ( .A1(n12839), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n12813) );
  INV_X1 U11999 ( .A(n17827), .ZN(n12830) );
  NAND2_X1 U12000 ( .A1(n12754), .A2(n12766), .ZN(n12995) );
  NOR2_X1 U12001 ( .A1(n18506), .A2(n10046), .ZN(n10045) );
  INV_X1 U12002 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n10046) );
  NOR2_X1 U12003 ( .A1(n18605), .A2(n18606), .ZN(n12988) );
  NAND2_X1 U12004 ( .A1(n12928), .A2(n9845), .ZN(n10096) );
  AND2_X1 U12005 ( .A1(n12931), .A2(n18919), .ZN(n12928) );
  AND2_X1 U12006 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n12910), .ZN(
        n12911) );
  NOR2_X1 U12007 ( .A1(n12995), .A2(n19494), .ZN(n14692) );
  AOI21_X1 U12008 ( .B1(n12998), .B2(n12997), .A(n12996), .ZN(n19492) );
  NAND2_X1 U12009 ( .A1(n12839), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n12678) );
  OAI211_X1 U12010 ( .C1(n17879), .C2(n17818), .A(n12715), .B(n12714), .ZN(
        n12759) );
  OAI211_X1 U12011 ( .C1(n17811), .C2(n17827), .A(n12753), .B(n12752), .ZN(
        n12945) );
  NOR2_X1 U12012 ( .A1(n12751), .A2(n9853), .ZN(n12752) );
  AOI211_X1 U12013 ( .C1(n17979), .C2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A(
        n12702), .B(n12701), .ZN(n12703) );
  NAND2_X1 U12014 ( .A1(n13953), .A2(n13945), .ZN(n20813) );
  OR2_X1 U12015 ( .A1(n21285), .A2(n13930), .ZN(n20845) );
  NAND2_X1 U12016 ( .A1(n15478), .A2(n10136), .ZN(n15184) );
  NOR2_X1 U12017 ( .A1(n13392), .A2(n21113), .ZN(n12631) );
  INV_X1 U12018 ( .A(n14735), .ZN(n10182) );
  AND2_X1 U12019 ( .A1(n12534), .A2(n10183), .ZN(n13015) );
  NAND2_X1 U12020 ( .A1(n12554), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n12577) );
  NOR2_X1 U12021 ( .A1(n12494), .A2(n12489), .ZN(n12495) );
  NOR2_X1 U12022 ( .A1(n12448), .A2(n12447), .ZN(n12449) );
  NAND2_X1 U12023 ( .A1(n12449), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n12494) );
  NAND2_X1 U12024 ( .A1(n12318), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12448) );
  AND2_X1 U12025 ( .A1(n12427), .A2(n9828), .ZN(n10179) );
  NOR2_X1 U12026 ( .A1(n12371), .A2(n15657), .ZN(n12372) );
  NOR2_X1 U12027 ( .A1(n12317), .A2(n12316), .ZN(n12408) );
  NOR2_X1 U12028 ( .A1(n12286), .A2(n16625), .ZN(n12302) );
  NOR2_X1 U12029 ( .A1(n12257), .A2(n14658), .ZN(n12282) );
  NOR2_X1 U12030 ( .A1(n12234), .A2(n12230), .ZN(n12235) );
  AND2_X1 U12031 ( .A1(n13819), .A2(n10171), .ZN(n10170) );
  AND2_X1 U12032 ( .A1(n13837), .A2(n10172), .ZN(n10171) );
  NOR2_X1 U12033 ( .A1(n14278), .A2(n10173), .ZN(n10172) );
  AND2_X1 U12034 ( .A1(n13819), .A2(n10168), .ZN(n10167) );
  AND2_X1 U12035 ( .A1(n13837), .A2(n10169), .ZN(n10168) );
  INV_X1 U12036 ( .A(n10173), .ZN(n10169) );
  AND2_X1 U12037 ( .A1(n13837), .A2(n13996), .ZN(n10174) );
  NAND2_X1 U12038 ( .A1(n13819), .A2(n13837), .ZN(n14081) );
  NOR2_X1 U12039 ( .A1(n12210), .A2(n15346), .ZN(n12211) );
  INV_X1 U12040 ( .A(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n15346) );
  NAND2_X1 U12041 ( .A1(n12205), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12210) );
  AND2_X1 U12042 ( .A1(n12196), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12205) );
  INV_X1 U12043 ( .A(n12164), .ZN(n12186) );
  AND2_X1 U12044 ( .A1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n12186), .ZN(
        n12196) );
  OAI21_X1 U12045 ( .B1(n13856), .B2(n12300), .A(n12168), .ZN(n12169) );
  NAND2_X1 U12046 ( .A1(n15478), .A2(n9780), .ZN(n12130) );
  INV_X1 U12047 ( .A(n9981), .ZN(n9912) );
  AND2_X1 U12048 ( .A1(n16673), .A2(n11661), .ZN(n10119) );
  NAND2_X1 U12049 ( .A1(n15478), .A2(n15479), .ZN(n15481) );
  NOR2_X1 U12050 ( .A1(n15627), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15629) );
  NAND2_X1 U12051 ( .A1(n16581), .A2(n15515), .ZN(n15514) );
  NOR2_X1 U12052 ( .A1(n15522), .A2(n15521), .ZN(n16579) );
  AND2_X1 U12053 ( .A1(n16579), .A2(n16578), .ZN(n16581) );
  INV_X1 U12054 ( .A(n9959), .ZN(n11458) );
  OR2_X1 U12055 ( .A1(n15431), .A2(n15432), .ZN(n15522) );
  NOR2_X1 U12056 ( .A1(n15538), .A2(n15537), .ZN(n15540) );
  OR2_X1 U12057 ( .A1(n14673), .A2(n14683), .ZN(n15445) );
  NAND2_X1 U12058 ( .A1(n10122), .A2(n10121), .ZN(n15538) );
  INV_X1 U12059 ( .A(n15444), .ZN(n10121) );
  INV_X1 U12060 ( .A(n15445), .ZN(n10122) );
  NAND2_X1 U12061 ( .A1(n16673), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n15666) );
  NOR2_X1 U12062 ( .A1(n14121), .A2(n10140), .ZN(n14675) );
  NAND2_X1 U12063 ( .A1(n14575), .A2(n10141), .ZN(n10140) );
  INV_X1 U12064 ( .A(n10142), .ZN(n10141) );
  OR2_X1 U12065 ( .A1(n14121), .A2(n13992), .ZN(n14293) );
  NAND2_X1 U12066 ( .A1(n16727), .A2(n9922), .ZN(n9921) );
  INV_X1 U12067 ( .A(n14352), .ZN(n9920) );
  AND2_X1 U12068 ( .A1(n10164), .A2(n11494), .ZN(n9958) );
  AND2_X1 U12069 ( .A1(n15738), .A2(n15784), .ZN(n15800) );
  AND2_X1 U12070 ( .A1(n14083), .A2(n14082), .ZN(n14119) );
  AND3_X1 U12071 ( .A1(n11610), .A2(n11649), .A3(n11609), .ZN(n13840) );
  NOR2_X1 U12072 ( .A1(n13841), .A2(n13840), .ZN(n14083) );
  INV_X1 U12073 ( .A(n10132), .ZN(n10131) );
  NOR2_X1 U12074 ( .A1(n10132), .A2(n13458), .ZN(n13725) );
  INV_X1 U12075 ( .A(n15788), .ZN(n15736) );
  AND2_X1 U12076 ( .A1(n11595), .A2(n11594), .ZN(n13457) );
  OR2_X1 U12077 ( .A1(n11589), .A2(P1_EBX_REG_2__SCAN_IN), .ZN(n11595) );
  INV_X1 U12078 ( .A(n13275), .ZN(n14817) );
  NAND2_X1 U12079 ( .A1(n11601), .A2(n12132), .ZN(n14818) );
  NAND2_X1 U12080 ( .A1(n10105), .A2(n10104), .ZN(n10103) );
  NAND2_X1 U12081 ( .A1(n11267), .A2(n11266), .ZN(n11275) );
  NOR2_X1 U12082 ( .A1(n13298), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11291) );
  NAND2_X1 U12083 ( .A1(n12175), .A2(n11260), .ZN(n11295) );
  INV_X1 U12084 ( .A(n20982), .ZN(n20940) );
  INV_X1 U12085 ( .A(n11554), .ZN(n11178) );
  NAND3_X1 U12086 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n9954), .A3(n13858), 
        .ZN(n13979) );
  NOR2_X1 U12087 ( .A1(n20954), .A2(n14095), .ZN(n21016) );
  AOI21_X1 U12088 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n21110), .A(n14095), 
        .ZN(n21120) );
  NAND2_X1 U12089 ( .A1(n9954), .A2(n13858), .ZN(n14095) );
  NOR2_X1 U12090 ( .A1(n13856), .A2(n14088), .ZN(n14318) );
  INV_X1 U12091 ( .A(n13897), .ZN(n14313) );
  INV_X1 U12092 ( .A(n21268), .ZN(n16498) );
  NAND2_X1 U12093 ( .A1(n10820), .A2(n10845), .ZN(n10834) );
  OR2_X1 U12094 ( .A1(n12082), .A2(n15841), .ZN(n12086) );
  NOR2_X1 U12095 ( .A1(n12086), .A2(n12085), .ZN(n12084) );
  NAND2_X1 U12096 ( .A1(n15840), .A2(n16055), .ZN(n15839) );
  OR2_X1 U12097 ( .A1(n12079), .A2(n16068), .ZN(n12082) );
  NAND2_X1 U12098 ( .A1(n10802), .A2(n9938), .ZN(n10822) );
  NOR2_X1 U12099 ( .A1(n9941), .A2(n9939), .ZN(n9938) );
  NAND2_X1 U12100 ( .A1(n10814), .A2(n9940), .ZN(n9939) );
  NOR2_X1 U12101 ( .A1(n9941), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n9937) );
  NAND2_X1 U12102 ( .A1(n10802), .A2(n10803), .ZN(n10813) );
  NAND2_X1 U12103 ( .A1(n10781), .A2(n10780), .ZN(n10782) );
  NOR2_X1 U12104 ( .A1(n12074), .A2(n10086), .ZN(n12078) );
  NAND2_X1 U12105 ( .A1(n13828), .A2(n9833), .ZN(n16021) );
  NOR2_X1 U12106 ( .A1(n12072), .A2(n16161), .ZN(n12075) );
  NAND2_X1 U12107 ( .A1(n12073), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12072) );
  AND3_X1 U12108 ( .A1(n11850), .A2(n11849), .A3(n11848), .ZN(n13403) );
  NOR2_X1 U12109 ( .A1(n10714), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n10720) );
  NAND2_X1 U12110 ( .A1(n10717), .A2(n9947), .ZN(n9946) );
  AND3_X1 U12111 ( .A1(n11812), .A2(n11811), .A3(n11810), .ZN(n14200) );
  XNOR2_X1 U12112 ( .A(n15052), .B(n10220), .ZN(n15914) );
  AND2_X1 U12113 ( .A1(n11963), .A2(n11966), .ZN(n10074) );
  XNOR2_X1 U12114 ( .A(n15927), .B(n14979), .ZN(n15922) );
  NAND2_X1 U12115 ( .A1(n15922), .A2(n15921), .ZN(n15920) );
  INV_X1 U12116 ( .A(n14482), .ZN(n10061) );
  AND2_X1 U12117 ( .A1(n11789), .A2(n11788), .ZN(n13400) );
  NAND2_X1 U12118 ( .A1(n13440), .A2(n13439), .ZN(n13698) );
  AOI21_X1 U12119 ( .B1(n13434), .B2(n13438), .A(n13437), .ZN(n13439) );
  XNOR2_X1 U12120 ( .A(n11760), .B(n11755), .ZN(n13264) );
  INV_X1 U12121 ( .A(n20727), .ZN(n13961) );
  INV_X1 U12122 ( .A(n13374), .ZN(n13369) );
  AND2_X1 U12123 ( .A1(n12099), .A2(n13106), .ZN(n14205) );
  NAND2_X1 U12124 ( .A1(n12084), .A2(n10079), .ZN(n12091) );
  NOR3_X1 U12125 ( .A1(n12074), .A2(n10086), .A3(n10084), .ZN(n12080) );
  NAND2_X1 U12126 ( .A1(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n10084) );
  NOR2_X1 U12127 ( .A1(n10014), .A2(n10018), .ZN(n10013) );
  INV_X1 U12128 ( .A(n15925), .ZN(n10018) );
  INV_X1 U12129 ( .A(n10015), .ZN(n10014) );
  AND2_X1 U12130 ( .A1(n10994), .A2(n10993), .ZN(n16107) );
  NAND2_X1 U12131 ( .A1(n14435), .A2(n10989), .ZN(n16108) );
  INV_X1 U12132 ( .A(n14435), .ZN(n16139) );
  NOR2_X1 U12133 ( .A1(n12074), .A2(n19768), .ZN(n12076) );
  AND2_X1 U12134 ( .A1(n12070), .A2(n10081), .ZN(n12073) );
  AND2_X1 U12135 ( .A1(n9773), .A2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n10081) );
  NAND2_X1 U12136 ( .A1(n12070), .A2(n9773), .ZN(n12071) );
  AND2_X1 U12137 ( .A1(n13640), .A2(n10966), .ZN(n16966) );
  NAND2_X1 U12138 ( .A1(n12070), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n12069) );
  NOR2_X1 U12139 ( .A1(n12067), .A2(n16986), .ZN(n12070) );
  NAND2_X1 U12140 ( .A1(n12068), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n12067) );
  AND3_X1 U12141 ( .A1(n10952), .A2(n10951), .A3(n10950), .ZN(n14240) );
  NOR2_X1 U12142 ( .A1(n12065), .A2(n17007), .ZN(n12068) );
  AND2_X1 U12143 ( .A1(n10087), .A2(n10089), .ZN(n12066) );
  NOR2_X1 U12144 ( .A1(n10088), .A2(n16200), .ZN(n10087) );
  INV_X1 U12145 ( .A(n10090), .ZN(n10088) );
  NAND2_X1 U12146 ( .A1(n12066), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12065) );
  NAND2_X1 U12147 ( .A1(n10089), .A2(n10090), .ZN(n12063) );
  NOR2_X1 U12148 ( .A1(n12061), .A2(n17014), .ZN(n12064) );
  NAND2_X1 U12149 ( .A1(n10930), .A2(n14267), .ZN(n14268) );
  NOR2_X1 U12150 ( .A1(n14786), .A2(n12060), .ZN(n12062) );
  NAND2_X1 U12151 ( .A1(n12062), .A2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12061) );
  NAND2_X1 U12152 ( .A1(n15894), .A2(n15893), .ZN(n15892) );
  NAND2_X1 U12153 ( .A1(n9933), .A2(n9932), .ZN(n16032) );
  AOI21_X1 U12154 ( .B1(n10832), .B2(n10833), .A(n9935), .ZN(n9932) );
  NAND2_X1 U12155 ( .A1(n13027), .A2(n9934), .ZN(n9933) );
  NAND2_X1 U12156 ( .A1(n9890), .A2(n13028), .ZN(n14800) );
  NAND2_X1 U12157 ( .A1(n10017), .A2(n10016), .ZN(n15855) );
  INV_X1 U12158 ( .A(n14750), .ZN(n10016) );
  INV_X1 U12159 ( .A(n14749), .ZN(n10017) );
  AND2_X1 U12160 ( .A1(n16095), .A2(n16094), .ZN(n16158) );
  NAND2_X1 U12161 ( .A1(n13640), .A2(n10008), .ZN(n16947) );
  NOR2_X1 U12162 ( .A1(n10009), .A2(n16945), .ZN(n10008) );
  INV_X1 U12163 ( .A(n10010), .ZN(n10009) );
  AND3_X1 U12164 ( .A1(n10977), .A2(n10976), .A3(n10975), .ZN(n14254) );
  NOR2_X1 U12165 ( .A1(n16947), .A2(n14254), .ZN(n16163) );
  OR2_X1 U12166 ( .A1(n19817), .A2(n10795), .ZN(n16941) );
  CLKBUF_X1 U12167 ( .A(n13573), .Z(n13574) );
  OR2_X1 U12168 ( .A1(n19853), .A2(n10735), .ZN(n16368) );
  AND3_X1 U12169 ( .A1(n11890), .A2(n11889), .A3(n11888), .ZN(n13501) );
  OR2_X1 U12170 ( .A1(n13402), .A2(n10064), .ZN(n13502) );
  INV_X1 U12171 ( .A(n10155), .ZN(n10154) );
  NAND2_X1 U12172 ( .A1(n9886), .A2(n10157), .ZN(n9883) );
  OAI21_X1 U12173 ( .B1(n10909), .B2(n11790), .A(n11984), .ZN(n10910) );
  NAND2_X1 U12174 ( .A1(n16198), .A2(n10936), .ZN(n10188) );
  NOR2_X1 U12175 ( .A1(n10004), .A2(n10003), .ZN(n10002) );
  INV_X1 U12176 ( .A(n13444), .ZN(n10003) );
  INV_X1 U12177 ( .A(n10005), .ZN(n10004) );
  AND3_X1 U12178 ( .A1(n11780), .A2(n11779), .A3(n11778), .ZN(n13702) );
  NAND2_X1 U12179 ( .A1(n9876), .A2(n9874), .ZN(n10368) );
  AND2_X1 U12180 ( .A1(n13428), .A2(n13427), .ZN(n13483) );
  AOI21_X1 U12181 ( .B1(n15888), .B2(n13419), .A(n13358), .ZN(n13363) );
  NAND2_X1 U12182 ( .A1(n13363), .A2(n13362), .ZN(n13428) );
  INV_X1 U12183 ( .A(n13132), .ZN(n13736) );
  INV_X1 U12184 ( .A(n20365), .ZN(n20363) );
  NAND2_X2 U12185 ( .A1(n10261), .A2(n10260), .ZN(n10325) );
  AND2_X1 U12186 ( .A1(n20701), .A2(n20727), .ZN(n20505) );
  INV_X1 U12187 ( .A(n20308), .ZN(n20555) );
  NOR2_X2 U12188 ( .A1(n14298), .A2(n13587), .ZN(n20118) );
  NAND2_X1 U12189 ( .A1(n10304), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10146) );
  NAND2_X1 U12190 ( .A1(n10305), .A2(n10291), .ZN(n10145) );
  INV_X1 U12191 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n13792) );
  INV_X1 U12192 ( .A(n14693), .ZN(n12757) );
  NOR2_X1 U12193 ( .A1(n17300), .A2(n17299), .ZN(n17298) );
  NOR2_X1 U12194 ( .A1(n17344), .A2(n18378), .ZN(n17343) );
  NOR2_X1 U12195 ( .A1(n17400), .A2(n17576), .ZN(n17389) );
  NAND2_X1 U12196 ( .A1(n17769), .A2(P3_EBX_REG_24__SCAN_IN), .ZN(n17756) );
  NAND2_X1 U12197 ( .A1(n17891), .A2(n9851), .ZN(n9852) );
  NOR2_X1 U12198 ( .A1(n17627), .A2(n17437), .ZN(n9851) );
  NOR2_X1 U12199 ( .A1(n12878), .A2(n12877), .ZN(n12879) );
  INV_X1 U12200 ( .A(n12875), .ZN(n12880) );
  AND2_X1 U12201 ( .A1(n17954), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n12877) );
  NOR2_X1 U12202 ( .A1(n19056), .A2(n18053), .ZN(n19516) );
  OAI211_X1 U12203 ( .C1(n17983), .C2(n17990), .A(n12694), .B(n12693), .ZN(
        n19700) );
  AOI211_X1 U12204 ( .C1(n17979), .C2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A(
        n12692), .B(n12691), .ZN(n12693) );
  NAND2_X1 U12205 ( .A1(n18355), .A2(n10039), .ZN(n17097) );
  NOR2_X1 U12206 ( .A1(n10041), .A2(n10042), .ZN(n10039) );
  NAND2_X1 U12207 ( .A1(n18355), .A2(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n18336) );
  NAND2_X1 U12208 ( .A1(n10030), .A2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n10029) );
  INV_X1 U12209 ( .A(n18410), .ZN(n10030) );
  AND2_X1 U12210 ( .A1(n17507), .A2(n10045), .ZN(n18526) );
  NAND2_X1 U12211 ( .A1(n17507), .A2(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n18554) );
  NAND2_X1 U12212 ( .A1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n18636) );
  OAI21_X1 U12213 ( .B1(n17092), .B2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n9902), .ZN(n9901) );
  AOI21_X1 U12214 ( .B1(n17093), .B2(n19661), .A(n9846), .ZN(n9902) );
  NOR2_X1 U12215 ( .A1(n17090), .A2(n18509), .ZN(n17092) );
  NAND2_X1 U12216 ( .A1(n17151), .A2(n17138), .ZN(n17093) );
  NOR2_X1 U12217 ( .A1(n18327), .A2(n16509), .ZN(n17126) );
  NOR2_X1 U12218 ( .A1(n16509), .A2(n17123), .ZN(n17124) );
  NAND2_X1 U12219 ( .A1(n18365), .A2(n18693), .ZN(n18327) );
  NOR2_X1 U12220 ( .A1(n12767), .A2(n12996), .ZN(n12994) );
  NOR2_X1 U12221 ( .A1(n18732), .A2(n18730), .ZN(n18365) );
  NAND2_X1 U12222 ( .A1(n18846), .A2(n18383), .ZN(n18732) );
  AOI21_X1 U12223 ( .B1(n18833), .B2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n12929), .ZN(n12930) );
  NOR2_X1 U12224 ( .A1(n12931), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12929) );
  INV_X1 U12225 ( .A(n18590), .ZN(n18575) );
  XNOR2_X1 U12226 ( .A(n9907), .B(n9906), .ZN(n18603) );
  INV_X1 U12227 ( .A(n12924), .ZN(n9906) );
  XNOR2_X1 U12228 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B(n12910), .ZN(
        n18613) );
  INV_X1 U12229 ( .A(n12895), .ZN(n10092) );
  INV_X1 U12230 ( .A(n17096), .ZN(n19484) );
  INV_X1 U12232 ( .A(n19505), .ZN(n19503) );
  NAND2_X1 U12233 ( .A1(n14692), .A2(n19711), .ZN(n19509) );
  NAND2_X1 U12234 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n19512) );
  NOR2_X1 U12235 ( .A1(n12663), .A2(n19512), .ZN(n19497) );
  INV_X1 U12236 ( .A(n19065), .ZN(n19388) );
  OR2_X1 U12237 ( .A1(n12736), .A2(n9860), .ZN(n9859) );
  INV_X1 U12238 ( .A(n12759), .ZN(n19048) );
  INV_X1 U12239 ( .A(n18143), .ZN(n19068) );
  OAI22_X1 U12240 ( .A1(n17096), .A2(n19483), .B1(n19480), .B2(n17149), .ZN(
        n19537) );
  CLKBUF_X1 U12241 ( .A(n13239), .Z(n14307) );
  CLKBUF_X1 U12242 ( .A(n12171), .Z(n12172) );
  INV_X1 U12243 ( .A(n14876), .ZN(n15595) );
  OR2_X1 U12244 ( .A1(n13391), .A2(n13390), .ZN(n15603) );
  OR2_X1 U12245 ( .A1(n15606), .A2(n13394), .ZN(n15605) );
  INV_X1 U12246 ( .A(n20894), .ZN(n20864) );
  INV_X1 U12247 ( .A(n20903), .ZN(n20869) );
  NOR2_X1 U12248 ( .A1(n20869), .A2(n21288), .ZN(n20894) );
  INV_X1 U12249 ( .A(n20864), .ZN(n20901) );
  OR2_X1 U12250 ( .A1(n12640), .A2(n15613), .ZN(n12641) );
  AOI21_X1 U12251 ( .B1(n15477), .B2(n9769), .A(n12534), .ZN(n16650) );
  NAND2_X1 U12252 ( .A1(n9957), .A2(n10113), .ZN(n15639) );
  INV_X1 U12253 ( .A(n16670), .ZN(n16734) );
  NOR2_X1 U12254 ( .A1(n16759), .A2(n9987), .ZN(n16751) );
  NOR2_X1 U12255 ( .A1(n15738), .A2(n9988), .ZN(n9987) );
  INV_X1 U12256 ( .A(n16763), .ZN(n9988) );
  NOR2_X1 U12257 ( .A1(n16774), .A2(n11581), .ZN(n16764) );
  AOI21_X1 U12258 ( .B1(n9986), .B2(n15763), .A(n15773), .ZN(n16786) );
  INV_X1 U12259 ( .A(n15738), .ZN(n9986) );
  OR2_X1 U12260 ( .A1(n9732), .A2(n16728), .ZN(n9918) );
  AND2_X1 U12261 ( .A1(n11679), .A2(n13303), .ZN(n15733) );
  AND2_X1 U12262 ( .A1(n11679), .A2(n11566), .ZN(n20934) );
  AND2_X1 U12263 ( .A1(n11679), .A2(n9997), .ZN(n20932) );
  INV_X1 U12264 ( .A(n12170), .ZN(n14398) );
  NAND2_X1 U12265 ( .A1(n11260), .A2(n11251), .ZN(n12177) );
  NOR2_X1 U12266 ( .A1(n20953), .A2(n13314), .ZN(n21268) );
  OAI21_X1 U12267 ( .B1(n14569), .B2(n20953), .A(n14541), .ZN(n14568) );
  INV_X1 U12268 ( .A(n21018), .ZN(n21050) );
  NAND2_X1 U12269 ( .A1(n16860), .A2(n16861), .ZN(n16859) );
  NAND2_X1 U12270 ( .A1(n16871), .A2(n16872), .ZN(n16870) );
  INV_X1 U12271 ( .A(n9936), .ZN(n13030) );
  NAND2_X1 U12272 ( .A1(n16894), .A2(n16895), .ZN(n16893) );
  NAND2_X1 U12273 ( .A1(n16903), .A2(n9718), .ZN(n15853) );
  NAND2_X1 U12274 ( .A1(n16904), .A2(n16905), .ZN(n16903) );
  AND2_X1 U12275 ( .A1(n13637), .A2(n13636), .ZN(n19960) );
  INV_X1 U12276 ( .A(n19959), .ZN(n16926) );
  INV_X1 U12277 ( .A(n20718), .ZN(n20074) );
  XNOR2_X1 U12278 ( .A(n15140), .B(n15139), .ZN(n15147) );
  OAI21_X1 U12279 ( .B1(n10055), .B2(n10053), .A(n10052), .ZN(n15140) );
  NAND2_X1 U12280 ( .A1(n10051), .A2(n15116), .ZN(n15891) );
  NAND2_X1 U12281 ( .A1(n10055), .A2(n10054), .ZN(n10051) );
  XNOR2_X1 U12282 ( .A(n15028), .B(n15027), .ZN(n15918) );
  AOI21_X1 U12283 ( .B1(n13367), .B2(n13366), .A(n17088), .ZN(n16020) );
  AND2_X1 U12284 ( .A1(n14308), .A2(n14298), .ZN(n16932) );
  AND2_X1 U12285 ( .A1(n16023), .A2(n19982), .ZN(n19988) );
  INV_X1 U12286 ( .A(n19982), .ZN(n16936) );
  OAI21_X1 U12287 ( .B1(n12097), .B2(n17048), .A(n12045), .ZN(n12046) );
  NOR2_X1 U12288 ( .A1(n12044), .A2(n10196), .ZN(n12045) );
  OR2_X1 U12289 ( .A1(n16281), .A2(n16280), .ZN(n16261) );
  INV_X1 U12290 ( .A(n16118), .ZN(n10152) );
  NAND2_X1 U12291 ( .A1(n10151), .A2(n16098), .ZN(n16115) );
  AND2_X1 U12292 ( .A1(n10160), .A2(n10711), .ZN(n16402) );
  AND2_X1 U12293 ( .A1(n10187), .A2(n10189), .ZN(n16197) );
  INV_X1 U12294 ( .A(n10905), .ZN(n10189) );
  INV_X1 U12295 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20710) );
  NAND2_X1 U12296 ( .A1(n13349), .A2(n13348), .ZN(n14878) );
  OAI21_X1 U12297 ( .B1(n13363), .B2(n13362), .A(n13428), .ZN(n20718) );
  AOI21_X1 U12298 ( .B1(n13773), .B2(n13412), .A(n13758), .ZN(n16437) );
  NOR2_X1 U12299 ( .A1(n13736), .A2(n20333), .ZN(n17082) );
  NOR2_X2 U12300 ( .A1(n20363), .A2(n20309), .ZN(n20182) );
  OR2_X1 U12301 ( .A1(n20165), .A2(n20551), .ZN(n20183) );
  INV_X1 U12302 ( .A(n20203), .ZN(n20213) );
  OAI21_X1 U12303 ( .B1(n20228), .B2(n20227), .A(n20226), .ZN(n20246) );
  INV_X1 U12304 ( .A(n20325), .ZN(n20327) );
  OR2_X1 U12305 ( .A1(n20303), .A2(n20302), .ZN(n20328) );
  OAI21_X1 U12306 ( .B1(n20357), .B2(n20336), .A(n20512), .ZN(n20359) );
  INV_X1 U12307 ( .A(n20395), .ZN(n20383) );
  OAI21_X1 U12308 ( .B1(n20405), .B2(n20420), .A(n20512), .ZN(n20423) );
  INV_X1 U12309 ( .A(n20386), .ZN(n20422) );
  INV_X1 U12310 ( .A(n20442), .ZN(n20445) );
  INV_X1 U12311 ( .A(n20537), .ZN(n20540) );
  OAI21_X1 U12312 ( .B1(n20518), .B2(n20517), .A(n20516), .ZN(n20541) );
  INV_X1 U12313 ( .A(n20521), .ZN(n20557) );
  INV_X1 U12314 ( .A(n20428), .ZN(n20561) );
  INV_X1 U12315 ( .A(n20433), .ZN(n20572) );
  NAND2_X1 U12316 ( .A1(n20505), .A2(n20555), .ZN(n20582) );
  INV_X1 U12317 ( .A(n20438), .ZN(n20586) );
  INV_X1 U12318 ( .A(n20582), .ZN(n20601) );
  INV_X1 U12319 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n20749) );
  INV_X1 U12320 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n20625) );
  AND3_X1 U12321 ( .A1(n20625), .A2(n20681), .A3(n20630), .ZN(n20756) );
  AOI21_X1 U12322 ( .B1(n19477), .B2(n19501), .A(n18204), .ZN(n19715) );
  OR2_X1 U12323 ( .A1(n17306), .A2(P3_EBX_REG_30__SCAN_IN), .ZN(n12791) );
  AND2_X1 U12324 ( .A1(n10025), .A2(n9842), .ZN(n13099) );
  AND2_X1 U12325 ( .A1(n10034), .A2(n9824), .ZN(n17351) );
  NOR2_X1 U12326 ( .A1(n17370), .A2(n18425), .ZN(n17369) );
  NOR2_X1 U12327 ( .A1(n18431), .A2(n17379), .ZN(n17378) );
  AND2_X1 U12328 ( .A1(n9843), .A2(n9778), .ZN(n17401) );
  NOR2_X2 U12329 ( .A1(n19538), .A2(n12784), .ZN(n17602) );
  INV_X1 U12330 ( .A(n17581), .ZN(n17619) );
  INV_X1 U12331 ( .A(n17586), .ZN(n17606) );
  NAND2_X1 U12332 ( .A1(n17759), .A2(P3_EBX_REG_26__SCAN_IN), .ZN(n17750) );
  NOR2_X1 U12333 ( .A1(n17756), .A2(n17737), .ZN(n17759) );
  NOR2_X1 U12334 ( .A1(n17765), .A2(n17736), .ZN(n17769) );
  NOR2_X1 U12335 ( .A1(n9754), .A2(n17830), .ZN(n17814) );
  NAND2_X1 U12336 ( .A1(P3_EBX_REG_19__SCAN_IN), .A2(n17846), .ZN(n17830) );
  INV_X1 U12337 ( .A(n17859), .ZN(n17832) );
  AND2_X1 U12338 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n17832), .ZN(n17846) );
  OR2_X1 U12339 ( .A1(n9852), .A2(n17412), .ZN(n17859) );
  NOR2_X1 U12340 ( .A1(n17909), .A2(n17905), .ZN(n17891) );
  NAND2_X1 U12341 ( .A1(n17891), .A2(P3_EBX_REG_15__SCAN_IN), .ZN(n17890) );
  NAND2_X1 U12342 ( .A1(n17927), .A2(P3_EBX_REG_13__SCAN_IN), .ZN(n17905) );
  AND2_X1 U12343 ( .A1(n17910), .A2(P3_EBX_REG_12__SCAN_IN), .ZN(n17927) );
  NOR2_X1 U12344 ( .A1(n18010), .A2(n18006), .ZN(n17987) );
  INV_X1 U12345 ( .A(n18048), .ZN(n18010) );
  INV_X2 U12346 ( .A(n18045), .ZN(n18039) );
  NAND2_X1 U12347 ( .A1(P3_EAX_REG_27__SCAN_IN), .A2(n18077), .ZN(n18073) );
  NOR2_X1 U12348 ( .A1(n18082), .A2(n18285), .ZN(n18077) );
  NAND2_X1 U12349 ( .A1(n18083), .A2(P3_EAX_REG_25__SCAN_IN), .ZN(n18082) );
  NOR3_X1 U12350 ( .A1(n18132), .A2(n18097), .A3(n18052), .ZN(n18093) );
  NOR2_X1 U12351 ( .A1(n9754), .A2(n18132), .ZN(n18126) );
  NAND2_X1 U12352 ( .A1(P3_EAX_REG_17__SCAN_IN), .A2(n18126), .ZN(n18125) );
  NOR2_X1 U12353 ( .A1(n18137), .A2(n18237), .ZN(n18133) );
  NAND2_X1 U12354 ( .A1(n18133), .A2(P3_EAX_REG_16__SCAN_IN), .ZN(n18132) );
  NOR2_X1 U12355 ( .A1(n18305), .A2(n18162), .ZN(n18158) );
  NOR2_X1 U12356 ( .A1(n18199), .A2(n18050), .ZN(n18051) );
  INV_X1 U12357 ( .A(n12980), .ZN(n18182) );
  NOR2_X1 U12358 ( .A1(n12844), .A2(n9893), .ZN(n9892) );
  AND2_X1 U12359 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(n18189), .ZN(n18194) );
  NAND2_X1 U12360 ( .A1(n16524), .A2(n18114), .ZN(n18195) );
  NOR2_X1 U12361 ( .A1(n12821), .A2(n12820), .ZN(n12827) );
  INV_X1 U12362 ( .A(n18269), .ZN(n18262) );
  BUF_X1 U12363 ( .A(n18289), .Z(n18318) );
  OR2_X1 U12364 ( .A1(n18332), .A2(n18331), .ZN(n18333) );
  NOR3_X1 U12365 ( .A1(n18446), .A2(n10031), .A3(n18410), .ZN(n18394) );
  NOR2_X1 U12366 ( .A1(n18586), .A2(n18811), .ZN(n18426) );
  NOR2_X1 U12367 ( .A1(n18446), .A2(n18447), .ZN(n18437) );
  NAND2_X1 U12368 ( .A1(n18630), .A2(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n18618) );
  INV_X1 U12369 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n18619) );
  NOR2_X1 U12370 ( .A1(n18636), .A2(n18650), .ZN(n18630) );
  INV_X1 U12371 ( .A(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n18650) );
  NAND2_X1 U12372 ( .A1(n18684), .A2(n19023), .ZN(n18677) );
  NOR2_X1 U12373 ( .A1(n17101), .A2(n17269), .ZN(n18674) );
  OAI21_X2 U12374 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n19693), .A(n17269), 
        .ZN(n18684) );
  INV_X1 U12375 ( .A(n18678), .ZN(n18687) );
  INV_X1 U12376 ( .A(n18674), .ZN(n18689) );
  XNOR2_X1 U12377 ( .A(n10097), .B(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n17119) );
  NAND2_X1 U12378 ( .A1(n17093), .A2(n10098), .ZN(n10097) );
  NAND2_X1 U12379 ( .A1(n17090), .A2(n12931), .ZN(n10098) );
  NAND2_X1 U12380 ( .A1(n10099), .A2(n18433), .ZN(n18385) );
  NOR2_X1 U12381 ( .A1(n18645), .A2(n18644), .ZN(n18643) );
  AND2_X1 U12382 ( .A1(n9905), .A2(n12863), .ZN(n18645) );
  INV_X1 U12383 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19527) );
  CLKBUF_X1 U12384 ( .A(n17255), .Z(n17253) );
  AND2_X1 U12385 ( .A1(n11196), .A2(n12132), .ZN(n13258) );
  AOI21_X1 U12386 ( .B1(n15161), .B2(n15162), .A(n10127), .ZN(n10126) );
  OAI21_X1 U12387 ( .B1(n15549), .B2(n16617), .A(n10128), .ZN(n10127) );
  OAI21_X1 U12388 ( .B1(n15699), .B2(n20773), .A(n9955), .ZN(P1_U2971) );
  NOR2_X1 U12389 ( .A1(n9794), .A2(n9956), .ZN(n9955) );
  INV_X1 U12390 ( .A(n13026), .ZN(n9956) );
  AOI211_X1 U12391 ( .C1(n14825), .C2(n16809), .A(n14824), .B(n14823), .ZN(
        n14829) );
  NAND2_X1 U12392 ( .A1(n9994), .A2(n9993), .ZN(P1_U3001) );
  AOI211_X1 U12393 ( .C1(n14827), .C2(n12136), .A(n12137), .B(n15615), .ZN(
        n9993) );
  AND2_X1 U12394 ( .A1(n13070), .A2(n13069), .ZN(n13071) );
  AND2_X1 U12395 ( .A1(n11682), .A2(n11681), .ZN(n11683) );
  INV_X1 U12396 ( .A(n19932), .ZN(n10076) );
  NOR2_X1 U12397 ( .A1(n14788), .A2(n10057), .ZN(n14789) );
  OR2_X1 U12398 ( .A1(n14787), .A2(n9830), .ZN(n10057) );
  NOR2_X1 U12399 ( .A1(n14768), .A2(n10056), .ZN(n14769) );
  AND2_X1 U12400 ( .A1(n19969), .A2(n13412), .ZN(n10056) );
  NAND2_X1 U12401 ( .A1(n9998), .A2(n11041), .ZN(n9966) );
  INV_X1 U12402 ( .A(n10194), .ZN(n10193) );
  OAI21_X1 U12403 ( .B1(n14846), .B2(n20043), .A(n10195), .ZN(n10194) );
  AOI21_X1 U12404 ( .B1(n16869), .B2(n20051), .A(n14847), .ZN(n10195) );
  AND2_X1 U12405 ( .A1(n20051), .A2(n13412), .ZN(n10058) );
  AOI211_X1 U12406 ( .C1(n20057), .C2(n15144), .A(n12025), .B(n12024), .ZN(
        n12026) );
  AOI21_X1 U12407 ( .B1(n14813), .B2(n17052), .A(n10067), .ZN(n14814) );
  OAI211_X1 U12408 ( .C1(n16867), .C2(n17048), .A(n10071), .B(n10068), .ZN(
        n10067) );
  OAI21_X1 U12409 ( .B1(n14798), .B2(n20068), .A(n13043), .ZN(n13044) );
  NAND2_X1 U12410 ( .A1(n17074), .A2(n13412), .ZN(n17058) );
  OR2_X1 U12411 ( .A1(n17586), .A2(n12659), .ZN(n10024) );
  INV_X1 U12412 ( .A(n17910), .ZN(n17941) );
  NAND2_X1 U12413 ( .A1(n18060), .A2(n9861), .ZN(n18054) );
  INV_X1 U12414 ( .A(n18083), .ZN(n18087) );
  OAI21_X1 U12415 ( .B1(n17148), .B2(n18877), .A(n9899), .ZN(P3_U2831) );
  AND2_X1 U12416 ( .A1(n17146), .A2(n17147), .ZN(n9899) );
  NAND2_X2 U12417 ( .A1(n12662), .A2(n12672), .ZN(n17913) );
  NAND2_X1 U12418 ( .A1(n12446), .A2(n10176), .ZN(n9769) );
  NAND2_X1 U12419 ( .A1(n9867), .A2(n9865), .ZN(n10326) );
  INV_X2 U12420 ( .A(n10326), .ZN(n10306) );
  OR2_X2 U12421 ( .A1(n19656), .A2(n12665), .ZN(n10201) );
  AND2_X2 U12422 ( .A1(n10556), .A2(n10555), .ZN(n11790) );
  OR3_X1 U12423 ( .A1(n18446), .A2(n10031), .A3(n10029), .ZN(n9770) );
  NOR2_X1 U12424 ( .A1(n10727), .A2(n10721), .ZN(n9771) );
  AND2_X1 U12425 ( .A1(n12446), .A2(n10177), .ZN(n15483) );
  NAND2_X1 U12426 ( .A1(n10167), .A2(n13995), .ZN(n13989) );
  INV_X1 U12427 ( .A(n16673), .ZN(n16645) );
  AND2_X1 U12428 ( .A1(n14664), .A2(n10180), .ZN(n9772) );
  AND2_X1 U12429 ( .A1(n10082), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n9773) );
  XNOR2_X1 U12430 ( .A(n13434), .B(n13435), .ZN(n13511) );
  NAND2_X1 U12431 ( .A1(n12446), .A2(n12445), .ZN(n15490) );
  AND2_X1 U12432 ( .A1(n13828), .A2(n9829), .ZN(n14579) );
  AND2_X1 U12433 ( .A1(n14299), .A2(n13436), .ZN(n9775) );
  INV_X1 U12434 ( .A(n10178), .ZN(n15428) );
  OR2_X1 U12435 ( .A1(n10096), .A2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n9776) );
  AND2_X1 U12436 ( .A1(n13637), .A2(n9823), .ZN(n14903) );
  AND2_X1 U12437 ( .A1(n10838), .A2(n10738), .ZN(n9777) );
  INV_X1 U12438 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n9954) );
  NAND2_X1 U12439 ( .A1(n17419), .A2(n17406), .ZN(n9778) );
  INV_X2 U12440 ( .A(n14928), .ZN(n10445) );
  NOR2_X1 U12441 ( .A1(n15504), .A2(n10139), .ZN(n9779) );
  AND2_X1 U12442 ( .A1(n10134), .A2(n14710), .ZN(n9780) );
  AND2_X1 U12443 ( .A1(n10079), .A2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n9781) );
  AND2_X1 U12444 ( .A1(n12938), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n9782) );
  NAND2_X2 U12445 ( .A1(n20765), .A2(P2_STATE_REG_2__SCAN_IN), .ZN(n20681) );
  INV_X4 U12446 ( .A(n17879), .ZN(n12839) );
  INV_X1 U12447 ( .A(n10306), .ZN(n10561) );
  NAND2_X1 U12448 ( .A1(n15856), .A2(n10021), .ZN(n13036) );
  OR2_X1 U12449 ( .A1(n14748), .A2(n9965), .ZN(n16053) );
  AND4_X1 U12450 ( .A1(n11056), .A2(n11055), .A3(n11054), .A4(n11053), .ZN(
        n9783) );
  AND3_X1 U12451 ( .A1(n10930), .A2(n14267), .A3(n10002), .ZN(n9784) );
  XOR2_X1 U12452 ( .A(n13062), .B(n13061), .Z(n9785) );
  OR2_X1 U12453 ( .A1(n15927), .A2(n15004), .ZN(n9786) );
  NAND2_X1 U12454 ( .A1(n10325), .A2(n20098), .ZN(n11715) );
  NAND2_X1 U12455 ( .A1(n13418), .A2(n13417), .ZN(n13434) );
  AND2_X1 U12456 ( .A1(n15858), .A2(n15837), .ZN(n15836) );
  NAND2_X1 U12457 ( .A1(n14664), .A2(n9828), .ZN(n10178) );
  AND2_X1 U12458 ( .A1(n15858), .A2(n10073), .ZN(n13038) );
  INV_X1 U12459 ( .A(n15180), .ZN(n12534) );
  NAND2_X1 U12460 ( .A1(n11057), .A2(n9783), .ZN(n11487) );
  NAND2_X1 U12461 ( .A1(n13412), .A2(n13420), .ZN(n10420) );
  XNOR2_X1 U12462 ( .A(n12041), .B(n12040), .ZN(n12097) );
  AND2_X1 U12463 ( .A1(n15478), .A2(n10134), .ZN(n9788) );
  OR2_X1 U12464 ( .A1(n16845), .A2(n20062), .ZN(n9789) );
  NAND2_X1 U12465 ( .A1(n10160), .A2(n10159), .ZN(n16401) );
  AND2_X2 U12466 ( .A1(n10230), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10448) );
  NOR2_X1 U12467 ( .A1(n16053), .A2(n10191), .ZN(n9790) );
  AND3_X1 U12468 ( .A1(n10276), .A2(n10291), .A3(n10275), .ZN(n9791) );
  INV_X1 U12469 ( .A(n10430), .ZN(n15873) );
  NOR2_X1 U12470 ( .A1(n14748), .A2(n9963), .ZN(n9792) );
  INV_X1 U12471 ( .A(n13468), .ZN(n10007) );
  AND2_X1 U12472 ( .A1(n11384), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n9793) );
  NOR2_X1 U12473 ( .A1(n14731), .A2(n16700), .ZN(n9794) );
  AND2_X1 U12474 ( .A1(n10232), .A2(n10291), .ZN(n9795) );
  INV_X1 U12475 ( .A(n9964), .ZN(n16065) );
  OR2_X1 U12476 ( .A1(n14748), .A2(n16262), .ZN(n9964) );
  NAND2_X1 U12477 ( .A1(n10802), .A2(n9937), .ZN(n9796) );
  NAND2_X1 U12478 ( .A1(n10149), .A2(n10147), .ZN(n10153) );
  OR2_X1 U12479 ( .A1(n11442), .A2(n11309), .ZN(n9797) );
  INV_X1 U12480 ( .A(n16508), .ZN(n17158) );
  XNOR2_X1 U12481 ( .A(n13431), .B(n13429), .ZN(n13482) );
  AND3_X1 U12482 ( .A1(n12749), .A2(n9855), .A3(n9854), .ZN(n9798) );
  OR2_X1 U12483 ( .A1(n10918), .A2(n10917), .ZN(n9799) );
  NAND2_X1 U12484 ( .A1(n13433), .A2(n13432), .ZN(n13512) );
  AND2_X1 U12485 ( .A1(n12836), .A2(n12835), .ZN(n9800) );
  INV_X1 U12486 ( .A(n17610), .ZN(n12662) );
  NAND2_X1 U12487 ( .A1(n10694), .A2(n10693), .ZN(n10877) );
  AND2_X1 U12488 ( .A1(n15629), .A2(n16673), .ZN(n9801) );
  AND2_X1 U12489 ( .A1(n14800), .A2(n14799), .ZN(n9802) );
  OR2_X1 U12490 ( .A1(n18967), .A2(n12881), .ZN(n9803) );
  NOR2_X1 U12491 ( .A1(n12814), .A2(n12813), .ZN(n9804) );
  AND2_X1 U12492 ( .A1(n11572), .A2(n11571), .ZN(n15784) );
  AND2_X1 U12493 ( .A1(n12939), .A2(n12938), .ZN(n9805) );
  NAND2_X1 U12494 ( .A1(n10903), .A2(n10902), .ZN(n14384) );
  INV_X1 U12495 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10573) );
  AND2_X1 U12496 ( .A1(n14241), .A2(n16387), .ZN(n13640) );
  NOR2_X1 U12497 ( .A1(n18446), .A2(n10031), .ZN(n9806) );
  NAND2_X1 U12498 ( .A1(n14563), .A2(n12256), .ZN(n14664) );
  NAND2_X1 U12499 ( .A1(n9885), .A2(n10703), .ZN(n16179) );
  NOR2_X1 U12500 ( .A1(n16099), .A2(n10150), .ZN(n9807) );
  AND2_X1 U12501 ( .A1(n13827), .A2(n13830), .ZN(n13828) );
  AND2_X1 U12502 ( .A1(n13828), .A2(n14303), .ZN(n14302) );
  AND2_X1 U12503 ( .A1(n13828), .A2(n10066), .ZN(n14371) );
  NOR2_X1 U12504 ( .A1(n16021), .A2(n16008), .ZN(n16000) );
  NAND2_X1 U12505 ( .A1(n14664), .A2(n12285), .ZN(n14663) );
  NOR2_X1 U12506 ( .A1(n14284), .A2(n14240), .ZN(n14241) );
  AND2_X1 U12507 ( .A1(n13721), .A2(n13818), .ZN(n13819) );
  AND3_X1 U12508 ( .A1(n13995), .A2(n10174), .A3(n13819), .ZN(n13988) );
  NOR2_X1 U12509 ( .A1(n13573), .A2(n16355), .ZN(n13827) );
  NAND2_X1 U12510 ( .A1(n13637), .A2(n10062), .ZN(n14481) );
  NAND2_X1 U12511 ( .A1(n15540), .A2(n15531), .ZN(n15431) );
  NOR2_X1 U12512 ( .A1(n13402), .A2(n13403), .ZN(n9808) );
  NAND2_X1 U12513 ( .A1(n14435), .A2(n10013), .ZN(n14749) );
  AND2_X1 U12514 ( .A1(n12070), .A2(n10082), .ZN(n9809) );
  AND2_X1 U12515 ( .A1(n10183), .A2(n13016), .ZN(n9810) );
  NAND2_X1 U12516 ( .A1(n13640), .A2(n10010), .ZN(n13714) );
  NAND2_X1 U12517 ( .A1(n18575), .A2(n12928), .ZN(n18519) );
  OR2_X1 U12518 ( .A1(n10064), .A2(n13501), .ZN(n9811) );
  NAND2_X1 U12519 ( .A1(n10112), .A2(n11362), .ZN(n13832) );
  AND2_X1 U12520 ( .A1(n15496), .A2(n15485), .ZN(n15478) );
  NAND2_X1 U12521 ( .A1(n9918), .A2(n16729), .ZN(n14351) );
  AND2_X1 U12522 ( .A1(n16163), .A2(n16162), .ZN(n14129) );
  AND2_X1 U12523 ( .A1(n14785), .A2(n17065), .ZN(n9812) );
  NAND2_X1 U12524 ( .A1(n16581), .A2(n9779), .ZN(n15493) );
  AND2_X1 U12525 ( .A1(n20850), .A2(P1_EBX_REG_30__SCAN_IN), .ZN(n9813) );
  AND2_X1 U12526 ( .A1(n11377), .A2(n11363), .ZN(n9814) );
  INV_X1 U12527 ( .A(n11442), .ZN(n10164) );
  AND2_X1 U12528 ( .A1(n13625), .A2(n13720), .ZN(n13721) );
  OR2_X1 U12529 ( .A1(n18590), .A2(n9776), .ZN(n18510) );
  OR2_X1 U12530 ( .A1(n10718), .A2(n10838), .ZN(n10824) );
  NOR2_X1 U12531 ( .A1(n17343), .A2(n17576), .ZN(n9815) );
  AND2_X1 U12532 ( .A1(n9814), .A2(n11399), .ZN(n9816) );
  INV_X1 U12533 ( .A(n14436), .ZN(n10989) );
  INV_X1 U12534 ( .A(n10041), .ZN(n10040) );
  AND2_X1 U12535 ( .A1(n11524), .A2(n11495), .ZN(n9817) );
  INV_X1 U12536 ( .A(n15182), .ZN(n12533) );
  AND2_X1 U12537 ( .A1(n10170), .A2(n13995), .ZN(n12254) );
  AND2_X1 U12538 ( .A1(n10599), .A2(n10598), .ZN(n11777) );
  NAND2_X1 U12539 ( .A1(n10075), .A2(n11963), .ZN(n15975) );
  OR2_X1 U12540 ( .A1(n11426), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n9818) );
  AND2_X1 U12541 ( .A1(n15856), .A2(n15846), .ZN(n15845) );
  AND2_X1 U12542 ( .A1(n14435), .A2(n10015), .ZN(n9819) );
  AND2_X1 U12543 ( .A1(n16098), .A2(n16100), .ZN(n9820) );
  AND2_X1 U12544 ( .A1(n11192), .A2(n10124), .ZN(n9821) );
  NOR2_X1 U12545 ( .A1(n13402), .A2(n9811), .ZN(n9822) );
  AND2_X1 U12546 ( .A1(n10062), .A2(n10061), .ZN(n9823) );
  AND2_X1 U12547 ( .A1(n10035), .A2(n10033), .ZN(n9824) );
  AND2_X1 U12548 ( .A1(n9810), .A2(n10182), .ZN(n9825) );
  OR2_X1 U12549 ( .A1(n9811), .A2(n10063), .ZN(n9826) );
  INV_X2 U12550 ( .A(n14992), .ZN(n10462) );
  INV_X1 U12551 ( .A(n11790), .ZN(n10826) );
  AND2_X1 U12552 ( .A1(n12084), .A2(n9781), .ZN(n9827) );
  INV_X1 U12553 ( .A(n14744), .ZN(n9997) );
  AND2_X1 U12554 ( .A1(n14857), .A2(n14856), .ZN(n14267) );
  INV_X1 U12555 ( .A(n10803), .ZN(n9941) );
  INV_X1 U12556 ( .A(n10763), .ZN(n9945) );
  AND2_X1 U12557 ( .A1(n10180), .A2(n15535), .ZN(n9828) );
  AND2_X1 U12558 ( .A1(n10066), .A2(n14580), .ZN(n9829) );
  INV_X1 U12559 ( .A(n9882), .ZN(n13365) );
  NAND2_X1 U12560 ( .A1(n12084), .A2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n12058) );
  AND2_X1 U12561 ( .A1(n13412), .A2(n19922), .ZN(n9830) );
  NOR2_X1 U12562 ( .A1(n17369), .A2(n17576), .ZN(n9831) );
  OR3_X1 U12563 ( .A1(n12074), .A2(n10086), .A3(n10085), .ZN(n9832) );
  AND2_X1 U12564 ( .A1(n9829), .A2(n16022), .ZN(n9833) );
  INV_X1 U12565 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n10124) );
  NOR2_X1 U12566 ( .A1(n15119), .A2(n15118), .ZN(n9834) );
  AND2_X1 U12567 ( .A1(n13142), .A2(n11996), .ZN(n9835) );
  NOR2_X1 U12568 ( .A1(n14121), .A2(n10142), .ZN(n9836) );
  AND3_X1 U12569 ( .A1(n10930), .A2(n14267), .A3(n10005), .ZN(n9837) );
  AND3_X1 U12570 ( .A1(n10930), .A2(n14267), .A3(n10007), .ZN(n9838) );
  AND2_X1 U12571 ( .A1(n10073), .A2(n13040), .ZN(n9839) );
  AND2_X1 U12572 ( .A1(n15494), .A2(n15502), .ZN(n9840) );
  NOR2_X1 U12573 ( .A1(n14778), .A2(n10058), .ZN(n9841) );
  AND2_X1 U12574 ( .A1(n10026), .A2(n10033), .ZN(n9842) );
  XOR2_X1 U12575 ( .A(n12660), .B(n12659), .Z(n9843) );
  INV_X1 U12576 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n10085) );
  NOR2_X1 U12577 ( .A1(n17097), .A2(n17615), .ZN(n12658) );
  NAND2_X1 U12578 ( .A1(n13299), .A2(n14703), .ZN(n11548) );
  INV_X1 U12579 ( .A(n13992), .ZN(n10143) );
  AND4_X1 U12580 ( .A1(P3_EAX_REG_14__SCAN_IN), .A2(P3_EAX_REG_11__SCAN_IN), 
        .A3(P3_EAX_REG_10__SCAN_IN), .A4(P3_EAX_REG_9__SCAN_IN), .ZN(n9844) );
  NOR2_X1 U12581 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n18520), .ZN(
        n9845) );
  AND2_X1 U12582 ( .A1(n18509), .A2(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n9846) );
  INV_X1 U12583 ( .A(n13458), .ZN(n11597) );
  INV_X1 U12584 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n9947) );
  INV_X1 U12585 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n10080) );
  INV_X1 U12586 ( .A(n18378), .ZN(n10028) );
  INV_X1 U12587 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n10042) );
  AND2_X1 U12588 ( .A1(n12119), .A2(n12118), .ZN(n9847) );
  NOR2_X1 U12589 ( .A1(n18618), .A2(n18619), .ZN(n17507) );
  AND2_X1 U12590 ( .A1(n18355), .A2(n10040), .ZN(n9848) );
  NAND2_X1 U12591 ( .A1(n15726), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n9849) );
  INV_X1 U12592 ( .A(P2_EBX_REG_23__SCAN_IN), .ZN(n9940) );
  INV_X1 U12593 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n10095) );
  INV_X1 U12594 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n9980) );
  INV_X1 U12595 ( .A(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n10091) );
  INV_X1 U12596 ( .A(n15690), .ZN(n9914) );
  AND2_X1 U12597 ( .A1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n9850) );
  NAND3_X2 U12598 ( .A1(n19713), .A2(n19542), .A3(n19712), .ZN(n19013) );
  AND2_X1 U12599 ( .A1(n13953), .A2(n13952), .ZN(n16609) );
  OAI22_X2 U12600 ( .A1(n20103), .A2(n20111), .B1(n20102), .B2(n20113), .ZN(
        n20492) );
  NOR3_X2 U12601 ( .A1(n19417), .A2(n19522), .A3(n19118), .ZN(n19134) );
  NOR2_X2 U12602 ( .A1(n13592), .A2(n20120), .ZN(n20548) );
  OAI21_X1 U12603 ( .B1(n15160), .B2(n20860), .A(n10126), .ZN(P1_U2810) );
  OAI211_X1 U12604 ( .C1(n12036), .C2(n17071), .A(n12026), .B(n10072), .ZN(
        P2_U3016) );
  AOI22_X2 U12605 ( .A1(BUF2_REG_17__SCAN_IN), .A2(n20118), .B1(
        BUF1_REG_17__SCAN_IN), .B2(n20119), .ZN(n20564) );
  NOR2_X2 U12606 ( .A1(n14307), .A2(n13587), .ZN(n20119) );
  NOR2_X2 U12607 ( .A1(n19059), .A2(n19354), .ZN(n19461) );
  OR2_X1 U12608 ( .A1(n11677), .A2(n9954), .ZN(n11277) );
  NOR4_X4 U12609 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(P3_STATE2_REG_0__SCAN_IN), .A3(P3_STATEBS16_REG_SCAN_IN), .A4(n19660), .ZN(n17608) );
  NOR2_X2 U12610 ( .A1(n20121), .A2(n20120), .ZN(n20596) );
  NOR2_X2 U12611 ( .A1(n11994), .A2(n20120), .ZN(n20576) );
  NAND2_X1 U12612 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n20512), .ZN(n20120) );
  INV_X1 U12613 ( .A(n9852), .ZN(n17875) );
  NAND3_X1 U12614 ( .A1(n12750), .A2(n12748), .A3(n9798), .ZN(n9853) );
  INV_X2 U12615 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n12663) );
  NOR2_X2 U12616 ( .A1(n16522), .A2(n9857), .ZN(n18048) );
  NOR2_X2 U12617 ( .A1(n12735), .A2(n9859), .ZN(n19044) );
  INV_X2 U12618 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n19666) );
  INV_X2 U12619 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n19674) );
  NAND2_X1 U12620 ( .A1(n9864), .A2(n10919), .ZN(n10000) );
  XNOR2_X2 U12621 ( .A(n9864), .B(n10919), .ZN(n10435) );
  NAND2_X2 U12622 ( .A1(n10001), .A2(n10388), .ZN(n9864) );
  NAND4_X1 U12623 ( .A1(n9866), .A2(n10293), .A3(n10294), .A4(n10292), .ZN(
        n9865) );
  NAND4_X1 U12624 ( .A1(n9868), .A2(n10287), .A3(n10288), .A4(n10289), .ZN(
        n9867) );
  NAND2_X1 U12625 ( .A1(n20032), .A2(n20030), .ZN(n10607) );
  NAND2_X1 U12626 ( .A1(n9873), .A2(n10582), .ZN(n20032) );
  NAND3_X1 U12627 ( .A1(n9878), .A2(n9879), .A3(n10363), .ZN(n9875) );
  NAND2_X1 U12628 ( .A1(n10364), .A2(n10362), .ZN(n9876) );
  NAND2_X1 U12629 ( .A1(n9877), .A2(n10362), .ZN(n10382) );
  NAND2_X1 U12630 ( .A1(n10345), .A2(n10344), .ZN(n9879) );
  NAND2_X1 U12631 ( .A1(n9882), .A2(n20098), .ZN(n9880) );
  NOR2_X1 U12632 ( .A1(n9882), .A2(n11715), .ZN(n10351) );
  MUX2_X1 U12633 ( .A(n11692), .B(n11992), .S(n9882), .Z(n11993) );
  NAND2_X1 U12634 ( .A1(n13772), .A2(n9882), .ZN(n12002) );
  NAND3_X1 U12635 ( .A1(n9884), .A2(n10154), .A3(n9883), .ZN(n16378) );
  NAND3_X1 U12636 ( .A1(n14382), .A2(n14381), .A3(n10157), .ZN(n9884) );
  NAND3_X2 U12637 ( .A1(n9887), .A2(n10442), .A3(n10443), .ZN(n10471) );
  NAND4_X1 U12638 ( .A1(n10492), .A2(n10490), .A3(n10489), .A4(n10491), .ZN(
        n10538) );
  NAND2_X1 U12639 ( .A1(n10471), .A2(n10470), .ZN(n9888) );
  NAND2_X1 U12640 ( .A1(n10538), .A2(n10537), .ZN(n9889) );
  OR2_X2 U12641 ( .A1(n16041), .A2(n10827), .ZN(n9890) );
  NOR2_X1 U12642 ( .A1(n9898), .A2(n9897), .ZN(n9896) );
  NAND2_X1 U12643 ( .A1(n12808), .A2(n12809), .ZN(n9897) );
  OAI21_X1 U12644 ( .B1(n18644), .B2(n12863), .A(n9803), .ZN(n9904) );
  INV_X1 U12645 ( .A(n9905), .ZN(n18651) );
  NOR2_X1 U12646 ( .A1(n18614), .A2(n18613), .ZN(n18612) );
  NAND2_X1 U12647 ( .A1(n9805), .A2(n18352), .ZN(n9908) );
  INV_X1 U12648 ( .A(n18354), .ZN(n9909) );
  NOR2_X2 U12649 ( .A1(n18418), .A2(n18705), .ZN(n18735) );
  NAND3_X1 U12650 ( .A1(n12662), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(
        n19656), .ZN(n12797) );
  AND2_X4 U12651 ( .A1(n11044), .A2(n13305), .ZN(n12606) );
  AND2_X4 U12652 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13305) );
  INV_X1 U12653 ( .A(n12116), .ZN(n9910) );
  NAND2_X1 U12654 ( .A1(n9910), .A2(n9981), .ZN(n9911) );
  OAI211_X1 U12655 ( .C1(n12117), .C2(n9912), .A(n16673), .B(n9911), .ZN(n9915) );
  NAND2_X1 U12656 ( .A1(n9916), .A2(n9981), .ZN(n12138) );
  INV_X1 U12657 ( .A(n9916), .ZN(n12139) );
  OR2_X2 U12658 ( .A1(n9916), .A2(n9914), .ZN(n9913) );
  NAND2_X1 U12659 ( .A1(n20978), .A2(n11267), .ZN(n14001) );
  NAND2_X2 U12660 ( .A1(n15675), .A2(n11428), .ZN(n15663) );
  OR2_X2 U12661 ( .A1(n14645), .A2(n11427), .ZN(n15675) );
  NAND2_X1 U12662 ( .A1(n16735), .A2(n16737), .ZN(n11409) );
  NAND2_X1 U12663 ( .A1(n9925), .A2(n9923), .ZN(n16735) );
  INV_X1 U12664 ( .A(n11362), .ZN(n9924) );
  NAND3_X1 U12665 ( .A1(n13729), .A2(n13833), .A3(n13730), .ZN(n9925) );
  XNOR2_X1 U12666 ( .A(n11314), .B(n11590), .ZN(n13456) );
  NAND2_X1 U12667 ( .A1(n11313), .A2(n9929), .ZN(n9928) );
  INV_X1 U12668 ( .A(n13476), .ZN(n9929) );
  NAND2_X1 U12669 ( .A1(n13449), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n9930) );
  INV_X2 U12670 ( .A(n11487), .ZN(n13880) );
  AOI21_X2 U12671 ( .B1(n16032), .B2(n16028), .A(n16030), .ZN(n11685) );
  NAND2_X1 U12672 ( .A1(n11487), .A2(n11553), .ZN(n9950) );
  NAND3_X1 U12673 ( .A1(n10166), .A2(n12171), .A3(n11307), .ZN(n10165) );
  XNOR2_X2 U12674 ( .A(n11254), .B(n11252), .ZN(n12171) );
  NAND2_X1 U12675 ( .A1(n11268), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n9952) );
  AND2_X4 U12676 ( .A1(n11411), .A2(n9958), .ZN(n16673) );
  NAND4_X1 U12677 ( .A1(n10234), .A2(n9795), .A3(n10231), .A4(n10233), .ZN(
        n9962) );
  NAND4_X1 U12678 ( .A1(n10538), .A2(n10471), .A3(n10537), .A4(n10470), .ZN(
        n10878) );
  NAND4_X1 U12679 ( .A1(n10538), .A2(n10471), .A3(n10537), .A4(n9968), .ZN(
        n10656) );
  XNOR2_X1 U12680 ( .A(n10909), .B(n11790), .ZN(n16198) );
  NAND2_X2 U12681 ( .A1(n9970), .A2(n10695), .ZN(n10909) );
  NAND2_X1 U12682 ( .A1(n11409), .A2(n16736), .ZN(n16727) );
  NOR2_X2 U12683 ( .A1(n11335), .A2(n14088), .ZN(n11364) );
  INV_X2 U12684 ( .A(n9974), .ZN(n11158) );
  NAND4_X1 U12685 ( .A1(n13316), .A2(n14745), .A3(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A4(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n9974) );
  AND2_X2 U12686 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11052) );
  NAND2_X1 U12687 ( .A1(n11158), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n9976) );
  AND2_X2 U12688 ( .A1(n11050), .A2(n11051), .ZN(n11159) );
  NOR2_X2 U12689 ( .A1(n15627), .A2(n9979), .ZN(n9981) );
  XNOR2_X1 U12690 ( .A(n11384), .B(n11383), .ZN(n13833) );
  OAI21_X2 U12691 ( .B1(n15663), .B2(n11458), .A(n11457), .ZN(n15660) );
  NAND2_X1 U12692 ( .A1(n11025), .A2(n11731), .ZN(n9999) );
  NAND3_X1 U12693 ( .A1(n17296), .A2(n17297), .A3(n10024), .ZN(P3_U2640) );
  NAND2_X1 U12694 ( .A1(n10025), .A2(n10026), .ZN(n17330) );
  NAND2_X1 U12695 ( .A1(n10034), .A2(n10035), .ZN(n17363) );
  INV_X1 U12696 ( .A(n17576), .ZN(n10033) );
  NAND3_X1 U12697 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n10041) );
  INV_X2 U12698 ( .A(n9843), .ZN(n17576) );
  NAND3_X1 U12699 ( .A1(n17507), .A2(n10212), .A3(n10045), .ZN(n18482) );
  INV_X2 U12700 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10291) );
  AND3_X2 U12701 ( .A1(n10047), .A2(n10307), .A3(n10308), .ZN(n13141) );
  INV_X1 U12702 ( .A(n10337), .ZN(n10047) );
  NAND2_X1 U12703 ( .A1(n10347), .A2(n10047), .ZN(n10861) );
  INV_X2 U12704 ( .A(n10920), .ZN(n10392) );
  NAND2_X2 U12705 ( .A1(n10048), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10920) );
  NAND2_X1 U12706 ( .A1(n10373), .A2(n11730), .ZN(n10049) );
  INV_X1 U12707 ( .A(n15899), .ZN(n10054) );
  INV_X1 U12708 ( .A(n10055), .ZN(n15904) );
  XNOR2_X1 U12709 ( .A(n15078), .B(n15077), .ZN(n15906) );
  OR2_X2 U12710 ( .A1(n13402), .A2(n9826), .ZN(n13573) );
  NAND2_X4 U12711 ( .A1(n10324), .A2(n10323), .ZN(n20755) );
  OR2_X1 U12712 ( .A1(n11748), .A2(n11953), .ZN(n11751) );
  NAND2_X1 U12713 ( .A1(n15858), .A2(n9839), .ZN(n13039) );
  INV_X1 U12714 ( .A(n13039), .ZN(n11976) );
  NAND2_X1 U12716 ( .A1(n10077), .A2(n10076), .ZN(n12113) );
  NAND2_X1 U12717 ( .A1(n16859), .A2(n9719), .ZN(n16848) );
  NOR2_X1 U12718 ( .A1(n18590), .A2(n10096), .ZN(n18498) );
  NAND3_X1 U12719 ( .A1(n10099), .A2(n18433), .A3(n18730), .ZN(n18374) );
  AND2_X4 U12720 ( .A1(n15828), .A2(n11052), .ZN(n12612) );
  INV_X1 U12721 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10100) );
  NAND2_X1 U12722 ( .A1(n10102), .A2(n10101), .ZN(n10106) );
  INV_X1 U12723 ( .A(n12171), .ZN(n10102) );
  NAND3_X1 U12724 ( .A1(n10108), .A2(n10106), .A3(n10103), .ZN(n12170) );
  INV_X1 U12725 ( .A(n11230), .ZN(n10107) );
  OAI211_X1 U12726 ( .C1(n12171), .C2(n10107), .A(n10110), .B(n10109), .ZN(
        n10108) );
  NAND2_X1 U12727 ( .A1(n11230), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10109) );
  INV_X1 U12728 ( .A(n11307), .ZN(n10110) );
  NAND2_X1 U12729 ( .A1(n13729), .A2(n13730), .ZN(n10112) );
  NAND2_X1 U12730 ( .A1(n11684), .A2(n11683), .ZN(P1_U3004) );
  NAND2_X1 U12731 ( .A1(n15663), .A2(n10114), .ZN(n10113) );
  OAI21_X1 U12732 ( .B1(n15663), .B2(n10118), .A(n10116), .ZN(n15645) );
  INV_X1 U12733 ( .A(n11457), .ZN(n10117) );
  NAND2_X1 U12734 ( .A1(n15629), .A2(n10119), .ZN(n16646) );
  NAND3_X1 U12735 ( .A1(n12132), .A2(n11196), .A3(n9724), .ZN(n10120) );
  NAND2_X1 U12736 ( .A1(n11201), .A2(n10120), .ZN(n11202) );
  AND2_X2 U12737 ( .A1(n11177), .A2(n11192), .ZN(n13275) );
  NAND2_X1 U12738 ( .A1(n12128), .A2(n10123), .ZN(n10125) );
  NAND3_X1 U12739 ( .A1(n10131), .A2(n11597), .A3(n13724), .ZN(n13823) );
  NAND2_X1 U12740 ( .A1(n11597), .A2(n11596), .ZN(n13558) );
  NAND2_X1 U12741 ( .A1(n14675), .A2(n14674), .ZN(n14673) );
  NAND2_X2 U12742 ( .A1(n10146), .A2(n10145), .ZN(n20750) );
  INV_X1 U12743 ( .A(n10656), .ZN(n10658) );
  NAND2_X1 U12744 ( .A1(n16157), .A2(n9807), .ZN(n10149) );
  AOI21_X1 U12745 ( .B1(n16157), .B2(n16158), .A(n16096), .ZN(n16146) );
  INV_X1 U12746 ( .A(n10433), .ZN(n10161) );
  NOR2_X1 U12747 ( .A1(n10162), .A2(n10433), .ZN(n10608) );
  NAND2_X1 U12748 ( .A1(n15888), .A2(n13420), .ZN(n10162) );
  NAND2_X1 U12749 ( .A1(n10165), .A2(n10163), .ZN(n11250) );
  NAND2_X1 U12750 ( .A1(n14664), .A2(n10179), .ZN(n15499) );
  AND2_X1 U12751 ( .A1(n11364), .A2(n9814), .ZN(n11400) );
  AND2_X2 U12753 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13746) );
  NAND3_X2 U12754 ( .A1(n10186), .A2(n10188), .A3(n10185), .ZN(n16119) );
  NAND3_X1 U12755 ( .A1(n9774), .A2(n10906), .A3(n14384), .ZN(n10186) );
  INV_X1 U12756 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n10192) );
  OAI21_X1 U12757 ( .B1(n14848), .B2(n16974), .A(n10193), .ZN(P2_U2986) );
  NAND2_X1 U12758 ( .A1(n14805), .A2(n16034), .ZN(n14846) );
  NAND2_X1 U12759 ( .A1(n14119), .A2(n14118), .ZN(n14121) );
  AND2_X1 U12760 ( .A1(n19979), .A2(n20121), .ZN(n16935) );
  NAND2_X1 U12761 ( .A1(n11608), .A2(n11607), .ZN(n13841) );
  AND2_X1 U12762 ( .A1(n14704), .A2(n11177), .ZN(n11494) );
  NOR2_X1 U12763 ( .A1(n11177), .A2(n11486), .ZN(n11180) );
  INV_X1 U12764 ( .A(n14760), .ZN(n14767) );
  NAND2_X1 U12765 ( .A1(n14760), .A2(n20927), .ZN(n11684) );
  INV_X1 U12766 ( .A(n13565), .ZN(n12184) );
  INV_X1 U12767 ( .A(n11400), .ZN(n11378) );
  NAND2_X1 U12768 ( .A1(n9725), .A2(n10327), .ZN(n10373) );
  AND2_X1 U12769 ( .A1(n10335), .A2(n13368), .ZN(n10329) );
  AOI22_X1 U12770 ( .A1(n9739), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(n9757), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10252) );
  OAI21_X1 U12771 ( .B1(n10402), .B2(n10398), .A(n10399), .ZN(n10377) );
  NAND2_X1 U12772 ( .A1(n9835), .A2(n9775), .ZN(n10327) );
  INV_X1 U12773 ( .A(n9722), .ZN(n13061) );
  CLKBUF_X1 U12774 ( .A(n11488), .Z(n13227) );
  OR2_X1 U12775 ( .A1(n10430), .A2(n15888), .ZN(n10431) );
  INV_X1 U12777 ( .A(n12254), .ZN(n14277) );
  INV_X1 U12778 ( .A(n10899), .ZN(n10901) );
  NAND2_X1 U12779 ( .A1(n10899), .A2(n10898), .ZN(n10903) );
  OAI22_X1 U12780 ( .A1(n13063), .A2(n12132), .B1(n12130), .B2(n12131), .ZN(
        n12133) );
  AOI21_X1 U12781 ( .B1(n10915), .B2(n10914), .A(n10913), .ZN(n16106) );
  CLKBUF_X1 U12782 ( .A(n14989), .Z(n15130) );
  AOI21_X2 U12783 ( .B1(n16170), .B2(n16169), .A(n16093), .ZN(n16157) );
  AND2_X1 U12784 ( .A1(n20845), .A2(n13943), .ZN(n16629) );
  NOR3_X1 U12785 ( .A1(n12027), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n12043), .ZN(n10196) );
  INV_X1 U12786 ( .A(n12846), .ZN(n12866) );
  AND2_X1 U12787 ( .A1(n12035), .A2(n10198), .ZN(n10197) );
  NOR2_X1 U12788 ( .A1(n12034), .A2(n12033), .ZN(n10198) );
  AND2_X1 U12789 ( .A1(n16102), .A2(n16100), .ZN(n10199) );
  AND2_X1 U12790 ( .A1(n12052), .A2(n12051), .ZN(n10200) );
  NAND2_X1 U12791 ( .A1(n18445), .A2(n18684), .ZN(n18430) );
  AND4_X1 U12792 ( .A1(n11067), .A2(n11066), .A3(n11065), .A4(n11064), .ZN(
        n10202) );
  OR2_X1 U12793 ( .A1(n12867), .A2(n19170), .ZN(n10203) );
  OR2_X1 U12794 ( .A1(n13649), .A2(n11129), .ZN(n10205) );
  AND2_X1 U12795 ( .A1(n11129), .A2(n13393), .ZN(n10206) );
  OR2_X1 U12796 ( .A1(n11553), .A2(n11192), .ZN(n10207) );
  AND2_X1 U12797 ( .A1(n10258), .A2(n10257), .ZN(n10208) );
  INV_X1 U12798 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n12027) );
  INV_X1 U12799 ( .A(n12333), .ZN(n12626) );
  NOR2_X1 U12800 ( .A1(n20476), .A2(n10474), .ZN(n10209) );
  OR2_X1 U12801 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n10210) );
  OR2_X1 U12802 ( .A1(n13058), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10211) );
  AND2_X1 U12803 ( .A1(n18524), .A2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n10212) );
  INV_X1 U12804 ( .A(n19815), .ZN(n19929) );
  AND2_X1 U12805 ( .A1(n10254), .A2(n10253), .ZN(n10214) );
  INV_X1 U12806 ( .A(n9713), .ZN(n11791) );
  INV_X1 U12807 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n10829) );
  AND2_X1 U12808 ( .A1(n15888), .A2(n13355), .ZN(n10215) );
  AND2_X1 U12809 ( .A1(n16674), .A2(n15716), .ZN(n10216) );
  AND3_X1 U12810 ( .A1(n10252), .A2(n10291), .A3(n10251), .ZN(n10217) );
  AND3_X1 U12811 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(P3_EAX_REG_8__SCAN_IN), 
        .A3(P3_EAX_REG_12__SCAN_IN), .ZN(n10218) );
  INV_X1 U12812 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n12659) );
  INV_X1 U12813 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n10828) );
  NOR2_X1 U12814 ( .A1(n12004), .A2(n16148), .ZN(n10219) );
  AND2_X1 U12815 ( .A1(n15055), .A2(n15050), .ZN(n10220) );
  OR2_X1 U12816 ( .A1(n16522), .A2(n16521), .ZN(n10221) );
  NOR2_X1 U12817 ( .A1(n17290), .A2(n12789), .ZN(n10222) );
  AND2_X1 U12818 ( .A1(n15518), .A2(n15517), .ZN(n10223) );
  AND2_X1 U12819 ( .A1(n16989), .A2(n16988), .ZN(n10224) );
  INV_X1 U12820 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n14745) );
  INV_X1 U12821 ( .A(n11677), .ZN(n11176) );
  AND2_X1 U12822 ( .A1(n11254), .A2(n11253), .ZN(n10228) );
  INV_X1 U12823 ( .A(n11257), .ZN(n11265) );
  AND2_X1 U12824 ( .A1(n21270), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11200) );
  NOR2_X1 U12825 ( .A1(n11429), .A2(n13951), .ZN(n11187) );
  AND2_X1 U12826 ( .A1(n11565), .A2(n11200), .ZN(n11201) );
  AND2_X1 U12827 ( .A1(n10349), .A2(n10353), .ZN(n11735) );
  NAND2_X1 U12828 ( .A1(n20082), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n10485) );
  OAI21_X1 U12829 ( .B1(n10931), .B2(n19736), .A(n10356), .ZN(n10357) );
  AND2_X1 U12830 ( .A1(n21110), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11501) );
  NAND2_X1 U12831 ( .A1(n12612), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n11116) );
  INV_X1 U12832 ( .A(n10455), .ZN(n14992) );
  AND4_X1 U12833 ( .A1(n10635), .A2(n10634), .A3(n10633), .A4(n10632), .ZN(
        n10639) );
  OAI22_X1 U12834 ( .A1(n14158), .A2(n10620), .B1(n20404), .B2(n10480), .ZN(
        n10481) );
  NAND2_X1 U12835 ( .A1(n13374), .A2(n10335), .ZN(n10333) );
  NOR2_X1 U12836 ( .A1(n10358), .A2(n10357), .ZN(n10359) );
  INV_X1 U12837 ( .A(n15500), .ZN(n12445) );
  OR2_X1 U12838 ( .A1(n14277), .A2(n12255), .ZN(n12256) );
  OR2_X1 U12839 ( .A1(n11374), .A2(n11373), .ZN(n11401) );
  AOI22_X1 U12840 ( .A1(n12588), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n9741), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11045) );
  AND4_X1 U12841 ( .A1(n10686), .A2(n10685), .A3(n10684), .A4(n10683), .ZN(
        n10690) );
  OAI211_X1 U12842 ( .C1(n10931), .C2(n10371), .A(n10370), .B(n10369), .ZN(
        n10372) );
  NOR2_X1 U12843 ( .A1(n19666), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12664) );
  NOR2_X1 U12844 ( .A1(n16521), .A2(n19068), .ZN(n12768) );
  NAND2_X1 U12845 ( .A1(n12209), .A2(n12144), .ZN(n12217) );
  INV_X1 U12846 ( .A(n13564), .ZN(n12183) );
  AND2_X1 U12847 ( .A1(n11418), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16728) );
  NAND2_X1 U12848 ( .A1(n13420), .A2(n13419), .ZN(n13426) );
  NAND2_X1 U12849 ( .A1(n15052), .A2(n10220), .ZN(n15053) );
  INV_X1 U12850 ( .A(n15989), .ZN(n11963) );
  NAND2_X1 U12851 ( .A1(n12048), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n12049) );
  NAND2_X1 U12852 ( .A1(n10342), .A2(n10341), .ZN(n11998) );
  AOI211_X1 U12853 ( .C1(n9740), .C2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A(
        n12872), .B(n12871), .ZN(n12873) );
  NOR2_X1 U12854 ( .A1(n12925), .A2(n12924), .ZN(n12926) );
  NAND2_X1 U12855 ( .A1(n12987), .A2(n18616), .ZN(n18606) );
  INV_X1 U12856 ( .A(n12801), .ZN(n12811) );
  AOI211_X1 U12857 ( .C1(n17979), .C2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A(
        n12713), .B(n12712), .ZN(n12714) );
  NAND2_X1 U12858 ( .A1(n11177), .A2(n11554), .ZN(n11195) );
  NOR2_X1 U12859 ( .A1(n12368), .A2(n16573), .ZN(n12318) );
  INV_X1 U12860 ( .A(n12228), .ZN(n12229) );
  NAND2_X1 U12861 ( .A1(n11273), .A2(n11272), .ZN(n11274) );
  AND2_X1 U12862 ( .A1(n11615), .A2(n11614), .ZN(n14082) );
  AND4_X1 U12863 ( .A1(n11171), .A2(n11170), .A3(n11169), .A4(n11168), .ZN(
        n11172) );
  AND2_X1 U12864 ( .A1(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n12553), .ZN(
        n12554) );
  INV_X1 U12865 ( .A(n12631), .ZN(n12333) );
  NAND2_X1 U12866 ( .A1(n12217), .A2(n12216), .ZN(n13837) );
  NAND2_X1 U12867 ( .A1(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n12164) );
  INV_X1 U12868 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20941) );
  INV_X1 U12869 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n21010) );
  INV_X1 U12870 ( .A(n15078), .ZN(n15075) );
  INV_X1 U12871 ( .A(n15976), .ZN(n11966) );
  NOR2_X1 U12872 ( .A1(n19961), .A2(n19962), .ZN(n13636) );
  AND2_X1 U12873 ( .A1(n10787), .A2(n10199), .ZN(n10788) );
  OR2_X1 U12874 ( .A1(n19769), .A2(n11790), .ZN(n16134) );
  AND2_X1 U12875 ( .A1(n10744), .A2(n10746), .ZN(n19782) );
  INV_X1 U12876 ( .A(n10348), .ZN(n10353) );
  NOR2_X1 U12877 ( .A1(n19656), .A2(n19666), .ZN(n12661) );
  OAI21_X1 U12878 ( .B1(n17615), .B2(n18430), .A(n19354), .ZN(n18523) );
  NAND2_X1 U12879 ( .A1(n19517), .A2(n19509), .ZN(n18873) );
  XNOR2_X1 U12880 ( .A(n12967), .B(n12912), .ZN(n12910) );
  NOR2_X1 U12881 ( .A1(n18662), .A2(n12850), .ZN(n12862) );
  NOR2_X1 U12882 ( .A1(n12995), .A2(n12944), .ZN(n12954) );
  NAND2_X1 U12883 ( .A1(n12229), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12234) );
  NAND2_X1 U12884 ( .A1(n11321), .A2(n11320), .ZN(n13860) );
  NOR2_X1 U12885 ( .A1(n13937), .A2(n13936), .ZN(n13953) );
  NAND2_X1 U12886 ( .A1(n13527), .A2(n13222), .ZN(n13651) );
  INV_X1 U12887 ( .A(n13047), .ZN(n13048) );
  NAND2_X1 U12888 ( .A1(n12282), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n12286) );
  NAND2_X1 U12889 ( .A1(n9722), .A2(n12140), .ZN(n12141) );
  AND2_X1 U12890 ( .A1(n16671), .A2(n11459), .ZN(n15659) );
  INV_X1 U12891 ( .A(n14533), .ZN(n14571) );
  NAND2_X1 U12892 ( .A1(n15813), .A2(n13856), .ZN(n20982) );
  NAND2_X1 U12893 ( .A1(n13857), .A2(n13896), .ZN(n14431) );
  INV_X1 U12894 ( .A(n13856), .ZN(n13892) );
  NAND2_X1 U12895 ( .A1(n14589), .A2(n13896), .ZN(n14639) );
  AND2_X1 U12896 ( .A1(n11334), .A2(n11333), .ZN(n14088) );
  INV_X1 U12897 ( .A(n14318), .ZN(n21119) );
  AND2_X1 U12898 ( .A1(n10867), .A2(n11706), .ZN(n13734) );
  OR2_X1 U12899 ( .A1(n19927), .A2(n20333), .ZN(n19815) );
  NAND2_X1 U12900 ( .A1(n19923), .A2(n13419), .ZN(n13349) );
  INV_X1 U12901 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n16200) );
  INV_X1 U12902 ( .A(n12050), .ZN(n12051) );
  NOR2_X1 U12903 ( .A1(n10818), .A2(n16243), .ZN(n16063) );
  AND3_X1 U12904 ( .A1(n12001), .A2(n12000), .A3(n11999), .ZN(n13772) );
  NAND2_X1 U12905 ( .A1(n20131), .A2(n13961), .ZN(n20309) );
  NAND2_X1 U12906 ( .A1(n19715), .A2(n9752), .ZN(n12784) );
  NOR2_X1 U12907 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12672) );
  INV_X1 U12908 ( .A(n18523), .ZN(n18483) );
  OR2_X1 U12909 ( .A1(n12931), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n12934) );
  NOR2_X1 U12910 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n18509), .ZN(
        n18463) );
  INV_X1 U12911 ( .A(n19515), .ZN(n18914) );
  XNOR2_X1 U12912 ( .A(n18967), .B(n12881), .ZN(n18644) );
  INV_X1 U12913 ( .A(n19501), .ZN(n14691) );
  INV_X1 U12914 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19522) );
  NAND2_X1 U12915 ( .A1(n12954), .A2(n12963), .ZN(n17149) );
  AND3_X1 U12916 ( .A1(n16548), .A2(P1_REIP_REG_22__SCAN_IN), .A3(
        P1_REIP_REG_23__SCAN_IN), .ZN(n16539) );
  NOR2_X1 U12917 ( .A1(n21227), .A2(n15436), .ZN(n16594) );
  NAND2_X1 U12918 ( .A1(n12235), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n12257) );
  AND2_X1 U12919 ( .A1(n20845), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20849) );
  OAI22_X1 U12920 ( .A1(n15160), .A2(n15543), .B1(n13054), .B2(n16644), .ZN(
        n13055) );
  INV_X1 U12921 ( .A(n11179), .ZN(n14703) );
  INV_X1 U12922 ( .A(n15603), .ZN(n15606) );
  NAND2_X1 U12923 ( .A1(n12495), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n12552) );
  NAND2_X1 U12924 ( .A1(n12372), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n12368) );
  NOR2_X1 U12925 ( .A1(n14667), .A2(n14666), .ZN(n16711) );
  NAND2_X1 U12926 ( .A1(n12211), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12228) );
  INV_X1 U12927 ( .A(n16743), .ZN(n16722) );
  OAI21_X1 U12928 ( .B1(n13060), .B2(n10211), .A(n12141), .ZN(n12142) );
  OR2_X1 U12929 ( .A1(n13068), .A2(n13067), .ZN(n13069) );
  NOR2_X1 U12930 ( .A1(n15736), .A2(n13450), .ZN(n15783) );
  INV_X1 U12931 ( .A(n20925), .ZN(n16809) );
  NOR2_X1 U12932 ( .A1(n20982), .A2(n14312), .ZN(n14533) );
  OAI21_X1 U12933 ( .B1(n21017), .B2(n21048), .A(n21016), .ZN(n21051) );
  INV_X1 U12934 ( .A(n14431), .ZN(n14228) );
  NOR2_X1 U12935 ( .A1(n15813), .A2(n13892), .ZN(n14589) );
  AND2_X1 U12936 ( .A1(n14589), .A2(n14588), .ZN(n21105) );
  AND2_X1 U12937 ( .A1(n14589), .A2(n14313), .ZN(n14218) );
  NOR2_X1 U12938 ( .A1(n21119), .A2(n14587), .ZN(n21169) );
  AND2_X1 U12939 ( .A1(n14318), .A2(n14313), .ZN(n20972) );
  NOR2_X1 U12940 ( .A1(n21119), .A2(n14312), .ZN(n14530) );
  OR2_X1 U12941 ( .A1(n12109), .A2(n12108), .ZN(n12110) );
  NAND2_X1 U12942 ( .A1(n15853), .A2(n16066), .ZN(n15852) );
  AND2_X1 U12943 ( .A1(n12102), .A2(n12094), .ZN(n19922) );
  INV_X1 U12944 ( .A(n19960), .ZN(n19953) );
  INV_X1 U12945 ( .A(n13696), .ZN(n14851) );
  AND2_X1 U12946 ( .A1(n14308), .A2(n14307), .ZN(n16933) );
  INV_X1 U12947 ( .A(n16020), .ZN(n19974) );
  INV_X1 U12948 ( .A(n20043), .ZN(n17010) );
  AOI21_X1 U12949 ( .B1(n14801), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n9802), .ZN(n14804) );
  AND2_X1 U12950 ( .A1(n12028), .A2(n13754), .ZN(n13319) );
  AND2_X1 U12951 ( .A1(n11729), .A2(n13139), .ZN(n12028) );
  XNOR2_X1 U12952 ( .A(n13511), .B(n13513), .ZN(n20701) );
  OAI21_X1 U12953 ( .B1(n20079), .B2(n20122), .A(n20512), .ZN(n20125) );
  INV_X1 U12954 ( .A(n20695), .ZN(n20187) );
  NOR2_X1 U12955 ( .A1(n20309), .A2(n20187), .ZN(n20245) );
  OR2_X1 U12956 ( .A1(n20701), .A2(n13961), .ZN(n20218) );
  NOR2_X1 U12957 ( .A1(n20309), .A2(n20473), .ZN(n20286) );
  INV_X1 U12958 ( .A(n20218), .ZN(n20075) );
  AND2_X1 U12959 ( .A1(n20706), .A2(n20074), .ZN(n20365) );
  AND2_X1 U12960 ( .A1(n20706), .A2(n20718), .ZN(n20695) );
  AND2_X1 U12961 ( .A1(n20505), .A2(n20482), .ZN(n20501) );
  INV_X1 U12962 ( .A(n20569), .ZN(n20524) );
  INV_X1 U12963 ( .A(n20605), .ZN(n20579) );
  INV_X1 U12964 ( .A(n20396), .ZN(n20600) );
  NAND2_X1 U12965 ( .A1(n12994), .A2(n19503), .ZN(n19501) );
  INV_X1 U12966 ( .A(n17583), .ZN(n17618) );
  INV_X1 U12967 ( .A(n17602), .ZN(n17609) );
  INV_X1 U12968 ( .A(n17621), .ZN(n17459) );
  NOR2_X1 U12969 ( .A1(n17801), .A2(n17802), .ZN(n17770) );
  OAI211_X1 U12970 ( .C1(n17913), .C2(n17781), .A(n12746), .B(n12745), .ZN(
        n18053) );
  NOR2_X1 U12971 ( .A1(n9754), .A2(n18092), .ZN(n18088) );
  NOR2_X1 U12972 ( .A1(n18097), .A2(n18125), .ZN(n18115) );
  NAND2_X1 U12973 ( .A1(n12880), .A2(n12879), .ZN(n12980) );
  AND2_X1 U12974 ( .A1(n18049), .A2(n9754), .ZN(n18114) );
  INV_X1 U12975 ( .A(n18540), .ZN(n18596) );
  NOR2_X1 U12976 ( .A1(n19040), .A2(n17269), .ZN(n18678) );
  INV_X1 U12977 ( .A(n13009), .ZN(n13010) );
  NAND2_X1 U12978 ( .A1(n18492), .A2(n18512), .ZN(n18513) );
  INV_X1 U12979 ( .A(n18877), .ZN(n18926) );
  INV_X1 U12980 ( .A(n20849), .ZN(n20818) );
  INV_X1 U12981 ( .A(n16629), .ZN(n20847) );
  INV_X1 U12982 ( .A(n16609), .ZN(n20860) );
  INV_X1 U12983 ( .A(n15612), .ZN(n15549) );
  OR2_X1 U12984 ( .A1(n15584), .A2(n15583), .ZN(n16677) );
  OR2_X1 U12985 ( .A1(n13529), .A2(n13528), .ZN(n20903) );
  INV_X1 U12986 ( .A(n20921), .ZN(n13693) );
  INV_X1 U12987 ( .A(n12643), .ZN(n12644) );
  NAND2_X1 U12988 ( .A1(n20773), .A2(n12637), .ZN(n16670) );
  NAND2_X1 U12989 ( .A1(n16670), .A2(n13477), .ZN(n16743) );
  INV_X1 U12990 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n21110) );
  AND2_X1 U12991 ( .A1(n13293), .A2(n13292), .ZN(n21275) );
  NAND2_X1 U12992 ( .A1(n20940), .A2(n21006), .ZN(n21005) );
  NAND2_X1 U12993 ( .A1(n20940), .A2(n14313), .ZN(n21018) );
  OR2_X1 U12994 ( .A1(n21008), .A2(n21007), .ZN(n21080) );
  NAND2_X1 U12995 ( .A1(n14589), .A2(n21006), .ZN(n21109) );
  NAND2_X1 U12996 ( .A1(n14318), .A2(n21006), .ZN(n21173) );
  INV_X1 U12997 ( .A(n21169), .ZN(n14532) );
  INV_X1 U12998 ( .A(n14530), .ZN(n14350) );
  NOR2_X1 U12999 ( .A1(n12111), .A2(n12110), .ZN(n12112) );
  OR2_X1 U13000 ( .A1(n12104), .A2(n12103), .ZN(n19919) );
  INV_X1 U13001 ( .A(n19927), .ZN(n19887) );
  XNOR2_X1 U13002 ( .A(n13482), .B(n13483), .ZN(n20706) );
  INV_X1 U13003 ( .A(n20701), .ZN(n20131) );
  INV_X1 U13004 ( .A(n16935), .ZN(n16023) );
  INV_X1 U13005 ( .A(n19974), .ZN(n19979) );
  NAND2_X1 U13006 ( .A1(n13118), .A2(n20756), .ZN(n20027) );
  NAND2_X1 U13007 ( .A1(n14791), .A2(n20046), .ZN(n14797) );
  INV_X1 U13008 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n17014) );
  INV_X1 U13009 ( .A(n17008), .ZN(n20045) );
  INV_X1 U13010 ( .A(n20051), .ZN(n16202) );
  INV_X1 U13011 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20732) );
  NAND2_X1 U13012 ( .A1(n20365), .A2(n20075), .ZN(n20156) );
  OR2_X1 U13013 ( .A1(n20218), .A2(n20187), .ZN(n20203) );
  OR2_X1 U13014 ( .A1(n20218), .A2(n20473), .ZN(n20276) );
  INV_X1 U13015 ( .A(n20286), .ZN(n20296) );
  NAND2_X1 U13016 ( .A1(n20555), .A2(n20075), .ZN(n20325) );
  INV_X1 U13017 ( .A(n20354), .ZN(n20362) );
  OR2_X1 U13018 ( .A1(n20474), .A2(n20363), .ZN(n20386) );
  NAND2_X1 U13019 ( .A1(n20505), .A2(n20365), .ZN(n20395) );
  NAND2_X1 U13020 ( .A1(n20505), .A2(n20695), .ZN(n20442) );
  AOI21_X1 U13021 ( .B1(n13812), .B2(n13813), .A(n13811), .ZN(n20472) );
  OR2_X1 U13022 ( .A1(n20474), .A2(n20473), .ZN(n20537) );
  INV_X1 U13023 ( .A(n20455), .ZN(n20575) );
  OR2_X1 U13024 ( .A1(n20474), .A2(n20308), .ZN(n20605) );
  NAND2_X1 U13025 ( .A1(n19694), .A2(n19537), .ZN(n17269) );
  AOI21_X1 U13026 ( .B1(n12794), .B2(n17608), .A(n12793), .ZN(n12795) );
  NAND2_X1 U13027 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n17459), .ZN(n17586) );
  NAND2_X1 U13028 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n17814), .ZN(n17802) );
  AND2_X1 U13029 ( .A1(n18048), .A2(n9754), .ZN(n18045) );
  AOI211_X1 U13030 ( .C1(n17954), .C2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A(
        n12908), .B(n12907), .ZN(n18175) );
  INV_X1 U13031 ( .A(n18196), .ZN(n18186) );
  OR2_X1 U13032 ( .A1(n19548), .A2(n18262), .ZN(n18264) );
  NAND2_X1 U13033 ( .A1(n18271), .A2(n18205), .ZN(n18269) );
  INV_X1 U13034 ( .A(n18317), .ZN(n18312) );
  NAND2_X1 U13035 ( .A1(n18948), .A2(P3_REIP_REG_29__SCAN_IN), .ZN(n17134) );
  INV_X1 U13036 ( .A(n18547), .ZN(n18529) );
  INV_X1 U13037 ( .A(n18426), .ZN(n18491) );
  NAND2_X1 U13038 ( .A1(n18678), .A2(n17103), .ZN(n18540) );
  INV_X1 U13039 ( .A(n18646), .ZN(n18681) );
  AND2_X1 U13040 ( .A1(n13011), .A2(n13010), .ZN(n13012) );
  NOR2_X1 U13041 ( .A1(n18513), .A2(n18819), .ZN(n18846) );
  INV_X1 U13042 ( .A(n18832), .ZN(n19017) );
  AND2_X1 U13043 ( .A1(n13081), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n14706)
         );
  NAND2_X1 U13044 ( .A1(n13057), .A2(n13056), .ZN(P1_U2842) );
  NAND2_X1 U13045 ( .A1(n12113), .A2(n12112), .ZN(P2_U2824) );
  INV_X1 U13046 ( .A(n12795), .ZN(P3_U2641) );
  NAND2_X1 U13047 ( .A1(n13013), .A2(n13012), .ZN(P3_U2833) );
  INV_X1 U13048 ( .A(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10409) );
  AND3_X4 U13049 ( .A1(n10230), .A2(n10229), .A3(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10316) );
  INV_X1 U13050 ( .A(n10316), .ZN(n15083) );
  AOI22_X1 U13051 ( .A1(n10316), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n10315), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10234) );
  AOI22_X1 U13053 ( .A1(n10444), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n10446), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10233) );
  AND2_X4 U13054 ( .A1(n10461), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10455) );
  AOI22_X1 U13055 ( .A1(n10455), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n9747), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10232) );
  AND2_X4 U13056 ( .A1(n10460), .A2(n13749), .ZN(n14927) );
  AND2_X4 U13057 ( .A1(n13748), .A2(n13749), .ZN(n14989) );
  AOI22_X1 U13058 ( .A1(n14927), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n14989), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10231) );
  AOI22_X1 U13059 ( .A1(n9739), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n9758), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10238) );
  AOI22_X1 U13060 ( .A1(n10316), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n9753), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10237) );
  AOI22_X1 U13061 ( .A1(n14927), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n14989), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n10236) );
  AOI22_X1 U13062 ( .A1(n10455), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n10317), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10235) );
  AOI22_X1 U13063 ( .A1(n9739), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(n9758), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n10242) );
  AOI22_X1 U13064 ( .A1(n10316), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n9753), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n10241) );
  AOI22_X1 U13065 ( .A1(n14927), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n14989), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10240) );
  AOI22_X1 U13066 ( .A1(n10455), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n9747), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10239) );
  NAND4_X1 U13067 ( .A1(n10242), .A2(n10241), .A3(n10240), .A4(n10239), .ZN(
        n10243) );
  NAND2_X1 U13068 ( .A1(n10243), .A2(n10291), .ZN(n10250) );
  AOI22_X1 U13069 ( .A1(n9739), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n9757), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10247) );
  AOI22_X1 U13070 ( .A1(n10455), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n10317), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n10246) );
  AOI22_X1 U13071 ( .A1(n14927), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n14989), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n10245) );
  AOI22_X1 U13072 ( .A1(n10316), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n10315), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10244) );
  NAND4_X1 U13073 ( .A1(n10247), .A2(n10246), .A3(n10245), .A4(n10244), .ZN(
        n10248) );
  NAND2_X4 U13074 ( .A1(n10250), .A2(n10249), .ZN(n13368) );
  INV_X2 U13075 ( .A(n14929), .ZN(n10446) );
  AOI22_X1 U13076 ( .A1(n10316), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n10315), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10251) );
  AOI22_X1 U13077 ( .A1(n14927), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n14989), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10254) );
  AOI22_X1 U13078 ( .A1(n10455), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n10317), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10253) );
  NAND2_X1 U13079 ( .A1(n10217), .A2(n10214), .ZN(n10261) );
  AOI22_X1 U13080 ( .A1(n10444), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n9757), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10256) );
  AOI22_X1 U13081 ( .A1(n10316), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n9753), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10255) );
  AOI22_X1 U13082 ( .A1(n14927), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n14989), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10258) );
  AOI22_X1 U13083 ( .A1(n10455), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n10317), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10257) );
  AOI22_X1 U13084 ( .A1(n10316), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n9753), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10262) );
  AOI22_X1 U13085 ( .A1(n10455), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n10317), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10265) );
  AOI22_X1 U13086 ( .A1(n14927), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n14989), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10264) );
  AOI22_X1 U13087 ( .A1(n9739), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(n9757), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10263) );
  NAND4_X1 U13088 ( .A1(n10266), .A2(n10265), .A3(n10264), .A4(n10263), .ZN(
        n10273) );
  AOI22_X1 U13089 ( .A1(n9739), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n9758), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10270) );
  AOI22_X1 U13090 ( .A1(n10316), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n9753), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10269) );
  AOI22_X1 U13091 ( .A1(n14927), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n14989), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10268) );
  AOI22_X1 U13092 ( .A1(n10455), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n9747), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10267) );
  AOI22_X1 U13093 ( .A1(n10455), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n10317), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10276) );
  AOI22_X1 U13094 ( .A1(n14927), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n14989), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10278) );
  AOI22_X1 U13095 ( .A1(n9739), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n10446), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10277) );
  NAND3_X1 U13096 ( .A1(n9791), .A2(n10278), .A3(n10277), .ZN(n10285) );
  AOI22_X1 U13097 ( .A1(n10455), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n9747), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10280) );
  AOI22_X1 U13098 ( .A1(n10315), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_9__6__SCAN_IN), .B2(n10316), .ZN(n10279) );
  AOI22_X1 U13099 ( .A1(n14927), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n14989), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10282) );
  AOI22_X1 U13100 ( .A1(n9739), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n9758), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10281) );
  NAND3_X1 U13101 ( .A1(n10283), .A2(n10282), .A3(n10281), .ZN(n10284) );
  NAND2_X2 U13102 ( .A1(n10285), .A2(n10284), .ZN(n13350) );
  AOI22_X1 U13103 ( .A1(n10444), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n10446), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10289) );
  AOI22_X1 U13104 ( .A1(n14927), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n14989), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10288) );
  AOI22_X1 U13105 ( .A1(n10455), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n9747), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10287) );
  AOI22_X1 U13106 ( .A1(n10316), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10315), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10286) );
  AOI22_X1 U13107 ( .A1(n10444), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10446), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10292) );
  AOI22_X1 U13108 ( .A1(n10316), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n9753), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10290) );
  AOI22_X1 U13109 ( .A1(n14927), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n14989), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10294) );
  AOI22_X1 U13110 ( .A1(n10455), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10317), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10293) );
  NAND2_X1 U13111 ( .A1(n13350), .A2(n10326), .ZN(n10331) );
  NOR2_X2 U13112 ( .A1(n10346), .A2(n10331), .ZN(n10348) );
  AOI22_X1 U13113 ( .A1(n9739), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10446), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10299) );
  AOI22_X1 U13114 ( .A1(n10316), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n10315), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10298) );
  AOI22_X1 U13115 ( .A1(n14927), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n14989), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10297) );
  AOI22_X1 U13116 ( .A1(n10455), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n10317), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10296) );
  NAND4_X1 U13117 ( .A1(n10299), .A2(n10298), .A3(n10297), .A4(n10296), .ZN(
        n10305) );
  AOI22_X1 U13118 ( .A1(n10444), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n9757), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10303) );
  AOI22_X1 U13119 ( .A1(n10316), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10315), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10302) );
  AOI22_X1 U13120 ( .A1(n14927), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n14989), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10301) );
  AOI22_X1 U13121 ( .A1(n10455), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n9747), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10300) );
  NAND4_X1 U13122 ( .A1(n10303), .A2(n10302), .A3(n10301), .A4(n10300), .ZN(
        n10304) );
  NAND2_X1 U13123 ( .A1(n10348), .A2(n20750), .ZN(n12098) );
  INV_X1 U13124 ( .A(n10325), .ZN(n11718) );
  AND2_X1 U13125 ( .A1(n11718), .A2(n13368), .ZN(n10307) );
  AOI21_X1 U13126 ( .B1(n9758), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A(n10309), .ZN(n10313) );
  AOI22_X1 U13127 ( .A1(n10444), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n10315), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10312) );
  AOI22_X1 U13128 ( .A1(n14927), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n14989), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10311) );
  AOI22_X1 U13129 ( .A1(n10455), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n10317), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10310) );
  NAND4_X1 U13130 ( .A1(n10313), .A2(n10312), .A3(n10311), .A4(n10310), .ZN(
        n10314) );
  NAND2_X1 U13131 ( .A1(n10314), .A2(n10291), .ZN(n10324) );
  AOI22_X1 U13132 ( .A1(n9739), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n9758), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10321) );
  AOI22_X1 U13133 ( .A1(n14927), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n14989), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10320) );
  AOI22_X1 U13134 ( .A1(n10316), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n10315), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10319) );
  AOI22_X1 U13135 ( .A1(n10455), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n9747), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10318) );
  NAND4_X1 U13136 ( .A1(n10321), .A2(n10320), .A3(n10319), .A4(n10318), .ZN(
        n10322) );
  NAND2_X1 U13137 ( .A1(n10322), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10323) );
  INV_X1 U13138 ( .A(n11715), .ZN(n11996) );
  NOR2_X1 U13139 ( .A1(n10331), .A2(n20755), .ZN(n10328) );
  NAND2_X2 U13140 ( .A1(n11692), .A2(n11730), .ZN(n13111) );
  AND3_X2 U13141 ( .A1(n10330), .A2(n10329), .A3(n13111), .ZN(n11736) );
  INV_X1 U13142 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n14877) );
  INV_X2 U13143 ( .A(n13368), .ZN(n20121) );
  NAND2_X1 U13144 ( .A1(n10331), .A2(n10337), .ZN(n11713) );
  NAND2_X1 U13145 ( .A1(n11713), .A2(n11994), .ZN(n10332) );
  INV_X1 U13146 ( .A(n10343), .ZN(n10334) );
  NAND3_X1 U13147 ( .A1(n10361), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n10334), 
        .ZN(n10350) );
  NAND2_X1 U13148 ( .A1(n13369), .A2(n11990), .ZN(n10340) );
  MUX2_X1 U13149 ( .A(n10336), .B(n13368), .S(n10335), .Z(n10339) );
  AND2_X1 U13150 ( .A1(n10325), .A2(n10337), .ZN(n10338) );
  NAND3_X1 U13151 ( .A1(n10340), .A2(n10339), .A3(n10338), .ZN(n10342) );
  INV_X1 U13152 ( .A(n13141), .ZN(n10341) );
  NAND2_X1 U13153 ( .A1(n10343), .A2(n11998), .ZN(n10345) );
  INV_X1 U13154 ( .A(n10346), .ZN(n10347) );
  NAND3_X1 U13155 ( .A1(n10861), .A2(n10325), .A3(n20755), .ZN(n10349) );
  INV_X1 U13156 ( .A(n20754), .ZN(n13119) );
  INV_X1 U13157 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n10352) );
  INV_X1 U13158 ( .A(n10353), .ZN(n13796) );
  INV_X1 U13159 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n19736) );
  NAND2_X1 U13160 ( .A1(n20749), .A2(n13792), .ZN(n13794) );
  NAND2_X1 U13161 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n10355) );
  AND2_X1 U13162 ( .A1(n13794), .A2(n10355), .ZN(n10356) );
  INV_X1 U13163 ( .A(n10361), .ZN(n10364) );
  INV_X1 U13164 ( .A(n13743), .ZN(n10366) );
  OAI21_X1 U13165 ( .B1(n13794), .B2(n20732), .A(n10925), .ZN(n10365) );
  AOI21_X1 U13166 ( .B1(n10366), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n10365), 
        .ZN(n10367) );
  NAND2_X1 U13167 ( .A1(n10368), .A2(n10367), .ZN(n10403) );
  NAND2_X1 U13168 ( .A1(n10404), .A2(n10403), .ZN(n10402) );
  INV_X1 U13169 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n10371) );
  NAND2_X1 U13170 ( .A1(n11019), .A2(P2_EBX_REG_1__SCAN_IN), .ZN(n10370) );
  NAND2_X1 U13171 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n10369) );
  NAND2_X1 U13172 ( .A1(n10382), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10375) );
  INV_X1 U13174 ( .A(n13794), .ZN(n10389) );
  AOI22_X1 U13175 ( .A1(n11732), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(n10389), 
        .B2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n10374) );
  NAND2_X1 U13176 ( .A1(n10402), .A2(n10398), .ZN(n10376) );
  NAND2_X1 U13177 ( .A1(n10377), .A2(n10376), .ZN(n10396) );
  INV_X1 U13178 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n10380) );
  NAND2_X1 U13179 ( .A1(n11019), .A2(P2_EBX_REG_2__SCAN_IN), .ZN(n10379) );
  NAND2_X1 U13180 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n10378) );
  NAND2_X1 U13181 ( .A1(n10382), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10384) );
  AOI21_X1 U13182 ( .B1(n20749), .B2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n10383) );
  INV_X1 U13183 ( .A(n10385), .ZN(n10387) );
  NAND2_X1 U13184 ( .A1(n10387), .A2(n10386), .ZN(n10388) );
  NAND2_X1 U13185 ( .A1(n10382), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10391) );
  NAND2_X1 U13186 ( .A1(n10389), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n10390) );
  INV_X1 U13187 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n14775) );
  NAND2_X1 U13188 ( .A1(n11026), .A2(P2_EBX_REG_3__SCAN_IN), .ZN(n10394) );
  NAND2_X1 U13189 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n10393) );
  OAI211_X1 U13190 ( .C1(n10931), .C2(n14775), .A(n10394), .B(n10393), .ZN(
        n10395) );
  BUF_X4 U13191 ( .A(n10435), .Z(n13412) );
  XNOR2_X2 U13192 ( .A(n10396), .B(n10397), .ZN(n10430) );
  INV_X1 U13193 ( .A(n10398), .ZN(n10401) );
  INV_X1 U13194 ( .A(n10399), .ZN(n10400) );
  XNOR2_X2 U13195 ( .A(n10401), .B(n10400), .ZN(n10411) );
  INV_X1 U13196 ( .A(n10411), .ZN(n10408) );
  INV_X1 U13197 ( .A(n10403), .ZN(n10406) );
  INV_X1 U13198 ( .A(n10404), .ZN(n10405) );
  NAND2_X1 U13199 ( .A1(n10406), .A2(n10405), .ZN(n10407) );
  NAND2_X1 U13200 ( .A1(n10408), .A2(n19923), .ZN(n10436) );
  NAND2_X1 U13201 ( .A1(n19923), .A2(n10411), .ZN(n10425) );
  INV_X1 U13202 ( .A(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n14472) );
  OAI22_X1 U13203 ( .A1(n10409), .A2(n20549), .B1(n20367), .B2(n14472), .ZN(
        n10414) );
  INV_X1 U13204 ( .A(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n14469) );
  INV_X1 U13205 ( .A(n10402), .ZN(n10410) );
  XNOR2_X2 U13206 ( .A(n10411), .B(n10410), .ZN(n15888) );
  OR2_X1 U13207 ( .A1(n15888), .A2(n19923), .ZN(n10421) );
  INV_X1 U13208 ( .A(n19923), .ZN(n13355) );
  INV_X1 U13209 ( .A(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11858) );
  OAI22_X1 U13210 ( .A1(n14469), .A2(n10616), .B1(n20514), .B2(n11858), .ZN(
        n10413) );
  NOR2_X1 U13211 ( .A1(n10414), .A2(n10413), .ZN(n10443) );
  INV_X1 U13212 ( .A(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10417) );
  INV_X1 U13213 ( .A(n10425), .ZN(n10415) );
  INV_X1 U13214 ( .A(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10416) );
  OAI22_X1 U13215 ( .A1(n10417), .A2(n10620), .B1(n20476), .B2(n10416), .ZN(
        n10424) );
  INV_X1 U13216 ( .A(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n14468) );
  INV_X1 U13217 ( .A(n10418), .ZN(n10419) );
  INV_X1 U13218 ( .A(n10421), .ZN(n10422) );
  INV_X1 U13219 ( .A(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n15037) );
  OAI22_X1 U13220 ( .A1(n14468), .A2(n20404), .B1(n13810), .B2(n15037), .ZN(
        n10423) );
  NOR2_X1 U13221 ( .A1(n10424), .A2(n10423), .ZN(n10442) );
  AOI22_X1 U13222 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n9763), .B1(
        n20162), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10441) );
  INV_X1 U13223 ( .A(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10429) );
  OR3_X2 U13224 ( .A1(n13412), .A2(n15873), .A3(n10425), .ZN(n10611) );
  INV_X1 U13225 ( .A(n13412), .ZN(n10427) );
  INV_X1 U13226 ( .A(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10428) );
  OAI22_X1 U13227 ( .A1(n10429), .A2(n10611), .B1(n20129), .B2(n10428), .ZN(
        n10439) );
  INV_X1 U13228 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10434) );
  OR2_X2 U13229 ( .A1(n10433), .A2(n10431), .ZN(n20077) );
  NAND2_X1 U13230 ( .A1(n13420), .A2(n13259), .ZN(n10432) );
  OR2_X2 U13231 ( .A1(n10433), .A2(n10432), .ZN(n20220) );
  INV_X1 U13232 ( .A(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n15029) );
  OAI22_X1 U13233 ( .A1(n10434), .A2(n20077), .B1(n20220), .B2(n15029), .ZN(
        n10438) );
  INV_X1 U13234 ( .A(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n15031) );
  INV_X1 U13235 ( .A(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10452) );
  OAI22_X1 U13236 ( .A1(n15031), .A2(n10659), .B1(n20300), .B2(n10452), .ZN(
        n10437) );
  NOR3_X1 U13237 ( .A1(n10439), .A2(n10438), .A3(n10437), .ZN(n10440) );
  INV_X1 U13238 ( .A(n10444), .ZN(n14928) );
  NAND2_X2 U13239 ( .A1(n10445), .A2(n10291), .ZN(n14919) );
  INV_X1 U13240 ( .A(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11857) );
  NAND2_X2 U13241 ( .A1(n13745), .A2(n10291), .ZN(n14917) );
  OAI22_X1 U13242 ( .A1(n14919), .A2(n11857), .B1(n14917), .B2(n14469), .ZN(
        n10454) );
  AND2_X2 U13243 ( .A1(n10447), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n14967) );
  NOR2_X4 U13244 ( .A1(n10870), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11881) );
  AOI22_X1 U13245 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n14967), .B1(
        n11881), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10451) );
  AND2_X2 U13246 ( .A1(n10448), .A2(n10449), .ZN(n14450) );
  NAND2_X1 U13247 ( .A1(n14450), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n10450) );
  OAI211_X1 U13248 ( .C1(n10452), .C2(n14473), .A(n10451), .B(n10450), .ZN(
        n10453) );
  NOR2_X1 U13249 ( .A1(n10454), .A2(n10453), .ZN(n10468) );
  AND2_X2 U13250 ( .A1(n10462), .A2(n10291), .ZN(n14908) );
  AOI22_X1 U13251 ( .A1(n14908), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n14910), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10467) );
  INV_X2 U13252 ( .A(n15083), .ZN(n15129) );
  NAND2_X1 U13253 ( .A1(n10631), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n10459) );
  NAND2_X1 U13254 ( .A1(n14951), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n10458) );
  AND2_X1 U13255 ( .A1(n10448), .A2(n14932), .ZN(n10500) );
  AOI22_X1 U13256 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n10500), .B1(
        n14885), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10457) );
  NAND2_X1 U13257 ( .A1(n10507), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(
        n10456) );
  AND4_X1 U13258 ( .A1(n10459), .A2(n10458), .A3(n10457), .A4(n10456), .ZN(
        n10466) );
  AOI22_X1 U13259 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n10498), .B1(
        n10499), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10464) );
  AND2_X2 U13260 ( .A1(n10462), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14909) );
  NAND2_X1 U13261 ( .A1(n14909), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n10463) );
  AND2_X1 U13262 ( .A1(n10464), .A2(n10463), .ZN(n10465) );
  NAND4_X1 U13263 ( .A1(n10468), .A2(n10467), .A3(n10466), .A4(n10465), .ZN(
        n10569) );
  INV_X1 U13264 ( .A(n10569), .ZN(n11776) );
  NAND2_X1 U13265 ( .A1(n11776), .A2(n9759), .ZN(n10470) );
  INV_X1 U13266 ( .A(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10472) );
  INV_X1 U13267 ( .A(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n14164) );
  AOI21_X1 U13268 ( .B1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n20162), .A(
        n10473), .ZN(n10492) );
  INV_X1 U13269 ( .A(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10474) );
  NAND2_X1 U13270 ( .A1(n9763), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n10478) );
  INV_X1 U13271 ( .A(n20300), .ZN(n10475) );
  NAND2_X1 U13272 ( .A1(n10475), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n10477) );
  INV_X1 U13273 ( .A(n10611), .ZN(n20252) );
  NAND2_X1 U13274 ( .A1(n20252), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n10476) );
  NAND4_X1 U13275 ( .A1(n10478), .A2(n20755), .A3(n10477), .A4(n10476), .ZN(
        n10479) );
  NOR2_X1 U13276 ( .A1(n10209), .A2(n10479), .ZN(n10491) );
  INV_X1 U13277 ( .A(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n14157) );
  INV_X1 U13278 ( .A(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n14991) );
  INV_X1 U13279 ( .A(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n14158) );
  INV_X1 U13280 ( .A(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10480) );
  NOR2_X1 U13281 ( .A1(n10482), .A2(n10481), .ZN(n10490) );
  INV_X1 U13282 ( .A(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n14981) );
  INV_X1 U13283 ( .A(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10483) );
  OAI22_X1 U13284 ( .A1(n14981), .A2(n20220), .B1(n20514), .B2(n10483), .ZN(
        n10488) );
  INV_X1 U13285 ( .A(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10486) );
  INV_X1 U13286 ( .A(n10659), .ZN(n20189) );
  NAND2_X1 U13287 ( .A1(n20189), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n10484) );
  OAI211_X1 U13288 ( .C1(n10486), .C2(n20129), .A(n10485), .B(n10484), .ZN(
        n10487) );
  NOR2_X1 U13289 ( .A1(n10488), .A2(n10487), .ZN(n10489) );
  AOI22_X1 U13290 ( .A1(n10631), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n14910), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10497) );
  AOI22_X1 U13291 ( .A1(n14956), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n10507), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10496) );
  AOI22_X1 U13292 ( .A1(n14908), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n14909), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10495) );
  INV_X1 U13293 ( .A(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n13971) );
  INV_X1 U13294 ( .A(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11802) );
  OAI22_X1 U13295 ( .A1(n14919), .A2(n13971), .B1(n14473), .B2(n11802), .ZN(
        n10493) );
  INV_X1 U13296 ( .A(n10493), .ZN(n10494) );
  NAND4_X1 U13297 ( .A1(n10497), .A2(n10496), .A3(n10495), .A4(n10494), .ZN(
        n10506) );
  AOI22_X1 U13298 ( .A1(n10498), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n10499), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10504) );
  AOI22_X1 U13299 ( .A1(n10500), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n11881), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10503) );
  AOI22_X1 U13300 ( .A1(n14450), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n14885), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10502) );
  AOI22_X1 U13301 ( .A1(n14951), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n14967), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10501) );
  NAND4_X1 U13302 ( .A1(n10504), .A2(n10503), .A3(n10502), .A4(n10501), .ZN(
        n10505) );
  AOI22_X1 U13303 ( .A1(n10631), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_9__1__SCAN_IN), .B2(n14910), .ZN(n10512) );
  AOI22_X1 U13304 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n14908), .B1(
        n14956), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10511) );
  AOI22_X1 U13305 ( .A1(n14957), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n14951), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10510) );
  INV_X1 U13306 ( .A(n14473), .ZN(n10508) );
  AOI22_X1 U13307 ( .A1(n10508), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n10507), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10509) );
  NAND4_X1 U13308 ( .A1(n10512), .A2(n10511), .A3(n10510), .A4(n10509), .ZN(
        n10518) );
  AOI22_X1 U13309 ( .A1(n10498), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n10499), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10516) );
  AOI22_X1 U13310 ( .A1(n10500), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n14885), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10515) );
  AOI22_X1 U13311 ( .A1(n14450), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_15__1__SCAN_IN), .B2(n11881), .ZN(n10514) );
  AOI22_X1 U13312 ( .A1(n14909), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__1__SCAN_IN), .B2(n14967), .ZN(n10513) );
  NAND4_X1 U13313 ( .A1(n10516), .A2(n10515), .A3(n10514), .A4(n10513), .ZN(
        n10517) );
  NOR2_X1 U13314 ( .A1(n11748), .A2(n11756), .ZN(n10519) );
  NAND2_X1 U13315 ( .A1(n9759), .A2(n10519), .ZN(n10882) );
  NAND2_X1 U13316 ( .A1(n10631), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n10523) );
  NAND2_X1 U13317 ( .A1(n14951), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n10522) );
  INV_X1 U13318 ( .A(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n15344) );
  AOI22_X1 U13319 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n10500), .B1(
        n14885), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10521) );
  NAND2_X1 U13320 ( .A1(n10507), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(
        n10520) );
  NAND4_X1 U13321 ( .A1(n10523), .A2(n10522), .A3(n10521), .A4(n10520), .ZN(
        n10529) );
  AOI22_X1 U13322 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n10498), .B1(
        n10499), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10527) );
  NAND2_X1 U13323 ( .A1(n14908), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(
        n10526) );
  NAND2_X1 U13324 ( .A1(n14909), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(
        n10525) );
  NAND2_X1 U13325 ( .A1(n14910), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n10524) );
  NAND4_X1 U13326 ( .A1(n10527), .A2(n10526), .A3(n10525), .A4(n10524), .ZN(
        n10528) );
  NOR2_X1 U13327 ( .A1(n10529), .A2(n10528), .ZN(n10536) );
  INV_X1 U13328 ( .A(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11838) );
  INV_X1 U13329 ( .A(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n14143) );
  OAI22_X1 U13330 ( .A1(n14919), .A2(n11838), .B1(n14917), .B2(n14143), .ZN(
        n10534) );
  INV_X1 U13331 ( .A(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10532) );
  AOI22_X1 U13332 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n14967), .B1(
        n11881), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10531) );
  NAND2_X1 U13333 ( .A1(n14450), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n10530) );
  OAI211_X1 U13334 ( .C1(n14473), .C2(n10532), .A(n10531), .B(n10530), .ZN(
        n10533) );
  NOR2_X1 U13335 ( .A1(n10534), .A2(n10533), .ZN(n10535) );
  NAND2_X1 U13336 ( .A1(n10882), .A2(n11762), .ZN(n10537) );
  NAND2_X1 U13337 ( .A1(n10631), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n10543) );
  NAND2_X1 U13338 ( .A1(n14951), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n10542) );
  AOI22_X1 U13339 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n10500), .B1(
        n14885), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10541) );
  NAND2_X1 U13340 ( .A1(n10507), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n10540) );
  NAND4_X1 U13341 ( .A1(n10543), .A2(n10542), .A3(n10541), .A4(n10540), .ZN(
        n10549) );
  AOI22_X1 U13342 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n10498), .B1(
        n10499), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10547) );
  NAND2_X1 U13343 ( .A1(n14908), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n10546) );
  NAND2_X1 U13344 ( .A1(n14909), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n10545) );
  NAND2_X1 U13345 ( .A1(n14910), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n10544) );
  NAND4_X1 U13346 ( .A1(n10547), .A2(n10546), .A3(n10545), .A4(n10544), .ZN(
        n10548) );
  NOR2_X1 U13347 ( .A1(n10549), .A2(n10548), .ZN(n10556) );
  INV_X1 U13348 ( .A(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n10550) );
  INV_X1 U13349 ( .A(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11946) );
  OAI22_X1 U13350 ( .A1(n14919), .A2(n10550), .B1(n14917), .B2(n11946), .ZN(
        n10554) );
  INV_X1 U13351 ( .A(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n14963) );
  AOI22_X1 U13352 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n14967), .B1(
        n11881), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10552) );
  NAND2_X1 U13353 ( .A1(n14450), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n10551) );
  OAI211_X1 U13354 ( .C1(n14963), .C2(n14473), .A(n10552), .B(n10551), .ZN(
        n10553) );
  NOR2_X1 U13355 ( .A1(n10554), .A2(n10553), .ZN(n10555) );
  INV_X1 U13356 ( .A(P2_EBX_REG_1__SCAN_IN), .ZN(n10557) );
  NAND2_X1 U13357 ( .A1(n10557), .A2(n10352), .ZN(n10558) );
  MUX2_X1 U13358 ( .A(n11756), .B(n10558), .S(n10561), .Z(n10578) );
  MUX2_X1 U13359 ( .A(n20721), .B(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .S(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Z(n10849) );
  NAND2_X1 U13360 ( .A1(n10849), .A2(n10865), .ZN(n10560) );
  NAND2_X1 U13361 ( .A1(n20721), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10559) );
  NAND2_X1 U13362 ( .A1(n10560), .A2(n10559), .ZN(n10564) );
  XNOR2_X1 U13363 ( .A(n20710), .B(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10562) );
  XNOR2_X1 U13364 ( .A(n10564), .B(n10562), .ZN(n11690) );
  INV_X1 U13365 ( .A(n11690), .ZN(n11699) );
  MUX2_X1 U13366 ( .A(n11762), .B(n11699), .S(n11730), .Z(n10850) );
  INV_X1 U13367 ( .A(n10562), .ZN(n10563) );
  NAND2_X1 U13368 ( .A1(n10564), .A2(n10563), .ZN(n10566) );
  NAND2_X1 U13369 ( .A1(n20710), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10565) );
  NAND2_X1 U13370 ( .A1(n10566), .A2(n10565), .ZN(n10602) );
  INV_X1 U13371 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n10567) );
  MUX2_X1 U13372 ( .A(n10567), .B(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n10601) );
  INV_X1 U13373 ( .A(n10601), .ZN(n10568) );
  XNOR2_X1 U13374 ( .A(n10602), .B(n10568), .ZN(n10863) );
  MUX2_X1 U13375 ( .A(n10569), .B(n10863), .S(n11730), .Z(n10854) );
  INV_X1 U13376 ( .A(P2_EBX_REG_3__SCAN_IN), .ZN(n10570) );
  MUX2_X1 U13377 ( .A(n10854), .B(n10570), .S(n10838), .Z(n10571) );
  OAI21_X1 U13378 ( .B1(n10572), .B2(n10571), .A(n10646), .ZN(n14785) );
  INV_X1 U13379 ( .A(n10865), .ZN(n10575) );
  NAND2_X1 U13380 ( .A1(n10573), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n10574) );
  NAND2_X1 U13381 ( .A1(n10575), .A2(n10574), .ZN(n11693) );
  MUX2_X1 U13382 ( .A(n11748), .B(n11693), .S(n11730), .Z(n10851) );
  MUX2_X1 U13383 ( .A(n10851), .B(n10352), .S(n10838), .Z(n19920) );
  OR2_X1 U13384 ( .A1(n19920), .A2(n14877), .ZN(n13250) );
  NAND3_X1 U13385 ( .A1(n10838), .A2(P2_EBX_REG_1__SCAN_IN), .A3(
        P2_EBX_REG_0__SCAN_IN), .ZN(n10576) );
  NAND2_X1 U13386 ( .A1(n10578), .A2(n10576), .ZN(n15880) );
  NOR2_X1 U13387 ( .A1(n13250), .A2(n15880), .ZN(n10577) );
  NAND2_X1 U13388 ( .A1(n13250), .A2(n15880), .ZN(n13122) );
  OAI21_X1 U13389 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n10577), .A(
        n13122), .ZN(n13332) );
  XNOR2_X1 U13390 ( .A(n10579), .B(n10578), .ZN(n15872) );
  INV_X1 U13391 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n13340) );
  XNOR2_X1 U13392 ( .A(n15872), .B(n13340), .ZN(n13331) );
  OR2_X1 U13393 ( .A1(n13332), .A2(n13331), .ZN(n20048) );
  INV_X1 U13394 ( .A(n15872), .ZN(n10580) );
  NAND2_X1 U13395 ( .A1(n10580), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10581) );
  NAND2_X1 U13396 ( .A1(n20048), .A2(n10581), .ZN(n14772) );
  NAND2_X1 U13397 ( .A1(n14774), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10582) );
  NAND2_X1 U13398 ( .A1(n10631), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n10586) );
  NAND2_X1 U13399 ( .A1(n14951), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n10585) );
  AOI22_X1 U13400 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n10500), .B1(
        n14885), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10584) );
  NAND2_X1 U13401 ( .A1(n10507), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n10583) );
  NAND4_X1 U13402 ( .A1(n10586), .A2(n10585), .A3(n10584), .A4(n10583), .ZN(
        n10592) );
  INV_X1 U13403 ( .A(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n15317) );
  AOI22_X1 U13404 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n10498), .B1(
        n10499), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10590) );
  NAND2_X1 U13405 ( .A1(n14908), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n10589) );
  NAND2_X1 U13406 ( .A1(n14909), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n10588) );
  NAND2_X1 U13407 ( .A1(n14910), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n10587) );
  NAND4_X1 U13408 ( .A1(n10590), .A2(n10589), .A3(n10588), .A4(n10587), .ZN(
        n10591) );
  NOR2_X1 U13409 ( .A1(n10592), .A2(n10591), .ZN(n10599) );
  INV_X1 U13410 ( .A(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10593) );
  INV_X1 U13411 ( .A(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n14449) );
  OAI22_X1 U13412 ( .A1(n14919), .A2(n10593), .B1(n14917), .B2(n14449), .ZN(
        n10597) );
  INV_X1 U13413 ( .A(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11880) );
  AOI22_X1 U13414 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n14967), .B1(
        n11881), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10595) );
  NAND2_X1 U13415 ( .A1(n14450), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n10594) );
  OAI211_X1 U13416 ( .C1(n14473), .C2(n11880), .A(n10595), .B(n10594), .ZN(
        n10596) );
  NOR2_X1 U13417 ( .A1(n10597), .A2(n10596), .ZN(n10598) );
  NOR2_X1 U13418 ( .A1(n10291), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n10600) );
  AOI21_X1 U13419 ( .B1(n10602), .B2(n10601), .A(n10600), .ZN(n10857) );
  INV_X1 U13420 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n16520) );
  NOR2_X1 U13421 ( .A1(n16520), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n10603) );
  NAND2_X1 U13422 ( .A1(n10857), .A2(n10603), .ZN(n10864) );
  INV_X1 U13423 ( .A(n10864), .ZN(n10604) );
  MUX2_X1 U13424 ( .A(n11777), .B(n10604), .S(n11730), .Z(n10852) );
  MUX2_X1 U13425 ( .A(n10852), .B(P2_EBX_REG_4__SCAN_IN), .S(n10838), .Z(
        n10645) );
  XNOR2_X1 U13426 ( .A(n10646), .B(n10645), .ZN(n10605) );
  XNOR2_X1 U13427 ( .A(n10605), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n20030) );
  INV_X1 U13428 ( .A(n10605), .ZN(n14868) );
  NAND2_X1 U13429 ( .A1(n14868), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10606) );
  NAND2_X1 U13430 ( .A1(n10607), .A2(n10606), .ZN(n14258) );
  AOI22_X1 U13431 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n9763), .B1(
        n20162), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10626) );
  INV_X1 U13432 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10609) );
  INV_X1 U13433 ( .A(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n15080) );
  OAI22_X1 U13434 ( .A1(n10609), .A2(n20077), .B1(n20220), .B2(n15080), .ZN(
        n10615) );
  INV_X1 U13435 ( .A(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10610) );
  INV_X1 U13436 ( .A(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n14893) );
  OAI22_X1 U13437 ( .A1(n10610), .A2(n20129), .B1(n20300), .B2(n14893), .ZN(
        n10613) );
  INV_X1 U13438 ( .A(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n15081) );
  INV_X1 U13439 ( .A(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n15082) );
  OAI22_X1 U13440 ( .A1(n15081), .A2(n10659), .B1(n10611), .B2(n15082), .ZN(
        n10612) );
  OR2_X1 U13441 ( .A1(n10613), .A2(n10612), .ZN(n10614) );
  NOR2_X1 U13442 ( .A1(n10615), .A2(n10614), .ZN(n10625) );
  INV_X1 U13443 ( .A(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n14892) );
  INV_X1 U13444 ( .A(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n15090) );
  OAI22_X1 U13445 ( .A1(n14892), .A2(n20549), .B1(n13810), .B2(n15090), .ZN(
        n10619) );
  INV_X1 U13446 ( .A(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11897) );
  INV_X1 U13447 ( .A(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10617) );
  OAI22_X1 U13448 ( .A1(n11897), .A2(n10616), .B1(n20476), .B2(n10617), .ZN(
        n10618) );
  NOR2_X1 U13449 ( .A1(n10619), .A2(n10618), .ZN(n10624) );
  INV_X1 U13450 ( .A(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11903) );
  INV_X1 U13451 ( .A(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n15092) );
  OAI22_X1 U13452 ( .A1(n11903), .A2(n20514), .B1(n20367), .B2(n15092), .ZN(
        n10622) );
  INV_X1 U13453 ( .A(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n15091) );
  INV_X1 U13454 ( .A(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11902) );
  OAI22_X1 U13455 ( .A1(n15091), .A2(n10620), .B1(n20404), .B2(n11902), .ZN(
        n10621) );
  NOR2_X1 U13456 ( .A1(n10622), .A2(n10621), .ZN(n10623) );
  NAND4_X1 U13457 ( .A1(n10626), .A2(n10625), .A3(n10624), .A4(n10623), .ZN(
        n10644) );
  INV_X1 U13458 ( .A(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11901) );
  OAI22_X1 U13459 ( .A1(n14919), .A2(n11901), .B1(n14917), .B2(n11897), .ZN(
        n10630) );
  AOI22_X1 U13460 ( .A1(n14967), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n11881), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10628) );
  NAND2_X1 U13461 ( .A1(n14450), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n10627) );
  OAI211_X1 U13462 ( .C1(n14893), .C2(n14473), .A(n10628), .B(n10627), .ZN(
        n10629) );
  NOR2_X1 U13463 ( .A1(n10630), .A2(n10629), .ZN(n10641) );
  AOI22_X1 U13464 ( .A1(n14908), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n14910), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10640) );
  NAND2_X1 U13465 ( .A1(n10631), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n10635) );
  NAND2_X1 U13466 ( .A1(n14951), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n10634) );
  AOI22_X1 U13467 ( .A1(n10500), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n14885), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10633) );
  NAND2_X1 U13468 ( .A1(n10507), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n10632) );
  AOI22_X1 U13469 ( .A1(n10498), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n10499), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10637) );
  NAND2_X1 U13470 ( .A1(n14909), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n10636) );
  AND2_X1 U13471 ( .A1(n10637), .A2(n10636), .ZN(n10638) );
  NAND4_X1 U13472 ( .A1(n10641), .A2(n10640), .A3(n10639), .A4(n10638), .ZN(
        n10647) );
  INV_X1 U13473 ( .A(n10647), .ZN(n10642) );
  NAND2_X1 U13474 ( .A1(n10642), .A2(n9759), .ZN(n10643) );
  NAND2_X1 U13475 ( .A1(n10892), .A2(n11790), .ZN(n10652) );
  NAND2_X1 U13476 ( .A1(n10306), .A2(n10647), .ZN(n11781) );
  INV_X1 U13477 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n14852) );
  NAND2_X1 U13478 ( .A1(n10838), .A2(n14852), .ZN(n10648) );
  NAND2_X1 U13479 ( .A1(n11781), .A2(n10648), .ZN(n10649) );
  NOR2_X1 U13480 ( .A1(n10650), .A2(n10649), .ZN(n10651) );
  OR2_X1 U13481 ( .A1(n10700), .A2(n10651), .ZN(n19903) );
  INV_X1 U13482 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n10926) );
  NAND2_X1 U13483 ( .A1(n14258), .A2(n14259), .ZN(n10655) );
  NAND2_X1 U13484 ( .A1(n10653), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10654) );
  NAND2_X1 U13485 ( .A1(n10655), .A2(n10654), .ZN(n14382) );
  NAND2_X1 U13486 ( .A1(n10658), .A2(n10657), .ZN(n10696) );
  AOI22_X1 U13487 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n9763), .B1(
        n20162), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10677) );
  INV_X1 U13488 ( .A(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n13506) );
  INV_X1 U13489 ( .A(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n15105) );
  OAI22_X1 U13490 ( .A1(n13506), .A2(n20077), .B1(n20220), .B2(n15105), .ZN(
        n10664) );
  INV_X1 U13491 ( .A(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11924) );
  INV_X1 U13492 ( .A(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n15107) );
  OAI22_X1 U13493 ( .A1(n11924), .A2(n20300), .B1(n20129), .B2(n15107), .ZN(
        n10662) );
  INV_X1 U13494 ( .A(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10660) );
  INV_X1 U13495 ( .A(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n15106) );
  OAI22_X1 U13496 ( .A1(n10660), .A2(n10611), .B1(n10659), .B2(n15106), .ZN(
        n10661) );
  OR2_X1 U13497 ( .A1(n10662), .A2(n10661), .ZN(n10663) );
  NOR2_X1 U13498 ( .A1(n10664), .A2(n10663), .ZN(n10676) );
  INV_X1 U13499 ( .A(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n14918) );
  INV_X1 U13500 ( .A(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10665) );
  OAI22_X1 U13501 ( .A1(n14918), .A2(n10616), .B1(n20549), .B2(n10665), .ZN(
        n10668) );
  INV_X1 U13502 ( .A(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10666) );
  INV_X1 U13503 ( .A(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n15104) );
  OAI22_X1 U13504 ( .A1(n10666), .A2(n10620), .B1(n20404), .B2(n15104), .ZN(
        n10667) );
  NOR2_X1 U13505 ( .A1(n10668), .A2(n10667), .ZN(n10675) );
  INV_X1 U13506 ( .A(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n14922) );
  INV_X1 U13507 ( .A(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10669) );
  OAI22_X1 U13508 ( .A1(n14922), .A2(n20367), .B1(n13810), .B2(n10669), .ZN(
        n10673) );
  INV_X1 U13509 ( .A(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10671) );
  INV_X1 U13510 ( .A(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10670) );
  OAI22_X1 U13511 ( .A1(n10671), .A2(n20514), .B1(n20476), .B2(n10670), .ZN(
        n10672) );
  NOR2_X1 U13512 ( .A1(n10673), .A2(n10672), .ZN(n10674) );
  NAND4_X1 U13513 ( .A1(n10677), .A2(n10676), .A3(n10675), .A4(n10674), .ZN(
        n10694) );
  INV_X1 U13514 ( .A(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10678) );
  OAI22_X1 U13515 ( .A1(n14919), .A2(n10678), .B1(n14917), .B2(n14918), .ZN(
        n10682) );
  AOI22_X1 U13516 ( .A1(n14967), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n11881), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10680) );
  NAND2_X1 U13517 ( .A1(n14450), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n10679) );
  OAI211_X1 U13518 ( .C1(n11924), .C2(n14473), .A(n10680), .B(n10679), .ZN(
        n10681) );
  NOR2_X1 U13519 ( .A1(n10682), .A2(n10681), .ZN(n10692) );
  AOI22_X1 U13520 ( .A1(n14908), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n14910), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10691) );
  NAND2_X1 U13521 ( .A1(n10631), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n10686) );
  NAND2_X1 U13522 ( .A1(n14951), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n10685) );
  AOI22_X1 U13523 ( .A1(n10500), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n14885), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10684) );
  NAND2_X1 U13524 ( .A1(n10507), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n10683) );
  AOI22_X1 U13525 ( .A1(n10498), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n10499), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10688) );
  NAND2_X1 U13526 ( .A1(n14909), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n10687) );
  AND2_X1 U13527 ( .A1(n10688), .A2(n10687), .ZN(n10689) );
  NAND4_X1 U13528 ( .A1(n10692), .A2(n10691), .A3(n10690), .A4(n10689), .ZN(
        n10698) );
  INV_X1 U13529 ( .A(n10698), .ZN(n11786) );
  NAND2_X1 U13530 ( .A1(n11786), .A2(n9759), .ZN(n10693) );
  INV_X1 U13531 ( .A(n10877), .ZN(n10695) );
  NAND2_X1 U13532 ( .A1(n10696), .A2(n10877), .ZN(n10697) );
  INV_X1 U13533 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n10932) );
  MUX2_X1 U13534 ( .A(n10698), .B(n10932), .S(n10838), .Z(n10699) );
  OR2_X1 U13535 ( .A1(n10700), .A2(n10699), .ZN(n10701) );
  NAND2_X1 U13536 ( .A1(n10707), .A2(n10701), .ZN(n19889) );
  INV_X1 U13537 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n14394) );
  NAND2_X1 U13538 ( .A1(n10702), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10703) );
  MUX2_X1 U13539 ( .A(n11790), .B(P2_EBX_REG_7__SCAN_IN), .S(n10838), .Z(
        n10705) );
  INV_X1 U13540 ( .A(n10712), .ZN(n10718) );
  NAND2_X1 U13541 ( .A1(n10838), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n10704) );
  XNOR2_X1 U13542 ( .A(n10718), .B(n10704), .ZN(n14208) );
  INV_X1 U13543 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n11984) );
  NOR2_X1 U13544 ( .A1(n11790), .A2(n11984), .ZN(n10907) );
  NAND2_X1 U13545 ( .A1(n14208), .A2(n10907), .ZN(n16181) );
  INV_X1 U13546 ( .A(n10705), .ZN(n10706) );
  XNOR2_X1 U13547 ( .A(n10707), .B(n10706), .ZN(n19878) );
  NAND2_X1 U13548 ( .A1(n19878), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16195) );
  NAND2_X1 U13549 ( .A1(n16181), .A2(n16195), .ZN(n10708) );
  NAND2_X1 U13550 ( .A1(n14208), .A2(n10826), .ZN(n10709) );
  NAND2_X1 U13551 ( .A1(n10709), .A2(n11984), .ZN(n16182) );
  INV_X1 U13552 ( .A(n19878), .ZN(n10710) );
  INV_X1 U13553 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n10936) );
  NAND2_X1 U13554 ( .A1(n10710), .A2(n10936), .ZN(n16194) );
  AND2_X1 U13555 ( .A1(n16182), .A2(n16194), .ZN(n10711) );
  NAND2_X1 U13556 ( .A1(n10838), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n10713) );
  MUX2_X1 U13557 ( .A(n10838), .B(n10713), .S(n10714), .Z(n10716) );
  INV_X1 U13558 ( .A(n10720), .ZN(n10715) );
  NAND2_X1 U13559 ( .A1(n10716), .A2(n10715), .ZN(n10724) );
  INV_X1 U13560 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n16407) );
  OAI21_X1 U13561 ( .B1(n10724), .B2(n11790), .A(n16407), .ZN(n16403) );
  INV_X1 U13562 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n10717) );
  NAND2_X1 U13563 ( .A1(n10838), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n10719) );
  OAI21_X1 U13564 ( .B1(n10720), .B2(n10719), .A(n10824), .ZN(n10721) );
  AOI21_X1 U13565 ( .B1(n9771), .B2(n10826), .A(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16991) );
  INV_X1 U13566 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n10722) );
  NOR2_X1 U13567 ( .A1(n11790), .A2(n10722), .ZN(n10723) );
  NAND2_X1 U13568 ( .A1(n9771), .A2(n10723), .ZN(n16989) );
  INV_X1 U13569 ( .A(n10724), .ZN(n14288) );
  NOR2_X1 U13570 ( .A1(n11790), .A2(n16407), .ZN(n10725) );
  NAND2_X1 U13571 ( .A1(n14288), .A2(n10725), .ZN(n16988) );
  INV_X1 U13572 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n19958) );
  NAND2_X1 U13573 ( .A1(n10838), .A2(P2_EBX_REG_11__SCAN_IN), .ZN(n10726) );
  NOR2_X1 U13574 ( .A1(n10727), .A2(n10726), .ZN(n10728) );
  NOR2_X1 U13575 ( .A1(n10730), .A2(n10728), .ZN(n19863) );
  NAND2_X1 U13576 ( .A1(n19863), .A2(n10826), .ZN(n10729) );
  NOR2_X1 U13577 ( .A1(n10729), .A2(n16393), .ZN(n16381) );
  NAND2_X1 U13578 ( .A1(n10729), .A2(n16393), .ZN(n16379) );
  OAI21_X1 U13579 ( .B1(n16378), .B2(n16381), .A(n16379), .ZN(n16367) );
  NAND2_X1 U13580 ( .A1(n10838), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n10731) );
  INV_X1 U13581 ( .A(n10736), .ZN(n10764) );
  INV_X1 U13582 ( .A(n10731), .ZN(n10732) );
  NAND2_X1 U13583 ( .A1(n10733), .A2(n10732), .ZN(n10734) );
  NAND2_X1 U13584 ( .A1(n10764), .A2(n10734), .ZN(n19853) );
  INV_X1 U13585 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n16373) );
  OR2_X1 U13586 ( .A1(n11790), .A2(n16373), .ZN(n10735) );
  NAND2_X1 U13587 ( .A1(n16367), .A2(n16368), .ZN(n16088) );
  NAND2_X1 U13588 ( .A1(n10838), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n10742) );
  NAND2_X1 U13589 ( .A1(n10838), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n10763) );
  INV_X1 U13590 ( .A(P2_EBX_REG_14__SCAN_IN), .ZN(n10757) );
  INV_X1 U13591 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n10737) );
  NAND2_X1 U13592 ( .A1(n10757), .A2(n10737), .ZN(n10738) );
  INV_X1 U13593 ( .A(P2_EBX_REG_16__SCAN_IN), .ZN(n14256) );
  INV_X1 U13594 ( .A(P2_EBX_REG_17__SCAN_IN), .ZN(n10739) );
  NAND2_X1 U13595 ( .A1(n14256), .A2(n10739), .ZN(n10740) );
  NAND2_X1 U13596 ( .A1(n10838), .A2(n10740), .ZN(n10741) );
  MUX2_X1 U13597 ( .A(n10838), .B(n10742), .S(n10770), .Z(n10744) );
  INV_X1 U13598 ( .A(n10770), .ZN(n10743) );
  INV_X1 U13599 ( .A(P2_EBX_REG_18__SCAN_IN), .ZN(n10748) );
  NAND2_X1 U13600 ( .A1(n10743), .A2(n10748), .ZN(n10746) );
  NAND2_X1 U13601 ( .A1(n19782), .A2(n10826), .ZN(n10745) );
  INV_X1 U13602 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n16320) );
  NAND2_X1 U13603 ( .A1(n10745), .A2(n16320), .ZN(n16145) );
  NAND3_X1 U13604 ( .A1(n10746), .A2(P2_EBX_REG_19__SCAN_IN), .A3(n10838), 
        .ZN(n10751) );
  INV_X1 U13605 ( .A(P2_EBX_REG_19__SCAN_IN), .ZN(n10747) );
  NAND2_X1 U13606 ( .A1(n10748), .A2(n10747), .ZN(n10749) );
  AND2_X1 U13607 ( .A1(n10838), .A2(n10749), .ZN(n10750) );
  INV_X1 U13608 ( .A(n10781), .ZN(n10785) );
  NAND2_X1 U13609 ( .A1(n10751), .A2(n10785), .ZN(n19769) );
  INV_X1 U13610 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n16307) );
  NAND2_X1 U13611 ( .A1(n16134), .A2(n16307), .ZN(n10752) );
  NAND2_X1 U13612 ( .A1(n16145), .A2(n10752), .ZN(n16097) );
  INV_X1 U13613 ( .A(n10754), .ZN(n10759) );
  AND2_X1 U13614 ( .A1(n10838), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n10753) );
  INV_X1 U13615 ( .A(n10824), .ZN(n10815) );
  AOI21_X1 U13616 ( .B1(n10759), .B2(n10753), .A(n10815), .ZN(n10755) );
  NAND2_X1 U13617 ( .A1(n10754), .A2(n14256), .ZN(n10769) );
  NAND2_X1 U13618 ( .A1(n10755), .A2(n10769), .ZN(n19806) );
  OR2_X1 U13619 ( .A1(n19806), .A2(n11790), .ZN(n10756) );
  XNOR2_X1 U13620 ( .A(n10756), .B(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n16169) );
  NAND2_X1 U13621 ( .A1(n10762), .A2(n10757), .ZN(n10775) );
  AND2_X1 U13622 ( .A1(n10838), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n10758) );
  NAND2_X1 U13623 ( .A1(n10775), .A2(n10758), .ZN(n10760) );
  NAND2_X1 U13624 ( .A1(n10760), .A2(n10759), .ZN(n19817) );
  OR2_X1 U13625 ( .A1(n19817), .A2(n11790), .ZN(n10761) );
  INV_X1 U13626 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n16340) );
  NAND2_X1 U13627 ( .A1(n10761), .A2(n16340), .ZN(n16942) );
  INV_X1 U13628 ( .A(n10762), .ZN(n10774) );
  NAND2_X1 U13629 ( .A1(n10764), .A2(n9945), .ZN(n10765) );
  NAND2_X1 U13630 ( .A1(n10774), .A2(n10765), .ZN(n19840) );
  OR2_X1 U13631 ( .A1(n19840), .A2(n11790), .ZN(n10766) );
  INV_X1 U13632 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n10796) );
  NAND2_X1 U13633 ( .A1(n10766), .A2(n10796), .ZN(n16959) );
  OR2_X1 U13634 ( .A1(n19853), .A2(n11790), .ZN(n10767) );
  NAND2_X1 U13635 ( .A1(n10767), .A2(n16373), .ZN(n16369) );
  AND3_X1 U13636 ( .A1(n16942), .A2(n16959), .A3(n16369), .ZN(n10778) );
  AND2_X1 U13637 ( .A1(n10838), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n10768) );
  NAND2_X1 U13638 ( .A1(n10769), .A2(n10768), .ZN(n10771) );
  NAND2_X1 U13639 ( .A1(n10771), .A2(n10770), .ZN(n19795) );
  OR2_X1 U13640 ( .A1(n19795), .A2(n11790), .ZN(n10772) );
  INV_X1 U13641 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n16159) );
  NAND2_X1 U13642 ( .A1(n10772), .A2(n16159), .ZN(n16095) );
  NAND2_X1 U13643 ( .A1(n10774), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n10773) );
  MUX2_X1 U13644 ( .A(n10774), .B(n10773), .S(n10838), .Z(n10776) );
  NAND2_X1 U13645 ( .A1(n10776), .A2(n10775), .ZN(n19831) );
  INV_X1 U13646 ( .A(n19831), .ZN(n10777) );
  NAND2_X1 U13647 ( .A1(n10777), .A2(n10826), .ZN(n10798) );
  INV_X1 U13648 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n16353) );
  NAND2_X1 U13649 ( .A1(n10798), .A2(n16353), .ZN(n16349) );
  NAND4_X1 U13650 ( .A1(n16169), .A2(n10778), .A3(n16095), .A4(n16349), .ZN(
        n10779) );
  NOR2_X1 U13651 ( .A1(n16097), .A2(n10779), .ZN(n10787) );
  INV_X1 U13652 ( .A(P2_EBX_REG_20__SCAN_IN), .ZN(n10780) );
  AND3_X1 U13653 ( .A1(n10782), .A2(P2_EBX_REG_21__SCAN_IN), .A3(n10838), .ZN(
        n10783) );
  OR2_X1 U13654 ( .A1(n10802), .A2(n10783), .ZN(n19747) );
  INV_X1 U13655 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n16280) );
  OAI21_X1 U13656 ( .B1(n19747), .B2(n11790), .A(n16280), .ZN(n16102) );
  NAND2_X1 U13657 ( .A1(n10838), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n10784) );
  XNOR2_X1 U13658 ( .A(n10785), .B(n10784), .ZN(n19757) );
  NAND2_X1 U13659 ( .A1(n19757), .A2(n10826), .ZN(n10786) );
  INV_X1 U13660 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n16297) );
  NAND2_X1 U13661 ( .A1(n10786), .A2(n16297), .ZN(n16100) );
  NAND2_X1 U13662 ( .A1(n16088), .A2(n10788), .ZN(n16078) );
  INV_X1 U13663 ( .A(n19747), .ZN(n10790) );
  NOR2_X1 U13664 ( .A1(n11790), .A2(n16280), .ZN(n10789) );
  NAND2_X1 U13665 ( .A1(n10790), .A2(n10789), .ZN(n16101) );
  NOR2_X1 U13666 ( .A1(n11790), .A2(n16320), .ZN(n10791) );
  NAND2_X1 U13667 ( .A1(n19782), .A2(n10791), .ZN(n16144) );
  OAI21_X1 U13668 ( .B1(n16134), .B2(n16307), .A(n16144), .ZN(n16099) );
  NOR2_X1 U13669 ( .A1(n11790), .A2(n16297), .ZN(n10792) );
  NOR2_X1 U13670 ( .A1(n16099), .A2(n16118), .ZN(n10801) );
  OR2_X1 U13671 ( .A1(n11790), .A2(n16159), .ZN(n10793) );
  OR2_X1 U13672 ( .A1(n19795), .A2(n10793), .ZN(n16094) );
  INV_X1 U13673 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n10974) );
  OR2_X1 U13674 ( .A1(n11790), .A2(n10974), .ZN(n10794) );
  OR2_X1 U13675 ( .A1(n19806), .A2(n10794), .ZN(n16092) );
  OR2_X1 U13676 ( .A1(n11790), .A2(n16340), .ZN(n10795) );
  OR2_X1 U13677 ( .A1(n11790), .A2(n10796), .ZN(n10797) );
  OR2_X1 U13678 ( .A1(n19840), .A2(n10797), .ZN(n16958) );
  AND4_X1 U13679 ( .A1(n16094), .A2(n16092), .A3(n16941), .A4(n16958), .ZN(
        n10800) );
  INV_X1 U13680 ( .A(n10798), .ZN(n10799) );
  NAND2_X1 U13681 ( .A1(n10799), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n16350) );
  AND4_X1 U13682 ( .A1(n16101), .A2(n10801), .A3(n10800), .A4(n16350), .ZN(
        n16077) );
  NAND2_X1 U13683 ( .A1(n10838), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n10803) );
  NAND2_X1 U13684 ( .A1(n10804), .A2(n9941), .ZN(n10805) );
  NAND2_X1 U13685 ( .A1(n10813), .A2(n10805), .ZN(n16459) );
  OR2_X1 U13686 ( .A1(n16459), .A2(n11790), .ZN(n10807) );
  INV_X1 U13687 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n16273) );
  OR2_X1 U13688 ( .A1(n10807), .A2(n16273), .ZN(n16076) );
  AND2_X1 U13689 ( .A1(n16077), .A2(n16076), .ZN(n10806) );
  NAND2_X1 U13690 ( .A1(n16078), .A2(n10806), .ZN(n14754) );
  NAND2_X1 U13691 ( .A1(n10807), .A2(n16273), .ZN(n16075) );
  NAND2_X1 U13692 ( .A1(n10838), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n10808) );
  XNOR2_X1 U13693 ( .A(n10813), .B(n10808), .ZN(n16900) );
  NAND2_X1 U13694 ( .A1(n16900), .A2(n10826), .ZN(n10810) );
  XNOR2_X1 U13695 ( .A(n10810), .B(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14755) );
  AND2_X1 U13696 ( .A1(n16075), .A2(n14755), .ZN(n10809) );
  INV_X1 U13697 ( .A(n10810), .ZN(n10811) );
  INV_X1 U13698 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n16258) );
  NAND2_X1 U13699 ( .A1(n10811), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n10812) );
  INV_X1 U13700 ( .A(P2_EBX_REG_24__SCAN_IN), .ZN(n10814) );
  AND2_X1 U13701 ( .A1(n10838), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n10816) );
  AOI21_X1 U13702 ( .B1(n9796), .B2(n10816), .A(n10815), .ZN(n10817) );
  NAND2_X1 U13703 ( .A1(n10822), .A2(n10817), .ZN(n15865) );
  INV_X1 U13704 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n16243) );
  NAND2_X1 U13705 ( .A1(n10818), .A2(n16243), .ZN(n16061) );
  AND2_X1 U13706 ( .A1(n10838), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n10819) );
  NAND2_X1 U13707 ( .A1(n10825), .A2(n10819), .ZN(n10820) );
  OR2_X1 U13708 ( .A1(n10834), .A2(n11790), .ZN(n10821) );
  INV_X1 U13709 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n16222) );
  XNOR2_X1 U13710 ( .A(n10821), .B(n16222), .ZN(n16044) );
  NAND3_X1 U13711 ( .A1(n10822), .A2(P2_EBX_REG_25__SCAN_IN), .A3(n10838), 
        .ZN(n10823) );
  AND3_X1 U13712 ( .A1(n10825), .A2(n10824), .A3(n10823), .ZN(n10835) );
  AOI21_X1 U13713 ( .B1(n10835), .B2(n10826), .A(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n16050) );
  NAND2_X1 U13714 ( .A1(n10829), .A2(n10828), .ZN(n10833) );
  INV_X1 U13715 ( .A(n10845), .ZN(n10830) );
  NAND2_X1 U13716 ( .A1(n10838), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n13029) );
  NAND2_X1 U13717 ( .A1(n10838), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n10831) );
  XNOR2_X1 U13718 ( .A(n13033), .B(n10831), .ZN(n16866) );
  NAND2_X1 U13719 ( .A1(n16866), .A2(n10826), .ZN(n14802) );
  INV_X1 U13720 ( .A(n14802), .ZN(n10832) );
  INV_X1 U13721 ( .A(n10834), .ZN(n16889) );
  NOR2_X1 U13722 ( .A1(n11790), .A2(n16222), .ZN(n10836) );
  INV_X1 U13723 ( .A(n10835), .ZN(n15851) );
  NOR3_X1 U13724 ( .A1(n15851), .A2(n11790), .A3(n10192), .ZN(n16051) );
  AOI21_X1 U13725 ( .B1(n16889), .B2(n10836), .A(n16051), .ZN(n13028) );
  AND2_X1 U13726 ( .A1(n10838), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n10837) );
  NAND2_X1 U13727 ( .A1(n10838), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n10839) );
  XNOR2_X1 U13728 ( .A(n10840), .B(n10839), .ZN(n16854) );
  INV_X1 U13729 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16206) );
  OAI21_X1 U13730 ( .B1(n16854), .B2(n11790), .A(n16206), .ZN(n16028) );
  NOR3_X1 U13731 ( .A1(n16854), .A2(n11790), .A3(n16206), .ZN(n16030) );
  NAND2_X1 U13732 ( .A1(n10838), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n10841) );
  NAND2_X1 U13733 ( .A1(n10840), .A2(n10839), .ZN(n10843) );
  XOR2_X1 U13734 ( .A(n10841), .B(n10843), .Z(n16843) );
  NOR2_X1 U13735 ( .A1(n16843), .A2(n11790), .ZN(n10842) );
  NOR2_X1 U13736 ( .A1(n10842), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11686) );
  NAND2_X1 U13737 ( .A1(n10842), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11687) );
  NOR2_X1 U13738 ( .A1(n10843), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n10844) );
  MUX2_X1 U13739 ( .A(n10845), .B(n10844), .S(n10838), .Z(n12105) );
  NAND2_X1 U13740 ( .A1(n12105), .A2(n10826), .ZN(n10846) );
  XNOR2_X1 U13741 ( .A(n10846), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n10847) );
  XNOR2_X1 U13742 ( .A(n10848), .B(n10847), .ZN(n12055) );
  INV_X1 U13743 ( .A(n10849), .ZN(n11694) );
  OAI21_X1 U13744 ( .B1(n10851), .B2(n11694), .A(n10850), .ZN(n10855) );
  INV_X1 U13745 ( .A(n10852), .ZN(n10853) );
  NAND3_X1 U13746 ( .A1(n10855), .A2(n10854), .A3(n10853), .ZN(n10860) );
  NAND2_X1 U13747 ( .A1(n16520), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n10856) );
  NAND2_X1 U13748 ( .A1(n10857), .A2(n10856), .ZN(n10859) );
  INV_X1 U13749 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n13144) );
  NAND2_X1 U13750 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n13144), .ZN(
        n10858) );
  NAND2_X1 U13751 ( .A1(n10859), .A2(n10858), .ZN(n11706) );
  AND2_X1 U13752 ( .A1(n10860), .A2(n11706), .ZN(n20740) );
  AND2_X1 U13753 ( .A1(n9759), .A2(n20750), .ZN(n12096) );
  INV_X1 U13754 ( .A(n12096), .ZN(n10862) );
  NOR2_X1 U13755 ( .A1(n13737), .A2(n10862), .ZN(n20734) );
  NAND2_X1 U13756 ( .A1(n20740), .A2(n20734), .ZN(n10874) );
  NAND2_X1 U13757 ( .A1(n10864), .A2(n10863), .ZN(n11702) );
  INV_X1 U13758 ( .A(n11693), .ZN(n11696) );
  NAND2_X1 U13759 ( .A1(n11690), .A2(n11696), .ZN(n10868) );
  XNOR2_X1 U13760 ( .A(n11694), .B(n10865), .ZN(n11695) );
  NAND2_X1 U13761 ( .A1(n11690), .A2(n11695), .ZN(n10866) );
  OR2_X1 U13762 ( .A1(n11702), .A2(n10866), .ZN(n10867) );
  OAI21_X1 U13763 ( .B1(n11702), .B2(n10868), .A(n13734), .ZN(n10869) );
  INV_X1 U13764 ( .A(n10869), .ZN(n10871) );
  NAND2_X1 U13765 ( .A1(n10870), .A2(n13144), .ZN(n13140) );
  INV_X1 U13766 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n13115) );
  OAI21_X1 U13767 ( .B1(n14450), .B2(n13140), .A(n13115), .ZN(n20723) );
  MUX2_X1 U13768 ( .A(n10871), .B(n20723), .S(P2_STATE2_REG_1__SCAN_IN), .Z(
        n17081) );
  NOR2_X1 U13769 ( .A1(n13737), .A2(n9759), .ZN(n10872) );
  NAND2_X1 U13770 ( .A1(n17081), .A2(n10872), .ZN(n10873) );
  NAND2_X1 U13771 ( .A1(n10874), .A2(n10873), .ZN(n11726) );
  NAND2_X1 U13772 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n13792), .ZN(n20616) );
  INV_X1 U13773 ( .A(n20616), .ZN(n10875) );
  NAND2_X1 U13774 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n10875), .ZN(n17088) );
  INV_X1 U13775 ( .A(n17088), .ZN(n13139) );
  AND2_X1 U13776 ( .A1(n20750), .A2(n13139), .ZN(n10876) );
  NAND2_X1 U13777 ( .A1(n11726), .A2(n10876), .ZN(n13114) );
  OR2_X1 U13778 ( .A1(n13114), .A2(n9759), .ZN(n16974) );
  NAND2_X1 U13779 ( .A1(n10892), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n14261) );
  OR2_X1 U13780 ( .A1(n14261), .A2(n10695), .ZN(n14383) );
  INV_X1 U13781 ( .A(n14383), .ZN(n10897) );
  INV_X1 U13782 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n10924) );
  NAND2_X1 U13783 ( .A1(n20034), .A2(n10924), .ZN(n10888) );
  INV_X1 U13784 ( .A(n11748), .ZN(n13248) );
  NOR2_X1 U13785 ( .A1(n14877), .A2(n13248), .ZN(n13247) );
  INV_X1 U13786 ( .A(n11756), .ZN(n10879) );
  NAND2_X1 U13787 ( .A1(n13247), .A2(n10879), .ZN(n10881) );
  NAND2_X1 U13788 ( .A1(n14877), .A2(n11748), .ZN(n10880) );
  XNOR2_X1 U13789 ( .A(n10880), .B(n11756), .ZN(n13125) );
  NAND2_X1 U13790 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n13125), .ZN(
        n13124) );
  NAND2_X1 U13791 ( .A1(n10881), .A2(n13124), .ZN(n10883) );
  XNOR2_X1 U13792 ( .A(n13340), .B(n10883), .ZN(n13324) );
  XNOR2_X1 U13793 ( .A(n10882), .B(n11762), .ZN(n13323) );
  NAND2_X1 U13794 ( .A1(n13324), .A2(n13323), .ZN(n10885) );
  NAND2_X1 U13795 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n10883), .ZN(
        n10884) );
  NAND2_X1 U13796 ( .A1(n10885), .A2(n10884), .ZN(n10886) );
  XNOR2_X1 U13797 ( .A(n10886), .B(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n14770) );
  NAND2_X1 U13798 ( .A1(n10886), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10887) );
  OAI21_X1 U13799 ( .B1(n14771), .B2(n14770), .A(n10887), .ZN(n20033) );
  NAND2_X1 U13800 ( .A1(n10888), .A2(n20033), .ZN(n10891) );
  INV_X1 U13801 ( .A(n20034), .ZN(n10889) );
  NAND2_X1 U13802 ( .A1(n10889), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10890) );
  INV_X1 U13803 ( .A(n10892), .ZN(n10893) );
  NAND2_X1 U13804 ( .A1(n10899), .A2(n14261), .ZN(n10895) );
  NAND2_X1 U13805 ( .A1(n10895), .A2(n10900), .ZN(n10904) );
  INV_X1 U13806 ( .A(n10904), .ZN(n10896) );
  NAND2_X1 U13807 ( .A1(n10900), .A2(n14261), .ZN(n10898) );
  INV_X1 U13808 ( .A(n16119), .ZN(n10915) );
  NAND2_X1 U13809 ( .A1(n16148), .A2(n10910), .ZN(n16185) );
  AND2_X1 U13810 ( .A1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n16314) );
  AND2_X1 U13811 ( .A1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n10911) );
  NAND2_X1 U13812 ( .A1(n16314), .A2(n10911), .ZN(n16290) );
  INV_X1 U13813 ( .A(n16290), .ZN(n10912) );
  INV_X1 U13814 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16393) );
  NOR2_X1 U13815 ( .A1(n10722), .A2(n16393), .ZN(n16386) );
  NAND4_X1 U13816 ( .A1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A4(n16386), .ZN(n16313) );
  INV_X1 U13817 ( .A(n16313), .ZN(n16149) );
  NAND3_X1 U13818 ( .A1(n10912), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A3(
        n16149), .ZN(n12004) );
  INV_X1 U13819 ( .A(n16106), .ZN(n16123) );
  NAND2_X1 U13820 ( .A1(n16123), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n14748) );
  NAND2_X1 U13821 ( .A1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n16262) );
  OR2_X1 U13822 ( .A1(n13114), .A2(n20755), .ZN(n20043) );
  INV_X1 U13823 ( .A(n10916), .ZN(n10918) );
  AOI22_X1 U13824 ( .A1(n11026), .A2(P2_EBX_REG_4__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10923) );
  INV_X1 U13825 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n10921) );
  OR2_X1 U13826 ( .A1(n11027), .A2(n10921), .ZN(n10922) );
  OAI211_X1 U13827 ( .C1(n10944), .C2(n10924), .A(n10923), .B(n10922), .ZN(
        n14856) );
  OAI22_X1 U13828 ( .A1(n10925), .A2(n14852), .B1(n13792), .B2(n17014), .ZN(
        n10928) );
  NOR2_X1 U13829 ( .A1(n10944), .A2(n10926), .ZN(n10927) );
  AOI211_X1 U13830 ( .C1(n10929), .C2(P2_REIP_REG_5__SCAN_IN), .A(n10928), .B(
        n10927), .ZN(n14270) );
  INV_X1 U13831 ( .A(n14270), .ZN(n10930) );
  INV_X1 U13832 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n14389) );
  OR2_X1 U13833 ( .A1(n10925), .A2(n10932), .ZN(n10934) );
  NAND2_X1 U13834 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n10933) );
  OAI211_X1 U13835 ( .C1(n11027), .C2(n14389), .A(n10934), .B(n10933), .ZN(
        n10935) );
  AOI21_X1 U13836 ( .B1(n10392), .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n10935), .ZN(n13468) );
  OR2_X1 U13837 ( .A1(n10944), .A2(n10936), .ZN(n10943) );
  INV_X1 U13838 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n10940) );
  INV_X1 U13839 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n10937) );
  OR2_X1 U13840 ( .A1(n10925), .A2(n10937), .ZN(n10939) );
  NAND2_X1 U13841 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n10938) );
  OAI211_X1 U13842 ( .C1(n11027), .C2(n10940), .A(n10939), .B(n10938), .ZN(
        n10941) );
  INV_X1 U13843 ( .A(n10941), .ZN(n10942) );
  NAND2_X1 U13844 ( .A1(n10943), .A2(n10942), .ZN(n13504) );
  AOI22_X1 U13845 ( .A1(n11026), .A2(P2_EBX_REG_8__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10947) );
  INV_X1 U13846 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n10945) );
  OR2_X1 U13847 ( .A1(n11027), .A2(n10945), .ZN(n10946) );
  OAI211_X1 U13848 ( .C1(n10944), .C2(n11984), .A(n10947), .B(n10946), .ZN(
        n13444) );
  INV_X1 U13849 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n14291) );
  NAND2_X1 U13850 ( .A1(n10392), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n10949) );
  AOI22_X1 U13851 ( .A1(n11026), .A2(P2_EBX_REG_9__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n10948) );
  OAI211_X1 U13852 ( .C1(n11027), .C2(n14291), .A(n10949), .B(n10948), .ZN(
        n14285) );
  OR2_X1 U13853 ( .A1(n10944), .A2(n10722), .ZN(n10952) );
  AOI22_X1 U13854 ( .A1(n11026), .A2(P2_EBX_REG_10__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), 
        .ZN(n10951) );
  INV_X1 U13855 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n14248) );
  OR2_X1 U13856 ( .A1(n11027), .A2(n14248), .ZN(n10950) );
  OR2_X1 U13857 ( .A1(n10944), .A2(n16393), .ZN(n10957) );
  OR2_X1 U13858 ( .A1(n10925), .A2(n19958), .ZN(n10954) );
  NAND2_X1 U13859 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n10953) );
  OAI211_X1 U13860 ( .C1(n11027), .C2(n20648), .A(n10954), .B(n10953), .ZN(
        n10955) );
  INV_X1 U13861 ( .A(n10955), .ZN(n10956) );
  NAND2_X1 U13862 ( .A1(n10957), .A2(n10956), .ZN(n16387) );
  INV_X1 U13863 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n11913) );
  INV_X1 U13864 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n10958) );
  OR2_X1 U13865 ( .A1(n10925), .A2(n10958), .ZN(n10960) );
  NAND2_X1 U13866 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n10959) );
  OAI211_X1 U13867 ( .C1(n11027), .C2(n11913), .A(n10960), .B(n10959), .ZN(
        n10961) );
  AOI21_X1 U13868 ( .B1(n10392), .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n10961), .ZN(n16964) );
  INV_X1 U13869 ( .A(n16964), .ZN(n10965) );
  AOI22_X1 U13870 ( .A1(n11026), .A2(P2_EBX_REG_12__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), 
        .ZN(n10964) );
  INV_X1 U13871 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n10962) );
  OR2_X1 U13872 ( .A1(n11027), .A2(n10962), .ZN(n10963) );
  OAI211_X1 U13873 ( .C1(n10944), .C2(n16373), .A(n10964), .B(n10963), .ZN(
        n13643) );
  AND2_X1 U13874 ( .A1(n10965), .A2(n13643), .ZN(n10966) );
  AOI22_X1 U13875 ( .A1(n11026), .A2(P2_EBX_REG_14__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), 
        .ZN(n10969) );
  INV_X1 U13876 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n10967) );
  OR2_X1 U13877 ( .A1(n11027), .A2(n10967), .ZN(n10968) );
  OAI211_X1 U13878 ( .C1(n10944), .C2(n16353), .A(n10969), .B(n10968), .ZN(
        n13715) );
  INV_X1 U13879 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n10972) );
  OR2_X1 U13880 ( .A1(n10925), .A2(n10737), .ZN(n10971) );
  NAND2_X1 U13881 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n10970) );
  OAI211_X1 U13882 ( .C1(n11027), .C2(n10972), .A(n10971), .B(n10970), .ZN(
        n10973) );
  AOI21_X1 U13883 ( .B1(n10392), .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n10973), .ZN(n16945) );
  OR2_X1 U13884 ( .A1(n10944), .A2(n10974), .ZN(n10977) );
  AOI22_X1 U13885 ( .A1(n11026), .A2(P2_EBX_REG_16__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), 
        .ZN(n10976) );
  INV_X1 U13886 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n20654) );
  OR2_X1 U13887 ( .A1(n11027), .A2(n20654), .ZN(n10975) );
  AOI22_X1 U13888 ( .A1(n11026), .A2(P2_EBX_REG_17__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), 
        .ZN(n10979) );
  INV_X1 U13889 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n20656) );
  OR2_X1 U13890 ( .A1(n11027), .A2(n20656), .ZN(n10978) );
  OAI211_X1 U13891 ( .C1(n10944), .C2(n16159), .A(n10979), .B(n10978), .ZN(
        n16162) );
  AOI22_X1 U13892 ( .A1(n11026), .A2(P2_EBX_REG_18__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), 
        .ZN(n10981) );
  INV_X1 U13893 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n20658) );
  OR2_X1 U13894 ( .A1(n11027), .A2(n20658), .ZN(n10980) );
  OAI211_X1 U13895 ( .C1(n10944), .C2(n16320), .A(n10981), .B(n10980), .ZN(
        n14130) );
  NAND2_X1 U13896 ( .A1(n14129), .A2(n14130), .ZN(n14128) );
  OR2_X1 U13897 ( .A1(n10944), .A2(n16307), .ZN(n10985) );
  INV_X1 U13898 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n20660) );
  NOR2_X1 U13899 ( .A1(n11027), .A2(n20660), .ZN(n10983) );
  INV_X1 U13900 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n19768) );
  OAI22_X1 U13901 ( .A1(n10925), .A2(n10747), .B1(n13792), .B2(n19768), .ZN(
        n10982) );
  NOR2_X1 U13902 ( .A1(n10983), .A2(n10982), .ZN(n10984) );
  AND2_X1 U13903 ( .A1(n10985), .A2(n10984), .ZN(n16137) );
  OR2_X1 U13904 ( .A1(n10944), .A2(n16297), .ZN(n10988) );
  AOI22_X1 U13905 ( .A1(n11026), .A2(P2_EBX_REG_20__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), 
        .ZN(n10987) );
  INV_X1 U13906 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n16124) );
  OR2_X1 U13907 ( .A1(n11027), .A2(n16124), .ZN(n10986) );
  AND3_X1 U13908 ( .A1(n10988), .A2(n10987), .A3(n10986), .ZN(n14436) );
  OR2_X1 U13909 ( .A1(n10944), .A2(n16280), .ZN(n10994) );
  INV_X1 U13910 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n20663) );
  NOR2_X1 U13911 ( .A1(n11027), .A2(n20663), .ZN(n10992) );
  INV_X1 U13912 ( .A(P2_EBX_REG_21__SCAN_IN), .ZN(n10990) );
  OAI22_X1 U13913 ( .A1(n10925), .A2(n10990), .B1(n13792), .B2(n10085), .ZN(
        n10991) );
  NOR2_X1 U13914 ( .A1(n10992), .A2(n10991), .ZN(n10993) );
  AOI22_X1 U13915 ( .A1(n11019), .A2(P2_EBX_REG_22__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), 
        .ZN(n10997) );
  INV_X1 U13916 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n10995) );
  OR2_X1 U13917 ( .A1(n11027), .A2(n10995), .ZN(n10996) );
  OAI211_X1 U13918 ( .C1(n10944), .C2(n16273), .A(n10997), .B(n10996), .ZN(
        n15925) );
  INV_X1 U13919 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n20666) );
  OR2_X1 U13920 ( .A1(n10925), .A2(n9940), .ZN(n10999) );
  NAND2_X1 U13921 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n10998) );
  OAI211_X1 U13922 ( .C1(n11027), .C2(n20666), .A(n10999), .B(n10998), .ZN(
        n11000) );
  AOI21_X1 U13923 ( .B1(n10392), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n11000), .ZN(n14750) );
  OR2_X1 U13924 ( .A1(n10944), .A2(n16243), .ZN(n11003) );
  AOI22_X1 U13925 ( .A1(n11026), .A2(P2_EBX_REG_24__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), 
        .ZN(n11002) );
  INV_X1 U13926 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n20668) );
  OR2_X1 U13927 ( .A1(n11027), .A2(n20668), .ZN(n11001) );
  AND3_X1 U13928 ( .A1(n11003), .A2(n11002), .A3(n11001), .ZN(n15854) );
  OR2_X1 U13929 ( .A1(n10944), .A2(n10192), .ZN(n11008) );
  INV_X1 U13930 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n20670) );
  NOR2_X1 U13931 ( .A1(n11027), .A2(n20670), .ZN(n11006) );
  INV_X1 U13932 ( .A(P2_EBX_REG_25__SCAN_IN), .ZN(n11004) );
  INV_X1 U13933 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n15841) );
  OAI22_X1 U13934 ( .A1(n10925), .A2(n11004), .B1(n13792), .B2(n15841), .ZN(
        n11005) );
  NOR2_X1 U13935 ( .A1(n11006), .A2(n11005), .ZN(n11007) );
  NAND2_X1 U13936 ( .A1(n11008), .A2(n11007), .ZN(n15846) );
  AOI22_X1 U13937 ( .A1(n11019), .A2(P2_EBX_REG_26__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), 
        .ZN(n11010) );
  INV_X1 U13938 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n20672) );
  OR2_X1 U13939 ( .A1(n11027), .A2(n20672), .ZN(n11009) );
  OAI211_X1 U13940 ( .C1(n10944), .C2(n16222), .A(n11010), .B(n11009), .ZN(
        n15910) );
  OR2_X1 U13941 ( .A1(n10944), .A2(n10829), .ZN(n11015) );
  INV_X1 U13942 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n20675) );
  NOR2_X1 U13943 ( .A1(n11027), .A2(n20675), .ZN(n11013) );
  INV_X1 U13944 ( .A(P2_EBX_REG_27__SCAN_IN), .ZN(n11011) );
  OAI22_X1 U13945 ( .A1(n10925), .A2(n11011), .B1(n13792), .B2(n10080), .ZN(
        n11012) );
  NOR2_X1 U13946 ( .A1(n11013), .A2(n11012), .ZN(n11014) );
  AND2_X1 U13947 ( .A1(n11015), .A2(n11014), .ZN(n13037) );
  OR2_X1 U13948 ( .A1(n10944), .A2(n10828), .ZN(n11018) );
  AOI22_X1 U13949 ( .A1(n11026), .A2(P2_EBX_REG_28__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), 
        .ZN(n11017) );
  INV_X1 U13950 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n20676) );
  OR2_X1 U13951 ( .A1(n11027), .A2(n20676), .ZN(n11016) );
  AND3_X1 U13952 ( .A1(n11018), .A2(n11017), .A3(n11016), .ZN(n14809) );
  AOI22_X1 U13953 ( .A1(n11019), .A2(P2_EBX_REG_29__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), 
        .ZN(n11021) );
  INV_X1 U13954 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n20678) );
  OR2_X1 U13955 ( .A1(n11027), .A2(n20678), .ZN(n11020) );
  OAI211_X1 U13956 ( .C1(n10944), .C2(n16206), .A(n11021), .B(n11020), .ZN(
        n15893) );
  INV_X1 U13957 ( .A(n15892), .ZN(n11025) );
  AOI22_X1 U13958 ( .A1(n11026), .A2(P2_EBX_REG_30__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), 
        .ZN(n11024) );
  INV_X1 U13959 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n11022) );
  OR2_X1 U13960 ( .A1(n11027), .A2(n11022), .ZN(n11023) );
  OAI211_X1 U13961 ( .C1(n10944), .C2(n12027), .A(n11024), .B(n11023), .ZN(
        n11731) );
  INV_X1 U13962 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n12057) );
  AOI22_X1 U13963 ( .A1(n11026), .A2(P2_EBX_REG_31__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n11029) );
  INV_X1 U13964 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n20683) );
  OR2_X1 U13965 ( .A1(n11027), .A2(n20683), .ZN(n11028) );
  OAI211_X1 U13966 ( .C1(n10944), .C2(n12057), .A(n11029), .B(n11028), .ZN(
        n11030) );
  INV_X1 U13967 ( .A(n11030), .ZN(n11031) );
  INV_X1 U13968 ( .A(n20699), .ZN(n20509) );
  NAND2_X1 U13969 ( .A1(n13792), .A2(n20333), .ZN(n20696) );
  NAND2_X1 U13970 ( .A1(n20509), .A2(n20696), .ZN(n20722) );
  NAND2_X1 U13971 ( .A1(n20722), .A2(n20749), .ZN(n11032) );
  AND2_X1 U13972 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n20713) );
  AND2_X1 U13973 ( .A1(n20749), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n13419) );
  INV_X1 U13974 ( .A(n13419), .ZN(n11035) );
  INV_X1 U13975 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n11033) );
  NAND2_X1 U13976 ( .A1(n11033), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n11034) );
  NAND2_X1 U13977 ( .A1(n11035), .A2(n11034), .ZN(n13252) );
  INV_X1 U13978 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n17007) );
  INV_X1 U13979 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n16986) );
  INV_X1 U13980 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n16971) );
  INV_X1 U13981 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n19816) );
  INV_X1 U13982 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n16161) );
  NAND2_X1 U13983 ( .A1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n12075), .ZN(
        n12074) );
  INV_X1 U13984 ( .A(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n16082) );
  NAND2_X1 U13985 ( .A1(n12080), .A2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n12079) );
  INV_X1 U13986 ( .A(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n16068) );
  INV_X1 U13987 ( .A(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n12085) );
  INV_X1 U13988 ( .A(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n12089) );
  INV_X1 U13989 ( .A(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n16035) );
  INV_X1 U13990 ( .A(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n11038) );
  INV_X1 U13991 ( .A(n12056), .ZN(n11040) );
  INV_X1 U13992 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n20607) );
  NAND2_X1 U13993 ( .A1(n20749), .A2(n20607), .ZN(n11037) );
  OR2_X1 U13994 ( .A1(n20696), .A2(n11037), .ZN(n12009) );
  INV_X1 U13995 ( .A(n12009), .ZN(n19905) );
  NAND2_X1 U13996 ( .A1(n19905), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n12042) );
  OAI21_X1 U13997 ( .B1(n20055), .B2(n11038), .A(n12042), .ZN(n11039) );
  AOI21_X1 U13998 ( .B1(n17008), .B2(n11040), .A(n11039), .ZN(n11041) );
  OAI21_X1 U13999 ( .B1(n12055), .B2(n16974), .A(n11042), .ZN(P2_U2983) );
  AND2_X4 U14000 ( .A1(n13599), .A2(n15828), .ZN(n11390) );
  AOI22_X1 U14001 ( .A1(n11390), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11098), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11048) );
  AND2_X2 U14002 ( .A1(n11049), .A2(n11044), .ZN(n11223) );
  AOI22_X1 U14003 ( .A1(n11223), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n9764), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11047) );
  AND2_X2 U14004 ( .A1(n11051), .A2(n11044), .ZN(n11153) );
  AOI22_X1 U14005 ( .A1(n11153), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n9749), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11046) );
  AOI22_X1 U14006 ( .A1(n11385), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n9756), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11056) );
  AOI22_X1 U14007 ( .A1(n11162), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11158), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11055) );
  AND2_X4 U14008 ( .A1(n11051), .A2(n13599), .ZN(n11222) );
  AOI22_X1 U14009 ( .A1(n11222), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12395), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11054) );
  AOI22_X1 U14010 ( .A1(n11159), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11163), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11053) );
  AOI22_X1 U14011 ( .A1(n12588), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12606), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11058) );
  INV_X1 U14012 ( .A(n11058), .ZN(n11063) );
  AOI22_X1 U14013 ( .A1(n11223), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n9764), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11061) );
  AOI22_X1 U14014 ( .A1(n11153), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n9749), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11060) );
  AOI22_X1 U14015 ( .A1(n11390), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11098), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11059) );
  NAND3_X1 U14016 ( .A1(n11061), .A2(n11060), .A3(n11059), .ZN(n11062) );
  AOI22_X1 U14017 ( .A1(n11385), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n9756), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11067) );
  AOI22_X1 U14018 ( .A1(n11162), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11158), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11066) );
  AOI22_X1 U14019 ( .A1(n11222), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12395), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11065) );
  AOI22_X1 U14020 ( .A1(n11159), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11163), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11064) );
  AOI22_X1 U14021 ( .A1(n11098), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12612), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11072) );
  AOI22_X1 U14022 ( .A1(n11385), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n9755), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11071) );
  AOI22_X1 U14023 ( .A1(n11153), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n12606), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11070) );
  AOI22_X1 U14024 ( .A1(n11159), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n9738), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11069) );
  AOI22_X1 U14025 ( .A1(n9743), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11158), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11076) );
  AOI22_X1 U14026 ( .A1(n11390), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11223), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11075) );
  AOI22_X1 U14027 ( .A1(n11238), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n12588), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11074) );
  AOI22_X1 U14028 ( .A1(n11222), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11163), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11073) );
  INV_X2 U14029 ( .A(n14704), .ZN(n13875) );
  NAND2_X1 U14030 ( .A1(n11385), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n11080) );
  NAND2_X1 U14031 ( .A1(n9756), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n11079) );
  NAND2_X1 U14032 ( .A1(n11162), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n11078) );
  NAND2_X1 U14033 ( .A1(n11158), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n11077) );
  NAND2_X1 U14034 ( .A1(n11222), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n11084) );
  NAND2_X1 U14035 ( .A1(n11159), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n11083) );
  NAND2_X1 U14036 ( .A1(n9738), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n11082) );
  NAND2_X1 U14037 ( .A1(n11163), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n11081) );
  NAND2_X1 U14038 ( .A1(n11390), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n11088) );
  NAND2_X1 U14039 ( .A1(n11223), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n11087) );
  NAND2_X1 U14040 ( .A1(n11098), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n11086) );
  NAND2_X1 U14041 ( .A1(n12612), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n11085) );
  NAND2_X1 U14042 ( .A1(n12588), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n11092) );
  NAND2_X1 U14043 ( .A1(n11153), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n11091) );
  NAND2_X1 U14044 ( .A1(n9750), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n11090) );
  NAND2_X1 U14045 ( .A1(n9741), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n11089) );
  NAND2_X1 U14046 ( .A1(n13875), .A2(n11129), .ZN(n11097) );
  AOI22_X1 U14047 ( .A1(n11153), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n11098), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11102) );
  AOI22_X1 U14048 ( .A1(n11158), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12395), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11101) );
  AOI22_X1 U14049 ( .A1(n11238), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n9741), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11100) );
  AOI22_X1 U14050 ( .A1(n11222), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11163), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11099) );
  AOI22_X1 U14051 ( .A1(n11385), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n9755), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11106) );
  AOI22_X1 U14052 ( .A1(n11159), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n9742), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11105) );
  AOI22_X1 U14053 ( .A1(n11390), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n9744), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11104) );
  AOI22_X1 U14054 ( .A1(n11223), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n12612), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11103) );
  NAND2_X2 U14055 ( .A1(n11107), .A2(n10227), .ZN(n13049) );
  NAND2_X1 U14056 ( .A1(n13875), .A2(n13049), .ZN(n11128) );
  NAND2_X1 U14057 ( .A1(n11385), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n11111) );
  NAND2_X1 U14058 ( .A1(n9756), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n11110) );
  NAND2_X1 U14059 ( .A1(n11162), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n11109) );
  NAND2_X1 U14060 ( .A1(n11158), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n11108) );
  NAND2_X1 U14061 ( .A1(n11153), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n11115) );
  NAND2_X1 U14062 ( .A1(n12588), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n11114) );
  NAND2_X1 U14063 ( .A1(n9750), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n11113) );
  NAND2_X1 U14064 ( .A1(n9741), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n11112) );
  NAND2_X1 U14065 ( .A1(n11390), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n11119) );
  NAND2_X1 U14066 ( .A1(n11098), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n11118) );
  NAND2_X1 U14067 ( .A1(n11223), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n11117) );
  NAND2_X1 U14068 ( .A1(n11222), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n11123) );
  NAND2_X1 U14069 ( .A1(n11159), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n11122) );
  NAND2_X1 U14070 ( .A1(n12395), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n11121) );
  NAND2_X1 U14071 ( .A1(n11163), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n11120) );
  AND2_X2 U14072 ( .A1(n11128), .A2(n13392), .ZN(n11191) );
  INV_X2 U14073 ( .A(n13049), .ZN(n11199) );
  NAND2_X2 U14074 ( .A1(n11199), .A2(n14704), .ZN(n13393) );
  INV_X1 U14075 ( .A(n13393), .ZN(n11130) );
  INV_X1 U14076 ( .A(n11677), .ZN(n11129) );
  NAND2_X1 U14077 ( .A1(n11130), .A2(n11129), .ZN(n11131) );
  AND2_X2 U14078 ( .A1(n11191), .A2(n11131), .ZN(n11561) );
  AND2_X2 U14079 ( .A1(n11132), .A2(n11561), .ZN(n11539) );
  NAND2_X1 U14080 ( .A1(n11385), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n11136) );
  NAND2_X1 U14081 ( .A1(n9756), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n11135) );
  NAND2_X1 U14082 ( .A1(n11162), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n11134) );
  NAND2_X1 U14083 ( .A1(n11158), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n11133) );
  NAND2_X1 U14084 ( .A1(n11222), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n11140) );
  NAND2_X1 U14085 ( .A1(n11159), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n11139) );
  NAND2_X1 U14086 ( .A1(n9738), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n11138) );
  NAND2_X1 U14087 ( .A1(n9737), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n11137) );
  NAND2_X1 U14088 ( .A1(n11390), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n11144) );
  NAND2_X1 U14089 ( .A1(n11098), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n11143) );
  NAND2_X1 U14090 ( .A1(n11223), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n11142) );
  NAND2_X1 U14091 ( .A1(n11153), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n11148) );
  NAND2_X1 U14092 ( .A1(n12588), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n11147) );
  NAND2_X1 U14093 ( .A1(n9749), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n11146) );
  NAND4_X4 U14094 ( .A1(n11152), .A2(n11151), .A3(n11150), .A4(n11149), .ZN(
        n11192) );
  NAND2_X1 U14095 ( .A1(n11539), .A2(n11192), .ZN(n11547) );
  NAND2_X1 U14096 ( .A1(n9755), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n11157) );
  NAND2_X1 U14097 ( .A1(n11153), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n11156) );
  NAND2_X1 U14098 ( .A1(n11223), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n11155) );
  NAND2_X1 U14099 ( .A1(n12612), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n11154) );
  NAND2_X1 U14100 ( .A1(n11222), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n11167) );
  NAND2_X1 U14101 ( .A1(n11162), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n11166) );
  NAND2_X1 U14102 ( .A1(n12588), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n11165) );
  NAND2_X1 U14103 ( .A1(n11163), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n11164) );
  NAND2_X1 U14104 ( .A1(n11390), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n11171) );
  NAND2_X1 U14105 ( .A1(n11098), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n11170) );
  NAND2_X1 U14106 ( .A1(n12606), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n11169) );
  NAND2_X1 U14107 ( .A1(n9750), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11168) );
  INV_X1 U14108 ( .A(P1_STATE_REG_1__SCAN_IN), .ZN(n21180) );
  XNOR2_X1 U14109 ( .A(n21180), .B(P1_STATE_REG_2__SCAN_IN), .ZN(n11486) );
  NAND2_X1 U14110 ( .A1(n13392), .A2(n11677), .ZN(n11185) );
  AND2_X1 U14111 ( .A1(n13049), .A2(n14704), .ZN(n11175) );
  NAND2_X2 U14112 ( .A1(n11176), .A2(n14704), .ZN(n11553) );
  NAND2_X1 U14113 ( .A1(n11488), .A2(n13951), .ZN(n11550) );
  NOR2_X2 U14114 ( .A1(n11177), .A2(n11192), .ZN(n11194) );
  OAI211_X1 U14115 ( .C1(n11547), .C2(n11180), .A(n11550), .B(n11548), .ZN(
        n11181) );
  NAND2_X1 U14116 ( .A1(n11181), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11257) );
  NAND2_X1 U14117 ( .A1(n11487), .A2(n11192), .ZN(n11555) );
  OAI211_X1 U14118 ( .C1(n11553), .C2(n11195), .A(n10205), .B(n11555), .ZN(
        n11183) );
  INV_X1 U14119 ( .A(n11183), .ZN(n11184) );
  NAND2_X1 U14120 ( .A1(n11191), .A2(n10206), .ZN(n11490) );
  NAND2_X1 U14121 ( .A1(n11206), .A2(n11186), .ZN(n11188) );
  NOR2_X1 U14122 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n21270) );
  NAND2_X1 U14123 ( .A1(n21270), .A2(n9954), .ZN(n12636) );
  MUX2_X1 U14124 ( .A(n11537), .B(n12636), .S(n21110), .Z(n11190) );
  AOI21_X1 U14125 ( .B1(n11191), .B2(n13951), .A(n11194), .ZN(n11204) );
  NAND2_X1 U14126 ( .A1(n11193), .A2(n13275), .ZN(n11203) );
  INV_X1 U14127 ( .A(n11194), .ZN(n11196) );
  INV_X1 U14128 ( .A(n11198), .ZN(n13306) );
  NAND2_X1 U14129 ( .A1(n13306), .A2(n11199), .ZN(n11565) );
  AOI22_X1 U14130 ( .A1(n12607), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n11278), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11210) );
  AOI22_X1 U14131 ( .A1(n9715), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12603), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11209) );
  AOI22_X1 U14132 ( .A1(n12413), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n12614), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11208) );
  AOI22_X1 U14133 ( .A1(n12588), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n12606), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11207) );
  NAND4_X1 U14134 ( .A1(n11210), .A2(n11209), .A3(n11208), .A4(n11207), .ZN(
        n11216) );
  AOI22_X1 U14135 ( .A1(n11390), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11098), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11214) );
  AOI22_X1 U14137 ( .A1(n9762), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n9756), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11213) );
  AOI22_X1 U14138 ( .A1(n12604), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n9764), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11212) );
  AOI22_X1 U14139 ( .A1(n9738), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n11163), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11211) );
  NAND4_X1 U14140 ( .A1(n11214), .A2(n11213), .A3(n11212), .A4(n11211), .ZN(
        n11215) );
  NOR2_X1 U14141 ( .A1(n11277), .A2(n11423), .ZN(n11245) );
  AOI22_X1 U14142 ( .A1(n12603), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11217), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11221) );
  AOI22_X1 U14143 ( .A1(n9715), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n9762), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11220) );
  AOI22_X1 U14144 ( .A1(n11390), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12539), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11219) );
  INV_X1 U14145 ( .A(n13597), .ZN(n12613) );
  AOI22_X1 U14146 ( .A1(n12613), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n9764), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11218) );
  NAND4_X1 U14147 ( .A1(n11221), .A2(n11220), .A3(n11219), .A4(n11218), .ZN(
        n11229) );
  BUF_X1 U14148 ( .A(n11222), .Z(n11278) );
  AOI22_X1 U14149 ( .A1(n11278), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12395), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11227) );
  AOI22_X1 U14150 ( .A1(n12413), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n11223), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11226) );
  BUF_X1 U14151 ( .A(n9750), .Z(n12614) );
  AOI22_X1 U14152 ( .A1(n12614), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n9741), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11225) );
  AOI22_X1 U14153 ( .A1(n12607), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n11163), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11224) );
  NAND4_X1 U14154 ( .A1(n11227), .A2(n11226), .A3(n11225), .A4(n11224), .ZN(
        n11228) );
  NAND2_X1 U14155 ( .A1(n11245), .A2(n11309), .ZN(n11230) );
  INV_X1 U14156 ( .A(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11233) );
  AOI21_X1 U14157 ( .B1(n11129), .B2(n11423), .A(n9954), .ZN(n11232) );
  NAND2_X1 U14158 ( .A1(n13936), .A2(n11309), .ZN(n11231) );
  OAI211_X1 U14159 ( .C1(n11520), .C2(n11233), .A(n11232), .B(n11231), .ZN(
        n11307) );
  INV_X1 U14160 ( .A(n11277), .ZN(n11258) );
  NAND2_X1 U14161 ( .A1(n11258), .A2(n11423), .ZN(n11442) );
  AOI22_X1 U14162 ( .A1(n12413), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n12605), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11237) );
  AOI22_X1 U14163 ( .A1(n9715), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12603), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11236) );
  AOI22_X1 U14164 ( .A1(n11217), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n12539), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11235) );
  AOI22_X1 U14165 ( .A1(n12607), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n11163), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11234) );
  NAND4_X1 U14166 ( .A1(n11237), .A2(n11236), .A3(n11235), .A4(n11234), .ZN(
        n11244) );
  AOI22_X1 U14167 ( .A1(n11278), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n9738), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11242) );
  AOI22_X1 U14168 ( .A1(n11223), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n9764), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11241) );
  AOI22_X1 U14169 ( .A1(n12613), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12614), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11240) );
  AOI22_X1 U14170 ( .A1(n9762), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12606), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11239) );
  NAND4_X1 U14171 ( .A1(n11242), .A2(n11241), .A3(n11240), .A4(n11239), .ZN(
        n11243) );
  INV_X1 U14172 ( .A(n11303), .ZN(n11248) );
  INV_X1 U14173 ( .A(n11245), .ZN(n11247) );
  NAND2_X1 U14174 ( .A1(n11529), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11246) );
  OAI211_X1 U14175 ( .C1(n11429), .C2(n11248), .A(n11247), .B(n11246), .ZN(
        n11249) );
  NAND2_X1 U14176 ( .A1(n11250), .A2(n11249), .ZN(n11251) );
  INV_X1 U14177 ( .A(n11252), .ZN(n11253) );
  INV_X1 U14178 ( .A(n12636), .ZN(n11319) );
  NAND2_X1 U14179 ( .A1(n21009), .A2(n21110), .ZN(n11255) );
  NAND2_X1 U14180 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n11270) );
  AND2_X1 U14181 ( .A1(n11255), .A2(n11270), .ZN(n14491) );
  INV_X1 U14182 ( .A(n11537), .ZN(n11318) );
  AND2_X1 U14183 ( .A1(n11318), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n11261) );
  AOI21_X1 U14184 ( .B1(n11319), .B2(n14491), .A(n11261), .ZN(n11256) );
  NAND2_X1 U14185 ( .A1(n11258), .A2(n11303), .ZN(n11259) );
  INV_X1 U14186 ( .A(n11295), .ZN(n11293) );
  INV_X1 U14187 ( .A(n11261), .ZN(n11263) );
  NAND2_X1 U14188 ( .A1(n11263), .A2(n11262), .ZN(n11264) );
  NAND2_X1 U14189 ( .A1(n11265), .A2(n11264), .ZN(n11266) );
  NAND2_X1 U14190 ( .A1(n11268), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11273) );
  INV_X1 U14191 ( .A(n11270), .ZN(n11269) );
  NAND2_X1 U14192 ( .A1(n11269), .A2(n20941), .ZN(n14057) );
  NAND2_X1 U14193 ( .A1(n11270), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n11271) );
  NAND2_X1 U14194 ( .A1(n14057), .A2(n11271), .ZN(n14007) );
  AOI22_X1 U14195 ( .A1(n11319), .A2(n14007), .B1(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n11318), .ZN(n11272) );
  AOI22_X1 U14196 ( .A1(n12413), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n12603), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11282) );
  AOI22_X1 U14197 ( .A1(n11278), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n9762), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11281) );
  AOI22_X1 U14198 ( .A1(n11390), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12604), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11280) );
  AOI22_X1 U14199 ( .A1(n12607), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11163), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11279) );
  NAND4_X1 U14200 ( .A1(n11282), .A2(n11281), .A3(n11280), .A4(n11279), .ZN(
        n11288) );
  AOI22_X1 U14201 ( .A1(n9715), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12395), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11286) );
  AOI22_X1 U14202 ( .A1(n11217), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12539), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11285) );
  AOI22_X1 U14203 ( .A1(n12613), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n9764), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11284) );
  AOI22_X1 U14204 ( .A1(n12614), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n9741), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11283) );
  NAND4_X1 U14205 ( .A1(n11286), .A2(n11285), .A3(n11284), .A4(n11283), .ZN(
        n11287) );
  OR2_X1 U14206 ( .A1(n11288), .A2(n11287), .ZN(n11297) );
  AOI22_X1 U14207 ( .A1(n11500), .A2(n11297), .B1(n11529), .B2(
        P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11289) );
  INV_X1 U14208 ( .A(n11289), .ZN(n11290) );
  INV_X1 U14209 ( .A(n11294), .ZN(n11292) );
  NAND2_X2 U14210 ( .A1(n11293), .A2(n11292), .ZN(n11335) );
  NAND2_X1 U14211 ( .A1(n11295), .A2(n11294), .ZN(n11296) );
  INV_X1 U14212 ( .A(n11494), .ZN(n11412) );
  INV_X1 U14213 ( .A(n11297), .ZN(n11299) );
  NAND2_X1 U14214 ( .A1(n11303), .A2(n11309), .ZN(n11298) );
  NAND2_X1 U14215 ( .A1(n11298), .A2(n11299), .ZN(n11356) );
  OAI21_X1 U14216 ( .B1(n11299), .B2(n11298), .A(n11356), .ZN(n11301) );
  INV_X1 U14217 ( .A(n13649), .ZN(n16495) );
  NAND2_X1 U14218 ( .A1(n13936), .A2(n11554), .ZN(n11308) );
  INV_X1 U14219 ( .A(n11308), .ZN(n11300) );
  AOI21_X1 U14220 ( .B1(n11301), .B2(n16495), .A(n11300), .ZN(n11302) );
  OAI21_X2 U14221 ( .B1(n13856), .B2(n11412), .A(n11302), .ZN(n13455) );
  XNOR2_X1 U14222 ( .A(n11303), .B(n11309), .ZN(n11304) );
  INV_X1 U14223 ( .A(n11567), .ZN(n11545) );
  OAI211_X1 U14224 ( .C1(n11304), .C2(n13649), .A(n11545), .B(n14704), .ZN(
        n11305) );
  INV_X1 U14225 ( .A(n11305), .ZN(n11306) );
  NAND2_X1 U14226 ( .A1(n12170), .A2(n11494), .ZN(n11312) );
  OAI21_X1 U14227 ( .B1(n13649), .B2(n11309), .A(n11308), .ZN(n11310) );
  INV_X1 U14228 ( .A(n11310), .ZN(n11311) );
  NAND2_X2 U14229 ( .A1(n13474), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13476) );
  INV_X1 U14230 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n11590) );
  NAND2_X1 U14231 ( .A1(n13455), .A2(n13456), .ZN(n11316) );
  NAND2_X1 U14232 ( .A1(n11314), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11315) );
  INV_X1 U14233 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n11317) );
  NAND2_X1 U14234 ( .A1(n11268), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11321) );
  NOR3_X1 U14235 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n20941), .A3(
        n21009), .ZN(n13868) );
  NAND2_X1 U14236 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n13868), .ZN(
        n13859) );
  NAND3_X1 U14237 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n14490) );
  NOR2_X1 U14238 ( .A1(n21110), .A2(n14490), .ZN(n14315) );
  AOI21_X1 U14239 ( .B1(n21010), .B2(n13859), .A(n14315), .ZN(n20947) );
  AOI22_X1 U14240 ( .A1(n11319), .A2(n20947), .B1(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n11318), .ZN(n11320) );
  XNOR2_X2 U14241 ( .A(n13294), .B(n13860), .ZN(n14055) );
  AOI22_X1 U14242 ( .A1(n12603), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11217), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11326) );
  AOI22_X1 U14243 ( .A1(n9715), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n9762), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11325) );
  AOI22_X1 U14244 ( .A1(n11278), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12395), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11324) );
  AOI22_X1 U14245 ( .A1(n12607), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n9737), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11323) );
  NAND4_X1 U14246 ( .A1(n11326), .A2(n11325), .A3(n11324), .A4(n11323), .ZN(
        n11332) );
  AOI22_X1 U14247 ( .A1(n11390), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12613), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11330) );
  AOI22_X1 U14248 ( .A1(n12604), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n9764), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11329) );
  AOI22_X1 U14249 ( .A1(n12413), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n12614), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11328) );
  AOI22_X1 U14250 ( .A1(n12539), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12606), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11327) );
  NAND4_X1 U14251 ( .A1(n11330), .A2(n11329), .A3(n11328), .A4(n11327), .ZN(
        n11331) );
  AOI22_X1 U14252 ( .A1(n11500), .A2(n11355), .B1(n11529), .B2(
        P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11333) );
  AND2_X1 U14253 ( .A1(n11335), .A2(n14088), .ZN(n11336) );
  XNOR2_X1 U14254 ( .A(n11356), .B(n11355), .ZN(n11337) );
  OAI22_X1 U14255 ( .A1(n15813), .A2(n11412), .B1(n13649), .B2(n11337), .ZN(
        n13554) );
  NAND2_X1 U14256 ( .A1(n13553), .A2(n13554), .ZN(n11340) );
  NAND2_X1 U14257 ( .A1(n11338), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11339) );
  INV_X1 U14258 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n11341) );
  AOI22_X1 U14259 ( .A1(n11385), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n11217), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11345) );
  AOI22_X1 U14260 ( .A1(n9715), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n9762), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11344) );
  AOI22_X1 U14261 ( .A1(n11278), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n9738), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11343) );
  AOI22_X1 U14262 ( .A1(n12607), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n11163), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11342) );
  NAND4_X1 U14263 ( .A1(n11345), .A2(n11344), .A3(n11343), .A4(n11342), .ZN(
        n11351) );
  AOI22_X1 U14264 ( .A1(n11390), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11098), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11349) );
  AOI22_X1 U14265 ( .A1(n12604), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n9745), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11348) );
  AOI22_X1 U14266 ( .A1(n12413), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n12614), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11347) );
  AOI22_X1 U14267 ( .A1(n12539), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n9741), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11346) );
  NAND4_X1 U14268 ( .A1(n11349), .A2(n11348), .A3(n11347), .A4(n11346), .ZN(
        n11350) );
  NAND2_X1 U14269 ( .A1(n11500), .A2(n11379), .ZN(n11353) );
  NAND2_X1 U14270 ( .A1(n11529), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n11352) );
  NAND2_X1 U14271 ( .A1(n11353), .A2(n11352), .ZN(n11363) );
  INV_X1 U14272 ( .A(n11363), .ZN(n11354) );
  XNOR2_X1 U14273 ( .A(n11364), .B(n11354), .ZN(n12193) );
  NAND2_X1 U14274 ( .A1(n12193), .A2(n11494), .ZN(n11360) );
  AND2_X1 U14275 ( .A1(n11356), .A2(n11355), .ZN(n11380) );
  INV_X1 U14276 ( .A(n11379), .ZN(n11357) );
  XNOR2_X1 U14277 ( .A(n11380), .B(n11357), .ZN(n11358) );
  NAND2_X1 U14278 ( .A1(n11358), .A2(n16495), .ZN(n11359) );
  NAND2_X1 U14279 ( .A1(n11360), .A2(n11359), .ZN(n13730) );
  NAND2_X1 U14280 ( .A1(n11361), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11362) );
  AOI22_X1 U14281 ( .A1(n12607), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11278), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11368) );
  AOI22_X1 U14282 ( .A1(n12605), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n9762), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11367) );
  AOI22_X1 U14283 ( .A1(n12603), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12539), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11366) );
  AOI22_X1 U14284 ( .A1(n12606), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11163), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11365) );
  NAND4_X1 U14285 ( .A1(n11368), .A2(n11367), .A3(n11366), .A4(n11365), .ZN(
        n11374) );
  AOI22_X1 U14286 ( .A1(n11217), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n9760), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11372) );
  AOI22_X1 U14287 ( .A1(n9715), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12604), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11371) );
  AOI22_X1 U14288 ( .A1(n12413), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n12614), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11370) );
  AOI22_X1 U14289 ( .A1(n12613), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n9764), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11369) );
  NAND4_X1 U14290 ( .A1(n11372), .A2(n11371), .A3(n11370), .A4(n11369), .ZN(
        n11373) );
  NAND2_X1 U14291 ( .A1(n11500), .A2(n11401), .ZN(n11376) );
  NAND2_X1 U14292 ( .A1(n11529), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n11375) );
  NAND2_X1 U14293 ( .A1(n11376), .A2(n11375), .ZN(n11377) );
  NAND2_X1 U14294 ( .A1(n11380), .A2(n11379), .ZN(n11402) );
  XNOR2_X1 U14295 ( .A(n11401), .B(n11402), .ZN(n11381) );
  NAND2_X1 U14296 ( .A1(n16495), .A2(n11381), .ZN(n11382) );
  OAI21_X1 U14297 ( .B1(n12208), .B2(n11412), .A(n11382), .ZN(n11384) );
  INV_X1 U14298 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n11383) );
  AOI22_X1 U14299 ( .A1(n11385), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11217), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11389) );
  AOI22_X1 U14300 ( .A1(n9715), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n9762), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11388) );
  AOI22_X1 U14301 ( .A1(n11278), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n9760), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11387) );
  AOI22_X1 U14302 ( .A1(n12607), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n9737), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11386) );
  NAND4_X1 U14303 ( .A1(n11389), .A2(n11388), .A3(n11387), .A4(n11386), .ZN(
        n11396) );
  AOI22_X1 U14304 ( .A1(n11390), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11098), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11394) );
  AOI22_X1 U14305 ( .A1(n12604), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n9745), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11393) );
  AOI22_X1 U14306 ( .A1(n12413), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n12614), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11392) );
  AOI22_X1 U14307 ( .A1(n12539), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n9741), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11391) );
  NAND4_X1 U14308 ( .A1(n11394), .A2(n11393), .A3(n11392), .A4(n11391), .ZN(
        n11395) );
  OR2_X1 U14309 ( .A1(n11396), .A2(n11395), .ZN(n11414) );
  NAND2_X1 U14310 ( .A1(n11500), .A2(n11414), .ZN(n11398) );
  NAND2_X1 U14311 ( .A1(n11529), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n11397) );
  NAND2_X1 U14312 ( .A1(n11398), .A2(n11397), .ZN(n11399) );
  NAND2_X1 U14313 ( .A1(n11444), .A2(n12209), .ZN(n11407) );
  INV_X1 U14314 ( .A(n11401), .ZN(n11403) );
  NOR2_X1 U14315 ( .A1(n11403), .A2(n11402), .ZN(n11413) );
  INV_X1 U14316 ( .A(n11413), .ZN(n11404) );
  XNOR2_X1 U14317 ( .A(n11414), .B(n11404), .ZN(n11405) );
  NAND2_X1 U14318 ( .A1(n16495), .A2(n11405), .ZN(n11406) );
  NAND2_X1 U14319 ( .A1(n11407), .A2(n11406), .ZN(n11408) );
  NAND2_X1 U14320 ( .A1(n11408), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n16736) );
  AOI22_X1 U14321 ( .A1(n11500), .A2(n11423), .B1(n11529), .B2(
        P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11410) );
  OR2_X1 U14322 ( .A1(n12143), .A2(n11412), .ZN(n11417) );
  NAND2_X1 U14323 ( .A1(n11414), .A2(n11413), .ZN(n11421) );
  XNOR2_X1 U14324 ( .A(n11423), .B(n11421), .ZN(n11415) );
  NAND2_X1 U14325 ( .A1(n16495), .A2(n11415), .ZN(n11416) );
  NAND2_X1 U14326 ( .A1(n11417), .A2(n11416), .ZN(n11418) );
  INV_X1 U14327 ( .A(n11418), .ZN(n11420) );
  INV_X1 U14328 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n11419) );
  NAND2_X1 U14329 ( .A1(n11420), .A2(n11419), .ZN(n16729) );
  INV_X1 U14330 ( .A(n11421), .ZN(n11422) );
  NAND2_X1 U14331 ( .A1(n11423), .A2(n11422), .ZN(n11424) );
  NOR2_X1 U14332 ( .A1(n13649), .A2(n11424), .ZN(n11425) );
  NOR2_X1 U14333 ( .A1(n16673), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n16707) );
  AND2_X1 U14334 ( .A1(n11429), .A2(n11520), .ZN(n11441) );
  AOI22_X1 U14335 ( .A1(n12603), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n11217), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11433) );
  AOI22_X1 U14336 ( .A1(n12607), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11278), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11432) );
  AOI22_X1 U14337 ( .A1(n9715), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n9762), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11431) );
  AOI22_X1 U14338 ( .A1(n12413), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n12539), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11430) );
  NAND4_X1 U14339 ( .A1(n11433), .A2(n11432), .A3(n11431), .A4(n11430), .ZN(
        n11439) );
  AOI22_X1 U14340 ( .A1(n12605), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12613), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11437) );
  AOI22_X1 U14341 ( .A1(n12604), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n9764), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11436) );
  AOI22_X1 U14342 ( .A1(n12614), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n12606), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11435) );
  AOI22_X1 U14343 ( .A1(n9760), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11163), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11434) );
  NAND4_X1 U14344 ( .A1(n11437), .A2(n11436), .A3(n11435), .A4(n11434), .ZN(
        n11438) );
  NOR2_X1 U14345 ( .A1(n11439), .A2(n11438), .ZN(n11440) );
  OR2_X1 U14346 ( .A1(n11441), .A2(n11440), .ZN(n11443) );
  NAND2_X1 U14347 ( .A1(n11443), .A2(n11442), .ZN(n12236) );
  NAND2_X1 U14348 ( .A1(n11444), .A2(n12236), .ZN(n11452) );
  INV_X1 U14349 ( .A(n11452), .ZN(n15676) );
  OAI22_X1 U14350 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n15676), .B1(
        n16673), .B2(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15778) );
  OAI21_X1 U14351 ( .B1(n16673), .B2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n15666), .ZN(n16709) );
  NOR3_X1 U14352 ( .A1(n16707), .A2(n15778), .A3(n16709), .ZN(n15665) );
  OR2_X1 U14353 ( .A1(n16673), .A2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11445) );
  NAND2_X1 U14354 ( .A1(n15665), .A2(n11445), .ZN(n15757) );
  INV_X1 U14355 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16796) );
  INV_X1 U14356 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n15763) );
  NAND2_X1 U14357 ( .A1(n16796), .A2(n15763), .ZN(n11446) );
  NAND2_X1 U14358 ( .A1(n16673), .A2(n11446), .ZN(n15759) );
  NAND2_X1 U14359 ( .A1(n16673), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n11447) );
  NAND2_X1 U14360 ( .A1(n15757), .A2(n11455), .ZN(n11449) );
  INV_X1 U14361 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n16785) );
  XNOR2_X1 U14362 ( .A(n16673), .B(n16785), .ZN(n16692) );
  OR2_X1 U14363 ( .A1(n16673), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n11448) );
  NAND2_X1 U14364 ( .A1(n11449), .A2(n16689), .ZN(n15746) );
  NOR2_X1 U14365 ( .A1(n16673), .A2(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n11450) );
  NAND2_X1 U14366 ( .A1(n16673), .A2(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n11454) );
  INV_X1 U14367 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n11451) );
  OR2_X1 U14368 ( .A1(n11452), .A2(n11451), .ZN(n11453) );
  NAND2_X1 U14369 ( .A1(n11454), .A2(n11453), .ZN(n15776) );
  AND2_X1 U14370 ( .A1(n16673), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n15779) );
  OAI21_X1 U14371 ( .B1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A(n16673), .ZN(n11456) );
  NAND2_X1 U14372 ( .A1(n16673), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n16671) );
  OR2_X1 U14373 ( .A1(n16673), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n11459) );
  AND2_X1 U14374 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15726) );
  INV_X1 U14375 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n11655) );
  INV_X1 U14376 ( .A(n15660), .ZN(n11461) );
  INV_X1 U14377 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n11460) );
  INV_X1 U14378 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n16674) );
  INV_X1 U14379 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15716) );
  NAND2_X2 U14380 ( .A1(n11463), .A2(n15637), .ZN(n15627) );
  INV_X1 U14381 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n11661) );
  NAND3_X1 U14382 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n12115) );
  INV_X1 U14383 ( .A(n12115), .ZN(n11465) );
  NAND2_X1 U14384 ( .A1(n16645), .A2(n11465), .ZN(n11464) );
  OAI21_X1 U14385 ( .B1(n16673), .B2(n11465), .A(n15627), .ZN(n13020) );
  NOR2_X1 U14386 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n12119) );
  INV_X1 U14387 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n12114) );
  NAND3_X1 U14388 ( .A1(n12119), .A2(n9980), .A3(n12114), .ZN(n11466) );
  AOI22_X1 U14389 ( .A1(n13020), .A2(n11466), .B1(n16645), .B2(n12114), .ZN(
        n13021) );
  XNOR2_X1 U14390 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n11482) );
  NAND2_X1 U14391 ( .A1(n11501), .A2(n11482), .ZN(n11469) );
  NAND2_X1 U14392 ( .A1(n21009), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11468) );
  NAND2_X1 U14393 ( .A1(n11469), .A2(n11468), .ZN(n11481) );
  NOR2_X1 U14394 ( .A1(n13316), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n11470) );
  OAI22_X1 U14395 ( .A1(n11481), .A2(n11470), .B1(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B2(n20941), .ZN(n11478) );
  NOR2_X1 U14396 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n21010), .ZN(
        n11471) );
  OR2_X1 U14397 ( .A1(n11478), .A2(n11471), .ZN(n11473) );
  NAND2_X1 U14398 ( .A1(n21010), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11472) );
  NAND2_X1 U14399 ( .A1(n11473), .A2(n11472), .ZN(n11477) );
  INV_X1 U14400 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n13297) );
  NOR2_X1 U14401 ( .A1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n13297), .ZN(
        n11474) );
  OR2_X1 U14402 ( .A1(n11477), .A2(n11474), .ZN(n11475) );
  INV_X1 U14403 ( .A(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n20939) );
  OR2_X1 U14404 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n20939), .ZN(
        n11476) );
  INV_X1 U14405 ( .A(n11495), .ZN(n11484) );
  NOR2_X1 U14406 ( .A1(n11477), .A2(n11476), .ZN(n11527) );
  XNOR2_X1 U14407 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n21010), .ZN(
        n11479) );
  XNOR2_X1 U14408 ( .A(n11479), .B(n11478), .ZN(n11523) );
  XNOR2_X1 U14409 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n11480) );
  XNOR2_X1 U14410 ( .A(n11481), .B(n11480), .ZN(n11499) );
  XNOR2_X1 U14411 ( .A(n11501), .B(n11482), .ZN(n11513) );
  OR4_X1 U14412 ( .A1(n11527), .A2(n11523), .A3(n11499), .A4(n11513), .ZN(
        n11483) );
  NAND2_X1 U14413 ( .A1(n11484), .A2(n11483), .ZN(n13281) );
  INV_X1 U14414 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n11485) );
  NAND2_X1 U14415 ( .A1(n11486), .A2(n11485), .ZN(n16516) );
  INV_X1 U14416 ( .A(n16516), .ZN(n13273) );
  NAND2_X1 U14417 ( .A1(READY1), .A2(READY11_REG_SCAN_IN), .ZN(n21287) );
  OAI211_X1 U14418 ( .C1(n13951), .C2(n13273), .A(n21287), .B(n11487), .ZN(
        n11536) );
  INV_X1 U14419 ( .A(n13227), .ZN(n11493) );
  NAND2_X1 U14420 ( .A1(n15821), .A2(n13936), .ZN(n11489) );
  NAND3_X1 U14421 ( .A1(n11561), .A2(n11545), .A3(n11489), .ZN(n11544) );
  INV_X1 U14422 ( .A(n11544), .ZN(n11491) );
  OAI211_X1 U14423 ( .C1(n13951), .C2(n13393), .A(n11490), .B(n11192), .ZN(
        n11559) );
  NAND2_X1 U14424 ( .A1(n11491), .A2(n11559), .ZN(n11492) );
  NAND2_X1 U14425 ( .A1(n11493), .A2(n11492), .ZN(n13286) );
  NAND2_X1 U14426 ( .A1(n11495), .A2(n11500), .ZN(n11534) );
  INV_X1 U14427 ( .A(n11499), .ZN(n11496) );
  NAND2_X1 U14428 ( .A1(n13875), .A2(n11192), .ZN(n11497) );
  NAND2_X1 U14429 ( .A1(n11497), .A2(n13951), .ZN(n11517) );
  INV_X1 U14430 ( .A(n11517), .ZN(n11498) );
  AOI211_X1 U14431 ( .C1(n11529), .C2(n11499), .A(n11516), .B(n11498), .ZN(
        n11519) );
  INV_X1 U14432 ( .A(n11501), .ZN(n11502) );
  OAI21_X1 U14433 ( .B1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n21110), .A(
        n11502), .ZN(n11503) );
  NOR2_X1 U14434 ( .A1(n11510), .A2(n11503), .ZN(n11506) );
  INV_X1 U14435 ( .A(n11503), .ZN(n11504) );
  OAI211_X1 U14436 ( .C1(n13936), .C2(n11553), .A(n11504), .B(n11517), .ZN(
        n11505) );
  INV_X1 U14437 ( .A(n11511), .ZN(n11515) );
  NAND2_X1 U14438 ( .A1(n13875), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11508) );
  OAI21_X1 U14439 ( .B1(n13951), .B2(n11510), .A(n11508), .ZN(n11507) );
  INV_X1 U14440 ( .A(n11512), .ZN(n11514) );
  AND2_X1 U14441 ( .A1(n11508), .A2(n11177), .ZN(n11509) );
  NAND2_X1 U14442 ( .A1(n11510), .A2(n11509), .ZN(n11526) );
  INV_X1 U14443 ( .A(n11516), .ZN(n11518) );
  NAND2_X1 U14444 ( .A1(n11523), .A2(n11520), .ZN(n11521) );
  AOI22_X1 U14445 ( .A1(n11524), .A2(n11523), .B1(n11522), .B2(n11521), .ZN(
        n11532) );
  INV_X1 U14446 ( .A(n11527), .ZN(n11525) );
  NOR2_X1 U14447 ( .A1(n11529), .A2(n11525), .ZN(n11531) );
  INV_X1 U14448 ( .A(n11526), .ZN(n11528) );
  NAND3_X1 U14449 ( .A1(n11529), .A2(n11528), .A3(n11527), .ZN(n11530) );
  OAI21_X1 U14450 ( .B1(n11532), .B2(n11531), .A(n11530), .ZN(n11533) );
  INV_X1 U14451 ( .A(n15821), .ZN(n12320) );
  OAI211_X1 U14452 ( .C1(n13281), .C2(n11536), .A(n13286), .B(n11535), .ZN(
        n11538) );
  NAND2_X1 U14453 ( .A1(n11537), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n20767) );
  INV_X1 U14454 ( .A(n20767), .ZN(n13289) );
  NAND2_X1 U14455 ( .A1(n11538), .A2(n13289), .ZN(n11543) );
  NAND2_X1 U14456 ( .A1(n13951), .A2(n16516), .ZN(n13939) );
  AND2_X1 U14457 ( .A1(n13939), .A2(n21287), .ZN(n11540) );
  NAND2_X1 U14458 ( .A1(n11539), .A2(n11540), .ZN(n16496) );
  NAND3_X1 U14459 ( .A1(n16496), .A2(n11192), .A3(n11179), .ZN(n11541) );
  NAND3_X1 U14460 ( .A1(n13527), .A2(n11541), .A3(n13880), .ZN(n11542) );
  NOR2_X1 U14461 ( .A1(n11544), .A2(n11553), .ZN(n16486) );
  NAND2_X1 U14462 ( .A1(n11545), .A2(n11194), .ZN(n11546) );
  NOR2_X1 U14463 ( .A1(n11546), .A2(n15821), .ZN(n13304) );
  NOR2_X1 U14464 ( .A1(n16486), .A2(n13304), .ZN(n13225) );
  OAI22_X1 U14465 ( .A1(n11547), .A2(n13951), .B1(n11129), .B2(n11548), .ZN(
        n11549) );
  INV_X1 U14466 ( .A(n11549), .ZN(n11551) );
  NAND3_X1 U14467 ( .A1(n13225), .A2(n11551), .A3(n11550), .ZN(n11552) );
  INV_X1 U14468 ( .A(n11553), .ZN(n11557) );
  OR2_X1 U14469 ( .A1(n13951), .A2(n11192), .ZN(n13283) );
  NAND2_X1 U14470 ( .A1(n11178), .A2(n11192), .ZN(n11601) );
  NAND2_X1 U14471 ( .A1(n14818), .A2(n11567), .ZN(n11556) );
  OAI211_X1 U14472 ( .C1(n11557), .C2(n13283), .A(n11556), .B(n11555), .ZN(
        n11558) );
  INV_X1 U14473 ( .A(n11558), .ZN(n11560) );
  OAI211_X1 U14474 ( .C1(n11561), .C2(n12132), .A(n11560), .B(n11559), .ZN(
        n11562) );
  INV_X1 U14475 ( .A(n11562), .ZN(n11564) );
  AND2_X1 U14476 ( .A1(n11564), .A2(n11563), .ZN(n13301) );
  NAND2_X1 U14477 ( .A1(n13301), .A2(n11565), .ZN(n11566) );
  NAND2_X1 U14478 ( .A1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15700) );
  OR2_X1 U14479 ( .A1(n14817), .A2(n11567), .ZN(n11568) );
  NOR2_X1 U14480 ( .A1(n11568), .A2(n15821), .ZN(n13303) );
  NAND2_X1 U14481 ( .A1(n13227), .A2(n11177), .ZN(n14744) );
  OAI21_X1 U14482 ( .B1(n15733), .B2(n20932), .A(n12115), .ZN(n11569) );
  INV_X1 U14483 ( .A(n11569), .ZN(n11575) );
  INV_X1 U14484 ( .A(n15733), .ZN(n20929) );
  NAND2_X1 U14485 ( .A1(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n16763) );
  INV_X1 U14486 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15765) );
  INV_X1 U14487 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15752) );
  NOR4_X1 U14488 ( .A1(n15765), .A2(n15763), .A3(n16785), .A4(n15752), .ZN(
        n15737) );
  NAND2_X1 U14489 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n15737), .ZN(
        n11574) );
  INV_X1 U14490 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16806) );
  INV_X1 U14491 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n14357) );
  INV_X1 U14492 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n16828) );
  NOR3_X1 U14493 ( .A1(n14357), .A2(n11419), .A3(n16828), .ZN(n15802) );
  NAND3_X1 U14494 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A3(n15802), .ZN(n16801) );
  NOR2_X1 U14495 ( .A1(n16806), .A2(n16801), .ZN(n15786) );
  NAND2_X1 U14496 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n15786), .ZN(
        n11570) );
  NAND2_X1 U14497 ( .A1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n13848) );
  INV_X1 U14498 ( .A(n13848), .ZN(n13847) );
  INV_X1 U14499 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n20930) );
  INV_X1 U14500 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n13460) );
  OAI21_X1 U14501 ( .B1(n20930), .B2(n13460), .A(n11590), .ZN(n13555) );
  NAND3_X1 U14502 ( .A1(n13847), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A3(
        n13555), .ZN(n15799) );
  NOR2_X1 U14503 ( .A1(n11570), .A2(n15799), .ZN(n11577) );
  NAND2_X1 U14504 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n11577), .ZN(
        n15769) );
  NAND4_X1 U14505 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A4(n13847), .ZN(n15789) );
  NOR2_X1 U14506 ( .A1(n15789), .A2(n11570), .ZN(n11579) );
  AND2_X1 U14507 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n11579), .ZN(
        n15735) );
  INV_X1 U14508 ( .A(n11574), .ZN(n11580) );
  NAND2_X1 U14509 ( .A1(n20934), .A2(n20930), .ZN(n11572) );
  INV_X2 U14510 ( .A(n16823), .ZN(n16782) );
  OR2_X1 U14511 ( .A1(n11679), .A2(n16782), .ZN(n11571) );
  OAI221_X1 U14512 ( .B1(n15736), .B2(n15735), .C1(n15736), .C2(n11580), .A(
        n15784), .ZN(n11573) );
  AOI221_X1 U14513 ( .B1(n11574), .B2(n15733), .C1(n15769), .C2(n15733), .A(
        n11573), .ZN(n15725) );
  INV_X1 U14514 ( .A(n15784), .ZN(n15732) );
  AOI21_X1 U14515 ( .B1(n15726), .B2(n15725), .A(n15800), .ZN(n16759) );
  OAI21_X1 U14516 ( .B1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n20929), .A(
        n16751), .ZN(n15708) );
  AOI211_X1 U14517 ( .C1(n20934), .C2(n15700), .A(n11575), .B(n15708), .ZN(
        n16750) );
  NAND2_X1 U14518 ( .A1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n16750), .ZN(
        n15701) );
  INV_X1 U14519 ( .A(n15701), .ZN(n11576) );
  AND2_X1 U14520 ( .A1(n16750), .A2(n15738), .ZN(n12134) );
  AOI21_X1 U14521 ( .B1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n11576), .A(
        n12134), .ZN(n15696) );
  NOR2_X1 U14522 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n20932), .ZN(
        n13450) );
  AND2_X1 U14523 ( .A1(n15733), .A2(n11577), .ZN(n11578) );
  AOI21_X1 U14524 ( .B1(n15783), .B2(n11579), .A(n11578), .ZN(n16787) );
  NOR2_X1 U14525 ( .A1(n16787), .A2(n16796), .ZN(n15741) );
  NAND2_X1 U14526 ( .A1(n11580), .A2(n15741), .ZN(n16774) );
  INV_X1 U14527 ( .A(n15726), .ZN(n11581) );
  NAND3_X1 U14528 ( .A1(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(n16764), .ZN(n16758) );
  NOR2_X1 U14529 ( .A1(n12115), .A2(n16758), .ZN(n15702) );
  NAND2_X1 U14530 ( .A1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n15702), .ZN(
        n15689) );
  INV_X1 U14531 ( .A(n15689), .ZN(n12135) );
  INV_X1 U14532 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15691) );
  INV_X1 U14533 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n21245) );
  NOR2_X1 U14534 ( .A1(n16823), .A2(n21245), .ZN(n11582) );
  AOI221_X1 U14535 ( .B1(n15696), .B2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), 
        .C1(n12135), .C2(n15691), .A(n11582), .ZN(n11682) );
  NAND2_X1 U14536 ( .A1(n11601), .A2(n13460), .ZN(n11584) );
  NAND2_X1 U14537 ( .A1(n13275), .A2(n10124), .ZN(n11583) );
  NAND3_X1 U14538 ( .A1(n11584), .A2(n12132), .A3(n11583), .ZN(n11585) );
  NAND2_X1 U14539 ( .A1(n11601), .A2(P1_EBX_REG_0__SCAN_IN), .ZN(n11587) );
  INV_X1 U14540 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n15459) );
  NAND2_X1 U14541 ( .A1(n12132), .A2(n15459), .ZN(n11586) );
  NAND2_X1 U14542 ( .A1(n11587), .A2(n11586), .ZN(n13342) );
  XNOR2_X1 U14543 ( .A(n11588), .B(n13342), .ZN(n13406) );
  NAND2_X1 U14544 ( .A1(n13406), .A2(n13275), .ZN(n13408) );
  NAND2_X1 U14545 ( .A1(n13408), .A2(n11588), .ZN(n13458) );
  NAND2_X1 U14546 ( .A1(n11601), .A2(n11590), .ZN(n11593) );
  INV_X1 U14547 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n11591) );
  NAND2_X1 U14548 ( .A1(n13275), .A2(n11591), .ZN(n11592) );
  NAND3_X1 U14549 ( .A1(n11593), .A2(n12132), .A3(n11592), .ZN(n11594) );
  MUX2_X1 U14550 ( .A(n11673), .B(n12132), .S(P1_EBX_REG_3__SCAN_IN), .Z(
        n11598) );
  OAI21_X1 U14551 ( .B1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n14818), .A(
        n11598), .ZN(n13559) );
  INV_X1 U14552 ( .A(n11601), .ZN(n11599) );
  NAND2_X1 U14553 ( .A1(n11599), .A2(n14817), .ZN(n11649) );
  NAND2_X1 U14554 ( .A1(n14817), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11600) );
  AND2_X1 U14555 ( .A1(n11649), .A2(n11600), .ZN(n11603) );
  MUX2_X1 U14556 ( .A(n11589), .B(n11601), .S(P1_EBX_REG_4__SCAN_IN), .Z(
        n11602) );
  NAND2_X1 U14557 ( .A1(n11603), .A2(n11602), .ZN(n13724) );
  INV_X1 U14558 ( .A(P1_EBX_REG_5__SCAN_IN), .ZN(n13825) );
  NAND2_X1 U14559 ( .A1(n13275), .A2(n13825), .ZN(n11605) );
  NAND2_X1 U14560 ( .A1(n12132), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11604) );
  NAND3_X1 U14561 ( .A1(n11601), .A2(n11605), .A3(n11604), .ZN(n11606) );
  OAI21_X1 U14562 ( .B1(n11673), .B2(P1_EBX_REG_5__SCAN_IN), .A(n11606), .ZN(
        n13824) );
  MUX2_X1 U14563 ( .A(n11589), .B(n11601), .S(P1_EBX_REG_6__SCAN_IN), .Z(
        n11610) );
  NAND2_X1 U14564 ( .A1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n14817), .ZN(
        n11609) );
  INV_X1 U14565 ( .A(n11673), .ZN(n11611) );
  INV_X1 U14566 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n14085) );
  NAND2_X1 U14567 ( .A1(n11611), .A2(n14085), .ZN(n11615) );
  NAND2_X1 U14568 ( .A1(n13275), .A2(n14085), .ZN(n11613) );
  NAND2_X1 U14569 ( .A1(n12132), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11612) );
  NAND3_X1 U14570 ( .A1(n11601), .A2(n11613), .A3(n11612), .ZN(n11614) );
  NAND2_X1 U14571 ( .A1(n14817), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11616) );
  AND2_X1 U14572 ( .A1(n11649), .A2(n11616), .ZN(n11618) );
  MUX2_X1 U14573 ( .A(n11589), .B(n11601), .S(P1_EBX_REG_8__SCAN_IN), .Z(
        n11617) );
  NAND2_X1 U14574 ( .A1(n11618), .A2(n11617), .ZN(n14118) );
  INV_X1 U14575 ( .A(P1_EBX_REG_9__SCAN_IN), .ZN(n11619) );
  NAND2_X1 U14576 ( .A1(n13275), .A2(n11619), .ZN(n11621) );
  NAND2_X1 U14577 ( .A1(n12132), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11620) );
  NAND3_X1 U14578 ( .A1(n11601), .A2(n11621), .A3(n11620), .ZN(n11622) );
  OAI21_X1 U14579 ( .B1(n11673), .B2(P1_EBX_REG_9__SCAN_IN), .A(n11622), .ZN(
        n13992) );
  MUX2_X1 U14580 ( .A(n11589), .B(n11601), .S(P1_EBX_REG_10__SCAN_IN), .Z(
        n11624) );
  NAND2_X1 U14581 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n14817), .ZN(
        n11623) );
  AND3_X1 U14582 ( .A1(n11624), .A2(n11649), .A3(n11623), .ZN(n14292) );
  MUX2_X1 U14583 ( .A(n11673), .B(n12132), .S(P1_EBX_REG_11__SCAN_IN), .Z(
        n11626) );
  OR2_X1 U14584 ( .A1(n14818), .A2(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n11625) );
  AND2_X1 U14585 ( .A1(n11626), .A2(n11625), .ZN(n14575) );
  NAND2_X1 U14586 ( .A1(n14817), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n11627) );
  AND2_X1 U14587 ( .A1(n11649), .A2(n11627), .ZN(n11629) );
  MUX2_X1 U14588 ( .A(n11589), .B(n11601), .S(P1_EBX_REG_12__SCAN_IN), .Z(
        n11628) );
  NAND2_X1 U14589 ( .A1(n11629), .A2(n11628), .ZN(n14674) );
  MUX2_X1 U14590 ( .A(n11673), .B(n12132), .S(P1_EBX_REG_13__SCAN_IN), .Z(
        n11630) );
  OAI21_X1 U14591 ( .B1(n14818), .B2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n11630), .ZN(n14683) );
  OR2_X1 U14592 ( .A1(n11589), .A2(P1_EBX_REG_14__SCAN_IN), .ZN(n11634) );
  NAND2_X1 U14593 ( .A1(n11601), .A2(n15763), .ZN(n11632) );
  INV_X1 U14594 ( .A(P1_EBX_REG_14__SCAN_IN), .ZN(n15542) );
  NAND2_X1 U14595 ( .A1(n13275), .A2(n15542), .ZN(n11631) );
  NAND3_X1 U14596 ( .A1(n11632), .A2(n12132), .A3(n11631), .ZN(n11633) );
  AND2_X1 U14597 ( .A1(n11634), .A2(n11633), .ZN(n15444) );
  MUX2_X1 U14598 ( .A(n11673), .B(n12132), .S(P1_EBX_REG_15__SCAN_IN), .Z(
        n11635) );
  OAI21_X1 U14599 ( .B1(n14818), .B2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n11635), .ZN(n15537) );
  OR2_X1 U14600 ( .A1(n11589), .A2(P1_EBX_REG_16__SCAN_IN), .ZN(n11639) );
  NAND2_X1 U14601 ( .A1(n11601), .A2(n16785), .ZN(n11637) );
  INV_X1 U14602 ( .A(P1_EBX_REG_16__SCAN_IN), .ZN(n16600) );
  NAND2_X1 U14603 ( .A1(n13275), .A2(n16600), .ZN(n11636) );
  NAND3_X1 U14604 ( .A1(n11637), .A2(n12132), .A3(n11636), .ZN(n11638) );
  NAND2_X1 U14605 ( .A1(n11639), .A2(n11638), .ZN(n15531) );
  MUX2_X1 U14606 ( .A(n11673), .B(n12132), .S(P1_EBX_REG_17__SCAN_IN), .Z(
        n11640) );
  OAI21_X1 U14607 ( .B1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n14818), .A(
        n11640), .ZN(n15432) );
  OR2_X1 U14608 ( .A1(n11589), .A2(P1_EBX_REG_18__SCAN_IN), .ZN(n11645) );
  INV_X1 U14609 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n11641) );
  NAND2_X1 U14610 ( .A1(n11601), .A2(n11641), .ZN(n11643) );
  INV_X1 U14611 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n15524) );
  NAND2_X1 U14612 ( .A1(n13275), .A2(n15524), .ZN(n11642) );
  NAND3_X1 U14613 ( .A1(n11643), .A2(n12132), .A3(n11642), .ZN(n11644) );
  AND2_X1 U14614 ( .A1(n11645), .A2(n11644), .ZN(n15521) );
  MUX2_X1 U14615 ( .A(n11673), .B(n12132), .S(P1_EBX_REG_19__SCAN_IN), .Z(
        n11647) );
  OR2_X1 U14616 ( .A1(n14818), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n11646) );
  AND2_X1 U14617 ( .A1(n11647), .A2(n11646), .ZN(n16578) );
  NAND2_X1 U14618 ( .A1(n14817), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n11648) );
  AND2_X1 U14619 ( .A1(n11649), .A2(n11648), .ZN(n11651) );
  MUX2_X1 U14620 ( .A(n11589), .B(n11601), .S(P1_EBX_REG_20__SCAN_IN), .Z(
        n11650) );
  NAND2_X1 U14621 ( .A1(n11651), .A2(n11650), .ZN(n15515) );
  MUX2_X1 U14622 ( .A(n11673), .B(n12132), .S(P1_EBX_REG_21__SCAN_IN), .Z(
        n11652) );
  OAI21_X1 U14623 ( .B1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n14818), .A(
        n11652), .ZN(n15504) );
  MUX2_X1 U14624 ( .A(n11673), .B(n12132), .S(P1_EBX_REG_23__SCAN_IN), .Z(
        n11654) );
  OR2_X1 U14625 ( .A1(n14818), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n11653) );
  AND2_X1 U14626 ( .A1(n11654), .A2(n11653), .ZN(n15494) );
  OR2_X1 U14627 ( .A1(n11589), .A2(P1_EBX_REG_22__SCAN_IN), .ZN(n11660) );
  NAND2_X1 U14628 ( .A1(n11601), .A2(n11655), .ZN(n11658) );
  INV_X1 U14629 ( .A(P1_EBX_REG_22__SCAN_IN), .ZN(n11656) );
  NAND2_X1 U14630 ( .A1(n13275), .A2(n11656), .ZN(n11657) );
  NAND3_X1 U14631 ( .A1(n11658), .A2(n12132), .A3(n11657), .ZN(n11659) );
  NAND2_X1 U14632 ( .A1(n11660), .A2(n11659), .ZN(n15502) );
  OR2_X1 U14633 ( .A1(n11589), .A2(P1_EBX_REG_24__SCAN_IN), .ZN(n11665) );
  NAND2_X1 U14634 ( .A1(n11601), .A2(n11661), .ZN(n11663) );
  INV_X1 U14635 ( .A(P1_EBX_REG_24__SCAN_IN), .ZN(n15487) );
  NAND2_X1 U14636 ( .A1(n13275), .A2(n15487), .ZN(n11662) );
  NAND3_X1 U14637 ( .A1(n11663), .A2(n12132), .A3(n11662), .ZN(n11664) );
  NAND2_X1 U14638 ( .A1(n11665), .A2(n11664), .ZN(n15485) );
  MUX2_X1 U14639 ( .A(n11673), .B(n12132), .S(P1_EBX_REG_25__SCAN_IN), .Z(
        n11667) );
  OR2_X1 U14640 ( .A1(n14818), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n11666) );
  AND2_X1 U14641 ( .A1(n11667), .A2(n11666), .ZN(n15479) );
  OR2_X1 U14642 ( .A1(n11589), .A2(P1_EBX_REG_26__SCAN_IN), .ZN(n11672) );
  NAND2_X1 U14643 ( .A1(n11601), .A2(n12114), .ZN(n11670) );
  INV_X1 U14644 ( .A(P1_EBX_REG_26__SCAN_IN), .ZN(n11668) );
  NAND2_X1 U14645 ( .A1(n13275), .A2(n11668), .ZN(n11669) );
  NAND3_X1 U14646 ( .A1(n11670), .A2(n12132), .A3(n11669), .ZN(n11671) );
  AND2_X1 U14647 ( .A1(n11672), .A2(n11671), .ZN(n15183) );
  MUX2_X1 U14648 ( .A(n11673), .B(n12132), .S(P1_EBX_REG_27__SCAN_IN), .Z(
        n11674) );
  OAI21_X1 U14649 ( .B1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n14818), .A(
        n11674), .ZN(n11675) );
  AND2_X1 U14650 ( .A1(n15184), .A2(n11675), .ZN(n11676) );
  OR2_X1 U14651 ( .A1(n9788), .A2(n11676), .ZN(n15473) );
  INV_X1 U14652 ( .A(n15473), .ZN(n11680) );
  INV_X1 U14653 ( .A(n11547), .ZN(n13222) );
  NAND2_X1 U14654 ( .A1(n13222), .A2(n13951), .ZN(n13272) );
  OAI21_X1 U14655 ( .B1(n11548), .B2(n11677), .A(n13272), .ZN(n11678) );
  NAND2_X1 U14656 ( .A1(n11680), .A2(n16809), .ZN(n11681) );
  INV_X1 U14657 ( .A(n11686), .ZN(n11688) );
  NAND2_X1 U14658 ( .A1(n11688), .A2(n11687), .ZN(n11689) );
  XNOR2_X1 U14659 ( .A(n11685), .B(n11689), .ZN(n12036) );
  NAND2_X1 U14660 ( .A1(n20754), .A2(n20755), .ZN(n11691) );
  MUX2_X1 U14661 ( .A(n11691), .B(n11730), .S(n11690), .Z(n11701) );
  INV_X1 U14662 ( .A(n11730), .ZN(n12093) );
  OAI21_X1 U14663 ( .B1(n11694), .B2(n11693), .A(n12093), .ZN(n11698) );
  OAI211_X1 U14664 ( .C1(n20755), .C2(n11696), .A(n13592), .B(n11695), .ZN(
        n11697) );
  OAI211_X1 U14665 ( .C1(n11692), .C2(n11699), .A(n11698), .B(n11697), .ZN(
        n11700) );
  NAND2_X1 U14666 ( .A1(n11701), .A2(n11700), .ZN(n11703) );
  MUX2_X1 U14667 ( .A(n11703), .B(n11730), .S(n11702), .Z(n11704) );
  NAND2_X1 U14668 ( .A1(n11704), .A2(n11706), .ZN(n11705) );
  MUX2_X1 U14669 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B(n11705), .S(
        P2_STATE2_REG_0__SCAN_IN), .Z(n11709) );
  INV_X1 U14670 ( .A(n11706), .ZN(n11707) );
  NAND2_X1 U14671 ( .A1(n11707), .A2(n13119), .ZN(n11708) );
  NAND2_X1 U14672 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n20625), .ZN(n20762) );
  INV_X2 U14673 ( .A(n20762), .ZN(n20765) );
  INV_X1 U14674 ( .A(P2_STATE_REG_1__SCAN_IN), .ZN(n19720) );
  INV_X1 U14675 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n20636) );
  NAND2_X1 U14676 ( .A1(n19720), .A2(n20636), .ZN(n20630) );
  NAND2_X1 U14677 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n20748) );
  NAND2_X1 U14678 ( .A1(n20756), .A2(n20748), .ZN(n12095) );
  INV_X1 U14679 ( .A(n12095), .ZN(n13112) );
  NAND2_X1 U14680 ( .A1(n13132), .A2(n13112), .ZN(n13136) );
  OAI22_X1 U14681 ( .A1(n13132), .A2(n13592), .B1(n20755), .B2(n11709), .ZN(
        n11710) );
  NAND2_X1 U14682 ( .A1(n11710), .A2(n10335), .ZN(n11728) );
  NAND2_X1 U14683 ( .A1(n11711), .A2(n10325), .ZN(n11717) );
  NAND2_X1 U14684 ( .A1(n11713), .A2(n13368), .ZN(n11714) );
  NAND2_X1 U14685 ( .A1(n11714), .A2(n12096), .ZN(n11989) );
  NAND2_X1 U14686 ( .A1(n11989), .A2(n11715), .ZN(n11716) );
  AOI21_X1 U14687 ( .B1(n11717), .B2(n11712), .A(n11716), .ZN(n11987) );
  NAND2_X1 U14688 ( .A1(n9759), .A2(n10335), .ZN(n11985) );
  AOI21_X1 U14689 ( .B1(n11985), .B2(n13592), .A(n20121), .ZN(n11720) );
  NAND3_X1 U14690 ( .A1(n13796), .A2(n13734), .A3(n13112), .ZN(n11719) );
  OAI21_X1 U14691 ( .B1(n11720), .B2(n11718), .A(n11719), .ZN(n11721) );
  INV_X1 U14692 ( .A(n11721), .ZN(n11722) );
  AND2_X1 U14693 ( .A1(n11987), .A2(n11722), .ZN(n13133) );
  MUX2_X1 U14694 ( .A(n13796), .B(n11718), .S(n9759), .Z(n11723) );
  NAND3_X1 U14695 ( .A1(n11723), .A2(n13734), .A3(n20748), .ZN(n11724) );
  NAND2_X1 U14696 ( .A1(n13133), .A2(n11724), .ZN(n11725) );
  NOR2_X1 U14697 ( .A1(n11726), .A2(n11725), .ZN(n11727) );
  OAI211_X1 U14698 ( .C1(n10325), .C2(n13136), .A(n11728), .B(n11727), .ZN(
        n11729) );
  NOR2_X1 U14699 ( .A1(n13737), .A2(n11730), .ZN(n20735) );
  NAND2_X1 U14700 ( .A1(n12028), .A2(n20735), .ZN(n17071) );
  NAND2_X1 U14701 ( .A1(n11732), .A2(n9759), .ZN(n11733) );
  NAND2_X1 U14702 ( .A1(n13743), .A2(n11733), .ZN(n11734) );
  NAND2_X1 U14703 ( .A1(n12028), .A2(n11734), .ZN(n20062) );
  INV_X1 U14704 ( .A(n11735), .ZN(n11737) );
  NAND2_X1 U14705 ( .A1(n11737), .A2(n11736), .ZN(n13752) );
  NAND2_X1 U14706 ( .A1(n11738), .A2(n20755), .ZN(n11739) );
  NAND2_X1 U14707 ( .A1(n13752), .A2(n11739), .ZN(n11740) );
  NAND2_X1 U14708 ( .A1(n12028), .A2(n11740), .ZN(n17048) );
  NAND2_X1 U14709 ( .A1(n12037), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n11742) );
  INV_X2 U14710 ( .A(n10213), .ZN(n11977) );
  AOI22_X1 U14711 ( .A1(n11977), .A2(P2_EAX_REG_30__SCAN_IN), .B1(n9713), .B2(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n11741) );
  NAND2_X1 U14712 ( .A1(n11742), .A2(n11741), .ZN(n11980) );
  INV_X1 U14713 ( .A(n11980), .ZN(n11983) );
  NAND2_X1 U14714 ( .A1(n12037), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n11747) );
  INV_X1 U14715 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n11744) );
  NAND2_X1 U14716 ( .A1(n20755), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n11743) );
  OAI211_X1 U14717 ( .C1(n13368), .C2(n11744), .A(n11743), .B(n20333), .ZN(
        n11745) );
  INV_X1 U14718 ( .A(n11745), .ZN(n11746) );
  NAND2_X1 U14719 ( .A1(n11747), .A2(n11746), .ZN(n13371) );
  MUX2_X1 U14720 ( .A(n13368), .B(n20732), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n11749) );
  NAND2_X1 U14721 ( .A1(n13374), .A2(n11752), .ZN(n11763) );
  AND2_X1 U14722 ( .A1(n11749), .A2(n11763), .ZN(n11750) );
  AND2_X2 U14723 ( .A1(n13371), .A2(n13372), .ZN(n11760) );
  NAND2_X1 U14724 ( .A1(n12037), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n11754) );
  AOI22_X1 U14725 ( .A1(n11977), .A2(P2_EAX_REG_1__SCAN_IN), .B1(n9713), .B2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n11753) );
  NAND2_X1 U14726 ( .A1(n11754), .A2(n11753), .ZN(n11761) );
  INV_X1 U14727 ( .A(n11761), .ZN(n11755) );
  OR2_X1 U14728 ( .A1(n11756), .A2(n11953), .ZN(n11759) );
  NAND2_X1 U14729 ( .A1(n13369), .A2(n13368), .ZN(n11757) );
  INV_X1 U14730 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20721) );
  MUX2_X1 U14731 ( .A(n11757), .B(n20721), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n11758) );
  NAND2_X1 U14732 ( .A1(n13264), .A2(n13263), .ZN(n11767) );
  OR2_X1 U14733 ( .A1(n11953), .A2(n11762), .ZN(n11764) );
  OAI211_X1 U14734 ( .C1(n20333), .C2(n20710), .A(n11764), .B(n11763), .ZN(
        n11765) );
  AND3_X1 U14735 ( .A1(n11767), .A2(n11766), .A3(n11765), .ZN(n11768) );
  AOI21_X2 U14736 ( .B1(n11767), .B2(n11766), .A(n11765), .ZN(n11771) );
  NAND2_X1 U14737 ( .A1(n12037), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n11770) );
  AOI22_X1 U14738 ( .A1(n11977), .A2(P2_EAX_REG_2__SCAN_IN), .B1(n9713), .B2(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n11769) );
  NAND2_X1 U14739 ( .A1(n11770), .A2(n11769), .ZN(n13326) );
  NOR2_X1 U14740 ( .A1(n13327), .A2(n13326), .ZN(n13328) );
  NOR2_X2 U14741 ( .A1(n13328), .A2(n11771), .ZN(n13515) );
  NAND2_X1 U14742 ( .A1(n12037), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n11775) );
  AOI22_X1 U14743 ( .A1(n9713), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B1(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n11773) );
  NAND2_X1 U14744 ( .A1(n11977), .A2(P2_EAX_REG_3__SCAN_IN), .ZN(n11772) );
  AND2_X1 U14745 ( .A1(n11773), .A2(n11772), .ZN(n11774) );
  OAI211_X1 U14746 ( .C1(n11953), .C2(n11776), .A(n11775), .B(n11774), .ZN(
        n13514) );
  NAND2_X1 U14747 ( .A1(n13515), .A2(n13514), .ZN(n13701) );
  NAND2_X1 U14748 ( .A1(n12037), .A2(P2_REIP_REG_4__SCAN_IN), .ZN(n11780) );
  AOI22_X1 U14749 ( .A1(n11977), .A2(P2_EAX_REG_4__SCAN_IN), .B1(n9713), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n11779) );
  OR2_X1 U14750 ( .A1(n11953), .A2(n11777), .ZN(n11778) );
  INV_X1 U14751 ( .A(n11781), .ZN(n11783) );
  AOI22_X1 U14752 ( .A1(n12037), .A2(P2_REIP_REG_5__SCAN_IN), .B1(n11783), 
        .B2(n11782), .ZN(n11785) );
  AOI22_X1 U14753 ( .A1(n11977), .A2(P2_EAX_REG_5__SCAN_IN), .B1(n9713), .B2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n11784) );
  NAND2_X1 U14754 ( .A1(n11785), .A2(n11784), .ZN(n14266) );
  NAND2_X1 U14755 ( .A1(n13703), .A2(n14266), .ZN(n14265) );
  OR2_X1 U14756 ( .A1(n11953), .A2(n11786), .ZN(n11787) );
  NAND2_X1 U14757 ( .A1(n12037), .A2(P2_REIP_REG_6__SCAN_IN), .ZN(n11789) );
  AOI22_X1 U14758 ( .A1(n11977), .A2(P2_EAX_REG_6__SCAN_IN), .B1(n9713), .B2(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n11788) );
  INV_X1 U14759 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n20007) );
  OAI222_X1 U14760 ( .A1(n11791), .A2(n10936), .B1(n10213), .B2(n20007), .C1(
        n11972), .C2(n10940), .ZN(n13398) );
  NAND2_X1 U14761 ( .A1(n13399), .A2(n13398), .ZN(n13397) );
  NAND2_X1 U14762 ( .A1(n12037), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n11812) );
  AOI22_X1 U14763 ( .A1(n11977), .A2(P2_EAX_REG_8__SCAN_IN), .B1(n9713), .B2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n11811) );
  NAND2_X1 U14764 ( .A1(n10631), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n11795) );
  NAND2_X1 U14765 ( .A1(n14951), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n11794) );
  AOI22_X1 U14766 ( .A1(n10500), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n14885), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11793) );
  NAND2_X1 U14767 ( .A1(n10507), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n11792) );
  NAND4_X1 U14768 ( .A1(n11795), .A2(n11794), .A3(n11793), .A4(n11792), .ZN(
        n11801) );
  AOI22_X1 U14769 ( .A1(n10498), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n10499), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11799) );
  NAND2_X1 U14770 ( .A1(n14908), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n11798) );
  NAND2_X1 U14771 ( .A1(n14909), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n11797) );
  NAND2_X1 U14772 ( .A1(n14910), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n11796) );
  NAND4_X1 U14773 ( .A1(n11799), .A2(n11798), .A3(n11797), .A4(n11796), .ZN(
        n11800) );
  NOR2_X1 U14774 ( .A1(n11801), .A2(n11800), .ZN(n11809) );
  INV_X1 U14775 ( .A(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n14182) );
  OAI22_X1 U14776 ( .A1(n14919), .A2(n11802), .B1(n14917), .B2(n14182), .ZN(
        n11807) );
  INV_X1 U14777 ( .A(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11805) );
  AOI22_X1 U14778 ( .A1(n14967), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n11881), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11804) );
  NAND2_X1 U14779 ( .A1(n14450), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n11803) );
  OAI211_X1 U14780 ( .C1(n11805), .C2(n14473), .A(n11804), .B(n11803), .ZN(
        n11806) );
  NOR2_X1 U14781 ( .A1(n11807), .A2(n11806), .ZN(n11808) );
  AND2_X1 U14782 ( .A1(n11809), .A2(n11808), .ZN(n19962) );
  OR2_X1 U14783 ( .A1(n11953), .A2(n19962), .ZN(n11810) );
  NOR2_X2 U14784 ( .A1(n13397), .A2(n14200), .ZN(n13404) );
  NAND2_X1 U14785 ( .A1(n10631), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n11816) );
  NAND2_X1 U14786 ( .A1(n14951), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n11815) );
  AOI22_X1 U14787 ( .A1(n10500), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n14885), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11814) );
  NAND2_X1 U14788 ( .A1(n10507), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n11813) );
  NAND4_X1 U14789 ( .A1(n11816), .A2(n11815), .A3(n11814), .A4(n11813), .ZN(
        n11822) );
  AOI22_X1 U14790 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n10498), .B1(
        n10499), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11820) );
  NAND2_X1 U14791 ( .A1(n14908), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n11819) );
  NAND2_X1 U14792 ( .A1(n14909), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n11818) );
  NAND2_X1 U14793 ( .A1(n14910), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n11817) );
  NAND4_X1 U14794 ( .A1(n11820), .A2(n11819), .A3(n11818), .A4(n11817), .ZN(
        n11821) );
  NOR2_X1 U14795 ( .A1(n11822), .A2(n11821), .ZN(n11828) );
  INV_X1 U14796 ( .A(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n14159) );
  AOI22_X1 U14797 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n14967), .B1(
        n11881), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11824) );
  NAND2_X1 U14798 ( .A1(n14450), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n11823) );
  OAI211_X1 U14799 ( .C1(n14919), .C2(n14159), .A(n11824), .B(n11823), .ZN(
        n11826) );
  OAI22_X1 U14800 ( .A1(n14164), .A2(n14917), .B1(n14473), .B2(n14991), .ZN(
        n11825) );
  NOR2_X1 U14801 ( .A1(n11826), .A2(n11825), .ZN(n11827) );
  AND2_X1 U14802 ( .A1(n11828), .A2(n11827), .ZN(n19961) );
  NAND2_X1 U14803 ( .A1(n12037), .A2(P2_REIP_REG_9__SCAN_IN), .ZN(n11830) );
  AOI22_X1 U14804 ( .A1(n11977), .A2(P2_EAX_REG_9__SCAN_IN), .B1(n9713), .B2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n11829) );
  OAI211_X1 U14805 ( .C1(n11953), .C2(n19961), .A(n11830), .B(n11829), .ZN(
        n13405) );
  NAND2_X1 U14806 ( .A1(n13404), .A2(n13405), .ZN(n13402) );
  NAND2_X1 U14807 ( .A1(n12037), .A2(P2_REIP_REG_10__SCAN_IN), .ZN(n11850) );
  AOI22_X1 U14808 ( .A1(n11977), .A2(P2_EAX_REG_10__SCAN_IN), .B1(n9713), .B2(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n11849) );
  NAND2_X1 U14809 ( .A1(n10631), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n11834) );
  NAND2_X1 U14810 ( .A1(n14951), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(
        n11833) );
  AOI22_X1 U14811 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n10500), .B1(
        n14885), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11832) );
  NAND2_X1 U14812 ( .A1(n10507), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(
        n11831) );
  AND4_X1 U14813 ( .A1(n11834), .A2(n11833), .A3(n11832), .A4(n11831), .ZN(
        n11847) );
  AOI22_X1 U14814 ( .A1(n14957), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n14956), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11846) );
  INV_X1 U14815 ( .A(n14909), .ZN(n14961) );
  INV_X1 U14816 ( .A(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11837) );
  NAND2_X1 U14817 ( .A1(n10499), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n11836) );
  NAND2_X1 U14818 ( .A1(n10498), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(
        n11835) );
  OAI211_X1 U14819 ( .C1(n14961), .C2(n11837), .A(n11836), .B(n11835), .ZN(
        n11840) );
  INV_X1 U14820 ( .A(n14908), .ZN(n14964) );
  INV_X1 U14821 ( .A(n14910), .ZN(n14962) );
  INV_X1 U14822 ( .A(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n14142) );
  OAI22_X1 U14823 ( .A1(n14964), .A2(n11838), .B1(n14962), .B2(n14142), .ZN(
        n11839) );
  NOR2_X1 U14824 ( .A1(n11840), .A2(n11839), .ZN(n11845) );
  AOI22_X1 U14825 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n14967), .B1(
        n11881), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11842) );
  NAND2_X1 U14826 ( .A1(n14450), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n11841) );
  OAI211_X1 U14827 ( .C1(n14473), .C2(n14143), .A(n11842), .B(n11841), .ZN(
        n11843) );
  INV_X1 U14828 ( .A(n11843), .ZN(n11844) );
  NAND4_X1 U14829 ( .A1(n11847), .A2(n11846), .A3(n11845), .A4(n11844), .ZN(
        n13639) );
  INV_X1 U14830 ( .A(n13639), .ZN(n19952) );
  OR2_X1 U14831 ( .A1(n11953), .A2(n19952), .ZN(n11848) );
  NAND2_X1 U14832 ( .A1(n10631), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n11854) );
  NAND2_X1 U14833 ( .A1(n14951), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(
        n11853) );
  AOI22_X1 U14834 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n14450), .B1(
        n10499), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11852) );
  NAND2_X1 U14835 ( .A1(n10507), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n11851) );
  AND4_X1 U14836 ( .A1(n11854), .A2(n11853), .A3(n11852), .A4(n11851), .ZN(
        n11867) );
  AOI22_X1 U14837 ( .A1(n14957), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n14956), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11866) );
  NAND2_X1 U14838 ( .A1(n10498), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(
        n11856) );
  NAND2_X1 U14839 ( .A1(n10500), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n11855) );
  OAI211_X1 U14840 ( .C1(n14964), .C2(n11857), .A(n11856), .B(n11855), .ZN(
        n11860) );
  OAI22_X1 U14841 ( .A1(n14961), .A2(n11858), .B1(n14962), .B2(n14468), .ZN(
        n11859) );
  NOR2_X1 U14842 ( .A1(n11860), .A2(n11859), .ZN(n11865) );
  AOI22_X1 U14843 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n14967), .B1(
        n11881), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11862) );
  NAND2_X1 U14844 ( .A1(n14885), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(
        n11861) );
  OAI211_X1 U14845 ( .C1(n14473), .C2(n14469), .A(n11862), .B(n11861), .ZN(
        n11863) );
  INV_X1 U14846 ( .A(n11863), .ZN(n11864) );
  NAND4_X1 U14847 ( .A1(n11867), .A2(n11866), .A3(n11865), .A4(n11864), .ZN(
        n13638) );
  INV_X1 U14848 ( .A(n13638), .ZN(n19951) );
  NAND2_X1 U14849 ( .A1(n12037), .A2(P2_REIP_REG_11__SCAN_IN), .ZN(n11869) );
  AOI22_X1 U14850 ( .A1(n11977), .A2(P2_EAX_REG_11__SCAN_IN), .B1(n9713), .B2(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n11868) );
  OAI211_X1 U14851 ( .C1(n11953), .C2(n19951), .A(n11869), .B(n11868), .ZN(
        n13473) );
  NAND2_X1 U14852 ( .A1(n12037), .A2(P2_REIP_REG_12__SCAN_IN), .ZN(n11890) );
  AOI22_X1 U14853 ( .A1(n11977), .A2(P2_EAX_REG_12__SCAN_IN), .B1(n9713), .B2(
        P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n11889) );
  NAND2_X1 U14854 ( .A1(n10631), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n11873) );
  NAND2_X1 U14855 ( .A1(n14951), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n11872) );
  AOI22_X1 U14856 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n10500), .B1(
        n14885), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11871) );
  NAND2_X1 U14857 ( .A1(n10507), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n11870) );
  NAND4_X1 U14858 ( .A1(n11873), .A2(n11872), .A3(n11871), .A4(n11870), .ZN(
        n11879) );
  AOI22_X1 U14859 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n10498), .B1(
        n10499), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11877) );
  NAND2_X1 U14860 ( .A1(n14908), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n11876) );
  NAND2_X1 U14861 ( .A1(n14909), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n11875) );
  NAND2_X1 U14862 ( .A1(n14910), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n11874) );
  NAND4_X1 U14863 ( .A1(n11877), .A2(n11876), .A3(n11875), .A4(n11874), .ZN(
        n11878) );
  NOR2_X1 U14864 ( .A1(n11879), .A2(n11878), .ZN(n11887) );
  INV_X1 U14865 ( .A(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n14453) );
  OAI22_X1 U14866 ( .A1(n14919), .A2(n11880), .B1(n14917), .B2(n14453), .ZN(
        n11885) );
  AOI22_X1 U14867 ( .A1(n14967), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n11881), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11883) );
  NAND2_X1 U14868 ( .A1(n14450), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n11882) );
  OAI211_X1 U14869 ( .C1(n14473), .C2(n14449), .A(n11883), .B(n11882), .ZN(
        n11884) );
  NOR2_X1 U14870 ( .A1(n11885), .A2(n11884), .ZN(n11886) );
  AND2_X1 U14871 ( .A1(n11887), .A2(n11886), .ZN(n13711) );
  OR2_X1 U14872 ( .A1(n11953), .A2(n13711), .ZN(n11888) );
  AOI22_X1 U14873 ( .A1(n11977), .A2(P2_EAX_REG_13__SCAN_IN), .B1(n9713), .B2(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n11912) );
  INV_X1 U14874 ( .A(n11953), .ZN(n11910) );
  AOI22_X1 U14875 ( .A1(n14957), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n10631), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11909) );
  NAND2_X1 U14876 ( .A1(n14951), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n11894) );
  AOI22_X1 U14877 ( .A1(n14450), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n10499), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11893) );
  NAND2_X1 U14878 ( .A1(n14956), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n11892) );
  NAND2_X1 U14879 ( .A1(n10507), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n11891) );
  AND4_X1 U14880 ( .A1(n11894), .A2(n11893), .A3(n11892), .A4(n11891), .ZN(
        n11908) );
  AOI22_X1 U14881 ( .A1(n14967), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11881), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11896) );
  NAND2_X1 U14882 ( .A1(n14885), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n11895) );
  OAI211_X1 U14883 ( .C1(n11897), .C2(n14473), .A(n11896), .B(n11895), .ZN(
        n11898) );
  INV_X1 U14884 ( .A(n11898), .ZN(n11907) );
  NAND2_X1 U14885 ( .A1(n10498), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n11900) );
  NAND2_X1 U14886 ( .A1(n10500), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n11899) );
  OAI211_X1 U14887 ( .C1(n14964), .C2(n11901), .A(n11900), .B(n11899), .ZN(
        n11905) );
  OAI22_X1 U14888 ( .A1(n14961), .A2(n11903), .B1(n14962), .B2(n11902), .ZN(
        n11904) );
  NOR2_X1 U14889 ( .A1(n11905), .A2(n11904), .ZN(n11906) );
  NAND4_X1 U14890 ( .A1(n11909), .A2(n11908), .A3(n11907), .A4(n11906), .ZN(
        n13713) );
  NAND2_X1 U14891 ( .A1(n11910), .A2(n13713), .ZN(n11911) );
  OAI211_X1 U14892 ( .C1(n11972), .C2(n11913), .A(n11912), .B(n11911), .ZN(
        n13575) );
  NAND2_X1 U14893 ( .A1(n12037), .A2(P2_REIP_REG_14__SCAN_IN), .ZN(n11933) );
  AOI22_X1 U14894 ( .A1(n11977), .A2(P2_EAX_REG_14__SCAN_IN), .B1(n9713), .B2(
        P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n11932) );
  NAND2_X1 U14895 ( .A1(n10631), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n11917) );
  NAND2_X1 U14896 ( .A1(n14951), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n11916) );
  AOI22_X1 U14897 ( .A1(n10500), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n14885), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11915) );
  NAND2_X1 U14898 ( .A1(n10507), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n11914) );
  NAND4_X1 U14899 ( .A1(n11917), .A2(n11916), .A3(n11915), .A4(n11914), .ZN(
        n11923) );
  AOI22_X1 U14900 ( .A1(n10498), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n10499), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11921) );
  NAND2_X1 U14901 ( .A1(n14908), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n11920) );
  NAND2_X1 U14902 ( .A1(n14909), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n11919) );
  NAND2_X1 U14903 ( .A1(n14910), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n11918) );
  NAND4_X1 U14904 ( .A1(n11921), .A2(n11920), .A3(n11919), .A4(n11918), .ZN(
        n11922) );
  NOR2_X1 U14905 ( .A1(n11923), .A2(n11922), .ZN(n11930) );
  OAI22_X1 U14906 ( .A1(n14919), .A2(n11924), .B1(n14917), .B2(n14922), .ZN(
        n11928) );
  AOI22_X1 U14907 ( .A1(n14967), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n11881), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11926) );
  NAND2_X1 U14908 ( .A1(n14450), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n11925) );
  OAI211_X1 U14909 ( .C1(n14918), .C2(n14473), .A(n11926), .B(n11925), .ZN(
        n11927) );
  NOR2_X1 U14910 ( .A1(n11928), .A2(n11927), .ZN(n11929) );
  AND2_X1 U14911 ( .A1(n11930), .A2(n11929), .ZN(n19934) );
  OR2_X1 U14912 ( .A1(n11953), .A2(n19934), .ZN(n11931) );
  AND3_X1 U14913 ( .A1(n11933), .A2(n11932), .A3(n11931), .ZN(n16355) );
  NAND2_X1 U14914 ( .A1(n10631), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n11937) );
  NAND2_X1 U14915 ( .A1(n14951), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n11936) );
  AOI22_X1 U14916 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n10500), .B1(
        n14885), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11935) );
  NAND2_X1 U14917 ( .A1(n10507), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n11934) );
  NAND4_X1 U14918 ( .A1(n11937), .A2(n11936), .A3(n11935), .A4(n11934), .ZN(
        n11943) );
  AOI22_X1 U14919 ( .A1(n10498), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n10499), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11941) );
  NAND2_X1 U14920 ( .A1(n14908), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n11940) );
  NAND2_X1 U14921 ( .A1(n14909), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n11939) );
  NAND2_X1 U14922 ( .A1(n14910), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n11938) );
  NAND4_X1 U14923 ( .A1(n11941), .A2(n11940), .A3(n11939), .A4(n11938), .ZN(
        n11942) );
  NOR2_X1 U14924 ( .A1(n11943), .A2(n11942), .ZN(n11950) );
  INV_X1 U14925 ( .A(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n14970) );
  OAI22_X1 U14926 ( .A1(n14919), .A2(n14963), .B1(n14917), .B2(n14970), .ZN(
        n11948) );
  AOI22_X1 U14927 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n14967), .B1(
        n11881), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11945) );
  NAND2_X1 U14928 ( .A1(n14450), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n11944) );
  OAI211_X1 U14929 ( .C1(n14473), .C2(n11946), .A(n11945), .B(n11944), .ZN(
        n11947) );
  NOR2_X1 U14930 ( .A1(n11948), .A2(n11947), .ZN(n11949) );
  AND2_X1 U14931 ( .A1(n11950), .A2(n11949), .ZN(n19937) );
  NAND2_X1 U14932 ( .A1(n12037), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n11952) );
  AOI22_X1 U14933 ( .A1(n11977), .A2(P2_EAX_REG_15__SCAN_IN), .B1(n9713), .B2(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n11951) );
  OAI211_X1 U14934 ( .C1(n19937), .C2(n11953), .A(n11952), .B(n11951), .ZN(
        n13830) );
  AOI22_X1 U14935 ( .A1(n11977), .A2(P2_EAX_REG_16__SCAN_IN), .B1(n9713), .B2(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n11954) );
  OAI21_X1 U14936 ( .B1(n11972), .B2(n20654), .A(n11954), .ZN(n14303) );
  AOI22_X1 U14937 ( .A1(n11977), .A2(P2_EAX_REG_17__SCAN_IN), .B1(n9713), .B2(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n11955) );
  OAI21_X1 U14938 ( .B1(n11972), .B2(n20656), .A(n11955), .ZN(n14372) );
  AOI22_X1 U14939 ( .A1(n11977), .A2(P2_EAX_REG_18__SCAN_IN), .B1(n9713), .B2(
        P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n11956) );
  OAI21_X1 U14940 ( .B1(n11972), .B2(n20658), .A(n11956), .ZN(n14580) );
  AOI22_X1 U14941 ( .A1(n11977), .A2(P2_EAX_REG_19__SCAN_IN), .B1(n9713), .B2(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n11957) );
  OAI21_X1 U14942 ( .B1(n11972), .B2(n20660), .A(n11957), .ZN(n16022) );
  NAND2_X1 U14943 ( .A1(n12037), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n11959) );
  AOI22_X1 U14944 ( .A1(n11977), .A2(P2_EAX_REG_20__SCAN_IN), .B1(n9713), .B2(
        P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n11958) );
  AND2_X1 U14945 ( .A1(n11959), .A2(n11958), .ZN(n16008) );
  AOI22_X1 U14946 ( .A1(n11977), .A2(P2_EAX_REG_21__SCAN_IN), .B1(n9713), .B2(
        P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n11960) );
  OAI21_X1 U14947 ( .B1(n11972), .B2(n20663), .A(n11960), .ZN(n16001) );
  NAND2_X1 U14948 ( .A1(n16000), .A2(n16001), .ZN(n15988) );
  NAND2_X1 U14949 ( .A1(n12037), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n11962) );
  AOI22_X1 U14950 ( .A1(n11977), .A2(P2_EAX_REG_22__SCAN_IN), .B1(n9713), .B2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n11961) );
  AND2_X1 U14951 ( .A1(n11962), .A2(n11961), .ZN(n15989) );
  NAND2_X1 U14952 ( .A1(n12037), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n11965) );
  AOI22_X1 U14953 ( .A1(n11977), .A2(P2_EAX_REG_23__SCAN_IN), .B1(n9713), .B2(
        P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n11964) );
  AND2_X1 U14954 ( .A1(n11965), .A2(n11964), .ZN(n15976) );
  NAND2_X1 U14955 ( .A1(n12037), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n11968) );
  AOI22_X1 U14956 ( .A1(n11977), .A2(P2_EAX_REG_24__SCAN_IN), .B1(n9713), .B2(
        P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n11967) );
  AND2_X1 U14957 ( .A1(n11968), .A2(n11967), .ZN(n15859) );
  NOR2_X4 U14958 ( .A1(n15978), .A2(n15859), .ZN(n15858) );
  AOI22_X1 U14959 ( .A1(n11977), .A2(P2_EAX_REG_25__SCAN_IN), .B1(n9713), .B2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n11969) );
  OAI21_X1 U14960 ( .B1(n11972), .B2(n20670), .A(n11969), .ZN(n15837) );
  AOI22_X1 U14961 ( .A1(n11977), .A2(P2_EAX_REG_26__SCAN_IN), .B1(n9713), .B2(
        P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n11970) );
  OAI21_X1 U14962 ( .B1(n11972), .B2(n20672), .A(n11970), .ZN(n15960) );
  AOI22_X1 U14963 ( .A1(n11977), .A2(P2_EAX_REG_27__SCAN_IN), .B1(n9713), .B2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n11971) );
  OAI21_X1 U14964 ( .B1(n11972), .B2(n20675), .A(n11971), .ZN(n13040) );
  NAND2_X1 U14965 ( .A1(n12037), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n11974) );
  AOI22_X1 U14966 ( .A1(n11977), .A2(P2_EAX_REG_28__SCAN_IN), .B1(n9713), .B2(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n11973) );
  AND2_X1 U14967 ( .A1(n11974), .A2(n11973), .ZN(n14810) );
  INV_X1 U14968 ( .A(n14810), .ZN(n11975) );
  NAND2_X1 U14969 ( .A1(n12037), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n11979) );
  AOI22_X1 U14970 ( .A1(n11977), .A2(P2_EAX_REG_29__SCAN_IN), .B1(n9713), .B2(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n11978) );
  AND2_X1 U14971 ( .A1(n11979), .A2(n11978), .ZN(n15933) );
  INV_X1 U14972 ( .A(n11981), .ZN(n11982) );
  AOI21_X1 U14973 ( .B1(n11983), .B2(n11982), .A(n12041), .ZN(n15144) );
  NAND2_X1 U14974 ( .A1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n14388) );
  NOR2_X1 U14975 ( .A1(n14394), .A2(n14388), .ZN(n16415) );
  NAND2_X1 U14976 ( .A1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n16415), .ZN(
        n17042) );
  NOR2_X1 U14977 ( .A1(n11984), .A2(n17042), .ZN(n12015) );
  INV_X1 U14978 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n17065) );
  NOR2_X1 U14979 ( .A1(n11985), .A2(n20121), .ZN(n11986) );
  INV_X1 U14980 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n16424) );
  NOR2_X1 U14981 ( .A1(n16424), .A2(n14877), .ZN(n13336) );
  INV_X1 U14982 ( .A(n13336), .ZN(n13321) );
  NOR2_X1 U14983 ( .A1(n13340), .A2(n13321), .ZN(n12012) );
  NOR2_X1 U14984 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n13336), .ZN(
        n12010) );
  INV_X1 U14985 ( .A(n12010), .ZN(n12003) );
  INV_X1 U14986 ( .A(n13319), .ZN(n16327) );
  NAND2_X1 U14987 ( .A1(n11988), .A2(n20755), .ZN(n13769) );
  NAND2_X1 U14988 ( .A1(n13769), .A2(n11989), .ZN(n11991) );
  NAND2_X1 U14989 ( .A1(n11991), .A2(n11990), .ZN(n12001) );
  NAND2_X1 U14990 ( .A1(n11993), .A2(n13111), .ZN(n11997) );
  NOR2_X1 U14991 ( .A1(n13111), .A2(n11994), .ZN(n11995) );
  AOI21_X1 U14992 ( .B1(n11997), .B2(n11996), .A(n11995), .ZN(n12000) );
  MUX2_X1 U14993 ( .A(n11998), .B(n10325), .S(n20750), .Z(n11999) );
  NAND2_X1 U14994 ( .A1(n12028), .A2(n12002), .ZN(n12011) );
  NAND2_X1 U14995 ( .A1(n16327), .A2(n12011), .ZN(n16289) );
  OAI211_X1 U14996 ( .C1(n13319), .C2(n12012), .A(n12003), .B(n16289), .ZN(
        n17064) );
  NOR2_X1 U14997 ( .A1(n17065), .A2(n17064), .ZN(n16414) );
  NAND2_X1 U14998 ( .A1(n12015), .A2(n16414), .ZN(n16408) );
  NOR2_X1 U14999 ( .A1(n16408), .A2(n12004), .ZN(n16308) );
  AND2_X1 U15000 ( .A1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n12005) );
  NAND2_X1 U15001 ( .A1(n16308), .A2(n12005), .ZN(n16281) );
  INV_X1 U15002 ( .A(n16262), .ZN(n12006) );
  NAND2_X1 U15003 ( .A1(n12006), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n12007) );
  NOR2_X1 U15004 ( .A1(n16261), .A2(n12007), .ZN(n16239) );
  NOR2_X1 U15005 ( .A1(n10192), .A2(n16222), .ZN(n16219) );
  NAND2_X1 U15006 ( .A1(n16239), .A2(n16219), .ZN(n14812) );
  NOR3_X1 U15007 ( .A1(n10828), .A2(n10829), .A3(n14812), .ZN(n16209) );
  NAND2_X1 U15008 ( .A1(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n16209), .ZN(
        n12043) );
  NAND2_X1 U15009 ( .A1(n19905), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n12032) );
  OAI21_X1 U15010 ( .B1(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n12043), .A(
        n12032), .ZN(n12025) );
  NAND2_X1 U15011 ( .A1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n12008) );
  OR2_X1 U15012 ( .A1(n16206), .A2(n12008), .ZN(n12023) );
  INV_X1 U15013 ( .A(n12009), .ZN(n20028) );
  NOR2_X1 U15014 ( .A1(n12028), .A2(n20028), .ZN(n17067) );
  NOR2_X1 U15015 ( .A1(n16289), .A2(n17067), .ZN(n16413) );
  INV_X1 U15016 ( .A(n16413), .ZN(n12021) );
  NOR2_X1 U15017 ( .A1(n17067), .A2(n17065), .ZN(n12014) );
  NAND2_X1 U15018 ( .A1(n13319), .A2(n12010), .ZN(n13325) );
  INV_X1 U15019 ( .A(n12011), .ZN(n16329) );
  INV_X1 U15020 ( .A(n12012), .ZN(n12013) );
  NAND2_X1 U15021 ( .A1(n16329), .A2(n12013), .ZN(n13322) );
  AND3_X1 U15022 ( .A1(n12014), .A2(n13325), .A3(n13322), .ZN(n17066) );
  NAND3_X1 U15023 ( .A1(n17066), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A3(
        n12015), .ZN(n12016) );
  NAND2_X1 U15024 ( .A1(n12021), .A2(n12016), .ZN(n17033) );
  OR2_X1 U15025 ( .A1(n16413), .A2(n16149), .ZN(n12017) );
  NAND2_X1 U15026 ( .A1(n17033), .A2(n12017), .ZN(n17019) );
  NAND2_X1 U15027 ( .A1(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n16291) );
  NOR2_X1 U15028 ( .A1(n16290), .A2(n16291), .ZN(n12018) );
  NOR2_X1 U15029 ( .A1(n16413), .A2(n12018), .ZN(n12019) );
  OR3_X1 U15030 ( .A1(n17019), .A2(n12019), .A3(n16280), .ZN(n16278) );
  NAND2_X1 U15031 ( .A1(n16278), .A2(n12021), .ZN(n16268) );
  AOI21_X1 U15032 ( .B1(n16289), .B2(n16262), .A(n16243), .ZN(n12020) );
  NAND2_X1 U15033 ( .A1(n16268), .A2(n12020), .ZN(n16251) );
  NAND2_X1 U15034 ( .A1(n16251), .A2(n12021), .ZN(n16234) );
  OR2_X1 U15035 ( .A1(n16413), .A2(n16219), .ZN(n12022) );
  NAND2_X1 U15036 ( .A1(n16234), .A2(n12022), .ZN(n14806) );
  AOI21_X1 U15037 ( .B1(n16289), .B2(n12023), .A(n14806), .ZN(n12047) );
  NOR2_X1 U15038 ( .A1(n12047), .A2(n12027), .ZN(n12024) );
  XNOR2_X1 U15039 ( .A(n16033), .B(n12027), .ZN(n12030) );
  NAND2_X1 U15040 ( .A1(n12028), .A2(n20734), .ZN(n20068) );
  NAND2_X1 U15041 ( .A1(n12030), .A2(n17052), .ZN(n12029) );
  NAND2_X1 U15042 ( .A1(n12030), .A2(n17010), .ZN(n12035) );
  NOR2_X1 U15043 ( .A1(n16845), .A2(n16202), .ZN(n12034) );
  XNOR2_X1 U15044 ( .A(n9827), .B(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16849) );
  INV_X1 U15045 ( .A(n20055), .ZN(n20029) );
  NAND2_X1 U15046 ( .A1(n20029), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12031) );
  OAI211_X1 U15047 ( .C1(n20045), .C2(n16849), .A(n12032), .B(n12031), .ZN(
        n12033) );
  OAI21_X1 U15048 ( .B1(n12036), .B2(n16974), .A(n10197), .ZN(P2_U2984) );
  NAND2_X1 U15049 ( .A1(n12037), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n12039) );
  AOI22_X1 U15050 ( .A1(n11977), .A2(P2_EAX_REG_31__SCAN_IN), .B1(n9713), .B2(
        P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n12038) );
  NAND2_X1 U15051 ( .A1(n12039), .A2(n12038), .ZN(n12040) );
  INV_X1 U15052 ( .A(n12042), .ZN(n12044) );
  INV_X1 U15053 ( .A(n12046), .ZN(n12052) );
  INV_X1 U15054 ( .A(n16289), .ZN(n17077) );
  OAI21_X1 U15055 ( .B1(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n17077), .A(
        n12047), .ZN(n12048) );
  OAI21_X1 U15056 ( .B1(n12092), .B2(n20062), .A(n12049), .ZN(n12050) );
  NAND2_X1 U15057 ( .A1(n12053), .A2(n17052), .ZN(n12054) );
  OAI211_X1 U15058 ( .C1(n12055), .C2(n17071), .A(n10200), .B(n12054), .ZN(
        P2_U3015) );
  OAI21_X1 U15059 ( .B1(n12084), .B2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n12058), .ZN(n16885) );
  AND2_X1 U15060 ( .A1(n9832), .A2(n16082), .ZN(n12059) );
  OR2_X1 U15061 ( .A1(n12059), .A2(n12080), .ZN(n16467) );
  OAI21_X1 U15062 ( .B1(n12078), .B2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        n9832), .ZN(n19751) );
  AOI21_X1 U15063 ( .B1(n12074), .B2(n19768), .A(n12076), .ZN(n19773) );
  AOI21_X1 U15064 ( .B1(n16161), .B2(n12072), .A(n12075), .ZN(n19798) );
  AOI21_X1 U15065 ( .B1(n19816), .B2(n12071), .A(n12073), .ZN(n19822) );
  AOI21_X1 U15066 ( .B1(n16971), .B2(n12069), .A(n9809), .ZN(n19844) );
  AOI21_X1 U15067 ( .B1(n16986), .B2(n12067), .A(n12070), .ZN(n19869) );
  AOI21_X1 U15068 ( .B1(n17007), .B2(n12065), .A(n12068), .ZN(n17000) );
  AOI21_X1 U15069 ( .B1(n16200), .B2(n12063), .A(n12066), .ZN(n19875) );
  AOI21_X1 U15070 ( .B1(n17014), .B2(n12061), .A(n12064), .ZN(n19908) );
  AOI21_X1 U15071 ( .B1(n14786), .B2(n12060), .A(n12062), .ZN(n14782) );
  OAI22_X1 U15072 ( .A1(n20749), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(P2_STATE2_REG_0__SCAN_IN), .ZN(
        n19933) );
  INV_X1 U15073 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n15883) );
  OAI22_X1 U15074 ( .A1(n20749), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(
        n15883), .B2(P2_STATE2_REG_0__SCAN_IN), .ZN(n15879) );
  AND2_X1 U15075 ( .A1(n19933), .A2(n15879), .ZN(n15866) );
  OAI21_X1 U15076 ( .B1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A(n12060), .ZN(n20044) );
  NAND2_X1 U15077 ( .A1(n15866), .A2(n20044), .ZN(n14780) );
  NOR2_X1 U15078 ( .A1(n14782), .A2(n14780), .ZN(n14861) );
  OAI21_X1 U15079 ( .B1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n12062), .A(
        n12061), .ZN(n20041) );
  NAND2_X1 U15080 ( .A1(n14861), .A2(n20041), .ZN(n19906) );
  NOR2_X1 U15081 ( .A1(n19908), .A2(n19906), .ZN(n19892) );
  OAI21_X1 U15082 ( .B1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n12064), .A(
        n12063), .ZN(n19893) );
  NAND2_X1 U15083 ( .A1(n19892), .A2(n19893), .ZN(n19874) );
  NOR2_X1 U15084 ( .A1(n19875), .A2(n19874), .ZN(n14198) );
  OAI21_X1 U15085 ( .B1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n12066), .A(
        n12065), .ZN(n16188) );
  NAND2_X1 U15086 ( .A1(n14198), .A2(n16188), .ZN(n14280) );
  NOR2_X1 U15087 ( .A1(n17000), .A2(n14280), .ZN(n14236) );
  OAI21_X1 U15088 ( .B1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n12068), .A(
        n12067), .ZN(n16999) );
  NAND2_X1 U15089 ( .A1(n14236), .A2(n16999), .ZN(n19867) );
  NOR2_X1 U15090 ( .A1(n19869), .A2(n19867), .ZN(n19850) );
  OAI21_X1 U15091 ( .B1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n12070), .A(
        n12069), .ZN(n19852) );
  NAND2_X1 U15092 ( .A1(n19850), .A2(n19852), .ZN(n19842) );
  NOR2_X1 U15093 ( .A1(n19844), .A2(n19842), .ZN(n19828) );
  OAI21_X1 U15094 ( .B1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n9809), .A(
        n12071), .ZN(n19829) );
  NAND2_X1 U15095 ( .A1(n19828), .A2(n19829), .ZN(n19820) );
  NOR2_X1 U15096 ( .A1(n19822), .A2(n19820), .ZN(n19803) );
  OAI21_X1 U15097 ( .B1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n12073), .A(
        n12072), .ZN(n19804) );
  NAND2_X1 U15098 ( .A1(n19803), .A2(n19804), .ZN(n19793) );
  NOR2_X1 U15099 ( .A1(n19798), .A2(n19793), .ZN(n19792) );
  OAI21_X1 U15100 ( .B1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n12075), .A(
        n12074), .ZN(n19780) );
  NAND2_X1 U15101 ( .A1(n19792), .A2(n19780), .ZN(n19772) );
  NOR2_X1 U15102 ( .A1(n19773), .A2(n19772), .ZN(n19755) );
  NOR2_X1 U15103 ( .A1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n12076), .ZN(
        n12077) );
  NOR2_X1 U15104 ( .A1(n12078), .A2(n12077), .ZN(n19760) );
  INV_X1 U15105 ( .A(n19760), .ZN(n16125) );
  NAND2_X1 U15106 ( .A1(n19755), .A2(n16125), .ZN(n19758) );
  NAND2_X1 U15107 ( .A1(n9718), .A2(n19758), .ZN(n19750) );
  NAND2_X1 U15108 ( .A1(n19751), .A2(n19750), .ZN(n19749) );
  NAND2_X1 U15109 ( .A1(n9718), .A2(n19749), .ZN(n16466) );
  NAND2_X1 U15110 ( .A1(n16467), .A2(n16466), .ZN(n16465) );
  NAND2_X1 U15111 ( .A1(n16465), .A2(n9718), .ZN(n16904) );
  OAI21_X1 U15112 ( .B1(n12080), .B2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n12079), .ZN(n16905) );
  NAND2_X1 U15113 ( .A1(n12079), .A2(n16068), .ZN(n12081) );
  NAND2_X1 U15114 ( .A1(n12082), .A2(n12081), .ZN(n16066) );
  NAND2_X1 U15115 ( .A1(n9718), .A2(n15852), .ZN(n15840) );
  NAND2_X1 U15116 ( .A1(n12082), .A2(n15841), .ZN(n12083) );
  NAND2_X1 U15117 ( .A1(n12086), .A2(n12083), .ZN(n16055) );
  NAND2_X1 U15118 ( .A1(n9718), .A2(n15839), .ZN(n16894) );
  INV_X1 U15119 ( .A(n12084), .ZN(n12088) );
  NAND2_X1 U15120 ( .A1(n12086), .A2(n12085), .ZN(n12087) );
  NAND2_X1 U15121 ( .A1(n12088), .A2(n12087), .ZN(n16895) );
  NAND2_X1 U15122 ( .A1(n9719), .A2(n16893), .ZN(n16884) );
  NAND2_X1 U15123 ( .A1(n16885), .A2(n16884), .ZN(n16883) );
  NAND2_X1 U15124 ( .A1(n16883), .A2(n9719), .ZN(n16871) );
  NAND2_X1 U15125 ( .A1(n12058), .A2(n12089), .ZN(n12090) );
  NAND2_X1 U15126 ( .A1(n12091), .A2(n12090), .ZN(n16872) );
  NAND2_X1 U15127 ( .A1(n9718), .A2(n16870), .ZN(n16860) );
  AOI21_X1 U15128 ( .B1(n16035), .B2(n12091), .A(n9827), .ZN(n16037) );
  INV_X1 U15129 ( .A(n16037), .ZN(n16861) );
  NOR4_X2 U15130 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(P2_STATEBS16_REG_SCAN_IN), .A4(n13792), .ZN(n19910) );
  NAND2_X1 U15131 ( .A1(n19897), .A2(n9719), .ZN(n19932) );
  AND2_X1 U15132 ( .A1(n13734), .A2(n13139), .ZN(n13106) );
  AND2_X1 U15133 ( .A1(n11738), .A2(n13106), .ZN(n20745) );
  AND2_X1 U15134 ( .A1(n20745), .A2(n12093), .ZN(n12102) );
  NAND2_X1 U15135 ( .A1(n11033), .A2(n20748), .ZN(n14204) );
  INV_X1 U15136 ( .A(n14204), .ZN(n12094) );
  INV_X1 U15137 ( .A(n19922), .ZN(n19880) );
  NOR2_X1 U15138 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n12095), .ZN(n12100) );
  AND2_X1 U15139 ( .A1(n12096), .A2(n12100), .ZN(n13795) );
  AND2_X1 U15140 ( .A1(n20745), .A2(n13795), .ZN(n19915) );
  INV_X1 U15141 ( .A(n19915), .ZN(n19914) );
  OAI22_X1 U15142 ( .A1(n12092), .A2(n19880), .B1(n12097), .B2(n19914), .ZN(
        n12111) );
  INV_X1 U15143 ( .A(n12098), .ZN(n12099) );
  NAND2_X1 U15144 ( .A1(n14205), .A2(n9759), .ZN(n13246) );
  INV_X1 U15145 ( .A(n13246), .ZN(n13214) );
  INV_X1 U15146 ( .A(n12100), .ZN(n12101) );
  NAND2_X1 U15147 ( .A1(n13214), .A2(n12101), .ZN(n14207) );
  INV_X1 U15148 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n12107) );
  INV_X1 U15149 ( .A(n12102), .ZN(n12104) );
  NAND2_X1 U15150 ( .A1(P2_EBX_REG_31__SCAN_IN), .A2(n14204), .ZN(n12103) );
  INV_X1 U15151 ( .A(n12105), .ZN(n12106) );
  NAND2_X1 U15152 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n20607), .ZN(n20128) );
  NOR2_X1 U15153 ( .A1(n20616), .A2(n20128), .ZN(n17078) );
  NOR4_X4 U15154 ( .A1(n19905), .A2(n19897), .A3(n20745), .A4(n17078), .ZN(
        n19927) );
  OAI222_X1 U15155 ( .A1(n14207), .A2(n12107), .B1(n19919), .B2(n12106), .C1(
        n20683), .C2(n19887), .ZN(n12109) );
  NOR2_X1 U15156 ( .A1(n19815), .A2(n11038), .ZN(n12108) );
  INV_X1 U15157 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n13067) );
  NAND2_X1 U15158 ( .A1(n16673), .A2(n13067), .ZN(n13058) );
  NOR2_X2 U15159 ( .A1(n16648), .A2(n12114), .ZN(n12117) );
  NAND2_X1 U15160 ( .A1(n15627), .A2(n12115), .ZN(n12116) );
  NOR2_X1 U15161 ( .A1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n12118) );
  AND2_X1 U15162 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15690) );
  NAND2_X1 U15163 ( .A1(n16645), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n13059) );
  INV_X1 U15164 ( .A(n13059), .ZN(n12120) );
  NAND3_X1 U15165 ( .A1(n12139), .A2(n15690), .A3(n12120), .ZN(n12121) );
  OAI21_X1 U15166 ( .B1(n13058), .B2(n12138), .A(n12121), .ZN(n12122) );
  XNOR2_X1 U15167 ( .A(n12122), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15619) );
  AOI22_X1 U15168 ( .A1(n14818), .A2(P1_EBX_REG_30__SCAN_IN), .B1(n14817), 
        .B2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14816) );
  OR2_X1 U15169 ( .A1(n11589), .A2(P1_EBX_REG_28__SCAN_IN), .ZN(n12126) );
  INV_X1 U15170 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15692) );
  NAND2_X1 U15171 ( .A1(n11601), .A2(n15692), .ZN(n12124) );
  INV_X1 U15172 ( .A(P1_EBX_REG_28__SCAN_IN), .ZN(n14725) );
  NAND2_X1 U15173 ( .A1(n13275), .A2(n14725), .ZN(n12123) );
  NAND3_X1 U15174 ( .A1(n12124), .A2(n12132), .A3(n12123), .ZN(n12125) );
  NAND2_X1 U15175 ( .A1(n12126), .A2(n12125), .ZN(n14710) );
  OR2_X1 U15176 ( .A1(n14818), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12127) );
  INV_X1 U15177 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n15471) );
  NAND2_X1 U15178 ( .A1(n13275), .A2(n15471), .ZN(n12129) );
  NAND2_X1 U15179 ( .A1(n12127), .A2(n12129), .ZN(n12131) );
  MUX2_X1 U15180 ( .A(n12131), .B(n12129), .S(n12128), .Z(n13064) );
  NOR2_X1 U15181 ( .A1(n15160), .A2(n20925), .ZN(n12137) );
  INV_X1 U15182 ( .A(n12134), .ZN(n14826) );
  AOI21_X1 U15183 ( .B1(n9914), .B2(n14826), .A(n15696), .ZN(n13068) );
  OAI211_X1 U15184 ( .C1(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n15738), .A(
        n13068), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14827) );
  INV_X1 U15185 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14821) );
  NAND3_X1 U15186 ( .A1(n12135), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n15690), .ZN(n14822) );
  NAND2_X1 U15187 ( .A1(n14821), .A2(n14822), .ZN(n12136) );
  INV_X1 U15188 ( .A(P1_REIP_REG_30__SCAN_IN), .ZN(n15158) );
  NOR2_X1 U15189 ( .A1(n16823), .A2(n15158), .ZN(n15615) );
  NOR2_X1 U15190 ( .A1(n13059), .A2(n14821), .ZN(n12140) );
  XNOR2_X1 U15191 ( .A(n12142), .B(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14830) );
  INV_X1 U15192 ( .A(n12143), .ZN(n12145) );
  NAND2_X1 U15193 ( .A1(n11199), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12300) );
  INV_X1 U15194 ( .A(n12300), .ZN(n12144) );
  NAND2_X1 U15195 ( .A1(n12145), .A2(n12144), .ZN(n12150) );
  INV_X2 U15196 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n21113) );
  INV_X1 U15197 ( .A(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n12147) );
  AND2_X1 U15198 ( .A1(n21113), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n12630) );
  INV_X1 U15199 ( .A(n12630), .ZN(n12240) );
  OAI21_X1 U15200 ( .B1(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n12211), .A(
        n12228), .ZN(n20799) );
  OR2_X1 U15201 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n12600) );
  INV_X1 U15202 ( .A(n12600), .ZN(n12557) );
  NAND2_X1 U15203 ( .A1(n20799), .A2(n12557), .ZN(n12146) );
  OAI21_X1 U15204 ( .B1(n12147), .B2(n12240), .A(n12146), .ZN(n12148) );
  AOI21_X1 U15205 ( .B1(n12626), .B2(P1_EAX_REG_7__SCAN_IN), .A(n12148), .ZN(
        n12149) );
  NAND2_X1 U15206 ( .A1(n12150), .A2(n12149), .ZN(n13995) );
  AOI22_X1 U15207 ( .A1(n12605), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11098), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12154) );
  AOI22_X1 U15208 ( .A1(n9762), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11217), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12153) );
  AOI22_X1 U15209 ( .A1(n12413), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n12539), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12152) );
  AOI22_X1 U15210 ( .A1(n12607), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n11163), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12151) );
  NAND4_X1 U15211 ( .A1(n12154), .A2(n12153), .A3(n12152), .A4(n12151), .ZN(
        n12160) );
  AOI22_X1 U15212 ( .A1(n9715), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12603), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12158) );
  AOI22_X1 U15213 ( .A1(n11278), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n9760), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12157) );
  AOI22_X1 U15214 ( .A1(n12604), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n9745), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12156) );
  AOI22_X1 U15215 ( .A1(n12614), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n12606), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12155) );
  NAND4_X1 U15216 ( .A1(n12158), .A2(n12157), .A3(n12156), .A4(n12155), .ZN(
        n12159) );
  OR2_X1 U15217 ( .A1(n12160), .A2(n12159), .ZN(n12161) );
  NAND2_X1 U15218 ( .A1(n12144), .A2(n12161), .ZN(n12163) );
  XOR2_X1 U15219 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B(n12228), .Z(n14362) );
  AOI22_X1 U15220 ( .A1(n12630), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(
        n12557), .B2(n14362), .ZN(n12162) );
  OAI211_X1 U15221 ( .C1(n12333), .C2(n20885), .A(n12163), .B(n12162), .ZN(
        n13996) );
  NOR2_X1 U15222 ( .A1(n11179), .A2(n21113), .ZN(n12185) );
  INV_X1 U15223 ( .A(n12185), .ZN(n12195) );
  NAND2_X1 U15224 ( .A1(n12626), .A2(P1_EAX_REG_2__SCAN_IN), .ZN(n12166) );
  OAI21_X1 U15225 ( .B1(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A(n12164), .ZN(n14834) );
  OAI21_X1 U15226 ( .B1(n14834), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n21113), 
        .ZN(n12165) );
  OAI211_X1 U15227 ( .C1(n12195), .C2(n13316), .A(n12166), .B(n12165), .ZN(
        n12167) );
  INV_X1 U15228 ( .A(n12167), .ZN(n12168) );
  NAND2_X1 U15229 ( .A1(n12630), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13622) );
  NAND2_X1 U15230 ( .A1(n12169), .A2(n13622), .ZN(n13565) );
  AOI21_X1 U15231 ( .B1(n14398), .B2(n11199), .A(n21113), .ZN(n13344) );
  AOI22_X1 U15232 ( .A1(n12631), .A2(P1_EAX_REG_0__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n21113), .ZN(n12173) );
  OAI21_X1 U15233 ( .B1(n12195), .B2(n10100), .A(n12173), .ZN(n12174) );
  AOI21_X1 U15234 ( .B1(n12172), .B2(n12144), .A(n12174), .ZN(n13345) );
  MUX2_X1 U15235 ( .A(n13344), .B(n12557), .S(n13345), .Z(n13385) );
  NAND2_X1 U15236 ( .A1(n12177), .A2(n12176), .ZN(n12178) );
  NAND2_X1 U15237 ( .A1(n15812), .A2(n12144), .ZN(n12182) );
  NAND2_X1 U15238 ( .A1(n12185), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12180) );
  AOI22_X1 U15239 ( .A1(n12626), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n21113), .ZN(n12179) );
  AND2_X1 U15240 ( .A1(n12180), .A2(n12179), .ZN(n12181) );
  NAND2_X1 U15241 ( .A1(n12182), .A2(n12181), .ZN(n13384) );
  NAND2_X1 U15242 ( .A1(n13385), .A2(n13384), .ZN(n13564) );
  NAND2_X1 U15243 ( .A1(n12184), .A2(n12183), .ZN(n13562) );
  NAND2_X1 U15244 ( .A1(n13562), .A2(n13622), .ZN(n12192) );
  NAND2_X1 U15245 ( .A1(n12185), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12190) );
  NOR2_X1 U15246 ( .A1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n12186), .ZN(
        n12187) );
  NOR2_X1 U15247 ( .A1(n12196), .A2(n12187), .ZN(n13944) );
  INV_X1 U15248 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n13948) );
  OAI22_X1 U15249 ( .A1(n13944), .A2(n12600), .B1(n12240), .B2(n13948), .ZN(
        n12188) );
  AOI21_X1 U15250 ( .B1(n12626), .B2(P1_EAX_REG_3__SCAN_IN), .A(n12188), .ZN(
        n12189) );
  AND2_X1 U15251 ( .A1(n12190), .A2(n12189), .ZN(n12191) );
  NAND2_X1 U15252 ( .A1(n12193), .A2(n12144), .ZN(n12204) );
  AOI22_X1 U15253 ( .A1(n12626), .A2(P1_EAX_REG_4__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n21113), .ZN(n12194) );
  OAI21_X1 U15254 ( .B1(n12195), .B2(n13297), .A(n12194), .ZN(n12202) );
  INV_X1 U15255 ( .A(n12205), .ZN(n12200) );
  INV_X1 U15256 ( .A(n12196), .ZN(n12198) );
  INV_X1 U15257 ( .A(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n12197) );
  NAND2_X1 U15258 ( .A1(n12198), .A2(n12197), .ZN(n12199) );
  NAND2_X1 U15259 ( .A1(n12200), .A2(n12199), .ZN(n20839) );
  AND2_X1 U15260 ( .A1(n20839), .A2(n12557), .ZN(n12201) );
  AOI21_X1 U15261 ( .B1(n12202), .B2(n12600), .A(n12201), .ZN(n12203) );
  NAND2_X1 U15262 ( .A1(n12204), .A2(n12203), .ZN(n13720) );
  OAI21_X1 U15263 ( .B1(n12205), .B2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A(
        n12210), .ZN(n20826) );
  AOI22_X1 U15264 ( .A1(n20826), .A2(n12557), .B1(n12630), .B2(
        P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n12207) );
  NAND2_X1 U15265 ( .A1(n12626), .A2(P1_EAX_REG_5__SCAN_IN), .ZN(n12206) );
  NAND2_X1 U15266 ( .A1(n12210), .A2(n15346), .ZN(n12213) );
  INV_X1 U15267 ( .A(n12211), .ZN(n12212) );
  NAND2_X1 U15268 ( .A1(n12213), .A2(n12212), .ZN(n20812) );
  NAND2_X1 U15269 ( .A1(n20812), .A2(n12557), .ZN(n12214) );
  OAI21_X1 U15270 ( .B1(n15346), .B2(n12240), .A(n12214), .ZN(n12215) );
  AOI21_X1 U15271 ( .B1(n12626), .B2(P1_EAX_REG_6__SCAN_IN), .A(n12215), .ZN(
        n12216) );
  AOI22_X1 U15272 ( .A1(n12603), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n9762), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12221) );
  AOI22_X1 U15273 ( .A1(n11278), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n9760), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12220) );
  AOI22_X1 U15274 ( .A1(n12613), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n9764), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12219) );
  AOI22_X1 U15275 ( .A1(n12413), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n12614), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12218) );
  NAND4_X1 U15276 ( .A1(n12221), .A2(n12220), .A3(n12219), .A4(n12218), .ZN(
        n12227) );
  AOI22_X1 U15277 ( .A1(n9715), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11217), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12225) );
  AOI22_X1 U15278 ( .A1(n12605), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12604), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12224) );
  AOI22_X1 U15279 ( .A1(n12539), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n12606), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12223) );
  AOI22_X1 U15280 ( .A1(n12607), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n11163), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12222) );
  NAND4_X1 U15281 ( .A1(n12225), .A2(n12224), .A3(n12223), .A4(n12222), .ZN(
        n12226) );
  NOR2_X1 U15282 ( .A1(n12227), .A2(n12226), .ZN(n12233) );
  INV_X1 U15283 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n12230) );
  XNOR2_X1 U15284 ( .A(n12234), .B(n12230), .ZN(n14647) );
  NAND2_X1 U15285 ( .A1(n14647), .A2(n12557), .ZN(n12232) );
  AOI22_X1 U15286 ( .A1(n12631), .A2(P1_EAX_REG_9__SCAN_IN), .B1(n12630), .B2(
        P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n12231) );
  OAI211_X1 U15287 ( .C1(n12233), .C2(n12300), .A(n12232), .B(n12231), .ZN(
        n13990) );
  OAI21_X1 U15288 ( .B1(n12235), .B2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n12257), .ZN(n16720) );
  NAND2_X1 U15289 ( .A1(n12236), .A2(n12144), .ZN(n12238) );
  AOI22_X1 U15290 ( .A1(n12626), .A2(P1_EAX_REG_10__SCAN_IN), .B1(n12630), 
        .B2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n12237) );
  NAND2_X1 U15291 ( .A1(n12238), .A2(n12237), .ZN(n12239) );
  AOI21_X1 U15292 ( .B1(n16720), .B2(n12557), .A(n12239), .ZN(n14278) );
  INV_X1 U15293 ( .A(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n14658) );
  XNOR2_X1 U15294 ( .A(n12257), .B(n14658), .ZN(n15682) );
  INV_X1 U15295 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n20879) );
  OAI22_X1 U15296 ( .A1(n12333), .A2(n20879), .B1(n12240), .B2(n14658), .ZN(
        n12241) );
  AOI21_X1 U15297 ( .B1(n15682), .B2(n12557), .A(n12241), .ZN(n12255) );
  INV_X1 U15298 ( .A(n12255), .ZN(n12242) );
  XNOR2_X1 U15299 ( .A(n12254), .B(n12242), .ZN(n14560) );
  AOI22_X1 U15300 ( .A1(n12413), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n12603), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12246) );
  AOI22_X1 U15301 ( .A1(n12613), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n9756), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12245) );
  AOI22_X1 U15302 ( .A1(n12607), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n9750), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12244) );
  AOI22_X1 U15303 ( .A1(n11158), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n9741), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12243) );
  NAND4_X1 U15304 ( .A1(n12246), .A2(n12245), .A3(n12244), .A4(n12243), .ZN(
        n12252) );
  AOI22_X1 U15305 ( .A1(n11222), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n9715), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12250) );
  AOI22_X1 U15306 ( .A1(n9760), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12604), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12249) );
  AOI22_X1 U15307 ( .A1(n12539), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n9737), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12248) );
  AOI22_X1 U15308 ( .A1(n12605), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12612), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12247) );
  NAND4_X1 U15309 ( .A1(n12250), .A2(n12249), .A3(n12248), .A4(n12247), .ZN(
        n12251) );
  OR2_X1 U15310 ( .A1(n12252), .A2(n12251), .ZN(n12253) );
  NAND2_X1 U15311 ( .A1(n12144), .A2(n12253), .ZN(n14561) );
  XNOR2_X1 U15312 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .B(n12286), .ZN(
        n16710) );
  AOI22_X1 U15313 ( .A1(n11278), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n9760), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12261) );
  AOI22_X1 U15314 ( .A1(n12613), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12604), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12260) );
  AOI22_X1 U15315 ( .A1(n12605), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12614), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12259) );
  AOI22_X1 U15316 ( .A1(n9715), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12606), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12258) );
  NAND4_X1 U15317 ( .A1(n12261), .A2(n12260), .A3(n12259), .A4(n12258), .ZN(
        n12267) );
  AOI22_X1 U15318 ( .A1(n12603), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n9762), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12265) );
  AOI22_X1 U15319 ( .A1(n11217), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12539), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12264) );
  AOI22_X1 U15320 ( .A1(n12413), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n9764), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12263) );
  AOI22_X1 U15321 ( .A1(n12607), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11163), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12262) );
  NAND4_X1 U15322 ( .A1(n12265), .A2(n12264), .A3(n12263), .A4(n12262), .ZN(
        n12266) );
  OR2_X1 U15323 ( .A1(n12267), .A2(n12266), .ZN(n12268) );
  AOI22_X1 U15324 ( .A1(n12144), .A2(n12268), .B1(n12630), .B2(
        P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n12270) );
  NAND2_X1 U15325 ( .A1(n12626), .A2(P1_EAX_REG_13__SCAN_IN), .ZN(n12269) );
  OAI211_X1 U15326 ( .C1(n16710), .C2(n12600), .A(n12270), .B(n12269), .ZN(
        n14665) );
  INV_X1 U15327 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n14687) );
  AOI22_X1 U15328 ( .A1(n9715), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n11158), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12274) );
  AOI22_X1 U15329 ( .A1(n11278), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n9760), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12273) );
  AOI22_X1 U15330 ( .A1(n9756), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n12539), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12272) );
  AOI22_X1 U15331 ( .A1(n12604), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n12606), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12271) );
  NAND4_X1 U15332 ( .A1(n12274), .A2(n12273), .A3(n12272), .A4(n12271), .ZN(
        n12280) );
  AOI22_X1 U15333 ( .A1(n12413), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n12605), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12278) );
  AOI22_X1 U15334 ( .A1(n12613), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n9764), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12277) );
  AOI22_X1 U15335 ( .A1(n12603), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n12614), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12276) );
  AOI22_X1 U15336 ( .A1(n12607), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n9737), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12275) );
  NAND4_X1 U15337 ( .A1(n12278), .A2(n12277), .A3(n12276), .A4(n12275), .ZN(
        n12279) );
  OR2_X1 U15338 ( .A1(n12280), .A2(n12279), .ZN(n12281) );
  NAND2_X1 U15339 ( .A1(n12144), .A2(n12281), .ZN(n12284) );
  XNOR2_X1 U15340 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B(n12282), .ZN(
        n16714) );
  AOI22_X1 U15341 ( .A1(n12557), .A2(n16714), .B1(n12630), .B2(
        P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n12283) );
  OAI211_X1 U15342 ( .C1(n12333), .C2(n14687), .A(n12284), .B(n12283), .ZN(
        n14669) );
  AND2_X1 U15343 ( .A1(n14665), .A2(n14669), .ZN(n12285) );
  INV_X1 U15344 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n16625) );
  XNOR2_X1 U15345 ( .A(n12302), .B(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n15671) );
  AOI22_X1 U15346 ( .A1(n12605), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12604), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12290) );
  AOI22_X1 U15347 ( .A1(n11278), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n9762), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12289) );
  AOI22_X1 U15348 ( .A1(n9756), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12539), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12288) );
  AOI22_X1 U15349 ( .A1(n12413), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n9749), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12287) );
  NAND4_X1 U15350 ( .A1(n12290), .A2(n12289), .A3(n12288), .A4(n12287), .ZN(
        n12296) );
  AOI22_X1 U15351 ( .A1(n9715), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n9760), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12294) );
  AOI22_X1 U15352 ( .A1(n12613), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n9745), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12293) );
  AOI22_X1 U15353 ( .A1(n12603), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n9741), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12292) );
  AOI22_X1 U15354 ( .A1(n12607), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n11163), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12291) );
  NAND4_X1 U15355 ( .A1(n12294), .A2(n12293), .A3(n12292), .A4(n12291), .ZN(
        n12295) );
  NOR2_X1 U15356 ( .A1(n12296), .A2(n12295), .ZN(n12299) );
  NAND2_X1 U15357 ( .A1(n12630), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12298) );
  NAND2_X1 U15358 ( .A1(n12626), .A2(P1_EAX_REG_14__SCAN_IN), .ZN(n12297) );
  OAI211_X1 U15359 ( .C1(n12300), .C2(n12299), .A(n12298), .B(n12297), .ZN(
        n12301) );
  AOI21_X1 U15360 ( .B1(n15671), .B2(n12557), .A(n12301), .ZN(n15440) );
  NAND2_X1 U15361 ( .A1(n12302), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12317) );
  XNOR2_X1 U15362 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B(n12317), .ZN(
        n16698) );
  AOI22_X1 U15363 ( .A1(n12413), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n11098), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12306) );
  AOI22_X1 U15364 ( .A1(n9715), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11158), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12305) );
  AOI22_X1 U15365 ( .A1(n12539), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n9749), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12304) );
  AOI22_X1 U15366 ( .A1(n12607), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n11163), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12303) );
  NAND4_X1 U15367 ( .A1(n12306), .A2(n12305), .A3(n12304), .A4(n12303), .ZN(
        n12312) );
  AOI22_X1 U15368 ( .A1(P1_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n12603), .B1(
        n9756), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12310) );
  AOI22_X1 U15369 ( .A1(n11222), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n9760), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12309) );
  AOI22_X1 U15370 ( .A1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n12604), .B1(
        n9745), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12308) );
  AOI22_X1 U15371 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n12605), .B1(
        n12606), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12307) );
  NAND4_X1 U15372 ( .A1(n12310), .A2(n12309), .A3(n12308), .A4(n12307), .ZN(
        n12311) );
  OR2_X1 U15373 ( .A1(n12312), .A2(n12311), .ZN(n12313) );
  AOI22_X1 U15374 ( .A1(n12144), .A2(n12313), .B1(n12630), .B2(
        P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n12315) );
  NAND2_X1 U15375 ( .A1(n12626), .A2(P1_EAX_REG_15__SCAN_IN), .ZN(n12314) );
  OAI211_X1 U15376 ( .C1(n16698), .C2(n12600), .A(n12315), .B(n12314), .ZN(
        n15535) );
  INV_X1 U15377 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n12316) );
  NAND2_X1 U15378 ( .A1(n12408), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12390) );
  INV_X1 U15379 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n15435) );
  INV_X1 U15380 ( .A(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n15657) );
  INV_X1 U15381 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n16573) );
  OR2_X1 U15382 ( .A1(n12318), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12319) );
  AND2_X1 U15383 ( .A1(n12319), .A2(n12448), .ZN(n16662) );
  NAND2_X1 U15384 ( .A1(n12320), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12597) );
  INV_X1 U15385 ( .A(n12597), .ZN(n12623) );
  AOI22_X1 U15386 ( .A1(n12607), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11222), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12324) );
  AOI22_X1 U15387 ( .A1(n9762), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n9760), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12323) );
  AOI22_X1 U15388 ( .A1(n12613), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n9764), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12322) );
  AOI22_X1 U15389 ( .A1(n12539), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n12606), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12321) );
  NAND4_X1 U15390 ( .A1(n12324), .A2(n12323), .A3(n12322), .A4(n12321), .ZN(
        n12330) );
  AOI22_X1 U15391 ( .A1(n12603), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n11217), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12328) );
  AOI22_X1 U15392 ( .A1(n12605), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12604), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12327) );
  AOI22_X1 U15393 ( .A1(n12413), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n9749), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12326) );
  AOI22_X1 U15394 ( .A1(n9715), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n9737), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12325) );
  NAND4_X1 U15395 ( .A1(n12328), .A2(n12327), .A3(n12326), .A4(n12325), .ZN(
        n12329) );
  OR2_X1 U15396 ( .A1(n12330), .A2(n12329), .ZN(n12335) );
  INV_X1 U15397 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n12332) );
  NAND2_X1 U15398 ( .A1(n21113), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12331) );
  OAI211_X1 U15399 ( .C1(n12333), .C2(n12332), .A(n12600), .B(n12331), .ZN(
        n12334) );
  AOI21_X1 U15400 ( .B1(n12623), .B2(n12335), .A(n12334), .ZN(n12336) );
  AOI21_X1 U15401 ( .B1(n16662), .B2(n12557), .A(n12336), .ZN(n15507) );
  NAND2_X1 U15402 ( .A1(n12597), .A2(n12600), .ZN(n12438) );
  AOI22_X1 U15403 ( .A1(n12603), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n9760), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12342) );
  AOI22_X1 U15404 ( .A1(n12613), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12606), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12341) );
  AOI22_X1 U15405 ( .A1(n9715), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n9750), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12340) );
  NAND2_X1 U15406 ( .A1(n9764), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n12338) );
  NAND2_X1 U15407 ( .A1(n11163), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n12337) );
  AND3_X1 U15408 ( .A1(n12338), .A2(n12600), .A3(n12337), .ZN(n12339) );
  NAND4_X1 U15409 ( .A1(n12342), .A2(n12341), .A3(n12340), .A4(n12339), .ZN(
        n12348) );
  AOI22_X1 U15410 ( .A1(n12605), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n9762), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12346) );
  AOI22_X1 U15411 ( .A1(n12607), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n9756), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12345) );
  AOI22_X1 U15412 ( .A1(n11222), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12413), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12344) );
  AOI22_X1 U15413 ( .A1(n12539), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n12604), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12343) );
  NAND4_X1 U15414 ( .A1(n12346), .A2(n12345), .A3(n12344), .A4(n12343), .ZN(
        n12347) );
  OR2_X1 U15415 ( .A1(n12348), .A2(n12347), .ZN(n12349) );
  NAND2_X1 U15416 ( .A1(n12438), .A2(n12349), .ZN(n12352) );
  AOI22_X1 U15417 ( .A1(n12631), .A2(P1_EAX_REG_20__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n21113), .ZN(n12351) );
  XNOR2_X1 U15418 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B(n12368), .ZN(
        n16563) );
  AND2_X1 U15419 ( .A1(n12557), .A2(n16563), .ZN(n12350) );
  AOI21_X1 U15420 ( .B1(n12352), .B2(n12351), .A(n12350), .ZN(n12353) );
  INV_X1 U15421 ( .A(n12353), .ZN(n15512) );
  AOI22_X1 U15422 ( .A1(n12607), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11278), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12357) );
  AOI22_X1 U15423 ( .A1(n9762), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11217), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12356) );
  AOI22_X1 U15424 ( .A1(n12605), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12604), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12355) );
  AOI22_X1 U15425 ( .A1(n12539), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n12614), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12354) );
  NAND4_X1 U15426 ( .A1(n12357), .A2(n12356), .A3(n12355), .A4(n12354), .ZN(
        n12363) );
  AOI22_X1 U15427 ( .A1(n9715), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12603), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12361) );
  AOI22_X1 U15428 ( .A1(n12613), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n9745), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12360) );
  AOI22_X1 U15429 ( .A1(n12413), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n9741), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12359) );
  AOI22_X1 U15430 ( .A1(n9760), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(n9737), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12358) );
  NAND4_X1 U15431 ( .A1(n12361), .A2(n12360), .A3(n12359), .A4(n12358), .ZN(
        n12362) );
  NOR2_X1 U15432 ( .A1(n12363), .A2(n12362), .ZN(n12367) );
  NAND2_X1 U15433 ( .A1(n21113), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n12364) );
  NAND2_X1 U15434 ( .A1(n12600), .A2(n12364), .ZN(n12365) );
  AOI21_X1 U15435 ( .B1(n12626), .B2(P1_EAX_REG_19__SCAN_IN), .A(n12365), .ZN(
        n12366) );
  OAI21_X1 U15436 ( .B1(n12597), .B2(n12367), .A(n12366), .ZN(n12370) );
  OAI21_X1 U15437 ( .B1(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n12372), .A(
        n12368), .ZN(n16681) );
  OR2_X1 U15438 ( .A1(n12600), .A2(n16681), .ZN(n12369) );
  AND2_X1 U15439 ( .A1(n12370), .A2(n12369), .ZN(n15581) );
  INV_X1 U15440 ( .A(n15581), .ZN(n12406) );
  NAND2_X1 U15441 ( .A1(n12371), .A2(n15657), .ZN(n12374) );
  INV_X1 U15442 ( .A(n12372), .ZN(n12373) );
  NAND2_X1 U15443 ( .A1(n12374), .A2(n12373), .ZN(n15655) );
  AOI22_X1 U15444 ( .A1(n12607), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12603), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12378) );
  AOI22_X1 U15445 ( .A1(n11278), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12605), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12377) );
  AOI22_X1 U15446 ( .A1(n11217), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12604), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12376) );
  AOI22_X1 U15447 ( .A1(n9760), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12614), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12375) );
  NAND4_X1 U15448 ( .A1(n12378), .A2(n12377), .A3(n12376), .A4(n12375), .ZN(
        n12386) );
  AOI22_X1 U15449 ( .A1(n12413), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n9762), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12384) );
  AOI22_X1 U15450 ( .A1(n9715), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12539), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12383) );
  AOI22_X1 U15451 ( .A1(n12613), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n9741), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12382) );
  NAND2_X1 U15452 ( .A1(n9764), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n12380) );
  NAND2_X1 U15453 ( .A1(n9737), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n12379) );
  AND3_X1 U15454 ( .A1(n12380), .A2(n12600), .A3(n12379), .ZN(n12381) );
  NAND4_X1 U15455 ( .A1(n12384), .A2(n12383), .A3(n12382), .A4(n12381), .ZN(
        n12385) );
  OAI21_X1 U15456 ( .B1(n12386), .B2(n12385), .A(n12438), .ZN(n12388) );
  AOI22_X1 U15457 ( .A1(n12631), .A2(P1_EAX_REG_18__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n21113), .ZN(n12387) );
  NAND2_X1 U15458 ( .A1(n12388), .A2(n12387), .ZN(n12389) );
  OAI21_X1 U15459 ( .B1(n15655), .B2(n12600), .A(n12389), .ZN(n15517) );
  XNOR2_X1 U15460 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B(n12390), .ZN(
        n16682) );
  INV_X1 U15461 ( .A(n16682), .ZN(n12405) );
  AOI22_X1 U15462 ( .A1(n12607), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n11278), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12394) );
  AOI22_X1 U15463 ( .A1(n12603), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n11217), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12393) );
  AOI22_X1 U15464 ( .A1(n12413), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n12604), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12392) );
  AOI22_X1 U15465 ( .A1(n12539), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n12614), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12391) );
  NAND4_X1 U15466 ( .A1(n12394), .A2(n12393), .A3(n12392), .A4(n12391), .ZN(
        n12401) );
  AOI22_X1 U15467 ( .A1(n9715), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11158), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12399) );
  AOI22_X1 U15468 ( .A1(n12613), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n9764), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12398) );
  AOI22_X1 U15469 ( .A1(n12605), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n9741), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12397) );
  AOI22_X1 U15470 ( .A1(n9760), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11163), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12396) );
  NAND4_X1 U15471 ( .A1(n12399), .A2(n12398), .A3(n12397), .A4(n12396), .ZN(
        n12400) );
  NOR2_X1 U15472 ( .A1(n12401), .A2(n12400), .ZN(n12403) );
  AOI22_X1 U15473 ( .A1(n12631), .A2(P1_EAX_REG_17__SCAN_IN), .B1(n12630), 
        .B2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n12402) );
  OAI21_X1 U15474 ( .B1(n12597), .B2(n12403), .A(n12402), .ZN(n12404) );
  AOI21_X1 U15475 ( .B1(n12405), .B2(n12557), .A(n12404), .ZN(n15430) );
  OR2_X1 U15476 ( .A1(n15517), .A2(n15430), .ZN(n15519) );
  INV_X1 U15477 ( .A(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n12407) );
  XNOR2_X1 U15478 ( .A(n12408), .B(n12407), .ZN(n16694) );
  NAND2_X1 U15479 ( .A1(n16694), .A2(n12557), .ZN(n12425) );
  AOI22_X1 U15480 ( .A1(n12605), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11217), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12412) );
  AOI22_X1 U15481 ( .A1(n12607), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12603), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12411) );
  AOI22_X1 U15482 ( .A1(n9762), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12539), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12410) );
  AOI22_X1 U15483 ( .A1(n9715), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12612), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12409) );
  NAND4_X1 U15484 ( .A1(n12412), .A2(n12411), .A3(n12410), .A4(n12409), .ZN(
        n12421) );
  AOI22_X1 U15485 ( .A1(n12613), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n9760), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12419) );
  NAND2_X1 U15486 ( .A1(n12413), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n12415) );
  NAND2_X1 U15487 ( .A1(n9737), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n12414) );
  AND3_X1 U15488 ( .A1(n12415), .A2(n12600), .A3(n12414), .ZN(n12418) );
  AOI22_X1 U15489 ( .A1(n12604), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12614), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12417) );
  AOI22_X1 U15490 ( .A1(n11278), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n9741), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12416) );
  NAND4_X1 U15491 ( .A1(n12419), .A2(n12418), .A3(n12417), .A4(n12416), .ZN(
        n12420) );
  OAI21_X1 U15492 ( .B1(n12421), .B2(n12420), .A(n12438), .ZN(n12423) );
  AOI22_X1 U15493 ( .A1(n12631), .A2(P1_EAX_REG_16__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n21113), .ZN(n12422) );
  NAND2_X1 U15494 ( .A1(n12423), .A2(n12422), .ZN(n12424) );
  NAND2_X1 U15495 ( .A1(n12425), .A2(n12424), .ZN(n15530) );
  NOR2_X1 U15496 ( .A1(n12426), .A2(n15530), .ZN(n15506) );
  AND2_X1 U15497 ( .A1(n15507), .A2(n15506), .ZN(n12427) );
  INV_X1 U15498 ( .A(n15499), .ZN(n12446) );
  AOI22_X1 U15499 ( .A1(n12413), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11158), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12431) );
  AOI22_X1 U15500 ( .A1(n12607), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12603), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12430) );
  AOI22_X1 U15501 ( .A1(n11222), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11098), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12429) );
  AOI22_X1 U15502 ( .A1(n12604), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n9741), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12428) );
  NAND4_X1 U15503 ( .A1(n12431), .A2(n12430), .A3(n12429), .A4(n12428), .ZN(
        n12440) );
  AOI22_X1 U15504 ( .A1(n11217), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n9760), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12437) );
  NAND2_X1 U15505 ( .A1(n12605), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n12433) );
  NAND2_X1 U15506 ( .A1(n11163), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n12432) );
  AND3_X1 U15507 ( .A1(n12433), .A2(n12600), .A3(n12432), .ZN(n12436) );
  AOI22_X1 U15508 ( .A1(n9715), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12614), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12435) );
  AOI22_X1 U15509 ( .A1(n12539), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n12612), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12434) );
  NAND4_X1 U15510 ( .A1(n12437), .A2(n12436), .A3(n12435), .A4(n12434), .ZN(
        n12439) );
  OAI21_X1 U15511 ( .B1(n12440), .B2(n12439), .A(n12438), .ZN(n12442) );
  AOI22_X1 U15512 ( .A1(n12626), .A2(P1_EAX_REG_22__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n21113), .ZN(n12441) );
  NAND2_X1 U15513 ( .A1(n12442), .A2(n12441), .ZN(n12444) );
  XNOR2_X1 U15514 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B(n12448), .ZN(
        n16549) );
  NAND2_X1 U15515 ( .A1(n16549), .A2(n12557), .ZN(n12443) );
  NAND2_X1 U15516 ( .A1(n12444), .A2(n12443), .ZN(n15500) );
  INV_X1 U15517 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n12447) );
  OR2_X1 U15518 ( .A1(n12449), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n12450) );
  NAND2_X1 U15519 ( .A1(n12450), .A2(n12494), .ZN(n16660) );
  AOI22_X1 U15520 ( .A1(n12605), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n9745), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12454) );
  AOI22_X1 U15521 ( .A1(n12413), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n12614), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12453) );
  AOI22_X1 U15522 ( .A1(n9762), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12606), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12452) );
  AOI22_X1 U15523 ( .A1(n11278), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n9737), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12451) );
  NAND4_X1 U15524 ( .A1(n12454), .A2(n12453), .A3(n12452), .A4(n12451), .ZN(
        n12460) );
  AOI22_X1 U15525 ( .A1(n9715), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12603), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12458) );
  AOI22_X1 U15526 ( .A1(n12607), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n9760), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12457) );
  AOI22_X1 U15527 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n12613), .B1(
        n12604), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12456) );
  AOI22_X1 U15528 ( .A1(n11217), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12539), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12455) );
  NAND4_X1 U15529 ( .A1(n12458), .A2(n12457), .A3(n12456), .A4(n12455), .ZN(
        n12459) );
  NOR2_X1 U15530 ( .A1(n12460), .A2(n12459), .ZN(n12476) );
  AOI22_X1 U15531 ( .A1(n12413), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12605), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12464) );
  AOI22_X1 U15532 ( .A1(n9762), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11217), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12463) );
  AOI22_X1 U15533 ( .A1(n12604), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n9764), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12462) );
  AOI22_X1 U15534 ( .A1(n9715), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n11163), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12461) );
  NAND4_X1 U15535 ( .A1(n12464), .A2(n12463), .A3(n12462), .A4(n12461), .ZN(
        n12470) );
  AOI22_X1 U15536 ( .A1(n12607), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11278), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12468) );
  AOI22_X1 U15537 ( .A1(n12603), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n9760), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12467) );
  AOI22_X1 U15538 ( .A1(n12613), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12614), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12466) );
  AOI22_X1 U15539 ( .A1(n12539), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n9741), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12465) );
  NAND4_X1 U15540 ( .A1(n12468), .A2(n12467), .A3(n12466), .A4(n12465), .ZN(
        n12469) );
  NOR2_X1 U15541 ( .A1(n12470), .A2(n12469), .ZN(n12475) );
  XNOR2_X1 U15542 ( .A(n12476), .B(n12475), .ZN(n12473) );
  INV_X1 U15543 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n15391) );
  AOI21_X1 U15544 ( .B1(n15391), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n12471) );
  AOI21_X1 U15545 ( .B1(n12626), .B2(P1_EAX_REG_23__SCAN_IN), .A(n12471), .ZN(
        n12472) );
  OAI21_X1 U15546 ( .B1(n12597), .B2(n12473), .A(n12472), .ZN(n12474) );
  OAI21_X1 U15547 ( .B1(n16660), .B2(n12600), .A(n12474), .ZN(n15491) );
  NOR2_X1 U15548 ( .A1(n12476), .A2(n12475), .ZN(n12508) );
  INV_X1 U15549 ( .A(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n15323) );
  AOI22_X1 U15550 ( .A1(n12603), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n11217), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12480) );
  AOI22_X1 U15551 ( .A1(n9715), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n9762), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12479) );
  AOI22_X1 U15552 ( .A1(n11278), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n9760), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12478) );
  AOI22_X1 U15553 ( .A1(n12607), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11163), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12477) );
  NAND4_X1 U15554 ( .A1(n12480), .A2(n12479), .A3(n12478), .A4(n12477), .ZN(
        n12486) );
  AOI22_X1 U15555 ( .A1(n12605), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12613), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12484) );
  AOI22_X1 U15556 ( .A1(n12604), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n9745), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12483) );
  AOI22_X1 U15557 ( .A1(n12413), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n12614), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12482) );
  AOI22_X1 U15558 ( .A1(n12539), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n9741), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12481) );
  NAND4_X1 U15559 ( .A1(n12484), .A2(n12483), .A3(n12482), .A4(n12481), .ZN(
        n12485) );
  OR2_X1 U15560 ( .A1(n12486), .A2(n12485), .ZN(n12507) );
  INV_X1 U15561 ( .A(n12507), .ZN(n12487) );
  XNOR2_X1 U15562 ( .A(n12508), .B(n12487), .ZN(n12488) );
  NAND2_X1 U15563 ( .A1(n12488), .A2(n12623), .ZN(n12493) );
  INV_X1 U15564 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n12489) );
  AOI21_X1 U15565 ( .B1(n12489), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n12490) );
  AOI21_X1 U15566 ( .B1(n12626), .B2(P1_EAX_REG_24__SCAN_IN), .A(n12490), .ZN(
        n12492) );
  XNOR2_X1 U15567 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .B(n12494), .ZN(
        n16532) );
  AND2_X1 U15568 ( .A1(n12557), .A2(n16532), .ZN(n12491) );
  AOI21_X1 U15569 ( .B1(n12493), .B2(n12492), .A(n12491), .ZN(n15484) );
  OR2_X1 U15570 ( .A1(n12495), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n12496) );
  NAND2_X1 U15571 ( .A1(n12496), .A2(n12552), .ZN(n16653) );
  AOI22_X1 U15572 ( .A1(n12603), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n11217), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12500) );
  AOI22_X1 U15573 ( .A1(n9715), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n9762), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12499) );
  AOI22_X1 U15574 ( .A1(n12613), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n9741), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12498) );
  AOI22_X1 U15575 ( .A1(n12607), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n9737), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12497) );
  NAND4_X1 U15576 ( .A1(n12500), .A2(n12499), .A3(n12498), .A4(n12497), .ZN(
        n12506) );
  AOI22_X1 U15577 ( .A1(n12413), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12605), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12504) );
  AOI22_X1 U15578 ( .A1(n11278), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n9760), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12503) );
  AOI22_X1 U15579 ( .A1(n12604), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n9745), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12502) );
  AOI22_X1 U15580 ( .A1(n12539), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n9750), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12501) );
  NAND4_X1 U15581 ( .A1(n12504), .A2(n12503), .A3(n12502), .A4(n12501), .ZN(
        n12505) );
  NOR2_X1 U15582 ( .A1(n12506), .A2(n12505), .ZN(n12516) );
  NAND2_X1 U15583 ( .A1(n12508), .A2(n12507), .ZN(n12515) );
  XNOR2_X1 U15584 ( .A(n12516), .B(n12515), .ZN(n12512) );
  INV_X1 U15585 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n12509) );
  AOI21_X1 U15586 ( .B1(n12509), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n12510) );
  AOI21_X1 U15587 ( .B1(n12631), .B2(P1_EAX_REG_25__SCAN_IN), .A(n12510), .ZN(
        n12511) );
  OAI21_X1 U15588 ( .B1(n12512), .B2(n12597), .A(n12511), .ZN(n12513) );
  OAI21_X1 U15589 ( .B1(n16653), .B2(n12600), .A(n12513), .ZN(n15477) );
  INV_X1 U15590 ( .A(n15477), .ZN(n12514) );
  NOR2_X1 U15591 ( .A1(n12516), .A2(n12515), .ZN(n12547) );
  AOI22_X1 U15592 ( .A1(n12603), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n9756), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12520) );
  AOI22_X1 U15593 ( .A1(n9715), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n9762), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12519) );
  AOI22_X1 U15594 ( .A1(n11222), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n9760), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12518) );
  AOI22_X1 U15595 ( .A1(n12607), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n9737), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12517) );
  NAND4_X1 U15596 ( .A1(n12520), .A2(n12519), .A3(n12518), .A4(n12517), .ZN(
        n12526) );
  AOI22_X1 U15597 ( .A1(n12605), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11098), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12524) );
  AOI22_X1 U15598 ( .A1(n12604), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n9745), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12523) );
  AOI22_X1 U15599 ( .A1(n12413), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12614), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12522) );
  AOI22_X1 U15600 ( .A1(n12539), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n9741), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12521) );
  NAND4_X1 U15601 ( .A1(n12524), .A2(n12523), .A3(n12522), .A4(n12521), .ZN(
        n12525) );
  OR2_X1 U15602 ( .A1(n12526), .A2(n12525), .ZN(n12546) );
  XNOR2_X1 U15603 ( .A(n12547), .B(n12546), .ZN(n12530) );
  NAND2_X1 U15604 ( .A1(n21113), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12527) );
  NAND2_X1 U15605 ( .A1(n12600), .A2(n12527), .ZN(n12528) );
  AOI21_X1 U15606 ( .B1(n12631), .B2(P1_EAX_REG_26__SCAN_IN), .A(n12528), .ZN(
        n12529) );
  OAI21_X1 U15607 ( .B1(n12530), .B2(n12597), .A(n12529), .ZN(n12532) );
  XNOR2_X1 U15608 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .B(n12552), .ZN(
        n15624) );
  NAND2_X1 U15609 ( .A1(n12557), .A2(n15624), .ZN(n12531) );
  NAND2_X1 U15610 ( .A1(n12532), .A2(n12531), .ZN(n15182) );
  AOI22_X1 U15611 ( .A1(n11278), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n9715), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12538) );
  AOI22_X1 U15612 ( .A1(n12613), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12612), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12537) );
  AOI22_X1 U15613 ( .A1(n11390), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n9749), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12536) );
  AOI22_X1 U15614 ( .A1(n12607), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11163), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12535) );
  NAND4_X1 U15615 ( .A1(n12538), .A2(n12537), .A3(n12536), .A4(n12535), .ZN(
        n12545) );
  AOI22_X1 U15616 ( .A1(n12603), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n11217), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12543) );
  AOI22_X1 U15617 ( .A1(n9762), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n9760), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12542) );
  AOI22_X1 U15618 ( .A1(n12413), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n12604), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12541) );
  AOI22_X1 U15619 ( .A1(n12539), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n12606), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12540) );
  NAND4_X1 U15620 ( .A1(n12543), .A2(n12542), .A3(n12541), .A4(n12540), .ZN(
        n12544) );
  NOR2_X1 U15621 ( .A1(n12545), .A2(n12544), .ZN(n12572) );
  NAND2_X1 U15622 ( .A1(n12547), .A2(n12546), .ZN(n12571) );
  XNOR2_X1 U15623 ( .A(n12572), .B(n12571), .ZN(n12551) );
  NAND2_X1 U15624 ( .A1(n21113), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n12548) );
  NAND2_X1 U15625 ( .A1(n12600), .A2(n12548), .ZN(n12549) );
  AOI21_X1 U15626 ( .B1(n12626), .B2(P1_EAX_REG_27__SCAN_IN), .A(n12549), .ZN(
        n12550) );
  OAI21_X1 U15627 ( .B1(n12551), .B2(n12597), .A(n12550), .ZN(n12559) );
  INV_X1 U15628 ( .A(n12552), .ZN(n12553) );
  INV_X1 U15629 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n14761) );
  INV_X1 U15630 ( .A(n12554), .ZN(n12555) );
  NAND2_X1 U15631 ( .A1(n14761), .A2(n12555), .ZN(n12556) );
  AND2_X1 U15632 ( .A1(n12577), .A2(n12556), .ZN(n15173) );
  NAND2_X1 U15633 ( .A1(n15173), .A2(n12557), .ZN(n12558) );
  NAND2_X1 U15634 ( .A1(n12559), .A2(n12558), .ZN(n14764) );
  AOI22_X1 U15635 ( .A1(n12603), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11217), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12564) );
  AOI22_X1 U15636 ( .A1(n9715), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n11158), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12563) );
  AOI22_X1 U15637 ( .A1(n11222), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n9760), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12562) );
  AOI22_X1 U15638 ( .A1(n12607), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11163), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12561) );
  NAND4_X1 U15639 ( .A1(n12564), .A2(n12563), .A3(n12562), .A4(n12561), .ZN(
        n12570) );
  AOI22_X1 U15640 ( .A1(n11390), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11098), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12568) );
  AOI22_X1 U15641 ( .A1(n12604), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12612), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12567) );
  AOI22_X1 U15642 ( .A1(n12413), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12614), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12566) );
  AOI22_X1 U15643 ( .A1(n12539), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n12606), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12565) );
  NAND4_X1 U15644 ( .A1(n12568), .A2(n12567), .A3(n12566), .A4(n12565), .ZN(
        n12569) );
  OR2_X1 U15645 ( .A1(n12570), .A2(n12569), .ZN(n12582) );
  NOR2_X1 U15646 ( .A1(n12572), .A2(n12571), .ZN(n12583) );
  XOR2_X1 U15647 ( .A(n12582), .B(n12583), .Z(n12573) );
  NAND2_X1 U15648 ( .A1(n12573), .A2(n12623), .ZN(n12576) );
  INV_X1 U15649 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n13024) );
  NOR2_X1 U15650 ( .A1(n13024), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12574) );
  AOI211_X1 U15651 ( .C1(n12626), .C2(P1_EAX_REG_28__SCAN_IN), .A(n12557), .B(
        n12574), .ZN(n12575) );
  XNOR2_X1 U15652 ( .A(n12577), .B(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14723) );
  AOI22_X1 U15653 ( .A1(n12576), .A2(n12575), .B1(n12557), .B2(n14723), .ZN(
        n13016) );
  NAND2_X1 U15654 ( .A1(n12578), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12640) );
  INV_X1 U15655 ( .A(n12578), .ZN(n12580) );
  INV_X1 U15656 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n12579) );
  NAND2_X1 U15657 ( .A1(n12580), .A2(n12579), .ZN(n12581) );
  NAND2_X1 U15658 ( .A1(n12640), .A2(n12581), .ZN(n15163) );
  NAND2_X1 U15659 ( .A1(n12583), .A2(n12582), .ZN(n12601) );
  AOI22_X1 U15660 ( .A1(n12413), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12605), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12587) );
  AOI22_X1 U15661 ( .A1(n9715), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n9760), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12586) );
  AOI22_X1 U15662 ( .A1(n9762), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12606), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12585) );
  AOI22_X1 U15663 ( .A1(n12607), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11163), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12584) );
  NAND4_X1 U15664 ( .A1(n12587), .A2(n12586), .A3(n12585), .A4(n12584), .ZN(
        n12594) );
  AOI22_X1 U15665 ( .A1(n11278), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12603), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12592) );
  AOI22_X1 U15666 ( .A1(n9756), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12539), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12591) );
  AOI22_X1 U15667 ( .A1(n12613), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n9749), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12590) );
  AOI22_X1 U15668 ( .A1(n12604), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12612), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12589) );
  NAND4_X1 U15669 ( .A1(n12592), .A2(n12591), .A3(n12590), .A4(n12589), .ZN(
        n12593) );
  NOR2_X1 U15670 ( .A1(n12594), .A2(n12593), .ZN(n12602) );
  XNOR2_X1 U15671 ( .A(n12601), .B(n12602), .ZN(n12598) );
  INV_X1 U15672 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n21118) );
  OAI21_X1 U15673 ( .B1(n21118), .B2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n21113), .ZN(n12596) );
  NAND2_X1 U15674 ( .A1(n12631), .A2(P1_EAX_REG_29__SCAN_IN), .ZN(n12595) );
  OAI211_X1 U15675 ( .C1(n12598), .C2(n12597), .A(n12596), .B(n12595), .ZN(
        n12599) );
  OAI21_X1 U15676 ( .B1(n12600), .B2(n15163), .A(n12599), .ZN(n14735) );
  NOR2_X1 U15677 ( .A1(n12602), .A2(n12601), .ZN(n12622) );
  AOI22_X1 U15678 ( .A1(n11222), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12603), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12611) );
  AOI22_X1 U15679 ( .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n12605), .B1(
        n12604), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12610) );
  AOI22_X1 U15680 ( .A1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n12539), .B1(
        n9741), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12609) );
  AOI22_X1 U15681 ( .A1(n12607), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11163), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12608) );
  NAND4_X1 U15682 ( .A1(n12611), .A2(n12610), .A3(n12609), .A4(n12608), .ZN(
        n12620) );
  AOI22_X1 U15683 ( .A1(P1_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n9762), .B1(
        n11217), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12618) );
  AOI22_X1 U15684 ( .A1(P1_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n9715), .B1(
        n9760), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12617) );
  AOI22_X1 U15685 ( .A1(n12613), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12612), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12616) );
  AOI22_X1 U15686 ( .A1(n12413), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n12614), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12615) );
  NAND4_X1 U15687 ( .A1(n12618), .A2(n12617), .A3(n12616), .A4(n12615), .ZN(
        n12619) );
  NOR2_X1 U15688 ( .A1(n12620), .A2(n12619), .ZN(n12621) );
  XNOR2_X1 U15689 ( .A(n12622), .B(n12621), .ZN(n12624) );
  NAND2_X1 U15690 ( .A1(n12624), .A2(n12623), .ZN(n12629) );
  INV_X1 U15691 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n15613) );
  AOI21_X1 U15692 ( .B1(n15613), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n12625) );
  AOI21_X1 U15693 ( .B1(n12626), .B2(P1_EAX_REG_30__SCAN_IN), .A(n12625), .ZN(
        n12628) );
  XNOR2_X1 U15694 ( .A(n12640), .B(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15616) );
  AND2_X1 U15695 ( .A1(n15616), .A2(n12557), .ZN(n12627) );
  AOI21_X1 U15696 ( .B1(n12629), .B2(n12628), .A(n12627), .ZN(n13047) );
  NAND2_X1 U15697 ( .A1(n14734), .A2(n13047), .ZN(n12634) );
  AOI22_X1 U15698 ( .A1(n12631), .A2(P1_EAX_REG_31__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n12630), .ZN(n12632) );
  INV_X1 U15699 ( .A(n12632), .ZN(n12633) );
  NAND3_X1 U15700 ( .A1(n9954), .A2(P1_STATEBS16_REG_SCAN_IN), .A3(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n16833) );
  INV_X1 U15701 ( .A(n16833), .ZN(n12635) );
  OR2_X1 U15702 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(P1_STATE2_REG_2__SCAN_IN), 
        .ZN(n21122) );
  INV_X1 U15703 ( .A(n21122), .ZN(n21085) );
  NAND2_X1 U15704 ( .A1(n12635), .A2(n21085), .ZN(n16700) );
  INV_X1 U15705 ( .A(n16700), .ZN(n16739) );
  NAND2_X1 U15706 ( .A1(n15148), .A2(n16739), .ZN(n12645) );
  NAND2_X1 U15707 ( .A1(n21122), .A2(n12636), .ZN(n21286) );
  NAND2_X1 U15708 ( .A1(n21286), .A2(n9954), .ZN(n12637) );
  NAND2_X1 U15709 ( .A1(n9954), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12639) );
  NAND2_X1 U15710 ( .A1(n21118), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n12638) );
  NAND2_X1 U15711 ( .A1(n12639), .A2(n12638), .ZN(n13477) );
  INV_X1 U15712 ( .A(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n15151) );
  XNOR2_X1 U15713 ( .A(n12641), .B(n15151), .ZN(n13942) );
  INV_X1 U15714 ( .A(P1_REIP_REG_31__SCAN_IN), .ZN(n21255) );
  NOR2_X1 U15715 ( .A1(n16823), .A2(n21255), .ZN(n14823) );
  AOI21_X1 U15716 ( .B1(n16734), .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n14823), .ZN(n12642) );
  OAI21_X1 U15717 ( .B1(n16743), .B2(n13942), .A(n12642), .ZN(n12643) );
  OAI211_X1 U15718 ( .C1(n14830), .C2(n20773), .A(n12645), .B(n12644), .ZN(
        P1_U2968) );
  NAND4_X1 U15719 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A4(
        P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n18506) );
  INV_X1 U15720 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n18542) );
  INV_X1 U15721 ( .A(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n18530) );
  NOR2_X1 U15722 ( .A1(n18542), .A2(n18530), .ZN(n18524) );
  NAND2_X1 U15723 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n18484) );
  NAND2_X1 U15724 ( .A1(n18468), .A2(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n18446) );
  NAND2_X1 U15725 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n18447) );
  NAND2_X1 U15726 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n18410) );
  NAND2_X1 U15727 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n18368) );
  INV_X1 U15728 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n18347) );
  INV_X1 U15729 ( .A(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n18337) );
  INV_X1 U15730 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n17615) );
  XOR2_X1 U15731 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B(n12658), .Z(
        n17289) );
  INV_X1 U15732 ( .A(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n13101) );
  NOR2_X1 U15733 ( .A1(n17615), .A2(n9770), .ZN(n12649) );
  NAND3_X1 U15734 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A3(n12649), .ZN(n18322) );
  NOR2_X1 U15735 ( .A1(n13101), .A2(n18322), .ZN(n12648) );
  NAND2_X1 U15736 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n12648), .ZN(
        n12647) );
  NOR2_X1 U15737 ( .A1(n18337), .A2(n12647), .ZN(n17098) );
  INV_X1 U15738 ( .A(n17098), .ZN(n12646) );
  AOI21_X1 U15739 ( .B1(n10042), .B2(n12646), .A(n12658), .ZN(n17300) );
  AOI21_X1 U15740 ( .B1(n18337), .B2(n12647), .A(n17098), .ZN(n18323) );
  OAI21_X1 U15741 ( .B1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n12648), .A(
        n12647), .ZN(n18344) );
  INV_X1 U15742 ( .A(n18344), .ZN(n17320) );
  AOI21_X1 U15743 ( .B1(n13101), .B2(n18322), .A(n12648), .ZN(n18356) );
  INV_X1 U15744 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n18380) );
  INV_X1 U15745 ( .A(n12649), .ZN(n12651) );
  NOR2_X1 U15746 ( .A1(n18380), .A2(n12651), .ZN(n12650) );
  OAI21_X1 U15747 ( .B1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n12650), .A(
        n18322), .ZN(n18370) );
  INV_X1 U15748 ( .A(n18370), .ZN(n17331) );
  AOI21_X1 U15749 ( .B1(n18380), .B2(n12651), .A(n12650), .ZN(n18378) );
  NAND2_X1 U15750 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n9806), .ZN(
        n12654) );
  NOR2_X1 U15751 ( .A1(n18410), .A2(n12654), .ZN(n18366) );
  OAI21_X1 U15752 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n18366), .A(
        n12651), .ZN(n12652) );
  INV_X1 U15753 ( .A(n12652), .ZN(n18395) );
  INV_X1 U15754 ( .A(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n18414) );
  INV_X1 U15755 ( .A(n12654), .ZN(n12655) );
  NAND2_X1 U15756 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n12655), .ZN(
        n12653) );
  AOI21_X1 U15757 ( .B1(n18414), .B2(n12653), .A(n18366), .ZN(n18412) );
  INV_X1 U15758 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n18422) );
  AOI22_X1 U15759 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n12655), .B1(
        n12654), .B2(n18422), .ZN(n18425) );
  INV_X1 U15760 ( .A(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n18409) );
  INV_X1 U15761 ( .A(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n17415) );
  NAND2_X1 U15762 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18468), .ZN(
        n17420) );
  NOR2_X1 U15763 ( .A1(n17415), .A2(n17420), .ZN(n17406) );
  INV_X1 U15764 ( .A(n17406), .ZN(n18444) );
  NOR2_X1 U15765 ( .A1(n18447), .A2(n18444), .ZN(n12656) );
  INV_X1 U15766 ( .A(n12656), .ZN(n18407) );
  AOI21_X1 U15767 ( .B1(n18409), .B2(n18407), .A(n12655), .ZN(n18431) );
  INV_X1 U15768 ( .A(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n18451) );
  NAND2_X1 U15769 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n17406), .ZN(
        n12657) );
  AOI21_X1 U15770 ( .B1(n18451), .B2(n12657), .A(n12656), .ZN(n18449) );
  NOR2_X1 U15771 ( .A1(n17615), .A2(n18482), .ZN(n18481) );
  NAND2_X1 U15772 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n18481), .ZN(
        n17433) );
  NOR2_X1 U15773 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n17433), .ZN(
        n17419) );
  INV_X1 U15774 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n18459) );
  AOI22_X1 U15775 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n17406), .B1(
        n18444), .B2(n18459), .ZN(n18462) );
  NOR2_X1 U15776 ( .A1(n18449), .A2(n17389), .ZN(n17388) );
  NOR2_X1 U15777 ( .A1(n17388), .A2(n17576), .ZN(n17379) );
  NOR2_X1 U15778 ( .A1(n17378), .A2(n17576), .ZN(n17370) );
  NOR2_X1 U15779 ( .A1(n18395), .A2(n17351), .ZN(n17350) );
  NOR2_X1 U15780 ( .A1(n17350), .A2(n17576), .ZN(n17344) );
  NOR2_X1 U15781 ( .A1(n18356), .A2(n13099), .ZN(n13098) );
  NOR2_X1 U15782 ( .A1(n13098), .A2(n17576), .ZN(n17319) );
  NOR2_X1 U15783 ( .A1(n17320), .A2(n17319), .ZN(n17318) );
  NOR2_X1 U15784 ( .A1(n17318), .A2(n17576), .ZN(n17311) );
  NOR2_X1 U15785 ( .A1(n18323), .A2(n17311), .ZN(n17310) );
  NOR2_X1 U15786 ( .A1(n17310), .A2(n17576), .ZN(n17299) );
  NOR2_X1 U15787 ( .A1(n17298), .A2(n17576), .ZN(n17288) );
  XOR2_X1 U15788 ( .A(n17289), .B(n17288), .Z(n12794) );
  INV_X1 U15789 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n19660) );
  INV_X1 U15790 ( .A(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n17848) );
  INV_X1 U15791 ( .A(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n17982) );
  OAI22_X1 U15792 ( .A1(n17827), .A2(n17848), .B1(n17958), .B2(n17982), .ZN(
        n12671) );
  AOI22_X1 U15793 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n17948), .B1(
        n17971), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12669) );
  AND2_X2 U15794 ( .A1(n12677), .A2(n12664), .ZN(n12882) );
  AOI22_X1 U15795 ( .A1(n12882), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n9714), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12668) );
  NAND3_X1 U15796 ( .A1(n19666), .A2(n19674), .A3(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n12665) );
  AOI22_X1 U15797 ( .A1(n17864), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12840), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12667) );
  NAND3_X1 U15798 ( .A1(n12669), .A2(n12668), .A3(n12667), .ZN(n12670) );
  AOI211_X1 U15799 ( .C1(n17979), .C2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A(
        n12671), .B(n12670), .ZN(n12683) );
  INV_X1 U15800 ( .A(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n17969) );
  AOI22_X1 U15801 ( .A1(n17970), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n17972), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12673) );
  OAI21_X1 U15802 ( .B1(n17969), .B2(n17983), .A(n12673), .ZN(n12681) );
  NOR3_X1 U15803 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n19506), .A3(
        n19666), .ZN(n12831) );
  INV_X4 U15804 ( .A(n12726), .ZN(n17989) );
  AOI22_X1 U15805 ( .A1(n17989), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n17967), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12679) );
  NOR2_X4 U15806 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n12676), .ZN(
        n12846) );
  INV_X1 U15807 ( .A(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n19170) );
  NAND3_X1 U15808 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(n12677), .ZN(n17879) );
  NAND3_X1 U15809 ( .A1(n12679), .A2(n10203), .A3(n12678), .ZN(n12680) );
  AND2_X2 U15810 ( .A1(n12683), .A2(n12682), .ZN(n19040) );
  INV_X1 U15811 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n19577) );
  INV_X1 U15812 ( .A(P3_STATE_REG_1__SCAN_IN), .ZN(n19565) );
  OR2_X1 U15813 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n19565), .ZN(n19708) );
  INV_X2 U15814 ( .A(n19708), .ZN(n19710) );
  OAI211_X1 U15815 ( .C1(P3_STATE_REG_1__SCAN_IN), .C2(P3_STATE_REG_2__SCAN_IN), .A(n19577), .B(n19640), .ZN(n19698) );
  NAND2_X1 U15816 ( .A1(READY22_REG_SCAN_IN), .A2(READY2), .ZN(n19701) );
  INV_X1 U15817 ( .A(n19701), .ZN(n19696) );
  AOI211_X1 U15818 ( .C1(n19040), .C2(n19698), .A(P3_STATEBS16_REG_SCAN_IN), 
        .B(n19696), .ZN(n12783) );
  INV_X1 U15819 ( .A(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n17990) );
  AOI22_X1 U15820 ( .A1(n18002), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n9714), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12694) );
  INV_X1 U15821 ( .A(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n19075) );
  AOI22_X1 U15822 ( .A1(n17972), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17948), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12686) );
  AOI22_X1 U15823 ( .A1(n12839), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17970), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12685) );
  OAI211_X1 U15824 ( .C1(n17975), .C2(n19075), .A(n12686), .B(n12685), .ZN(
        n12692) );
  AOI22_X1 U15825 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n12882), .B1(
        P3_INSTQUEUE_REG_7__0__SCAN_IN), .B2(n17989), .ZN(n12690) );
  INV_X4 U15826 ( .A(n17827), .ZN(n17991) );
  AOI22_X1 U15827 ( .A1(n17991), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17971), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12689) );
  AOI22_X1 U15828 ( .A1(n17967), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n17864), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12688) );
  NAND2_X1 U15829 ( .A1(n12846), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n12687) );
  NAND4_X1 U15830 ( .A1(n12690), .A2(n12689), .A3(n12688), .A4(n12687), .ZN(
        n12691) );
  INV_X1 U15831 ( .A(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n17789) );
  AOI22_X1 U15832 ( .A1(n12846), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17971), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12704) );
  INV_X1 U15833 ( .A(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n17708) );
  AOI22_X1 U15834 ( .A1(n17972), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17948), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12696) );
  AOI22_X1 U15835 ( .A1(n17991), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12882), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12695) );
  OAI211_X1 U15836 ( .C1(n10201), .C2(n17708), .A(n12696), .B(n12695), .ZN(
        n12702) );
  AOI22_X1 U15837 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n17989), .B1(
        P3_INSTQUEUE_REG_2__5__SCAN_IN), .B2(n9714), .ZN(n12700) );
  AOI22_X1 U15838 ( .A1(P3_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n17970), .B1(
        n17954), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12699) );
  AOI22_X1 U15839 ( .A1(n12839), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n18002), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12698) );
  NAND2_X1 U15840 ( .A1(n12840), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n12697) );
  NAND4_X1 U15841 ( .A1(n12700), .A2(n12699), .A3(n12698), .A4(n12697), .ZN(
        n12701) );
  INV_X1 U15842 ( .A(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n17818) );
  AOI22_X1 U15843 ( .A1(n18002), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12899), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12715) );
  INV_X1 U15844 ( .A(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n17819) );
  AOI22_X1 U15845 ( .A1(n17989), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17967), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12707) );
  AOI22_X1 U15846 ( .A1(n17971), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n9714), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12706) );
  OAI211_X1 U15847 ( .C1(n10201), .C2(n17819), .A(n12707), .B(n12706), .ZN(
        n12713) );
  AOI22_X1 U15848 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n17954), .B1(
        n17972), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12711) );
  AOI22_X1 U15849 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n17991), .B1(
        n17970), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12710) );
  AOI22_X1 U15850 ( .A1(n12846), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17948), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12709) );
  NAND2_X1 U15851 ( .A1(n12840), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n12708) );
  NAND4_X1 U15852 ( .A1(n12711), .A2(n12710), .A3(n12709), .A4(n12708), .ZN(
        n12712) );
  INV_X1 U15853 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n18014) );
  AOI22_X1 U15854 ( .A1(n12846), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17864), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12725) );
  INV_X1 U15855 ( .A(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n17887) );
  AOI22_X1 U15856 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n12839), .B1(
        n12899), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12717) );
  AOI22_X1 U15857 ( .A1(n9740), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n9714), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12716) );
  OAI211_X1 U15858 ( .C1(n17887), .C2(n17995), .A(n12717), .B(n12716), .ZN(
        n12723) );
  AOI22_X1 U15859 ( .A1(n17972), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n17991), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12721) );
  AOI22_X1 U15860 ( .A1(n17989), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n17967), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12720) );
  AOI22_X1 U15861 ( .A1(n17954), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n17948), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12719) );
  NAND2_X1 U15862 ( .A1(n18002), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n12718) );
  NAND4_X1 U15863 ( .A1(n12721), .A2(n12720), .A3(n12719), .A4(n12718), .ZN(
        n12722) );
  NAND2_X1 U15864 ( .A1(n12759), .A2(n9754), .ZN(n12997) );
  INV_X1 U15865 ( .A(n12997), .ZN(n12754) );
  INV_X1 U15866 ( .A(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n17947) );
  AOI22_X1 U15867 ( .A1(n12882), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n9714), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12727) );
  OAI21_X1 U15868 ( .B1(n12726), .B2(n17947), .A(n12727), .ZN(n12736) );
  INV_X1 U15869 ( .A(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n17659) );
  AOI22_X1 U15870 ( .A1(n17972), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n17967), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12734) );
  INV_X1 U15871 ( .A(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n17957) );
  INV_X1 U15872 ( .A(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n17945) );
  OAI22_X1 U15873 ( .A1(n17995), .A2(n17957), .B1(n12838), .B2(n17945), .ZN(
        n12732) );
  AOI22_X1 U15874 ( .A1(n17970), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n17991), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12730) );
  AOI22_X1 U15875 ( .A1(n17954), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17948), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12729) );
  AOI22_X1 U15876 ( .A1(n17864), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12840), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12728) );
  NAND3_X1 U15877 ( .A1(n12730), .A2(n12729), .A3(n12728), .ZN(n12731) );
  AOI211_X1 U15878 ( .C1(n12846), .C2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A(
        n12732), .B(n12731), .ZN(n12733) );
  OAI211_X1 U15879 ( .C1(n17958), .C2(n17659), .A(n12734), .B(n12733), .ZN(
        n12735) );
  NAND2_X1 U15880 ( .A1(n19044), .A2(n12755), .ZN(n12956) );
  INV_X1 U15881 ( .A(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17781) );
  AOI22_X1 U15882 ( .A1(n17967), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n18002), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12746) );
  INV_X1 U15883 ( .A(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n17642) );
  AOI22_X1 U15884 ( .A1(n12839), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17948), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12738) );
  AOI22_X1 U15885 ( .A1(n17989), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n9740), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12737) );
  OAI211_X1 U15886 ( .C1(n10201), .C2(n17642), .A(n12738), .B(n12737), .ZN(
        n12744) );
  AOI22_X1 U15887 ( .A1(n17972), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n9714), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12742) );
  AOI22_X1 U15888 ( .A1(n17954), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17991), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12741) );
  AOI22_X1 U15889 ( .A1(n12840), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n12882), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12740) );
  NAND2_X1 U15890 ( .A1(n12846), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(
        n12739) );
  NAND4_X1 U15891 ( .A1(n12742), .A2(n12741), .A3(n12740), .A4(n12739), .ZN(
        n12743) );
  AOI211_X1 U15892 ( .C1(n17979), .C2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A(
        n12744), .B(n12743), .ZN(n12745) );
  INV_X1 U15893 ( .A(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n17811) );
  AOI22_X1 U15894 ( .A1(n18002), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17948), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12753) );
  INV_X1 U15895 ( .A(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n17923) );
  AOI22_X1 U15896 ( .A1(n17972), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n9714), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12747) );
  OAI21_X1 U15897 ( .B1(n17923), .B2(n12705), .A(n12747), .ZN(n12751) );
  INV_X1 U15898 ( .A(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n17918) );
  AOI22_X1 U15899 ( .A1(n12846), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17989), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12750) );
  INV_X1 U15900 ( .A(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n17915) );
  AOI22_X1 U15901 ( .A1(n17967), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n17971), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12749) );
  AOI22_X1 U15902 ( .A1(n17954), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17970), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12748) );
  NAND2_X1 U15903 ( .A1(n19061), .A2(n12945), .ZN(n19494) );
  NAND2_X1 U15904 ( .A1(n19056), .A2(n18053), .ZN(n12769) );
  NAND3_X1 U15905 ( .A1(n19044), .A2(n19494), .A3(n12769), .ZN(n12758) );
  NOR4_X1 U15906 ( .A1(n9752), .A2(n12945), .A3(n12759), .A4(n12946), .ZN(
        n12756) );
  NAND2_X1 U15907 ( .A1(n12756), .A2(n9754), .ZN(n12767) );
  NAND2_X1 U15908 ( .A1(n12760), .A2(n17263), .ZN(n14693) );
  OAI211_X1 U15909 ( .C1(n19068), .C2(n19516), .A(n19040), .B(n9752), .ZN(
        n12953) );
  INV_X1 U15910 ( .A(n12758), .ZN(n12765) );
  NOR3_X1 U15911 ( .A1(n12760), .A2(n12768), .A3(n12759), .ZN(n12764) );
  INV_X1 U15912 ( .A(n19516), .ZN(n16524) );
  NAND2_X1 U15913 ( .A1(n9754), .A2(n12946), .ZN(n12761) );
  NAND2_X1 U15914 ( .A1(n12945), .A2(n12761), .ZN(n12762) );
  AOI211_X2 U15915 ( .C1(n12765), .C2(n9751), .A(n12764), .B(n12763), .ZN(
        n12943) );
  OAI211_X1 U15916 ( .C1(n19048), .C2(n12766), .A(n12953), .B(n12943), .ZN(
        n12996) );
  INV_X1 U15917 ( .A(n12768), .ZN(n12770) );
  NAND2_X1 U15918 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n19660), .ZN(n19549) );
  INV_X1 U15919 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n19712) );
  NOR2_X1 U15920 ( .A1(n19549), .A2(n19712), .ZN(n19694) );
  NOR2_X1 U15921 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n12663), .ZN(
        n12948) );
  AOI22_X1 U15922 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n19522), .B1(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n19674), .ZN(n12950) );
  XNOR2_X1 U15923 ( .A(n12948), .B(n12950), .ZN(n12781) );
  AOI21_X1 U15924 ( .B1(n19522), .B2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n12771), .ZN(n12777) );
  OAI22_X1 U15925 ( .A1(n19666), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B1(
        n19527), .B2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n12776) );
  INV_X1 U15926 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n19531) );
  OR2_X1 U15927 ( .A1(n12776), .A2(n12777), .ZN(n12772) );
  OAI21_X1 U15928 ( .B1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n19666), .A(
        n12772), .ZN(n12773) );
  OAI22_X1 U15929 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n19531), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n12773), .ZN(n12778) );
  NOR2_X1 U15930 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n19531), .ZN(
        n12774) );
  NAND2_X1 U15931 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n12773), .ZN(
        n12779) );
  AOI22_X1 U15932 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n12778), .B1(
        n12774), .B2(n12779), .ZN(n12949) );
  NAND2_X1 U15933 ( .A1(n12777), .A2(n12776), .ZN(n12775) );
  OAI211_X1 U15934 ( .C1(n12777), .C2(n12776), .A(n12949), .B(n12775), .ZN(
        n12962) );
  AOI21_X1 U15935 ( .B1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n12779), .A(
        n12778), .ZN(n12780) );
  AOI21_X1 U15936 ( .B1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n19531), .A(
        n12780), .ZN(n12952) );
  OAI21_X1 U15937 ( .B1(n12781), .B2(n12962), .A(n12952), .ZN(n19479) );
  INV_X1 U15938 ( .A(n19479), .ZN(n12960) );
  NAND2_X1 U15939 ( .A1(n19694), .A2(n12960), .ZN(n18204) );
  AOI211_X4 U15940 ( .C1(P3_EBX_REG_31__SCAN_IN), .C2(n17101), .A(n12783), .B(
        n12784), .ZN(n17581) );
  NOR2_X1 U15941 ( .A1(P3_STATEBS16_REG_SCAN_IN), .A2(n19696), .ZN(n12782) );
  INV_X1 U15942 ( .A(P3_EBX_REG_31__SCAN_IN), .ZN(n17631) );
  NOR4_X4 U15943 ( .A1(n12782), .A2(n19040), .A3(n17631), .A4(n12784), .ZN(
        n17583) );
  NOR3_X1 U15944 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n17591) );
  INV_X1 U15945 ( .A(P3_EBX_REG_3__SCAN_IN), .ZN(n18026) );
  NAND2_X1 U15946 ( .A1(n17591), .A2(n18026), .ZN(n17582) );
  NOR2_X1 U15947 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n17582), .ZN(n17565) );
  INV_X1 U15948 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n18011) );
  NAND2_X1 U15949 ( .A1(n17565), .A2(n18011), .ZN(n17555) );
  NOR2_X1 U15950 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n17555), .ZN(n17540) );
  INV_X1 U15951 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n18012) );
  NAND2_X1 U15952 ( .A1(n17540), .A2(n18012), .ZN(n17528) );
  NOR2_X1 U15953 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n17528), .ZN(n17519) );
  INV_X1 U15954 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n17511) );
  NAND2_X1 U15955 ( .A1(n17519), .A2(n17511), .ZN(n17510) );
  NOR2_X1 U15956 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n17510), .ZN(n17495) );
  INV_X1 U15957 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n17490) );
  NAND2_X1 U15958 ( .A1(n17495), .A2(n17490), .ZN(n17482) );
  NOR2_X1 U15959 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n17482), .ZN(n17467) );
  INV_X1 U15960 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n17462) );
  NAND2_X1 U15961 ( .A1(n17467), .A2(n17462), .ZN(n17461) );
  NOR2_X1 U15962 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n17461), .ZN(n17444) );
  INV_X1 U15963 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n17437) );
  NAND2_X1 U15964 ( .A1(n17444), .A2(n17437), .ZN(n17436) );
  NOR2_X1 U15965 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n17436), .ZN(n17422) );
  INV_X1 U15966 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n17412) );
  NAND2_X1 U15967 ( .A1(n17422), .A2(n17412), .ZN(n17411) );
  NOR2_X1 U15968 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n17411), .ZN(n17398) );
  INV_X1 U15969 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n17392) );
  NAND2_X1 U15970 ( .A1(n17398), .A2(n17392), .ZN(n17390) );
  NOR2_X1 U15971 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n17390), .ZN(n17380) );
  INV_X1 U15972 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n17801) );
  NAND2_X1 U15973 ( .A1(n17380), .A2(n17801), .ZN(n17374) );
  NOR2_X1 U15974 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n17374), .ZN(n17362) );
  INV_X1 U15975 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n17736) );
  NAND2_X1 U15976 ( .A1(n17362), .A2(n17736), .ZN(n17357) );
  NOR2_X1 U15977 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n17357), .ZN(n17342) );
  INV_X1 U15978 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n17737) );
  NAND2_X1 U15979 ( .A1(n17342), .A2(n17737), .ZN(n17336) );
  NOR2_X1 U15980 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n17336), .ZN(n17326) );
  INV_X1 U15981 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n17325) );
  NAND2_X1 U15982 ( .A1(n17326), .A2(n17325), .ZN(n17324) );
  NOR2_X1 U15983 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n17324), .ZN(n17309) );
  INV_X1 U15984 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n17743) );
  NAND2_X1 U15985 ( .A1(n17309), .A2(n17743), .ZN(n12790) );
  NOR2_X1 U15986 ( .A1(n17618), .A2(n12790), .ZN(n17295) );
  OAI21_X1 U15987 ( .B1(n17581), .B2(n17295), .A(P3_EBX_REG_30__SCAN_IN), .ZN(
        n12792) );
  INV_X1 U15988 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n19628) );
  INV_X1 U15989 ( .A(n12783), .ZN(n19538) );
  INV_X1 U15990 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n19623) );
  INV_X1 U15991 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n19611) );
  INV_X1 U15992 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n19606) );
  INV_X1 U15993 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n19602) );
  INV_X1 U15994 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n19598) );
  INV_X1 U15995 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n19590) );
  INV_X1 U15996 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n19588) );
  INV_X1 U15997 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n19582) );
  NAND2_X1 U15998 ( .A1(P3_REIP_REG_2__SCAN_IN), .A2(P3_REIP_REG_1__SCAN_IN), 
        .ZN(n17601) );
  NOR2_X1 U15999 ( .A1(n19582), .A2(n17601), .ZN(n17548) );
  NAND3_X1 U16000 ( .A1(P3_REIP_REG_5__SCAN_IN), .A2(P3_REIP_REG_4__SCAN_IN), 
        .A3(n17548), .ZN(n17537) );
  NOR3_X1 U16001 ( .A1(n19590), .A2(n19588), .A3(n17537), .ZN(n17521) );
  NAND2_X1 U16002 ( .A1(P3_REIP_REG_8__SCAN_IN), .A2(n17521), .ZN(n17491) );
  NAND2_X1 U16003 ( .A1(P3_REIP_REG_10__SCAN_IN), .A2(P3_REIP_REG_9__SCAN_IN), 
        .ZN(n17500) );
  NOR3_X1 U16004 ( .A1(n19598), .A2(n17491), .A3(n17500), .ZN(n17470) );
  NAND2_X1 U16005 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n17470), .ZN(n17454) );
  NOR2_X1 U16006 ( .A1(n19602), .A2(n17454), .ZN(n17446) );
  NAND2_X1 U16007 ( .A1(P3_REIP_REG_14__SCAN_IN), .A2(n17446), .ZN(n17430) );
  NOR2_X1 U16008 ( .A1(n19606), .A2(n17430), .ZN(n17423) );
  NAND2_X1 U16009 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(n17423), .ZN(n17408) );
  NOR2_X1 U16010 ( .A1(n19611), .A2(n17408), .ZN(n17387) );
  NAND4_X1 U16011 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(n17387), .A3(
        P3_REIP_REG_19__SCAN_IN), .A4(P3_REIP_REG_18__SCAN_IN), .ZN(n17361) );
  NAND2_X1 U16012 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(P3_REIP_REG_21__SCAN_IN), 
        .ZN(n17349) );
  NOR3_X1 U16013 ( .A1(n19623), .A2(n17361), .A3(n17349), .ZN(n17341) );
  NAND2_X1 U16014 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n17341), .ZN(n12786) );
  NOR2_X1 U16015 ( .A1(n17609), .A2(n12786), .ZN(n17335) );
  NAND2_X1 U16016 ( .A1(P3_REIP_REG_25__SCAN_IN), .A2(n17335), .ZN(n13097) );
  NOR2_X1 U16017 ( .A1(n19628), .A2(n13097), .ZN(n17308) );
  NAND4_X1 U16018 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .A4(n17308), .ZN(n17286) );
  NOR2_X1 U16019 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n17286), .ZN(n17290) );
  NAND3_X1 U16020 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .ZN(n12788) );
  NAND2_X1 U16021 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n19712), .ZN(n19550) );
  INV_X1 U16022 ( .A(n17608), .ZN(n19555) );
  NOR2_X1 U16023 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n19713) );
  INV_X1 U16024 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n19542) );
  OAI211_X1 U16025 ( .C1(n19549), .C2(n19550), .A(n19555), .B(n19013), .ZN(
        n12785) );
  INV_X1 U16026 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n19626) );
  NOR3_X1 U16027 ( .A1(n17621), .A2(n12786), .A3(n19626), .ZN(n12787) );
  NOR2_X1 U16028 ( .A1(n17602), .A2(n17621), .ZN(n17617) );
  AOI21_X1 U16029 ( .B1(P3_REIP_REG_26__SCAN_IN), .B2(n12787), .A(n17617), 
        .ZN(n13096) );
  AOI21_X1 U16030 ( .B1(n17602), .B2(n12788), .A(n13096), .ZN(n17301) );
  INV_X1 U16031 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n19639) );
  INV_X1 U16032 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n17109) );
  OAI22_X1 U16033 ( .A1(n17301), .A2(n19639), .B1(n17109), .B2(n17586), .ZN(
        n12789) );
  NAND2_X1 U16034 ( .A1(n17583), .A2(n12790), .ZN(n17306) );
  NAND3_X1 U16035 ( .A1(n12792), .A2(n10222), .A3(n12791), .ZN(n12793) );
  NAND2_X1 U16036 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n13000) );
  INV_X1 U16037 ( .A(n13000), .ZN(n18800) );
  INV_X1 U16038 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n18040) );
  AOI22_X1 U16039 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n9748), .B1(
        n12831), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12800) );
  INV_X1 U16040 ( .A(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12796) );
  OAI22_X1 U16041 ( .A1(n19170), .A2(n12797), .B1(n17983), .B2(n12796), .ZN(
        n12798) );
  INV_X1 U16042 ( .A(n12798), .ZN(n12799) );
  OAI211_X1 U16043 ( .C1(n18040), .C2(n17995), .A(n12800), .B(n12799), .ZN(
        n12801) );
  AOI22_X1 U16044 ( .A1(n17970), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_13__1__SCAN_IN), .B2(n17971), .ZN(n12810) );
  INV_X1 U16045 ( .A(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12802) );
  INV_X1 U16046 ( .A(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n17851) );
  AND2_X1 U16047 ( .A1(n12805), .A2(n12804), .ZN(n12806) );
  OAI21_X1 U16048 ( .B1(n17975), .B2(n17851), .A(n12806), .ZN(n12807) );
  INV_X1 U16049 ( .A(n12807), .ZN(n12808) );
  INV_X1 U16050 ( .A(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n17976) );
  AOI22_X1 U16051 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n17948), .B1(
        n12830), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12812) );
  OAI21_X1 U16052 ( .B1(n17976), .B2(n12829), .A(n12812), .ZN(n12814) );
  INV_X1 U16053 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n19662) );
  NOR2_X1 U16054 ( .A1(n9895), .A2(n19662), .ZN(n12828) );
  XNOR2_X1 U16055 ( .A(n12847), .B(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18676) );
  AOI22_X1 U16056 ( .A1(n12839), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17972), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12818) );
  AOI22_X1 U16057 ( .A1(n17992), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12830), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12817) );
  AOI22_X1 U16058 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n12882), .B1(
        n17971), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12816) );
  NAND2_X1 U16059 ( .A1(n18002), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n12815) );
  NAND4_X1 U16060 ( .A1(n12818), .A2(n12817), .A3(n12816), .A4(n12815), .ZN(
        n12821) );
  AOI22_X1 U16061 ( .A1(n17967), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n17948), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12819) );
  INV_X1 U16062 ( .A(n12819), .ZN(n12820) );
  AOI22_X1 U16063 ( .A1(n17989), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n9714), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12826) );
  AOI22_X1 U16064 ( .A1(n17864), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12840), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12825) );
  INV_X1 U16065 ( .A(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n15307) );
  INV_X1 U16066 ( .A(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n17863) );
  OAI22_X1 U16067 ( .A1(n15307), .A2(n12866), .B1(n17995), .B2(n17863), .ZN(
        n12822) );
  INV_X1 U16068 ( .A(n12822), .ZN(n12824) );
  NAND2_X1 U16069 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n18683), .ZN(
        n18682) );
  NOR2_X1 U16070 ( .A1(n12828), .A2(n18675), .ZN(n18664) );
  INV_X1 U16071 ( .A(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n17842) );
  AOI22_X1 U16072 ( .A1(n12831), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12830), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12832) );
  OAI21_X1 U16073 ( .B1(n12829), .B2(n17842), .A(n12832), .ZN(n12837) );
  AOI22_X1 U16074 ( .A1(n9748), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n18002), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12836) );
  INV_X1 U16075 ( .A(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n19081) );
  AOI21_X1 U16076 ( .B1(n17972), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A(
        n12834), .ZN(n12835) );
  INV_X1 U16077 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n18038) );
  INV_X1 U16078 ( .A(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n17837) );
  OAI22_X1 U16079 ( .A1(n17995), .A2(n18038), .B1(n17966), .B2(n17837), .ZN(
        n12845) );
  AOI22_X1 U16080 ( .A1(n12839), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n17971), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12843) );
  AOI22_X1 U16081 ( .A1(n17992), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12882), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12842) );
  AOI22_X1 U16082 ( .A1(n17864), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12840), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12841) );
  NAND3_X1 U16083 ( .A1(n12843), .A2(n12842), .A3(n12841), .ZN(n12844) );
  NAND2_X1 U16084 ( .A1(n12847), .A2(n18191), .ZN(n12848) );
  INV_X1 U16085 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18999) );
  XNOR2_X1 U16086 ( .A(n12849), .B(n18999), .ZN(n18663) );
  NOR2_X1 U16087 ( .A1(n18999), .A2(n12849), .ZN(n12850) );
  INV_X1 U16088 ( .A(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n17930) );
  AOI22_X1 U16089 ( .A1(n12846), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17971), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12860) );
  INV_X1 U16090 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n18031) );
  AOI22_X1 U16091 ( .A1(n17970), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n17948), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12852) );
  AOI22_X1 U16092 ( .A1(n17954), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17972), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12851) );
  OAI211_X1 U16093 ( .C1(n17995), .C2(n18031), .A(n12852), .B(n12851), .ZN(
        n12858) );
  AOI22_X1 U16094 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n17967), .B1(
        n12839), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12856) );
  AOI22_X1 U16095 ( .A1(n12882), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n9714), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12855) );
  AOI22_X1 U16096 ( .A1(n17991), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n18002), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12854) );
  NAND2_X1 U16097 ( .A1(n17864), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n12853) );
  NAND4_X1 U16098 ( .A1(n12856), .A2(n12855), .A3(n12854), .A4(n12853), .ZN(
        n12857) );
  AOI211_X1 U16099 ( .C1(n12840), .C2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A(
        n12858), .B(n12857), .ZN(n12859) );
  OAI211_X1 U16100 ( .C1(n17930), .C2(n12726), .A(n12860), .B(n12859), .ZN(
        n12865) );
  INV_X1 U16101 ( .A(n12865), .ZN(n18185) );
  XNOR2_X1 U16102 ( .A(n18185), .B(n12864), .ZN(n12861) );
  XNOR2_X1 U16103 ( .A(n12862), .B(n12861), .ZN(n18652) );
  INV_X1 U16104 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n18976) );
  INV_X1 U16105 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n18967) );
  NAND2_X1 U16106 ( .A1(n12974), .A2(n12865), .ZN(n12894) );
  INV_X1 U16107 ( .A(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n17645) );
  AOI22_X1 U16108 ( .A1(n12840), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n12899), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12874) );
  OAI22_X1 U16109 ( .A1(n17923), .A2(n12867), .B1(n17811), .B2(n12726), .ZN(
        n12872) );
  AOI22_X1 U16110 ( .A1(n17991), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17948), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12870) );
  AOI22_X1 U16111 ( .A1(n12839), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n9748), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12869) );
  AOI22_X1 U16112 ( .A1(n17979), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n17864), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12868) );
  NAND3_X1 U16113 ( .A1(n12870), .A2(n12869), .A3(n12868), .ZN(n12871) );
  OAI211_X1 U16114 ( .C1(n17958), .C2(n17645), .A(n12874), .B(n12873), .ZN(
        n12875) );
  AOI22_X1 U16115 ( .A1(n17972), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n9714), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12876) );
  OAI21_X1 U16116 ( .B1(n17918), .B2(n17913), .A(n12876), .ZN(n12878) );
  INV_X2 U16117 ( .A(n17983), .ZN(n17954) );
  INV_X1 U16118 ( .A(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12893) );
  AOI22_X1 U16119 ( .A1(n17967), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n9714), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12892) );
  INV_X1 U16120 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n18021) );
  AOI22_X1 U16121 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n12882), .B1(
        n17991), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12884) );
  AOI22_X1 U16122 ( .A1(n17972), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17948), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12883) );
  OAI211_X1 U16123 ( .C1(n18021), .C2(n17995), .A(n12884), .B(n12883), .ZN(
        n12890) );
  AOI22_X1 U16124 ( .A1(n12839), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17971), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12888) );
  AOI22_X1 U16125 ( .A1(n17970), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n17989), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12887) );
  AOI22_X1 U16126 ( .A1(n17954), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n18002), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12886) );
  NAND2_X1 U16127 ( .A1(n17864), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n12885) );
  NAND4_X1 U16128 ( .A1(n12888), .A2(n12887), .A3(n12886), .A4(n12885), .ZN(
        n12889) );
  AOI211_X1 U16129 ( .C1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .C2(n12840), .A(
        n12890), .B(n12889), .ZN(n12891) );
  OAI211_X1 U16130 ( .C1(n12867), .C2(n12893), .A(n12892), .B(n12891), .ZN(
        n12969) );
  INV_X1 U16131 ( .A(n12969), .ZN(n18178) );
  XOR2_X1 U16132 ( .A(n18178), .B(n12909), .Z(n12895) );
  INV_X1 U16133 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n18629) );
  NOR2_X1 U16134 ( .A1(n12896), .A2(n12895), .ZN(n12897) );
  NOR2_X1 U16135 ( .A1(n18627), .A2(n12897), .ZN(n18614) );
  INV_X1 U16136 ( .A(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n17894) );
  AOI22_X1 U16137 ( .A1(n17972), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n9740), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12898) );
  OAI21_X1 U16138 ( .B1(n17879), .B2(n17894), .A(n12898), .ZN(n12908) );
  INV_X1 U16139 ( .A(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n17893) );
  AOI22_X1 U16140 ( .A1(n17970), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n12899), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12906) );
  INV_X1 U16141 ( .A(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n17776) );
  AOI22_X1 U16142 ( .A1(n12846), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n9714), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12900) );
  OAI21_X1 U16143 ( .B1(n17975), .B2(n17776), .A(n12900), .ZN(n12904) );
  AOI22_X1 U16144 ( .A1(n17967), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17948), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12902) );
  AOI22_X1 U16145 ( .A1(n17989), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17991), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12901) );
  OAI211_X1 U16146 ( .C1(n17995), .C2(n17781), .A(n12902), .B(n12901), .ZN(
        n12903) );
  AOI211_X1 U16147 ( .C1(n17864), .C2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A(
        n12904), .B(n12903), .ZN(n12905) );
  OAI211_X1 U16148 ( .C1(n17958), .C2(n17893), .A(n12906), .B(n12905), .ZN(
        n12907) );
  NAND2_X1 U16149 ( .A1(n12909), .A2(n12969), .ZN(n12912) );
  NOR2_X1 U16150 ( .A1(n18175), .A2(n12912), .ZN(n12923) );
  INV_X1 U16151 ( .A(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n17720) );
  AOI22_X1 U16152 ( .A1(n17954), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n17989), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12922) );
  AOI22_X1 U16153 ( .A1(n12899), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n9714), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12914) );
  AOI22_X1 U16154 ( .A1(n17970), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n17971), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12913) );
  OAI211_X1 U16155 ( .C1(n17995), .C2(n18014), .A(n12914), .B(n12913), .ZN(
        n12920) );
  AOI22_X1 U16156 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n12839), .B1(
        n17991), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12918) );
  AOI22_X1 U16157 ( .A1(n17967), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n17948), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12917) );
  AOI22_X1 U16158 ( .A1(n17972), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n12846), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12916) );
  NAND2_X1 U16159 ( .A1(n17864), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n12915) );
  NAND4_X1 U16160 ( .A1(n12918), .A2(n12917), .A3(n12916), .A4(n12915), .ZN(
        n12919) );
  AOI211_X1 U16161 ( .C1(n12840), .C2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A(
        n12920), .B(n12919), .ZN(n12921) );
  OAI21_X1 U16162 ( .B1(n12923), .B2(n17103), .A(n12931), .ZN(n12924) );
  INV_X1 U16163 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n18946) );
  INV_X1 U16164 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n18932) );
  NOR2_X2 U16165 ( .A1(n12927), .A2(n18932), .ZN(n17112) );
  INV_X1 U16166 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n18919) );
  INV_X1 U16167 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18906) );
  NOR2_X1 U16168 ( .A1(n18919), .A2(n18906), .ZN(n18895) );
  NAND2_X1 U16169 ( .A1(n18895), .A2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n18879) );
  INV_X1 U16170 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n18880) );
  NOR2_X1 U16171 ( .A1(n18879), .A2(n18880), .ZN(n18872) );
  NAND3_X1 U16172 ( .A1(n18872), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n18821) );
  INV_X1 U16173 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n18819) );
  NOR2_X1 U16174 ( .A1(n18821), .A2(n18819), .ZN(n18816) );
  NAND2_X1 U16175 ( .A1(n12927), .A2(n18932), .ZN(n18590) );
  OR2_X1 U16176 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18520) );
  INV_X1 U16177 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n18855) );
  NAND2_X1 U16178 ( .A1(n18855), .A2(n18819), .ZN(n18836) );
  INV_X1 U16179 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n18829) );
  NAND2_X1 U16180 ( .A1(n12930), .A2(n18479), .ZN(n18474) );
  INV_X1 U16181 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n18758) );
  INV_X1 U16182 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n18767) );
  INV_X1 U16183 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n18787) );
  INV_X1 U16184 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n18435) );
  NOR2_X1 U16185 ( .A1(n18787), .A2(n18435), .ZN(n18771) );
  NAND2_X1 U16186 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n18771), .ZN(
        n18759) );
  OR2_X1 U16187 ( .A1(n18767), .A2(n18759), .ZN(n18749) );
  NOR2_X1 U16188 ( .A1(n18758), .A2(n18749), .ZN(n17164) );
  NAND2_X1 U16189 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n17164), .ZN(
        n18705) );
  NAND2_X1 U16190 ( .A1(n18463), .A2(n18787), .ZN(n12932) );
  NOR2_X1 U16191 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n12932), .ZN(
        n18419) );
  INV_X1 U16192 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n18768) );
  NAND2_X1 U16193 ( .A1(n18419), .A2(n18768), .ZN(n18405) );
  NOR3_X1 U16194 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(n18405), .ZN(n12933) );
  NOR3_X1 U16195 ( .A1(n18465), .A2(n18384), .A3(n18705), .ZN(n12937) );
  INV_X1 U16196 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n18721) );
  NAND2_X1 U16197 ( .A1(n12931), .A2(n18374), .ZN(n12935) );
  OAI211_X1 U16198 ( .C1(n12937), .C2(n18721), .A(n12935), .B(n12934), .ZN(
        n18354) );
  INV_X1 U16199 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n12936) );
  NOR2_X1 U16200 ( .A1(n12937), .A2(n12931), .ZN(n18373) );
  INV_X1 U16201 ( .A(n18373), .ZN(n12939) );
  NAND2_X1 U16202 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n12999) );
  NAND2_X1 U16203 ( .A1(n18509), .A2(n12999), .ZN(n12938) );
  INV_X1 U16204 ( .A(n17151), .ZN(n12941) );
  INV_X1 U16205 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n18328) );
  NAND2_X1 U16206 ( .A1(n17158), .A2(n18328), .ZN(n12940) );
  NOR2_X1 U16207 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n12931), .ZN(
        n17160) );
  INV_X1 U16208 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n17128) );
  XNOR2_X1 U16209 ( .A(n12942), .B(n17128), .ZN(n17131) );
  INV_X1 U16210 ( .A(n12943), .ZN(n12944) );
  NAND2_X1 U16211 ( .A1(n19044), .A2(n17101), .ZN(n12955) );
  NOR2_X1 U16212 ( .A1(n19061), .A2(n12955), .ZN(n12963) );
  INV_X1 U16213 ( .A(n12945), .ZN(n19052) );
  OAI21_X1 U16214 ( .B1(n12947), .B2(n12946), .A(n19052), .ZN(n12958) );
  AOI21_X1 U16215 ( .B1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n12663), .A(
        n12948), .ZN(n12959) );
  NAND3_X1 U16216 ( .A1(n12950), .A2(n12949), .A3(n12959), .ZN(n12951) );
  NAND3_X1 U16217 ( .A1(n12952), .A2(n12962), .A3(n12951), .ZN(n17096) );
  OAI21_X1 U16218 ( .B1(n17263), .B2(n12954), .A(n12953), .ZN(n14690) );
  NOR2_X1 U16219 ( .A1(n19696), .A2(n19479), .ZN(n14694) );
  OAI211_X1 U16220 ( .C1(n19044), .C2(n17101), .A(n12955), .B(n19698), .ZN(
        n17268) );
  AND3_X1 U16221 ( .A1(n14694), .A2(n12956), .A3(n17268), .ZN(n12957) );
  AOI211_X1 U16222 ( .C1(n12958), .C2(n19484), .A(n14690), .B(n12957), .ZN(
        n12965) );
  INV_X1 U16223 ( .A(n12959), .ZN(n12961) );
  OAI21_X1 U16224 ( .B1(n12962), .B2(n12961), .A(n12960), .ZN(n19480) );
  INV_X1 U16225 ( .A(n12963), .ZN(n12964) );
  INV_X1 U16226 ( .A(n19694), .ZN(n19546) );
  AOI221_X4 U16227 ( .B1(n12965), .B2(n19480), .C1(n12965), .C2(n12964), .A(
        n19546), .ZN(n18995) );
  NAND2_X1 U16228 ( .A1(n17131), .A2(n18926), .ZN(n13013) );
  NAND2_X1 U16229 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n17152) );
  NOR2_X1 U16230 ( .A1(n17152), .A2(n17128), .ZN(n17138) );
  INV_X1 U16231 ( .A(n17138), .ZN(n16509) );
  INV_X1 U16232 ( .A(n12999), .ZN(n18693) );
  NAND3_X1 U16233 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n18693), .A3(
        n18735), .ZN(n17123) );
  INV_X1 U16234 ( .A(n17149), .ZN(n19481) );
  INV_X1 U16235 ( .A(n17103), .ZN(n18171) );
  NAND2_X1 U16236 ( .A1(n19481), .A2(n18171), .ZN(n18871) );
  NOR2_X1 U16237 ( .A1(n19014), .A2(n18871), .ZN(n18862) );
  INV_X1 U16238 ( .A(n18862), .ZN(n18922) );
  INV_X1 U16239 ( .A(n18821), .ZN(n18492) );
  NOR2_X1 U16240 ( .A1(n18185), .A2(n12973), .ZN(n12981) );
  NAND2_X1 U16241 ( .A1(n12981), .A2(n12980), .ZN(n12970) );
  NOR2_X1 U16242 ( .A1(n18178), .A2(n12970), .ZN(n12968) );
  NAND2_X1 U16243 ( .A1(n12968), .A2(n12967), .ZN(n12966) );
  NOR2_X1 U16244 ( .A1(n18171), .A2(n12966), .ZN(n12992) );
  XNOR2_X1 U16245 ( .A(n12966), .B(n17103), .ZN(n18605) );
  XOR2_X1 U16246 ( .A(n12968), .B(n12967), .Z(n12985) );
  XNOR2_X1 U16247 ( .A(n12970), .B(n12969), .ZN(n12971) );
  NAND2_X1 U16248 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n12971), .ZN(
        n12984) );
  XNOR2_X1 U16249 ( .A(n18629), .B(n12971), .ZN(n18626) );
  XOR2_X1 U16250 ( .A(n12973), .B(n18185), .Z(n12972) );
  NAND2_X1 U16251 ( .A1(n12972), .A2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12979) );
  XNOR2_X1 U16252 ( .A(n18976), .B(n12972), .ZN(n18655) );
  AOI21_X1 U16253 ( .B1(n18683), .B2(n12974), .A(n12973), .ZN(n12977) );
  OR2_X1 U16254 ( .A1(n18999), .A2(n12977), .ZN(n12978) );
  AOI21_X1 U16255 ( .B1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n9895), .A(
        n18683), .ZN(n12976) );
  INV_X1 U16256 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n19677) );
  NOR2_X1 U16257 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n9895), .ZN(
        n12975) );
  AOI221_X1 U16258 ( .B1(n18683), .B2(n9895), .C1(n12976), .C2(n19677), .A(
        n12975), .ZN(n18667) );
  XNOR2_X1 U16259 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n12977), .ZN(
        n18666) );
  NAND2_X1 U16260 ( .A1(n18667), .A2(n18666), .ZN(n18665) );
  NAND2_X1 U16261 ( .A1(n12978), .A2(n18665), .ZN(n18654) );
  NAND2_X1 U16262 ( .A1(n18655), .A2(n18654), .ZN(n18653) );
  NAND2_X1 U16263 ( .A1(n12979), .A2(n18653), .ZN(n12982) );
  NAND2_X1 U16264 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n12982), .ZN(
        n12983) );
  XOR2_X1 U16265 ( .A(n12981), .B(n12980), .Z(n18640) );
  XOR2_X1 U16266 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B(n12982), .Z(
        n18639) );
  NAND2_X1 U16267 ( .A1(n18640), .A2(n18639), .ZN(n18638) );
  NAND2_X1 U16268 ( .A1(n12983), .A2(n18638), .ZN(n18625) );
  NAND2_X1 U16269 ( .A1(n18626), .A2(n18625), .ZN(n18624) );
  NAND2_X1 U16270 ( .A1(n12984), .A2(n18624), .ZN(n12986) );
  NAND2_X1 U16271 ( .A1(n12985), .A2(n12986), .ZN(n12987) );
  XOR2_X1 U16272 ( .A(n12986), .B(n12985), .Z(n18617) );
  NAND2_X1 U16273 ( .A1(n18617), .A2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n18616) );
  NAND2_X1 U16274 ( .A1(n12992), .A2(n12989), .ZN(n12993) );
  INV_X1 U16275 ( .A(n12989), .ZN(n12991) );
  NAND2_X1 U16276 ( .A1(n18605), .A2(n18606), .ZN(n18604) );
  NAND2_X1 U16277 ( .A1(n12992), .A2(n12991), .ZN(n12990) );
  OAI211_X1 U16278 ( .C1(n12992), .C2(n12991), .A(n18604), .B(n12990), .ZN(
        n18593) );
  NAND2_X1 U16279 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n18593), .ZN(
        n18592) );
  NOR2_X1 U16280 ( .A1(n13000), .A2(n18705), .ZN(n18383) );
  INV_X1 U16281 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n18730) );
  NOR2_X2 U16282 ( .A1(n12994), .A2(n19505), .ZN(n19517) );
  NAND2_X1 U16283 ( .A1(n17101), .A2(n9752), .ZN(n16456) );
  NAND2_X1 U16284 ( .A1(n16521), .A2(n16456), .ZN(n19711) );
  NOR2_X1 U16285 ( .A1(n19040), .A2(n19505), .ZN(n12998) );
  NOR2_X1 U16286 ( .A1(n19483), .A2(n19014), .ZN(n18832) );
  OAI22_X1 U16287 ( .A1(n17124), .A2(n18922), .B1(n17126), .B2(n19017), .ZN(
        n16512) );
  INV_X2 U16288 ( .A(n19013), .ZN(n18948) );
  NAND2_X1 U16289 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n18716) );
  NOR2_X1 U16290 ( .A1(n12999), .A2(n18716), .ZN(n17113) );
  INV_X1 U16291 ( .A(n17164), .ZN(n18390) );
  INV_X1 U16292 ( .A(n18816), .ZN(n18811) );
  NOR2_X1 U16293 ( .A1(n13000), .A2(n18811), .ZN(n18456) );
  INV_X1 U16294 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n18950) );
  NOR2_X1 U16295 ( .A1(n18946), .A2(n18950), .ZN(n18933) );
  NAND2_X1 U16296 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n18933), .ZN(
        n13001) );
  NOR3_X1 U16297 ( .A1(n18629), .A2(n18967), .A3(n18976), .ZN(n18795) );
  OAI21_X1 U16298 ( .B1(n19677), .B2(n19662), .A(n18999), .ZN(n18986) );
  NAND2_X1 U16299 ( .A1(n18795), .A2(n18986), .ZN(n18930) );
  NOR2_X1 U16300 ( .A1(n13001), .A2(n18930), .ZN(n18867) );
  NAND2_X1 U16301 ( .A1(n18456), .A2(n18867), .ZN(n18802) );
  NOR2_X1 U16302 ( .A1(n18390), .A2(n18802), .ZN(n18714) );
  AOI21_X1 U16303 ( .B1(n17113), .B2(n18714), .A(n19509), .ZN(n18698) );
  NAND2_X1 U16304 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18964) );
  INV_X1 U16305 ( .A(n18964), .ZN(n18793) );
  AND2_X1 U16306 ( .A1(n18793), .A2(n18795), .ZN(n18927) );
  INV_X1 U16307 ( .A(n13001), .ZN(n18796) );
  NAND2_X1 U16308 ( .A1(n18927), .A2(n18796), .ZN(n18849) );
  NAND2_X1 U16309 ( .A1(n17164), .A2(n18456), .ZN(n18393) );
  NOR2_X1 U16310 ( .A1(n18849), .A2(n18393), .ZN(n18690) );
  INV_X1 U16311 ( .A(n19517), .ZN(n19499) );
  NOR2_X1 U16312 ( .A1(n19499), .A2(n19515), .ZN(n18928) );
  AOI21_X1 U16313 ( .B1(n18690), .B2(n17113), .A(n18928), .ZN(n13003) );
  AOI21_X1 U16314 ( .B1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A(n18914), .ZN(n13002) );
  NOR4_X1 U16315 ( .A1(n18698), .A2(n13003), .A3(n19014), .A4(n13002), .ZN(
        n16511) );
  INV_X1 U16316 ( .A(n16511), .ZN(n13004) );
  AOI21_X1 U16317 ( .B1(n18873), .B2(n10095), .A(n13004), .ZN(n17154) );
  INV_X1 U16318 ( .A(n18931), .ZN(n18824) );
  NAND2_X1 U16319 ( .A1(n18995), .A2(n18824), .ZN(n19001) );
  OAI22_X1 U16320 ( .A1(n18948), .A2(n17154), .B1(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n19001), .ZN(n13005) );
  OAI21_X1 U16321 ( .B1(n16512), .B2(n13005), .A(
        P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n13011) );
  INV_X1 U16322 ( .A(n17123), .ZN(n18694) );
  INV_X1 U16323 ( .A(n18849), .ZN(n18820) );
  OAI21_X1 U16324 ( .B1(n18914), .B2(n19677), .A(n19517), .ZN(n18989) );
  NAND3_X1 U16325 ( .A1(n18820), .A2(n18456), .A3(n18989), .ZN(n13006) );
  OAI21_X1 U16326 ( .B1(n18802), .B2(n19509), .A(n13006), .ZN(n17161) );
  NAND2_X1 U16327 ( .A1(n17164), .A2(n17161), .ZN(n18713) );
  NAND2_X1 U16328 ( .A1(n18995), .A2(n17113), .ZN(n17165) );
  NOR2_X1 U16329 ( .A1(n18713), .A2(n17165), .ZN(n17137) );
  AOI21_X1 U16330 ( .B1(n18862), .B2(n18694), .A(n17137), .ZN(n13007) );
  OAI21_X1 U16331 ( .B1(n18327), .B2(n19017), .A(n13007), .ZN(n16510) );
  NAND2_X1 U16332 ( .A1(n17128), .A2(n16510), .ZN(n13008) );
  OAI21_X1 U16333 ( .B1(n13008), .B2(n17152), .A(n17134), .ZN(n13009) );
  INV_X1 U16334 ( .A(n13015), .ZN(n13018) );
  INV_X1 U16335 ( .A(n13016), .ZN(n13017) );
  NAND2_X1 U16336 ( .A1(n13018), .A2(n13017), .ZN(n13019) );
  NAND2_X1 U16337 ( .A1(n13014), .A2(n13019), .ZN(n14731) );
  MUX2_X1 U16338 ( .A(n13020), .B(n16645), .S(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .Z(n13022) );
  NAND2_X1 U16339 ( .A1(n13022), .A2(n13021), .ZN(n13023) );
  NAND2_X1 U16340 ( .A1(n16782), .A2(P1_REIP_REG_28__SCAN_IN), .ZN(n15688) );
  OAI21_X1 U16341 ( .B1(n16670), .B2(n13024), .A(n15688), .ZN(n13025) );
  INV_X1 U16342 ( .A(n13029), .ZN(n13031) );
  NAND2_X1 U16343 ( .A1(n13031), .A2(n13030), .ZN(n13032) );
  NAND2_X1 U16344 ( .A1(n13033), .A2(n13032), .ZN(n16880) );
  NOR2_X1 U16345 ( .A1(n16880), .A2(n11790), .ZN(n14799) );
  XNOR2_X1 U16346 ( .A(n14801), .B(n10829), .ZN(n14791) );
  INV_X1 U16347 ( .A(n17071), .ZN(n20059) );
  NAND2_X1 U16348 ( .A1(n14791), .A2(n20059), .ZN(n13046) );
  NOR2_X1 U16349 ( .A1(n9790), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n13035) );
  XNOR2_X1 U16350 ( .A(n13036), .B(n13037), .ZN(n15909) );
  INV_X1 U16351 ( .A(n15909), .ZN(n16882) );
  OAI21_X1 U16352 ( .B1(n13038), .B2(n13040), .A(n13039), .ZN(n16888) );
  NAND2_X1 U16353 ( .A1(n14806), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n13041) );
  NAND2_X1 U16354 ( .A1(n19905), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n14792) );
  OAI211_X1 U16355 ( .C1(n17048), .C2(n16888), .A(n13041), .B(n14792), .ZN(
        n13042) );
  NOR2_X1 U16356 ( .A1(n14812), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14807) );
  AOI211_X1 U16357 ( .C1(n17074), .C2(n16882), .A(n13042), .B(n14807), .ZN(
        n13043) );
  INV_X1 U16358 ( .A(n13044), .ZN(n13045) );
  NAND2_X1 U16359 ( .A1(n13046), .A2(n13045), .ZN(P2_U3019) );
  NAND2_X1 U16360 ( .A1(n13314), .A2(n13303), .ZN(n13285) );
  INV_X1 U16361 ( .A(n13392), .ZN(n14873) );
  AND3_X1 U16362 ( .A1(n11129), .A2(n14873), .A3(n13049), .ZN(n13050) );
  AND2_X1 U16363 ( .A1(n13051), .A2(n13050), .ZN(n13386) );
  NAND2_X1 U16364 ( .A1(n13386), .A2(n13275), .ZN(n13052) );
  NAND2_X1 U16365 ( .A1(n13285), .A2(n13052), .ZN(n13053) );
  AND2_X2 U16366 ( .A1(n13053), .A2(n13289), .ZN(n16644) );
  AND2_X1 U16367 ( .A1(n16644), .A2(n13392), .ZN(n15545) );
  INV_X2 U16368 ( .A(n15545), .ZN(n16640) );
  NAND2_X1 U16369 ( .A1(n15612), .A2(n15545), .ZN(n13057) );
  NAND2_X2 U16370 ( .A1(n16644), .A2(n14873), .ZN(n15543) );
  INV_X1 U16371 ( .A(P1_EBX_REG_30__SCAN_IN), .ZN(n13054) );
  INV_X1 U16372 ( .A(n13055), .ZN(n13056) );
  NAND2_X1 U16373 ( .A1(n13059), .A2(n13058), .ZN(n13062) );
  INV_X1 U16374 ( .A(n13063), .ZN(n14815) );
  NAND2_X1 U16375 ( .A1(n12130), .A2(n13064), .ZN(n13065) );
  INV_X1 U16376 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n21251) );
  NOR2_X1 U16377 ( .A1(n16823), .A2(n21251), .ZN(n14736) );
  NOR3_X1 U16378 ( .A1(n15689), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n9914), .ZN(n13066) );
  AOI211_X1 U16379 ( .C1(n15469), .C2(n16809), .A(n14736), .B(n13066), .ZN(
        n13070) );
  OAI21_X1 U16380 ( .B1(n9785), .B2(n16792), .A(n13071), .ZN(P1_U3002) );
  NOR2_X1 U16381 ( .A1(P1_ADDRESS_REG_8__SCAN_IN), .A2(
        P1_ADDRESS_REG_24__SCAN_IN), .ZN(n15208) );
  NOR3_X1 U16382 ( .A1(P1_ADDRESS_REG_2__SCAN_IN), .A2(
        P1_ADDRESS_REG_1__SCAN_IN), .A3(P1_ADDRESS_REG_0__SCAN_IN), .ZN(n13074) );
  NOR4_X1 U16383 ( .A1(P1_ADDRESS_REG_25__SCAN_IN), .A2(
        P1_ADDRESS_REG_23__SCAN_IN), .A3(P1_ADDRESS_REG_22__SCAN_IN), .A4(
        P1_ADDRESS_REG_21__SCAN_IN), .ZN(n13073) );
  NOR4_X1 U16384 ( .A1(P1_ADDRESS_REG_5__SCAN_IN), .A2(
        P1_ADDRESS_REG_28__SCAN_IN), .A3(P1_ADDRESS_REG_27__SCAN_IN), .A4(
        P1_ADDRESS_REG_26__SCAN_IN), .ZN(n13072) );
  AND4_X1 U16385 ( .A1(n15208), .A2(n13074), .A3(n13073), .A4(n13072), .ZN(
        n13080) );
  NOR4_X1 U16386 ( .A1(P1_ADDRESS_REG_16__SCAN_IN), .A2(
        P1_ADDRESS_REG_15__SCAN_IN), .A3(P1_ADDRESS_REG_14__SCAN_IN), .A4(
        P1_ADDRESS_REG_13__SCAN_IN), .ZN(n13078) );
  NOR4_X1 U16387 ( .A1(P1_ADDRESS_REG_20__SCAN_IN), .A2(
        P1_ADDRESS_REG_19__SCAN_IN), .A3(P1_ADDRESS_REG_18__SCAN_IN), .A4(
        P1_ADDRESS_REG_17__SCAN_IN), .ZN(n13077) );
  NOR4_X1 U16388 ( .A1(P1_ADDRESS_REG_7__SCAN_IN), .A2(
        P1_ADDRESS_REG_6__SCAN_IN), .A3(P1_ADDRESS_REG_4__SCAN_IN), .A4(
        P1_ADDRESS_REG_3__SCAN_IN), .ZN(n13076) );
  NOR4_X1 U16389 ( .A1(P1_ADDRESS_REG_12__SCAN_IN), .A2(
        P1_ADDRESS_REG_11__SCAN_IN), .A3(P1_ADDRESS_REG_10__SCAN_IN), .A4(
        P1_ADDRESS_REG_9__SCAN_IN), .ZN(n13075) );
  AND4_X1 U16390 ( .A1(n13078), .A2(n13077), .A3(n13076), .A4(n13075), .ZN(
        n13079) );
  NAND2_X1 U16391 ( .A1(n13080), .A2(n13079), .ZN(n13081) );
  INV_X1 U16392 ( .A(P1_BE_N_REG_3__SCAN_IN), .ZN(n21256) );
  INV_X1 U16393 ( .A(P1_D_C_N_REG_SCAN_IN), .ZN(n15321) );
  AND4_X1 U16394 ( .A1(P1_M_IO_N_REG_SCAN_IN), .A2(P1_W_R_N_REG_SCAN_IN), .A3(
        n21256), .A4(n15321), .ZN(n13083) );
  NOR4_X1 U16395 ( .A1(P1_BE_N_REG_0__SCAN_IN), .A2(P1_BE_N_REG_1__SCAN_IN), 
        .A3(P1_BE_N_REG_2__SCAN_IN), .A4(P1_ADS_N_REG_SCAN_IN), .ZN(n13082) );
  NAND3_X1 U16396 ( .A1(n14706), .A2(n13083), .A3(n13082), .ZN(U214) );
  NOR2_X1 U16397 ( .A1(P2_BE_N_REG_0__SCAN_IN), .A2(P2_BE_N_REG_1__SCAN_IN), 
        .ZN(n13085) );
  NOR4_X1 U16398 ( .A1(P2_BE_N_REG_2__SCAN_IN), .A2(P2_BE_N_REG_3__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n13084) );
  NAND4_X1 U16399 ( .A1(P2_M_IO_N_REG_SCAN_IN), .A2(P2_W_R_N_REG_SCAN_IN), 
        .A3(n13085), .A4(n13084), .ZN(n13095) );
  NOR2_X1 U16400 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n13095), .ZN(n17255)
         );
  NOR4_X1 U16401 ( .A1(P2_ADDRESS_REG_18__SCAN_IN), .A2(
        P2_ADDRESS_REG_15__SCAN_IN), .A3(P2_ADDRESS_REG_14__SCAN_IN), .A4(
        P2_ADDRESS_REG_13__SCAN_IN), .ZN(n13089) );
  NOR4_X1 U16402 ( .A1(P2_ADDRESS_REG_23__SCAN_IN), .A2(
        P2_ADDRESS_REG_22__SCAN_IN), .A3(P2_ADDRESS_REG_20__SCAN_IN), .A4(
        P2_ADDRESS_REG_19__SCAN_IN), .ZN(n13088) );
  NOR4_X1 U16403 ( .A1(P2_ADDRESS_REG_7__SCAN_IN), .A2(
        P2_ADDRESS_REG_6__SCAN_IN), .A3(P2_ADDRESS_REG_5__SCAN_IN), .A4(
        P2_ADDRESS_REG_4__SCAN_IN), .ZN(n13087) );
  NOR4_X1 U16404 ( .A1(P2_ADDRESS_REG_11__SCAN_IN), .A2(
        P2_ADDRESS_REG_10__SCAN_IN), .A3(P2_ADDRESS_REG_9__SCAN_IN), .A4(
        P2_ADDRESS_REG_8__SCAN_IN), .ZN(n13086) );
  NAND4_X1 U16405 ( .A1(n13089), .A2(n13088), .A3(n13087), .A4(n13086), .ZN(
        n13094) );
  NOR2_X1 U16406 ( .A1(P2_ADDRESS_REG_12__SCAN_IN), .A2(
        P2_ADDRESS_REG_2__SCAN_IN), .ZN(n15206) );
  NOR3_X1 U16407 ( .A1(P2_ADDRESS_REG_3__SCAN_IN), .A2(
        P2_ADDRESS_REG_1__SCAN_IN), .A3(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n13092) );
  NOR4_X1 U16408 ( .A1(P2_ADDRESS_REG_27__SCAN_IN), .A2(
        P2_ADDRESS_REG_26__SCAN_IN), .A3(P2_ADDRESS_REG_25__SCAN_IN), .A4(
        P2_ADDRESS_REG_24__SCAN_IN), .ZN(n13091) );
  NOR4_X1 U16409 ( .A1(P2_ADDRESS_REG_17__SCAN_IN), .A2(
        P2_ADDRESS_REG_16__SCAN_IN), .A3(P2_ADDRESS_REG_21__SCAN_IN), .A4(
        P2_ADDRESS_REG_28__SCAN_IN), .ZN(n13090) );
  NAND4_X1 U16410 ( .A1(n15206), .A2(n13092), .A3(n13091), .A4(n13090), .ZN(
        n13093) );
  OAI21_X1 U16411 ( .B1(n13094), .B2(n13093), .A(P2_ADDRESS_REG_29__SCAN_IN), 
        .ZN(n13239) );
  NOR2_X1 U16412 ( .A1(n14307), .A2(n13095), .ZN(n17172) );
  NAND2_X1 U16413 ( .A1(n17172), .A2(U214), .ZN(U212) );
  AOI211_X1 U16414 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n17336), .A(n17326), .B(
        n17618), .ZN(n13105) );
  INV_X1 U16415 ( .A(n13096), .ZN(n17321) );
  AOI21_X1 U16416 ( .B1(n19628), .B2(n13097), .A(n17321), .ZN(n13104) );
  AOI211_X1 U16417 ( .C1(n18356), .C2(n13099), .A(n13098), .B(n19555), .ZN(
        n13103) );
  INV_X1 U16418 ( .A(P3_EBX_REG_26__SCAN_IN), .ZN(n13100) );
  OAI22_X1 U16419 ( .A1(n13101), .A2(n17586), .B1(n17619), .B2(n13100), .ZN(
        n13102) );
  OR4_X1 U16420 ( .A1(n13105), .A2(n13104), .A3(n13103), .A4(n13102), .ZN(
        P3_U2645) );
  INV_X1 U16421 ( .A(n11712), .ZN(n13116) );
  NAND2_X1 U16422 ( .A1(n13116), .A2(n13106), .ZN(n19925) );
  INV_X1 U16423 ( .A(n19925), .ZN(n13107) );
  INV_X1 U16424 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .ZN(n20764) );
  INV_X1 U16425 ( .A(n20696), .ZN(n16433) );
  AOI21_X1 U16426 ( .B1(n16433), .B2(n20607), .A(n14205), .ZN(n13110) );
  OAI21_X1 U16427 ( .B1(n13107), .B2(n20764), .A(n13110), .ZN(P2_U2814) );
  NOR2_X1 U16428 ( .A1(n13107), .A2(P2_READREQUEST_REG_SCAN_IN), .ZN(n13109)
         );
  INV_X1 U16429 ( .A(n13111), .ZN(n13108) );
  AOI22_X1 U16430 ( .A1(n13110), .A2(n13109), .B1(n13108), .B2(n20745), .ZN(
        P2_U3612) );
  AND2_X1 U16431 ( .A1(n13111), .A2(n20748), .ZN(n13130) );
  INV_X1 U16432 ( .A(n13734), .ZN(n13113) );
  NOR4_X1 U16433 ( .A1(n9721), .A2(n13130), .A3(n13113), .A4(n13112), .ZN(
        n13740) );
  NOR2_X1 U16434 ( .A1(n13740), .A2(n17088), .ZN(n20741) );
  OAI21_X1 U16435 ( .B1(n20741), .B2(n13115), .A(n13114), .ZN(P2_U2819) );
  NAND3_X1 U16436 ( .A1(n13116), .A2(n13139), .A3(n20755), .ZN(n13117) );
  OAI21_X1 U16437 ( .B1(n13736), .B2(n13117), .A(n13246), .ZN(n13118) );
  INV_X1 U16438 ( .A(n20027), .ZN(n13120) );
  NAND2_X1 U16439 ( .A1(n13120), .A2(n13119), .ZN(n13159) );
  INV_X1 U16440 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n16019) );
  OR2_X1 U16441 ( .A1(n20607), .A2(n13792), .ZN(n20724) );
  NOR2_X1 U16442 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n20724), .ZN(n20025) );
  INV_X1 U16443 ( .A(n20025), .ZN(n20743) );
  NAND2_X1 U16444 ( .A1(n20027), .A2(n20743), .ZN(n20020) );
  INV_X1 U16445 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n17242) );
  INV_X1 U16446 ( .A(P2_UWORD_REG_3__SCAN_IN), .ZN(n15285) );
  OAI222_X1 U16447 ( .A1(n13159), .A2(n16019), .B1(n20020), .B2(n17242), .C1(
        n15285), .C2(n20743), .ZN(P2_U2932) );
  INV_X1 U16448 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n14370) );
  INV_X1 U16449 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n17240) );
  INV_X1 U16450 ( .A(P2_UWORD_REG_1__SCAN_IN), .ZN(n13121) );
  OAI222_X1 U16451 ( .A1(n13159), .A2(n14370), .B1(n20020), .B2(n17240), .C1(
        n13121), .C2(n20743), .ZN(P2_U2934) );
  OAI21_X1 U16452 ( .B1(n13250), .B2(n15880), .A(n13122), .ZN(n13123) );
  XNOR2_X1 U16453 ( .A(n13123), .B(n16424), .ZN(n13260) );
  NOR2_X1 U16454 ( .A1(n20055), .A2(n15883), .ZN(n13127) );
  OAI21_X1 U16455 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n13125), .A(
        n13124), .ZN(n13267) );
  NAND2_X1 U16456 ( .A1(n19905), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n13261) );
  OAI21_X1 U16457 ( .B1(n20043), .B2(n13267), .A(n13261), .ZN(n13126) );
  AOI211_X1 U16458 ( .C1(n17008), .C2(n15883), .A(n13127), .B(n13126), .ZN(
        n13129) );
  NAND2_X1 U16459 ( .A1(n15888), .A2(n20051), .ZN(n13128) );
  OAI211_X1 U16460 ( .C1(n13260), .C2(n16974), .A(n13129), .B(n13128), .ZN(
        P2_U3013) );
  AND2_X1 U16461 ( .A1(n11738), .A2(n13130), .ZN(n13131) );
  AOI22_X1 U16462 ( .A1(n13132), .A2(n13754), .B1(n13131), .B2(n13734), .ZN(
        n13367) );
  NOR2_X1 U16463 ( .A1(n13132), .A2(n13752), .ZN(n13353) );
  INV_X1 U16464 ( .A(n13133), .ZN(n13134) );
  NOR2_X1 U16465 ( .A1(n13353), .A2(n13134), .ZN(n13135) );
  OAI211_X1 U16466 ( .C1(n11712), .C2(n13136), .A(n13367), .B(n13135), .ZN(
        n13779) );
  NAND2_X1 U16467 ( .A1(n20749), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n13800) );
  NOR2_X1 U16468 ( .A1(n20749), .A2(n20724), .ZN(n17080) );
  NAND2_X1 U16469 ( .A1(P2_FLUSH_REG_SCAN_IN), .A2(n17080), .ZN(n13137) );
  NAND2_X1 U16470 ( .A1(n13800), .A2(n13137), .ZN(n13138) );
  AOI21_X1 U16471 ( .B1(n13779), .B2(n13139), .A(n13138), .ZN(n16439) );
  INV_X1 U16472 ( .A(n16439), .ZN(n13145) );
  AND3_X1 U16473 ( .A1(n13142), .A2(n13141), .A3(n13140), .ZN(n13738) );
  NAND3_X1 U16474 ( .A1(n13145), .A2(n16433), .A3(n13738), .ZN(n13143) );
  OAI21_X1 U16475 ( .B1(n13145), .B2(n13144), .A(n13143), .ZN(P2_U3595) );
  INV_X1 U16476 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n15942) );
  INV_X2 U16477 ( .A(n20020), .ZN(n20024) );
  AOI22_X1 U16478 ( .A1(n20025), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(n20024), 
        .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n13146) );
  OAI21_X1 U16479 ( .B1(n15942), .B2(n13159), .A(n13146), .ZN(P2_U2923) );
  INV_X1 U16480 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n14300) );
  AOI22_X1 U16481 ( .A1(n20025), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(n20024), 
        .B2(P2_DATAO_REG_16__SCAN_IN), .ZN(n13147) );
  OAI21_X1 U16482 ( .B1(n14300), .B2(n13159), .A(n13147), .ZN(P2_U2935) );
  INV_X1 U16483 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n16007) );
  INV_X1 U16484 ( .A(n20743), .ZN(n20021) );
  AOI22_X1 U16485 ( .A1(P2_DATAO_REG_20__SCAN_IN), .A2(n20024), .B1(n20021), 
        .B2(P2_UWORD_REG_4__SCAN_IN), .ZN(n13148) );
  OAI21_X1 U16486 ( .B1(n16007), .B2(n13159), .A(n13148), .ZN(P2_U2931) );
  INV_X1 U16487 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n14578) );
  AOI22_X1 U16488 ( .A1(n20021), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n20024), 
        .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n13149) );
  OAI21_X1 U16489 ( .B1(n14578), .B2(n13159), .A(n13149), .ZN(P2_U2933) );
  INV_X1 U16490 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n15991) );
  AOI22_X1 U16491 ( .A1(n20021), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(n20024), 
        .B2(P2_DATAO_REG_22__SCAN_IN), .ZN(n13150) );
  OAI21_X1 U16492 ( .B1(n15991), .B2(n13159), .A(n13150), .ZN(P2_U2929) );
  INV_X1 U16493 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n15979) );
  AOI22_X1 U16494 ( .A1(n20021), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n20024), 
        .B2(P2_DATAO_REG_23__SCAN_IN), .ZN(n13151) );
  OAI21_X1 U16495 ( .B1(n15979), .B2(n13159), .A(n13151), .ZN(P2_U2928) );
  INV_X1 U16496 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n13242) );
  AOI22_X1 U16497 ( .A1(n20021), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n20024), 
        .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n13152) );
  OAI21_X1 U16498 ( .B1(n13242), .B2(n13159), .A(n13152), .ZN(P2_U2927) );
  INV_X1 U16499 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n15967) );
  AOI22_X1 U16500 ( .A1(n20021), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(n20024), 
        .B2(P2_DATAO_REG_25__SCAN_IN), .ZN(n13153) );
  OAI21_X1 U16501 ( .B1(n15967), .B2(n13159), .A(n13153), .ZN(P2_U2926) );
  INV_X1 U16502 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n15958) );
  AOI22_X1 U16503 ( .A1(n20021), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(n20024), 
        .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n13154) );
  OAI21_X1 U16504 ( .B1(n15958), .B2(n13159), .A(n13154), .ZN(P2_U2925) );
  INV_X1 U16505 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n15950) );
  AOI22_X1 U16506 ( .A1(n20021), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(n20024), 
        .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n13155) );
  OAI21_X1 U16507 ( .B1(n15950), .B2(n13159), .A(n13155), .ZN(P2_U2924) );
  INV_X1 U16508 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n15999) );
  AOI22_X1 U16509 ( .A1(n20021), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n20024), 
        .B2(P2_DATAO_REG_21__SCAN_IN), .ZN(n13156) );
  OAI21_X1 U16510 ( .B1(n15999), .B2(n13159), .A(n13156), .ZN(P2_U2930) );
  INV_X1 U16511 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n15934) );
  AOI22_X1 U16512 ( .A1(n20021), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(n20024), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n13157) );
  OAI21_X1 U16513 ( .B1(n15934), .B2(n13159), .A(n13157), .ZN(P2_U2922) );
  INV_X1 U16514 ( .A(P2_EAX_REG_30__SCAN_IN), .ZN(n13238) );
  AOI22_X1 U16515 ( .A1(n20021), .A2(P2_UWORD_REG_14__SCAN_IN), .B1(n20024), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .ZN(n13158) );
  OAI21_X1 U16516 ( .B1(n13238), .B2(n13159), .A(n13158), .ZN(P2_U2921) );
  INV_X1 U16517 ( .A(n13281), .ZN(n13160) );
  AND2_X1 U16518 ( .A1(n13227), .A2(n13160), .ZN(n13223) );
  NAND2_X1 U16519 ( .A1(n13223), .A2(n13289), .ZN(n13255) );
  AND2_X1 U16520 ( .A1(n21085), .A2(n16839), .ZN(n14049) );
  INV_X1 U16521 ( .A(n13651), .ZN(n13161) );
  AOI211_X1 U16522 ( .C1(P1_MEMORYFETCH_REG_SCAN_IN), .C2(n13255), .A(n14049), 
        .B(n13161), .ZN(n13162) );
  INV_X1 U16523 ( .A(n13162), .ZN(P1_U2801) );
  INV_X1 U16524 ( .A(n14205), .ZN(n13163) );
  INV_X1 U16525 ( .A(n20748), .ZN(n20744) );
  NOR3_X1 U16526 ( .A1(n13163), .A2(n9759), .A3(n20744), .ZN(n13164) );
  CLKBUF_X1 U16527 ( .A(n13164), .Z(n13240) );
  INV_X1 U16528 ( .A(n13240), .ZN(n13166) );
  INV_X1 U16529 ( .A(n13239), .ZN(n14298) );
  AOI22_X1 U16530 ( .A1(n14298), .A2(BUF1_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n14307), .ZN(n13831) );
  INV_X1 U16531 ( .A(n13246), .ZN(n13219) );
  OAI21_X1 U16532 ( .B1(n9759), .B2(n20748), .A(n14205), .ZN(n13213) );
  CLKBUF_X1 U16533 ( .A(n13213), .Z(n13243) );
  AOI22_X1 U16534 ( .A1(P2_EAX_REG_15__SCAN_IN), .A2(n13219), .B1(n13243), 
        .B2(P2_LWORD_REG_15__SCAN_IN), .ZN(n13165) );
  OAI21_X1 U16535 ( .B1(n13166), .B2(n13831), .A(n13165), .ZN(P2_U2982) );
  AOI22_X1 U16536 ( .A1(n14298), .A2(BUF1_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n14307), .ZN(n14301) );
  INV_X1 U16537 ( .A(n14301), .ZN(n13167) );
  NAND2_X1 U16538 ( .A1(n13240), .A2(n13167), .ZN(n13192) );
  AOI22_X1 U16539 ( .A1(P2_EAX_REG_16__SCAN_IN), .A2(n13219), .B1(n13243), 
        .B2(P2_UWORD_REG_0__SCAN_IN), .ZN(n13168) );
  NAND2_X1 U16540 ( .A1(n13192), .A2(n13168), .ZN(P2_U2952) );
  AOI22_X1 U16541 ( .A1(n14298), .A2(BUF1_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n13239), .ZN(n20088) );
  INV_X1 U16542 ( .A(n20088), .ZN(n13169) );
  NAND2_X1 U16543 ( .A1(n13240), .A2(n13169), .ZN(n13190) );
  AOI22_X1 U16544 ( .A1(n13214), .A2(P2_EAX_REG_17__SCAN_IN), .B1(n13243), 
        .B2(P2_UWORD_REG_1__SCAN_IN), .ZN(n13170) );
  NAND2_X1 U16545 ( .A1(n13190), .A2(n13170), .ZN(P2_U2953) );
  AOI22_X1 U16546 ( .A1(n14298), .A2(BUF1_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n14307), .ZN(n20092) );
  INV_X1 U16547 ( .A(n20092), .ZN(n13171) );
  NAND2_X1 U16548 ( .A1(n13240), .A2(n13171), .ZN(n13188) );
  AOI22_X1 U16549 ( .A1(P2_EAX_REG_18__SCAN_IN), .A2(n13219), .B1(n13213), 
        .B2(P2_UWORD_REG_2__SCAN_IN), .ZN(n13172) );
  NAND2_X1 U16550 ( .A1(n13188), .A2(n13172), .ZN(P2_U2954) );
  AOI22_X1 U16551 ( .A1(n14298), .A2(BUF1_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n14307), .ZN(n20099) );
  INV_X1 U16552 ( .A(n20099), .ZN(n13173) );
  NAND2_X1 U16553 ( .A1(n13240), .A2(n13173), .ZN(n13186) );
  AOI22_X1 U16554 ( .A1(n13214), .A2(P2_EAX_REG_19__SCAN_IN), .B1(n13243), 
        .B2(P2_UWORD_REG_3__SCAN_IN), .ZN(n13174) );
  NAND2_X1 U16555 ( .A1(n13186), .A2(n13174), .ZN(P2_U2955) );
  AOI22_X1 U16556 ( .A1(n14298), .A2(BUF1_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n14307), .ZN(n20105) );
  INV_X1 U16557 ( .A(n20105), .ZN(n13175) );
  NAND2_X1 U16558 ( .A1(n13240), .A2(n13175), .ZN(n13184) );
  AOI22_X1 U16559 ( .A1(P2_EAX_REG_20__SCAN_IN), .A2(n13219), .B1(n13213), 
        .B2(P2_UWORD_REG_4__SCAN_IN), .ZN(n13176) );
  NAND2_X1 U16560 ( .A1(n13184), .A2(n13176), .ZN(P2_U2956) );
  AOI22_X1 U16561 ( .A1(n14298), .A2(BUF1_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n14307), .ZN(n20108) );
  INV_X1 U16562 ( .A(n20108), .ZN(n13177) );
  NAND2_X1 U16563 ( .A1(n13240), .A2(n13177), .ZN(n13198) );
  AOI22_X1 U16564 ( .A1(n13219), .A2(P2_EAX_REG_21__SCAN_IN), .B1(n13213), 
        .B2(P2_UWORD_REG_5__SCAN_IN), .ZN(n13178) );
  NAND2_X1 U16565 ( .A1(n13198), .A2(n13178), .ZN(P2_U2957) );
  AOI22_X1 U16566 ( .A1(n14298), .A2(BUF1_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n14307), .ZN(n20115) );
  INV_X1 U16567 ( .A(n20115), .ZN(n13179) );
  NAND2_X1 U16568 ( .A1(n13240), .A2(n13179), .ZN(n13210) );
  AOI22_X1 U16569 ( .A1(P2_EAX_REG_22__SCAN_IN), .A2(n13219), .B1(n13213), 
        .B2(P2_UWORD_REG_6__SCAN_IN), .ZN(n13180) );
  NAND2_X1 U16570 ( .A1(n13210), .A2(n13180), .ZN(P2_U2958) );
  AOI22_X1 U16571 ( .A1(n14298), .A2(BUF1_REG_13__SCAN_IN), .B1(
        BUF2_REG_13__SCAN_IN), .B2(n13239), .ZN(n15935) );
  INV_X1 U16572 ( .A(n15935), .ZN(n13181) );
  NAND2_X1 U16573 ( .A1(n13240), .A2(n13181), .ZN(n13196) );
  AOI22_X1 U16574 ( .A1(n13214), .A2(P2_EAX_REG_13__SCAN_IN), .B1(n13213), 
        .B2(P2_LWORD_REG_13__SCAN_IN), .ZN(n13182) );
  NAND2_X1 U16575 ( .A1(n13196), .A2(n13182), .ZN(P2_U2980) );
  AOI22_X1 U16576 ( .A1(n13214), .A2(P2_EAX_REG_4__SCAN_IN), .B1(n13243), .B2(
        P2_LWORD_REG_4__SCAN_IN), .ZN(n13183) );
  NAND2_X1 U16577 ( .A1(n13184), .A2(n13183), .ZN(P2_U2971) );
  AOI22_X1 U16578 ( .A1(n13214), .A2(P2_EAX_REG_3__SCAN_IN), .B1(n13243), .B2(
        P2_LWORD_REG_3__SCAN_IN), .ZN(n13185) );
  NAND2_X1 U16579 ( .A1(n13186), .A2(n13185), .ZN(P2_U2970) );
  AOI22_X1 U16580 ( .A1(n13214), .A2(P2_EAX_REG_2__SCAN_IN), .B1(n13243), .B2(
        P2_LWORD_REG_2__SCAN_IN), .ZN(n13187) );
  NAND2_X1 U16581 ( .A1(n13188), .A2(n13187), .ZN(P2_U2969) );
  AOI22_X1 U16582 ( .A1(n13219), .A2(P2_EAX_REG_1__SCAN_IN), .B1(n13243), .B2(
        P2_LWORD_REG_1__SCAN_IN), .ZN(n13189) );
  NAND2_X1 U16583 ( .A1(n13190), .A2(n13189), .ZN(P2_U2968) );
  AOI22_X1 U16584 ( .A1(n13219), .A2(P2_EAX_REG_0__SCAN_IN), .B1(n13243), .B2(
        P2_LWORD_REG_0__SCAN_IN), .ZN(n13191) );
  NAND2_X1 U16585 ( .A1(n13192), .A2(n13191), .ZN(P2_U2967) );
  AOI22_X1 U16586 ( .A1(n14298), .A2(BUF1_REG_9__SCAN_IN), .B1(
        BUF2_REG_9__SCAN_IN), .B2(n13239), .ZN(n15968) );
  INV_X1 U16587 ( .A(n15968), .ZN(n13193) );
  NAND2_X1 U16588 ( .A1(n13240), .A2(n13193), .ZN(n13221) );
  AOI22_X1 U16589 ( .A1(P2_EAX_REG_9__SCAN_IN), .A2(n13219), .B1(n13213), .B2(
        P2_LWORD_REG_9__SCAN_IN), .ZN(n13194) );
  NAND2_X1 U16590 ( .A1(n13221), .A2(n13194), .ZN(P2_U2976) );
  AOI22_X1 U16591 ( .A1(P2_EAX_REG_29__SCAN_IN), .A2(n13219), .B1(n13243), 
        .B2(P2_UWORD_REG_13__SCAN_IN), .ZN(n13195) );
  NAND2_X1 U16592 ( .A1(n13196), .A2(n13195), .ZN(P2_U2965) );
  AOI22_X1 U16593 ( .A1(n13214), .A2(P2_EAX_REG_5__SCAN_IN), .B1(n13243), .B2(
        P2_LWORD_REG_5__SCAN_IN), .ZN(n13197) );
  NAND2_X1 U16594 ( .A1(n13198), .A2(n13197), .ZN(P2_U2972) );
  AOI22_X1 U16595 ( .A1(n14298), .A2(BUF1_REG_11__SCAN_IN), .B1(
        BUF2_REG_11__SCAN_IN), .B2(n13239), .ZN(n15951) );
  INV_X1 U16596 ( .A(n15951), .ZN(n13199) );
  NAND2_X1 U16597 ( .A1(n13240), .A2(n13199), .ZN(n13206) );
  AOI22_X1 U16598 ( .A1(P2_EAX_REG_27__SCAN_IN), .A2(n13219), .B1(n13243), 
        .B2(P2_UWORD_REG_11__SCAN_IN), .ZN(n13200) );
  NAND2_X1 U16599 ( .A1(n13206), .A2(n13200), .ZN(P2_U2963) );
  AOI22_X1 U16600 ( .A1(n14298), .A2(BUF1_REG_10__SCAN_IN), .B1(
        BUF2_REG_10__SCAN_IN), .B2(n13239), .ZN(n15959) );
  INV_X1 U16601 ( .A(n15959), .ZN(n13201) );
  NAND2_X1 U16602 ( .A1(n13240), .A2(n13201), .ZN(n13208) );
  AOI22_X1 U16603 ( .A1(P2_EAX_REG_26__SCAN_IN), .A2(n13219), .B1(n13243), 
        .B2(P2_UWORD_REG_10__SCAN_IN), .ZN(n13202) );
  NAND2_X1 U16604 ( .A1(n13208), .A2(n13202), .ZN(P2_U2962) );
  AOI22_X1 U16605 ( .A1(n14298), .A2(BUF1_REG_12__SCAN_IN), .B1(
        BUF2_REG_12__SCAN_IN), .B2(n13239), .ZN(n15943) );
  INV_X1 U16606 ( .A(n15943), .ZN(n13203) );
  NAND2_X1 U16607 ( .A1(n13240), .A2(n13203), .ZN(n13218) );
  AOI22_X1 U16608 ( .A1(P2_EAX_REG_12__SCAN_IN), .A2(n13219), .B1(n13213), 
        .B2(P2_LWORD_REG_12__SCAN_IN), .ZN(n13204) );
  NAND2_X1 U16609 ( .A1(n13218), .A2(n13204), .ZN(P2_U2979) );
  AOI22_X1 U16610 ( .A1(P2_EAX_REG_11__SCAN_IN), .A2(n13219), .B1(n13243), 
        .B2(P2_LWORD_REG_11__SCAN_IN), .ZN(n13205) );
  NAND2_X1 U16611 ( .A1(n13206), .A2(n13205), .ZN(P2_U2978) );
  AOI22_X1 U16612 ( .A1(P2_EAX_REG_10__SCAN_IN), .A2(n13219), .B1(n13213), 
        .B2(P2_LWORD_REG_10__SCAN_IN), .ZN(n13207) );
  NAND2_X1 U16613 ( .A1(n13208), .A2(n13207), .ZN(P2_U2977) );
  AOI22_X1 U16614 ( .A1(n13214), .A2(P2_EAX_REG_6__SCAN_IN), .B1(n13213), .B2(
        P2_LWORD_REG_6__SCAN_IN), .ZN(n13209) );
  NAND2_X1 U16615 ( .A1(n13210), .A2(n13209), .ZN(P2_U2973) );
  AOI22_X1 U16616 ( .A1(n14298), .A2(BUF1_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n14307), .ZN(n20123) );
  INV_X1 U16617 ( .A(n20123), .ZN(n13211) );
  NAND2_X1 U16618 ( .A1(n13240), .A2(n13211), .ZN(n13216) );
  AOI22_X1 U16619 ( .A1(n13219), .A2(P2_EAX_REG_23__SCAN_IN), .B1(n13213), 
        .B2(P2_UWORD_REG_7__SCAN_IN), .ZN(n13212) );
  NAND2_X1 U16620 ( .A1(n13216), .A2(n13212), .ZN(P2_U2959) );
  AOI22_X1 U16621 ( .A1(n13214), .A2(P2_EAX_REG_7__SCAN_IN), .B1(n13213), .B2(
        P2_LWORD_REG_7__SCAN_IN), .ZN(n13215) );
  NAND2_X1 U16622 ( .A1(n13216), .A2(n13215), .ZN(P2_U2974) );
  AOI22_X1 U16623 ( .A1(P2_EAX_REG_28__SCAN_IN), .A2(n13219), .B1(n13243), 
        .B2(P2_UWORD_REG_12__SCAN_IN), .ZN(n13217) );
  NAND2_X1 U16624 ( .A1(n13218), .A2(n13217), .ZN(P2_U2964) );
  AOI22_X1 U16625 ( .A1(P2_EAX_REG_25__SCAN_IN), .A2(n13219), .B1(n13243), 
        .B2(P2_UWORD_REG_9__SCAN_IN), .ZN(n13220) );
  NAND2_X1 U16626 ( .A1(n13221), .A2(n13220), .ZN(P2_U2961) );
  INV_X1 U16627 ( .A(n13314), .ZN(n13279) );
  OAI22_X1 U16628 ( .A1(n13223), .A2(n13222), .B1(n11194), .B2(n13279), .ZN(
        n20768) );
  NOR3_X1 U16629 ( .A1(n11194), .A2(n13275), .A3(n13273), .ZN(n13224) );
  INV_X1 U16630 ( .A(n21287), .ZN(n21190) );
  NOR2_X1 U16631 ( .A1(n13224), .A2(n21190), .ZN(n21290) );
  NOR2_X1 U16632 ( .A1(n20768), .A2(n21290), .ZN(n16488) );
  NOR2_X1 U16633 ( .A1(n16488), .A2(n20767), .ZN(n20775) );
  INV_X1 U16634 ( .A(P1_MORE_REG_SCAN_IN), .ZN(n13231) );
  NAND2_X1 U16635 ( .A1(n13225), .A2(n11547), .ZN(n13226) );
  NAND2_X1 U16636 ( .A1(n13226), .A2(n13314), .ZN(n13229) );
  AOI22_X1 U16637 ( .A1(n13303), .A2(n13279), .B1(n13227), .B2(n13281), .ZN(
        n13228) );
  NAND2_X1 U16638 ( .A1(n13229), .A2(n13228), .ZN(n16487) );
  NAND2_X1 U16639 ( .A1(n20775), .A2(n16487), .ZN(n13230) );
  OAI21_X1 U16640 ( .B1(n20775), .B2(n13231), .A(n13230), .ZN(P1_U3484) );
  INV_X1 U16641 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n19993) );
  INV_X1 U16642 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n17200) );
  OR2_X1 U16643 ( .A1(n13239), .A2(n17200), .ZN(n13233) );
  NAND2_X1 U16644 ( .A1(n13239), .A2(BUF2_REG_14__SCAN_IN), .ZN(n13232) );
  AND2_X1 U16645 ( .A1(n13233), .A2(n13232), .ZN(n19970) );
  INV_X1 U16646 ( .A(n19970), .ZN(n13234) );
  NAND2_X1 U16647 ( .A1(n13240), .A2(n13234), .ZN(n13237) );
  NAND2_X1 U16648 ( .A1(n13243), .A2(P2_LWORD_REG_14__SCAN_IN), .ZN(n13235) );
  OAI211_X1 U16649 ( .C1(n19993), .C2(n13246), .A(n13237), .B(n13235), .ZN(
        P2_U2981) );
  NAND2_X1 U16650 ( .A1(n13243), .A2(P2_UWORD_REG_14__SCAN_IN), .ZN(n13236) );
  OAI211_X1 U16651 ( .C1(n13238), .C2(n13246), .A(n13237), .B(n13236), .ZN(
        P2_U2966) );
  INV_X1 U16652 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n17207) );
  INV_X1 U16653 ( .A(BUF2_REG_8__SCAN_IN), .ZN(n18301) );
  AOI22_X1 U16654 ( .A1(n14298), .A2(n17207), .B1(n18301), .B2(n13239), .ZN(
        n19975) );
  NAND2_X1 U16655 ( .A1(n13240), .A2(n19975), .ZN(n13245) );
  NAND2_X1 U16656 ( .A1(n13243), .A2(P2_UWORD_REG_8__SCAN_IN), .ZN(n13241) );
  OAI211_X1 U16657 ( .C1(n13242), .C2(n13246), .A(n13245), .B(n13241), .ZN(
        P2_U2960) );
  INV_X1 U16658 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n20005) );
  NAND2_X1 U16659 ( .A1(n13243), .A2(P2_LWORD_REG_8__SCAN_IN), .ZN(n13244) );
  OAI211_X1 U16660 ( .C1(n20005), .C2(n13246), .A(n13245), .B(n13244), .ZN(
        P2_U2975) );
  AOI21_X1 U16661 ( .B1(n14877), .B2(n13248), .A(n13247), .ZN(n17068) );
  NOR2_X1 U16662 ( .A1(n20073), .A2(n19736), .ZN(n17073) );
  NAND2_X1 U16663 ( .A1(n19920), .A2(n14877), .ZN(n13249) );
  NAND2_X1 U16664 ( .A1(n13250), .A2(n13249), .ZN(n17070) );
  NOR2_X1 U16665 ( .A1(n16974), .A2(n17070), .ZN(n13251) );
  AOI211_X1 U16666 ( .C1(n17010), .C2(n17068), .A(n17073), .B(n13251), .ZN(
        n13254) );
  OAI21_X1 U16667 ( .B1(n20029), .B2(n13252), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13253) );
  OAI211_X1 U16668 ( .C1(n16202), .C2(n13355), .A(n13254), .B(n13253), .ZN(
        P2_U3014) );
  INV_X1 U16669 ( .A(n21285), .ZN(n13257) );
  OAI21_X1 U16670 ( .B1(n14049), .B2(P1_READREQUEST_REG_SCAN_IN), .A(n13257), 
        .ZN(n13256) );
  OAI21_X1 U16671 ( .B1(n13258), .B2(n13257), .A(n13256), .ZN(P1_U3487) );
  INV_X1 U16672 ( .A(n13260), .ZN(n13270) );
  INV_X1 U16673 ( .A(n17067), .ZN(n13262) );
  OAI21_X1 U16674 ( .B1(n13262), .B2(n16424), .A(n13261), .ZN(n13269) );
  OAI211_X1 U16675 ( .C1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(n16289), .B(n13321), .ZN(n13266) );
  OAI21_X1 U16676 ( .B1(n13264), .B2(n13263), .A(n11767), .ZN(n20712) );
  NAND2_X1 U16677 ( .A1(n20057), .A2(n20712), .ZN(n13265) );
  OAI211_X1 U16678 ( .C1(n13267), .C2(n20068), .A(n13266), .B(n13265), .ZN(
        n13268) );
  AOI211_X1 U16679 ( .C1(n20059), .C2(n13270), .A(n13269), .B(n13268), .ZN(
        n13271) );
  OAI21_X1 U16680 ( .B1(n13259), .B2(n20062), .A(n13271), .ZN(P2_U3045) );
  NAND2_X1 U16681 ( .A1(n13272), .A2(n14744), .ZN(n13274) );
  NAND2_X1 U16682 ( .A1(n13274), .A2(n13273), .ZN(n13529) );
  NAND3_X1 U16683 ( .A1(n11539), .A2(n13275), .A3(n21287), .ZN(n13277) );
  INV_X1 U16684 ( .A(n13304), .ZN(n13276) );
  NAND2_X1 U16685 ( .A1(n13277), .A2(n13276), .ZN(n13389) );
  INV_X1 U16686 ( .A(n13389), .ZN(n13278) );
  OAI21_X1 U16687 ( .B1(n13529), .B2(n21190), .A(n13278), .ZN(n13280) );
  NAND2_X1 U16688 ( .A1(n13280), .A2(n13279), .ZN(n13288) );
  INV_X1 U16689 ( .A(n11550), .ZN(n13611) );
  NOR2_X1 U16690 ( .A1(n13281), .A2(n21190), .ZN(n13282) );
  NAND2_X1 U16691 ( .A1(n13611), .A2(n13282), .ZN(n13388) );
  INV_X1 U16692 ( .A(n13283), .ZN(n13931) );
  NAND2_X1 U16693 ( .A1(n13931), .A2(n13880), .ZN(n13284) );
  AND4_X1 U16694 ( .A1(n13388), .A2(n13286), .A3(n13285), .A4(n13284), .ZN(
        n13287) );
  NAND2_X1 U16695 ( .A1(n13288), .A2(n13287), .ZN(n16475) );
  NAND2_X1 U16696 ( .A1(n16475), .A2(n13289), .ZN(n13293) );
  INV_X1 U16697 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n20774) );
  NOR2_X1 U16698 ( .A1(n21113), .A2(n16839), .ZN(n16835) );
  NAND2_X1 U16699 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n16835), .ZN(n13617) );
  NOR2_X1 U16700 ( .A1(n20774), .A2(n13617), .ZN(n13291) );
  INV_X1 U16701 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n20953) );
  NOR2_X1 U16702 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n20953), .ZN(n13290) );
  NOR2_X1 U16703 ( .A1(n13291), .A2(n13290), .ZN(n13292) );
  INV_X1 U16704 ( .A(n21275), .ZN(n15834) );
  INV_X1 U16705 ( .A(n13860), .ZN(n14091) );
  OR2_X1 U16706 ( .A1(n13294), .A2(n14091), .ZN(n13295) );
  XNOR2_X1 U16707 ( .A(n13295), .B(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n20838) );
  NAND4_X1 U16708 ( .A1(n20838), .A2(n21270), .A3(n13611), .A4(n15834), .ZN(
        n13296) );
  OAI21_X1 U16709 ( .B1(n13297), .B2(n15834), .A(n13296), .ZN(P1_U3468) );
  NOR2_X1 U16710 ( .A1(n11539), .A2(n13299), .ZN(n13300) );
  AND3_X1 U16711 ( .A1(n13301), .A2(n13300), .A3(n11550), .ZN(n14740) );
  OR2_X1 U16712 ( .A1(n9734), .A2(n14740), .ZN(n13312) );
  NOR2_X1 U16713 ( .A1(n14744), .A2(n11262), .ZN(n13302) );
  NOR2_X1 U16714 ( .A1(n14744), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n15823) );
  MUX2_X1 U16715 ( .A(n13302), .B(n15823), .S(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n13310) );
  NOR2_X1 U16716 ( .A1(n13304), .A2(n13303), .ZN(n13602) );
  XNOR2_X1 U16717 ( .A(n13305), .B(n13316), .ZN(n13315) );
  NAND2_X1 U16718 ( .A1(n11194), .A2(n13306), .ZN(n13307) );
  NOR2_X1 U16719 ( .A1(n15821), .A2(n13307), .ZN(n13598) );
  NAND2_X1 U16720 ( .A1(n13598), .A2(n13315), .ZN(n13308) );
  OAI21_X1 U16721 ( .B1(n13602), .B2(n13315), .A(n13308), .ZN(n13309) );
  NOR2_X1 U16722 ( .A1(n13310), .A2(n13309), .ZN(n13311) );
  NAND2_X1 U16723 ( .A1(n13312), .A2(n13311), .ZN(n13595) );
  NOR2_X1 U16724 ( .A1(n16839), .A2(n20930), .ZN(n15827) );
  INV_X1 U16725 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n13313) );
  AOI22_X1 U16726 ( .A1(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n13460), .B2(n13313), .ZN(
        n15825) );
  AOI222_X1 U16727 ( .A1(n13595), .A2(n21270), .B1(n15827), .B2(n15825), .C1(
        n13315), .C2(n21268), .ZN(n13317) );
  MUX2_X1 U16728 ( .A(n13317), .B(n13316), .S(n21275), .Z(n13318) );
  INV_X1 U16729 ( .A(n13318), .ZN(P1_U3472) );
  AND2_X1 U16730 ( .A1(n13319), .A2(n13336), .ZN(n13320) );
  AOI211_X1 U16731 ( .C1(n16329), .C2(n13321), .A(n17067), .B(n13320), .ZN(
        n13341) );
  INV_X1 U16732 ( .A(n13322), .ZN(n13337) );
  XNOR2_X1 U16733 ( .A(n13324), .B(n13323), .ZN(n20042) );
  NAND2_X1 U16734 ( .A1(P2_REIP_REG_2__SCAN_IN), .A2(n19905), .ZN(n20052) );
  OAI211_X1 U16735 ( .C1(n20068), .C2(n20042), .A(n13325), .B(n20052), .ZN(
        n13335) );
  NAND2_X1 U16736 ( .A1(n13327), .A2(n13326), .ZN(n13330) );
  INV_X1 U16737 ( .A(n13328), .ZN(n13329) );
  NAND2_X1 U16738 ( .A1(n13330), .A2(n13329), .ZN(n20708) );
  INV_X1 U16739 ( .A(n20708), .ZN(n13519) );
  NAND2_X1 U16740 ( .A1(n13332), .A2(n13331), .ZN(n20047) );
  NAND3_X1 U16741 ( .A1(n20048), .A2(n20059), .A3(n20047), .ZN(n13333) );
  OAI21_X1 U16742 ( .B1(n13519), .B2(n17048), .A(n13333), .ZN(n13334) );
  AOI211_X1 U16743 ( .C1(n13337), .C2(n13336), .A(n13335), .B(n13334), .ZN(
        n13339) );
  NAND2_X1 U16744 ( .A1(n10430), .A2(n17074), .ZN(n13338) );
  OAI211_X1 U16745 ( .C1(n13341), .C2(n13340), .A(n13339), .B(n13338), .ZN(
        P2_U3044) );
  OR2_X1 U16746 ( .A1(n14818), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13343) );
  NAND2_X1 U16747 ( .A1(n13343), .A2(n13342), .ZN(n20924) );
  XOR2_X1 U16748 ( .A(n13345), .B(n13344), .Z(n15454) );
  OAI222_X1 U16749 ( .A1(n20924), .A2(n15543), .B1(n15459), .B2(n16644), .C1(
        n16640), .C2(n15454), .ZN(P1_U2872) );
  NAND2_X1 U16750 ( .A1(n13436), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n13346) );
  NAND2_X1 U16751 ( .A1(n13346), .A2(n20333), .ZN(n13424) );
  NOR2_X1 U16752 ( .A1(n20509), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n13347) );
  AOI21_X1 U16753 ( .B1(n13424), .B2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n13347), .ZN(n13348) );
  NAND2_X1 U16754 ( .A1(n20755), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n13351) );
  AND4_X1 U16755 ( .A1(n13350), .A2(n13351), .A3(P2_STATE2_REG_0__SCAN_IN), 
        .A4(n20333), .ZN(n13352) );
  INV_X1 U16756 ( .A(n13353), .ZN(n13354) );
  NAND2_X1 U16757 ( .A1(n13772), .A2(n13365), .ZN(n13744) );
  NAND2_X1 U16758 ( .A1(n19969), .A2(n13368), .ZN(n19959) );
  MUX2_X1 U16759 ( .A(n10352), .B(n13355), .S(n19965), .Z(n13356) );
  OAI21_X1 U16760 ( .B1(n20727), .B2(n19959), .A(n13356), .ZN(P2_U2887) );
  NAND2_X1 U16761 ( .A1(n13424), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13357) );
  NAND2_X1 U16762 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20721), .ZN(
        n20364) );
  NAND2_X1 U16763 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20732), .ZN(
        n20397) );
  NAND2_X1 U16764 ( .A1(n20364), .A2(n20397), .ZN(n13806) );
  NAND2_X1 U16765 ( .A1(n20699), .A2(n13806), .ZN(n20400) );
  NAND2_X1 U16766 ( .A1(n13357), .A2(n20400), .ZN(n13358) );
  AND3_X1 U16767 ( .A1(n13350), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n20755), 
        .ZN(n15073) );
  INV_X1 U16768 ( .A(n15073), .ZN(n15047) );
  INV_X1 U16769 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n13359) );
  NOR2_X1 U16770 ( .A1(n15047), .A2(n13359), .ZN(n13360) );
  NAND2_X1 U16771 ( .A1(n14878), .A2(n13360), .ZN(n13361) );
  MUX2_X1 U16772 ( .A(n10557), .B(n13259), .S(n19965), .Z(n13364) );
  OAI21_X1 U16773 ( .B1(n20074), .B2(n19959), .A(n13364), .ZN(P2_U2886) );
  NAND2_X1 U16774 ( .A1(n9835), .A2(n13365), .ZN(n13366) );
  NAND2_X1 U16775 ( .A1(n19979), .A2(n13368), .ZN(n14297) );
  INV_X1 U16776 ( .A(n14297), .ZN(n13370) );
  NAND2_X1 U16777 ( .A1(n13370), .A2(n13369), .ZN(n19980) );
  NOR2_X1 U16778 ( .A1(n13372), .A2(n13371), .ZN(n13373) );
  NOR2_X1 U16779 ( .A1(n11760), .A2(n13373), .ZN(n19916) );
  NAND2_X1 U16780 ( .A1(n19979), .A2(n13374), .ZN(n19982) );
  NOR3_X1 U16781 ( .A1(n20727), .A2(n19916), .A3(n19982), .ZN(n13375) );
  AOI21_X1 U16782 ( .B1(P2_EAX_REG_0__SCAN_IN), .B2(n19974), .A(n13375), .ZN(
        n13378) );
  OAI21_X1 U16783 ( .B1(n13961), .B2(n19982), .A(n16023), .ZN(n13376) );
  NAND2_X1 U16784 ( .A1(n13376), .A2(n19916), .ZN(n13377) );
  OAI211_X1 U16785 ( .C1(n14301), .C2(n19980), .A(n13378), .B(n13377), .ZN(
        P2_U2919) );
  XNOR2_X1 U16786 ( .A(n20074), .B(n20712), .ZN(n13380) );
  NAND2_X1 U16787 ( .A1(n13961), .A2(n19916), .ZN(n13379) );
  NAND2_X1 U16788 ( .A1(n13380), .A2(n13379), .ZN(n13485) );
  OAI21_X1 U16789 ( .B1(n13380), .B2(n13379), .A(n13485), .ZN(n13381) );
  NAND2_X1 U16790 ( .A1(n13381), .A2(n16936), .ZN(n13383) );
  AOI22_X1 U16791 ( .A1(n16935), .A2(n20712), .B1(n19974), .B2(
        P2_EAX_REG_1__SCAN_IN), .ZN(n13382) );
  OAI211_X1 U16792 ( .C1(n20088), .C2(n19980), .A(n13383), .B(n13382), .ZN(
        P2_U2918) );
  OAI21_X1 U16793 ( .B1(n13385), .B2(n13384), .A(n13564), .ZN(n20844) );
  NAND2_X1 U16794 ( .A1(n13386), .A2(n11194), .ZN(n13387) );
  AOI21_X1 U16795 ( .B1(n13388), .B2(n13387), .A(n20767), .ZN(n13391) );
  AND2_X1 U16796 ( .A1(n13527), .A2(n13389), .ZN(n13390) );
  NAND2_X1 U16797 ( .A1(n13393), .A2(n13392), .ZN(n13394) );
  INV_X1 U16798 ( .A(n14706), .ZN(n13855) );
  NAND2_X1 U16799 ( .A1(n13855), .A2(DATAI_1_), .ZN(n13396) );
  NAND2_X1 U16800 ( .A1(n14706), .A2(BUF1_REG_1__SCAN_IN), .ZN(n13395) );
  AND2_X1 U16801 ( .A1(n13396), .A2(n13395), .ZN(n13888) );
  INV_X1 U16802 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n20900) );
  OAI222_X1 U16803 ( .A1(n20844), .A2(n15610), .B1(n15605), .B2(n13888), .C1(
        n15603), .C2(n20900), .ZN(P1_U2903) );
  OAI21_X1 U16804 ( .B1(n13399), .B2(n13398), .A(n13397), .ZN(n19882) );
  OAI222_X1 U16805 ( .A1(n19980), .A2(n20123), .B1(n19882), .B2(n19988), .C1(
        n20007), .C2(n19979), .ZN(P2_U2912) );
  XNOR2_X1 U16806 ( .A(n13401), .B(n13400), .ZN(n19901) );
  INV_X1 U16807 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n20010) );
  OAI222_X1 U16808 ( .A1(n19980), .A2(n20115), .B1(n19901), .B2(n19988), .C1(
        n20010), .C2(n19979), .ZN(P2_U2913) );
  AOI21_X1 U16809 ( .B1(n13403), .B2(n13402), .A(n9808), .ZN(n14239) );
  INV_X1 U16810 ( .A(n14239), .ZN(n17035) );
  INV_X1 U16811 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n20001) );
  OAI222_X1 U16812 ( .A1(n19980), .A2(n15959), .B1(n17035), .B2(n19988), .C1(
        n20001), .C2(n19979), .ZN(P2_U2909) );
  INV_X1 U16813 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n20003) );
  INV_X1 U16814 ( .A(n13404), .ZN(n14201) );
  XNOR2_X1 U16815 ( .A(n13405), .B(n14201), .ZN(n14283) );
  INV_X1 U16816 ( .A(n14283), .ZN(n16409) );
  OAI222_X1 U16817 ( .A1(n19980), .A2(n15968), .B1(n19979), .B2(n20003), .C1(
        n19988), .C2(n16409), .ZN(P2_U2910) );
  INV_X1 U16818 ( .A(n15543), .ZN(n15528) );
  INV_X1 U16819 ( .A(n13406), .ZN(n13407) );
  NAND2_X1 U16820 ( .A1(n13407), .A2(n14817), .ZN(n13409) );
  AND2_X1 U16821 ( .A1(n13409), .A2(n13408), .ZN(n20861) );
  INV_X1 U16822 ( .A(n20861), .ZN(n13410) );
  INV_X1 U16823 ( .A(n16644), .ZN(n15527) );
  AOI22_X1 U16824 ( .A1(n15528), .A2(n13410), .B1(P1_EBX_REG_1__SCAN_IN), .B2(
        n15527), .ZN(n13411) );
  OAI21_X1 U16825 ( .B1(n20844), .B2(n16640), .A(n13411), .ZN(P1_U2871) );
  NAND2_X1 U16826 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20545) );
  INV_X1 U16827 ( .A(n20545), .ZN(n13413) );
  NAND2_X1 U16828 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n13413), .ZN(
        n13421) );
  INV_X1 U16829 ( .A(n13421), .ZN(n13414) );
  NAND2_X1 U16830 ( .A1(n13414), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20080) );
  OAI211_X1 U16831 ( .C1(n13414), .C2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(
        n20080), .B(n20699), .ZN(n13415) );
  INV_X1 U16832 ( .A(n13415), .ZN(n13416) );
  AOI21_X1 U16833 ( .B1(n13424), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n13416), .ZN(n13417) );
  NAND2_X1 U16834 ( .A1(n15073), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n13435) );
  NAND2_X1 U16835 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20186) );
  NAND2_X1 U16836 ( .A1(n20186), .A2(n20710), .ZN(n13422) );
  NAND2_X1 U16837 ( .A1(n13422), .A2(n13421), .ZN(n13807) );
  NOR2_X1 U16838 ( .A1(n13807), .A2(n20509), .ZN(n13423) );
  AOI21_X1 U16839 ( .B1(n13424), .B2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n13423), .ZN(n13425) );
  NAND2_X1 U16840 ( .A1(n15073), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n13429) );
  NAND2_X1 U16841 ( .A1(n13482), .A2(n13483), .ZN(n13433) );
  INV_X1 U16842 ( .A(n13429), .ZN(n13430) );
  NAND2_X1 U16843 ( .A1(n13431), .A2(n13430), .ZN(n13432) );
  NAND2_X1 U16844 ( .A1(n13511), .A2(n13512), .ZN(n13440) );
  INV_X1 U16845 ( .A(n13435), .ZN(n13438) );
  AND2_X1 U16846 ( .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n13436), .ZN(
        n13437) );
  INV_X1 U16847 ( .A(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13441) );
  NOR2_X1 U16848 ( .A1(n15047), .A2(n13441), .ZN(n13697) );
  AND2_X1 U16849 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n13442) );
  AND2_X1 U16850 ( .A1(n13442), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n13443) );
  XNOR2_X1 U16851 ( .A(n19963), .B(n19962), .ZN(n13448) );
  INV_X1 U16852 ( .A(P2_EBX_REG_8__SCAN_IN), .ZN(n13446) );
  NOR2_X1 U16853 ( .A1(n9837), .A2(n13444), .ZN(n13445) );
  NOR2_X1 U16854 ( .A1(n9784), .A2(n13445), .ZN(n17051) );
  INV_X1 U16855 ( .A(n17051), .ZN(n16190) );
  MUX2_X1 U16856 ( .A(n13446), .B(n16190), .S(n19965), .Z(n13447) );
  OAI21_X1 U16857 ( .B1(n13448), .B2(n19959), .A(n13447), .ZN(P2_U2879) );
  XNOR2_X1 U16858 ( .A(n13449), .B(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13496) );
  NOR2_X1 U16859 ( .A1(n15738), .A2(n13450), .ZN(n13453) );
  OAI21_X1 U16860 ( .B1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n20929), .A(
        n15784), .ZN(n20931) );
  AOI22_X1 U16861 ( .A1(n16782), .A2(P1_REIP_REG_1__SCAN_IN), .B1(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n20931), .ZN(n13451) );
  OAI21_X1 U16862 ( .B1(n20925), .B2(n20861), .A(n13451), .ZN(n13452) );
  AOI21_X1 U16863 ( .B1(n13453), .B2(n13460), .A(n13452), .ZN(n13454) );
  OAI21_X1 U16864 ( .B1(n13496), .B2(n16792), .A(n13454), .ZN(P1_U3030) );
  XNOR2_X1 U16865 ( .A(n13456), .B(n13455), .ZN(n13572) );
  NOR2_X1 U16866 ( .A1(n11590), .A2(n13460), .ZN(n13556) );
  OAI21_X1 U16867 ( .B1(n15736), .B2(n13556), .A(n15784), .ZN(n15798) );
  NAND2_X1 U16868 ( .A1(n13458), .A2(n13457), .ZN(n13459) );
  NAND2_X1 U16869 ( .A1(n13558), .A2(n13459), .ZN(n13566) );
  NAND3_X1 U16870 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n15783), .A3(
        n11590), .ZN(n13465) );
  NOR2_X1 U16871 ( .A1(n20930), .A2(n13460), .ZN(n13461) );
  INV_X1 U16872 ( .A(n13555), .ZN(n13557) );
  AOI21_X1 U16873 ( .B1(n13461), .B2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A(
        n13557), .ZN(n13462) );
  INV_X1 U16874 ( .A(n13462), .ZN(n13463) );
  AND2_X1 U16875 ( .A1(n16782), .A2(P1_REIP_REG_2__SCAN_IN), .ZN(n13568) );
  AOI21_X1 U16876 ( .B1(n15733), .B2(n13463), .A(n13568), .ZN(n13464) );
  OAI211_X1 U16877 ( .C1(n20925), .C2(n13566), .A(n13465), .B(n13464), .ZN(
        n13466) );
  AOI21_X1 U16878 ( .B1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n15798), .A(
        n13466), .ZN(n13467) );
  OAI21_X1 U16879 ( .B1(n16792), .B2(n13572), .A(n13467), .ZN(P1_U3029) );
  AND2_X1 U16880 ( .A1(n13696), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n13505) );
  XNOR2_X1 U16881 ( .A(n13505), .B(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n13472) );
  NAND2_X1 U16882 ( .A1(n13468), .A2(n14268), .ZN(n13470) );
  INV_X1 U16883 ( .A(n9838), .ZN(n13469) );
  NAND2_X1 U16884 ( .A1(n13470), .A2(n13469), .ZN(n19895) );
  MUX2_X1 U16885 ( .A(n10932), .B(n19895), .S(n19965), .Z(n13471) );
  OAI21_X1 U16886 ( .B1(n13472), .B2(n19959), .A(n13471), .ZN(P2_U2881) );
  OAI21_X1 U16887 ( .B1(n13473), .B2(n9808), .A(n13502), .ZN(n19873) );
  INV_X1 U16888 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n19999) );
  OAI222_X1 U16889 ( .A1(n19980), .A2(n15951), .B1(n19873), .B2(n19988), .C1(
        n19999), .C2(n19979), .ZN(P2_U2908) );
  OR2_X1 U16890 ( .A1(n13474), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13475) );
  AND2_X1 U16891 ( .A1(n13476), .A2(n13475), .ZN(n20928) );
  INV_X1 U16892 ( .A(n20773), .ZN(n16740) );
  OAI21_X1 U16893 ( .B1(n16734), .B2(n13477), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13479) );
  INV_X1 U16894 ( .A(P1_REIP_REG_0__SCAN_IN), .ZN(n13478) );
  OR2_X1 U16895 ( .A1(n16823), .A2(n13478), .ZN(n20936) );
  NAND2_X1 U16896 ( .A1(n13479), .A2(n20936), .ZN(n13480) );
  AOI21_X1 U16897 ( .B1(n20928), .B2(n16740), .A(n13480), .ZN(n13481) );
  OAI21_X1 U16898 ( .B1(n15454), .B2(n16700), .A(n13481), .ZN(P1_U2999) );
  XNOR2_X1 U16899 ( .A(n20706), .B(n20708), .ZN(n13488) );
  INV_X1 U16900 ( .A(n20712), .ZN(n13484) );
  NAND2_X1 U16901 ( .A1(n20074), .A2(n13484), .ZN(n13486) );
  NAND2_X1 U16902 ( .A1(n13486), .A2(n13485), .ZN(n13487) );
  NAND2_X1 U16903 ( .A1(n13488), .A2(n13487), .ZN(n13520) );
  OAI21_X1 U16904 ( .B1(n13488), .B2(n13487), .A(n13520), .ZN(n13489) );
  NAND2_X1 U16905 ( .A1(n13489), .A2(n16936), .ZN(n13491) );
  AOI22_X1 U16906 ( .A1(n20708), .A2(n16935), .B1(n19974), .B2(
        P2_EAX_REG_2__SCAN_IN), .ZN(n13490) );
  OAI211_X1 U16907 ( .C1(n20092), .C2(n19980), .A(n13491), .B(n13490), .ZN(
        P2_U2917) );
  INV_X1 U16908 ( .A(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13494) );
  INV_X1 U16909 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n20846) );
  OAI22_X1 U16910 ( .A1(n16670), .A2(n13494), .B1(n16823), .B2(n20846), .ZN(
        n13493) );
  NOR2_X1 U16911 ( .A1(n20844), .A2(n16700), .ZN(n13492) );
  AOI211_X1 U16912 ( .C1(n16722), .C2(n13494), .A(n13493), .B(n13492), .ZN(
        n13495) );
  OAI21_X1 U16913 ( .B1(n13496), .B2(n20773), .A(n13495), .ZN(P1_U2998) );
  INV_X1 U16914 ( .A(n20706), .ZN(n16430) );
  MUX2_X1 U16915 ( .A(P2_EBX_REG_2__SCAN_IN), .B(n10430), .S(n19965), .Z(
        n13497) );
  AOI21_X1 U16916 ( .B1(n16430), .B2(n16926), .A(n13497), .ZN(n13498) );
  INV_X1 U16917 ( .A(n13498), .ZN(P2_U2885) );
  NAND2_X1 U16918 ( .A1(n13855), .A2(DATAI_0_), .ZN(n13500) );
  NAND2_X1 U16919 ( .A1(n14706), .A2(BUF1_REG_0__SCAN_IN), .ZN(n13499) );
  AND2_X1 U16920 ( .A1(n13500), .A2(n13499), .ZN(n13863) );
  INV_X1 U16921 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n20904) );
  OAI222_X1 U16922 ( .A1(n15610), .A2(n15454), .B1(n15605), .B2(n13863), .C1(
        n15603), .C2(n20904), .ZN(P1_U2904) );
  XNOR2_X1 U16923 ( .A(n13502), .B(n13501), .ZN(n19857) );
  INV_X1 U16924 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n19997) );
  OAI222_X1 U16925 ( .A1(n19980), .A2(n15943), .B1(n19857), .B2(n19988), .C1(
        n19997), .C2(n19979), .ZN(P2_U2907) );
  INV_X1 U16926 ( .A(n9837), .ZN(n13503) );
  OAI21_X1 U16927 ( .B1(n9838), .B2(n13504), .A(n13503), .ZN(n19881) );
  INV_X2 U16928 ( .A(n19969), .ZN(n19947) );
  INV_X1 U16929 ( .A(n13505), .ZN(n13507) );
  NOR2_X1 U16930 ( .A1(n13507), .A2(n13506), .ZN(n13508) );
  OAI211_X1 U16931 ( .C1(n13508), .C2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A(
        n16926), .B(n19963), .ZN(n13510) );
  NAND2_X1 U16932 ( .A1(n19947), .A2(P2_EBX_REG_7__SCAN_IN), .ZN(n13509) );
  OAI211_X1 U16933 ( .C1(n19881), .C2(n19947), .A(n13510), .B(n13509), .ZN(
        P2_U2880) );
  INV_X1 U16934 ( .A(n13514), .ZN(n13517) );
  INV_X1 U16935 ( .A(n13515), .ZN(n13516) );
  NAND2_X1 U16936 ( .A1(n13517), .A2(n13516), .ZN(n13518) );
  AND2_X1 U16937 ( .A1(n13518), .A2(n13701), .ZN(n20700) );
  INV_X1 U16938 ( .A(n20700), .ZN(n13700) );
  XNOR2_X1 U16939 ( .A(n20701), .B(n13700), .ZN(n13523) );
  NAND2_X1 U16940 ( .A1(n20706), .A2(n13519), .ZN(n13521) );
  NAND2_X1 U16941 ( .A1(n13521), .A2(n13520), .ZN(n13522) );
  NAND2_X1 U16942 ( .A1(n13523), .A2(n13522), .ZN(n13706) );
  OAI21_X1 U16943 ( .B1(n13523), .B2(n13522), .A(n13706), .ZN(n13524) );
  NAND2_X1 U16944 ( .A1(n13524), .A2(n16936), .ZN(n13526) );
  AOI22_X1 U16945 ( .A1(n16935), .A2(n20700), .B1(n19974), .B2(
        P2_EAX_REG_3__SCAN_IN), .ZN(n13525) );
  OAI211_X1 U16946 ( .C1(n20099), .C2(n19980), .A(n13526), .B(n13525), .ZN(
        P2_U2916) );
  INV_X1 U16947 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n13531) );
  INV_X1 U16948 ( .A(n13527), .ZN(n13528) );
  NAND2_X1 U16949 ( .A1(n20869), .A2(n11192), .ZN(n20862) );
  INV_X1 U16950 ( .A(n16835), .ZN(n16841) );
  OR2_X1 U16951 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n16841), .ZN(n20871) );
  INV_X2 U16952 ( .A(n20871), .ZN(n21288) );
  AOI22_X1 U16953 ( .A1(P1_UWORD_REG_7__SCAN_IN), .A2(n21288), .B1(n20901), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n13530) );
  OAI21_X1 U16954 ( .B1(n13531), .B2(n20862), .A(n13530), .ZN(P1_U2913) );
  INV_X1 U16955 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n13533) );
  AOI22_X1 U16956 ( .A1(P1_UWORD_REG_9__SCAN_IN), .A2(n21288), .B1(n20901), 
        .B2(P1_DATAO_REG_25__SCAN_IN), .ZN(n13532) );
  OAI21_X1 U16957 ( .B1(n13533), .B2(n20862), .A(n13532), .ZN(P1_U2911) );
  AOI22_X1 U16958 ( .A1(P1_UWORD_REG_5__SCAN_IN), .A2(n21288), .B1(n20901), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n13534) );
  OAI21_X1 U16959 ( .B1(n12332), .B2(n20862), .A(n13534), .ZN(P1_U2915) );
  INV_X1 U16960 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n13536) );
  AOI22_X1 U16961 ( .A1(P1_UWORD_REG_4__SCAN_IN), .A2(n21288), .B1(n20901), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n13535) );
  OAI21_X1 U16962 ( .B1(n13536), .B2(n20862), .A(n13535), .ZN(P1_U2916) );
  INV_X1 U16963 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n13538) );
  AOI22_X1 U16964 ( .A1(P1_UWORD_REG_0__SCAN_IN), .A2(n21288), .B1(n20901), 
        .B2(P1_DATAO_REG_16__SCAN_IN), .ZN(n13537) );
  OAI21_X1 U16965 ( .B1(n13538), .B2(n20862), .A(n13537), .ZN(P1_U2920) );
  INV_X1 U16966 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n13540) );
  AOI22_X1 U16967 ( .A1(P1_UWORD_REG_12__SCAN_IN), .A2(n21288), .B1(n20901), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n13539) );
  OAI21_X1 U16968 ( .B1(n13540), .B2(n20862), .A(n13539), .ZN(P1_U2908) );
  INV_X1 U16969 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n13542) );
  AOI22_X1 U16970 ( .A1(P1_UWORD_REG_2__SCAN_IN), .A2(n21288), .B1(n20901), 
        .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n13541) );
  OAI21_X1 U16971 ( .B1(n13542), .B2(n20862), .A(n13541), .ZN(P1_U2918) );
  INV_X1 U16972 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n13544) );
  AOI22_X1 U16973 ( .A1(P1_UWORD_REG_10__SCAN_IN), .A2(n21288), .B1(n20901), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n13543) );
  OAI21_X1 U16974 ( .B1(n13544), .B2(n20862), .A(n13543), .ZN(P1_U2910) );
  INV_X1 U16975 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n15283) );
  AOI22_X1 U16976 ( .A1(P1_UWORD_REG_3__SCAN_IN), .A2(n21288), .B1(n20901), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n13545) );
  OAI21_X1 U16977 ( .B1(n15283), .B2(n20862), .A(n13545), .ZN(P1_U2917) );
  INV_X1 U16978 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n13547) );
  AOI22_X1 U16979 ( .A1(P1_UWORD_REG_8__SCAN_IN), .A2(n21288), .B1(n20901), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n13546) );
  OAI21_X1 U16980 ( .B1(n13547), .B2(n20862), .A(n13546), .ZN(P1_U2912) );
  INV_X1 U16981 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n13549) );
  AOI22_X1 U16982 ( .A1(P1_UWORD_REG_1__SCAN_IN), .A2(n21288), .B1(n20901), 
        .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n13548) );
  OAI21_X1 U16983 ( .B1(n13549), .B2(n20862), .A(n13548), .ZN(P1_U2919) );
  INV_X1 U16984 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n15366) );
  AOI22_X1 U16985 ( .A1(P1_UWORD_REG_14__SCAN_IN), .A2(n21288), .B1(n20901), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .ZN(n13550) );
  OAI21_X1 U16986 ( .B1(n15366), .B2(n20862), .A(n13550), .ZN(P1_U2906) );
  INV_X1 U16987 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n13552) );
  AOI22_X1 U16988 ( .A1(P1_UWORD_REG_13__SCAN_IN), .A2(n21288), .B1(n20901), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n13551) );
  OAI21_X1 U16989 ( .B1(n13552), .B2(n20862), .A(n13551), .ZN(P1_U2907) );
  XNOR2_X1 U16990 ( .A(n9733), .B(n13554), .ZN(n13632) );
  INV_X1 U16991 ( .A(n15798), .ZN(n13846) );
  OAI21_X1 U16992 ( .B1(n20929), .B2(n13555), .A(n13846), .ZN(n13802) );
  AOI21_X1 U16993 ( .B1(n13556), .B2(n15783), .A(n15733), .ZN(n15770) );
  NOR2_X1 U16994 ( .A1(n13557), .A2(n15770), .ZN(n13849) );
  AOI22_X1 U16995 ( .A1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n13802), .B1(
        n13849), .B2(n11317), .ZN(n13561) );
  AOI21_X1 U16996 ( .B1(n13559), .B2(n13558), .A(n13725), .ZN(n13954) );
  INV_X1 U16997 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n21200) );
  NOR2_X1 U16998 ( .A1(n16823), .A2(n21200), .ZN(n13629) );
  AOI21_X1 U16999 ( .B1(n13954), .B2(n16809), .A(n13629), .ZN(n13560) );
  OAI211_X1 U17000 ( .C1(n16792), .C2(n13632), .A(n13561), .B(n13560), .ZN(
        P1_U3028) );
  INV_X1 U17001 ( .A(n13562), .ZN(n13563) );
  AOI21_X1 U17002 ( .B1(n13565), .B2(n13564), .A(n13563), .ZN(n14831) );
  INV_X1 U17003 ( .A(n14831), .ZN(n13578) );
  INV_X1 U17004 ( .A(n13566), .ZN(n14841) );
  AOI22_X1 U17005 ( .A1(n14841), .A2(n15528), .B1(P1_EBX_REG_2__SCAN_IN), .B2(
        n15527), .ZN(n13567) );
  OAI21_X1 U17006 ( .B1(n13578), .B2(n16640), .A(n13567), .ZN(P1_U2870) );
  AOI21_X1 U17007 ( .B1(n16734), .B2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .A(
        n13568), .ZN(n13569) );
  OAI21_X1 U17008 ( .B1(n14834), .B2(n16743), .A(n13569), .ZN(n13570) );
  AOI21_X1 U17009 ( .B1(n14831), .B2(n16739), .A(n13570), .ZN(n13571) );
  OAI21_X1 U17010 ( .B1(n20773), .B2(n13572), .A(n13571), .ZN(P1_U2997) );
  OAI21_X1 U17011 ( .B1(n13575), .B2(n9822), .A(n13574), .ZN(n19849) );
  INV_X1 U17012 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n19995) );
  OAI222_X1 U17013 ( .A1(n19980), .A2(n15935), .B1(n19849), .B2(n19988), .C1(
        n19995), .C2(n19979), .ZN(P2_U2906) );
  NAND2_X1 U17014 ( .A1(n13855), .A2(DATAI_2_), .ZN(n13577) );
  NAND2_X1 U17015 ( .A1(n14706), .A2(BUF1_REG_2__SCAN_IN), .ZN(n13576) );
  AND2_X1 U17016 ( .A1(n13577), .A2(n13576), .ZN(n13881) );
  INV_X1 U17017 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n20898) );
  OAI222_X1 U17018 ( .A1(n13578), .A2(n15610), .B1(n15605), .B2(n13881), .C1(
        n15603), .C2(n20898), .ZN(P1_U2902) );
  AND2_X1 U17019 ( .A1(n20701), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n20554) );
  NAND2_X1 U17020 ( .A1(n20554), .A2(n20695), .ZN(n13579) );
  NOR2_X1 U17021 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n10567), .ZN(
        n20331) );
  NAND2_X1 U17022 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20331), .ZN(
        n13590) );
  NAND2_X1 U17023 ( .A1(n13579), .A2(n13590), .ZN(n13586) );
  OR2_X1 U17024 ( .A1(n10620), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n13584) );
  INV_X1 U17025 ( .A(n20331), .ZN(n20401) );
  NOR2_X1 U17026 ( .A1(n20186), .A2(n20401), .ZN(n20443) );
  NOR2_X1 U17027 ( .A1(n20443), .A2(n20699), .ZN(n13583) );
  OAI21_X1 U17028 ( .B1(P2_STATE2_REG_2__SCAN_IN), .B2(
        P2_STATE2_REG_1__SCAN_IN), .A(n20749), .ZN(n20753) );
  INV_X1 U17029 ( .A(n20753), .ZN(n13580) );
  NAND2_X1 U17030 ( .A1(n20724), .A2(n13580), .ZN(n13581) );
  AOI21_X1 U17031 ( .B1(n13584), .B2(n13583), .A(n20551), .ZN(n13585) );
  NAND2_X1 U17032 ( .A1(n13586), .A2(n13585), .ZN(n20439) );
  INV_X1 U17033 ( .A(n20439), .ZN(n20449) );
  INV_X1 U17034 ( .A(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n14177) );
  AND2_X1 U17035 ( .A1(n20699), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n20711) );
  AOI22_X1 U17036 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n20119), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n20118), .ZN(n20521) );
  NAND2_X1 U17037 ( .A1(n20701), .A2(n13961), .ZN(n20474) );
  NOR2_X2 U17038 ( .A1(n20474), .A2(n20187), .ZN(n20467) );
  AOI22_X1 U17039 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n20119), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n20118), .ZN(n20560) );
  INV_X1 U17040 ( .A(n20560), .ZN(n20506) );
  AOI22_X1 U17041 ( .A1(n20445), .A2(n20557), .B1(n20467), .B2(n20506), .ZN(
        n13594) );
  INV_X1 U17042 ( .A(n10620), .ZN(n13588) );
  OAI21_X1 U17043 ( .B1(n13588), .B2(n20443), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n13589) );
  OAI21_X1 U17044 ( .B1(n13590), .B2(n20509), .A(n13589), .ZN(n20444) );
  AOI22_X1 U17045 ( .A1(n20444), .A2(n13591), .B1(n20548), .B2(n20443), .ZN(
        n13593) );
  OAI211_X1 U17046 ( .C1(n20449), .C2(n14177), .A(n13594), .B(n13593), .ZN(
        P2_U3136) );
  NOR2_X1 U17047 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n16839), .ZN(n13612) );
  MUX2_X1 U17048 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n13595), .S(
        n16475), .Z(n16472) );
  AOI22_X1 U17049 ( .A1(n13612), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n16839), .B2(n16472), .ZN(n13609) );
  INV_X1 U17050 ( .A(n14055), .ZN(n15819) );
  OAI21_X1 U17051 ( .B1(n13602), .B2(n13305), .A(n14744), .ZN(n13600) );
  INV_X1 U17052 ( .A(n13599), .ZN(n13596) );
  OAI211_X1 U17053 ( .C1(n13305), .C2(n11043), .A(n13597), .B(n13596), .ZN(
        n21269) );
  AOI22_X1 U17054 ( .A1(n13600), .A2(n13599), .B1(n13598), .B2(n21269), .ZN(
        n13607) );
  NAND2_X1 U17055 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13603) );
  NOR2_X1 U17056 ( .A1(n13305), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13601) );
  OAI22_X1 U17057 ( .A1(n13603), .A2(n14744), .B1(n13602), .B2(n13601), .ZN(
        n13604) );
  MUX2_X1 U17058 ( .A(n13604), .B(n15823), .S(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n13605) );
  INV_X1 U17059 ( .A(n13605), .ZN(n13606) );
  OAI211_X1 U17060 ( .C1(n15819), .C2(n14740), .A(n13607), .B(n13606), .ZN(
        n21271) );
  MUX2_X1 U17061 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n21271), .S(
        n16475), .Z(n16484) );
  AOI22_X1 U17062 ( .A1(n13612), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n16484), .B2(n16839), .ZN(n13608) );
  NOR2_X1 U17063 ( .A1(n13609), .A2(n13608), .ZN(n16494) );
  INV_X1 U17064 ( .A(n16494), .ZN(n13610) );
  NOR2_X1 U17065 ( .A1(n13610), .A2(n15828), .ZN(n13619) );
  NAND3_X1 U17066 ( .A1(n20838), .A2(n13611), .A3(n16839), .ZN(n13616) );
  INV_X1 U17067 ( .A(n13612), .ZN(n13613) );
  OAI21_X1 U17068 ( .B1(n16475), .B2(P1_STATE2_REG_1__SCAN_IN), .A(n13613), 
        .ZN(n13614) );
  NAND2_X1 U17069 ( .A1(n13614), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n13615) );
  NAND2_X1 U17070 ( .A1(n13616), .A2(n13615), .ZN(n16493) );
  NOR3_X1 U17071 ( .A1(n13619), .A2(n16493), .A3(P1_FLUSH_REG_SCAN_IN), .ZN(
        n13618) );
  NOR2_X1 U17072 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n21291) );
  OAI21_X1 U17073 ( .B1(n13618), .B2(n13617), .A(n14095), .ZN(n20938) );
  NOR3_X1 U17074 ( .A1(n13619), .A2(n16493), .A3(n16841), .ZN(n16502) );
  AND2_X1 U17075 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n20953), .ZN(n15818) );
  OAI22_X1 U17076 ( .A1(n14398), .A2(n21122), .B1(n10102), .B2(n15818), .ZN(
        n13620) );
  OAI21_X1 U17077 ( .B1(n16502), .B2(n13620), .A(n20938), .ZN(n13621) );
  OAI21_X1 U17078 ( .B1(n20938), .B2(n21110), .A(n13621), .ZN(P1_U3478) );
  INV_X1 U17079 ( .A(n13622), .ZN(n13623) );
  NOR2_X1 U17080 ( .A1(n13624), .A2(n13623), .ZN(n13626) );
  AOI21_X1 U17081 ( .B1(n13626), .B2(n13562), .A(n13625), .ZN(n13935) );
  INV_X1 U17082 ( .A(n13935), .ZN(n13635) );
  AOI22_X1 U17083 ( .A1(n13954), .A2(n15528), .B1(P1_EBX_REG_3__SCAN_IN), .B2(
        n15527), .ZN(n13627) );
  OAI21_X1 U17084 ( .B1(n13635), .B2(n16640), .A(n13627), .ZN(P1_U2869) );
  NOR2_X1 U17085 ( .A1(n16670), .A2(n13948), .ZN(n13628) );
  AOI211_X1 U17086 ( .C1(n16722), .C2(n13944), .A(n13629), .B(n13628), .ZN(
        n13631) );
  NAND2_X1 U17087 ( .A1(n13935), .A2(n16739), .ZN(n13630) );
  OAI211_X1 U17088 ( .C1(n13632), .C2(n20773), .A(n13631), .B(n13630), .ZN(
        P1_U2996) );
  NAND2_X1 U17089 ( .A1(n13855), .A2(DATAI_3_), .ZN(n13634) );
  NAND2_X1 U17090 ( .A1(n14706), .A2(BUF1_REG_3__SCAN_IN), .ZN(n13633) );
  AND2_X1 U17091 ( .A1(n13634), .A2(n13633), .ZN(n13871) );
  INV_X1 U17092 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n20896) );
  OAI222_X1 U17093 ( .A1(n13635), .A2(n15610), .B1(n15605), .B2(n13871), .C1(
        n15603), .C2(n20896), .ZN(P1_U2901) );
  NAND2_X1 U17094 ( .A1(n13639), .A2(n13638), .ZN(n13712) );
  OR2_X1 U17095 ( .A1(n19953), .A2(n13712), .ZN(n19949) );
  XNOR2_X1 U17096 ( .A(n19949), .B(n13711), .ZN(n13648) );
  INV_X1 U17097 ( .A(n13640), .ZN(n13642) );
  INV_X1 U17098 ( .A(n13643), .ZN(n13641) );
  NAND2_X1 U17099 ( .A1(n13642), .A2(n13641), .ZN(n13644) );
  NAND2_X1 U17100 ( .A1(n13640), .A2(n13643), .ZN(n16965) );
  AND2_X1 U17101 ( .A1(n13644), .A2(n16965), .ZN(n19856) );
  INV_X1 U17102 ( .A(P2_EBX_REG_12__SCAN_IN), .ZN(n13645) );
  NOR2_X1 U17103 ( .A1(n19969), .A2(n13645), .ZN(n13646) );
  AOI21_X1 U17104 ( .B1(n19856), .B2(n19969), .A(n13646), .ZN(n13647) );
  OAI21_X1 U17105 ( .B1(n13648), .B2(n19959), .A(n13647), .ZN(P2_U2875) );
  AND2_X1 U17106 ( .A1(n13649), .A2(n21190), .ZN(n13650) );
  OR2_X2 U17107 ( .A1(n13651), .A2(n13650), .ZN(n20921) );
  OR2_X1 U17108 ( .A1(n20921), .A2(n11177), .ZN(n13695) );
  AOI22_X1 U17109 ( .A1(n9717), .A2(P1_EAX_REG_25__SCAN_IN), .B1(
        P1_UWORD_REG_9__SCAN_IN), .B2(n20921), .ZN(n13653) );
  MUX2_X1 U17110 ( .A(DATAI_9_), .B(BUF1_REG_9__SCAN_IN), .S(n14706), .Z(
        n15561) );
  NAND2_X1 U17111 ( .A1(n13652), .A2(n15561), .ZN(n20913) );
  NAND2_X1 U17112 ( .A1(n13653), .A2(n20913), .ZN(P1_U2946) );
  AOI22_X1 U17113 ( .A1(n9717), .A2(P1_EAX_REG_29__SCAN_IN), .B1(
        P1_UWORD_REG_13__SCAN_IN), .B2(n20921), .ZN(n13654) );
  MUX2_X1 U17114 ( .A(DATAI_13_), .B(BUF1_REG_13__SCAN_IN), .S(n14706), .Z(
        n15550) );
  NAND2_X1 U17115 ( .A1(n13652), .A2(n15550), .ZN(n20919) );
  NAND2_X1 U17116 ( .A1(n13654), .A2(n20919), .ZN(P1_U2950) );
  AOI22_X1 U17117 ( .A1(n9717), .A2(P1_EAX_REG_21__SCAN_IN), .B1(
        P1_UWORD_REG_5__SCAN_IN), .B2(n20921), .ZN(n13657) );
  NAND2_X1 U17118 ( .A1(n13855), .A2(DATAI_5_), .ZN(n13656) );
  NAND2_X1 U17119 ( .A1(n14706), .A2(BUF1_REG_5__SCAN_IN), .ZN(n13655) );
  AND2_X1 U17120 ( .A1(n13656), .A2(n13655), .ZN(n13876) );
  INV_X1 U17121 ( .A(n13876), .ZN(n15575) );
  NAND2_X1 U17122 ( .A1(n13652), .A2(n15575), .ZN(n13679) );
  NAND2_X1 U17123 ( .A1(n13657), .A2(n13679), .ZN(P1_U2942) );
  AOI22_X1 U17124 ( .A1(n9717), .A2(P1_EAX_REG_20__SCAN_IN), .B1(
        P1_UWORD_REG_4__SCAN_IN), .B2(n20921), .ZN(n13660) );
  NAND2_X1 U17125 ( .A1(n13855), .A2(DATAI_4_), .ZN(n13659) );
  NAND2_X1 U17126 ( .A1(n14706), .A2(BUF1_REG_4__SCAN_IN), .ZN(n13658) );
  AND2_X1 U17127 ( .A1(n13659), .A2(n13658), .ZN(n13972) );
  INV_X1 U17128 ( .A(n13972), .ZN(n15578) );
  NAND2_X1 U17129 ( .A1(n13652), .A2(n15578), .ZN(n13681) );
  NAND2_X1 U17130 ( .A1(n13660), .A2(n13681), .ZN(P1_U2941) );
  AOI22_X1 U17131 ( .A1(n9717), .A2(P1_EAX_REG_17__SCAN_IN), .B1(
        P1_UWORD_REG_1__SCAN_IN), .B2(n20921), .ZN(n13661) );
  INV_X1 U17132 ( .A(n13888), .ZN(n15591) );
  NAND2_X1 U17133 ( .A1(n13652), .A2(n15591), .ZN(n13666) );
  NAND2_X1 U17134 ( .A1(n13661), .A2(n13666), .ZN(P1_U2938) );
  AOI22_X1 U17135 ( .A1(n9717), .A2(P1_EAX_REG_23__SCAN_IN), .B1(
        P1_UWORD_REG_7__SCAN_IN), .B2(n20921), .ZN(n13664) );
  NAND2_X1 U17136 ( .A1(n13855), .A2(DATAI_7_), .ZN(n13663) );
  NAND2_X1 U17137 ( .A1(n14706), .A2(BUF1_REG_7__SCAN_IN), .ZN(n13662) );
  AND2_X1 U17138 ( .A1(n13663), .A2(n13662), .ZN(n14233) );
  INV_X1 U17139 ( .A(n14233), .ZN(n15567) );
  NAND2_X1 U17140 ( .A1(n13652), .A2(n15567), .ZN(n13673) );
  NAND2_X1 U17141 ( .A1(n13664), .A2(n13673), .ZN(P1_U2944) );
  AOI22_X1 U17142 ( .A1(n9717), .A2(P1_EAX_REG_0__SCAN_IN), .B1(
        P1_LWORD_REG_0__SCAN_IN), .B2(n20921), .ZN(n13665) );
  INV_X1 U17143 ( .A(n13863), .ZN(n15597) );
  NAND2_X1 U17144 ( .A1(n13652), .A2(n15597), .ZN(n13677) );
  NAND2_X1 U17145 ( .A1(n13665), .A2(n13677), .ZN(P1_U2952) );
  AOI22_X1 U17146 ( .A1(n9717), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_LWORD_REG_1__SCAN_IN), .B2(n20921), .ZN(n13667) );
  NAND2_X1 U17147 ( .A1(n13667), .A2(n13666), .ZN(P1_U2953) );
  AOI22_X1 U17148 ( .A1(n9717), .A2(P1_EAX_REG_2__SCAN_IN), .B1(
        P1_LWORD_REG_2__SCAN_IN), .B2(n20921), .ZN(n13668) );
  INV_X1 U17149 ( .A(n13881), .ZN(n15588) );
  NAND2_X1 U17150 ( .A1(n13652), .A2(n15588), .ZN(n13683) );
  NAND2_X1 U17151 ( .A1(n13668), .A2(n13683), .ZN(P1_U2954) );
  AOI22_X1 U17152 ( .A1(n9717), .A2(P1_EAX_REG_6__SCAN_IN), .B1(
        P1_LWORD_REG_6__SCAN_IN), .B2(n20921), .ZN(n13671) );
  NAND2_X1 U17153 ( .A1(n13855), .A2(DATAI_6_), .ZN(n13670) );
  NAND2_X1 U17154 ( .A1(n14706), .A2(BUF1_REG_6__SCAN_IN), .ZN(n13669) );
  AND2_X1 U17155 ( .A1(n13670), .A2(n13669), .ZN(n13980) );
  INV_X1 U17156 ( .A(n13980), .ZN(n15571) );
  NAND2_X1 U17157 ( .A1(n13652), .A2(n15571), .ZN(n13675) );
  NAND2_X1 U17158 ( .A1(n13671), .A2(n13675), .ZN(P1_U2958) );
  AOI22_X1 U17159 ( .A1(n9717), .A2(P1_EAX_REG_19__SCAN_IN), .B1(
        P1_UWORD_REG_3__SCAN_IN), .B2(n20921), .ZN(n13672) );
  INV_X1 U17160 ( .A(n13871), .ZN(n15585) );
  NAND2_X1 U17161 ( .A1(n13652), .A2(n15585), .ZN(n13685) );
  NAND2_X1 U17162 ( .A1(n13672), .A2(n13685), .ZN(P1_U2940) );
  AOI22_X1 U17163 ( .A1(n9717), .A2(P1_EAX_REG_7__SCAN_IN), .B1(
        P1_LWORD_REG_7__SCAN_IN), .B2(n20921), .ZN(n13674) );
  NAND2_X1 U17164 ( .A1(n13674), .A2(n13673), .ZN(P1_U2959) );
  AOI22_X1 U17165 ( .A1(n9717), .A2(P1_EAX_REG_22__SCAN_IN), .B1(
        P1_UWORD_REG_6__SCAN_IN), .B2(n20921), .ZN(n13676) );
  NAND2_X1 U17166 ( .A1(n13676), .A2(n13675), .ZN(P1_U2943) );
  AOI22_X1 U17167 ( .A1(n9717), .A2(P1_EAX_REG_16__SCAN_IN), .B1(
        P1_UWORD_REG_0__SCAN_IN), .B2(n20921), .ZN(n13678) );
  NAND2_X1 U17168 ( .A1(n13678), .A2(n13677), .ZN(P1_U2937) );
  AOI22_X1 U17169 ( .A1(n9717), .A2(P1_EAX_REG_5__SCAN_IN), .B1(
        P1_LWORD_REG_5__SCAN_IN), .B2(n20921), .ZN(n13680) );
  NAND2_X1 U17170 ( .A1(n13680), .A2(n13679), .ZN(P1_U2957) );
  AOI22_X1 U17171 ( .A1(n9717), .A2(P1_EAX_REG_4__SCAN_IN), .B1(
        P1_LWORD_REG_4__SCAN_IN), .B2(n20921), .ZN(n13682) );
  NAND2_X1 U17172 ( .A1(n13682), .A2(n13681), .ZN(P1_U2956) );
  AOI22_X1 U17173 ( .A1(n9717), .A2(P1_EAX_REG_18__SCAN_IN), .B1(
        P1_UWORD_REG_2__SCAN_IN), .B2(n20921), .ZN(n13684) );
  NAND2_X1 U17174 ( .A1(n13684), .A2(n13683), .ZN(P1_U2939) );
  AOI22_X1 U17175 ( .A1(n9717), .A2(P1_EAX_REG_3__SCAN_IN), .B1(
        P1_LWORD_REG_3__SCAN_IN), .B2(n20921), .ZN(n13686) );
  NAND2_X1 U17176 ( .A1(n13686), .A2(n13685), .ZN(P1_U2955) );
  AOI22_X1 U17177 ( .A1(n9717), .A2(P1_EAX_REG_27__SCAN_IN), .B1(
        P1_UWORD_REG_11__SCAN_IN), .B2(n20921), .ZN(n13687) );
  MUX2_X1 U17178 ( .A(DATAI_11_), .B(BUF1_REG_11__SCAN_IN), .S(n14706), .Z(
        n15554) );
  NAND2_X1 U17179 ( .A1(n13652), .A2(n15554), .ZN(n13688) );
  NAND2_X1 U17180 ( .A1(n13687), .A2(n13688), .ZN(P1_U2948) );
  AOI22_X1 U17181 ( .A1(n9717), .A2(P1_EAX_REG_11__SCAN_IN), .B1(
        P1_LWORD_REG_11__SCAN_IN), .B2(n20921), .ZN(n13689) );
  NAND2_X1 U17182 ( .A1(n13689), .A2(n13688), .ZN(P1_U2963) );
  NAND2_X1 U17183 ( .A1(n20921), .A2(P1_UWORD_REG_14__SCAN_IN), .ZN(n13690) );
  MUX2_X1 U17184 ( .A(DATAI_14_), .B(BUF1_REG_14__SCAN_IN), .S(n14706), .Z(
        n15607) );
  NAND2_X1 U17185 ( .A1(n13652), .A2(n15607), .ZN(n20922) );
  OAI211_X1 U17186 ( .C1(n13695), .C2(n15366), .A(n13690), .B(n20922), .ZN(
        P1_U2951) );
  INV_X1 U17187 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n15602) );
  INV_X1 U17188 ( .A(n13652), .ZN(n13694) );
  INV_X1 U17189 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n13691) );
  NOR2_X1 U17190 ( .A1(n13855), .A2(n13691), .ZN(n13692) );
  AOI21_X1 U17191 ( .B1(DATAI_15_), .B2(n13855), .A(n13692), .ZN(n15604) );
  INV_X1 U17192 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n20872) );
  OAI222_X1 U17193 ( .A1(n13695), .A2(n15602), .B1(n13694), .B2(n15604), .C1(
        n13693), .C2(n20872), .ZN(P1_U2967) );
  OR2_X1 U17194 ( .A1(n13698), .A2(n13697), .ZN(n13699) );
  NAND2_X1 U17195 ( .A1(n14851), .A2(n13699), .ZN(n19983) );
  NAND2_X1 U17196 ( .A1(n20131), .A2(n13700), .ZN(n13707) );
  NAND2_X1 U17197 ( .A1(n13702), .A2(n13701), .ZN(n13705) );
  INV_X1 U17198 ( .A(n13703), .ZN(n13704) );
  AND2_X1 U17199 ( .A1(n13705), .A2(n13704), .ZN(n20056) );
  AOI21_X1 U17200 ( .B1(n13707), .B2(n13706), .A(n20056), .ZN(n19984) );
  XOR2_X1 U17201 ( .A(n19983), .B(n19984), .Z(n13708) );
  NAND2_X1 U17202 ( .A1(n13708), .A2(n16936), .ZN(n13710) );
  AOI22_X1 U17203 ( .A1(n16935), .A2(n20056), .B1(n19974), .B2(
        P2_EAX_REG_4__SCAN_IN), .ZN(n13709) );
  OAI211_X1 U17204 ( .C1(n20105), .C2(n19980), .A(n13710), .B(n13709), .ZN(
        P2_U2915) );
  OR2_X1 U17205 ( .A1(n13712), .A2(n13711), .ZN(n19941) );
  INV_X1 U17206 ( .A(n13713), .ZN(n19942) );
  OR2_X1 U17207 ( .A1(n19941), .A2(n19942), .ZN(n14190) );
  NOR2_X1 U17208 ( .A1(n19953), .A2(n14190), .ZN(n14251) );
  INV_X1 U17209 ( .A(n14251), .ZN(n19944) );
  XNOR2_X1 U17210 ( .A(n19944), .B(n19934), .ZN(n13719) );
  OR2_X1 U17211 ( .A1(n16966), .A2(n13715), .ZN(n13716) );
  AND2_X1 U17212 ( .A1(n13714), .A2(n13716), .ZN(n19835) );
  NOR2_X1 U17213 ( .A1(n19969), .A2(n10757), .ZN(n13717) );
  AOI21_X1 U17214 ( .B1(n19835), .B2(n19969), .A(n13717), .ZN(n13718) );
  OAI21_X1 U17215 ( .B1(n13719), .B2(n19959), .A(n13718), .ZN(P2_U2873) );
  INV_X1 U17216 ( .A(n13720), .ZN(n13723) );
  INV_X1 U17217 ( .A(n13625), .ZN(n13722) );
  AOI21_X1 U17218 ( .B1(n13723), .B2(n13722), .A(n13721), .ZN(n20841) );
  INV_X1 U17219 ( .A(n20841), .ZN(n13728) );
  INV_X1 U17220 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n13727) );
  OR2_X1 U17221 ( .A1(n13725), .A2(n13724), .ZN(n13726) );
  NAND2_X1 U17222 ( .A1(n13823), .A2(n13726), .ZN(n20835) );
  OAI222_X1 U17223 ( .A1(n13728), .A2(n16640), .B1(n13727), .B2(n16644), .C1(
        n20835), .C2(n15543), .ZN(P1_U2868) );
  INV_X1 U17224 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n20893) );
  OAI222_X1 U17225 ( .A1(n13728), .A2(n15610), .B1(n15605), .B2(n13972), .C1(
        n15603), .C2(n20893), .ZN(P1_U2900) );
  XNOR2_X1 U17226 ( .A(n13729), .B(n13730), .ZN(n13805) );
  AOI22_X1 U17227 ( .A1(n16734), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B1(
        n16782), .B2(P1_REIP_REG_4__SCAN_IN), .ZN(n13731) );
  OAI21_X1 U17228 ( .B1(n20839), .B2(n16743), .A(n13731), .ZN(n13732) );
  AOI21_X1 U17229 ( .B1(n20841), .B2(n16739), .A(n13732), .ZN(n13733) );
  OAI21_X1 U17230 ( .B1(n13805), .B2(n20773), .A(n13733), .ZN(P1_U2995) );
  INV_X1 U17231 ( .A(n13779), .ZN(n13791) );
  OAI22_X1 U17232 ( .A1(n13736), .A2(n13752), .B1(n9721), .B2(n13734), .ZN(
        n13735) );
  AOI21_X1 U17233 ( .B1(n13736), .B2(n13754), .A(n13735), .ZN(n20738) );
  INV_X1 U17234 ( .A(n13737), .ZN(n13739) );
  AOI21_X1 U17235 ( .B1(n13739), .B2(n20750), .A(n13738), .ZN(n13742) );
  OAI21_X1 U17236 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(P2_MORE_REG_SCAN_IN), .A(
        n13740), .ZN(n13741) );
  NAND3_X1 U17237 ( .A1(n20738), .A2(n13742), .A3(n13741), .ZN(n13790) );
  INV_X1 U17238 ( .A(n13772), .ZN(n13773) );
  NAND2_X1 U17239 ( .A1(n13744), .A2(n13743), .ZN(n13765) );
  INV_X1 U17240 ( .A(n13745), .ZN(n15122) );
  INV_X1 U17241 ( .A(n13746), .ZN(n13747) );
  NAND2_X1 U17242 ( .A1(n11732), .A2(n13747), .ZN(n13761) );
  INV_X1 U17243 ( .A(n13748), .ZN(n13750) );
  NAND2_X1 U17244 ( .A1(n13750), .A2(n13749), .ZN(n13759) );
  NAND2_X1 U17245 ( .A1(n13761), .A2(n13759), .ZN(n13751) );
  AOI21_X1 U17246 ( .B1(n13765), .B2(n15122), .A(n13751), .ZN(n13756) );
  INV_X1 U17247 ( .A(n13752), .ZN(n13753) );
  OR2_X1 U17248 ( .A1(n13754), .A2(n13753), .ZN(n13760) );
  AOI22_X1 U17249 ( .A1(n13760), .A2(n13759), .B1(n13746), .B2(n11732), .ZN(
        n13755) );
  MUX2_X1 U17250 ( .A(n13756), .B(n13755), .S(n10291), .Z(n13757) );
  NAND2_X1 U17251 ( .A1(n13757), .A2(n14917), .ZN(n13758) );
  MUX2_X1 U17252 ( .A(n10291), .B(n16437), .S(n13779), .Z(n13788) );
  AND2_X1 U17253 ( .A1(n15122), .A2(n13759), .ZN(n13766) );
  INV_X1 U17254 ( .A(n13760), .ZN(n13763) );
  OAI22_X1 U17255 ( .A1(n13763), .A2(n13766), .B1(n13762), .B2(n13761), .ZN(
        n13764) );
  AOI21_X1 U17256 ( .B1(n13766), .B2(n13765), .A(n13764), .ZN(n13767) );
  OAI21_X1 U17257 ( .B1(n15873), .B2(n13772), .A(n13767), .ZN(n16434) );
  AOI22_X1 U17258 ( .A1(n13791), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n16434), .B2(n13779), .ZN(n13787) );
  INV_X1 U17259 ( .A(n13788), .ZN(n13785) );
  NAND2_X1 U17260 ( .A1(n11732), .A2(n10230), .ZN(n13771) );
  INV_X1 U17261 ( .A(n11736), .ZN(n13768) );
  NAND2_X1 U17262 ( .A1(n13769), .A2(n13768), .ZN(n13774) );
  OAI21_X1 U17263 ( .B1(n10460), .B2(n10448), .A(n13774), .ZN(n13770) );
  OAI211_X1 U17264 ( .C1(n13259), .C2(n13772), .A(n13771), .B(n13770), .ZN(
        n16427) );
  INV_X1 U17265 ( .A(n16427), .ZN(n13778) );
  NAND2_X1 U17266 ( .A1(n19923), .A2(n13773), .ZN(n13776) );
  NAND2_X1 U17267 ( .A1(n13774), .A2(n14882), .ZN(n13775) );
  NAND2_X1 U17268 ( .A1(n13776), .A2(n13775), .ZN(n14879) );
  AOI211_X1 U17269 ( .C1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .C2(n11732), .A(
        n20732), .B(n14879), .ZN(n13777) );
  OAI21_X1 U17270 ( .B1(n13778), .B2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(
        n13777), .ZN(n13780) );
  OAI211_X1 U17271 ( .C1(n20721), .C2(n16427), .A(n13780), .B(n13779), .ZN(
        n13783) );
  OR2_X1 U17272 ( .A1(n13787), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n13782) );
  OAI21_X1 U17273 ( .B1(n10567), .B2(n13785), .A(n20710), .ZN(n13781) );
  AOI222_X1 U17274 ( .A1(n13783), .A2(n13782), .B1(n13783), .B2(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .C1(n13782), .C2(n13781), .ZN(
        n13784) );
  AOI21_X1 U17275 ( .B1(n10567), .B2(n13785), .A(n13784), .ZN(n13786) );
  OAI22_X1 U17276 ( .A1(n13788), .A2(n13787), .B1(
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(n13786), .ZN(n13789) );
  AOI211_X1 U17277 ( .C1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .C2(n13791), .A(
        n13790), .B(n13789), .ZN(n17089) );
  AOI21_X1 U17278 ( .B1(n17089), .B2(n13792), .A(n20749), .ZN(n13793) );
  INV_X1 U17279 ( .A(n13793), .ZN(n13798) );
  NAND2_X1 U17280 ( .A1(n13794), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n20747) );
  AOI21_X1 U17281 ( .B1(n13796), .B2(n13795), .A(n20747), .ZN(n13797) );
  NAND2_X1 U17282 ( .A1(n13798), .A2(n13797), .ZN(n20609) );
  INV_X1 U17283 ( .A(n17080), .ZN(n13799) );
  OAI211_X1 U17284 ( .C1(n20609), .C2(n20333), .A(n13800), .B(n13799), .ZN(
        P2_U3593) );
  OAI211_X1 U17285 ( .C1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A(n13849), .B(n13848), .ZN(n13804) );
  INV_X1 U17286 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n21202) );
  OAI22_X1 U17287 ( .A1(n20835), .A2(n20925), .B1(n21202), .B2(n16823), .ZN(
        n13801) );
  AOI21_X1 U17288 ( .B1(n13802), .B2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A(
        n13801), .ZN(n13803) );
  OAI211_X1 U17289 ( .C1(n13805), .C2(n16792), .A(n13804), .B(n13803), .ZN(
        P1_U3027) );
  INV_X1 U17290 ( .A(n20473), .ZN(n20482) );
  OAI21_X1 U17291 ( .B1(n20501), .B2(n20467), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n13812) );
  NOR2_X1 U17292 ( .A1(n13807), .A2(n13806), .ZN(n20219) );
  NAND2_X1 U17293 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n20219), .ZN(
        n13813) );
  NOR3_X1 U17294 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20710), .A3(
        n10567), .ZN(n20483) );
  INV_X1 U17295 ( .A(n20483), .ZN(n20475) );
  NOR2_X1 U17296 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20475), .ZN(
        n20465) );
  INV_X1 U17297 ( .A(n20465), .ZN(n13808) );
  AND2_X1 U17298 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n13808), .ZN(n13809) );
  NAND2_X1 U17299 ( .A1(n13810), .A2(n13809), .ZN(n13815) );
  OAI211_X1 U17300 ( .C1(n20465), .C2(n20333), .A(n13815), .B(n20512), .ZN(
        n13811) );
  INV_X1 U17301 ( .A(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n14943) );
  AOI22_X1 U17302 ( .A1(n20467), .A2(n20557), .B1(n20501), .B2(n20506), .ZN(
        n13817) );
  OAI21_X1 U17303 ( .B1(n13813), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n20607), 
        .ZN(n13814) );
  AND2_X1 U17304 ( .A1(n13815), .A2(n13814), .ZN(n20466) );
  AOI22_X1 U17305 ( .A1(n20466), .A2(n13591), .B1(n20548), .B2(n20465), .ZN(
        n13816) );
  OAI211_X1 U17306 ( .C1(n20472), .C2(n14943), .A(n13817), .B(n13816), .ZN(
        P2_U3144) );
  INV_X1 U17307 ( .A(n13818), .ZN(n13821) );
  INV_X1 U17308 ( .A(n13721), .ZN(n13820) );
  AOI21_X1 U17309 ( .B1(n13821), .B2(n13820), .A(n13819), .ZN(n20824) );
  INV_X1 U17310 ( .A(n20824), .ZN(n13826) );
  INV_X1 U17311 ( .A(n13841), .ZN(n13822) );
  AOI21_X1 U17312 ( .B1(n13824), .B2(n13823), .A(n13822), .ZN(n13851) );
  INV_X1 U17313 ( .A(n13851), .ZN(n20821) );
  OAI222_X1 U17314 ( .A1(n13826), .A2(n16640), .B1(n13825), .B2(n16644), .C1(
        n20821), .C2(n15543), .ZN(P1_U2867) );
  INV_X1 U17315 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n20891) );
  OAI222_X1 U17316 ( .A1(n13826), .A2(n15610), .B1(n15605), .B2(n13876), .C1(
        n15603), .C2(n20891), .ZN(P1_U2899) );
  INV_X1 U17317 ( .A(n13828), .ZN(n13829) );
  OAI21_X1 U17318 ( .B1(n13827), .B2(n13830), .A(n13829), .ZN(n19827) );
  INV_X1 U17319 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n19991) );
  OAI222_X1 U17320 ( .A1(n19827), .A2(n19988), .B1(n19980), .B2(n13831), .C1(
        n19991), .C2(n19979), .ZN(P2_U2904) );
  XNOR2_X1 U17321 ( .A(n13832), .B(n13833), .ZN(n13854) );
  INV_X1 U17322 ( .A(P1_REIP_REG_5__SCAN_IN), .ZN(n21205) );
  NOR2_X1 U17323 ( .A1(n16823), .A2(n21205), .ZN(n13850) );
  AOI21_X1 U17324 ( .B1(n16734), .B2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A(
        n13850), .ZN(n13834) );
  OAI21_X1 U17325 ( .B1(n20826), .B2(n16743), .A(n13834), .ZN(n13835) );
  AOI21_X1 U17326 ( .B1(n20824), .B2(n16739), .A(n13835), .ZN(n13836) );
  OAI21_X1 U17327 ( .B1(n13854), .B2(n20773), .A(n13836), .ZN(P1_U2994) );
  INV_X1 U17328 ( .A(n13837), .ZN(n13839) );
  INV_X1 U17329 ( .A(n13819), .ZN(n13838) );
  INV_X1 U17330 ( .A(n14081), .ZN(n13997) );
  AOI21_X1 U17331 ( .B1(n13839), .B2(n13838), .A(n13997), .ZN(n20809) );
  INV_X1 U17332 ( .A(n20809), .ZN(n13844) );
  INV_X1 U17333 ( .A(P1_EBX_REG_6__SCAN_IN), .ZN(n13843) );
  AND2_X1 U17334 ( .A1(n13841), .A2(n13840), .ZN(n13842) );
  OR2_X1 U17335 ( .A1(n13842), .A2(n14083), .ZN(n20802) );
  OAI222_X1 U17336 ( .A1(n13844), .A2(n16640), .B1(n13843), .B2(n16644), .C1(
        n20802), .C2(n15543), .ZN(P1_U2866) );
  INV_X1 U17337 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n20889) );
  OAI222_X1 U17338 ( .A1(n13844), .A2(n15610), .B1(n15605), .B2(n13980), .C1(
        n15603), .C2(n20889), .ZN(P1_U2898) );
  NAND2_X1 U17339 ( .A1(n15733), .A2(n15799), .ZN(n13845) );
  OAI211_X1 U17340 ( .C1(n15736), .C2(n13847), .A(n13846), .B(n13845), .ZN(
        n14354) );
  NOR2_X1 U17341 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n13848), .ZN(
        n14355) );
  AOI22_X1 U17342 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n14354), .B1(
        n14355), .B2(n13849), .ZN(n13853) );
  AOI21_X1 U17343 ( .B1(n13851), .B2(n16809), .A(n13850), .ZN(n13852) );
  OAI211_X1 U17344 ( .C1(n13854), .C2(n16792), .A(n13853), .B(n13852), .ZN(
        P1_U3026) );
  NOR2_X2 U17345 ( .A1(n14706), .A2(n16700), .ZN(n13977) );
  NOR2_X2 U17346 ( .A1(n16700), .A2(n13855), .ZN(n13978) );
  AOI22_X1 U17347 ( .A1(DATAI_16_), .A2(n13977), .B1(BUF1_REG_16__SCAN_IN), 
        .B2(n13978), .ZN(n21022) );
  NAND2_X1 U17348 ( .A1(n13892), .A2(n14088), .ZN(n21008) );
  NAND2_X1 U17349 ( .A1(n15812), .A2(n12170), .ZN(n13897) );
  OR2_X1 U17350 ( .A1(n21008), .A2(n13897), .ZN(n14232) );
  INV_X1 U17351 ( .A(n21008), .ZN(n13857) );
  NAND2_X1 U17352 ( .A1(n15812), .A2(n14398), .ZN(n14312) );
  INV_X1 U17353 ( .A(n14312), .ZN(n13896) );
  AOI22_X1 U17354 ( .A1(DATAI_24_), .A2(n13977), .B1(BUF1_REG_24__SCAN_IN), 
        .B2(n13978), .ZN(n21127) );
  INV_X1 U17355 ( .A(n21127), .ZN(n21019) );
  NOR2_X2 U17356 ( .A1(n13979), .A2(n13936), .ZN(n21115) );
  INV_X1 U17357 ( .A(n21115), .ZN(n14509) );
  NOR2_X1 U17358 ( .A1(n9734), .A2(n13860), .ZN(n21055) );
  INV_X1 U17359 ( .A(n21055), .ZN(n13862) );
  NAND2_X1 U17360 ( .A1(n13861), .A2(n12172), .ZN(n14056) );
  OAI21_X1 U17361 ( .B1(n13862), .B2(n14056), .A(n13859), .ZN(n13865) );
  INV_X1 U17362 ( .A(n13868), .ZN(n14401) );
  AOI22_X1 U17363 ( .A1(n13865), .A2(n21085), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n13868), .ZN(n14226) );
  INV_X1 U17364 ( .A(n21114), .ZN(n14617) );
  OAI22_X1 U17365 ( .A1(n14509), .A2(n13859), .B1(n14226), .B2(n14617), .ZN(
        n13864) );
  AOI21_X1 U17366 ( .B1(n14228), .B2(n21019), .A(n13864), .ZN(n13870) );
  NAND2_X1 U17367 ( .A1(n15812), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n15809) );
  INV_X1 U17368 ( .A(n13865), .ZN(n13866) );
  OAI211_X1 U17369 ( .C1(n21008), .C2(n15809), .A(n21085), .B(n13866), .ZN(
        n13867) );
  OAI211_X1 U17370 ( .C1(n21085), .C2(n13868), .A(n13867), .B(n21120), .ZN(
        n14229) );
  NAND2_X1 U17371 ( .A1(n14229), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n13869) );
  OAI211_X1 U17372 ( .C1(n21022), .C2(n14232), .A(n13870), .B(n13869), .ZN(
        P1_U3089) );
  AOI22_X1 U17373 ( .A1(DATAI_19_), .A2(n13977), .B1(BUF1_REG_19__SCAN_IN), 
        .B2(n13978), .ZN(n21034) );
  AOI22_X1 U17374 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n13978), .B1(DATAI_27_), 
        .B2(n13977), .ZN(n21145) );
  INV_X1 U17375 ( .A(n21145), .ZN(n21031) );
  NOR2_X2 U17376 ( .A1(n13979), .A2(n11178), .ZN(n21141) );
  INV_X1 U17377 ( .A(n21141), .ZN(n14513) );
  INV_X1 U17378 ( .A(n21140), .ZN(n14602) );
  OAI22_X1 U17379 ( .A1(n14513), .A2(n13859), .B1(n14226), .B2(n14602), .ZN(
        n13872) );
  AOI21_X1 U17380 ( .B1(n14228), .B2(n21031), .A(n13872), .ZN(n13874) );
  NAND2_X1 U17381 ( .A1(n14229), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n13873) );
  OAI211_X1 U17382 ( .C1(n21034), .C2(n14232), .A(n13874), .B(n13873), .ZN(
        P1_U3092) );
  AOI22_X1 U17383 ( .A1(DATAI_21_), .A2(n13977), .B1(BUF1_REG_21__SCAN_IN), 
        .B2(n13978), .ZN(n21042) );
  AOI22_X1 U17384 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n13978), .B1(DATAI_29_), 
        .B2(n13977), .ZN(n21157) );
  INV_X1 U17385 ( .A(n21157), .ZN(n21039) );
  NOR2_X2 U17386 ( .A1(n13979), .A2(n13875), .ZN(n21153) );
  INV_X1 U17387 ( .A(n21153), .ZN(n14505) );
  INV_X1 U17388 ( .A(n21152), .ZN(n14622) );
  OAI22_X1 U17389 ( .A1(n14505), .A2(n13859), .B1(n14226), .B2(n14622), .ZN(
        n13877) );
  AOI21_X1 U17390 ( .B1(n14228), .B2(n21039), .A(n13877), .ZN(n13879) );
  NAND2_X1 U17391 ( .A1(n14229), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n13878) );
  OAI211_X1 U17392 ( .C1(n21042), .C2(n14232), .A(n13879), .B(n13878), .ZN(
        P1_U3094) );
  AOI22_X1 U17393 ( .A1(DATAI_18_), .A2(n13977), .B1(BUF1_REG_18__SCAN_IN), 
        .B2(n13978), .ZN(n21030) );
  AOI22_X1 U17394 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n13978), .B1(DATAI_26_), 
        .B2(n13977), .ZN(n21139) );
  INV_X1 U17395 ( .A(n21139), .ZN(n21027) );
  NOR2_X2 U17396 ( .A1(n13979), .A2(n13880), .ZN(n21135) );
  INV_X1 U17397 ( .A(n21135), .ZN(n14501) );
  INV_X1 U17398 ( .A(n21134), .ZN(n14632) );
  OAI22_X1 U17399 ( .A1(n14501), .A2(n13859), .B1(n14226), .B2(n14632), .ZN(
        n13882) );
  AOI21_X1 U17400 ( .B1(n14228), .B2(n21027), .A(n13882), .ZN(n13884) );
  NAND2_X1 U17401 ( .A1(n14229), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n13883) );
  OAI211_X1 U17402 ( .C1(n21030), .C2(n14232), .A(n13884), .B(n13883), .ZN(
        P1_U3091) );
  AOI22_X1 U17403 ( .A1(DATAI_23_), .A2(n13977), .B1(BUF1_REG_23__SCAN_IN), 
        .B2(n13978), .ZN(n21054) );
  AOI22_X1 U17404 ( .A1(DATAI_31_), .A2(n13977), .B1(BUF1_REG_31__SCAN_IN), 
        .B2(n13978), .ZN(n21174) );
  INV_X1 U17405 ( .A(n21174), .ZN(n21049) );
  NOR2_X2 U17406 ( .A1(n13979), .A2(n14873), .ZN(n21167) );
  INV_X1 U17407 ( .A(n21167), .ZN(n14528) );
  INV_X1 U17408 ( .A(n21165), .ZN(n14607) );
  OAI22_X1 U17409 ( .A1(n14528), .A2(n13859), .B1(n14226), .B2(n14607), .ZN(
        n13885) );
  AOI21_X1 U17410 ( .B1(n14228), .B2(n21049), .A(n13885), .ZN(n13887) );
  NAND2_X1 U17411 ( .A1(n14229), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n13886) );
  OAI211_X1 U17412 ( .C1(n21054), .C2(n14232), .A(n13887), .B(n13886), .ZN(
        P1_U3096) );
  AOI22_X1 U17413 ( .A1(DATAI_17_), .A2(n13977), .B1(BUF1_REG_17__SCAN_IN), 
        .B2(n13978), .ZN(n21026) );
  AOI22_X1 U17414 ( .A1(DATAI_25_), .A2(n13977), .B1(BUF1_REG_25__SCAN_IN), 
        .B2(n13978), .ZN(n21133) );
  INV_X1 U17415 ( .A(n21133), .ZN(n21023) );
  NOR2_X2 U17416 ( .A1(n13979), .A2(n13951), .ZN(n21129) );
  INV_X1 U17417 ( .A(n21129), .ZN(n14521) );
  INV_X1 U17418 ( .A(n21128), .ZN(n14612) );
  OAI22_X1 U17419 ( .A1(n14521), .A2(n13859), .B1(n14226), .B2(n14612), .ZN(
        n13889) );
  AOI21_X1 U17420 ( .B1(n14228), .B2(n21023), .A(n13889), .ZN(n13891) );
  NAND2_X1 U17421 ( .A1(n14229), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n13890) );
  OAI211_X1 U17422 ( .C1(n21026), .C2(n14232), .A(n13891), .B(n13890), .ZN(
        P1_U3090) );
  NAND3_X1 U17423 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n20941), .ZN(n14590) );
  INV_X1 U17424 ( .A(n14590), .ZN(n13901) );
  INV_X1 U17425 ( .A(n14589), .ZN(n21086) );
  NAND2_X1 U17426 ( .A1(n14055), .A2(n9734), .ZN(n21081) );
  OR2_X1 U17427 ( .A1(n21081), .A2(n14056), .ZN(n13894) );
  INV_X1 U17428 ( .A(n14057), .ZN(n13893) );
  NAND2_X1 U17429 ( .A1(n13893), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n13898) );
  AND2_X1 U17430 ( .A1(n13894), .A2(n13898), .ZN(n13899) );
  OAI211_X1 U17431 ( .C1(n21086), .C2(n15809), .A(n21085), .B(n13899), .ZN(
        n13895) );
  OAI211_X1 U17432 ( .C1(n21085), .C2(n13901), .A(n13895), .B(n21120), .ZN(
        n13986) );
  INV_X1 U17433 ( .A(n21034), .ZN(n21142) );
  NAND2_X1 U17434 ( .A1(n14218), .A2(n21142), .ZN(n13905) );
  INV_X1 U17435 ( .A(n13898), .ZN(n13982) );
  INV_X1 U17436 ( .A(n13899), .ZN(n13900) );
  NAND2_X1 U17437 ( .A1(n13900), .A2(n21085), .ZN(n13903) );
  NAND2_X1 U17438 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n13901), .ZN(n13902) );
  NAND2_X1 U17439 ( .A1(n13903), .A2(n13902), .ZN(n13981) );
  AOI22_X1 U17440 ( .A1(n21141), .A2(n13982), .B1(n21140), .B2(n13981), .ZN(
        n13904) );
  OAI211_X1 U17441 ( .C1(n21145), .C2(n14639), .A(n13905), .B(n13904), .ZN(
        n13906) );
  AOI21_X1 U17442 ( .B1(n13986), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .A(
        n13906), .ZN(n13907) );
  INV_X1 U17443 ( .A(n13907), .ZN(P1_U3124) );
  INV_X1 U17444 ( .A(n21022), .ZN(n21124) );
  NAND2_X1 U17445 ( .A1(n14218), .A2(n21124), .ZN(n13909) );
  AOI22_X1 U17446 ( .A1(n21115), .A2(n13982), .B1(n21114), .B2(n13981), .ZN(
        n13908) );
  OAI211_X1 U17447 ( .C1(n21127), .C2(n14639), .A(n13909), .B(n13908), .ZN(
        n13910) );
  AOI21_X1 U17448 ( .B1(n13986), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A(
        n13910), .ZN(n13911) );
  INV_X1 U17449 ( .A(n13911), .ZN(P1_U3121) );
  INV_X1 U17450 ( .A(n21042), .ZN(n21154) );
  NAND2_X1 U17451 ( .A1(n14218), .A2(n21154), .ZN(n13913) );
  AOI22_X1 U17452 ( .A1(n21153), .A2(n13982), .B1(n21152), .B2(n13981), .ZN(
        n13912) );
  OAI211_X1 U17453 ( .C1(n21157), .C2(n14639), .A(n13913), .B(n13912), .ZN(
        n13914) );
  AOI21_X1 U17454 ( .B1(n13986), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .A(
        n13914), .ZN(n13915) );
  INV_X1 U17455 ( .A(n13915), .ZN(P1_U3126) );
  INV_X1 U17456 ( .A(n21026), .ZN(n21130) );
  NAND2_X1 U17457 ( .A1(n14218), .A2(n21130), .ZN(n13917) );
  AOI22_X1 U17458 ( .A1(n21129), .A2(n13982), .B1(n21128), .B2(n13981), .ZN(
        n13916) );
  OAI211_X1 U17459 ( .C1(n21133), .C2(n14639), .A(n13917), .B(n13916), .ZN(
        n13918) );
  AOI21_X1 U17460 ( .B1(n13986), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .A(
        n13918), .ZN(n13919) );
  INV_X1 U17461 ( .A(n13919), .ZN(P1_U3122) );
  INV_X1 U17462 ( .A(n21030), .ZN(n21136) );
  NAND2_X1 U17463 ( .A1(n14218), .A2(n21136), .ZN(n13921) );
  AOI22_X1 U17464 ( .A1(n21135), .A2(n13982), .B1(n21134), .B2(n13981), .ZN(
        n13920) );
  OAI211_X1 U17465 ( .C1(n21139), .C2(n14639), .A(n13921), .B(n13920), .ZN(
        n13922) );
  AOI21_X1 U17466 ( .B1(n13986), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .A(
        n13922), .ZN(n13923) );
  INV_X1 U17467 ( .A(n13923), .ZN(P1_U3123) );
  INV_X1 U17468 ( .A(n21054), .ZN(n21168) );
  NAND2_X1 U17469 ( .A1(n14218), .A2(n21168), .ZN(n13925) );
  AOI22_X1 U17470 ( .A1(n21167), .A2(n13982), .B1(n21165), .B2(n13981), .ZN(
        n13924) );
  OAI211_X1 U17471 ( .C1(n21174), .C2(n14639), .A(n13925), .B(n13924), .ZN(
        n13926) );
  AOI21_X1 U17472 ( .B1(n13986), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A(
        n13926), .ZN(n13927) );
  INV_X1 U17473 ( .A(n13927), .ZN(P1_U3128) );
  NAND2_X1 U17474 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n21291), .ZN(n16500) );
  AND2_X1 U17475 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n9954), .ZN(n13928) );
  NAND2_X1 U17476 ( .A1(n12557), .A2(n13928), .ZN(n13929) );
  OAI211_X1 U17477 ( .C1(n16500), .C2(n9954), .A(n16823), .B(n13929), .ZN(
        n13930) );
  INV_X1 U17478 ( .A(n13937), .ZN(n13932) );
  NAND2_X1 U17479 ( .A1(n13932), .A2(n13931), .ZN(n20853) );
  NAND2_X1 U17480 ( .A1(n13932), .A2(n11194), .ZN(n13934) );
  NOR2_X1 U17481 ( .A1(n13942), .A2(n16839), .ZN(n13933) );
  NAND2_X1 U17482 ( .A1(n13934), .A2(n16617), .ZN(n20855) );
  NAND2_X1 U17483 ( .A1(n13935), .A2(n20855), .ZN(n13960) );
  NAND2_X1 U17484 ( .A1(n21287), .A2(n21118), .ZN(n13949) );
  INV_X1 U17485 ( .A(n13949), .ZN(n13938) );
  AND2_X1 U17486 ( .A1(n13939), .A2(n13938), .ZN(n13945) );
  INV_X1 U17487 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n15466) );
  NOR2_X1 U17488 ( .A1(n13951), .A2(n15466), .ZN(n13940) );
  NOR2_X1 U17489 ( .A1(n13945), .A2(n13940), .ZN(n13941) );
  NAND2_X1 U17490 ( .A1(n13953), .A2(n13941), .ZN(n16622) );
  AND2_X1 U17491 ( .A1(n13942), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13943) );
  NAND2_X1 U17492 ( .A1(n16629), .A2(n13944), .ZN(n13947) );
  NOR2_X1 U17493 ( .A1(P1_REIP_REG_2__SCAN_IN), .A2(n20813), .ZN(n14833) );
  OAI21_X1 U17494 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n20813), .A(n20845), .ZN(
        n14832) );
  OAI21_X1 U17495 ( .B1(n14833), .B2(n14832), .A(P1_REIP_REG_3__SCAN_IN), .ZN(
        n13946) );
  OAI211_X1 U17496 ( .C1(n20818), .C2(n13948), .A(n13947), .B(n13946), .ZN(
        n13958) );
  NAND2_X1 U17497 ( .A1(n13949), .A2(P1_EBX_REG_31__SCAN_IN), .ZN(n13950) );
  NOR2_X1 U17498 ( .A1(n13951), .A2(n13950), .ZN(n13952) );
  INV_X1 U17499 ( .A(n13954), .ZN(n13956) );
  INV_X1 U17500 ( .A(n20813), .ZN(n20857) );
  NAND4_X1 U17501 ( .A1(n20857), .A2(n21200), .A3(P1_REIP_REG_1__SCAN_IN), 
        .A4(P1_REIP_REG_2__SCAN_IN), .ZN(n13955) );
  OAI21_X1 U17502 ( .B1(n20860), .B2(n13956), .A(n13955), .ZN(n13957) );
  AOI211_X1 U17503 ( .C1(n20850), .C2(P1_EBX_REG_3__SCAN_IN), .A(n13958), .B(
        n13957), .ZN(n13959) );
  OAI211_X1 U17504 ( .C1(n15819), .C2(n20853), .A(n13960), .B(n13959), .ZN(
        P1_U2837) );
  OAI21_X1 U17505 ( .B1(n20286), .B2(n20327), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n13963) );
  NAND3_X1 U17506 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n10567), .A3(
        n20721), .ZN(n20254) );
  NOR2_X1 U17507 ( .A1(n20732), .A2(n20254), .ZN(n20271) );
  NOR2_X1 U17508 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n20545), .ZN(
        n20298) );
  INV_X1 U17509 ( .A(n20298), .ZN(n20307) );
  NOR2_X1 U17510 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20307), .ZN(
        n20291) );
  NOR2_X1 U17511 ( .A1(n20271), .A2(n20291), .ZN(n13965) );
  AOI211_X1 U17512 ( .C1(n13963), .C2(n13965), .A(n20551), .B(n13962), .ZN(
        n20277) );
  OAI21_X1 U17513 ( .B1(n9763), .B2(n20291), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n13964) );
  OAI21_X1 U17514 ( .B1(n13965), .B2(n20509), .A(n13964), .ZN(n20292) );
  INV_X1 U17515 ( .A(n20548), .ZN(n13968) );
  INV_X1 U17516 ( .A(n20291), .ZN(n13967) );
  AOI22_X1 U17517 ( .A1(n20286), .A2(n20557), .B1(n20327), .B2(n20506), .ZN(
        n13966) );
  OAI21_X1 U17518 ( .B1(n13968), .B2(n13967), .A(n13966), .ZN(n13969) );
  AOI21_X1 U17519 ( .B1(n20292), .B2(n13591), .A(n13969), .ZN(n13970) );
  OAI21_X1 U17520 ( .B1(n20277), .B2(n13971), .A(n13970), .ZN(P2_U3096) );
  AOI22_X1 U17521 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n13978), .B1(DATAI_28_), 
        .B2(n13977), .ZN(n21151) );
  AOI22_X1 U17522 ( .A1(DATAI_20_), .A2(n13977), .B1(BUF1_REG_20__SCAN_IN), 
        .B2(n13978), .ZN(n21038) );
  INV_X1 U17523 ( .A(n21038), .ZN(n21148) );
  NAND2_X1 U17524 ( .A1(n14218), .A2(n21148), .ZN(n13974) );
  NOR2_X2 U17525 ( .A1(n13979), .A2(n11129), .ZN(n21147) );
  AOI22_X1 U17526 ( .A1(n21147), .A2(n13982), .B1(n21146), .B2(n13981), .ZN(
        n13973) );
  OAI211_X1 U17527 ( .C1(n21151), .C2(n14639), .A(n13974), .B(n13973), .ZN(
        n13975) );
  AOI21_X1 U17528 ( .B1(n13986), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A(
        n13975), .ZN(n13976) );
  INV_X1 U17529 ( .A(n13976), .ZN(P1_U3125) );
  AOI22_X1 U17530 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n13978), .B1(DATAI_30_), 
        .B2(n13977), .ZN(n21163) );
  AOI22_X1 U17531 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n13978), .B1(DATAI_22_), 
        .B2(n13977), .ZN(n21046) );
  INV_X1 U17532 ( .A(n21046), .ZN(n21160) );
  NAND2_X1 U17533 ( .A1(n14218), .A2(n21160), .ZN(n13984) );
  NOR2_X2 U17534 ( .A1(n13979), .A2(n11199), .ZN(n21159) );
  AOI22_X1 U17535 ( .A1(n21159), .A2(n13982), .B1(n21158), .B2(n13981), .ZN(
        n13983) );
  OAI211_X1 U17536 ( .C1(n21163), .C2(n14639), .A(n13984), .B(n13983), .ZN(
        n13985) );
  AOI21_X1 U17537 ( .B1(n13986), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A(
        n13985), .ZN(n13987) );
  INV_X1 U17538 ( .A(n13987), .ZN(P1_U3127) );
  OAI21_X1 U17539 ( .B1(n13988), .B2(n13990), .A(n13989), .ZN(n14651) );
  INV_X1 U17540 ( .A(n15605), .ZN(n15608) );
  AOI22_X1 U17541 ( .A1(n15608), .A2(n15561), .B1(P1_EAX_REG_9__SCAN_IN), .B2(
        n15606), .ZN(n13991) );
  OAI21_X1 U17542 ( .B1(n14651), .B2(n15610), .A(n13991), .ZN(P1_U2895) );
  INV_X1 U17543 ( .A(n14121), .ZN(n13993) );
  OAI21_X1 U17544 ( .B1(n13993), .B2(n10143), .A(n14293), .ZN(n14046) );
  INV_X1 U17545 ( .A(n14046), .ZN(n16810) );
  AOI22_X1 U17546 ( .A1(n16810), .A2(n15528), .B1(P1_EBX_REG_9__SCAN_IN), .B2(
        n15527), .ZN(n13994) );
  OAI21_X1 U17547 ( .B1(n14651), .B2(n16640), .A(n13994), .ZN(P1_U2863) );
  AOI21_X1 U17548 ( .B1(n13997), .B2(n13995), .A(n13996), .ZN(n13998) );
  NOR2_X1 U17549 ( .A1(n13998), .A2(n13988), .ZN(n14364) );
  INV_X1 U17550 ( .A(n14364), .ZN(n14235) );
  MUX2_X1 U17551 ( .A(DATAI_8_), .B(BUF1_REG_8__SCAN_IN), .S(n14706), .Z(
        n20905) );
  INV_X1 U17552 ( .A(n20905), .ZN(n13999) );
  OAI222_X1 U17553 ( .A1(n14235), .A2(n15610), .B1(n15605), .B2(n13999), .C1(
        n20885), .C2(n15603), .ZN(P1_U2896) );
  NAND3_X1 U17554 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n20941), .A3(
        n21009), .ZN(n21083) );
  NOR2_X1 U17555 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21083), .ZN(
        n14039) );
  INV_X1 U17556 ( .A(n14095), .ZN(n14000) );
  NAND2_X1 U17557 ( .A1(n14007), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n21012) );
  NAND2_X1 U17558 ( .A1(n14000), .A2(n21012), .ZN(n14594) );
  INV_X1 U17559 ( .A(n14594), .ZN(n20952) );
  AOI21_X1 U17560 ( .B1(n21109), .B2(n14232), .A(n21118), .ZN(n14004) );
  INV_X1 U17561 ( .A(n14001), .ZN(n20945) );
  OR2_X1 U17562 ( .A1(n21081), .A2(n20945), .ZN(n14003) );
  INV_X1 U17563 ( .A(n14039), .ZN(n14002) );
  NAND2_X1 U17564 ( .A1(n14003), .A2(n14002), .ZN(n14006) );
  OR2_X1 U17565 ( .A1(n14004), .A2(n14006), .ZN(n14005) );
  OAI211_X1 U17566 ( .C1(n14039), .C2(n20953), .A(n20952), .B(n14005), .ZN(
        n14044) );
  NAND2_X1 U17567 ( .A1(n14006), .A2(n21085), .ZN(n14009) );
  INV_X1 U17568 ( .A(n14491), .ZN(n20949) );
  NAND2_X1 U17569 ( .A1(n20949), .A2(n20947), .ZN(n14096) );
  INV_X1 U17570 ( .A(n14096), .ZN(n14092) );
  NOR2_X1 U17571 ( .A1(n14007), .A2(n21113), .ZN(n20954) );
  NAND2_X1 U17572 ( .A1(n14092), .A2(n20954), .ZN(n14008) );
  NAND2_X1 U17573 ( .A1(n14009), .A2(n14008), .ZN(n14038) );
  AOI22_X1 U17574 ( .A1(n21115), .A2(n14039), .B1(n21114), .B2(n14038), .ZN(
        n14011) );
  INV_X1 U17575 ( .A(n14232), .ZN(n14040) );
  NAND2_X1 U17576 ( .A1(n14040), .A2(n21019), .ZN(n14010) );
  OAI211_X1 U17577 ( .C1(n21109), .C2(n21022), .A(n14011), .B(n14010), .ZN(
        n14012) );
  AOI21_X1 U17578 ( .B1(n14044), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A(
        n14012), .ZN(n14013) );
  INV_X1 U17579 ( .A(n14013), .ZN(P1_U3097) );
  AOI22_X1 U17580 ( .A1(n21167), .A2(n14039), .B1(n21165), .B2(n14038), .ZN(
        n14015) );
  NAND2_X1 U17581 ( .A1(n14040), .A2(n21049), .ZN(n14014) );
  OAI211_X1 U17582 ( .C1(n21109), .C2(n21054), .A(n14015), .B(n14014), .ZN(
        n14016) );
  AOI21_X1 U17583 ( .B1(n14044), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .A(
        n14016), .ZN(n14017) );
  INV_X1 U17584 ( .A(n14017), .ZN(P1_U3104) );
  AOI22_X1 U17585 ( .A1(n21135), .A2(n14039), .B1(n21134), .B2(n14038), .ZN(
        n14019) );
  NAND2_X1 U17586 ( .A1(n14040), .A2(n21027), .ZN(n14018) );
  OAI211_X1 U17587 ( .C1(n21109), .C2(n21030), .A(n14019), .B(n14018), .ZN(
        n14020) );
  AOI21_X1 U17588 ( .B1(n14044), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .A(
        n14020), .ZN(n14021) );
  INV_X1 U17589 ( .A(n14021), .ZN(P1_U3099) );
  AOI22_X1 U17590 ( .A1(n21129), .A2(n14039), .B1(n21128), .B2(n14038), .ZN(
        n14023) );
  NAND2_X1 U17591 ( .A1(n14040), .A2(n21023), .ZN(n14022) );
  OAI211_X1 U17592 ( .C1(n21109), .C2(n21026), .A(n14023), .B(n14022), .ZN(
        n14024) );
  AOI21_X1 U17593 ( .B1(n14044), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .A(
        n14024), .ZN(n14025) );
  INV_X1 U17594 ( .A(n14025), .ZN(P1_U3098) );
  AOI22_X1 U17595 ( .A1(n21153), .A2(n14039), .B1(n21152), .B2(n14038), .ZN(
        n14027) );
  NAND2_X1 U17596 ( .A1(n14040), .A2(n21039), .ZN(n14026) );
  OAI211_X1 U17597 ( .C1(n21109), .C2(n21042), .A(n14027), .B(n14026), .ZN(
        n14028) );
  AOI21_X1 U17598 ( .B1(n14044), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .A(
        n14028), .ZN(n14029) );
  INV_X1 U17599 ( .A(n14029), .ZN(P1_U3102) );
  AOI22_X1 U17600 ( .A1(n21147), .A2(n14039), .B1(n21146), .B2(n14038), .ZN(
        n14031) );
  INV_X1 U17601 ( .A(n21151), .ZN(n21035) );
  NAND2_X1 U17602 ( .A1(n14040), .A2(n21035), .ZN(n14030) );
  OAI211_X1 U17603 ( .C1(n21109), .C2(n21038), .A(n14031), .B(n14030), .ZN(
        n14032) );
  AOI21_X1 U17604 ( .B1(n14044), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A(
        n14032), .ZN(n14033) );
  INV_X1 U17605 ( .A(n14033), .ZN(P1_U3101) );
  AOI22_X1 U17606 ( .A1(n21159), .A2(n14039), .B1(n21158), .B2(n14038), .ZN(
        n14035) );
  INV_X1 U17607 ( .A(n21163), .ZN(n21043) );
  NAND2_X1 U17608 ( .A1(n14040), .A2(n21043), .ZN(n14034) );
  OAI211_X1 U17609 ( .C1(n21109), .C2(n21046), .A(n14035), .B(n14034), .ZN(
        n14036) );
  AOI21_X1 U17610 ( .B1(n14044), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .A(
        n14036), .ZN(n14037) );
  INV_X1 U17611 ( .A(n14037), .ZN(P1_U3103) );
  AOI22_X1 U17612 ( .A1(n21141), .A2(n14039), .B1(n21140), .B2(n14038), .ZN(
        n14042) );
  NAND2_X1 U17613 ( .A1(n14040), .A2(n21031), .ZN(n14041) );
  OAI211_X1 U17614 ( .C1(n21109), .C2(n21034), .A(n14042), .B(n14041), .ZN(
        n14043) );
  AOI21_X1 U17615 ( .B1(n14044), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .A(
        n14043), .ZN(n14045) );
  INV_X1 U17616 ( .A(n14045), .ZN(P1_U3100) );
  NAND4_X1 U17617 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_2__SCAN_IN), 
        .A3(P1_REIP_REG_3__SCAN_IN), .A4(P1_REIP_REG_4__SCAN_IN), .ZN(n20827)
         );
  INV_X1 U17618 ( .A(P1_REIP_REG_6__SCAN_IN), .ZN(n21206) );
  NOR3_X1 U17619 ( .A1(n20827), .A2(n21206), .A3(n21205), .ZN(n20792) );
  NAND3_X1 U17620 ( .A1(n20792), .A2(P1_REIP_REG_7__SCAN_IN), .A3(
        P1_REIP_REG_8__SCAN_IN), .ZN(n14712) );
  NOR2_X1 U17621 ( .A1(n20813), .A2(n14712), .ZN(n14654) );
  INV_X1 U17622 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n21213) );
  OAI22_X1 U17623 ( .A1(n14046), .A2(n20860), .B1(n14647), .B2(n20847), .ZN(
        n14052) );
  INV_X1 U17624 ( .A(n20845), .ZN(n20805) );
  NOR2_X1 U17625 ( .A1(n20805), .A2(n14712), .ZN(n14670) );
  NAND2_X1 U17626 ( .A1(n20813), .A2(n20845), .ZN(n15461) );
  NAND2_X1 U17627 ( .A1(n15461), .A2(P1_REIP_REG_9__SCAN_IN), .ZN(n14047) );
  OAI22_X1 U17628 ( .A1(n14670), .A2(n14047), .B1(n16622), .B2(n11619), .ZN(
        n14048) );
  INV_X1 U17629 ( .A(n14048), .ZN(n14050) );
  NAND2_X1 U17630 ( .A1(n20845), .A2(n14049), .ZN(n20816) );
  OAI211_X1 U17631 ( .C1(n20818), .C2(n12230), .A(n14050), .B(n20816), .ZN(
        n14051) );
  AOI211_X1 U17632 ( .C1(n14654), .C2(n21213), .A(n14052), .B(n14051), .ZN(
        n14053) );
  OAI21_X1 U17633 ( .B1(n16617), .B2(n14651), .A(n14053), .ZN(P1_U2831) );
  INV_X1 U17634 ( .A(n9734), .ZN(n14054) );
  OR2_X1 U17635 ( .A1(n14055), .A2(n14054), .ZN(n20946) );
  INV_X1 U17636 ( .A(n20946), .ZN(n20979) );
  INV_X1 U17637 ( .A(n14056), .ZN(n14316) );
  NOR2_X1 U17638 ( .A1(n14057), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n14078) );
  AOI21_X1 U17639 ( .B1(n20979), .B2(n14316), .A(n14078), .ZN(n14060) );
  INV_X1 U17640 ( .A(n15809), .ZN(n14317) );
  AOI21_X1 U17641 ( .B1(n20940), .B2(n14317), .A(n21122), .ZN(n14059) );
  NAND3_X1 U17642 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n21010), .A3(
        n20941), .ZN(n14536) );
  AOI22_X1 U17643 ( .A1(n14060), .A2(n14059), .B1(n21122), .B2(n14536), .ZN(
        n14058) );
  NAND2_X1 U17644 ( .A1(n21120), .A2(n14058), .ZN(n14077) );
  INV_X1 U17645 ( .A(n14059), .ZN(n14061) );
  OAI22_X1 U17646 ( .A1(n14061), .A2(n14060), .B1(n21113), .B2(n14536), .ZN(
        n14076) );
  AOI22_X1 U17647 ( .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n14077), .B1(
        n21140), .B2(n14076), .ZN(n14063) );
  AOI22_X1 U17648 ( .A1(n14533), .A2(n21031), .B1(n14078), .B2(n21141), .ZN(
        n14062) );
  OAI211_X1 U17649 ( .C1(n21034), .C2(n21018), .A(n14063), .B(n14062), .ZN(
        P1_U3060) );
  AOI22_X1 U17650 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n14077), .B1(
        n21114), .B2(n14076), .ZN(n14065) );
  AOI22_X1 U17651 ( .A1(n14533), .A2(n21019), .B1(n14078), .B2(n21115), .ZN(
        n14064) );
  OAI211_X1 U17652 ( .C1(n21022), .C2(n21018), .A(n14065), .B(n14064), .ZN(
        P1_U3057) );
  AOI22_X1 U17653 ( .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n14077), .B1(
        n21152), .B2(n14076), .ZN(n14067) );
  AOI22_X1 U17654 ( .A1(n14533), .A2(n21039), .B1(n14078), .B2(n21153), .ZN(
        n14066) );
  OAI211_X1 U17655 ( .C1(n21042), .C2(n21018), .A(n14067), .B(n14066), .ZN(
        P1_U3062) );
  AOI22_X1 U17656 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n14077), .B1(
        n21146), .B2(n14076), .ZN(n14069) );
  AOI22_X1 U17657 ( .A1(n14533), .A2(n21035), .B1(n14078), .B2(n21147), .ZN(
        n14068) );
  OAI211_X1 U17658 ( .C1(n21038), .C2(n21018), .A(n14069), .B(n14068), .ZN(
        P1_U3061) );
  AOI22_X1 U17659 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n14077), .B1(
        n21158), .B2(n14076), .ZN(n14071) );
  AOI22_X1 U17660 ( .A1(n14533), .A2(n21043), .B1(n14078), .B2(n21159), .ZN(
        n14070) );
  OAI211_X1 U17661 ( .C1(n21046), .C2(n21018), .A(n14071), .B(n14070), .ZN(
        P1_U3063) );
  AOI22_X1 U17662 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n14077), .B1(
        n21165), .B2(n14076), .ZN(n14073) );
  AOI22_X1 U17663 ( .A1(n14533), .A2(n21049), .B1(n14078), .B2(n21167), .ZN(
        n14072) );
  OAI211_X1 U17664 ( .C1(n21054), .C2(n21018), .A(n14073), .B(n14072), .ZN(
        P1_U3064) );
  AOI22_X1 U17665 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n14077), .B1(
        n21134), .B2(n14076), .ZN(n14075) );
  AOI22_X1 U17666 ( .A1(n14533), .A2(n21027), .B1(n14078), .B2(n21135), .ZN(
        n14074) );
  OAI211_X1 U17667 ( .C1(n21030), .C2(n21018), .A(n14075), .B(n14074), .ZN(
        P1_U3059) );
  AOI22_X1 U17668 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n14077), .B1(
        n21128), .B2(n14076), .ZN(n14080) );
  AOI22_X1 U17669 ( .A1(n14533), .A2(n21023), .B1(n14078), .B2(n21129), .ZN(
        n14079) );
  OAI211_X1 U17670 ( .C1(n21026), .C2(n21018), .A(n14080), .B(n14079), .ZN(
        P1_U3058) );
  XNOR2_X1 U17671 ( .A(n14081), .B(n13995), .ZN(n20797) );
  NOR2_X1 U17672 ( .A1(n14083), .A2(n14082), .ZN(n14084) );
  OR2_X1 U17673 ( .A1(n14119), .A2(n14084), .ZN(n20795) );
  OAI22_X1 U17674 ( .A1(n20795), .A2(n15543), .B1(n14085), .B2(n16644), .ZN(
        n14086) );
  AOI21_X1 U17675 ( .B1(n20797), .B2(n15545), .A(n14086), .ZN(n14087) );
  INV_X1 U17676 ( .A(n14087), .ZN(P1_U2865) );
  INV_X1 U17677 ( .A(n21173), .ZN(n14089) );
  OAI21_X1 U17678 ( .B1(n14218), .B2(n14089), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n14090) );
  NAND2_X1 U17679 ( .A1(n14090), .A2(n21085), .ZN(n14099) );
  INV_X1 U17680 ( .A(n14099), .ZN(n14093) );
  OR2_X1 U17681 ( .A1(n9734), .A2(n14091), .ZN(n14314) );
  NOR2_X1 U17682 ( .A1(n14314), .A2(n20945), .ZN(n14098) );
  INV_X1 U17683 ( .A(n21012), .ZN(n14400) );
  AOI22_X1 U17684 ( .A1(n14093), .A2(n14098), .B1(n14092), .B2(n14400), .ZN(
        n14222) );
  NAND3_X1 U17685 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n21009), .ZN(n21116) );
  OR2_X1 U17686 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21116), .ZN(
        n14216) );
  OAI22_X1 U17687 ( .A1(n14509), .A2(n14216), .B1(n21022), .B2(n21173), .ZN(
        n14094) );
  AOI21_X1 U17688 ( .B1(n14218), .B2(n21019), .A(n14094), .ZN(n14101) );
  AOI22_X1 U17689 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n14096), .B1(
        P1_STATE2_REG_3__SCAN_IN), .B2(n14216), .ZN(n14097) );
  OAI211_X1 U17690 ( .C1(n14099), .C2(n14098), .A(n21016), .B(n14097), .ZN(
        n14219) );
  NAND2_X1 U17691 ( .A1(n14219), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n14100) );
  OAI211_X1 U17692 ( .C1(n14222), .C2(n14617), .A(n14101), .B(n14100), .ZN(
        P1_U3129) );
  OAI22_X1 U17693 ( .A1(n14521), .A2(n14216), .B1(n21026), .B2(n21173), .ZN(
        n14102) );
  AOI21_X1 U17694 ( .B1(n14218), .B2(n21023), .A(n14102), .ZN(n14104) );
  NAND2_X1 U17695 ( .A1(n14219), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n14103) );
  OAI211_X1 U17696 ( .C1(n14222), .C2(n14612), .A(n14104), .B(n14103), .ZN(
        P1_U3130) );
  OAI22_X1 U17697 ( .A1(n14528), .A2(n14216), .B1(n21054), .B2(n21173), .ZN(
        n14105) );
  AOI21_X1 U17698 ( .B1(n14218), .B2(n21049), .A(n14105), .ZN(n14107) );
  NAND2_X1 U17699 ( .A1(n14219), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n14106) );
  OAI211_X1 U17700 ( .C1(n14222), .C2(n14607), .A(n14107), .B(n14106), .ZN(
        P1_U3136) );
  OAI22_X1 U17701 ( .A1(n14505), .A2(n14216), .B1(n21042), .B2(n21173), .ZN(
        n14108) );
  AOI21_X1 U17702 ( .B1(n14218), .B2(n21039), .A(n14108), .ZN(n14110) );
  NAND2_X1 U17703 ( .A1(n14219), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n14109) );
  OAI211_X1 U17704 ( .C1(n14222), .C2(n14622), .A(n14110), .B(n14109), .ZN(
        P1_U3134) );
  OAI22_X1 U17705 ( .A1(n14501), .A2(n14216), .B1(n21030), .B2(n21173), .ZN(
        n14111) );
  AOI21_X1 U17706 ( .B1(n14218), .B2(n21027), .A(n14111), .ZN(n14113) );
  NAND2_X1 U17707 ( .A1(n14219), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(
        n14112) );
  OAI211_X1 U17708 ( .C1(n14222), .C2(n14632), .A(n14113), .B(n14112), .ZN(
        P1_U3131) );
  OAI22_X1 U17709 ( .A1(n14513), .A2(n14216), .B1(n21034), .B2(n21173), .ZN(
        n14114) );
  AOI21_X1 U17710 ( .B1(n14218), .B2(n21031), .A(n14114), .ZN(n14116) );
  NAND2_X1 U17711 ( .A1(n14219), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(
        n14115) );
  OAI211_X1 U17712 ( .C1(n14222), .C2(n14602), .A(n14116), .B(n14115), .ZN(
        P1_U3132) );
  NAND2_X1 U17713 ( .A1(n20849), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n14117) );
  OAI211_X1 U17714 ( .C1(n20847), .C2(n14362), .A(n20816), .B(n14117), .ZN(
        n14123) );
  OR2_X1 U17715 ( .A1(n14119), .A2(n14118), .ZN(n14120) );
  NAND2_X1 U17716 ( .A1(n14121), .A2(n14120), .ZN(n14356) );
  NOR2_X1 U17717 ( .A1(n14356), .A2(n20860), .ZN(n14122) );
  AOI211_X1 U17718 ( .C1(n20850), .C2(P1_EBX_REG_8__SCAN_IN), .A(n14123), .B(
        n14122), .ZN(n14127) );
  INV_X1 U17719 ( .A(P1_REIP_REG_7__SCAN_IN), .ZN(n21208) );
  NAND2_X1 U17720 ( .A1(n20857), .A2(n20792), .ZN(n20789) );
  INV_X1 U17721 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n21210) );
  OAI21_X1 U17722 ( .B1(n21208), .B2(n20789), .A(n21210), .ZN(n14125) );
  INV_X1 U17723 ( .A(n14670), .ZN(n14124) );
  NAND3_X1 U17724 ( .A1(n14125), .A2(n15461), .A3(n14124), .ZN(n14126) );
  OAI211_X1 U17725 ( .C1(n14235), .C2(n16617), .A(n14127), .B(n14126), .ZN(
        P1_U2832) );
  OR2_X1 U17726 ( .A1(n14129), .A2(n14130), .ZN(n14131) );
  NAND2_X1 U17727 ( .A1(n14128), .A2(n14131), .ZN(n19787) );
  NAND2_X1 U17728 ( .A1(n10631), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(
        n14135) );
  NAND2_X1 U17729 ( .A1(n14951), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(
        n14134) );
  AOI22_X1 U17730 ( .A1(n10500), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n14885), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n14133) );
  NAND2_X1 U17731 ( .A1(n10507), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n14132) );
  NAND4_X1 U17732 ( .A1(n14135), .A2(n14134), .A3(n14133), .A4(n14132), .ZN(
        n14141) );
  AOI22_X1 U17733 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n10498), .B1(
        n10499), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n14139) );
  NAND2_X1 U17734 ( .A1(n14908), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n14138) );
  NAND2_X1 U17735 ( .A1(n14909), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n14137) );
  NAND2_X1 U17736 ( .A1(n14910), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n14136) );
  NAND4_X1 U17737 ( .A1(n14139), .A2(n14138), .A3(n14137), .A4(n14136), .ZN(
        n14140) );
  NOR2_X1 U17738 ( .A1(n14141), .A2(n14140), .ZN(n14150) );
  OAI22_X1 U17739 ( .A1(n14919), .A2(n14143), .B1(n14917), .B2(n14142), .ZN(
        n14148) );
  INV_X1 U17740 ( .A(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n14146) );
  AOI22_X1 U17741 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n14967), .B1(
        n11881), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n14145) );
  NAND2_X1 U17742 ( .A1(n14450), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n14144) );
  OAI211_X1 U17743 ( .C1(n14473), .C2(n14146), .A(n14145), .B(n14144), .ZN(
        n14147) );
  NOR2_X1 U17744 ( .A1(n14148), .A2(n14147), .ZN(n14149) );
  AND2_X1 U17745 ( .A1(n14150), .A2(n14149), .ZN(n14194) );
  NAND2_X1 U17746 ( .A1(n10631), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n14154) );
  NAND2_X1 U17747 ( .A1(n14951), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n14153) );
  AOI22_X1 U17748 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n10500), .B1(
        n14885), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n14152) );
  NAND2_X1 U17749 ( .A1(n10507), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n14151) );
  AND4_X1 U17750 ( .A1(n14154), .A2(n14153), .A3(n14152), .A4(n14151), .ZN(
        n14169) );
  AOI22_X1 U17751 ( .A1(n14957), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n14956), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n14168) );
  NAND2_X1 U17752 ( .A1(n10499), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n14156) );
  NAND2_X1 U17753 ( .A1(n10498), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n14155) );
  OAI211_X1 U17754 ( .C1(n14961), .C2(n14157), .A(n14156), .B(n14155), .ZN(
        n14161) );
  OAI22_X1 U17755 ( .A1(n14964), .A2(n14159), .B1(n14962), .B2(n14158), .ZN(
        n14160) );
  NOR2_X1 U17756 ( .A1(n14161), .A2(n14160), .ZN(n14167) );
  AOI22_X1 U17757 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n14967), .B1(
        n11881), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n14163) );
  NAND2_X1 U17758 ( .A1(n14450), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n14162) );
  OAI211_X1 U17759 ( .C1(n14473), .C2(n14164), .A(n14163), .B(n14162), .ZN(
        n14165) );
  INV_X1 U17760 ( .A(n14165), .ZN(n14166) );
  NAND4_X1 U17761 ( .A1(n14169), .A2(n14168), .A3(n14167), .A4(n14166), .ZN(
        n14368) );
  NAND2_X1 U17762 ( .A1(n10631), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n14173) );
  NAND2_X1 U17763 ( .A1(n14951), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n14172) );
  AOI22_X1 U17764 ( .A1(n10500), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n14885), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n14171) );
  NAND2_X1 U17765 ( .A1(n10507), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n14170) );
  AND4_X1 U17766 ( .A1(n14173), .A2(n14172), .A3(n14171), .A4(n14170), .ZN(
        n14187) );
  AOI22_X1 U17767 ( .A1(n14957), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n14956), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n14186) );
  INV_X1 U17768 ( .A(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n14176) );
  NAND2_X1 U17769 ( .A1(n10499), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n14175) );
  NAND2_X1 U17770 ( .A1(n10498), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n14174) );
  OAI211_X1 U17771 ( .C1(n14961), .C2(n14176), .A(n14175), .B(n14174), .ZN(
        n14179) );
  OAI22_X1 U17772 ( .A1(n14964), .A2(n11802), .B1(n14962), .B2(n14177), .ZN(
        n14178) );
  NOR2_X1 U17773 ( .A1(n14179), .A2(n14178), .ZN(n14185) );
  AOI22_X1 U17774 ( .A1(n14967), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n11881), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n14181) );
  NAND2_X1 U17775 ( .A1(n14450), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n14180) );
  OAI211_X1 U17776 ( .C1(n14182), .C2(n14473), .A(n14181), .B(n14180), .ZN(
        n14183) );
  INV_X1 U17777 ( .A(n14183), .ZN(n14184) );
  NAND4_X1 U17778 ( .A1(n14187), .A2(n14186), .A3(n14185), .A4(n14184), .ZN(
        n14253) );
  INV_X1 U17779 ( .A(n14253), .ZN(n14188) );
  OR2_X1 U17780 ( .A1(n19937), .A2(n19934), .ZN(n14249) );
  NOR2_X1 U17781 ( .A1(n14188), .A2(n14249), .ZN(n14250) );
  NAND2_X1 U17782 ( .A1(n14368), .A2(n14250), .ZN(n14189) );
  NOR2_X1 U17783 ( .A1(n14190), .A2(n14189), .ZN(n14192) );
  NAND2_X1 U17784 ( .A1(n19960), .A2(n14192), .ZN(n14367) );
  INV_X1 U17785 ( .A(n14194), .ZN(n14191) );
  AND2_X1 U17786 ( .A1(n14192), .A2(n14191), .ZN(n14479) );
  NAND2_X1 U17787 ( .A1(n19960), .A2(n14479), .ZN(n16017) );
  INV_X1 U17788 ( .A(n16017), .ZN(n14193) );
  AOI21_X1 U17789 ( .B1(n14194), .B2(n14367), .A(n14193), .ZN(n14577) );
  NAND2_X1 U17790 ( .A1(n14577), .A2(n16926), .ZN(n14196) );
  NAND2_X1 U17791 ( .A1(n19947), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n14195) );
  OAI211_X1 U17792 ( .C1(n19787), .C2(n19947), .A(n14196), .B(n14195), .ZN(
        P2_U2869) );
  NOR2_X1 U17793 ( .A1(n9766), .A2(n14198), .ZN(n14199) );
  XNOR2_X1 U17794 ( .A(n14199), .B(n16188), .ZN(n14203) );
  NAND2_X1 U17795 ( .A1(n14200), .A2(n13397), .ZN(n14202) );
  AND2_X1 U17796 ( .A1(n14202), .A2(n14201), .ZN(n17047) );
  AOI22_X1 U17797 ( .A1(n19897), .A2(n14203), .B1(n19915), .B2(n17047), .ZN(
        n14212) );
  INV_X1 U17798 ( .A(n19919), .ZN(n19877) );
  NAND3_X1 U17799 ( .A1(n14205), .A2(n14204), .A3(n12107), .ZN(n14206) );
  NAND2_X1 U17800 ( .A1(n14207), .A2(n14206), .ZN(n19917) );
  AOI22_X1 U17801 ( .A1(n14208), .A2(n19877), .B1(P2_EBX_REG_8__SCAN_IN), .B2(
        n19917), .ZN(n14209) );
  INV_X1 U17802 ( .A(n19905), .ZN(n20073) );
  OAI211_X1 U17803 ( .C1(n10945), .C2(n19887), .A(n14209), .B(n20073), .ZN(
        n14210) );
  AOI21_X1 U17804 ( .B1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n19929), .A(
        n14210), .ZN(n14211) );
  OAI211_X1 U17805 ( .C1(n16190), .C2(n19880), .A(n14212), .B(n14211), .ZN(
        P2_U2847) );
  INV_X1 U17806 ( .A(n21158), .ZN(n14640) );
  INV_X1 U17807 ( .A(n21159), .ZN(n14497) );
  OAI22_X1 U17808 ( .A1(n14497), .A2(n14216), .B1(n21046), .B2(n21173), .ZN(
        n14213) );
  AOI21_X1 U17809 ( .B1(n14218), .B2(n21043), .A(n14213), .ZN(n14215) );
  NAND2_X1 U17810 ( .A1(n14219), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n14214) );
  OAI211_X1 U17811 ( .C1(n14222), .C2(n14640), .A(n14215), .B(n14214), .ZN(
        P1_U3135) );
  INV_X1 U17812 ( .A(n21146), .ZN(n14627) );
  INV_X1 U17813 ( .A(n21147), .ZN(n14517) );
  OAI22_X1 U17814 ( .A1(n14517), .A2(n14216), .B1(n21038), .B2(n21173), .ZN(
        n14217) );
  AOI21_X1 U17815 ( .B1(n14218), .B2(n21035), .A(n14217), .ZN(n14221) );
  NAND2_X1 U17816 ( .A1(n14219), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n14220) );
  OAI211_X1 U17817 ( .C1(n14222), .C2(n14627), .A(n14221), .B(n14220), .ZN(
        P1_U3133) );
  OAI22_X1 U17818 ( .A1(n14497), .A2(n13859), .B1(n14226), .B2(n14640), .ZN(
        n14223) );
  AOI21_X1 U17819 ( .B1(n14228), .B2(n21043), .A(n14223), .ZN(n14225) );
  NAND2_X1 U17820 ( .A1(n14229), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n14224) );
  OAI211_X1 U17821 ( .C1(n21046), .C2(n14232), .A(n14225), .B(n14224), .ZN(
        P1_U3095) );
  OAI22_X1 U17822 ( .A1(n14517), .A2(n13859), .B1(n14226), .B2(n14627), .ZN(
        n14227) );
  AOI21_X1 U17823 ( .B1(n14228), .B2(n21035), .A(n14227), .ZN(n14231) );
  NAND2_X1 U17824 ( .A1(n14229), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n14230) );
  OAI211_X1 U17825 ( .C1(n21038), .C2(n14232), .A(n14231), .B(n14230), .ZN(
        P1_U3093) );
  INV_X1 U17826 ( .A(n20797), .ZN(n14234) );
  INV_X1 U17827 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n20887) );
  OAI222_X1 U17828 ( .A1(n15610), .A2(n14234), .B1(n15605), .B2(n14233), .C1(
        n15603), .C2(n20887), .ZN(P1_U2897) );
  INV_X1 U17829 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n15336) );
  OAI222_X1 U17830 ( .A1(n14356), .A2(n15543), .B1(n16644), .B2(n15336), .C1(
        n14235), .C2(n16640), .ZN(P1_U2864) );
  NOR2_X1 U17831 ( .A1(n9766), .A2(n14236), .ZN(n14237) );
  XNOR2_X1 U17832 ( .A(n14237), .B(n16999), .ZN(n14238) );
  AOI22_X1 U17833 ( .A1(n14239), .A2(n19915), .B1(n19910), .B2(n14238), .ZN(
        n14247) );
  NAND2_X1 U17834 ( .A1(n14240), .A2(n14284), .ZN(n14243) );
  INV_X1 U17835 ( .A(n14241), .ZN(n14242) );
  AND2_X1 U17836 ( .A1(n14243), .A2(n14242), .ZN(n16996) );
  INV_X1 U17837 ( .A(n16996), .ZN(n17036) );
  AOI22_X1 U17838 ( .A1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n19929), .B1(
        P2_EBX_REG_10__SCAN_IN), .B2(n19917), .ZN(n14244) );
  OAI211_X1 U17839 ( .C1(n17036), .C2(n19880), .A(n14244), .B(n20073), .ZN(
        n14245) );
  AOI21_X1 U17840 ( .B1(n9771), .B2(n19877), .A(n14245), .ZN(n14246) );
  OAI211_X1 U17841 ( .C1(n14248), .C2(n19887), .A(n14247), .B(n14246), .ZN(
        P2_U2845) );
  NOR2_X1 U17842 ( .A1(n19944), .A2(n14249), .ZN(n19935) );
  AND2_X1 U17843 ( .A1(n14251), .A2(n14250), .ZN(n14369) );
  INV_X1 U17844 ( .A(n14369), .ZN(n14252) );
  OAI21_X1 U17845 ( .B1(n19935), .B2(n14253), .A(n14252), .ZN(n14311) );
  AND2_X1 U17846 ( .A1(n16947), .A2(n14254), .ZN(n14255) );
  OR2_X1 U17847 ( .A1(n14255), .A2(n16163), .ZN(n19810) );
  MUX2_X1 U17848 ( .A(n19810), .B(n14256), .S(n19947), .Z(n14257) );
  OAI21_X1 U17849 ( .B1(n14311), .B2(n19959), .A(n14257), .ZN(P2_U2871) );
  XOR2_X1 U17850 ( .A(n14259), .B(n14258), .Z(n17009) );
  INV_X1 U17851 ( .A(n17009), .ZN(n14276) );
  NAND2_X1 U17852 ( .A1(n14261), .A2(n14260), .ZN(n14262) );
  XNOR2_X1 U17853 ( .A(n14263), .B(n14262), .ZN(n17011) );
  NOR2_X1 U17854 ( .A1(n16413), .A2(n17066), .ZN(n20058) );
  AOI21_X1 U17855 ( .B1(n16414), .B2(n14388), .A(n20058), .ZN(n14395) );
  AOI21_X1 U17856 ( .B1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n16414), .A(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n14264) );
  NOR2_X1 U17857 ( .A1(n14395), .A2(n14264), .ZN(n14274) );
  OAI21_X1 U17858 ( .B1(n13703), .B2(n14266), .A(n14265), .ZN(n19987) );
  INV_X1 U17859 ( .A(n14267), .ZN(n14271) );
  INV_X1 U17860 ( .A(n14268), .ZN(n14269) );
  AOI21_X1 U17861 ( .B1(n14271), .B2(n14270), .A(n14269), .ZN(n19909) );
  AOI22_X1 U17862 ( .A1(n19909), .A2(n17074), .B1(n19905), .B2(
        P2_REIP_REG_5__SCAN_IN), .ZN(n14272) );
  OAI21_X1 U17863 ( .B1(n19987), .B2(n17048), .A(n14272), .ZN(n14273) );
  AOI211_X1 U17864 ( .C1(n17011), .C2(n17052), .A(n14274), .B(n14273), .ZN(
        n14275) );
  OAI21_X1 U17865 ( .B1(n14276), .B2(n17071), .A(n14275), .ZN(P2_U3041) );
  AOI21_X1 U17866 ( .B1(n14278), .B2(n13989), .A(n12254), .ZN(n16723) );
  INV_X1 U17867 ( .A(n16723), .ZN(n14296) );
  MUX2_X1 U17868 ( .A(DATAI_10_), .B(BUF1_REG_10__SCAN_IN), .S(n14706), .Z(
        n20907) );
  AOI22_X1 U17869 ( .A1(n15608), .A2(n20907), .B1(P1_EAX_REG_10__SCAN_IN), 
        .B2(n15606), .ZN(n14279) );
  OAI21_X1 U17870 ( .B1(n14296), .B2(n15610), .A(n14279), .ZN(P1_U2894) );
  NAND2_X1 U17871 ( .A1(n9718), .A2(n14280), .ZN(n14281) );
  XNOR2_X1 U17872 ( .A(n17000), .B(n14281), .ZN(n14282) );
  AOI22_X1 U17873 ( .A1(n14283), .A2(n19915), .B1(n19910), .B2(n14282), .ZN(
        n14290) );
  OAI21_X1 U17874 ( .B1(n9784), .B2(n14285), .A(n14284), .ZN(n17002) );
  AOI22_X1 U17875 ( .A1(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n19929), .B1(
        P2_EBX_REG_9__SCAN_IN), .B2(n19917), .ZN(n14286) );
  OAI211_X1 U17876 ( .C1(n17002), .C2(n19880), .A(n14286), .B(n20073), .ZN(
        n14287) );
  AOI21_X1 U17877 ( .B1(n14288), .B2(n19877), .A(n14287), .ZN(n14289) );
  OAI211_X1 U17878 ( .C1(n14291), .C2(n19887), .A(n14290), .B(n14289), .ZN(
        P2_U2846) );
  INV_X1 U17879 ( .A(P1_EBX_REG_10__SCAN_IN), .ZN(n14295) );
  AND2_X1 U17880 ( .A1(n14293), .A2(n14292), .ZN(n14294) );
  OR2_X1 U17881 ( .A1(n14294), .A2(n9836), .ZN(n16635) );
  OAI222_X1 U17882 ( .A1(n14296), .A2(n16640), .B1(n14295), .B2(n16644), .C1(
        n16635), .C2(n15543), .ZN(P1_U2862) );
  NOR2_X1 U17883 ( .A1(n14297), .A2(n13350), .ZN(n14308) );
  NAND2_X1 U17884 ( .A1(n19979), .A2(n14299), .ZN(n16930) );
  OAI22_X1 U17885 ( .A1(n16930), .A2(n14301), .B1(n19979), .B2(n14300), .ZN(
        n14306) );
  NOR2_X1 U17886 ( .A1(n13828), .A2(n14303), .ZN(n14304) );
  NOR2_X1 U17887 ( .A1(n14302), .A2(n14304), .ZN(n16342) );
  INV_X1 U17888 ( .A(n16342), .ZN(n19809) );
  NOR2_X1 U17889 ( .A1(n16023), .A2(n19809), .ZN(n14305) );
  AOI211_X1 U17890 ( .C1(BUF1_REG_16__SCAN_IN), .C2(n16932), .A(n14306), .B(
        n14305), .ZN(n14310) );
  NAND2_X1 U17891 ( .A1(n16933), .A2(BUF2_REG_16__SCAN_IN), .ZN(n14309) );
  OAI211_X1 U17892 ( .C1(n14311), .C2(n19982), .A(n14310), .B(n14309), .ZN(
        P2_U2903) );
  INV_X1 U17893 ( .A(n14315), .ZN(n14347) );
  INV_X1 U17894 ( .A(n14314), .ZN(n21112) );
  AOI21_X1 U17895 ( .B1(n21112), .B2(n14316), .A(n14315), .ZN(n14319) );
  OAI22_X1 U17896 ( .A1(n14319), .A2(n21122), .B1(n14490), .B2(n21113), .ZN(
        n14345) );
  INV_X1 U17897 ( .A(n14490), .ZN(n14322) );
  NAND2_X1 U17898 ( .A1(n14318), .A2(n14317), .ZN(n15815) );
  NAND2_X1 U17899 ( .A1(n14319), .A2(n15815), .ZN(n14320) );
  OR2_X1 U17900 ( .A1(n21122), .A2(n14320), .ZN(n14321) );
  OAI211_X1 U17901 ( .C1(n21085), .C2(n14322), .A(n14321), .B(n21120), .ZN(
        n14344) );
  AOI22_X1 U17902 ( .A1(n14345), .A2(n21134), .B1(
        P1_INSTQUEUE_REG_15__2__SCAN_IN), .B2(n14344), .ZN(n14323) );
  OAI21_X1 U17903 ( .B1(n14501), .B2(n14347), .A(n14323), .ZN(n14324) );
  AOI21_X1 U17904 ( .B1(n20972), .B2(n21136), .A(n14324), .ZN(n14325) );
  OAI21_X1 U17905 ( .B1(n21139), .B2(n14350), .A(n14325), .ZN(P1_U3155) );
  AOI22_X1 U17906 ( .A1(n14345), .A2(n21114), .B1(
        P1_INSTQUEUE_REG_15__0__SCAN_IN), .B2(n14344), .ZN(n14326) );
  OAI21_X1 U17907 ( .B1(n14509), .B2(n14347), .A(n14326), .ZN(n14327) );
  AOI21_X1 U17908 ( .B1(n20972), .B2(n21124), .A(n14327), .ZN(n14328) );
  OAI21_X1 U17909 ( .B1(n21127), .B2(n14350), .A(n14328), .ZN(P1_U3153) );
  AOI22_X1 U17910 ( .A1(n14345), .A2(n21128), .B1(
        P1_INSTQUEUE_REG_15__1__SCAN_IN), .B2(n14344), .ZN(n14329) );
  OAI21_X1 U17911 ( .B1(n14521), .B2(n14347), .A(n14329), .ZN(n14330) );
  AOI21_X1 U17912 ( .B1(n20972), .B2(n21130), .A(n14330), .ZN(n14331) );
  OAI21_X1 U17913 ( .B1(n21133), .B2(n14350), .A(n14331), .ZN(P1_U3154) );
  AOI22_X1 U17914 ( .A1(n14345), .A2(n21152), .B1(
        P1_INSTQUEUE_REG_15__5__SCAN_IN), .B2(n14344), .ZN(n14332) );
  OAI21_X1 U17915 ( .B1(n14505), .B2(n14347), .A(n14332), .ZN(n14333) );
  AOI21_X1 U17916 ( .B1(n20972), .B2(n21154), .A(n14333), .ZN(n14334) );
  OAI21_X1 U17917 ( .B1(n21157), .B2(n14350), .A(n14334), .ZN(P1_U3158) );
  AOI22_X1 U17918 ( .A1(n14345), .A2(n21140), .B1(
        P1_INSTQUEUE_REG_15__3__SCAN_IN), .B2(n14344), .ZN(n14335) );
  OAI21_X1 U17919 ( .B1(n14513), .B2(n14347), .A(n14335), .ZN(n14336) );
  AOI21_X1 U17920 ( .B1(n20972), .B2(n21142), .A(n14336), .ZN(n14337) );
  OAI21_X1 U17921 ( .B1(n21145), .B2(n14350), .A(n14337), .ZN(P1_U3156) );
  AOI22_X1 U17922 ( .A1(n14345), .A2(n21165), .B1(
        P1_INSTQUEUE_REG_15__7__SCAN_IN), .B2(n14344), .ZN(n14338) );
  OAI21_X1 U17923 ( .B1(n14528), .B2(n14347), .A(n14338), .ZN(n14339) );
  AOI21_X1 U17924 ( .B1(n20972), .B2(n21168), .A(n14339), .ZN(n14340) );
  OAI21_X1 U17925 ( .B1(n21174), .B2(n14350), .A(n14340), .ZN(P1_U3160) );
  AOI22_X1 U17926 ( .A1(n14345), .A2(n21158), .B1(
        P1_INSTQUEUE_REG_15__6__SCAN_IN), .B2(n14344), .ZN(n14341) );
  OAI21_X1 U17927 ( .B1(n14497), .B2(n14347), .A(n14341), .ZN(n14342) );
  AOI21_X1 U17928 ( .B1(n20972), .B2(n21160), .A(n14342), .ZN(n14343) );
  OAI21_X1 U17929 ( .B1(n21163), .B2(n14350), .A(n14343), .ZN(P1_U3159) );
  AOI22_X1 U17930 ( .A1(n14345), .A2(n21146), .B1(
        P1_INSTQUEUE_REG_15__4__SCAN_IN), .B2(n14344), .ZN(n14346) );
  OAI21_X1 U17931 ( .B1(n14517), .B2(n14347), .A(n14346), .ZN(n14348) );
  AOI21_X1 U17932 ( .B1(n20972), .B2(n21148), .A(n14348), .ZN(n14349) );
  OAI21_X1 U17933 ( .B1(n21151), .B2(n14350), .A(n14349), .ZN(P1_U3157) );
  NAND2_X1 U17934 ( .A1(n9818), .A2(n14352), .ZN(n14353) );
  XNOR2_X1 U17935 ( .A(n14351), .B(n14353), .ZN(n14366) );
  AOI21_X1 U17936 ( .B1(n15783), .B2(n14355), .A(n14354), .ZN(n16827) );
  OAI21_X1 U17937 ( .B1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n15738), .A(
        n16827), .ZN(n16817) );
  OAI22_X1 U17938 ( .A1(n14356), .A2(n20925), .B1(n21210), .B2(n16823), .ZN(
        n14359) );
  NOR2_X1 U17939 ( .A1(n15770), .A2(n15799), .ZN(n16822) );
  NAND2_X1 U17940 ( .A1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n16822), .ZN(
        n16821) );
  AOI221_X1 U17941 ( .B1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .C1(n14357), .C2(n11419), .A(
        n16821), .ZN(n14358) );
  AOI211_X1 U17942 ( .C1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .C2(n16817), .A(
        n14359), .B(n14358), .ZN(n14360) );
  OAI21_X1 U17943 ( .B1(n14366), .B2(n16792), .A(n14360), .ZN(P1_U3023) );
  AOI22_X1 U17944 ( .A1(n16734), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(
        n16782), .B2(P1_REIP_REG_8__SCAN_IN), .ZN(n14361) );
  OAI21_X1 U17945 ( .B1(n16743), .B2(n14362), .A(n14361), .ZN(n14363) );
  AOI21_X1 U17946 ( .B1(n14364), .B2(n16739), .A(n14363), .ZN(n14365) );
  OAI21_X1 U17947 ( .B1(n14366), .B2(n20773), .A(n14365), .ZN(P1_U2991) );
  OAI21_X1 U17948 ( .B1(n14369), .B2(n14368), .A(n14367), .ZN(n16925) );
  OAI22_X1 U17949 ( .A1(n16930), .A2(n20088), .B1(n19979), .B2(n14370), .ZN(
        n14378) );
  INV_X1 U17950 ( .A(n14371), .ZN(n14376) );
  INV_X1 U17951 ( .A(n14302), .ZN(n14374) );
  INV_X1 U17952 ( .A(n14372), .ZN(n14373) );
  NAND2_X1 U17953 ( .A1(n14374), .A2(n14373), .ZN(n14375) );
  NAND2_X1 U17954 ( .A1(n14376), .A2(n14375), .ZN(n19802) );
  NOR2_X1 U17955 ( .A1(n16023), .A2(n19802), .ZN(n14377) );
  AOI211_X1 U17956 ( .C1(BUF1_REG_17__SCAN_IN), .C2(n16932), .A(n14378), .B(
        n14377), .ZN(n14380) );
  NAND2_X1 U17957 ( .A1(n16933), .A2(BUF2_REG_17__SCAN_IN), .ZN(n14379) );
  OAI211_X1 U17958 ( .C1(n16925), .C2(n19982), .A(n14380), .B(n14379), .ZN(
        P2_U2902) );
  XNOR2_X1 U17959 ( .A(n14381), .B(n14382), .ZN(n14489) );
  NAND2_X1 U17960 ( .A1(n14384), .A2(n14383), .ZN(n14386) );
  NAND2_X1 U17961 ( .A1(n14386), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n14385) );
  OAI21_X1 U17962 ( .B1(n14386), .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n14385), .ZN(n14387) );
  INV_X1 U17963 ( .A(n14387), .ZN(n14487) );
  INV_X1 U17964 ( .A(n16414), .ZN(n20061) );
  OR3_X1 U17965 ( .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n14388), .A3(
        n20061), .ZN(n14393) );
  INV_X1 U17966 ( .A(n19901), .ZN(n14391) );
  OAI22_X1 U17967 ( .A1(n20062), .A2(n19895), .B1(n12009), .B2(n14389), .ZN(
        n14390) );
  AOI21_X1 U17968 ( .B1(n14391), .B2(n20057), .A(n14390), .ZN(n14392) );
  OAI211_X1 U17969 ( .C1(n14395), .C2(n14394), .A(n14393), .B(n14392), .ZN(
        n14396) );
  AOI21_X1 U17970 ( .B1(n14487), .B2(n17052), .A(n14396), .ZN(n14397) );
  OAI21_X1 U17971 ( .B1(n17071), .B2(n14489), .A(n14397), .ZN(P2_U3040) );
  NAND2_X1 U17972 ( .A1(n14431), .A2(n21085), .ZN(n14399) );
  NOR2_X2 U17973 ( .A1(n21008), .A2(n14587), .ZN(n21076) );
  NAND2_X1 U17974 ( .A1(n21085), .A2(n21118), .ZN(n20942) );
  OAI21_X1 U17975 ( .B1(n14399), .B2(n21076), .A(n20942), .ZN(n14405) );
  AND2_X1 U17976 ( .A1(n21055), .A2(n20945), .ZN(n14402) );
  NAND2_X1 U17977 ( .A1(n14491), .A2(n21010), .ZN(n14403) );
  INV_X1 U17978 ( .A(n14403), .ZN(n14535) );
  AOI22_X1 U17979 ( .A1(n14405), .A2(n14402), .B1(n14400), .B2(n14535), .ZN(
        n14434) );
  NOR2_X1 U17980 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n14401), .ZN(
        n14429) );
  INV_X1 U17981 ( .A(n14402), .ZN(n14404) );
  AND2_X1 U17982 ( .A1(n14403), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n14538) );
  AOI21_X1 U17983 ( .B1(n14405), .B2(n14404), .A(n14538), .ZN(n14406) );
  OAI211_X1 U17984 ( .C1(n14429), .C2(n20953), .A(n21016), .B(n14406), .ZN(
        n14428) );
  AOI22_X1 U17985 ( .A1(n21167), .A2(n14429), .B1(
        P1_INSTQUEUE_REG_6__7__SCAN_IN), .B2(n14428), .ZN(n14407) );
  OAI21_X1 U17986 ( .B1(n21054), .B2(n14431), .A(n14407), .ZN(n14408) );
  AOI21_X1 U17987 ( .B1(n21076), .B2(n21049), .A(n14408), .ZN(n14409) );
  OAI21_X1 U17988 ( .B1(n14434), .B2(n14607), .A(n14409), .ZN(P1_U3088) );
  AOI22_X1 U17989 ( .A1(n21153), .A2(n14429), .B1(
        P1_INSTQUEUE_REG_6__5__SCAN_IN), .B2(n14428), .ZN(n14410) );
  OAI21_X1 U17990 ( .B1(n21042), .B2(n14431), .A(n14410), .ZN(n14411) );
  AOI21_X1 U17991 ( .B1(n21076), .B2(n21039), .A(n14411), .ZN(n14412) );
  OAI21_X1 U17992 ( .B1(n14434), .B2(n14622), .A(n14412), .ZN(P1_U3086) );
  AOI22_X1 U17993 ( .A1(n21115), .A2(n14429), .B1(
        P1_INSTQUEUE_REG_6__0__SCAN_IN), .B2(n14428), .ZN(n14413) );
  OAI21_X1 U17994 ( .B1(n21022), .B2(n14431), .A(n14413), .ZN(n14414) );
  AOI21_X1 U17995 ( .B1(n21076), .B2(n21019), .A(n14414), .ZN(n14415) );
  OAI21_X1 U17996 ( .B1(n14434), .B2(n14617), .A(n14415), .ZN(P1_U3081) );
  AOI22_X1 U17997 ( .A1(n21141), .A2(n14429), .B1(
        P1_INSTQUEUE_REG_6__3__SCAN_IN), .B2(n14428), .ZN(n14416) );
  OAI21_X1 U17998 ( .B1(n21034), .B2(n14431), .A(n14416), .ZN(n14417) );
  AOI21_X1 U17999 ( .B1(n21076), .B2(n21031), .A(n14417), .ZN(n14418) );
  OAI21_X1 U18000 ( .B1(n14434), .B2(n14602), .A(n14418), .ZN(P1_U3084) );
  AOI22_X1 U18001 ( .A1(n21135), .A2(n14429), .B1(
        P1_INSTQUEUE_REG_6__2__SCAN_IN), .B2(n14428), .ZN(n14419) );
  OAI21_X1 U18002 ( .B1(n21030), .B2(n14431), .A(n14419), .ZN(n14420) );
  AOI21_X1 U18003 ( .B1(n21076), .B2(n21027), .A(n14420), .ZN(n14421) );
  OAI21_X1 U18004 ( .B1(n14434), .B2(n14632), .A(n14421), .ZN(P1_U3083) );
  AOI22_X1 U18005 ( .A1(n21129), .A2(n14429), .B1(
        P1_INSTQUEUE_REG_6__1__SCAN_IN), .B2(n14428), .ZN(n14422) );
  OAI21_X1 U18006 ( .B1(n21026), .B2(n14431), .A(n14422), .ZN(n14423) );
  AOI21_X1 U18007 ( .B1(n21076), .B2(n21023), .A(n14423), .ZN(n14424) );
  OAI21_X1 U18008 ( .B1(n14434), .B2(n14612), .A(n14424), .ZN(P1_U3082) );
  AOI22_X1 U18009 ( .A1(n21147), .A2(n14429), .B1(
        P1_INSTQUEUE_REG_6__4__SCAN_IN), .B2(n14428), .ZN(n14425) );
  OAI21_X1 U18010 ( .B1(n21038), .B2(n14431), .A(n14425), .ZN(n14426) );
  AOI21_X1 U18011 ( .B1(n21076), .B2(n21035), .A(n14426), .ZN(n14427) );
  OAI21_X1 U18012 ( .B1(n14434), .B2(n14627), .A(n14427), .ZN(P1_U3085) );
  AOI22_X1 U18013 ( .A1(n21159), .A2(n14429), .B1(
        P1_INSTQUEUE_REG_6__6__SCAN_IN), .B2(n14428), .ZN(n14430) );
  OAI21_X1 U18014 ( .B1(n21046), .B2(n14431), .A(n14430), .ZN(n14432) );
  AOI21_X1 U18015 ( .B1(n21076), .B2(n21043), .A(n14432), .ZN(n14433) );
  OAI21_X1 U18016 ( .B1(n14434), .B2(n14640), .A(n14433), .ZN(P1_U3087) );
  NAND2_X1 U18017 ( .A1(n16139), .A2(n14436), .ZN(n14437) );
  NAND2_X1 U18018 ( .A1(n16108), .A2(n14437), .ZN(n19762) );
  NAND2_X1 U18019 ( .A1(n10631), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n14441) );
  NAND2_X1 U18020 ( .A1(n14951), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n14440) );
  AOI22_X1 U18021 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n10500), .B1(
        n14885), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n14439) );
  NAND2_X1 U18022 ( .A1(n10507), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n14438) );
  NAND4_X1 U18023 ( .A1(n14441), .A2(n14440), .A3(n14439), .A4(n14438), .ZN(
        n14447) );
  AOI22_X1 U18024 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n10498), .B1(
        n10499), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n14445) );
  NAND2_X1 U18025 ( .A1(n14908), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n14444) );
  NAND2_X1 U18026 ( .A1(n14909), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n14443) );
  NAND2_X1 U18027 ( .A1(n14910), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n14442) );
  NAND4_X1 U18028 ( .A1(n14445), .A2(n14444), .A3(n14443), .A4(n14442), .ZN(
        n14446) );
  NOR2_X1 U18029 ( .A1(n14447), .A2(n14446), .ZN(n14457) );
  INV_X1 U18030 ( .A(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n14448) );
  OAI22_X1 U18031 ( .A1(n14919), .A2(n14449), .B1(n14917), .B2(n14448), .ZN(
        n14455) );
  AOI22_X1 U18032 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n14967), .B1(
        n11881), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n14452) );
  NAND2_X1 U18033 ( .A1(n14450), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n14451) );
  OAI211_X1 U18034 ( .C1(n14473), .C2(n14453), .A(n14452), .B(n14451), .ZN(
        n14454) );
  NOR2_X1 U18035 ( .A1(n14455), .A2(n14454), .ZN(n14456) );
  AND2_X1 U18036 ( .A1(n14457), .A2(n14456), .ZN(n14482) );
  NAND2_X1 U18037 ( .A1(n10631), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(
        n14461) );
  NAND2_X1 U18038 ( .A1(n14951), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n14460) );
  AOI22_X1 U18039 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n10500), .B1(
        n14885), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n14459) );
  NAND2_X1 U18040 ( .A1(n10507), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n14458) );
  NAND4_X1 U18041 ( .A1(n14461), .A2(n14460), .A3(n14459), .A4(n14458), .ZN(
        n14467) );
  AOI22_X1 U18042 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n10498), .B1(
        n10499), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n14465) );
  NAND2_X1 U18043 ( .A1(n14908), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n14464) );
  NAND2_X1 U18044 ( .A1(n14909), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n14463) );
  NAND2_X1 U18045 ( .A1(n14910), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n14462) );
  NAND4_X1 U18046 ( .A1(n14465), .A2(n14464), .A3(n14463), .A4(n14462), .ZN(
        n14466) );
  NOR2_X1 U18047 ( .A1(n14467), .A2(n14466), .ZN(n14477) );
  OAI22_X1 U18048 ( .A1(n14919), .A2(n14469), .B1(n14917), .B2(n14468), .ZN(
        n14475) );
  AOI22_X1 U18049 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n14967), .B1(
        n11881), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n14471) );
  NAND2_X1 U18050 ( .A1(n14450), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n14470) );
  OAI211_X1 U18051 ( .C1(n14473), .C2(n14472), .A(n14471), .B(n14470), .ZN(
        n14474) );
  NOR2_X1 U18052 ( .A1(n14475), .A2(n14474), .ZN(n14476) );
  AND2_X1 U18053 ( .A1(n14477), .A2(n14476), .ZN(n16016) );
  INV_X1 U18054 ( .A(n16016), .ZN(n14478) );
  AND2_X1 U18055 ( .A1(n14479), .A2(n14478), .ZN(n14480) );
  AOI21_X1 U18056 ( .B1(n14482), .B2(n14481), .A(n14903), .ZN(n16006) );
  NAND2_X1 U18057 ( .A1(n16006), .A2(n16926), .ZN(n14484) );
  NAND2_X1 U18058 ( .A1(n19947), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n14483) );
  OAI211_X1 U18059 ( .C1(n19762), .C2(n19947), .A(n14484), .B(n14483), .ZN(
        P2_U2867) );
  OAI22_X1 U18060 ( .A1(n14389), .A2(n20073), .B1(n20045), .B2(n19893), .ZN(
        n14486) );
  OAI22_X1 U18061 ( .A1(n16202), .A2(n19895), .B1(n20055), .B2(n10091), .ZN(
        n14485) );
  AOI211_X1 U18062 ( .C1(n14487), .C2(n17010), .A(n14486), .B(n14485), .ZN(
        n14488) );
  OAI21_X1 U18063 ( .B1(n16974), .B2(n14489), .A(n14488), .ZN(P2_U3008) );
  NOR2_X1 U18064 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n14490), .ZN(
        n14495) );
  INV_X1 U18065 ( .A(n14495), .ZN(n14527) );
  NAND2_X1 U18066 ( .A1(n21112), .A2(n20945), .ZN(n14493) );
  NAND2_X1 U18067 ( .A1(n14491), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n14598) );
  OAI22_X1 U18068 ( .A1(n14493), .A2(n21122), .B1(n21012), .B2(n14598), .ZN(
        n14525) );
  OAI21_X1 U18069 ( .B1(n21169), .B2(n14530), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n14492) );
  AOI21_X1 U18070 ( .B1(n14493), .B2(n14492), .A(P1_STATE2_REG_3__SCAN_IN), 
        .ZN(n14494) );
  NAND2_X1 U18071 ( .A1(n14598), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n14592) );
  OAI211_X1 U18072 ( .C1(n14495), .C2(n14494), .A(n21016), .B(n14592), .ZN(
        n14524) );
  AOI22_X1 U18073 ( .A1(n14525), .A2(n21158), .B1(
        P1_INSTQUEUE_REG_14__6__SCAN_IN), .B2(n14524), .ZN(n14496) );
  OAI21_X1 U18074 ( .B1(n14497), .B2(n14527), .A(n14496), .ZN(n14498) );
  AOI21_X1 U18075 ( .B1(n14530), .B2(n21160), .A(n14498), .ZN(n14499) );
  OAI21_X1 U18076 ( .B1(n21163), .B2(n14532), .A(n14499), .ZN(P1_U3151) );
  AOI22_X1 U18077 ( .A1(n14525), .A2(n21134), .B1(
        P1_INSTQUEUE_REG_14__2__SCAN_IN), .B2(n14524), .ZN(n14500) );
  OAI21_X1 U18078 ( .B1(n14501), .B2(n14527), .A(n14500), .ZN(n14502) );
  AOI21_X1 U18079 ( .B1(n14530), .B2(n21136), .A(n14502), .ZN(n14503) );
  OAI21_X1 U18080 ( .B1(n21139), .B2(n14532), .A(n14503), .ZN(P1_U3147) );
  AOI22_X1 U18081 ( .A1(n14525), .A2(n21152), .B1(
        P1_INSTQUEUE_REG_14__5__SCAN_IN), .B2(n14524), .ZN(n14504) );
  OAI21_X1 U18082 ( .B1(n14505), .B2(n14527), .A(n14504), .ZN(n14506) );
  AOI21_X1 U18083 ( .B1(n14530), .B2(n21154), .A(n14506), .ZN(n14507) );
  OAI21_X1 U18084 ( .B1(n21157), .B2(n14532), .A(n14507), .ZN(P1_U3150) );
  AOI22_X1 U18085 ( .A1(n14525), .A2(n21114), .B1(
        P1_INSTQUEUE_REG_14__0__SCAN_IN), .B2(n14524), .ZN(n14508) );
  OAI21_X1 U18086 ( .B1(n14509), .B2(n14527), .A(n14508), .ZN(n14510) );
  AOI21_X1 U18087 ( .B1(n14530), .B2(n21124), .A(n14510), .ZN(n14511) );
  OAI21_X1 U18088 ( .B1(n21127), .B2(n14532), .A(n14511), .ZN(P1_U3145) );
  AOI22_X1 U18089 ( .A1(n14525), .A2(n21140), .B1(
        P1_INSTQUEUE_REG_14__3__SCAN_IN), .B2(n14524), .ZN(n14512) );
  OAI21_X1 U18090 ( .B1(n14513), .B2(n14527), .A(n14512), .ZN(n14514) );
  AOI21_X1 U18091 ( .B1(n14530), .B2(n21142), .A(n14514), .ZN(n14515) );
  OAI21_X1 U18092 ( .B1(n21145), .B2(n14532), .A(n14515), .ZN(P1_U3148) );
  AOI22_X1 U18093 ( .A1(n14525), .A2(n21146), .B1(
        P1_INSTQUEUE_REG_14__4__SCAN_IN), .B2(n14524), .ZN(n14516) );
  OAI21_X1 U18094 ( .B1(n14517), .B2(n14527), .A(n14516), .ZN(n14518) );
  AOI21_X1 U18095 ( .B1(n14530), .B2(n21148), .A(n14518), .ZN(n14519) );
  OAI21_X1 U18096 ( .B1(n21151), .B2(n14532), .A(n14519), .ZN(P1_U3149) );
  AOI22_X1 U18097 ( .A1(n14525), .A2(n21128), .B1(
        P1_INSTQUEUE_REG_14__1__SCAN_IN), .B2(n14524), .ZN(n14520) );
  OAI21_X1 U18098 ( .B1(n14521), .B2(n14527), .A(n14520), .ZN(n14522) );
  AOI21_X1 U18099 ( .B1(n14530), .B2(n21130), .A(n14522), .ZN(n14523) );
  OAI21_X1 U18100 ( .B1(n21133), .B2(n14532), .A(n14523), .ZN(P1_U3146) );
  AOI22_X1 U18101 ( .A1(n14525), .A2(n21165), .B1(
        P1_INSTQUEUE_REG_14__7__SCAN_IN), .B2(n14524), .ZN(n14526) );
  OAI21_X1 U18102 ( .B1(n14528), .B2(n14527), .A(n14526), .ZN(n14529) );
  AOI21_X1 U18103 ( .B1(n14530), .B2(n21168), .A(n14529), .ZN(n14531) );
  OAI21_X1 U18104 ( .B1(n21174), .B2(n14532), .A(n14531), .ZN(P1_U3152) );
  NAND2_X1 U18105 ( .A1(n14571), .A2(n21085), .ZN(n14534) );
  NOR2_X2 U18106 ( .A1(n20982), .A2(n14587), .ZN(n21001) );
  OAI21_X1 U18107 ( .B1(n14534), .B2(n21001), .A(n20942), .ZN(n14540) );
  NOR2_X1 U18108 ( .A1(n20946), .A2(n14001), .ZN(n14537) );
  AOI22_X1 U18109 ( .A1(n14540), .A2(n14537), .B1(n20954), .B2(n14535), .ZN(
        n14574) );
  NOR2_X1 U18110 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n14536), .ZN(
        n14569) );
  INV_X1 U18111 ( .A(n14537), .ZN(n14539) );
  AOI211_X1 U18112 ( .C1(n14540), .C2(n14539), .A(n14538), .B(n14594), .ZN(
        n14541) );
  AOI22_X1 U18113 ( .A1(n21167), .A2(n14569), .B1(
        P1_INSTQUEUE_REG_2__7__SCAN_IN), .B2(n14568), .ZN(n14542) );
  OAI21_X1 U18114 ( .B1(n14571), .B2(n21054), .A(n14542), .ZN(n14543) );
  AOI21_X1 U18115 ( .B1(n21001), .B2(n21049), .A(n14543), .ZN(n14544) );
  OAI21_X1 U18116 ( .B1(n14574), .B2(n14607), .A(n14544), .ZN(P1_U3056) );
  AOI22_X1 U18117 ( .A1(n21115), .A2(n14569), .B1(
        P1_INSTQUEUE_REG_2__0__SCAN_IN), .B2(n14568), .ZN(n14545) );
  OAI21_X1 U18118 ( .B1(n14571), .B2(n21022), .A(n14545), .ZN(n14546) );
  AOI21_X1 U18119 ( .B1(n21001), .B2(n21019), .A(n14546), .ZN(n14547) );
  OAI21_X1 U18120 ( .B1(n14574), .B2(n14617), .A(n14547), .ZN(P1_U3049) );
  AOI22_X1 U18121 ( .A1(n21135), .A2(n14569), .B1(
        P1_INSTQUEUE_REG_2__2__SCAN_IN), .B2(n14568), .ZN(n14548) );
  OAI21_X1 U18122 ( .B1(n14571), .B2(n21030), .A(n14548), .ZN(n14549) );
  AOI21_X1 U18123 ( .B1(n21001), .B2(n21027), .A(n14549), .ZN(n14550) );
  OAI21_X1 U18124 ( .B1(n14574), .B2(n14632), .A(n14550), .ZN(P1_U3051) );
  AOI22_X1 U18125 ( .A1(n21141), .A2(n14569), .B1(
        P1_INSTQUEUE_REG_2__3__SCAN_IN), .B2(n14568), .ZN(n14551) );
  OAI21_X1 U18126 ( .B1(n14571), .B2(n21034), .A(n14551), .ZN(n14552) );
  AOI21_X1 U18127 ( .B1(n21001), .B2(n21031), .A(n14552), .ZN(n14553) );
  OAI21_X1 U18128 ( .B1(n14574), .B2(n14602), .A(n14553), .ZN(P1_U3052) );
  AOI22_X1 U18129 ( .A1(n21129), .A2(n14569), .B1(
        P1_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n14568), .ZN(n14554) );
  OAI21_X1 U18130 ( .B1(n14571), .B2(n21026), .A(n14554), .ZN(n14555) );
  AOI21_X1 U18131 ( .B1(n21001), .B2(n21023), .A(n14555), .ZN(n14556) );
  OAI21_X1 U18132 ( .B1(n14574), .B2(n14612), .A(n14556), .ZN(P1_U3050) );
  AOI22_X1 U18133 ( .A1(n21153), .A2(n14569), .B1(
        P1_INSTQUEUE_REG_2__5__SCAN_IN), .B2(n14568), .ZN(n14557) );
  OAI21_X1 U18134 ( .B1(n14571), .B2(n21042), .A(n14557), .ZN(n14558) );
  AOI21_X1 U18135 ( .B1(n21001), .B2(n21039), .A(n14558), .ZN(n14559) );
  OAI21_X1 U18136 ( .B1(n14574), .B2(n14622), .A(n14559), .ZN(P1_U3054) );
  NAND2_X1 U18137 ( .A1(n14560), .A2(n14561), .ZN(n14562) );
  NAND2_X1 U18138 ( .A1(n14563), .A2(n14562), .ZN(n15686) );
  INV_X1 U18139 ( .A(n15554), .ZN(n14564) );
  OAI222_X1 U18140 ( .A1(n15686), .A2(n15610), .B1(n15605), .B2(n14564), .C1(
        n20879), .C2(n15603), .ZN(P1_U2893) );
  AOI22_X1 U18141 ( .A1(n21159), .A2(n14569), .B1(
        P1_INSTQUEUE_REG_2__6__SCAN_IN), .B2(n14568), .ZN(n14565) );
  OAI21_X1 U18142 ( .B1(n14571), .B2(n21046), .A(n14565), .ZN(n14566) );
  AOI21_X1 U18143 ( .B1(n21001), .B2(n21043), .A(n14566), .ZN(n14567) );
  OAI21_X1 U18144 ( .B1(n14574), .B2(n14640), .A(n14567), .ZN(P1_U3055) );
  AOI22_X1 U18145 ( .A1(n21147), .A2(n14569), .B1(
        P1_INSTQUEUE_REG_2__4__SCAN_IN), .B2(n14568), .ZN(n14570) );
  OAI21_X1 U18146 ( .B1(n14571), .B2(n21038), .A(n14570), .ZN(n14572) );
  AOI21_X1 U18147 ( .B1(n21001), .B2(n21035), .A(n14572), .ZN(n14573) );
  OAI21_X1 U18148 ( .B1(n14574), .B2(n14627), .A(n14573), .ZN(P1_U3053) );
  NOR2_X1 U18149 ( .A1(n9836), .A2(n14575), .ZN(n14576) );
  OR2_X1 U18150 ( .A1(n14675), .A2(n14576), .ZN(n16798) );
  INV_X1 U18151 ( .A(P1_EBX_REG_11__SCAN_IN), .ZN(n14655) );
  OAI222_X1 U18152 ( .A1(n16798), .A2(n15543), .B1(n14655), .B2(n16644), .C1(
        n15686), .C2(n16640), .ZN(P1_U2861) );
  INV_X1 U18153 ( .A(n16933), .ZN(n16015) );
  INV_X1 U18154 ( .A(BUF2_REG_18__SCAN_IN), .ZN(n14586) );
  NAND2_X1 U18155 ( .A1(n14577), .A2(n16936), .ZN(n14585) );
  OAI22_X1 U18156 ( .A1(n16930), .A2(n20092), .B1(n16020), .B2(n14578), .ZN(
        n14583) );
  NOR2_X1 U18157 ( .A1(n14371), .A2(n14580), .ZN(n14581) );
  NOR2_X1 U18158 ( .A1(n14579), .A2(n14581), .ZN(n16318) );
  INV_X1 U18159 ( .A(n16318), .ZN(n19786) );
  NOR2_X1 U18160 ( .A1(n16023), .A2(n19786), .ZN(n14582) );
  AOI211_X1 U18161 ( .C1(BUF1_REG_18__SCAN_IN), .C2(n16932), .A(n14583), .B(
        n14582), .ZN(n14584) );
  OAI211_X1 U18162 ( .C1(n16015), .C2(n14586), .A(n14585), .B(n14584), .ZN(
        P2_U2901) );
  INV_X1 U18163 ( .A(n14587), .ZN(n14588) );
  NOR2_X1 U18164 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n14590), .ZN(
        n14637) );
  NAND2_X1 U18165 ( .A1(n14639), .A2(n21085), .ZN(n14591) );
  OAI21_X1 U18166 ( .B1(n14591), .B2(n21105), .A(n20942), .ZN(n14601) );
  NOR2_X1 U18167 ( .A1(n21081), .A2(n14001), .ZN(n14600) );
  INV_X1 U18168 ( .A(n14600), .ZN(n14595) );
  INV_X1 U18169 ( .A(n14592), .ZN(n14593) );
  AOI211_X1 U18170 ( .C1(n14601), .C2(n14595), .A(n14594), .B(n14593), .ZN(
        n14596) );
  OAI21_X1 U18171 ( .B1(n14637), .B2(n20953), .A(n14596), .ZN(n14636) );
  AOI22_X1 U18172 ( .A1(n21141), .A2(n14637), .B1(
        P1_INSTQUEUE_REG_10__3__SCAN_IN), .B2(n14636), .ZN(n14597) );
  OAI21_X1 U18173 ( .B1(n14639), .B2(n21034), .A(n14597), .ZN(n14604) );
  INV_X1 U18174 ( .A(n14598), .ZN(n14599) );
  AOI22_X1 U18175 ( .A1(n14601), .A2(n14600), .B1(n20954), .B2(n14599), .ZN(
        n14641) );
  NOR2_X1 U18176 ( .A1(n14641), .A2(n14602), .ZN(n14603) );
  AOI211_X1 U18177 ( .C1(n21105), .C2(n21031), .A(n14604), .B(n14603), .ZN(
        n14605) );
  INV_X1 U18178 ( .A(n14605), .ZN(P1_U3116) );
  AOI22_X1 U18179 ( .A1(n21167), .A2(n14637), .B1(
        P1_INSTQUEUE_REG_10__7__SCAN_IN), .B2(n14636), .ZN(n14606) );
  OAI21_X1 U18180 ( .B1(n14639), .B2(n21054), .A(n14606), .ZN(n14609) );
  NOR2_X1 U18181 ( .A1(n14641), .A2(n14607), .ZN(n14608) );
  AOI211_X1 U18182 ( .C1(n21105), .C2(n21049), .A(n14609), .B(n14608), .ZN(
        n14610) );
  INV_X1 U18183 ( .A(n14610), .ZN(P1_U3120) );
  AOI22_X1 U18184 ( .A1(n21129), .A2(n14637), .B1(
        P1_INSTQUEUE_REG_10__1__SCAN_IN), .B2(n14636), .ZN(n14611) );
  OAI21_X1 U18185 ( .B1(n14639), .B2(n21026), .A(n14611), .ZN(n14614) );
  NOR2_X1 U18186 ( .A1(n14641), .A2(n14612), .ZN(n14613) );
  AOI211_X1 U18187 ( .C1(n21105), .C2(n21023), .A(n14614), .B(n14613), .ZN(
        n14615) );
  INV_X1 U18188 ( .A(n14615), .ZN(P1_U3114) );
  AOI22_X1 U18189 ( .A1(n21115), .A2(n14637), .B1(
        P1_INSTQUEUE_REG_10__0__SCAN_IN), .B2(n14636), .ZN(n14616) );
  OAI21_X1 U18190 ( .B1(n14639), .B2(n21022), .A(n14616), .ZN(n14619) );
  NOR2_X1 U18191 ( .A1(n14641), .A2(n14617), .ZN(n14618) );
  AOI211_X1 U18192 ( .C1(n21105), .C2(n21019), .A(n14619), .B(n14618), .ZN(
        n14620) );
  INV_X1 U18193 ( .A(n14620), .ZN(P1_U3113) );
  AOI22_X1 U18194 ( .A1(n21153), .A2(n14637), .B1(
        P1_INSTQUEUE_REG_10__5__SCAN_IN), .B2(n14636), .ZN(n14621) );
  OAI21_X1 U18195 ( .B1(n14639), .B2(n21042), .A(n14621), .ZN(n14624) );
  NOR2_X1 U18196 ( .A1(n14641), .A2(n14622), .ZN(n14623) );
  AOI211_X1 U18197 ( .C1(n21105), .C2(n21039), .A(n14624), .B(n14623), .ZN(
        n14625) );
  INV_X1 U18198 ( .A(n14625), .ZN(P1_U3118) );
  AOI22_X1 U18199 ( .A1(n21147), .A2(n14637), .B1(
        P1_INSTQUEUE_REG_10__4__SCAN_IN), .B2(n14636), .ZN(n14626) );
  OAI21_X1 U18200 ( .B1(n14639), .B2(n21038), .A(n14626), .ZN(n14629) );
  NOR2_X1 U18201 ( .A1(n14641), .A2(n14627), .ZN(n14628) );
  AOI211_X1 U18202 ( .C1(n21105), .C2(n21035), .A(n14629), .B(n14628), .ZN(
        n14630) );
  INV_X1 U18203 ( .A(n14630), .ZN(P1_U3117) );
  AOI22_X1 U18204 ( .A1(n21135), .A2(n14637), .B1(
        P1_INSTQUEUE_REG_10__2__SCAN_IN), .B2(n14636), .ZN(n14631) );
  OAI21_X1 U18205 ( .B1(n14639), .B2(n21030), .A(n14631), .ZN(n14634) );
  NOR2_X1 U18206 ( .A1(n14641), .A2(n14632), .ZN(n14633) );
  AOI211_X1 U18207 ( .C1(n21105), .C2(n21027), .A(n14634), .B(n14633), .ZN(
        n14635) );
  INV_X1 U18208 ( .A(n14635), .ZN(P1_U3115) );
  AOI22_X1 U18209 ( .A1(n21159), .A2(n14637), .B1(
        P1_INSTQUEUE_REG_10__6__SCAN_IN), .B2(n14636), .ZN(n14638) );
  OAI21_X1 U18210 ( .B1(n14639), .B2(n21046), .A(n14638), .ZN(n14643) );
  NOR2_X1 U18211 ( .A1(n14641), .A2(n14640), .ZN(n14642) );
  AOI211_X1 U18212 ( .C1(n21105), .C2(n21043), .A(n14643), .B(n14642), .ZN(
        n14644) );
  INV_X1 U18213 ( .A(n14644), .ZN(P1_U3119) );
  XNOR2_X1 U18214 ( .A(n16673), .B(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n14646) );
  XNOR2_X1 U18215 ( .A(n14645), .B(n14646), .ZN(n16812) );
  NAND2_X1 U18216 ( .A1(n16812), .A2(n16740), .ZN(n14650) );
  NOR2_X1 U18217 ( .A1(n16823), .A2(n21213), .ZN(n16808) );
  NOR2_X1 U18218 ( .A1(n16743), .A2(n14647), .ZN(n14648) );
  AOI211_X1 U18219 ( .C1(n16734), .C2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .A(
        n16808), .B(n14648), .ZN(n14649) );
  OAI211_X1 U18220 ( .C1(n16700), .C2(n14651), .A(n14650), .B(n14649), .ZN(
        P1_U2990) );
  INV_X1 U18221 ( .A(n15686), .ZN(n14652) );
  NAND2_X1 U18222 ( .A1(n14652), .A2(n20808), .ZN(n14662) );
  INV_X1 U18223 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n21215) );
  NOR2_X1 U18224 ( .A1(n21215), .A2(n21213), .ZN(n14653) );
  INV_X1 U18225 ( .A(n15461), .ZN(n15149) );
  AOI21_X1 U18226 ( .B1(n14670), .B2(n14653), .A(n15149), .ZN(n16637) );
  INV_X1 U18227 ( .A(n14654), .ZN(n16632) );
  NOR4_X1 U18228 ( .A1(P1_REIP_REG_11__SCAN_IN), .A2(n21213), .A3(n21215), 
        .A4(n16632), .ZN(n14660) );
  OAI22_X1 U18229 ( .A1(n16798), .A2(n20860), .B1(n16622), .B2(n14655), .ZN(
        n14656) );
  INV_X1 U18230 ( .A(n14656), .ZN(n14657) );
  OAI211_X1 U18231 ( .C1(n20818), .C2(n14658), .A(n14657), .B(n20816), .ZN(
        n14659) );
  AOI211_X1 U18232 ( .C1(P1_REIP_REG_11__SCAN_IN), .C2(n16637), .A(n14660), 
        .B(n14659), .ZN(n14661) );
  OAI211_X1 U18233 ( .C1(n15682), .C2(n20847), .A(n14662), .B(n14661), .ZN(
        P1_U2829) );
  INV_X1 U18234 ( .A(n14663), .ZN(n14667) );
  AOI21_X1 U18235 ( .B1(n14664), .B2(n14669), .A(n14665), .ZN(n14666) );
  INV_X1 U18236 ( .A(n16711), .ZN(n14685) );
  AOI22_X1 U18237 ( .A1(n15608), .A2(n15550), .B1(P1_EAX_REG_13__SCAN_IN), 
        .B2(n15606), .ZN(n14668) );
  OAI21_X1 U18238 ( .B1(n14685), .B2(n15610), .A(n14668), .ZN(P1_U2891) );
  XOR2_X1 U18239 ( .A(n14669), .B(n14664), .Z(n16716) );
  INV_X1 U18240 ( .A(n16716), .ZN(n14689) );
  NAND4_X1 U18241 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(P1_REIP_REG_9__SCAN_IN), 
        .A3(P1_REIP_REG_11__SCAN_IN), .A4(P1_REIP_REG_12__SCAN_IN), .ZN(n15441) );
  INV_X1 U18242 ( .A(n15441), .ZN(n14671) );
  AOI21_X1 U18243 ( .B1(n14671), .B2(n14670), .A(n15149), .ZN(n16628) );
  NAND3_X1 U18244 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(P1_REIP_REG_9__SCAN_IN), 
        .A3(P1_REIP_REG_11__SCAN_IN), .ZN(n14672) );
  INV_X1 U18245 ( .A(P1_REIP_REG_12__SCAN_IN), .ZN(n21217) );
  OAI21_X1 U18246 ( .B1(n14672), .B2(n16632), .A(n21217), .ZN(n14681) );
  OR2_X1 U18247 ( .A1(n14675), .A2(n14674), .ZN(n14676) );
  NAND2_X1 U18248 ( .A1(n14673), .A2(n14676), .ZN(n15791) );
  INV_X1 U18249 ( .A(n20816), .ZN(n20831) );
  AOI21_X1 U18250 ( .B1(n20849), .B2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n20831), .ZN(n14677) );
  OAI21_X1 U18251 ( .B1(n16714), .B2(n20847), .A(n14677), .ZN(n14678) );
  AOI21_X1 U18252 ( .B1(P1_EBX_REG_12__SCAN_IN), .B2(n20850), .A(n14678), .ZN(
        n14679) );
  OAI21_X1 U18253 ( .B1(n15791), .B2(n20860), .A(n14679), .ZN(n14680) );
  AOI21_X1 U18254 ( .B1(n16628), .B2(n14681), .A(n14680), .ZN(n14682) );
  OAI21_X1 U18255 ( .B1(n14689), .B2(n16617), .A(n14682), .ZN(P1_U2828) );
  INV_X1 U18256 ( .A(P1_EBX_REG_13__SCAN_IN), .ZN(n16621) );
  NAND2_X1 U18257 ( .A1(n14673), .A2(n14683), .ZN(n14684) );
  NAND2_X1 U18258 ( .A1(n15445), .A2(n14684), .ZN(n16788) );
  OAI222_X1 U18259 ( .A1(n14685), .A2(n16640), .B1(n16621), .B2(n16644), .C1(
        n16788), .C2(n15543), .ZN(P1_U2859) );
  INV_X1 U18260 ( .A(P1_EBX_REG_12__SCAN_IN), .ZN(n14686) );
  OAI222_X1 U18261 ( .A1(n14689), .A2(n16640), .B1(n16644), .B2(n14686), .C1(
        n15791), .C2(n15543), .ZN(P1_U2860) );
  MUX2_X1 U18262 ( .A(DATAI_12_), .B(BUF1_REG_12__SCAN_IN), .S(n14706), .Z(
        n20909) );
  INV_X1 U18263 ( .A(n20909), .ZN(n14688) );
  OAI222_X1 U18264 ( .A1(n14689), .A2(n15610), .B1(n15605), .B2(n14688), .C1(
        n14687), .C2(n15603), .ZN(P1_U2892) );
  INV_X1 U18265 ( .A(n19713), .ZN(n14700) );
  INV_X1 U18266 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n19488) );
  OAI21_X1 U18267 ( .B1(n19512), .B2(n19656), .A(n19488), .ZN(n14699) );
  NAND2_X1 U18268 ( .A1(n14691), .A2(n14699), .ZN(n19487) );
  NOR2_X1 U18269 ( .A1(n14700), .A2(n19487), .ZN(n14698) );
  INV_X1 U18270 ( .A(n14690), .ZN(n14696) );
  NAND2_X1 U18271 ( .A1(n19040), .A2(n18272), .ZN(n19539) );
  AOI21_X1 U18272 ( .B1(n14693), .B2(n19539), .A(n19698), .ZN(n18205) );
  NAND2_X1 U18273 ( .A1(n14694), .A2(n18205), .ZN(n14695) );
  NAND4_X1 U18274 ( .A1(n14696), .A2(n16523), .A3(n16455), .A4(n14695), .ZN(
        n19514) );
  INV_X1 U18275 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n19651) );
  NOR2_X1 U18276 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n19651), .ZN(n19036) );
  INV_X1 U18277 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n17270) );
  NAND3_X1 U18278 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_0__SCAN_IN), .A3(P3_STATE2_REG_2__SCAN_IN), .ZN(n19649)
         );
  NOR2_X1 U18279 ( .A1(n17270), .A2(n19649), .ZN(n14697) );
  AOI211_X2 U18280 ( .C1(n19694), .C2(n19514), .A(n19036), .B(n14697), .ZN(
        n19680) );
  MUX2_X1 U18281 ( .A(n14698), .B(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .S(
        n19680), .Z(P3_U3284) );
  NOR2_X1 U18282 ( .A1(n18002), .A2(n14699), .ZN(n19019) );
  NOR2_X1 U18283 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n19651), .ZN(
        n19675) );
  NOR2_X1 U18284 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n19703) );
  AOI21_X1 U18285 ( .B1(P3_STATE2_REG_2__SCAN_IN), .B2(
        P3_STATE2_REG_1__SCAN_IN), .A(n19703), .ZN(n19556) );
  OR2_X1 U18286 ( .A1(n19675), .A2(n19556), .ZN(n19035) );
  NAND2_X1 U18287 ( .A1(n19542), .A2(n19035), .ZN(n19065) );
  OAI221_X1 U18288 ( .B1(n19649), .B2(n19019), .C1(n19649), .C2(n17270), .A(
        n19065), .ZN(n19032) );
  INV_X1 U18289 ( .A(n19032), .ZN(n19022) );
  NAND2_X1 U18290 ( .A1(n19712), .A2(n19651), .ZN(n17265) );
  NAND2_X1 U18291 ( .A1(n14700), .A2(n17265), .ZN(n19020) );
  NAND2_X1 U18292 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n19023) );
  AOI22_X1 U18293 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P3_STATE2_REG_3__SCAN_IN), .B1(n19020), .B2(n19023), .ZN(n19027) );
  NOR2_X1 U18294 ( .A1(n19022), .A2(n19027), .ZN(n14702) );
  INV_X1 U18295 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n19699) );
  NOR3_X1 U18296 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .A3(n19699), .ZN(n19116) );
  INV_X1 U18297 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19325) );
  NAND2_X1 U18298 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n19325), .ZN(n19072) );
  NAND2_X1 U18299 ( .A1(n19072), .A2(n19032), .ZN(n19025) );
  OR2_X1 U18300 ( .A1(n19116), .A2(n19025), .ZN(n14701) );
  MUX2_X1 U18301 ( .A(n14702), .B(n14701), .S(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .Z(P3_U2864) );
  NAND3_X1 U18302 ( .A1(n15603), .A2(n14703), .A3(n14706), .ZN(n14876) );
  AOI22_X1 U18303 ( .A1(n15595), .A2(BUF1_REG_28__SCAN_IN), .B1(
        P1_EAX_REG_28__SCAN_IN), .B2(n15606), .ZN(n14709) );
  NOR3_X1 U18304 ( .A1(n15606), .A2(n14873), .A3(n14704), .ZN(n14705) );
  NOR3_X1 U18305 ( .A1(n15606), .A2(n14706), .A3(n11179), .ZN(n14707) );
  AOI22_X1 U18306 ( .A1(n15598), .A2(n20909), .B1(n15596), .B2(DATAI_28_), 
        .ZN(n14708) );
  OAI211_X1 U18307 ( .C1(n14731), .C2(n15610), .A(n14709), .B(n14708), .ZN(
        P1_U2876) );
  OR2_X1 U18308 ( .A1(n9788), .A2(n14710), .ZN(n14711) );
  NAND2_X1 U18309 ( .A1(n12130), .A2(n14711), .ZN(n15687) );
  OAI222_X1 U18310 ( .A1(n16640), .A2(n14731), .B1(n14725), .B2(n16644), .C1(
        n15687), .C2(n15543), .ZN(P1_U2844) );
  INV_X1 U18311 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n21234) );
  INV_X1 U18312 ( .A(P1_REIP_REG_17__SCAN_IN), .ZN(n21227) );
  INV_X1 U18313 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n21219) );
  INV_X1 U18314 ( .A(P1_REIP_REG_14__SCAN_IN), .ZN(n21222) );
  NOR4_X1 U18315 ( .A1(n14712), .A2(n15441), .A3(n21219), .A4(n21222), .ZN(
        n15442) );
  NAND2_X1 U18316 ( .A1(n15442), .A2(P1_REIP_REG_15__SCAN_IN), .ZN(n14715) );
  NOR2_X1 U18317 ( .A1(n20813), .A2(n14715), .ZN(n16598) );
  NAND2_X1 U18318 ( .A1(P1_REIP_REG_16__SCAN_IN), .A2(n16598), .ZN(n15436) );
  NAND4_X1 U18319 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(P1_REIP_REG_18__SCAN_IN), 
        .A3(P1_REIP_REG_20__SCAN_IN), .A4(n16594), .ZN(n16551) );
  NOR2_X1 U18320 ( .A1(n21234), .A2(n16551), .ZN(n16548) );
  NAND2_X1 U18321 ( .A1(P1_REIP_REG_24__SCAN_IN), .A2(P1_REIP_REG_25__SCAN_IN), 
        .ZN(n16527) );
  INV_X1 U18322 ( .A(n16527), .ZN(n14713) );
  NAND2_X1 U18323 ( .A1(n16539), .A2(n14713), .ZN(n15192) );
  INV_X1 U18324 ( .A(P1_REIP_REG_26__SCAN_IN), .ZN(n21242) );
  NOR2_X1 U18325 ( .A1(n15192), .A2(n21242), .ZN(n15152) );
  INV_X1 U18326 ( .A(n15152), .ZN(n15179) );
  NOR3_X1 U18327 ( .A1(n15179), .A2(P1_REIP_REG_28__SCAN_IN), .A3(n21245), 
        .ZN(n14729) );
  NAND2_X1 U18328 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(P1_REIP_REG_18__SCAN_IN), 
        .ZN(n16565) );
  INV_X1 U18329 ( .A(P1_REIP_REG_20__SCAN_IN), .ZN(n21232) );
  NOR2_X1 U18330 ( .A1(n16565), .A2(n21232), .ZN(n14716) );
  NAND3_X1 U18331 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(P1_REIP_REG_16__SCAN_IN), 
        .A3(n20845), .ZN(n14714) );
  OAI21_X1 U18332 ( .B1(n14715), .B2(n14714), .A(n15461), .ZN(n16574) );
  OAI21_X1 U18333 ( .B1(n14716), .B2(n20813), .A(n16574), .ZN(n16570) );
  NAND2_X1 U18334 ( .A1(P1_REIP_REG_22__SCAN_IN), .A2(P1_REIP_REG_23__SCAN_IN), 
        .ZN(n14717) );
  OAI21_X1 U18335 ( .B1(n21234), .B2(n14717), .A(n15461), .ZN(n14718) );
  INV_X1 U18336 ( .A(n14718), .ZN(n14719) );
  NOR2_X1 U18337 ( .A1(n16570), .A2(n14719), .ZN(n16547) );
  OAI21_X1 U18338 ( .B1(n21242), .B2(n16527), .A(n15461), .ZN(n14720) );
  AND2_X1 U18339 ( .A1(n16547), .A2(n14720), .ZN(n15172) );
  NAND2_X1 U18340 ( .A1(P1_REIP_REG_28__SCAN_IN), .A2(P1_REIP_REG_27__SCAN_IN), 
        .ZN(n14721) );
  NAND2_X1 U18341 ( .A1(n15461), .A2(n14721), .ZN(n14722) );
  AND2_X1 U18342 ( .A1(n15172), .A2(n14722), .ZN(n15166) );
  INV_X1 U18343 ( .A(P1_REIP_REG_28__SCAN_IN), .ZN(n21247) );
  NOR2_X1 U18344 ( .A1(n15166), .A2(n21247), .ZN(n14728) );
  NOR2_X1 U18345 ( .A1(n15687), .A2(n20860), .ZN(n14727) );
  AOI22_X1 U18346 ( .A1(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n20849), .B1(
        n16629), .B2(n14723), .ZN(n14724) );
  OAI21_X1 U18347 ( .B1(n16622), .B2(n14725), .A(n14724), .ZN(n14726) );
  NOR4_X1 U18348 ( .A1(n14729), .A2(n14728), .A3(n14727), .A4(n14726), .ZN(
        n14730) );
  OAI21_X1 U18349 ( .B1(n14731), .B2(n16617), .A(n14730), .ZN(P1_U2812) );
  AOI22_X1 U18350 ( .A1(n16933), .A2(BUF2_REG_31__SCAN_IN), .B1(
        P2_EAX_REG_31__SCAN_IN), .B2(n19974), .ZN(n14733) );
  NAND2_X1 U18351 ( .A1(n16932), .A2(BUF1_REG_31__SCAN_IN), .ZN(n14732) );
  OAI211_X1 U18352 ( .C1(n12097), .C2(n16023), .A(n14733), .B(n14732), .ZN(
        P2_U2888) );
  AOI21_X1 U18353 ( .B1(n14735), .B2(n13014), .A(n14734), .ZN(n15468) );
  AOI21_X1 U18354 ( .B1(n16734), .B2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n14736), .ZN(n14737) );
  OAI21_X1 U18355 ( .B1(n15163), .B2(n16743), .A(n14737), .ZN(n14738) );
  AOI21_X1 U18356 ( .B1(n15468), .B2(n16739), .A(n14738), .ZN(n14739) );
  OAI21_X1 U18357 ( .B1(n20773), .B2(n9785), .A(n14739), .ZN(P1_U2970) );
  INV_X1 U18358 ( .A(n14740), .ZN(n15824) );
  NOR2_X1 U18359 ( .A1(n15821), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n14741) );
  AOI21_X1 U18360 ( .B1(n12172), .B2(n15824), .A(n14741), .ZN(n16474) );
  INV_X1 U18361 ( .A(n16474), .ZN(n14743) );
  OAI22_X1 U18362 ( .A1(n16839), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n16498), .ZN(n14742) );
  AOI21_X1 U18363 ( .B1(n14743), .B2(n21270), .A(n14742), .ZN(n14747) );
  AOI21_X1 U18364 ( .B1(n9997), .B2(n21270), .A(n21275), .ZN(n14746) );
  OAI22_X1 U18365 ( .A1(n14747), .A2(n21275), .B1(n14746), .B2(n10100), .ZN(
        P1_U3474) );
  NOR2_X1 U18366 ( .A1(n14748), .A2(n16273), .ZN(n16081) );
  OAI21_X1 U18367 ( .B1(n16081), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n9964), .ZN(n16254) );
  NAND2_X1 U18368 ( .A1(n14749), .A2(n14750), .ZN(n14751) );
  AND2_X1 U18369 ( .A1(n15855), .A2(n14751), .ZN(n16902) );
  NOR2_X1 U18370 ( .A1(n12009), .A2(n20666), .ZN(n16255) );
  AOI21_X1 U18371 ( .B1(n20029), .B2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n16255), .ZN(n14752) );
  OAI21_X1 U18372 ( .B1(n20045), .B2(n16905), .A(n14752), .ZN(n14753) );
  AOI21_X1 U18373 ( .B1(n16902), .B2(n20051), .A(n14753), .ZN(n14759) );
  AND2_X1 U18374 ( .A1(n14754), .A2(n16075), .ZN(n14756) );
  OR2_X1 U18375 ( .A1(n14756), .A2(n14755), .ZN(n16260) );
  INV_X1 U18376 ( .A(n16974), .ZN(n20046) );
  NAND3_X1 U18377 ( .A1(n16260), .A2(n14757), .A3(n20046), .ZN(n14758) );
  OAI211_X1 U18378 ( .C1(n16254), .C2(n20043), .A(n14759), .B(n14758), .ZN(
        P2_U2991) );
  OAI22_X1 U18379 ( .A1(n16670), .A2(n14761), .B1(n16823), .B2(n21245), .ZN(
        n14762) );
  AOI21_X1 U18380 ( .B1(n16722), .B2(n15173), .A(n14762), .ZN(n14766) );
  AOI21_X1 U18381 ( .B1(n14764), .B2(n14763), .A(n13015), .ZN(n15472) );
  NAND2_X1 U18382 ( .A1(n15472), .A2(n16739), .ZN(n14765) );
  OAI211_X1 U18383 ( .C1(n14767), .C2(n20773), .A(n14766), .B(n14765), .ZN(
        P1_U2972) );
  NOR2_X1 U18384 ( .A1(n19969), .A2(n10570), .ZN(n14768) );
  OAI21_X1 U18385 ( .B1(n20131), .B2(n19959), .A(n14769), .ZN(P2_U2884) );
  XNOR2_X1 U18386 ( .A(n14771), .B(n14770), .ZN(n17060) );
  XNOR2_X1 U18387 ( .A(n14772), .B(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n14773) );
  XNOR2_X1 U18388 ( .A(n14774), .B(n14773), .ZN(n17062) );
  NAND2_X1 U18389 ( .A1(n17062), .A2(n20046), .ZN(n14779) );
  NAND2_X1 U18390 ( .A1(n17008), .A2(n14782), .ZN(n14777) );
  NOR2_X1 U18391 ( .A1(n20073), .A2(n14775), .ZN(n17057) );
  INV_X1 U18392 ( .A(n17057), .ZN(n14776) );
  OAI211_X1 U18393 ( .C1(n14786), .C2(n20055), .A(n14777), .B(n14776), .ZN(
        n14778) );
  OAI211_X1 U18394 ( .C1(n17060), .C2(n20043), .A(n14779), .B(n9841), .ZN(
        P2_U3011) );
  NAND2_X1 U18395 ( .A1(n9719), .A2(n14780), .ZN(n14781) );
  XNOR2_X1 U18396 ( .A(n14782), .B(n14781), .ZN(n14783) );
  NAND2_X1 U18397 ( .A1(n14783), .A2(n19897), .ZN(n14790) );
  AOI22_X1 U18398 ( .A1(n19917), .A2(P2_EBX_REG_3__SCAN_IN), .B1(n20700), .B2(
        n19915), .ZN(n14784) );
  OAI21_X1 U18399 ( .B1(n14785), .B2(n19919), .A(n14784), .ZN(n14788) );
  OAI22_X1 U18400 ( .A1(n14786), .A2(n19815), .B1(n14775), .B2(n19887), .ZN(
        n14787) );
  OAI211_X1 U18401 ( .C1(n19925), .C2(n20131), .A(n14790), .B(n14789), .ZN(
        P2_U2852) );
  INV_X1 U18402 ( .A(n16885), .ZN(n14795) );
  OAI21_X1 U18403 ( .B1(n20055), .B2(n10080), .A(n14792), .ZN(n14794) );
  NOR2_X1 U18404 ( .A1(n15909), .A2(n16202), .ZN(n14793) );
  AOI211_X1 U18405 ( .C1(n17008), .C2(n14795), .A(n14794), .B(n14793), .ZN(
        n14796) );
  OAI211_X1 U18406 ( .C1(n20043), .C2(n14798), .A(n14797), .B(n14796), .ZN(
        P2_U2987) );
  XOR2_X1 U18407 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .B(n14802), .Z(
        n14803) );
  XNOR2_X1 U18408 ( .A(n14804), .B(n14803), .ZN(n14848) );
  INV_X1 U18409 ( .A(n14846), .ZN(n14813) );
  NOR2_X1 U18410 ( .A1(n14807), .A2(n14806), .ZN(n16208) );
  AOI21_X1 U18411 ( .B1(n14809), .B2(n14808), .A(n15894), .ZN(n16869) );
  NOR2_X1 U18412 ( .A1(n12009), .A2(n20676), .ZN(n14844) );
  NAND2_X1 U18413 ( .A1(n13039), .A2(n14810), .ZN(n14811) );
  NAND2_X1 U18414 ( .A1(n15932), .A2(n14811), .ZN(n16867) );
  OR3_X1 U18415 ( .A1(n14812), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        n10829), .ZN(n16207) );
  OAI21_X1 U18416 ( .B1(n14848), .B2(n17071), .A(n14814), .ZN(P2_U3018) );
  MUX2_X1 U18417 ( .A(n14816), .B(n12132), .S(n14815), .Z(n14820) );
  AOI22_X1 U18418 ( .A1(n14818), .A2(P1_EBX_REG_31__SCAN_IN), .B1(n14817), 
        .B2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14819) );
  INV_X1 U18419 ( .A(n15467), .ZN(n14825) );
  NOR3_X1 U18420 ( .A1(n14822), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n14821), .ZN(n14824) );
  NAND3_X1 U18421 ( .A1(n14827), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n14826), .ZN(n14828) );
  OAI211_X1 U18422 ( .C1(n14830), .C2(n16792), .A(n14829), .B(n14828), .ZN(
        P1_U3000) );
  NAND2_X1 U18423 ( .A1(n14831), .A2(n20855), .ZN(n14843) );
  NAND2_X1 U18424 ( .A1(n20850), .A2(P1_EBX_REG_2__SCAN_IN), .ZN(n14839) );
  AOI22_X1 U18425 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(n14833), .B1(
        P1_REIP_REG_2__SCAN_IN), .B2(n14832), .ZN(n14838) );
  INV_X1 U18426 ( .A(n14834), .ZN(n14835) );
  NAND2_X1 U18427 ( .A1(n16629), .A2(n14835), .ZN(n14837) );
  NAND2_X1 U18428 ( .A1(n20849), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n14836) );
  NAND4_X1 U18429 ( .A1(n14839), .A2(n14838), .A3(n14837), .A4(n14836), .ZN(
        n14840) );
  AOI21_X1 U18430 ( .B1(n16609), .B2(n14841), .A(n14840), .ZN(n14842) );
  OAI211_X1 U18431 ( .C1(n20853), .C2(n9734), .A(n14843), .B(n14842), .ZN(
        P1_U2838) );
  AOI21_X1 U18432 ( .B1(n20029), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n14844), .ZN(n14845) );
  OAI21_X1 U18433 ( .B1(n20045), .B2(n16872), .A(n14845), .ZN(n14847) );
  XNOR2_X1 U18434 ( .A(n19953), .B(n19952), .ZN(n14850) );
  MUX2_X1 U18435 ( .A(n10717), .B(n17036), .S(n19969), .Z(n14849) );
  OAI21_X1 U18436 ( .B1(n14850), .B2(n19959), .A(n14849), .ZN(P2_U2877) );
  XOR2_X1 U18437 ( .A(n14851), .B(P2_INSTQUEUE_REG_0__5__SCAN_IN), .Z(n14855)
         );
  NOR2_X1 U18438 ( .A1(n19969), .A2(n14852), .ZN(n14853) );
  AOI21_X1 U18439 ( .B1(n19909), .B2(n19969), .A(n14853), .ZN(n14854) );
  OAI21_X1 U18440 ( .B1(n14855), .B2(n19959), .A(n14854), .ZN(P2_U2882) );
  NOR2_X1 U18441 ( .A1(n14857), .A2(n14856), .ZN(n14858) );
  OR2_X1 U18442 ( .A1(n14267), .A2(n14858), .ZN(n20063) );
  NOR2_X1 U18443 ( .A1(n20063), .A2(n19947), .ZN(n14859) );
  AOI21_X1 U18444 ( .B1(P2_EBX_REG_4__SCAN_IN), .B2(n19947), .A(n14859), .ZN(
        n14860) );
  OAI21_X1 U18445 ( .B1(n19983), .B2(n19959), .A(n14860), .ZN(P2_U2883) );
  INV_X1 U18446 ( .A(n20041), .ZN(n14864) );
  NOR2_X1 U18447 ( .A1(n9766), .A2(n14861), .ZN(n14863) );
  INV_X1 U18448 ( .A(n19910), .ZN(n20613) );
  AOI21_X1 U18449 ( .B1(n14864), .B2(n14863), .A(n20613), .ZN(n14862) );
  OAI21_X1 U18450 ( .B1(n14864), .B2(n14863), .A(n14862), .ZN(n14872) );
  INV_X1 U18451 ( .A(n20063), .ZN(n20038) );
  INV_X1 U18452 ( .A(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n14866) );
  AOI22_X1 U18453 ( .A1(P2_EBX_REG_4__SCAN_IN), .A2(n19917), .B1(n19915), .B2(
        n20056), .ZN(n14865) );
  OAI211_X1 U18454 ( .C1(n14866), .C2(n19815), .A(n20073), .B(n14865), .ZN(
        n14867) );
  AOI21_X1 U18455 ( .B1(n14868), .B2(n19877), .A(n14867), .ZN(n14869) );
  OAI21_X1 U18456 ( .B1(n19887), .B2(n10921), .A(n14869), .ZN(n14870) );
  AOI21_X1 U18457 ( .B1(n19922), .B2(n20038), .A(n14870), .ZN(n14871) );
  OAI211_X1 U18458 ( .C1(n19925), .C2(n19983), .A(n14872), .B(n14871), .ZN(
        P2_U2851) );
  INV_X1 U18459 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n17173) );
  NAND3_X1 U18460 ( .A1(n15148), .A2(n14873), .A3(n15603), .ZN(n14875) );
  AOI22_X1 U18461 ( .A1(n15596), .A2(DATAI_31_), .B1(P1_EAX_REG_31__SCAN_IN), 
        .B2(n15606), .ZN(n14874) );
  OAI211_X1 U18462 ( .C1(n14876), .C2(n17173), .A(n14875), .B(n14874), .ZN(
        P1_U2873) );
  OAI22_X1 U18463 ( .A1(n9719), .A2(n14877), .B1(n19933), .B2(n9766), .ZN(
        n16425) );
  INV_X1 U18464 ( .A(n16425), .ZN(n14881) );
  INV_X1 U18465 ( .A(n14878), .ZN(n14880) );
  AOI222_X1 U18466 ( .A1(n14881), .A2(P2_STATE2_REG_1__SCAN_IN), .B1(n14880), 
        .B2(n17082), .C1(n14879), .C2(n16433), .ZN(n14884) );
  AOI21_X1 U18467 ( .B1(n16433), .B2(n11732), .A(n16439), .ZN(n14883) );
  OAI22_X1 U18468 ( .A1(n14884), .A2(n16439), .B1(n14883), .B2(n14882), .ZN(
        P2_U3601) );
  NAND2_X1 U18469 ( .A1(n10631), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n14889) );
  NAND2_X1 U18470 ( .A1(n14951), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n14888) );
  AOI22_X1 U18471 ( .A1(n10500), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n14885), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n14887) );
  NAND2_X1 U18472 ( .A1(n10507), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n14886) );
  AND4_X1 U18473 ( .A1(n14889), .A2(n14888), .A3(n14887), .A4(n14886), .ZN(
        n14902) );
  AOI22_X1 U18474 ( .A1(n14957), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n14956), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n14901) );
  NAND2_X1 U18475 ( .A1(n10499), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n14891) );
  NAND2_X1 U18476 ( .A1(n10498), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n14890) );
  OAI211_X1 U18477 ( .C1(n14961), .C2(n14892), .A(n14891), .B(n14890), .ZN(
        n14895) );
  OAI22_X1 U18478 ( .A1(n14964), .A2(n14893), .B1(n14962), .B2(n15091), .ZN(
        n14894) );
  NOR2_X1 U18479 ( .A1(n14895), .A2(n14894), .ZN(n14900) );
  AOI22_X1 U18480 ( .A1(n14967), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n11881), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n14897) );
  NAND2_X1 U18481 ( .A1(n14450), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n14896) );
  OAI211_X1 U18482 ( .C1(n15092), .C2(n14473), .A(n14897), .B(n14896), .ZN(
        n14898) );
  INV_X1 U18483 ( .A(n14898), .ZN(n14899) );
  NAND4_X1 U18484 ( .A1(n14902), .A2(n14901), .A3(n14900), .A4(n14899), .ZN(
        n15998) );
  NAND2_X1 U18485 ( .A1(n10631), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n14907) );
  NAND2_X1 U18486 ( .A1(n14951), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n14906) );
  AOI22_X1 U18487 ( .A1(n10500), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n14885), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n14905) );
  NAND2_X1 U18488 ( .A1(n10507), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n14904) );
  NAND4_X1 U18489 ( .A1(n14907), .A2(n14906), .A3(n14905), .A4(n14904), .ZN(
        n14916) );
  AOI22_X1 U18490 ( .A1(n10498), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n10499), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n14914) );
  NAND2_X1 U18491 ( .A1(n14908), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n14913) );
  NAND2_X1 U18492 ( .A1(n14909), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n14912) );
  NAND2_X1 U18493 ( .A1(n14910), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n14911) );
  NAND4_X1 U18494 ( .A1(n14914), .A2(n14913), .A3(n14912), .A4(n14911), .ZN(
        n14915) );
  NOR2_X1 U18495 ( .A1(n14916), .A2(n14915), .ZN(n14926) );
  OAI22_X1 U18496 ( .A1(n14919), .A2(n14918), .B1(n14917), .B2(n15104), .ZN(
        n14924) );
  AOI22_X1 U18497 ( .A1(n14967), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n11881), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n14921) );
  NAND2_X1 U18498 ( .A1(n14450), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n14920) );
  OAI211_X1 U18499 ( .C1(n14922), .C2(n14473), .A(n14921), .B(n14920), .ZN(
        n14923) );
  NOR2_X1 U18500 ( .A1(n14924), .A2(n14923), .ZN(n14925) );
  AND2_X1 U18501 ( .A1(n14926), .A2(n14925), .ZN(n15929) );
  AOI22_X1 U18502 ( .A1(n9761), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10462), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n14941) );
  AOI22_X1 U18503 ( .A1(n15129), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n14989), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n14940) );
  AOI22_X1 U18504 ( .A1(n10445), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n13745), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n14939) );
  INV_X1 U18505 ( .A(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n14936) );
  INV_X1 U18506 ( .A(n10317), .ZN(n15127) );
  INV_X1 U18507 ( .A(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n14931) );
  OR2_X1 U18508 ( .A1(n15127), .A2(n14931), .ZN(n14935) );
  INV_X1 U18509 ( .A(n14932), .ZN(n14934) );
  NAND2_X1 U18510 ( .A1(n14934), .A2(n14933), .ZN(n15125) );
  OAI211_X1 U18511 ( .C1(n14929), .C2(n14936), .A(n14935), .B(n15125), .ZN(
        n14937) );
  INV_X1 U18512 ( .A(n14937), .ZN(n14938) );
  NAND4_X1 U18513 ( .A1(n14941), .A2(n14940), .A3(n14939), .A4(n14938), .ZN(
        n14950) );
  AOI22_X1 U18514 ( .A1(n9761), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n10462), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n14948) );
  AOI22_X1 U18515 ( .A1(n15129), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n14989), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n14947) );
  AOI22_X1 U18516 ( .A1(n10445), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n13745), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n14946) );
  NAND2_X1 U18517 ( .A1(n10446), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n14942) );
  INV_X1 U18518 ( .A(n15125), .ZN(n15089) );
  OAI211_X1 U18519 ( .C1(n15127), .C2(n14943), .A(n14942), .B(n15089), .ZN(
        n14944) );
  INV_X1 U18520 ( .A(n14944), .ZN(n14945) );
  NAND4_X1 U18521 ( .A1(n14948), .A2(n14947), .A3(n14946), .A4(n14945), .ZN(
        n14949) );
  NAND2_X1 U18522 ( .A1(n14950), .A2(n14949), .ZN(n14980) );
  NOR2_X1 U18523 ( .A1(n9759), .A2(n14980), .ZN(n14978) );
  NAND2_X1 U18524 ( .A1(n10631), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n14955) );
  NAND2_X1 U18525 ( .A1(n14951), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n14954) );
  AOI22_X1 U18526 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n10500), .B1(
        n14885), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n14953) );
  NAND2_X1 U18527 ( .A1(n10507), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n14952) );
  AND4_X1 U18528 ( .A1(n14955), .A2(n14954), .A3(n14953), .A4(n14952), .ZN(
        n14975) );
  AOI22_X1 U18529 ( .A1(n14957), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n14956), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n14974) );
  INV_X1 U18530 ( .A(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n14960) );
  NAND2_X1 U18531 ( .A1(n10499), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n14959) );
  NAND2_X1 U18532 ( .A1(n10498), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n14958) );
  OAI211_X1 U18533 ( .C1(n14961), .C2(n14960), .A(n14959), .B(n14958), .ZN(
        n14966) );
  INV_X1 U18534 ( .A(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n20448) );
  OAI22_X1 U18535 ( .A1(n14964), .A2(n14963), .B1(n14962), .B2(n20448), .ZN(
        n14965) );
  NOR2_X1 U18536 ( .A1(n14966), .A2(n14965), .ZN(n14973) );
  AOI22_X1 U18537 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n14967), .B1(
        n11881), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n14969) );
  NAND2_X1 U18538 ( .A1(n14450), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n14968) );
  OAI211_X1 U18539 ( .C1(n14473), .C2(n14970), .A(n14969), .B(n14968), .ZN(
        n14971) );
  INV_X1 U18540 ( .A(n14971), .ZN(n14972) );
  NAND4_X1 U18541 ( .A1(n14975), .A2(n14974), .A3(n14973), .A4(n14972), .ZN(
        n14977) );
  INV_X1 U18542 ( .A(n14980), .ZN(n14976) );
  NAND2_X1 U18543 ( .A1(n14977), .A2(n14976), .ZN(n15002) );
  OAI22_X1 U18544 ( .A1(n14978), .A2(n14977), .B1(n9759), .B2(n15002), .ZN(
        n15004) );
  INV_X1 U18545 ( .A(n15004), .ZN(n14979) );
  NOR2_X1 U18546 ( .A1(n20755), .A2(n14980), .ZN(n15921) );
  AOI22_X1 U18547 ( .A1(n9761), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n10462), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n14988) );
  AOI22_X1 U18548 ( .A1(n15129), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n14989), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n14987) );
  AOI22_X1 U18549 ( .A1(n10445), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n9758), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n14986) );
  INV_X1 U18550 ( .A(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n14983) );
  OR2_X1 U18551 ( .A1(n15127), .A2(n14981), .ZN(n14982) );
  OAI211_X1 U18552 ( .C1(n15122), .C2(n14983), .A(n14982), .B(n15125), .ZN(
        n14984) );
  INV_X1 U18553 ( .A(n14984), .ZN(n14985) );
  NAND4_X1 U18554 ( .A1(n14988), .A2(n14987), .A3(n14986), .A4(n14985), .ZN(
        n14999) );
  AOI22_X1 U18555 ( .A1(n15129), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n15130), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n14997) );
  AOI22_X1 U18556 ( .A1(n10445), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n13745), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n14996) );
  AOI22_X1 U18557 ( .A1(n9761), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n9747), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n14995) );
  NAND2_X1 U18558 ( .A1(n10446), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n14990) );
  OAI211_X1 U18559 ( .C1(n14992), .C2(n14991), .A(n14990), .B(n15089), .ZN(
        n14993) );
  INV_X1 U18560 ( .A(n14993), .ZN(n14994) );
  NAND4_X1 U18561 ( .A1(n14997), .A2(n14996), .A3(n14995), .A4(n14994), .ZN(
        n14998) );
  AND2_X1 U18562 ( .A1(n14999), .A2(n14998), .ZN(n15000) );
  INV_X1 U18563 ( .A(n15000), .ZN(n16910) );
  INV_X1 U18564 ( .A(n15002), .ZN(n15001) );
  AND2_X1 U18565 ( .A1(n15001), .A2(n15000), .ZN(n15006) );
  AOI211_X1 U18566 ( .C1(n16910), .C2(n15002), .A(n15047), .B(n15006), .ZN(
        n16912) );
  INV_X1 U18567 ( .A(n15921), .ZN(n15003) );
  NOR3_X1 U18568 ( .A1(n15004), .A2(n16910), .A3(n15003), .ZN(n15005) );
  INV_X1 U18569 ( .A(n15006), .ZN(n15023) );
  AOI22_X1 U18570 ( .A1(n9761), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n10462), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n15013) );
  AOI22_X1 U18571 ( .A1(n15129), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n15130), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n15012) );
  AOI22_X1 U18572 ( .A1(n10445), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n13745), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n15011) );
  INV_X1 U18573 ( .A(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n15008) );
  NAND2_X1 U18574 ( .A1(n9747), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(
        n15007) );
  OAI211_X1 U18575 ( .C1(n14930), .C2(n15008), .A(n15007), .B(n15125), .ZN(
        n15009) );
  INV_X1 U18576 ( .A(n15009), .ZN(n15010) );
  NAND4_X1 U18577 ( .A1(n15013), .A2(n15012), .A3(n15011), .A4(n15010), .ZN(
        n15022) );
  AOI22_X1 U18578 ( .A1(n9761), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n10462), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n15020) );
  AOI22_X1 U18579 ( .A1(n15129), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n15130), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n15019) );
  AOI22_X1 U18580 ( .A1(n10445), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n13745), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n15018) );
  INV_X1 U18581 ( .A(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n15015) );
  NAND2_X1 U18582 ( .A1(n9757), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n15014) );
  OAI211_X1 U18583 ( .C1(n15127), .C2(n15015), .A(n15014), .B(n15089), .ZN(
        n15016) );
  INV_X1 U18584 ( .A(n15016), .ZN(n15017) );
  NAND4_X1 U18585 ( .A1(n15020), .A2(n15019), .A3(n15018), .A4(n15017), .ZN(
        n15021) );
  NAND2_X1 U18586 ( .A1(n15022), .A2(n15021), .ZN(n15025) );
  OR2_X1 U18587 ( .A1(n15023), .A2(n15025), .ZN(n15049) );
  NAND2_X1 U18588 ( .A1(n15023), .A2(n15025), .ZN(n15024) );
  NAND3_X1 U18589 ( .A1(n15049), .A2(n15073), .A3(n15024), .ZN(n15027) );
  INV_X1 U18590 ( .A(n15025), .ZN(n15026) );
  NAND2_X1 U18591 ( .A1(n9759), .A2(n15026), .ZN(n15917) );
  INV_X1 U18592 ( .A(n15049), .ZN(n15046) );
  AOI22_X1 U18593 ( .A1(n9761), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n10462), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n15036) );
  AOI22_X1 U18594 ( .A1(n15129), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n15130), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n15035) );
  AOI22_X1 U18595 ( .A1(n10445), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n9757), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n15034) );
  OR2_X1 U18596 ( .A1(n15127), .A2(n15029), .ZN(n15030) );
  OAI211_X1 U18597 ( .C1(n15122), .C2(n15031), .A(n15030), .B(n15125), .ZN(
        n15032) );
  INV_X1 U18598 ( .A(n15032), .ZN(n15033) );
  NAND4_X1 U18599 ( .A1(n15036), .A2(n15035), .A3(n15034), .A4(n15033), .ZN(
        n15045) );
  OR2_X1 U18600 ( .A1(n15127), .A2(n15037), .ZN(n15038) );
  OAI211_X1 U18601 ( .C1(n15083), .C2(n10416), .A(n15089), .B(n15038), .ZN(
        n15039) );
  INV_X1 U18602 ( .A(n15039), .ZN(n15043) );
  AOI22_X1 U18603 ( .A1(n10445), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n10446), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n15042) );
  AOI22_X1 U18604 ( .A1(n9761), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n13745), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n15041) );
  AOI22_X1 U18605 ( .A1(n10462), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n15130), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n15040) );
  NAND4_X1 U18606 ( .A1(n15043), .A2(n15042), .A3(n15041), .A4(n15040), .ZN(
        n15044) );
  AND2_X1 U18607 ( .A1(n15045), .A2(n15044), .ZN(n15051) );
  NAND2_X1 U18608 ( .A1(n15046), .A2(n15051), .ZN(n15055) );
  INV_X1 U18609 ( .A(n15051), .ZN(n15048) );
  AOI21_X1 U18610 ( .B1(n15049), .B2(n15048), .A(n15047), .ZN(n15050) );
  NAND2_X1 U18611 ( .A1(n9759), .A2(n15051), .ZN(n15913) );
  INV_X1 U18612 ( .A(n15912), .ZN(n15054) );
  INV_X1 U18613 ( .A(n15055), .ZN(n15074) );
  AOI22_X1 U18614 ( .A1(n9761), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n10462), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n15063) );
  AOI22_X1 U18615 ( .A1(n15129), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n15130), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n15062) );
  AOI22_X1 U18616 ( .A1(n10445), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n13745), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n15061) );
  INV_X1 U18617 ( .A(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n15058) );
  INV_X1 U18618 ( .A(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n15056) );
  OR2_X1 U18619 ( .A1(n15127), .A2(n15056), .ZN(n15057) );
  OAI211_X1 U18620 ( .C1(n14930), .C2(n15058), .A(n15057), .B(n15125), .ZN(
        n15059) );
  INV_X1 U18621 ( .A(n15059), .ZN(n15060) );
  NAND4_X1 U18622 ( .A1(n15063), .A2(n15062), .A3(n15061), .A4(n15060), .ZN(
        n15072) );
  AOI22_X1 U18623 ( .A1(n9761), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n10462), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n15070) );
  AOI22_X1 U18624 ( .A1(n15129), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n15130), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n15069) );
  AOI22_X1 U18625 ( .A1(n10445), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n13745), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n15068) );
  INV_X1 U18626 ( .A(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n15065) );
  NAND2_X1 U18627 ( .A1(n10446), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n15064) );
  OAI211_X1 U18628 ( .C1(n15127), .C2(n15065), .A(n15064), .B(n15089), .ZN(
        n15066) );
  INV_X1 U18629 ( .A(n15066), .ZN(n15067) );
  NAND4_X1 U18630 ( .A1(n15070), .A2(n15069), .A3(n15068), .A4(n15067), .ZN(
        n15071) );
  AND2_X1 U18631 ( .A1(n15072), .A2(n15071), .ZN(n15079) );
  NAND2_X1 U18632 ( .A1(n15074), .A2(n15079), .ZN(n15897) );
  OAI211_X1 U18633 ( .C1(n15074), .C2(n15079), .A(n15073), .B(n15897), .ZN(
        n15076) );
  INV_X1 U18634 ( .A(n15076), .ZN(n15077) );
  NAND2_X1 U18635 ( .A1(n9759), .A2(n15079), .ZN(n15905) );
  OAI21_X1 U18636 ( .B1(n15127), .B2(n15080), .A(n15125), .ZN(n15085) );
  OAI22_X1 U18637 ( .A1(n15083), .A2(n15082), .B1(n15122), .B2(n15081), .ZN(
        n15084) );
  AOI211_X1 U18638 ( .C1(n9757), .C2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A(
        n15085), .B(n15084), .ZN(n15088) );
  AOI22_X1 U18639 ( .A1(n9761), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10462), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n15087) );
  AOI22_X1 U18640 ( .A1(n10445), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n15130), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n15086) );
  NAND3_X1 U18641 ( .A1(n15088), .A2(n15087), .A3(n15086), .ZN(n15099) );
  OAI21_X1 U18642 ( .B1(n15127), .B2(n15090), .A(n15089), .ZN(n15094) );
  OAI22_X1 U18643 ( .A1(n14928), .A2(n15092), .B1(n15122), .B2(n15091), .ZN(
        n15093) );
  AOI211_X1 U18644 ( .C1(n9758), .C2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A(
        n15094), .B(n15093), .ZN(n15097) );
  AOI22_X1 U18645 ( .A1(n9761), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n10462), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n15096) );
  AOI22_X1 U18646 ( .A1(n15129), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n15130), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n15095) );
  NAND3_X1 U18647 ( .A1(n15097), .A2(n15096), .A3(n15095), .ZN(n15098) );
  AND2_X1 U18648 ( .A1(n15099), .A2(n15098), .ZN(n15116) );
  AOI22_X1 U18649 ( .A1(n9761), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n10462), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n15101) );
  AOI22_X1 U18650 ( .A1(n15129), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n15130), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n15100) );
  NAND2_X1 U18651 ( .A1(n15101), .A2(n15100), .ZN(n15115) );
  AOI22_X1 U18652 ( .A1(n10445), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n13745), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n15103) );
  AOI21_X1 U18653 ( .B1(n10317), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A(
        n15125), .ZN(n15102) );
  OAI211_X1 U18654 ( .C1(n14930), .C2(n15104), .A(n15103), .B(n15102), .ZN(
        n15114) );
  OAI21_X1 U18655 ( .B1(n15127), .B2(n15105), .A(n15125), .ZN(n15109) );
  OAI22_X1 U18656 ( .A1(n14928), .A2(n15107), .B1(n15122), .B2(n15106), .ZN(
        n15108) );
  AOI211_X1 U18657 ( .C1(n10446), .C2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A(
        n15109), .B(n15108), .ZN(n15112) );
  AOI22_X1 U18658 ( .A1(n9761), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n10462), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n15111) );
  AOI22_X1 U18659 ( .A1(n15129), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n15130), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n15110) );
  NAND3_X1 U18660 ( .A1(n15112), .A2(n15111), .A3(n15110), .ZN(n15113) );
  OAI21_X1 U18661 ( .B1(n15115), .B2(n15114), .A(n15113), .ZN(n15118) );
  INV_X1 U18662 ( .A(n15116), .ZN(n15900) );
  NOR3_X1 U18663 ( .A1(n15897), .A2(n9759), .A3(n15900), .ZN(n15117) );
  XOR2_X1 U18664 ( .A(n15118), .B(n15117), .Z(n15890) );
  INV_X1 U18665 ( .A(n15117), .ZN(n15119) );
  AOI22_X1 U18666 ( .A1(n10445), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n9758), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n15121) );
  AOI21_X1 U18667 ( .B1(n9747), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A(
        n15125), .ZN(n15120) );
  OAI211_X1 U18668 ( .C1(n15122), .C2(n20448), .A(n15121), .B(n15120), .ZN(
        n15137) );
  AOI22_X1 U18669 ( .A1(n9761), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n10462), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n15124) );
  AOI22_X1 U18670 ( .A1(n15129), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n15130), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n15123) );
  NAND2_X1 U18671 ( .A1(n15124), .A2(n15123), .ZN(n15136) );
  INV_X1 U18672 ( .A(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n15126) );
  OAI21_X1 U18673 ( .B1(n15127), .B2(n15126), .A(n15125), .ZN(n15128) );
  AOI21_X1 U18674 ( .B1(n10445), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A(
        n15128), .ZN(n15134) );
  AOI22_X1 U18675 ( .A1(n15129), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n9761), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n15133) );
  AOI22_X1 U18676 ( .A1(n10462), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n15130), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n15132) );
  AOI22_X1 U18677 ( .A1(n13745), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n10446), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n15131) );
  NAND4_X1 U18678 ( .A1(n15134), .A2(n15133), .A3(n15132), .A4(n15131), .ZN(
        n15135) );
  OAI21_X1 U18679 ( .B1(n15137), .B2(n15136), .A(n15135), .ZN(n15138) );
  INV_X1 U18680 ( .A(n15138), .ZN(n15139) );
  NOR2_X1 U18681 ( .A1(n16845), .A2(n19947), .ZN(n15141) );
  AOI21_X1 U18682 ( .B1(P2_EBX_REG_30__SCAN_IN), .B2(n19947), .A(n15141), .ZN(
        n15142) );
  OAI21_X1 U18683 ( .B1(n15147), .B2(n19959), .A(n15142), .ZN(P2_U2857) );
  OAI22_X1 U18684 ( .A1(n16930), .A2(n19970), .B1(n19979), .B2(n13238), .ZN(
        n15143) );
  AOI21_X1 U18685 ( .B1(n16932), .B2(BUF1_REG_30__SCAN_IN), .A(n15143), .ZN(
        n15146) );
  AOI22_X1 U18686 ( .A1(n15144), .A2(n16935), .B1(n16933), .B2(
        BUF2_REG_30__SCAN_IN), .ZN(n15145) );
  OAI211_X1 U18687 ( .C1(n15147), .C2(n19982), .A(n15146), .B(n15145), .ZN(
        P2_U2889) );
  NAND2_X1 U18688 ( .A1(n15148), .A2(n20808), .ZN(n15157) );
  NAND2_X1 U18689 ( .A1(P1_REIP_REG_29__SCAN_IN), .A2(P1_REIP_REG_30__SCAN_IN), 
        .ZN(n15153) );
  INV_X1 U18690 ( .A(n15153), .ZN(n15150) );
  OAI21_X1 U18691 ( .B1(n15150), .B2(n15149), .A(n15166), .ZN(n15162) );
  OAI22_X1 U18692 ( .A1(n16622), .A2(n15466), .B1(n15151), .B2(n20818), .ZN(
        n15155) );
  NAND3_X1 U18693 ( .A1(n15152), .A2(P1_REIP_REG_27__SCAN_IN), .A3(
        P1_REIP_REG_28__SCAN_IN), .ZN(n15171) );
  NOR3_X1 U18694 ( .A1(n15171), .A2(P1_REIP_REG_31__SCAN_IN), .A3(n15153), 
        .ZN(n15154) );
  AOI211_X1 U18695 ( .C1(P1_REIP_REG_31__SCAN_IN), .C2(n15162), .A(n15155), 
        .B(n15154), .ZN(n15156) );
  OAI211_X1 U18696 ( .C1(n15467), .C2(n20860), .A(n15157), .B(n15156), .ZN(
        P1_U2809) );
  OAI21_X1 U18697 ( .B1(n15171), .B2(n21251), .A(n15158), .ZN(n15161) );
  AOI22_X1 U18698 ( .A1(n15616), .A2(n16629), .B1(n20849), .B2(
        P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n15159) );
  NAND2_X1 U18699 ( .A1(n15468), .A2(n20808), .ZN(n15170) );
  INV_X1 U18700 ( .A(n15163), .ZN(n15164) );
  AOI22_X1 U18701 ( .A1(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n20849), .B1(
        n16629), .B2(n15164), .ZN(n15165) );
  OAI21_X1 U18702 ( .B1(n16622), .B2(n15471), .A(n15165), .ZN(n15168) );
  NOR2_X1 U18703 ( .A1(n15166), .A2(n21251), .ZN(n15167) );
  AOI211_X1 U18704 ( .C1(n15469), .C2(n16609), .A(n15168), .B(n15167), .ZN(
        n15169) );
  OAI211_X1 U18705 ( .C1(P1_REIP_REG_29__SCAN_IN), .C2(n15171), .A(n15170), 
        .B(n15169), .ZN(P1_U2811) );
  NAND2_X1 U18706 ( .A1(n15472), .A2(n20808), .ZN(n15178) );
  INV_X1 U18707 ( .A(n15172), .ZN(n15190) );
  INV_X1 U18708 ( .A(P1_EBX_REG_27__SCAN_IN), .ZN(n15474) );
  AOI22_X1 U18709 ( .A1(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n20849), .B1(
        n16629), .B2(n15173), .ZN(n15174) );
  OAI21_X1 U18710 ( .B1(n16622), .B2(n15474), .A(n15174), .ZN(n15176) );
  NOR2_X1 U18711 ( .A1(n15473), .A2(n20860), .ZN(n15175) );
  AOI211_X1 U18712 ( .C1(P1_REIP_REG_27__SCAN_IN), .C2(n15190), .A(n15176), 
        .B(n15175), .ZN(n15177) );
  OAI211_X1 U18713 ( .C1(P1_REIP_REG_27__SCAN_IN), .C2(n15179), .A(n15178), 
        .B(n15177), .ZN(P1_U2813) );
  INV_X1 U18714 ( .A(n14763), .ZN(n15181) );
  AOI21_X1 U18715 ( .B1(n15182), .B2(n15180), .A(n15181), .ZN(n15621) );
  INV_X1 U18716 ( .A(n15481), .ZN(n15186) );
  INV_X1 U18717 ( .A(n15183), .ZN(n15185) );
  OAI21_X1 U18718 ( .B1(n15186), .B2(n15185), .A(n15184), .ZN(n15475) );
  AOI22_X1 U18719 ( .A1(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n20849), .B1(
        n16629), .B2(n15624), .ZN(n15188) );
  NAND2_X1 U18720 ( .A1(n20850), .A2(P1_EBX_REG_26__SCAN_IN), .ZN(n15187) );
  OAI211_X1 U18721 ( .C1(n15475), .C2(n20860), .A(n15188), .B(n15187), .ZN(
        n15189) );
  AOI21_X1 U18722 ( .B1(P1_REIP_REG_26__SCAN_IN), .B2(n15190), .A(n15189), 
        .ZN(n15191) );
  OAI21_X1 U18723 ( .B1(P1_REIP_REG_26__SCAN_IN), .B2(n15192), .A(n15191), 
        .ZN(n15193) );
  AOI21_X1 U18724 ( .B1(n15621), .B2(n20808), .A(n15193), .ZN(n15427) );
  NAND4_X1 U18725 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_4__7__SCAN_IN), .A3(P2_ADDRESS_REG_21__SCAN_IN), .A4(
        P1_D_C_N_REG_SCAN_IN), .ZN(n15197) );
  NAND4_X1 U18726 ( .A1(P2_DATAO_REG_17__SCAN_IN), .A2(
        P3_INSTQUEUE_REG_7__5__SCAN_IN), .A3(BUF2_REG_22__SCAN_IN), .A4(
        P3_EBX_REG_16__SCAN_IN), .ZN(n15196) );
  NAND4_X1 U18727 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(
        READY22_REG_SCAN_IN), .A3(P3_INSTQUEUE_REG_0__5__SCAN_IN), .A4(
        P3_UWORD_REG_6__SCAN_IN), .ZN(n15195) );
  NAND4_X1 U18728 ( .A1(P2_LWORD_REG_7__SCAN_IN), .A2(P3_EBX_REG_23__SCAN_IN), 
        .A3(P3_DATAWIDTH_REG_23__SCAN_IN), .A4(P1_UWORD_REG_6__SCAN_IN), .ZN(
        n15194) );
  OR4_X1 U18729 ( .A1(n15197), .A2(n15196), .A3(n15195), .A4(n15194), .ZN(
        n15201) );
  NAND4_X1 U18730 ( .A1(P1_ADDRESS_REG_5__SCAN_IN), .A2(DATAI_14_), .A3(
        P3_REIP_REG_2__SCAN_IN), .A4(BUF2_REG_17__SCAN_IN), .ZN(n15200) );
  NAND4_X1 U18731 ( .A1(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_23__SCAN_IN), .A3(
        P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A4(P1_REIP_REG_24__SCAN_IN), .ZN(
        n15199) );
  NAND4_X1 U18732 ( .A1(BUF1_REG_8__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A3(P3_DATAO_REG_16__SCAN_IN), 
        .A4(P1_BE_N_REG_3__SCAN_IN), .ZN(n15198) );
  NOR4_X1 U18733 ( .A1(n15201), .A2(n15200), .A3(n15199), .A4(n15198), .ZN(
        n15227) );
  NAND4_X1 U18734 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(P1_REIP_REG_4__SCAN_IN), 
        .A3(P1_REIP_REG_12__SCAN_IN), .A4(n15283), .ZN(n15204) );
  NAND4_X1 U18735 ( .A1(P2_INSTQUEUE_REG_6__0__SCAN_IN), .A2(
        P2_EBX_REG_18__SCAN_IN), .A3(BUF1_REG_5__SCAN_IN), .A4(
        P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n15203) );
  NAND4_X1 U18736 ( .A1(P2_EBX_REG_28__SCAN_IN), .A2(
        P2_ADDRESS_REG_16__SCAN_IN), .A3(P2_DATAWIDTH_REG_8__SCAN_IN), .A4(
        P3_EBX_REG_31__SCAN_IN), .ZN(n15202) );
  NOR3_X1 U18737 ( .A1(n15204), .A2(n15203), .A3(n15202), .ZN(n15226) );
  NOR4_X1 U18738 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(
        P1_INSTQUEUE_REG_5__0__SCAN_IN), .A3(P2_DATAWIDTH_REG_2__SCAN_IN), 
        .A4(P2_DATAWIDTH_REG_11__SCAN_IN), .ZN(n15205) );
  NAND4_X1 U18739 ( .A1(n15206), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A3(
        P1_INSTQUEUE_REG_8__0__SCAN_IN), .A4(n15205), .ZN(n15210) );
  NOR4_X1 U18740 ( .A1(P2_EAX_REG_7__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_26__SCAN_IN), .A3(DATAI_20_), .A4(
        P2_UWORD_REG_3__SCAN_IN), .ZN(n15207) );
  NAND4_X1 U18741 ( .A1(n15208), .A2(n15207), .A3(n9947), .A4(n20333), .ZN(
        n15209) );
  NOR2_X1 U18742 ( .A1(n15210), .A2(n15209), .ZN(n15225) );
  NOR4_X1 U18743 ( .A1(P1_INSTQUEUE_REG_8__2__SCAN_IN), .A2(
        P1_INSTQUEUE_REG_14__2__SCAN_IN), .A3(P1_INSTQUEUE_REG_0__2__SCAN_IN), 
        .A4(n15336), .ZN(n15214) );
  INV_X1 U18744 ( .A(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n15381) );
  NOR4_X1 U18745 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(P1_EBX_REG_19__SCAN_IN), .A4(
        n15381), .ZN(n15213) );
  NOR4_X1 U18746 ( .A1(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(
        P1_INSTQUEUE_REG_12__7__SCAN_IN), .A3(P1_EBX_REG_31__SCAN_IN), .A4(
        n9954), .ZN(n15212) );
  INV_X1 U18747 ( .A(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n15347) );
  NOR4_X1 U18748 ( .A1(P1_INSTQUEUE_REG_13__5__SCAN_IN), .A2(
        P1_INSTQUEUE_REG_0__5__SCAN_IN), .A3(P1_INSTQUEUE_REG_4__7__SCAN_IN), 
        .A4(n15347), .ZN(n15211) );
  NAND4_X1 U18749 ( .A1(n15214), .A2(n15213), .A3(n15212), .A4(n15211), .ZN(
        n15223) );
  NOR4_X1 U18750 ( .A1(P3_UWORD_REG_5__SCAN_IN), .A2(P3_EAX_REG_13__SCAN_IN), 
        .A3(BUF2_REG_15__SCAN_IN), .A4(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n15218) );
  NOR4_X1 U18751 ( .A1(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A4(P3_DATAO_REG_1__SCAN_IN), .ZN(
        n15217) );
  NOR4_X1 U18752 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(
        P3_INSTQUEUE_REG_1__4__SCAN_IN), .A3(P3_INSTQUEUE_REG_8__4__SCAN_IN), 
        .A4(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n15216) );
  NOR4_X1 U18753 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(
        P3_INSTQUEUE_REG_11__1__SCAN_IN), .A3(P3_INSTQUEUE_REG_3__1__SCAN_IN), 
        .A4(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n15215) );
  NAND4_X1 U18754 ( .A1(n15218), .A2(n15217), .A3(n15216), .A4(n15215), .ZN(
        n15222) );
  NOR2_X1 U18755 ( .A1(P1_EAX_REG_2__SCAN_IN), .A2(
        P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n15220) );
  NOR4_X1 U18756 ( .A1(P2_ADDRESS_REG_17__SCAN_IN), .A2(
        P2_DATAO_REG_20__SCAN_IN), .A3(P3_ADDRESS_REG_22__SCAN_IN), .A4(
        P3_DATAO_REG_31__SCAN_IN), .ZN(n15219) );
  NAND4_X1 U18757 ( .A1(P1_EAX_REG_5__SCAN_IN), .A2(P1_EAX_REG_1__SCAN_IN), 
        .A3(n15220), .A4(n15219), .ZN(n15221) );
  NOR3_X1 U18758 ( .A1(n15223), .A2(n15222), .A3(n15221), .ZN(n15224) );
  NAND4_X1 U18759 ( .A1(n15227), .A2(n15226), .A3(n15225), .A4(n15224), .ZN(
        n15239) );
  NAND4_X1 U18760 ( .A1(BUF1_REG_1__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A3(P2_DATAO_REG_2__SCAN_IN), 
        .A4(P1_DATAWIDTH_REG_9__SCAN_IN), .ZN(n15228) );
  NOR3_X1 U18761 ( .A1(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(DATAI_31_), 
        .A3(n15228), .ZN(n15237) );
  NAND4_X1 U18762 ( .A1(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_2__7__SCAN_IN), .A3(P2_PHYADDRPOINTER_REG_0__SCAN_IN), 
        .A4(P2_REIP_REG_29__SCAN_IN), .ZN(n15235) );
  NAND4_X1 U18763 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(
        P3_INSTQUEUE_REG_5__1__SCAN_IN), .A3(P3_INSTQUEUE_REG_8__3__SCAN_IN), 
        .A4(P3_EAX_REG_12__SCAN_IN), .ZN(n15234) );
  NOR4_X1 U18764 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_14__3__SCAN_IN), .A3(P2_INSTQUEUE_REG_7__0__SCAN_IN), 
        .A4(P3_D_C_N_REG_SCAN_IN), .ZN(n15232) );
  NOR4_X1 U18765 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A3(P3_EBX_REG_25__SCAN_IN), .A4(
        P3_EBX_REG_27__SCAN_IN), .ZN(n15231) );
  NOR4_X1 U18766 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A3(P1_EAX_REG_30__SCAN_IN), .A4(
        DATAI_17_), .ZN(n15230) );
  NOR4_X1 U18767 ( .A1(P2_EBX_REG_1__SCAN_IN), .A2(P2_REIP_REG_30__SCAN_IN), 
        .A3(BUF2_REG_30__SCAN_IN), .A4(BUF1_REG_28__SCAN_IN), .ZN(n15229) );
  NAND4_X1 U18768 ( .A1(n15232), .A2(n15231), .A3(n15230), .A4(n15229), .ZN(
        n15233) );
  NOR3_X1 U18769 ( .A1(n15235), .A2(n15234), .A3(n15233), .ZN(n15236) );
  NAND4_X1 U18770 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(
        P1_DATAO_REG_27__SCAN_IN), .A3(n15237), .A4(n15236), .ZN(n15238) );
  NOR2_X1 U18771 ( .A1(n15239), .A2(n15238), .ZN(n15425) );
  INV_X1 U18772 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n18671) );
  INV_X1 U18773 ( .A(P1_ADDRESS_REG_8__SCAN_IN), .ZN(n21212) );
  AOI22_X1 U18774 ( .A1(n18671), .A2(keyinput43), .B1(n21212), .B2(keyinput21), 
        .ZN(n15240) );
  OAI221_X1 U18775 ( .B1(n18671), .B2(keyinput43), .C1(n21212), .C2(keyinput21), .A(n15240), .ZN(n15248) );
  INV_X1 U18776 ( .A(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n17799) );
  AOI22_X1 U18777 ( .A1(n17799), .A2(keyinput98), .B1(n10748), .B2(keyinput12), 
        .ZN(n15241) );
  OAI221_X1 U18778 ( .B1(n17799), .B2(keyinput98), .C1(n10748), .C2(keyinput12), .A(n15241), .ZN(n15247) );
  INV_X1 U18779 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n19622) );
  AOI22_X1 U18780 ( .A1(n17976), .A2(keyinput99), .B1(n19622), .B2(keyinput16), 
        .ZN(n15242) );
  OAI221_X1 U18781 ( .B1(n17976), .B2(keyinput99), .C1(n19622), .C2(keyinput16), .A(n15242), .ZN(n15246) );
  INV_X1 U18782 ( .A(P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n15244) );
  AOI22_X1 U18783 ( .A1(n11022), .A2(keyinput41), .B1(n15244), .B2(keyinput105), .ZN(n15243) );
  OAI221_X1 U18784 ( .B1(n11022), .B2(keyinput41), .C1(n15244), .C2(
        keyinput105), .A(n15243), .ZN(n15245) );
  NOR4_X1 U18785 ( .A1(n15248), .A2(n15247), .A3(n15246), .A4(n15245), .ZN(
        n15260) );
  XOR2_X1 U18786 ( .A(keyinput87), .B(n18459), .Z(n15259) );
  XOR2_X1 U18787 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B(keyinput92), .Z(
        n15257) );
  XNOR2_X1 U18788 ( .A(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B(keyinput46), .ZN(
        n15252) );
  XNOR2_X1 U18789 ( .A(P2_REIP_REG_29__SCAN_IN), .B(keyinput101), .ZN(n15251)
         );
  XNOR2_X1 U18790 ( .A(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B(keyinput93), .ZN(
        n15250) );
  XNOR2_X1 U18791 ( .A(keyinput97), .B(BUF1_REG_5__SCAN_IN), .ZN(n15249) );
  NAND4_X1 U18792 ( .A1(n15252), .A2(n15251), .A3(n15250), .A4(n15249), .ZN(
        n15256) );
  XNOR2_X1 U18793 ( .A(n10291), .B(keyinput120), .ZN(n15255) );
  INV_X1 U18794 ( .A(DATAI_17_), .ZN(n15253) );
  XNOR2_X1 U18795 ( .A(keyinput35), .B(n15253), .ZN(n15254) );
  NOR4_X1 U18796 ( .A1(n15257), .A2(n15256), .A3(n15255), .A4(n15254), .ZN(
        n15258) );
  AND3_X1 U18797 ( .A1(n15260), .A2(n15259), .A3(n15258), .ZN(n15293) );
  INV_X1 U18798 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n20103) );
  INV_X1 U18799 ( .A(BUF2_REG_22__SCAN_IN), .ZN(n19059) );
  AOI22_X1 U18800 ( .A1(n20103), .A2(keyinput24), .B1(keyinput61), .B2(n19059), 
        .ZN(n15261) );
  OAI221_X1 U18801 ( .B1(n20103), .B2(keyinput24), .C1(n19059), .C2(keyinput61), .A(n15261), .ZN(n15271) );
  INV_X1 U18802 ( .A(DATAI_31_), .ZN(n15263) );
  AOI22_X1 U18803 ( .A1(n15263), .A2(keyinput26), .B1(keyinput78), .B2(n17325), 
        .ZN(n15262) );
  OAI221_X1 U18804 ( .B1(n15263), .B2(keyinput26), .C1(n17325), .C2(keyinput78), .A(n15262), .ZN(n15270) );
  INV_X1 U18805 ( .A(P3_D_C_N_REG_SCAN_IN), .ZN(n15265) );
  AOI22_X1 U18806 ( .A1(n16159), .A2(keyinput116), .B1(keyinput67), .B2(n15265), .ZN(n15264) );
  OAI221_X1 U18807 ( .B1(n16159), .B2(keyinput116), .C1(n15265), .C2(
        keyinput67), .A(n15264), .ZN(n15269) );
  INV_X1 U18808 ( .A(P3_EBX_REG_16__SCAN_IN), .ZN(n17627) );
  INV_X1 U18809 ( .A(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n15267) );
  AOI22_X1 U18810 ( .A1(n17627), .A2(keyinput47), .B1(n15267), .B2(keyinput110), .ZN(n15266) );
  OAI221_X1 U18811 ( .B1(n17627), .B2(keyinput47), .C1(n15267), .C2(
        keyinput110), .A(n15266), .ZN(n15268) );
  NOR4_X1 U18812 ( .A1(n15271), .A2(n15270), .A3(n15269), .A4(n15268), .ZN(
        n15292) );
  INV_X1 U18813 ( .A(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n17933) );
  AOI22_X1 U18814 ( .A1(n17933), .A2(keyinput96), .B1(n20891), .B2(keyinput108), .ZN(n15272) );
  OAI221_X1 U18815 ( .B1(n17933), .B2(keyinput96), .C1(n20891), .C2(
        keyinput108), .A(n15272), .ZN(n15279) );
  AOI22_X1 U18816 ( .A1(n17720), .A2(keyinput48), .B1(n9947), .B2(keyinput127), 
        .ZN(n15273) );
  OAI221_X1 U18817 ( .B1(n17720), .B2(keyinput48), .C1(n9947), .C2(keyinput127), .A(n15273), .ZN(n15278) );
  INV_X1 U18818 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n21257) );
  INV_X1 U18819 ( .A(P3_UWORD_REG_5__SCAN_IN), .ZN(n18224) );
  AOI22_X1 U18820 ( .A1(n21257), .A2(keyinput118), .B1(keyinput109), .B2(
        n18224), .ZN(n15274) );
  OAI221_X1 U18821 ( .B1(n21257), .B2(keyinput118), .C1(n18224), .C2(
        keyinput109), .A(n15274), .ZN(n15277) );
  INV_X1 U18822 ( .A(P2_DATAWIDTH_REG_11__SCAN_IN), .ZN(n20617) );
  AOI22_X1 U18823 ( .A1(n17811), .A2(keyinput77), .B1(n20617), .B2(keyinput27), 
        .ZN(n15275) );
  OAI221_X1 U18824 ( .B1(n17811), .B2(keyinput77), .C1(n20617), .C2(keyinput27), .A(n15275), .ZN(n15276) );
  NOR4_X1 U18825 ( .A1(n15279), .A2(n15278), .A3(n15277), .A4(n15276), .ZN(
        n15291) );
  INV_X1 U18826 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n20865) );
  INV_X1 U18827 ( .A(BUF1_REG_1__SCAN_IN), .ZN(n17219) );
  AOI22_X1 U18828 ( .A1(n20865), .A2(keyinput51), .B1(keyinput20), .B2(n17219), 
        .ZN(n15280) );
  OAI221_X1 U18829 ( .B1(n20865), .B2(keyinput51), .C1(n17219), .C2(keyinput20), .A(n15280), .ZN(n15289) );
  AOI22_X1 U18830 ( .A1(n17631), .A2(keyinput79), .B1(keyinput5), .B2(n17207), 
        .ZN(n15281) );
  OAI221_X1 U18831 ( .B1(n17631), .B2(keyinput79), .C1(n17207), .C2(keyinput5), 
        .A(n15281), .ZN(n15288) );
  AOI22_X1 U18832 ( .A1(n15283), .A2(keyinput49), .B1(keyinput19), .B2(n20900), 
        .ZN(n15282) );
  OAI221_X1 U18833 ( .B1(n15283), .B2(keyinput49), .C1(n20900), .C2(keyinput19), .A(n15282), .ZN(n15287) );
  AOI22_X1 U18834 ( .A1(n14761), .A2(keyinput44), .B1(keyinput28), .B2(n15285), 
        .ZN(n15284) );
  OAI221_X1 U18835 ( .B1(n14761), .B2(keyinput44), .C1(n15285), .C2(keyinput28), .A(n15284), .ZN(n15286) );
  NOR4_X1 U18836 ( .A1(n15289), .A2(n15288), .A3(n15287), .A4(n15286), .ZN(
        n15290) );
  AND4_X1 U18837 ( .A1(n15293), .A2(n15292), .A3(n15291), .A4(n15290), .ZN(
        n15331) );
  INV_X1 U18838 ( .A(BUF2_REG_15__SCAN_IN), .ZN(n17236) );
  AOI22_X1 U18839 ( .A1(n17737), .A2(keyinput113), .B1(n17236), .B2(keyinput91), .ZN(n15294) );
  OAI221_X1 U18840 ( .B1(n17737), .B2(keyinput113), .C1(n17236), .C2(
        keyinput91), .A(n15294), .ZN(n15302) );
  INV_X1 U18841 ( .A(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n15296) );
  AOI22_X1 U18842 ( .A1(n15296), .A2(keyinput31), .B1(n10085), .B2(keyinput75), 
        .ZN(n15295) );
  OAI221_X1 U18843 ( .B1(n15296), .B2(keyinput31), .C1(n10085), .C2(keyinput75), .A(n15295), .ZN(n15301) );
  INV_X1 U18844 ( .A(P1_DATAWIDTH_REG_26__SCAN_IN), .ZN(n21177) );
  INV_X1 U18845 ( .A(P1_DATAWIDTH_REG_9__SCAN_IN), .ZN(n21178) );
  AOI22_X1 U18846 ( .A1(n21177), .A2(keyinput73), .B1(keyinput36), .B2(n21178), 
        .ZN(n15297) );
  OAI221_X1 U18847 ( .B1(n21177), .B2(keyinput73), .C1(n21178), .C2(keyinput36), .A(n15297), .ZN(n15300) );
  INV_X1 U18848 ( .A(P3_DATAO_REG_1__SCAN_IN), .ZN(n18265) );
  AOI22_X1 U18849 ( .A1(n18265), .A2(keyinput53), .B1(keyinput74), .B2(n18337), 
        .ZN(n15298) );
  OAI221_X1 U18850 ( .B1(n18265), .B2(keyinput53), .C1(n18337), .C2(keyinput74), .A(n15298), .ZN(n15299) );
  NOR4_X1 U18851 ( .A1(n15302), .A2(n15301), .A3(n15300), .A4(n15299), .ZN(
        n15330) );
  INV_X1 U18852 ( .A(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n15305) );
  INV_X1 U18853 ( .A(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n15304) );
  AOI22_X1 U18854 ( .A1(n15305), .A2(keyinput11), .B1(n15304), .B2(keyinput119), .ZN(n15303) );
  OAI221_X1 U18855 ( .B1(n15305), .B2(keyinput11), .C1(n15304), .C2(
        keyinput119), .A(n15303), .ZN(n15315) );
  AOI22_X1 U18856 ( .A1(n15307), .A2(keyinput95), .B1(n15126), .B2(keyinput111), .ZN(n15306) );
  OAI221_X1 U18857 ( .B1(n15307), .B2(keyinput95), .C1(n15126), .C2(
        keyinput111), .A(n15306), .ZN(n15314) );
  INV_X1 U18858 ( .A(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n15310) );
  INV_X1 U18859 ( .A(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n15309) );
  AOI22_X1 U18860 ( .A1(n15310), .A2(keyinput125), .B1(n15309), .B2(
        keyinput122), .ZN(n15308) );
  OAI221_X1 U18861 ( .B1(n15310), .B2(keyinput125), .C1(n15309), .C2(
        keyinput122), .A(n15308), .ZN(n15313) );
  INV_X1 U18862 ( .A(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n17788) );
  AOI22_X1 U18863 ( .A1(n17240), .A2(keyinput71), .B1(keyinput65), .B2(n17788), 
        .ZN(n15311) );
  OAI221_X1 U18864 ( .B1(n17240), .B2(keyinput71), .C1(n17788), .C2(keyinput65), .A(n15311), .ZN(n15312) );
  NOR4_X1 U18865 ( .A1(n15315), .A2(n15314), .A3(n15313), .A4(n15312), .ZN(
        n15329) );
  INV_X1 U18866 ( .A(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n15318) );
  AOI22_X1 U18867 ( .A1(n15318), .A2(keyinput102), .B1(n15317), .B2(
        keyinput100), .ZN(n15316) );
  OAI221_X1 U18868 ( .B1(n15318), .B2(keyinput102), .C1(n15317), .C2(
        keyinput100), .A(n15316), .ZN(n15327) );
  INV_X1 U18869 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n17243) );
  INV_X1 U18870 ( .A(P3_DATAO_REG_16__SCAN_IN), .ZN(n18235) );
  AOI22_X1 U18871 ( .A1(n17243), .A2(keyinput40), .B1(keyinput94), .B2(n18235), 
        .ZN(n15319) );
  OAI221_X1 U18872 ( .B1(n17243), .B2(keyinput40), .C1(n18235), .C2(keyinput94), .A(n15319), .ZN(n15326) );
  AOI22_X1 U18873 ( .A1(n21256), .A2(keyinput59), .B1(keyinput66), .B2(n15321), 
        .ZN(n15320) );
  OAI221_X1 U18874 ( .B1(n21256), .B2(keyinput59), .C1(n15321), .C2(keyinput66), .A(n15320), .ZN(n15325) );
  AOI22_X1 U18875 ( .A1(n19666), .A2(keyinput52), .B1(n15323), .B2(keyinput123), .ZN(n15322) );
  OAI221_X1 U18876 ( .B1(n19666), .B2(keyinput52), .C1(n15323), .C2(
        keyinput123), .A(n15322), .ZN(n15324) );
  NOR4_X1 U18877 ( .A1(n15327), .A2(n15326), .A3(n15325), .A4(n15324), .ZN(
        n15328) );
  NAND4_X1 U18878 ( .A1(n15331), .A2(n15330), .A3(n15329), .A4(n15328), .ZN(
        n15423) );
  AOI22_X1 U18879 ( .A1(n17887), .A2(keyinput0), .B1(keyinput7), .B2(n19170), 
        .ZN(n15332) );
  OAI221_X1 U18880 ( .B1(n17887), .B2(keyinput0), .C1(n19170), .C2(keyinput7), 
        .A(n15332), .ZN(n15340) );
  AOI22_X1 U18881 ( .A1(n20007), .A2(keyinput13), .B1(keyinput68), .B2(n17930), 
        .ZN(n15333) );
  OAI221_X1 U18882 ( .B1(n20007), .B2(keyinput13), .C1(n17930), .C2(keyinput68), .A(n15333), .ZN(n15339) );
  INV_X1 U18883 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n18242) );
  AOI22_X1 U18884 ( .A1(n18242), .A2(keyinput1), .B1(n16785), .B2(keyinput23), 
        .ZN(n15334) );
  OAI221_X1 U18885 ( .B1(n18242), .B2(keyinput1), .C1(n16785), .C2(keyinput23), 
        .A(n15334), .ZN(n15338) );
  INV_X1 U18886 ( .A(P1_EBX_REG_19__SCAN_IN), .ZN(n16643) );
  AOI22_X1 U18887 ( .A1(n15336), .A2(keyinput58), .B1(n16643), .B2(keyinput18), 
        .ZN(n15335) );
  OAI221_X1 U18888 ( .B1(n15336), .B2(keyinput58), .C1(n16643), .C2(keyinput18), .A(n15335), .ZN(n15337) );
  NOR4_X1 U18889 ( .A1(n15340), .A2(n15339), .A3(n15338), .A4(n15337), .ZN(
        n15377) );
  INV_X1 U18890 ( .A(READY22_REG_SCAN_IN), .ZN(n15342) );
  AOI22_X1 U18891 ( .A1(n15342), .A2(keyinput89), .B1(keyinput9), .B2(n18021), 
        .ZN(n15341) );
  OAI221_X1 U18892 ( .B1(n15342), .B2(keyinput89), .C1(n18021), .C2(keyinput9), 
        .A(n15341), .ZN(n15354) );
  AOI22_X1 U18893 ( .A1(n15344), .A2(keyinput4), .B1(n20749), .B2(keyinput15), 
        .ZN(n15343) );
  OAI221_X1 U18894 ( .B1(n15344), .B2(keyinput4), .C1(n20749), .C2(keyinput15), 
        .A(n15343), .ZN(n15353) );
  AOI22_X1 U18895 ( .A1(n15347), .A2(keyinput106), .B1(keyinput69), .B2(n15346), .ZN(n15345) );
  OAI221_X1 U18896 ( .B1(n15347), .B2(keyinput106), .C1(n15346), .C2(
        keyinput69), .A(n15345), .ZN(n15352) );
  INV_X1 U18897 ( .A(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n15350) );
  INV_X1 U18898 ( .A(P3_UWORD_REG_6__SCAN_IN), .ZN(n15349) );
  AOI22_X1 U18899 ( .A1(n15350), .A2(keyinput10), .B1(keyinput55), .B2(n15349), 
        .ZN(n15348) );
  OAI221_X1 U18900 ( .B1(n15350), .B2(keyinput10), .C1(n15349), .C2(keyinput55), .A(n15348), .ZN(n15351) );
  NOR4_X1 U18901 ( .A1(n15354), .A2(n15353), .A3(n15352), .A4(n15351), .ZN(
        n15376) );
  INV_X1 U18902 ( .A(BUF2_REG_17__SCAN_IN), .ZN(n17239) );
  AOI22_X1 U18903 ( .A1(n17239), .A2(keyinput107), .B1(n17969), .B2(keyinput34), .ZN(n15355) );
  OAI221_X1 U18904 ( .B1(n17239), .B2(keyinput107), .C1(n17969), .C2(
        keyinput34), .A(n15355), .ZN(n15363) );
  INV_X1 U18905 ( .A(P1_ADDRESS_REG_5__SCAN_IN), .ZN(n21207) );
  INV_X1 U18906 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n20657) );
  AOI22_X1 U18907 ( .A1(n21207), .A2(keyinput114), .B1(n20657), .B2(keyinput6), 
        .ZN(n15356) );
  OAI221_X1 U18908 ( .B1(n21207), .B2(keyinput114), .C1(n20657), .C2(keyinput6), .A(n15356), .ZN(n15362) );
  INV_X1 U18909 ( .A(P2_EBX_REG_28__SCAN_IN), .ZN(n15358) );
  INV_X1 U18910 ( .A(P2_DATAWIDTH_REG_8__SCAN_IN), .ZN(n20618) );
  AOI22_X1 U18911 ( .A1(n15358), .A2(keyinput115), .B1(keyinput88), .B2(n20618), .ZN(n15357) );
  OAI221_X1 U18912 ( .B1(n15358), .B2(keyinput115), .C1(n20618), .C2(
        keyinput88), .A(n15357), .ZN(n15361) );
  INV_X1 U18913 ( .A(P1_REIP_REG_19__SCAN_IN), .ZN(n21229) );
  AOI22_X1 U18914 ( .A1(n21229), .A2(keyinput83), .B1(n15657), .B2(keyinput63), 
        .ZN(n15359) );
  OAI221_X1 U18915 ( .B1(n21229), .B2(keyinput83), .C1(n15657), .C2(keyinput63), .A(n15359), .ZN(n15360) );
  NOR4_X1 U18916 ( .A1(n15363), .A2(n15362), .A3(n15361), .A4(n15360), .ZN(
        n15375) );
  INV_X1 U18917 ( .A(P3_DATAWIDTH_REG_23__SCAN_IN), .ZN(n19561) );
  AOI22_X1 U18918 ( .A1(n17736), .A2(keyinput8), .B1(keyinput60), .B2(n19561), 
        .ZN(n15364) );
  OAI221_X1 U18919 ( .B1(n17736), .B2(keyinput8), .C1(n19561), .C2(keyinput60), 
        .A(n15364), .ZN(n15373) );
  INV_X1 U18920 ( .A(P2_DATAWIDTH_REG_2__SCAN_IN), .ZN(n20620) );
  AOI22_X1 U18921 ( .A1(n15366), .A2(keyinput25), .B1(keyinput33), .B2(n20620), 
        .ZN(n15365) );
  OAI221_X1 U18922 ( .B1(n15366), .B2(keyinput25), .C1(n20620), .C2(keyinput33), .A(n15365), .ZN(n15372) );
  INV_X1 U18923 ( .A(P1_UWORD_REG_6__SCAN_IN), .ZN(n20868) );
  AOI22_X1 U18924 ( .A1(n20333), .A2(keyinput39), .B1(keyinput54), .B2(n20868), 
        .ZN(n15367) );
  OAI221_X1 U18925 ( .B1(n20333), .B2(keyinput39), .C1(n20868), .C2(keyinput54), .A(n15367), .ZN(n15371) );
  INV_X1 U18926 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n19580) );
  INV_X1 U18927 ( .A(DATAI_14_), .ZN(n15369) );
  AOI22_X1 U18928 ( .A1(n19580), .A2(keyinput30), .B1(n15369), .B2(keyinput76), 
        .ZN(n15368) );
  OAI221_X1 U18929 ( .B1(n19580), .B2(keyinput30), .C1(n15369), .C2(keyinput76), .A(n15368), .ZN(n15370) );
  NOR4_X1 U18930 ( .A1(n15373), .A2(n15372), .A3(n15371), .A4(n15370), .ZN(
        n15374) );
  NAND4_X1 U18931 ( .A1(n15377), .A2(n15376), .A3(n15375), .A4(n15374), .ZN(
        n15422) );
  INV_X1 U18932 ( .A(DATAI_20_), .ZN(n15379) );
  INV_X1 U18933 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n18808) );
  AOI22_X1 U18934 ( .A1(n15379), .A2(keyinput62), .B1(keyinput72), .B2(n18808), 
        .ZN(n15378) );
  OAI221_X1 U18935 ( .B1(n15379), .B2(keyinput62), .C1(n18808), .C2(keyinput72), .A(n15378), .ZN(n15387) );
  AOI22_X1 U18936 ( .A1(n9954), .A2(keyinput3), .B1(keyinput112), .B2(n15381), 
        .ZN(n15380) );
  OAI221_X1 U18937 ( .B1(n9954), .B2(keyinput3), .C1(n15381), .C2(keyinput112), 
        .A(n15380), .ZN(n15386) );
  AOI22_X1 U18938 ( .A1(n11802), .A2(keyinput90), .B1(keyinput126), .B2(n10557), .ZN(n15382) );
  OAI221_X1 U18939 ( .B1(n11802), .B2(keyinput90), .C1(n10557), .C2(
        keyinput126), .A(n15382), .ZN(n15385) );
  INV_X1 U18940 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n20019) );
  INV_X1 U18941 ( .A(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n17478) );
  AOI22_X1 U18942 ( .A1(n20019), .A2(keyinput85), .B1(n17478), .B2(keyinput104), .ZN(n15383) );
  OAI221_X1 U18943 ( .B1(n20019), .B2(keyinput85), .C1(n17478), .C2(
        keyinput104), .A(n15383), .ZN(n15384) );
  NOR4_X1 U18944 ( .A1(n15387), .A2(n15386), .A3(n15385), .A4(n15384), .ZN(
        n15420) );
  INV_X1 U18945 ( .A(BUF2_REG_30__SCAN_IN), .ZN(n20114) );
  AOI22_X1 U18946 ( .A1(n21217), .A2(keyinput84), .B1(n20114), .B2(keyinput14), 
        .ZN(n15388) );
  OAI221_X1 U18947 ( .B1(n21217), .B2(keyinput84), .C1(n20114), .C2(keyinput14), .A(n15388), .ZN(n15397) );
  INV_X1 U18948 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n20659) );
  INV_X1 U18949 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n21239) );
  AOI22_X1 U18950 ( .A1(n20659), .A2(keyinput80), .B1(keyinput56), .B2(n21239), 
        .ZN(n15389) );
  OAI221_X1 U18951 ( .B1(n20659), .B2(keyinput80), .C1(n21239), .C2(keyinput56), .A(n15389), .ZN(n15396) );
  INV_X1 U18952 ( .A(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n17999) );
  AOI22_X1 U18953 ( .A1(n17999), .A2(keyinput64), .B1(n15391), .B2(keyinput50), 
        .ZN(n15390) );
  OAI221_X1 U18954 ( .B1(n17999), .B2(keyinput64), .C1(n15391), .C2(keyinput50), .A(n15390), .ZN(n15395) );
  INV_X1 U18955 ( .A(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n15393) );
  AOI22_X1 U18956 ( .A1(n15393), .A2(keyinput32), .B1(n10660), .B2(keyinput38), 
        .ZN(n15392) );
  OAI221_X1 U18957 ( .B1(n15393), .B2(keyinput32), .C1(n10660), .C2(keyinput38), .A(n15392), .ZN(n15394) );
  NOR4_X1 U18958 ( .A1(n15397), .A2(n15396), .A3(n15395), .A4(n15394), .ZN(
        n15419) );
  INV_X1 U18959 ( .A(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n15399) );
  AOI22_X1 U18960 ( .A1(n15399), .A2(keyinput103), .B1(keyinput37), .B2(n17923), .ZN(n15398) );
  OAI221_X1 U18961 ( .B1(n15399), .B2(keyinput103), .C1(n17923), .C2(
        keyinput37), .A(n15398), .ZN(n15406) );
  INV_X1 U18962 ( .A(P1_ADDRESS_REG_24__SCAN_IN), .ZN(n21240) );
  AOI22_X1 U18963 ( .A1(n21240), .A2(keyinput82), .B1(n20898), .B2(keyinput117), .ZN(n15400) );
  OAI221_X1 U18964 ( .B1(n21240), .B2(keyinput82), .C1(n20898), .C2(
        keyinput117), .A(n15400), .ZN(n15405) );
  INV_X1 U18965 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n20651) );
  INV_X1 U18966 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n18240) );
  AOI22_X1 U18967 ( .A1(n20651), .A2(keyinput45), .B1(keyinput121), .B2(n18240), .ZN(n15401) );
  OAI221_X1 U18968 ( .B1(n20651), .B2(keyinput45), .C1(n18240), .C2(
        keyinput121), .A(n15401), .ZN(n15404) );
  INV_X1 U18969 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n20639) );
  INV_X1 U18970 ( .A(P2_LWORD_REG_7__SCAN_IN), .ZN(n20008) );
  AOI22_X1 U18971 ( .A1(n20639), .A2(keyinput81), .B1(keyinput57), .B2(n20008), 
        .ZN(n15402) );
  OAI221_X1 U18972 ( .B1(n20639), .B2(keyinput81), .C1(n20008), .C2(keyinput57), .A(n15402), .ZN(n15403) );
  NOR4_X1 U18973 ( .A1(n15406), .A2(n15405), .A3(n15404), .A4(n15403), .ZN(
        n15418) );
  AOI22_X1 U18974 ( .A1(n15466), .A2(keyinput124), .B1(n10829), .B2(keyinput42), .ZN(n15407) );
  OAI221_X1 U18975 ( .B1(n15466), .B2(keyinput124), .C1(n10829), .C2(
        keyinput42), .A(n15407), .ZN(n15416) );
  INV_X1 U18976 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n18206) );
  AOI22_X1 U18977 ( .A1(n18206), .A2(keyinput17), .B1(n21202), .B2(keyinput22), 
        .ZN(n15408) );
  OAI221_X1 U18978 ( .B1(n18206), .B2(keyinput17), .C1(n21202), .C2(keyinput22), .A(n15408), .ZN(n15415) );
  INV_X1 U18979 ( .A(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n15411) );
  INV_X1 U18980 ( .A(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n15410) );
  AOI22_X1 U18981 ( .A1(n15411), .A2(keyinput86), .B1(n15410), .B2(keyinput29), 
        .ZN(n15409) );
  OAI221_X1 U18982 ( .B1(n15411), .B2(keyinput86), .C1(n15410), .C2(keyinput29), .A(n15409), .ZN(n15414) );
  INV_X1 U18983 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n20665) );
  AOI22_X1 U18984 ( .A1(n17918), .A2(keyinput70), .B1(n20665), .B2(keyinput2), 
        .ZN(n15412) );
  OAI221_X1 U18985 ( .B1(n17918), .B2(keyinput70), .C1(n20665), .C2(keyinput2), 
        .A(n15412), .ZN(n15413) );
  NOR4_X1 U18986 ( .A1(n15416), .A2(n15415), .A3(n15414), .A4(n15413), .ZN(
        n15417) );
  NAND4_X1 U18987 ( .A1(n15420), .A2(n15419), .A3(n15418), .A4(n15417), .ZN(
        n15421) );
  NOR3_X1 U18988 ( .A1(n15423), .A2(n15422), .A3(n15421), .ZN(n15424) );
  XOR2_X1 U18989 ( .A(n15425), .B(n15424), .Z(n15426) );
  XNOR2_X1 U18990 ( .A(n15427), .B(n15426), .ZN(P1_U2814) );
  INV_X1 U18991 ( .A(n15518), .ZN(n15429) );
  AOI21_X1 U18992 ( .B1(n15430), .B2(n15520), .A(n15429), .ZN(n16683) );
  INV_X1 U18993 ( .A(n16683), .ZN(n15594) );
  NAND2_X1 U18994 ( .A1(n15431), .A2(n15432), .ZN(n15433) );
  AND2_X1 U18995 ( .A1(n15522), .A2(n15433), .ZN(n15751) );
  AOI22_X1 U18996 ( .A1(n20850), .A2(P1_EBX_REG_17__SCAN_IN), .B1(n16629), 
        .B2(n16682), .ZN(n15434) );
  OAI211_X1 U18997 ( .C1(n20818), .C2(n15435), .A(n15434), .B(n20816), .ZN(
        n15438) );
  AOI21_X1 U18998 ( .B1(n21227), .B2(n15436), .A(n16574), .ZN(n15437) );
  AOI211_X1 U18999 ( .C1(n15751), .C2(n16609), .A(n15438), .B(n15437), .ZN(
        n15439) );
  OAI21_X1 U19000 ( .B1(n15594), .B2(n16617), .A(n15439), .ZN(P1_U2823) );
  AOI21_X1 U19001 ( .B1(n15440), .B2(n14663), .A(n9772), .ZN(n15673) );
  INV_X1 U19002 ( .A(n15673), .ZN(n15611) );
  NOR2_X1 U19003 ( .A1(n15441), .A2(n16632), .ZN(n16627) );
  NAND2_X1 U19004 ( .A1(P1_REIP_REG_13__SCAN_IN), .A2(n16627), .ZN(n16605) );
  NAND2_X1 U19005 ( .A1(n21222), .A2(n16605), .ZN(n15452) );
  OR2_X1 U19006 ( .A1(n20813), .A2(n15442), .ZN(n15443) );
  NAND2_X1 U19007 ( .A1(n15443), .A2(n20845), .ZN(n16613) );
  NAND2_X1 U19008 ( .A1(n15445), .A2(n15444), .ZN(n15446) );
  NAND2_X1 U19009 ( .A1(n15538), .A2(n15446), .ZN(n15768) );
  INV_X1 U19010 ( .A(n15671), .ZN(n15449) );
  NAND2_X1 U19011 ( .A1(n20849), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n15447) );
  OAI211_X1 U19012 ( .C1(n16622), .C2(n15542), .A(n15447), .B(n20816), .ZN(
        n15448) );
  AOI21_X1 U19013 ( .B1(n15449), .B2(n16629), .A(n15448), .ZN(n15450) );
  OAI21_X1 U19014 ( .B1(n15768), .B2(n20860), .A(n15450), .ZN(n15451) );
  AOI21_X1 U19015 ( .B1(n15452), .B2(n16613), .A(n15451), .ZN(n15453) );
  OAI21_X1 U19016 ( .B1(n15611), .B2(n16617), .A(n15453), .ZN(P1_U2826) );
  INV_X1 U19017 ( .A(n15454), .ZN(n15455) );
  NAND2_X1 U19018 ( .A1(n15455), .A2(n20855), .ZN(n15465) );
  INV_X1 U19019 ( .A(n20924), .ZN(n15456) );
  NAND2_X1 U19020 ( .A1(n16609), .A2(n15456), .ZN(n15458) );
  OAI21_X1 U19021 ( .B1(n20849), .B2(n16629), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n15457) );
  OAI211_X1 U19022 ( .C1(n15459), .C2(n16622), .A(n15458), .B(n15457), .ZN(
        n15460) );
  INV_X1 U19023 ( .A(n15460), .ZN(n15464) );
  INV_X1 U19024 ( .A(n20853), .ZN(n20837) );
  NAND2_X1 U19025 ( .A1(n20837), .A2(n12172), .ZN(n15463) );
  NAND2_X1 U19026 ( .A1(n15461), .A2(P1_REIP_REG_0__SCAN_IN), .ZN(n15462) );
  NAND4_X1 U19027 ( .A1(n15465), .A2(n15464), .A3(n15463), .A4(n15462), .ZN(
        P1_U2840) );
  OAI22_X1 U19028 ( .A1(n15467), .A2(n15543), .B1(n16644), .B2(n15466), .ZN(
        P1_U2841) );
  INV_X1 U19029 ( .A(n15468), .ZN(n15553) );
  INV_X1 U19030 ( .A(n15469), .ZN(n15470) );
  OAI222_X1 U19031 ( .A1(n16640), .A2(n15553), .B1(n15471), .B2(n16644), .C1(
        n15470), .C2(n15543), .ZN(P1_U2843) );
  INV_X1 U19032 ( .A(n15472), .ZN(n15557) );
  OAI222_X1 U19033 ( .A1(n16640), .A2(n15557), .B1(n15474), .B2(n16644), .C1(
        n15473), .C2(n15543), .ZN(P1_U2845) );
  INV_X1 U19034 ( .A(n15621), .ZN(n15560) );
  INV_X1 U19035 ( .A(n15475), .ZN(n15704) );
  AOI22_X1 U19036 ( .A1(n15704), .A2(n15528), .B1(P1_EBX_REG_26__SCAN_IN), 
        .B2(n15527), .ZN(n15476) );
  OAI21_X1 U19037 ( .B1(n15560), .B2(n16640), .A(n15476), .ZN(P1_U2846) );
  INV_X1 U19038 ( .A(n16650), .ZN(n15564) );
  OR2_X1 U19039 ( .A1(n15478), .A2(n15479), .ZN(n15480) );
  AND2_X1 U19040 ( .A1(n15481), .A2(n15480), .ZN(n16745) );
  AOI22_X1 U19041 ( .A1(n16745), .A2(n15528), .B1(P1_EBX_REG_25__SCAN_IN), 
        .B2(n15527), .ZN(n15482) );
  OAI21_X1 U19042 ( .B1(n15564), .B2(n16640), .A(n15482), .ZN(P1_U2847) );
  OAI21_X1 U19043 ( .B1(n15483), .B2(n15484), .A(n9769), .ZN(n16537) );
  NOR2_X1 U19044 ( .A1(n15496), .A2(n15485), .ZN(n15486) );
  OR2_X1 U19045 ( .A1(n15478), .A2(n15486), .ZN(n16541) );
  OAI22_X1 U19046 ( .A1(n16541), .A2(n15543), .B1(n15487), .B2(n16644), .ZN(
        n15488) );
  INV_X1 U19047 ( .A(n15488), .ZN(n15489) );
  OAI21_X1 U19048 ( .B1(n16537), .B2(n16640), .A(n15489), .ZN(P1_U2848) );
  AND2_X1 U19049 ( .A1(n15490), .A2(n15491), .ZN(n15492) );
  NOR2_X1 U19050 ( .A1(n15483), .A2(n15492), .ZN(n16657) );
  INV_X1 U19051 ( .A(n16657), .ZN(n15570) );
  INV_X1 U19052 ( .A(P1_EBX_REG_23__SCAN_IN), .ZN(n15498) );
  INV_X1 U19053 ( .A(n15493), .ZN(n15495) );
  AOI21_X1 U19054 ( .B1(n15495), .B2(n15502), .A(n15494), .ZN(n15497) );
  OR2_X1 U19055 ( .A1(n15497), .A2(n15496), .ZN(n16753) );
  OAI222_X1 U19056 ( .A1(n16640), .A2(n15570), .B1(n15498), .B2(n16644), .C1(
        n16753), .C2(n15543), .ZN(P1_U2849) );
  NAND2_X1 U19057 ( .A1(n15499), .A2(n15500), .ZN(n15501) );
  AND2_X1 U19058 ( .A1(n15490), .A2(n15501), .ZN(n16550) );
  INV_X1 U19059 ( .A(n16550), .ZN(n15574) );
  XNOR2_X1 U19060 ( .A(n15493), .B(n15502), .ZN(n16761) );
  AOI22_X1 U19061 ( .A1(n16761), .A2(n15528), .B1(P1_EBX_REG_22__SCAN_IN), 
        .B2(n15527), .ZN(n15503) );
  OAI21_X1 U19062 ( .B1(n15574), .B2(n16640), .A(n15503), .ZN(P1_U2850) );
  NAND2_X1 U19063 ( .A1(n15514), .A2(n15504), .ZN(n15505) );
  NAND2_X1 U19064 ( .A1(n15493), .A2(n15505), .ZN(n16556) );
  INV_X1 U19065 ( .A(P1_EBX_REG_21__SCAN_IN), .ZN(n15509) );
  AND2_X1 U19066 ( .A1(n15428), .A2(n15506), .ZN(n15511) );
  OR2_X1 U19067 ( .A1(n15511), .A2(n15507), .ZN(n15508) );
  NAND2_X1 U19068 ( .A1(n15499), .A2(n15508), .ZN(n16665) );
  OAI222_X1 U19069 ( .A1(n15543), .A2(n16556), .B1(n15509), .B2(n16644), .C1(
        n16665), .C2(n16640), .ZN(P1_U2851) );
  NOR2_X1 U19070 ( .A1(n15520), .A2(n15510), .ZN(n15584) );
  INV_X1 U19071 ( .A(n15584), .ZN(n15513) );
  AOI21_X1 U19072 ( .B1(n15513), .B2(n15512), .A(n15511), .ZN(n15653) );
  INV_X1 U19073 ( .A(n15653), .ZN(n16567) );
  INV_X1 U19074 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n15516) );
  OAI21_X1 U19075 ( .B1(n16581), .B2(n15515), .A(n15514), .ZN(n16566) );
  OAI222_X1 U19076 ( .A1(n16567), .A2(n16640), .B1(n16644), .B2(n15516), .C1(
        n16566), .C2(n15543), .ZN(P1_U2852) );
  NOR2_X1 U19077 ( .A1(n15520), .A2(n15519), .ZN(n15582) );
  AND2_X1 U19078 ( .A1(n15522), .A2(n15521), .ZN(n15523) );
  OR2_X1 U19079 ( .A1(n15523), .A2(n16579), .ZN(n16597) );
  OAI22_X1 U19080 ( .A1(n16597), .A2(n15543), .B1(n15524), .B2(n16644), .ZN(
        n15525) );
  INV_X1 U19081 ( .A(n15525), .ZN(n15526) );
  OAI21_X1 U19082 ( .B1(n16591), .B2(n16640), .A(n15526), .ZN(P1_U2854) );
  AOI22_X1 U19083 ( .A1(n15751), .A2(n15528), .B1(P1_EBX_REG_17__SCAN_IN), 
        .B2(n15527), .ZN(n15529) );
  OAI21_X1 U19084 ( .B1(n15594), .B2(n16640), .A(n15529), .ZN(P1_U2855) );
  XOR2_X1 U19085 ( .A(n15530), .B(n10178), .Z(n16695) );
  INV_X1 U19086 ( .A(n16695), .ZN(n15601) );
  OR2_X1 U19087 ( .A1(n15540), .A2(n15531), .ZN(n15532) );
  NAND2_X1 U19088 ( .A1(n15431), .A2(n15532), .ZN(n16777) );
  OAI22_X1 U19089 ( .A1(n16777), .A2(n15543), .B1(n16600), .B2(n16644), .ZN(
        n15533) );
  INV_X1 U19090 ( .A(n15533), .ZN(n15534) );
  OAI21_X1 U19091 ( .B1(n15601), .B2(n16640), .A(n15534), .ZN(P1_U2856) );
  OR2_X1 U19092 ( .A1(n9772), .A2(n15535), .ZN(n15536) );
  NAND2_X1 U19093 ( .A1(n10178), .A2(n15536), .ZN(n16701) );
  INV_X1 U19094 ( .A(P1_EBX_REG_15__SCAN_IN), .ZN(n16611) );
  AND2_X1 U19095 ( .A1(n15538), .A2(n15537), .ZN(n15539) );
  NOR2_X1 U19096 ( .A1(n15540), .A2(n15539), .ZN(n16608) );
  INV_X1 U19097 ( .A(n16608), .ZN(n15541) );
  OAI222_X1 U19098 ( .A1(n16701), .A2(n16640), .B1(n16611), .B2(n16644), .C1(
        n15541), .C2(n15543), .ZN(P1_U2857) );
  OAI22_X1 U19099 ( .A1(n15768), .A2(n15543), .B1(n15542), .B2(n16644), .ZN(
        n15544) );
  AOI21_X1 U19100 ( .B1(n15673), .B2(n15545), .A(n15544), .ZN(n15546) );
  INV_X1 U19101 ( .A(n15546), .ZN(P1_U2858) );
  AOI22_X1 U19102 ( .A1(n15595), .A2(BUF1_REG_30__SCAN_IN), .B1(
        P1_EAX_REG_30__SCAN_IN), .B2(n15606), .ZN(n15548) );
  AOI22_X1 U19103 ( .A1(n15598), .A2(n15607), .B1(n15596), .B2(DATAI_30_), 
        .ZN(n15547) );
  OAI211_X1 U19104 ( .C1(n15549), .C2(n15610), .A(n15548), .B(n15547), .ZN(
        P1_U2874) );
  AOI22_X1 U19105 ( .A1(n15595), .A2(BUF1_REG_29__SCAN_IN), .B1(
        P1_EAX_REG_29__SCAN_IN), .B2(n15606), .ZN(n15552) );
  AOI22_X1 U19106 ( .A1(n15598), .A2(n15550), .B1(n15596), .B2(DATAI_29_), 
        .ZN(n15551) );
  OAI211_X1 U19107 ( .C1(n15553), .C2(n15610), .A(n15552), .B(n15551), .ZN(
        P1_U2875) );
  AOI22_X1 U19108 ( .A1(n15595), .A2(BUF1_REG_27__SCAN_IN), .B1(
        P1_EAX_REG_27__SCAN_IN), .B2(n15606), .ZN(n15556) );
  AOI22_X1 U19109 ( .A1(n15598), .A2(n15554), .B1(n15596), .B2(DATAI_27_), 
        .ZN(n15555) );
  OAI211_X1 U19110 ( .C1(n15557), .C2(n15610), .A(n15556), .B(n15555), .ZN(
        P1_U2877) );
  AOI22_X1 U19111 ( .A1(n15595), .A2(BUF1_REG_26__SCAN_IN), .B1(
        P1_EAX_REG_26__SCAN_IN), .B2(n15606), .ZN(n15559) );
  AOI22_X1 U19112 ( .A1(n15598), .A2(n20907), .B1(n15596), .B2(DATAI_26_), 
        .ZN(n15558) );
  OAI211_X1 U19113 ( .C1(n15560), .C2(n15610), .A(n15559), .B(n15558), .ZN(
        P1_U2878) );
  AOI22_X1 U19114 ( .A1(n15595), .A2(BUF1_REG_25__SCAN_IN), .B1(
        P1_EAX_REG_25__SCAN_IN), .B2(n15606), .ZN(n15563) );
  AOI22_X1 U19115 ( .A1(n15598), .A2(n15561), .B1(n15596), .B2(DATAI_25_), 
        .ZN(n15562) );
  OAI211_X1 U19116 ( .C1(n15564), .C2(n15610), .A(n15563), .B(n15562), .ZN(
        P1_U2879) );
  AOI22_X1 U19117 ( .A1(n15595), .A2(BUF1_REG_24__SCAN_IN), .B1(
        P1_EAX_REG_24__SCAN_IN), .B2(n15606), .ZN(n15566) );
  AOI22_X1 U19118 ( .A1(n15598), .A2(n20905), .B1(n15596), .B2(DATAI_24_), 
        .ZN(n15565) );
  OAI211_X1 U19119 ( .C1(n16537), .C2(n15610), .A(n15566), .B(n15565), .ZN(
        P1_U2880) );
  AOI22_X1 U19120 ( .A1(n15595), .A2(BUF1_REG_23__SCAN_IN), .B1(
        P1_EAX_REG_23__SCAN_IN), .B2(n15606), .ZN(n15569) );
  AOI22_X1 U19121 ( .A1(n15598), .A2(n15567), .B1(n15596), .B2(DATAI_23_), 
        .ZN(n15568) );
  OAI211_X1 U19122 ( .C1(n15570), .C2(n15610), .A(n15569), .B(n15568), .ZN(
        P1_U2881) );
  AOI22_X1 U19123 ( .A1(n15595), .A2(BUF1_REG_22__SCAN_IN), .B1(
        P1_EAX_REG_22__SCAN_IN), .B2(n15606), .ZN(n15573) );
  AOI22_X1 U19124 ( .A1(n15598), .A2(n15571), .B1(n15596), .B2(DATAI_22_), 
        .ZN(n15572) );
  OAI211_X1 U19125 ( .C1(n15574), .C2(n15610), .A(n15573), .B(n15572), .ZN(
        P1_U2882) );
  AOI22_X1 U19126 ( .A1(n15595), .A2(BUF1_REG_21__SCAN_IN), .B1(
        P1_EAX_REG_21__SCAN_IN), .B2(n15606), .ZN(n15577) );
  AOI22_X1 U19127 ( .A1(n15598), .A2(n15575), .B1(n15596), .B2(DATAI_21_), 
        .ZN(n15576) );
  OAI211_X1 U19128 ( .C1(n16665), .C2(n15610), .A(n15577), .B(n15576), .ZN(
        P1_U2883) );
  AOI22_X1 U19129 ( .A1(n15595), .A2(BUF1_REG_20__SCAN_IN), .B1(
        P1_EAX_REG_20__SCAN_IN), .B2(n15606), .ZN(n15580) );
  AOI22_X1 U19130 ( .A1(n15598), .A2(n15578), .B1(n15596), .B2(DATAI_20_), 
        .ZN(n15579) );
  OAI211_X1 U19131 ( .C1(n16567), .C2(n15610), .A(n15580), .B(n15579), .ZN(
        P1_U2884) );
  NOR2_X1 U19132 ( .A1(n15582), .A2(n15581), .ZN(n15583) );
  AOI22_X1 U19133 ( .A1(n15595), .A2(BUF1_REG_19__SCAN_IN), .B1(
        P1_EAX_REG_19__SCAN_IN), .B2(n15606), .ZN(n15587) );
  AOI22_X1 U19134 ( .A1(n15598), .A2(n15585), .B1(n15596), .B2(DATAI_19_), 
        .ZN(n15586) );
  OAI211_X1 U19135 ( .C1(n16677), .C2(n15610), .A(n15587), .B(n15586), .ZN(
        P1_U2885) );
  AOI22_X1 U19136 ( .A1(n15595), .A2(BUF1_REG_18__SCAN_IN), .B1(
        P1_EAX_REG_18__SCAN_IN), .B2(n15606), .ZN(n15590) );
  AOI22_X1 U19137 ( .A1(n15598), .A2(n15588), .B1(n15596), .B2(DATAI_18_), 
        .ZN(n15589) );
  OAI211_X1 U19138 ( .C1(n16591), .C2(n15610), .A(n15590), .B(n15589), .ZN(
        P1_U2886) );
  AOI22_X1 U19139 ( .A1(n15595), .A2(BUF1_REG_17__SCAN_IN), .B1(
        P1_EAX_REG_17__SCAN_IN), .B2(n15606), .ZN(n15593) );
  AOI22_X1 U19140 ( .A1(n15598), .A2(n15591), .B1(n15596), .B2(DATAI_17_), 
        .ZN(n15592) );
  OAI211_X1 U19141 ( .C1(n15594), .C2(n15610), .A(n15593), .B(n15592), .ZN(
        P1_U2887) );
  AOI22_X1 U19142 ( .A1(n15595), .A2(BUF1_REG_16__SCAN_IN), .B1(
        P1_EAX_REG_16__SCAN_IN), .B2(n15606), .ZN(n15600) );
  AOI22_X1 U19143 ( .A1(n15598), .A2(n15597), .B1(n15596), .B2(DATAI_16_), 
        .ZN(n15599) );
  OAI211_X1 U19144 ( .C1(n15601), .C2(n15610), .A(n15600), .B(n15599), .ZN(
        P1_U2888) );
  OAI222_X1 U19145 ( .A1(n16701), .A2(n15610), .B1(n15605), .B2(n15604), .C1(
        n15603), .C2(n15602), .ZN(P1_U2889) );
  AOI22_X1 U19146 ( .A1(n15608), .A2(n15607), .B1(P1_EAX_REG_14__SCAN_IN), 
        .B2(n15606), .ZN(n15609) );
  OAI21_X1 U19147 ( .B1(n15611), .B2(n15610), .A(n15609), .ZN(P1_U2890) );
  NAND2_X1 U19148 ( .A1(n15612), .A2(n16739), .ZN(n15618) );
  NOR2_X1 U19149 ( .A1(n16670), .A2(n15613), .ZN(n15614) );
  AOI211_X1 U19150 ( .C1(n16722), .C2(n15616), .A(n15615), .B(n15614), .ZN(
        n15617) );
  OAI211_X1 U19151 ( .C1(n15619), .C2(n20773), .A(n15618), .B(n15617), .ZN(
        P1_U2969) );
  XNOR2_X1 U19152 ( .A(n15620), .B(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15707) );
  NAND2_X1 U19153 ( .A1(n15621), .A2(n16739), .ZN(n15626) );
  NOR2_X1 U19154 ( .A1(n16823), .A2(n21242), .ZN(n15703) );
  INV_X1 U19155 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n15622) );
  NOR2_X1 U19156 ( .A1(n16670), .A2(n15622), .ZN(n15623) );
  AOI211_X1 U19157 ( .C1(n16722), .C2(n15624), .A(n15703), .B(n15623), .ZN(
        n15625) );
  OAI211_X1 U19158 ( .C1(n15707), .C2(n20773), .A(n15626), .B(n15625), .ZN(
        P1_U2973) );
  AOI21_X1 U19159 ( .B1(n15627), .B2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n16673), .ZN(n15628) );
  NOR2_X1 U19160 ( .A1(n15629), .A2(n15628), .ZN(n15631) );
  AOI22_X1 U19161 ( .A1(n16673), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .B1(
        n11661), .B2(n16645), .ZN(n15630) );
  XNOR2_X1 U19162 ( .A(n15631), .B(n15630), .ZN(n15714) );
  INV_X1 U19163 ( .A(n16537), .ZN(n15635) );
  INV_X1 U19164 ( .A(n16532), .ZN(n15633) );
  AOI22_X1 U19165 ( .A1(n16734), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .B1(
        n16782), .B2(P1_REIP_REG_24__SCAN_IN), .ZN(n15632) );
  OAI21_X1 U19166 ( .B1(n15633), .B2(n16743), .A(n15632), .ZN(n15634) );
  AOI21_X1 U19167 ( .B1(n15635), .B2(n16739), .A(n15634), .ZN(n15636) );
  OAI21_X1 U19168 ( .B1(n20773), .B2(n15714), .A(n15636), .ZN(P1_U2975) );
  INV_X1 U19169 ( .A(n15637), .ZN(n15638) );
  NOR2_X1 U19170 ( .A1(n15639), .A2(n15638), .ZN(n15640) );
  XNOR2_X1 U19171 ( .A(n15640), .B(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n16760) );
  INV_X1 U19172 ( .A(n16549), .ZN(n15642) );
  AOI22_X1 U19173 ( .A1(n16734), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B1(
        n16782), .B2(P1_REIP_REG_22__SCAN_IN), .ZN(n15641) );
  OAI21_X1 U19174 ( .B1(n15642), .B2(n16743), .A(n15641), .ZN(n15643) );
  AOI21_X1 U19175 ( .B1(n16550), .B2(n16739), .A(n15643), .ZN(n15644) );
  OAI21_X1 U19176 ( .B1(n20773), .B2(n16760), .A(n15644), .ZN(P1_U2977) );
  NOR2_X1 U19177 ( .A1(n16673), .A2(n16674), .ZN(n15646) );
  NAND2_X1 U19178 ( .A1(n15645), .A2(n15646), .ZN(n15715) );
  NOR2_X1 U19179 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15647) );
  AND2_X1 U19180 ( .A1(n16673), .A2(n15647), .ZN(n15648) );
  NAND2_X1 U19181 ( .A1(n11461), .A2(n15648), .ZN(n15717) );
  NAND2_X1 U19182 ( .A1(n15715), .A2(n15717), .ZN(n15649) );
  XOR2_X1 U19183 ( .A(n15716), .B(n15649), .Z(n15730) );
  INV_X1 U19184 ( .A(n16563), .ZN(n15651) );
  AOI22_X1 U19185 ( .A1(n16734), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B1(
        n16782), .B2(P1_REIP_REG_20__SCAN_IN), .ZN(n15650) );
  OAI21_X1 U19186 ( .B1(n15651), .B2(n16743), .A(n15650), .ZN(n15652) );
  AOI21_X1 U19187 ( .B1(n15653), .B2(n16739), .A(n15652), .ZN(n15654) );
  OAI21_X1 U19188 ( .B1(n20773), .B2(n15730), .A(n15654), .ZN(P1_U2979) );
  INV_X1 U19189 ( .A(n15655), .ZN(n16588) );
  INV_X1 U19190 ( .A(P1_REIP_REG_18__SCAN_IN), .ZN(n15656) );
  NOR2_X1 U19191 ( .A1(n16823), .A2(n15656), .ZN(n15739) );
  NOR2_X1 U19192 ( .A1(n16670), .A2(n15657), .ZN(n15658) );
  AOI211_X1 U19193 ( .C1(n16588), .C2(n16722), .A(n15739), .B(n15658), .ZN(
        n15662) );
  INV_X1 U19194 ( .A(n15645), .ZN(n16672) );
  OR2_X1 U19195 ( .A1(n15660), .A2(n15659), .ZN(n15731) );
  NAND3_X1 U19196 ( .A1(n16672), .A2(n16740), .A3(n15731), .ZN(n15661) );
  OAI211_X1 U19197 ( .C1(n16591), .C2(n16700), .A(n15662), .B(n15661), .ZN(
        P1_U2981) );
  INV_X1 U19198 ( .A(n15663), .ZN(n15677) );
  NOR2_X1 U19199 ( .A1(n15677), .A2(n15664), .ZN(n15758) );
  INV_X1 U19200 ( .A(n15665), .ZN(n15667) );
  OAI21_X1 U19201 ( .B1(n15758), .B2(n15667), .A(n15666), .ZN(n15669) );
  AOI22_X1 U19202 ( .A1(n16673), .A2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B1(
        n15763), .B2(n16645), .ZN(n15668) );
  XNOR2_X1 U19203 ( .A(n15669), .B(n15668), .ZN(n15775) );
  AOI22_X1 U19204 ( .A1(n16734), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        n16782), .B2(P1_REIP_REG_14__SCAN_IN), .ZN(n15670) );
  OAI21_X1 U19205 ( .B1(n15671), .B2(n16743), .A(n15670), .ZN(n15672) );
  AOI21_X1 U19206 ( .B1(n15673), .B2(n16739), .A(n15672), .ZN(n15674) );
  OAI21_X1 U19207 ( .B1(n15775), .B2(n20773), .A(n15674), .ZN(P1_U2985) );
  INV_X1 U19208 ( .A(n15675), .ZN(n15678) );
  MUX2_X1 U19209 ( .A(n15677), .B(n15678), .S(n15676), .Z(n15797) );
  NAND2_X1 U19210 ( .A1(n15797), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n15796) );
  NAND3_X1 U19211 ( .A1(n15678), .A2(n16673), .A3(n15796), .ZN(n15679) );
  OAI21_X1 U19212 ( .B1(n16673), .B2(n15796), .A(n15679), .ZN(n15680) );
  XNOR2_X1 U19213 ( .A(n15680), .B(n16806), .ZN(n16803) );
  NAND2_X1 U19214 ( .A1(n16803), .A2(n16740), .ZN(n15685) );
  INV_X1 U19215 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n15681) );
  NOR2_X1 U19216 ( .A1(n16823), .A2(n15681), .ZN(n16799) );
  NOR2_X1 U19217 ( .A1(n16743), .A2(n15682), .ZN(n15683) );
  AOI211_X1 U19218 ( .C1(n16734), .C2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n16799), .B(n15683), .ZN(n15684) );
  OAI211_X1 U19219 ( .C1(n16700), .C2(n15686), .A(n15685), .B(n15684), .ZN(
        P1_U2988) );
  INV_X1 U19220 ( .A(n15687), .ZN(n15695) );
  INV_X1 U19221 ( .A(n15688), .ZN(n15694) );
  AOI211_X1 U19222 ( .C1(n15692), .C2(n15691), .A(n15690), .B(n15689), .ZN(
        n15693) );
  AOI211_X1 U19223 ( .C1(n15695), .C2(n16809), .A(n15694), .B(n15693), .ZN(
        n15698) );
  NAND2_X1 U19224 ( .A1(n15696), .A2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15697) );
  OAI211_X1 U19225 ( .C1(n15699), .C2(n16792), .A(n15698), .B(n15697), .ZN(
        P1_U3003) );
  NOR3_X1 U19226 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n15700), .A3(
        n16758), .ZN(n16744) );
  OAI22_X1 U19227 ( .A1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n15702), .B1(
        n16744), .B2(n15701), .ZN(n15706) );
  AOI21_X1 U19228 ( .B1(n15704), .B2(n16809), .A(n15703), .ZN(n15705) );
  OAI211_X1 U19229 ( .C1(n15707), .C2(n16792), .A(n15706), .B(n15705), .ZN(
        P1_U3005) );
  INV_X1 U19230 ( .A(n16541), .ZN(n15712) );
  OAI221_X1 U19231 ( .B1(n15708), .B2(n15783), .C1(n15708), .C2(n9980), .A(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15709) );
  OAI21_X1 U19232 ( .B1(n16823), .B2(n21239), .A(n15709), .ZN(n15711) );
  NOR3_X1 U19233 ( .A1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n9980), .A3(
        n16758), .ZN(n15710) );
  AOI211_X1 U19234 ( .C1(n16809), .C2(n15712), .A(n15711), .B(n15710), .ZN(
        n15713) );
  OAI21_X1 U19235 ( .B1(n15714), .B2(n16792), .A(n15713), .ZN(P1_U3007) );
  NAND2_X1 U19236 ( .A1(n15715), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15719) );
  NAND2_X1 U19237 ( .A1(n15717), .A2(n15716), .ZN(n15718) );
  NAND2_X1 U19238 ( .A1(n15719), .A2(n15718), .ZN(n15720) );
  XNOR2_X1 U19239 ( .A(n15720), .B(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n16661) );
  INV_X1 U19240 ( .A(n16661), .ZN(n15724) );
  OAI22_X1 U19241 ( .A1(n16556), .A2(n20925), .B1(n16823), .B2(n21234), .ZN(
        n15721) );
  AOI21_X1 U19242 ( .B1(n11460), .B2(n16764), .A(n15721), .ZN(n15723) );
  NAND2_X1 U19243 ( .A1(n16759), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15722) );
  OAI211_X1 U19244 ( .C1(n15724), .C2(n16792), .A(n15723), .B(n15722), .ZN(
        P1_U3010) );
  INV_X1 U19245 ( .A(n15725), .ZN(n16768) );
  OAI22_X1 U19246 ( .A1(n16566), .A2(n20925), .B1(n21232), .B2(n16823), .ZN(
        n15728) );
  NOR3_X1 U19247 ( .A1(n16774), .A2(n15726), .A3(n10216), .ZN(n15727) );
  AOI211_X1 U19248 ( .C1(n16768), .C2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n15728), .B(n15727), .ZN(n15729) );
  OAI21_X1 U19249 ( .B1(n15730), .B2(n16792), .A(n15729), .ZN(P1_U3011) );
  NAND3_X1 U19250 ( .A1(n16672), .A2(n20927), .A3(n15731), .ZN(n15745) );
  AOI21_X1 U19251 ( .B1(n15733), .B2(n15769), .A(n15732), .ZN(n15734) );
  OAI21_X1 U19252 ( .B1(n15736), .B2(n15735), .A(n15734), .ZN(n15773) );
  INV_X1 U19253 ( .A(n15773), .ZN(n16797) );
  OAI21_X1 U19254 ( .B1(n15738), .B2(n15737), .A(n16797), .ZN(n15753) );
  INV_X1 U19255 ( .A(n15739), .ZN(n15740) );
  OAI21_X1 U19256 ( .B1(n16597), .B2(n20925), .A(n15740), .ZN(n15743) );
  NAND2_X1 U19257 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n16780) );
  NAND2_X1 U19258 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n15741), .ZN(
        n16775) );
  NOR4_X1 U19259 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n15752), .A3(
        n16780), .A4(n16775), .ZN(n15742) );
  AOI211_X1 U19260 ( .C1(n15753), .C2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n15743), .B(n15742), .ZN(n15744) );
  NAND2_X1 U19261 ( .A1(n15745), .A2(n15744), .ZN(P1_U3013) );
  NOR2_X1 U19262 ( .A1(n16645), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15749) );
  AOI21_X1 U19263 ( .B1(n15747), .B2(n15663), .A(n15746), .ZN(n15748) );
  MUX2_X1 U19264 ( .A(n15749), .B(n16645), .S(n15748), .Z(n15750) );
  XNOR2_X1 U19265 ( .A(n15750), .B(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n16686) );
  AOI22_X1 U19266 ( .A1(n15751), .A2(n16809), .B1(n16782), .B2(
        P1_REIP_REG_17__SCAN_IN), .ZN(n15756) );
  OAI21_X1 U19267 ( .B1(n16780), .B2(n16775), .A(n15752), .ZN(n15754) );
  NAND2_X1 U19268 ( .A1(n15754), .A2(n15753), .ZN(n15755) );
  OAI211_X1 U19269 ( .C1(n16686), .C2(n16792), .A(n15756), .B(n15755), .ZN(
        P1_U3014) );
  NOR2_X1 U19270 ( .A1(n15758), .A2(n15757), .ZN(n16688) );
  INV_X1 U19271 ( .A(n15759), .ZN(n15760) );
  NOR2_X1 U19272 ( .A1(n16688), .A2(n15760), .ZN(n15762) );
  AOI22_X1 U19273 ( .A1(n16673), .A2(n15765), .B1(
        P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n16645), .ZN(n15761) );
  XNOR2_X1 U19274 ( .A(n15762), .B(n15761), .ZN(n16705) );
  NAND2_X1 U19275 ( .A1(n16782), .A2(P1_REIP_REG_15__SCAN_IN), .ZN(n15764) );
  OAI221_X1 U19276 ( .B1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n16775), 
        .C1(n15765), .C2(n16786), .A(n15764), .ZN(n15766) );
  AOI21_X1 U19277 ( .B1(n16608), .B2(n16809), .A(n15766), .ZN(n15767) );
  OAI21_X1 U19278 ( .B1(n16705), .B2(n16792), .A(n15767), .ZN(P1_U3016) );
  OAI22_X1 U19279 ( .A1(n15768), .A2(n20925), .B1(n21222), .B2(n16823), .ZN(
        n15772) );
  NOR3_X1 U19280 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n15770), .A3(
        n15769), .ZN(n15771) );
  AOI211_X1 U19281 ( .C1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n15773), .A(
        n15772), .B(n15771), .ZN(n15774) );
  OAI21_X1 U19282 ( .B1(n15775), .B2(n16792), .A(n15774), .ZN(P1_U3017) );
  INV_X1 U19283 ( .A(n15776), .ZN(n15777) );
  OAI21_X1 U19284 ( .B1(n15663), .B2(n15778), .A(n15777), .ZN(n15781) );
  OR2_X1 U19285 ( .A1(n16707), .A2(n15779), .ZN(n15780) );
  NOR2_X1 U19286 ( .A1(n15781), .A2(n15780), .ZN(n16706) );
  AOI21_X1 U19287 ( .B1(n15781), .B2(n15780), .A(n16706), .ZN(n16719) );
  INV_X1 U19288 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n15782) );
  NAND3_X1 U19289 ( .A1(n15786), .A2(n16822), .A3(n15782), .ZN(n15795) );
  INV_X1 U19290 ( .A(n15783), .ZN(n15790) );
  INV_X1 U19291 ( .A(n15799), .ZN(n15785) );
  OAI221_X1 U19292 ( .B1(n20929), .B2(n15786), .C1(n20929), .C2(n15785), .A(
        n15784), .ZN(n15787) );
  AOI221_X1 U19293 ( .B1(n15789), .B2(n15788), .C1(n16801), .C2(n15788), .A(
        n15787), .ZN(n16807) );
  OAI21_X1 U19294 ( .B1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n15790), .A(
        n16807), .ZN(n15793) );
  OAI22_X1 U19295 ( .A1(n15791), .A2(n20925), .B1(n21217), .B2(n16823), .ZN(
        n15792) );
  AOI21_X1 U19296 ( .B1(n15793), .B2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n15792), .ZN(n15794) );
  OAI211_X1 U19297 ( .C1(n16719), .C2(n16792), .A(n15795), .B(n15794), .ZN(
        P1_U3019) );
  OAI21_X1 U19298 ( .B1(n15797), .B2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n15796), .ZN(n16726) );
  NOR2_X1 U19299 ( .A1(n15799), .A2(n15798), .ZN(n15801) );
  AOI21_X1 U19300 ( .B1(n15801), .B2(n15802), .A(n15800), .ZN(n16811) );
  OAI22_X1 U19301 ( .A1(n16635), .A2(n20925), .B1(n21215), .B2(n16823), .ZN(
        n15805) );
  INV_X1 U19302 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15803) );
  NAND2_X1 U19303 ( .A1(n15802), .A2(n16822), .ZN(n16815) );
  AOI221_X1 U19304 ( .B1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .C1(n11451), .C2(n15803), .A(
        n16815), .ZN(n15804) );
  AOI211_X1 U19305 ( .C1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .C2(n16811), .A(
        n15805), .B(n15804), .ZN(n15806) );
  OAI21_X1 U19306 ( .B1(n16726), .B2(n16792), .A(n15806), .ZN(P1_U3021) );
  OAI211_X1 U19307 ( .C1(P1_STATEBS16_REG_SCAN_IN), .C2(n15812), .A(n15809), 
        .B(n21085), .ZN(n15807) );
  OAI21_X1 U19308 ( .B1(n14001), .B2(n15818), .A(n15807), .ZN(n15808) );
  MUX2_X1 U19309 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n15808), .S(
        n20938), .Z(P1_U3477) );
  XNOR2_X1 U19310 ( .A(n13856), .B(n15809), .ZN(n15810) );
  OAI22_X1 U19311 ( .A1(n15810), .A2(n21122), .B1(n9734), .B2(n15818), .ZN(
        n15811) );
  MUX2_X1 U19312 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n15811), .S(
        n20938), .Z(P1_U3476) );
  NOR3_X1 U19313 ( .A1(n21008), .A2(n21122), .A3(n21118), .ZN(n21058) );
  NAND2_X1 U19314 ( .A1(n21058), .A2(n15812), .ZN(n15817) );
  INV_X1 U19315 ( .A(n15813), .ZN(n15814) );
  NAND3_X1 U19316 ( .A1(n15815), .A2(n15814), .A3(n21085), .ZN(n15816) );
  OAI211_X1 U19317 ( .C1(n15819), .C2(n15818), .A(n15817), .B(n15816), .ZN(
        n15820) );
  MUX2_X1 U19318 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B(n15820), .S(
        n20938), .Z(P1_U3475) );
  NOR3_X1 U19319 ( .A1(n15821), .A2(n15828), .A3(n13305), .ZN(n15822) );
  AOI211_X1 U19320 ( .C1(n20945), .C2(n15824), .A(n15823), .B(n15822), .ZN(
        n16476) );
  INV_X1 U19321 ( .A(n21270), .ZN(n15833) );
  INV_X1 U19322 ( .A(n15825), .ZN(n15826) );
  NAND2_X1 U19323 ( .A1(n15827), .A2(n15826), .ZN(n15832) );
  INV_X1 U19324 ( .A(n15828), .ZN(n15830) );
  INV_X1 U19325 ( .A(n13305), .ZN(n15829) );
  NAND3_X1 U19326 ( .A1(n15830), .A2(n21268), .A3(n15829), .ZN(n15831) );
  OAI211_X1 U19327 ( .C1(n16476), .C2(n15833), .A(n15832), .B(n15831), .ZN(
        n15835) );
  MUX2_X1 U19328 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n15835), .S(
        n15834), .Z(P1_U3473) );
  NOR2_X1 U19329 ( .A1(n15858), .A2(n15837), .ZN(n15838) );
  OR2_X1 U19330 ( .A1(n15836), .A2(n15838), .ZN(n15969) );
  INV_X1 U19331 ( .A(n15969), .ZN(n16233) );
  INV_X1 U19332 ( .A(n19917), .ZN(n19888) );
  OAI211_X1 U19333 ( .C1(n16055), .C2(n15840), .A(n19910), .B(n15839), .ZN(
        n15844) );
  OAI22_X1 U19334 ( .A1(n15841), .A2(n19815), .B1(n20670), .B2(n19887), .ZN(
        n15842) );
  INV_X1 U19335 ( .A(n15842), .ZN(n15843) );
  OAI211_X1 U19336 ( .C1(n19888), .C2(n11004), .A(n15844), .B(n15843), .ZN(
        n15849) );
  NOR2_X1 U19337 ( .A1(n15856), .A2(n15846), .ZN(n15847) );
  OR2_X1 U19338 ( .A1(n15845), .A2(n15847), .ZN(n16237) );
  NOR2_X1 U19339 ( .A1(n16237), .A2(n19880), .ZN(n15848) );
  AOI211_X1 U19340 ( .C1(n19915), .C2(n16233), .A(n15849), .B(n15848), .ZN(
        n15850) );
  OAI21_X1 U19341 ( .B1(n15851), .B2(n19919), .A(n15850), .ZN(P2_U2830) );
  OAI211_X1 U19342 ( .C1(n15853), .C2(n16066), .A(n19897), .B(n15852), .ZN(
        n15864) );
  AND2_X1 U19343 ( .A1(n15855), .A2(n15854), .ZN(n15857) );
  OR2_X1 U19344 ( .A1(n15857), .A2(n15856), .ZN(n16246) );
  INV_X1 U19345 ( .A(n16246), .ZN(n16915) );
  OAI22_X1 U19346 ( .A1(n16068), .A2(n19815), .B1(n20668), .B2(n19887), .ZN(
        n15862) );
  AOI21_X1 U19347 ( .B1(n15859), .B2(n15978), .A(n15858), .ZN(n16934) );
  INV_X1 U19348 ( .A(n16934), .ZN(n15860) );
  OAI22_X1 U19349 ( .A1(n15860), .A2(n19914), .B1(n19888), .B2(n10814), .ZN(
        n15861) );
  AOI211_X1 U19350 ( .C1(n16915), .C2(n19922), .A(n15862), .B(n15861), .ZN(
        n15863) );
  OAI211_X1 U19351 ( .C1(n15865), .C2(n19919), .A(n15864), .B(n15863), .ZN(
        P2_U2831) );
  INV_X1 U19352 ( .A(n20044), .ZN(n15868) );
  NOR2_X1 U19353 ( .A1(n9766), .A2(n15866), .ZN(n15878) );
  INV_X1 U19354 ( .A(n15878), .ZN(n15867) );
  AOI221_X1 U19355 ( .B1(n15868), .B2(n15878), .C1(n20044), .C2(n15867), .A(
        n20613), .ZN(n15869) );
  INV_X1 U19356 ( .A(n15869), .ZN(n15877) );
  NAND2_X1 U19357 ( .A1(n19917), .A2(P2_EBX_REG_2__SCAN_IN), .ZN(n15871) );
  AOI22_X1 U19358 ( .A1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n19929), .B1(
        P2_REIP_REG_2__SCAN_IN), .B2(n19927), .ZN(n15870) );
  OAI211_X1 U19359 ( .C1(n19919), .C2(n15872), .A(n15871), .B(n15870), .ZN(
        n15875) );
  NOR2_X1 U19360 ( .A1(n15873), .A2(n19880), .ZN(n15874) );
  AOI211_X1 U19361 ( .C1(n19915), .C2(n20708), .A(n15875), .B(n15874), .ZN(
        n15876) );
  OAI211_X1 U19362 ( .C1(n20706), .C2(n19925), .A(n15877), .B(n15876), .ZN(
        P2_U2853) );
  OAI21_X1 U19363 ( .B1(n19933), .B2(n15879), .A(n15878), .ZN(n16423) );
  NOR2_X1 U19364 ( .A1(n9719), .A2(n20613), .ZN(n19928) );
  OAI22_X1 U19365 ( .A1(n15883), .A2(n19815), .B1(n10371), .B2(n19887), .ZN(
        n15882) );
  NOR2_X1 U19366 ( .A1(n19919), .A2(n15880), .ZN(n15881) );
  AOI211_X1 U19367 ( .C1(n19928), .C2(n15883), .A(n15882), .B(n15881), .ZN(
        n15885) );
  NAND2_X1 U19368 ( .A1(n20712), .A2(n19915), .ZN(n15884) );
  OAI211_X1 U19369 ( .C1(n19888), .C2(n10557), .A(n15885), .B(n15884), .ZN(
        n15887) );
  NOR2_X1 U19370 ( .A1(n20074), .A2(n19925), .ZN(n15886) );
  AOI211_X1 U19371 ( .C1(n19922), .C2(n15888), .A(n15887), .B(n15886), .ZN(
        n15889) );
  OAI21_X1 U19372 ( .B1(n16423), .B2(n20613), .A(n15889), .ZN(P2_U2854) );
  XNOR2_X1 U19373 ( .A(n15891), .B(n15890), .ZN(n15941) );
  OAI21_X1 U19374 ( .B1(n15894), .B2(n15893), .A(n15892), .ZN(n16856) );
  NOR2_X1 U19375 ( .A1(n16856), .A2(n19947), .ZN(n15895) );
  AOI21_X1 U19376 ( .B1(P2_EBX_REG_29__SCAN_IN), .B2(n19947), .A(n15895), .ZN(
        n15896) );
  OAI21_X1 U19377 ( .B1(n15941), .B2(n19959), .A(n15896), .ZN(P2_U2858) );
  INV_X1 U19378 ( .A(n15897), .ZN(n15898) );
  NOR2_X1 U19379 ( .A1(n15899), .A2(n15898), .ZN(n15901) );
  XNOR2_X1 U19380 ( .A(n15901), .B(n15900), .ZN(n15948) );
  NAND2_X1 U19381 ( .A1(n19947), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n15903) );
  NAND2_X1 U19382 ( .A1(n16869), .A2(n19969), .ZN(n15902) );
  OAI211_X1 U19383 ( .C1(n15948), .C2(n19959), .A(n15903), .B(n15902), .ZN(
        P2_U2859) );
  AOI21_X1 U19384 ( .B1(n15906), .B2(n15905), .A(n15904), .ZN(n15949) );
  NAND2_X1 U19385 ( .A1(n15949), .A2(n16926), .ZN(n15908) );
  NAND2_X1 U19386 ( .A1(n19947), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n15907) );
  OAI211_X1 U19387 ( .C1(n15909), .C2(n19947), .A(n15908), .B(n15907), .ZN(
        P2_U2860) );
  OR2_X1 U19388 ( .A1(n15845), .A2(n15910), .ZN(n15911) );
  NAND2_X1 U19389 ( .A1(n13036), .A2(n15911), .ZN(n16890) );
  AOI21_X1 U19390 ( .B1(n15914), .B2(n15913), .A(n15912), .ZN(n15957) );
  NAND2_X1 U19391 ( .A1(n15957), .A2(n16926), .ZN(n15916) );
  NAND2_X1 U19392 ( .A1(n19947), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n15915) );
  OAI211_X1 U19393 ( .C1(n19947), .C2(n16890), .A(n15916), .B(n15915), .ZN(
        P2_U2861) );
  XNOR2_X1 U19394 ( .A(n15918), .B(n15917), .ZN(n15974) );
  MUX2_X1 U19395 ( .A(n16237), .B(n11004), .S(n19947), .Z(n15919) );
  OAI21_X1 U19396 ( .B1(n15974), .B2(n19959), .A(n15919), .ZN(P2_U2862) );
  OAI21_X1 U19397 ( .B1(n15922), .B2(n15921), .A(n15920), .ZN(n15986) );
  NAND2_X1 U19398 ( .A1(n19947), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n15924) );
  NAND2_X1 U19399 ( .A1(n16902), .A2(n19969), .ZN(n15923) );
  OAI211_X1 U19400 ( .C1(n15986), .C2(n19959), .A(n15924), .B(n15923), .ZN(
        P2_U2864) );
  OR2_X1 U19401 ( .A1(n9819), .A2(n15925), .ZN(n15926) );
  NAND2_X1 U19402 ( .A1(n14749), .A2(n15926), .ZN(n16463) );
  INV_X1 U19403 ( .A(n15927), .ZN(n15928) );
  AOI21_X1 U19404 ( .B1(n15929), .B2(n15997), .A(n15928), .ZN(n15987) );
  NAND2_X1 U19405 ( .A1(n15987), .A2(n16926), .ZN(n15931) );
  NAND2_X1 U19406 ( .A1(n19947), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n15930) );
  OAI211_X1 U19407 ( .C1(n16463), .C2(n19947), .A(n15931), .B(n15930), .ZN(
        P2_U2865) );
  XOR2_X1 U19408 ( .A(n15933), .B(n15932), .Z(n16857) );
  INV_X1 U19409 ( .A(BUF2_REG_29__SCAN_IN), .ZN(n15938) );
  OAI22_X1 U19410 ( .A1(n16930), .A2(n15935), .B1(n19979), .B2(n15934), .ZN(
        n15936) );
  AOI21_X1 U19411 ( .B1(n16932), .B2(BUF1_REG_29__SCAN_IN), .A(n15936), .ZN(
        n15937) );
  OAI21_X1 U19412 ( .B1(n16015), .B2(n15938), .A(n15937), .ZN(n15939) );
  AOI21_X1 U19413 ( .B1(n16857), .B2(n16935), .A(n15939), .ZN(n15940) );
  OAI21_X1 U19414 ( .B1(n15941), .B2(n19982), .A(n15940), .ZN(P2_U2890) );
  OAI22_X1 U19415 ( .A1(n16930), .A2(n15943), .B1(n16020), .B2(n15942), .ZN(
        n15945) );
  NOR2_X1 U19416 ( .A1(n16867), .A2(n16023), .ZN(n15944) );
  AOI211_X1 U19417 ( .C1(BUF1_REG_28__SCAN_IN), .C2(n16932), .A(n15945), .B(
        n15944), .ZN(n15947) );
  NAND2_X1 U19418 ( .A1(n16933), .A2(BUF2_REG_28__SCAN_IN), .ZN(n15946) );
  OAI211_X1 U19419 ( .C1(n15948), .C2(n19982), .A(n15947), .B(n15946), .ZN(
        P2_U2891) );
  INV_X1 U19420 ( .A(BUF2_REG_27__SCAN_IN), .ZN(n15956) );
  NAND2_X1 U19421 ( .A1(n15949), .A2(n16936), .ZN(n15955) );
  OAI22_X1 U19422 ( .A1(n16930), .A2(n15951), .B1(n16020), .B2(n15950), .ZN(
        n15953) );
  NOR2_X1 U19423 ( .A1(n16888), .A2(n16023), .ZN(n15952) );
  AOI211_X1 U19424 ( .C1(BUF1_REG_27__SCAN_IN), .C2(n16932), .A(n15953), .B(
        n15952), .ZN(n15954) );
  OAI211_X1 U19425 ( .C1(n16015), .C2(n15956), .A(n15955), .B(n15954), .ZN(
        P2_U2892) );
  INV_X1 U19426 ( .A(BUF2_REG_26__SCAN_IN), .ZN(n15966) );
  NAND2_X1 U19427 ( .A1(n15957), .A2(n16936), .ZN(n15965) );
  OAI22_X1 U19428 ( .A1(n16930), .A2(n15959), .B1(n16020), .B2(n15958), .ZN(
        n15963) );
  NOR2_X1 U19429 ( .A1(n15836), .A2(n15960), .ZN(n15961) );
  OR2_X1 U19430 ( .A1(n13038), .A2(n15961), .ZN(n16220) );
  NOR2_X1 U19431 ( .A1(n16220), .A2(n16023), .ZN(n15962) );
  AOI211_X1 U19432 ( .C1(BUF1_REG_26__SCAN_IN), .C2(n16932), .A(n15963), .B(
        n15962), .ZN(n15964) );
  OAI211_X1 U19433 ( .C1(n16015), .C2(n15966), .A(n15965), .B(n15964), .ZN(
        P2_U2893) );
  OAI22_X1 U19434 ( .A1(n16930), .A2(n15968), .B1(n16020), .B2(n15967), .ZN(
        n15971) );
  NOR2_X1 U19435 ( .A1(n15969), .A2(n16023), .ZN(n15970) );
  AOI211_X1 U19436 ( .C1(BUF1_REG_25__SCAN_IN), .C2(n16932), .A(n15971), .B(
        n15970), .ZN(n15973) );
  NAND2_X1 U19437 ( .A1(n16933), .A2(BUF2_REG_25__SCAN_IN), .ZN(n15972) );
  OAI211_X1 U19438 ( .C1(n15974), .C2(n19982), .A(n15973), .B(n15972), .ZN(
        P2_U2894) );
  INV_X1 U19439 ( .A(BUF2_REG_23__SCAN_IN), .ZN(n15983) );
  NAND2_X1 U19440 ( .A1(n15975), .A2(n15976), .ZN(n15977) );
  AND2_X1 U19441 ( .A1(n15978), .A2(n15977), .ZN(n16901) );
  OAI22_X1 U19442 ( .A1(n16930), .A2(n20123), .B1(n16020), .B2(n15979), .ZN(
        n15980) );
  AOI21_X1 U19443 ( .B1(n16901), .B2(n16935), .A(n15980), .ZN(n15982) );
  NAND2_X1 U19444 ( .A1(n16932), .A2(BUF1_REG_23__SCAN_IN), .ZN(n15981) );
  OAI211_X1 U19445 ( .C1(n16015), .C2(n15983), .A(n15982), .B(n15981), .ZN(
        n15984) );
  INV_X1 U19446 ( .A(n15984), .ZN(n15985) );
  OAI21_X1 U19447 ( .B1(n15986), .B2(n19982), .A(n15985), .ZN(P2_U2896) );
  NAND2_X1 U19448 ( .A1(n15987), .A2(n16936), .ZN(n15996) );
  NAND2_X1 U19449 ( .A1(n15988), .A2(n15989), .ZN(n15990) );
  AND2_X1 U19450 ( .A1(n15975), .A2(n15990), .ZN(n16461) );
  OAI22_X1 U19451 ( .A1(n16930), .A2(n20115), .B1(n16020), .B2(n15991), .ZN(
        n15992) );
  AOI21_X1 U19452 ( .B1(n16461), .B2(n16935), .A(n15992), .ZN(n15995) );
  NAND2_X1 U19453 ( .A1(n16933), .A2(BUF2_REG_22__SCAN_IN), .ZN(n15994) );
  NAND2_X1 U19454 ( .A1(n16932), .A2(BUF1_REG_22__SCAN_IN), .ZN(n15993) );
  NAND4_X1 U19455 ( .A1(n15996), .A2(n15995), .A3(n15994), .A4(n15993), .ZN(
        P2_U2897) );
  OAI21_X1 U19456 ( .B1(n14903), .B2(n15998), .A(n15997), .ZN(n16917) );
  OAI22_X1 U19457 ( .A1(n16930), .A2(n20108), .B1(n16020), .B2(n15999), .ZN(
        n16003) );
  OAI21_X1 U19458 ( .B1(n16000), .B2(n16001), .A(n15988), .ZN(n19754) );
  NOR2_X1 U19459 ( .A1(n16023), .A2(n19754), .ZN(n16002) );
  AOI211_X1 U19460 ( .C1(BUF1_REG_21__SCAN_IN), .C2(n16932), .A(n16003), .B(
        n16002), .ZN(n16005) );
  NAND2_X1 U19461 ( .A1(n16933), .A2(BUF2_REG_21__SCAN_IN), .ZN(n16004) );
  OAI211_X1 U19462 ( .C1(n16917), .C2(n19982), .A(n16005), .B(n16004), .ZN(
        P2_U2898) );
  INV_X1 U19463 ( .A(BUF2_REG_20__SCAN_IN), .ZN(n16014) );
  NAND2_X1 U19464 ( .A1(n16006), .A2(n16936), .ZN(n16013) );
  OAI22_X1 U19465 ( .A1(n16930), .A2(n20105), .B1(n16020), .B2(n16007), .ZN(
        n16011) );
  AND2_X1 U19466 ( .A1(n16021), .A2(n16008), .ZN(n16009) );
  NOR2_X1 U19467 ( .A1(n16000), .A2(n16009), .ZN(n16294) );
  INV_X1 U19468 ( .A(n16294), .ZN(n19761) );
  NOR2_X1 U19469 ( .A1(n19761), .A2(n16023), .ZN(n16010) );
  AOI211_X1 U19470 ( .C1(BUF1_REG_20__SCAN_IN), .C2(n16932), .A(n16011), .B(
        n16010), .ZN(n16012) );
  OAI211_X1 U19471 ( .C1(n16015), .C2(n16014), .A(n16013), .B(n16012), .ZN(
        P2_U2899) );
  NAND2_X1 U19472 ( .A1(n16017), .A2(n16016), .ZN(n16018) );
  NAND2_X1 U19473 ( .A1(n14481), .A2(n16018), .ZN(n16921) );
  OAI22_X1 U19474 ( .A1(n16930), .A2(n20099), .B1(n16020), .B2(n16019), .ZN(
        n16025) );
  OAI21_X1 U19475 ( .B1(n14579), .B2(n16022), .A(n16021), .ZN(n19779) );
  NOR2_X1 U19476 ( .A1(n16023), .A2(n19779), .ZN(n16024) );
  AOI211_X1 U19477 ( .C1(BUF1_REG_19__SCAN_IN), .C2(n16932), .A(n16025), .B(
        n16024), .ZN(n16027) );
  NAND2_X1 U19478 ( .A1(n16933), .A2(BUF2_REG_19__SCAN_IN), .ZN(n16026) );
  OAI211_X1 U19479 ( .C1(n16921), .C2(n19982), .A(n16027), .B(n16026), .ZN(
        P2_U2900) );
  INV_X1 U19480 ( .A(n16028), .ZN(n16029) );
  NOR2_X1 U19481 ( .A1(n16030), .A2(n16029), .ZN(n16031) );
  XNOR2_X1 U19482 ( .A(n16032), .B(n16031), .ZN(n16218) );
  AOI21_X1 U19483 ( .B1(n16206), .B2(n16034), .A(n16033), .ZN(n16216) );
  NAND2_X1 U19484 ( .A1(n19905), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n16210) );
  OAI21_X1 U19485 ( .B1(n20055), .B2(n16035), .A(n16210), .ZN(n16036) );
  AOI21_X1 U19486 ( .B1(n17008), .B2(n16037), .A(n16036), .ZN(n16038) );
  OAI21_X1 U19487 ( .B1(n16856), .B2(n16202), .A(n16038), .ZN(n16039) );
  AOI21_X1 U19488 ( .B1(n16216), .B2(n17010), .A(n16039), .ZN(n16040) );
  OAI21_X1 U19489 ( .B1(n16218), .B2(n16974), .A(n16040), .ZN(P2_U2985) );
  INV_X1 U19490 ( .A(n16051), .ZN(n16042) );
  OAI21_X1 U19491 ( .B1(n16041), .B2(n16050), .A(n16042), .ZN(n16043) );
  XOR2_X1 U19492 ( .A(n16044), .B(n16043), .Z(n16230) );
  AOI21_X1 U19493 ( .B1(n16222), .B2(n16045), .A(n9790), .ZN(n16227) );
  NOR2_X1 U19494 ( .A1(n12009), .A2(n20672), .ZN(n16221) );
  NOR2_X1 U19495 ( .A1(n20045), .A2(n16895), .ZN(n16046) );
  AOI211_X1 U19496 ( .C1(n20029), .C2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n16221), .B(n16046), .ZN(n16047) );
  OAI21_X1 U19497 ( .B1(n16890), .B2(n16202), .A(n16047), .ZN(n16048) );
  AOI21_X1 U19498 ( .B1(n16227), .B2(n17010), .A(n16048), .ZN(n16049) );
  OAI21_X1 U19499 ( .B1(n16230), .B2(n16974), .A(n16049), .ZN(P2_U2988) );
  NOR2_X1 U19500 ( .A1(n16051), .A2(n16050), .ZN(n16052) );
  XOR2_X1 U19501 ( .A(n16052), .B(n16041), .Z(n16242) );
  INV_X1 U19502 ( .A(n16045), .ZN(n16054) );
  AOI21_X1 U19503 ( .B1(n10192), .B2(n16053), .A(n16054), .ZN(n16231) );
  NOR2_X1 U19504 ( .A1(n12009), .A2(n20670), .ZN(n16232) );
  NOR2_X1 U19505 ( .A1(n20045), .A2(n16055), .ZN(n16056) );
  AOI211_X1 U19506 ( .C1(n20029), .C2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n16232), .B(n16056), .ZN(n16057) );
  OAI21_X1 U19507 ( .B1(n16237), .B2(n16202), .A(n16057), .ZN(n16058) );
  AOI21_X1 U19508 ( .B1(n16231), .B2(n17010), .A(n16058), .ZN(n16059) );
  OAI21_X1 U19509 ( .B1(n16974), .B2(n16242), .A(n16059), .ZN(P2_U2989) );
  INV_X1 U19510 ( .A(n16061), .ZN(n16062) );
  NOR2_X1 U19511 ( .A1(n16063), .A2(n16062), .ZN(n16064) );
  XNOR2_X1 U19512 ( .A(n16060), .B(n16064), .ZN(n16253) );
  OAI21_X1 U19513 ( .B1(n16065), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n16053), .ZN(n16247) );
  INV_X1 U19514 ( .A(n16247), .ZN(n16073) );
  INV_X1 U19515 ( .A(n16066), .ZN(n16070) );
  NOR2_X1 U19516 ( .A1(n12009), .A2(n20668), .ZN(n16244) );
  INV_X1 U19517 ( .A(n16244), .ZN(n16067) );
  OAI21_X1 U19518 ( .B1(n20055), .B2(n16068), .A(n16067), .ZN(n16069) );
  AOI21_X1 U19519 ( .B1(n17008), .B2(n16070), .A(n16069), .ZN(n16071) );
  OAI21_X1 U19520 ( .B1(n16246), .B2(n16202), .A(n16071), .ZN(n16072) );
  AOI21_X1 U19521 ( .B1(n16073), .B2(n17010), .A(n16072), .ZN(n16074) );
  OAI21_X1 U19522 ( .B1(n16253), .B2(n16974), .A(n16074), .ZN(P2_U2990) );
  NAND2_X1 U19523 ( .A1(n16076), .A2(n16075), .ZN(n16080) );
  NAND2_X1 U19524 ( .A1(n16078), .A2(n16077), .ZN(n16079) );
  XOR2_X1 U19525 ( .A(n16080), .B(n16079), .Z(n16277) );
  AOI21_X1 U19526 ( .B1(n16273), .B2(n14748), .A(n16081), .ZN(n16267) );
  INV_X1 U19527 ( .A(n16467), .ZN(n16084) );
  NAND2_X1 U19528 ( .A1(n19905), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n16270) );
  OAI21_X1 U19529 ( .B1(n20055), .B2(n16082), .A(n16270), .ZN(n16083) );
  AOI21_X1 U19530 ( .B1(n17008), .B2(n16084), .A(n16083), .ZN(n16085) );
  OAI21_X1 U19531 ( .B1(n16463), .B2(n16202), .A(n16085), .ZN(n16086) );
  AOI21_X1 U19532 ( .B1(n16267), .B2(n17010), .A(n16086), .ZN(n16087) );
  OAI21_X1 U19533 ( .B1(n16277), .B2(n16974), .A(n16087), .ZN(P2_U2992) );
  NAND2_X1 U19534 ( .A1(n16088), .A2(n16369), .ZN(n16957) );
  INV_X1 U19535 ( .A(n16959), .ZN(n16089) );
  OAI21_X2 U19536 ( .B1(n16957), .B2(n16089), .A(n16958), .ZN(n16351) );
  INV_X1 U19537 ( .A(n16350), .ZN(n16090) );
  INV_X1 U19538 ( .A(n16942), .ZN(n16091) );
  INV_X1 U19539 ( .A(n16092), .ZN(n16093) );
  INV_X1 U19540 ( .A(n16095), .ZN(n16096) );
  INV_X1 U19541 ( .A(n16097), .ZN(n16098) );
  INV_X1 U19542 ( .A(n16100), .ZN(n16116) );
  NAND2_X1 U19543 ( .A1(n16102), .A2(n16101), .ZN(n16103) );
  XNOR2_X1 U19544 ( .A(n16104), .B(n16103), .ZN(n16288) );
  INV_X1 U19545 ( .A(n14748), .ZN(n16105) );
  AOI21_X1 U19546 ( .B1(n16280), .B2(n16106), .A(n16105), .ZN(n16286) );
  AND2_X1 U19547 ( .A1(n16108), .A2(n16107), .ZN(n16109) );
  OR2_X1 U19548 ( .A1(n16109), .A2(n9819), .ZN(n16920) );
  INV_X1 U19549 ( .A(n19751), .ZN(n16111) );
  NAND2_X1 U19550 ( .A1(n20028), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n16282) );
  OAI21_X1 U19551 ( .B1(n20055), .B2(n10085), .A(n16282), .ZN(n16110) );
  AOI21_X1 U19552 ( .B1(n17008), .B2(n16111), .A(n16110), .ZN(n16112) );
  OAI21_X1 U19553 ( .B1(n16920), .B2(n16202), .A(n16112), .ZN(n16113) );
  AOI21_X1 U19554 ( .B1(n16286), .B2(n17010), .A(n16113), .ZN(n16114) );
  OAI21_X1 U19555 ( .B1(n16288), .B2(n16974), .A(n16114), .ZN(P2_U2993) );
  OAI21_X1 U19556 ( .B1(n16116), .B2(n16118), .A(n16115), .ZN(n16117) );
  OAI21_X1 U19557 ( .B1(n10153), .B2(n16118), .A(n16117), .ZN(n16301) );
  NOR2_X1 U19558 ( .A1(n16119), .A2(n16120), .ZN(n16122) );
  NOR2_X1 U19559 ( .A1(n16122), .A2(n16121), .ZN(n16132) );
  AOI21_X1 U19560 ( .B1(n16297), .B2(n16132), .A(n16123), .ZN(n16299) );
  NOR2_X1 U19561 ( .A1(n12009), .A2(n16124), .ZN(n16293) );
  NOR2_X1 U19562 ( .A1(n20045), .A2(n16125), .ZN(n16126) );
  AOI211_X1 U19563 ( .C1(n20029), .C2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n16293), .B(n16126), .ZN(n16127) );
  OAI21_X1 U19564 ( .B1(n19762), .B2(n16202), .A(n16127), .ZN(n16128) );
  AOI21_X1 U19565 ( .B1(n16299), .B2(n17010), .A(n16128), .ZN(n16129) );
  OAI21_X1 U19566 ( .B1(n16301), .B2(n16974), .A(n16129), .ZN(P2_U2994) );
  NOR2_X1 U19567 ( .A1(n16119), .A2(n16130), .ZN(n16131) );
  OR2_X1 U19568 ( .A1(n16131), .A2(n10219), .ZN(n16151) );
  OAI21_X1 U19569 ( .B1(n16151), .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n16132), .ZN(n16311) );
  INV_X1 U19570 ( .A(n16144), .ZN(n16133) );
  OAI21_X1 U19571 ( .B1(n16146), .B2(n16133), .A(n16145), .ZN(n16136) );
  XNOR2_X1 U19572 ( .A(n16134), .B(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n16135) );
  XNOR2_X1 U19573 ( .A(n16136), .B(n16135), .ZN(n16302) );
  NAND2_X1 U19574 ( .A1(n16302), .A2(n20046), .ZN(n16143) );
  NAND2_X1 U19575 ( .A1(n19905), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n16303) );
  OAI21_X1 U19576 ( .B1(n20055), .B2(n19768), .A(n16303), .ZN(n16141) );
  NAND2_X1 U19577 ( .A1(n14128), .A2(n16137), .ZN(n16138) );
  NAND2_X1 U19578 ( .A1(n16139), .A2(n16138), .ZN(n16924) );
  NOR2_X1 U19579 ( .A1(n16924), .A2(n16202), .ZN(n16140) );
  AOI211_X1 U19580 ( .C1(n17008), .C2(n19773), .A(n16141), .B(n16140), .ZN(
        n16142) );
  OAI211_X1 U19581 ( .C1(n20043), .C2(n16311), .A(n16143), .B(n16142), .ZN(
        P2_U2995) );
  NAND2_X1 U19582 ( .A1(n16145), .A2(n16144), .ZN(n16147) );
  XOR2_X1 U19583 ( .A(n16147), .B(n16146), .Z(n16325) );
  NAND2_X2 U19584 ( .A1(n16187), .A2(n16148), .ZN(n16400) );
  AND2_X1 U19585 ( .A1(n16149), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n16150) );
  NAND2_X2 U19586 ( .A1(n16400), .A2(n16150), .ZN(n16948) );
  INV_X1 U19587 ( .A(n16314), .ZN(n16331) );
  NOR2_X2 U19588 ( .A1(n16948), .A2(n16331), .ZN(n16326) );
  AOI21_X1 U19589 ( .B1(n16326), .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n16152) );
  NOR2_X1 U19590 ( .A1(n16152), .A2(n16151), .ZN(n16323) );
  NOR2_X1 U19591 ( .A1(n12009), .A2(n20658), .ZN(n16312) );
  NOR2_X1 U19592 ( .A1(n19780), .A2(n20045), .ZN(n16153) );
  AOI211_X1 U19593 ( .C1(n20029), .C2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n16312), .B(n16153), .ZN(n16154) );
  OAI21_X1 U19594 ( .B1(n16202), .B2(n19787), .A(n16154), .ZN(n16155) );
  AOI21_X1 U19595 ( .B1(n16323), .B2(n17010), .A(n16155), .ZN(n16156) );
  OAI21_X1 U19596 ( .B1(n16325), .B2(n16974), .A(n16156), .ZN(P2_U2996) );
  XOR2_X1 U19597 ( .A(n16158), .B(n16157), .Z(n16338) );
  XNOR2_X1 U19598 ( .A(n16326), .B(n16159), .ZN(n16167) );
  INV_X1 U19599 ( .A(n19798), .ZN(n16160) );
  OAI22_X1 U19600 ( .A1(n16161), .A2(n20055), .B1(n20045), .B2(n16160), .ZN(
        n16166) );
  NOR2_X1 U19601 ( .A1(n16163), .A2(n16162), .ZN(n16164) );
  OR2_X1 U19602 ( .A1(n14129), .A2(n16164), .ZN(n16929) );
  NAND2_X1 U19603 ( .A1(n19905), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n16332) );
  OAI21_X1 U19604 ( .B1(n16929), .B2(n16202), .A(n16332), .ZN(n16165) );
  AOI211_X1 U19605 ( .C1(n16167), .C2(n17010), .A(n16166), .B(n16165), .ZN(
        n16168) );
  OAI21_X1 U19606 ( .B1(n16338), .B2(n16974), .A(n16168), .ZN(P2_U2997) );
  XNOR2_X1 U19607 ( .A(n16170), .B(n16169), .ZN(n16348) );
  INV_X1 U19608 ( .A(n19810), .ZN(n16174) );
  NOR2_X1 U19609 ( .A1(n20654), .A2(n12009), .ZN(n16173) );
  INV_X1 U19610 ( .A(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n16171) );
  OAI22_X1 U19611 ( .A1(n16171), .A2(n20055), .B1(n20045), .B2(n19804), .ZN(
        n16172) );
  AOI211_X1 U19612 ( .C1(n20051), .C2(n16174), .A(n16173), .B(n16172), .ZN(
        n16178) );
  NOR2_X1 U19613 ( .A1(n16948), .A2(n16340), .ZN(n16176) );
  INV_X1 U19614 ( .A(n16326), .ZN(n16175) );
  OAI211_X1 U19615 ( .C1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .C2(n16176), .A(
        n16175), .B(n17010), .ZN(n16177) );
  OAI211_X1 U19616 ( .C1(n16348), .C2(n16974), .A(n16178), .B(n16177), .ZN(
        P2_U2998) );
  INV_X1 U19617 ( .A(n16195), .ZN(n16180) );
  AOI21_X1 U19618 ( .B1(n16179), .B2(n16194), .A(n16180), .ZN(n16184) );
  NAND2_X1 U19619 ( .A1(n16182), .A2(n16181), .ZN(n16183) );
  XNOR2_X1 U19620 ( .A(n16184), .B(n16183), .ZN(n17056) );
  NAND2_X1 U19621 ( .A1(n16119), .A2(n16185), .ZN(n16186) );
  AND2_X1 U19622 ( .A1(n16187), .A2(n16186), .ZN(n17053) );
  OAI22_X1 U19623 ( .A1(n10945), .A2(n20073), .B1(n20045), .B2(n16188), .ZN(
        n16192) );
  INV_X1 U19624 ( .A(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n16189) );
  OAI22_X1 U19625 ( .A1(n16190), .A2(n16202), .B1(n20055), .B2(n16189), .ZN(
        n16191) );
  AOI211_X1 U19626 ( .C1(n17053), .C2(n17010), .A(n16192), .B(n16191), .ZN(
        n16193) );
  OAI21_X1 U19627 ( .B1(n17056), .B2(n16974), .A(n16193), .ZN(P2_U3006) );
  NAND2_X1 U19628 ( .A1(n16195), .A2(n16194), .ZN(n16196) );
  XOR2_X1 U19629 ( .A(n16196), .B(n16179), .Z(n16422) );
  XNOR2_X1 U19630 ( .A(n16198), .B(n10936), .ZN(n16199) );
  XNOR2_X1 U19631 ( .A(n16197), .B(n16199), .ZN(n16420) );
  OAI22_X1 U19632 ( .A1(n16200), .A2(n20055), .B1(n10940), .B2(n20073), .ZN(
        n16204) );
  INV_X1 U19633 ( .A(n19875), .ZN(n16201) );
  OAI22_X1 U19634 ( .A1(n16202), .A2(n19881), .B1(n20045), .B2(n16201), .ZN(
        n16203) );
  AOI211_X1 U19635 ( .C1(n16420), .C2(n17010), .A(n16204), .B(n16203), .ZN(
        n16205) );
  OAI21_X1 U19636 ( .B1(n16422), .B2(n16974), .A(n16205), .ZN(P2_U3007) );
  AOI21_X1 U19637 ( .B1(n16208), .B2(n16207), .A(n16206), .ZN(n16215) );
  INV_X1 U19638 ( .A(n16209), .ZN(n16211) );
  OAI21_X1 U19639 ( .B1(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n16211), .A(
        n16210), .ZN(n16212) );
  AOI21_X1 U19640 ( .B1(n16857), .B2(n20057), .A(n16212), .ZN(n16213) );
  OAI21_X1 U19641 ( .B1(n16856), .B2(n20062), .A(n16213), .ZN(n16214) );
  OAI21_X1 U19642 ( .B1(n16218), .B2(n17071), .A(n16217), .ZN(P2_U3017) );
  AOI21_X1 U19643 ( .B1(n16222), .B2(n10192), .A(n16219), .ZN(n16226) );
  INV_X1 U19644 ( .A(n16220), .ZN(n16891) );
  AOI21_X1 U19645 ( .B1(n16891), .B2(n20057), .A(n16221), .ZN(n16224) );
  OR2_X1 U19646 ( .A1(n16234), .A2(n16222), .ZN(n16223) );
  OAI211_X1 U19647 ( .C1(n16890), .C2(n20062), .A(n16224), .B(n16223), .ZN(
        n16225) );
  AOI21_X1 U19648 ( .B1(n16239), .B2(n16226), .A(n16225), .ZN(n16229) );
  NAND2_X1 U19649 ( .A1(n16227), .A2(n17052), .ZN(n16228) );
  OAI211_X1 U19650 ( .C1(n16230), .C2(n17071), .A(n16229), .B(n16228), .ZN(
        P2_U3020) );
  NAND2_X1 U19651 ( .A1(n16231), .A2(n17052), .ZN(n16241) );
  AOI21_X1 U19652 ( .B1(n16233), .B2(n20057), .A(n16232), .ZN(n16236) );
  OR2_X1 U19653 ( .A1(n16234), .A2(n10192), .ZN(n16235) );
  OAI211_X1 U19654 ( .C1(n16237), .C2(n20062), .A(n16236), .B(n16235), .ZN(
        n16238) );
  AOI21_X1 U19655 ( .B1(n16239), .B2(n10192), .A(n16238), .ZN(n16240) );
  OAI211_X1 U19656 ( .C1(n16242), .C2(n17071), .A(n16241), .B(n16240), .ZN(
        P2_U3021) );
  OAI21_X1 U19657 ( .B1(n16261), .B2(n16262), .A(n16243), .ZN(n16250) );
  AOI21_X1 U19658 ( .B1(n16934), .B2(n20057), .A(n16244), .ZN(n16245) );
  OAI21_X1 U19659 ( .B1(n16246), .B2(n20062), .A(n16245), .ZN(n16249) );
  NOR2_X1 U19660 ( .A1(n16247), .A2(n20068), .ZN(n16248) );
  AOI211_X1 U19661 ( .C1(n16251), .C2(n16250), .A(n16249), .B(n16248), .ZN(
        n16252) );
  OAI21_X1 U19662 ( .B1(n16253), .B2(n17071), .A(n16252), .ZN(P2_U3022) );
  OR2_X1 U19663 ( .A1(n16254), .A2(n20068), .ZN(n16266) );
  NAND2_X1 U19664 ( .A1(n16902), .A2(n17074), .ZN(n16257) );
  AOI21_X1 U19665 ( .B1(n16901), .B2(n20057), .A(n16255), .ZN(n16256) );
  OAI211_X1 U19666 ( .C1(n16268), .C2(n16258), .A(n16257), .B(n16256), .ZN(
        n16259) );
  INV_X1 U19667 ( .A(n16259), .ZN(n16265) );
  NAND3_X1 U19668 ( .A1(n16260), .A2(n14757), .A3(n20059), .ZN(n16264) );
  INV_X1 U19669 ( .A(n16261), .ZN(n16274) );
  OAI211_X1 U19670 ( .C1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(n16274), .B(n16262), .ZN(
        n16263) );
  NAND4_X1 U19671 ( .A1(n16266), .A2(n16265), .A3(n16264), .A4(n16263), .ZN(
        P2_U3023) );
  NAND2_X1 U19672 ( .A1(n16267), .A2(n17052), .ZN(n16276) );
  NOR2_X1 U19673 ( .A1(n16268), .A2(n16273), .ZN(n16272) );
  NAND2_X1 U19674 ( .A1(n20057), .A2(n16461), .ZN(n16269) );
  OAI211_X1 U19675 ( .C1(n16463), .C2(n20062), .A(n16270), .B(n16269), .ZN(
        n16271) );
  AOI211_X1 U19676 ( .C1(n16274), .C2(n16273), .A(n16272), .B(n16271), .ZN(
        n16275) );
  OAI211_X1 U19677 ( .C1(n16277), .C2(n17071), .A(n16276), .B(n16275), .ZN(
        P2_U3024) );
  INV_X1 U19678 ( .A(n16278), .ZN(n16279) );
  AOI21_X1 U19679 ( .B1(n16281), .B2(n16280), .A(n16279), .ZN(n16285) );
  INV_X1 U19680 ( .A(n16920), .ZN(n19745) );
  NAND2_X1 U19681 ( .A1(n19745), .A2(n17074), .ZN(n16283) );
  OAI211_X1 U19682 ( .C1(n17048), .C2(n19754), .A(n16283), .B(n16282), .ZN(
        n16284) );
  AOI211_X1 U19683 ( .C1(n16286), .C2(n17052), .A(n16285), .B(n16284), .ZN(
        n16287) );
  OAI21_X1 U19684 ( .B1(n16288), .B2(n17071), .A(n16287), .ZN(P2_U3025) );
  AOI21_X1 U19685 ( .B1(n16290), .B2(n16289), .A(n17019), .ZN(n16321) );
  OAI211_X1 U19686 ( .C1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(n16308), .B(n16291), .ZN(
        n16296) );
  NOR2_X1 U19687 ( .A1(n19762), .A2(n20062), .ZN(n16292) );
  AOI211_X1 U19688 ( .C1(n20057), .C2(n16294), .A(n16293), .B(n16292), .ZN(
        n16295) );
  OAI211_X1 U19689 ( .C1(n16321), .C2(n16297), .A(n16296), .B(n16295), .ZN(
        n16298) );
  AOI21_X1 U19690 ( .B1(n16299), .B2(n17052), .A(n16298), .ZN(n16300) );
  OAI21_X1 U19691 ( .B1(n16301), .B2(n17071), .A(n16300), .ZN(P2_U3026) );
  NAND2_X1 U19692 ( .A1(n16302), .A2(n20059), .ZN(n16310) );
  INV_X1 U19693 ( .A(n16924), .ZN(n19775) );
  OAI21_X1 U19694 ( .B1(n17048), .B2(n19779), .A(n16303), .ZN(n16304) );
  AOI21_X1 U19695 ( .B1(n19775), .B2(n17074), .A(n16304), .ZN(n16305) );
  OAI21_X1 U19696 ( .B1(n16321), .B2(n16307), .A(n16305), .ZN(n16306) );
  AOI21_X1 U19697 ( .B1(n16308), .B2(n16307), .A(n16306), .ZN(n16309) );
  OAI211_X1 U19698 ( .C1(n16311), .C2(n20068), .A(n16310), .B(n16309), .ZN(
        P2_U3027) );
  INV_X1 U19699 ( .A(n16312), .ZN(n16316) );
  NOR2_X1 U19700 ( .A1(n16407), .A2(n16408), .ZN(n16357) );
  INV_X1 U19701 ( .A(n16357), .ZN(n17034) );
  NOR2_X1 U19702 ( .A1(n16313), .A2(n17034), .ZN(n17015) );
  NAND4_X1 U19703 ( .A1(n17015), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A3(
        n16314), .A4(n16320), .ZN(n16315) );
  OAI211_X1 U19704 ( .C1(n19787), .C2(n20062), .A(n16316), .B(n16315), .ZN(
        n16317) );
  AOI21_X1 U19705 ( .B1(n20057), .B2(n16318), .A(n16317), .ZN(n16319) );
  OAI21_X1 U19706 ( .B1(n16321), .B2(n16320), .A(n16319), .ZN(n16322) );
  AOI21_X1 U19707 ( .B1(n16323), .B2(n17052), .A(n16322), .ZN(n16324) );
  OAI21_X1 U19708 ( .B1(n16325), .B2(n17071), .A(n16324), .ZN(P2_U3028) );
  AOI21_X1 U19709 ( .B1(n20068), .B2(n16327), .A(n16326), .ZN(n16328) );
  AOI211_X1 U19710 ( .C1(n16329), .C2(n16340), .A(n17019), .B(n16328), .ZN(
        n16339) );
  OAI21_X1 U19711 ( .B1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n17077), .A(
        n16339), .ZN(n16336) );
  INV_X1 U19712 ( .A(n16948), .ZN(n16330) );
  AOI21_X1 U19713 ( .B1(n16330), .B2(n17052), .A(n17015), .ZN(n16341) );
  NOR3_X1 U19714 ( .A1(n16341), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A3(
        n16331), .ZN(n16335) );
  INV_X1 U19715 ( .A(n16929), .ZN(n19799) );
  NAND2_X1 U19716 ( .A1(n19799), .A2(n17074), .ZN(n16333) );
  OAI211_X1 U19717 ( .C1(n17048), .C2(n19802), .A(n16333), .B(n16332), .ZN(
        n16334) );
  AOI211_X1 U19718 ( .C1(n16336), .C2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n16335), .B(n16334), .ZN(n16337) );
  OAI21_X1 U19719 ( .B1(n16338), .B2(n17071), .A(n16337), .ZN(P2_U3029) );
  INV_X1 U19720 ( .A(n16339), .ZN(n16346) );
  NOR3_X1 U19721 ( .A1(n16341), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        n16340), .ZN(n16345) );
  AOI22_X1 U19722 ( .A1(n20057), .A2(n16342), .B1(P2_REIP_REG_16__SCAN_IN), 
        .B2(n20028), .ZN(n16343) );
  OAI21_X1 U19723 ( .B1(n19810), .B2(n20062), .A(n16343), .ZN(n16344) );
  AOI211_X1 U19724 ( .C1(n16346), .C2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n16345), .B(n16344), .ZN(n16347) );
  OAI21_X1 U19725 ( .B1(n17071), .B2(n16348), .A(n16347), .ZN(P2_U3030) );
  NAND2_X1 U19726 ( .A1(n16350), .A2(n16349), .ZN(n16352) );
  XOR2_X1 U19727 ( .A(n16352), .B(n16351), .Z(n16953) );
  NAND2_X2 U19728 ( .A1(n16987), .A2(n16386), .ZN(n16384) );
  NOR2_X2 U19729 ( .A1(n16384), .A2(n16373), .ZN(n16961) );
  NAND2_X1 U19730 ( .A1(n16961), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n16963) );
  NAND2_X1 U19731 ( .A1(n16963), .A2(n16353), .ZN(n16354) );
  NAND2_X1 U19732 ( .A1(n16354), .A2(n16948), .ZN(n16952) );
  AOI21_X1 U19733 ( .B1(n16355), .B2(n13574), .A(n13827), .ZN(n19834) );
  INV_X1 U19734 ( .A(n19834), .ZN(n19973) );
  OAI22_X1 U19735 ( .A1(n17048), .A2(n19973), .B1(n10967), .B2(n20073), .ZN(
        n16356) );
  AOI21_X1 U19736 ( .B1(n17074), .B2(n19835), .A(n16356), .ZN(n16364) );
  NAND2_X1 U19737 ( .A1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16359) );
  NAND2_X1 U19738 ( .A1(n16386), .A2(n16357), .ZN(n16358) );
  NOR2_X1 U19739 ( .A1(n16359), .A2(n16358), .ZN(n16361) );
  INV_X1 U19740 ( .A(n16358), .ZN(n17024) );
  OAI21_X1 U19741 ( .B1(n16386), .B2(n17077), .A(n17033), .ZN(n16372) );
  AOI21_X1 U19742 ( .B1(n17024), .B2(n16359), .A(n16372), .ZN(n17026) );
  INV_X1 U19743 ( .A(n17026), .ZN(n16360) );
  MUX2_X1 U19744 ( .A(n16361), .B(n16360), .S(
        P2_INSTADDRPOINTER_REG_14__SCAN_IN), .Z(n16362) );
  INV_X1 U19745 ( .A(n16362), .ZN(n16363) );
  OAI211_X1 U19746 ( .C1(n16952), .C2(n20068), .A(n16364), .B(n16363), .ZN(
        n16365) );
  INV_X1 U19747 ( .A(n16365), .ZN(n16366) );
  OAI21_X1 U19748 ( .B1(n16953), .B2(n17071), .A(n16366), .ZN(P2_U3032) );
  NAND2_X1 U19749 ( .A1(n16369), .A2(n16368), .ZN(n16370) );
  XNOR2_X1 U19750 ( .A(n16367), .B(n16370), .ZN(n16973) );
  AOI21_X1 U19751 ( .B1(n16373), .B2(n16384), .A(n16961), .ZN(n16972) );
  NOR2_X1 U19752 ( .A1(n10962), .A2(n20073), .ZN(n16371) );
  AOI221_X1 U19753 ( .B1(n17024), .B2(n16373), .C1(n16372), .C2(
        P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A(n16371), .ZN(n16375) );
  NAND2_X1 U19754 ( .A1(n17074), .A2(n19856), .ZN(n16374) );
  OAI211_X1 U19755 ( .C1(n17048), .C2(n19857), .A(n16375), .B(n16374), .ZN(
        n16376) );
  AOI21_X1 U19756 ( .B1(n16972), .B2(n17052), .A(n16376), .ZN(n16377) );
  OAI21_X1 U19757 ( .B1(n17071), .B2(n16973), .A(n16377), .ZN(P2_U3034) );
  INV_X1 U19758 ( .A(n16379), .ZN(n16380) );
  OR2_X1 U19759 ( .A1(n16381), .A2(n16380), .ZN(n16382) );
  XNOR2_X1 U19760 ( .A(n16378), .B(n16382), .ZN(n16979) );
  INV_X1 U19761 ( .A(n16979), .ZN(n16398) );
  NAND2_X1 U19762 ( .A1(n16987), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n16383) );
  NAND2_X1 U19763 ( .A1(n16383), .A2(n16393), .ZN(n16385) );
  NAND2_X1 U19764 ( .A1(n16385), .A2(n16384), .ZN(n16982) );
  INV_X1 U19765 ( .A(n16982), .ZN(n16396) );
  AOI211_X1 U19766 ( .C1(n10722), .C2(n16393), .A(n16386), .B(n17034), .ZN(
        n16395) );
  OAI22_X1 U19767 ( .A1(n17048), .A2(n19873), .B1(n20648), .B2(n20073), .ZN(
        n16391) );
  NOR2_X1 U19768 ( .A1(n16387), .A2(n14241), .ZN(n16388) );
  NOR2_X1 U19769 ( .A1(n13640), .A2(n16388), .ZN(n19954) );
  INV_X1 U19770 ( .A(n19954), .ZN(n16389) );
  NOR2_X1 U19771 ( .A1(n20062), .A2(n16389), .ZN(n16390) );
  NOR2_X1 U19772 ( .A1(n16391), .A2(n16390), .ZN(n16392) );
  OAI21_X1 U19773 ( .B1(n17033), .B2(n16393), .A(n16392), .ZN(n16394) );
  AOI211_X1 U19774 ( .C1(n16396), .C2(n17052), .A(n16395), .B(n16394), .ZN(
        n16397) );
  OAI21_X1 U19775 ( .B1(n16398), .B2(n17071), .A(n16397), .ZN(P2_U3035) );
  INV_X1 U19776 ( .A(n16987), .ZN(n16399) );
  OAI21_X1 U19777 ( .B1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n16400), .A(
        n16399), .ZN(n17001) );
  INV_X1 U19778 ( .A(n16401), .ZN(n16405) );
  AOI21_X1 U19779 ( .B1(n16403), .B2(n16988), .A(n16402), .ZN(n16404) );
  AOI21_X1 U19780 ( .B1(n16405), .B2(n16988), .A(n16404), .ZN(n17003) );
  NAND2_X1 U19781 ( .A1(P2_REIP_REG_9__SCAN_IN), .A2(n19905), .ZN(n16406) );
  OAI221_X1 U19782 ( .B1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n16408), .C1(
        n16407), .C2(n17033), .A(n16406), .ZN(n16411) );
  OAI22_X1 U19783 ( .A1(n16409), .A2(n17048), .B1(n20062), .B2(n17002), .ZN(
        n16410) );
  AOI211_X1 U19784 ( .C1(n17003), .C2(n20059), .A(n16411), .B(n16410), .ZN(
        n16412) );
  OAI21_X1 U19785 ( .B1(n20068), .B2(n17001), .A(n16412), .ZN(P2_U3037) );
  AOI21_X1 U19786 ( .B1(n17066), .B2(n16415), .A(n16413), .ZN(n17043) );
  AND3_X1 U19787 ( .A1(n10936), .A2(n16415), .A3(n16414), .ZN(n17044) );
  NOR2_X1 U19788 ( .A1(n10940), .A2(n20073), .ZN(n16416) );
  AOI211_X1 U19789 ( .C1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .C2(n17043), .A(
        n17044), .B(n16416), .ZN(n16417) );
  INV_X1 U19790 ( .A(n16417), .ZN(n16419) );
  OAI22_X1 U19791 ( .A1(n19882), .A2(n17048), .B1(n20062), .B2(n19881), .ZN(
        n16418) );
  AOI211_X1 U19792 ( .C1(n16420), .C2(n17052), .A(n16419), .B(n16418), .ZN(
        n16421) );
  OAI21_X1 U19793 ( .B1(n16422), .B2(n17071), .A(n16421), .ZN(P2_U3039) );
  OAI21_X1 U19794 ( .B1(n9719), .B2(n16424), .A(n16423), .ZN(n16432) );
  INV_X1 U19795 ( .A(n16432), .ZN(n16426) );
  AND2_X1 U19796 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n16425), .ZN(n16431) );
  AOI222_X1 U19797 ( .A1(n16427), .A2(n16433), .B1(n20718), .B2(n17082), .C1(
        n16426), .C2(n16431), .ZN(n16429) );
  NAND2_X1 U19798 ( .A1(n16439), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n16428) );
  OAI21_X1 U19799 ( .B1(n16429), .B2(n16439), .A(n16428), .ZN(P2_U3600) );
  AOI222_X1 U19800 ( .A1(n16434), .A2(n16433), .B1(n16432), .B2(n16431), .C1(
        n16430), .C2(n17082), .ZN(n16436) );
  NAND2_X1 U19801 ( .A1(n16439), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n16435) );
  OAI21_X1 U19802 ( .B1(n16436), .B2(n16439), .A(n16435), .ZN(P2_U3599) );
  INV_X1 U19803 ( .A(n17082), .ZN(n16438) );
  OAI22_X1 U19804 ( .A1(n20131), .A2(n16438), .B1(n16437), .B2(n20696), .ZN(
        n16440) );
  MUX2_X1 U19805 ( .A(n16440), .B(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n16439), .Z(P2_U3596) );
  AOI22_X1 U19806 ( .A1(n17948), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n9714), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n16441) );
  OAI21_X1 U19807 ( .B1(n17827), .B2(n17789), .A(n16441), .ZN(n16451) );
  AOI22_X1 U19808 ( .A1(n17992), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n18002), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n16449) );
  INV_X1 U19809 ( .A(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n16442) );
  OAI22_X1 U19810 ( .A1(n17788), .A2(n12867), .B1(n10201), .B2(n16442), .ZN(
        n16447) );
  AOI22_X1 U19811 ( .A1(P3_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n12839), .B1(
        n12899), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n16445) );
  AOI22_X1 U19812 ( .A1(n17972), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n9740), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n16444) );
  AOI22_X1 U19813 ( .A1(n17979), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n12840), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n16443) );
  NAND3_X1 U19814 ( .A1(n16445), .A2(n16444), .A3(n16443), .ZN(n16446) );
  AOI211_X1 U19815 ( .C1(n17967), .C2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A(
        n16447), .B(n16446), .ZN(n16448) );
  OAI211_X1 U19816 ( .C1(n17799), .C2(n17913), .A(n16449), .B(n16448), .ZN(
        n16450) );
  AOI211_X1 U19817 ( .C1(n17989), .C2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A(
        n16451), .B(n16450), .ZN(n18148) );
  INV_X1 U19818 ( .A(n16452), .ZN(n16453) );
  NAND3_X1 U19819 ( .A1(n19052), .A2(n19068), .A3(n16453), .ZN(n16454) );
  INV_X1 U19820 ( .A(P3_EBX_REG_10__SCAN_IN), .ZN(n17962) );
  INV_X1 U19821 ( .A(P3_EBX_REG_6__SCAN_IN), .ZN(n18019) );
  INV_X1 U19822 ( .A(P3_EBX_REG_2__SCAN_IN), .ZN(n17605) );
  NAND2_X1 U19823 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n18034) );
  NOR2_X1 U19824 ( .A1(n17605), .A2(n18034), .ZN(n18025) );
  NAND3_X1 U19825 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(P3_EBX_REG_3__SCAN_IN), 
        .A3(n18025), .ZN(n18024) );
  NOR4_X1 U19826 ( .A1(n18012), .A2(n18019), .A3(n18011), .A4(n18024), .ZN(
        n18007) );
  NAND2_X1 U19827 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n18007), .ZN(n18006) );
  NOR2_X1 U19828 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(n17927), .ZN(n16457) );
  NAND2_X1 U19829 ( .A1(n18039), .A2(n17905), .ZN(n17908) );
  OAI22_X1 U19830 ( .A1(n18148), .A2(n18039), .B1(n16457), .B2(n17908), .ZN(
        P3_U2690) );
  AOI22_X1 U19831 ( .A1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n19929), .B1(
        P2_REIP_REG_22__SCAN_IN), .B2(n19927), .ZN(n16471) );
  INV_X1 U19832 ( .A(P2_EBX_REG_22__SCAN_IN), .ZN(n16458) );
  OAI22_X1 U19833 ( .A1(n16459), .A2(n19919), .B1(n19888), .B2(n16458), .ZN(
        n16460) );
  INV_X1 U19834 ( .A(n16460), .ZN(n16470) );
  INV_X1 U19835 ( .A(n16461), .ZN(n16462) );
  OAI22_X1 U19836 ( .A1(n16463), .A2(n19880), .B1(n16462), .B2(n19914), .ZN(
        n16464) );
  INV_X1 U19837 ( .A(n16464), .ZN(n16469) );
  OAI211_X1 U19838 ( .C1(n16467), .C2(n16466), .A(n19897), .B(n16465), .ZN(
        n16468) );
  NAND4_X1 U19839 ( .A1(n16471), .A2(n16470), .A3(n16469), .A4(n16468), .ZN(
        P2_U2833) );
  INV_X1 U19840 ( .A(n16472), .ZN(n16482) );
  AOI21_X1 U19841 ( .B1(n9997), .B2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n21110), .ZN(n16473) );
  AND2_X1 U19842 ( .A1(n16474), .A2(n16473), .ZN(n16478) );
  INV_X1 U19843 ( .A(n16478), .ZN(n16480) );
  INV_X1 U19844 ( .A(n16475), .ZN(n16477) );
  OAI22_X1 U19845 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n16478), .B1(
        n16477), .B2(n16476), .ZN(n16479) );
  OAI21_X1 U19846 ( .B1(n16480), .B2(n21009), .A(n16479), .ZN(n16481) );
  AOI222_X1 U19847 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n16482), 
        .B1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n16481), .C1(n16482), 
        .C2(n16481), .ZN(n16483) );
  OR2_X1 U19848 ( .A1(n16484), .A2(n16483), .ZN(n16485) );
  AOI22_X1 U19849 ( .A1(n16485), .A2(n21010), .B1(n16484), .B2(n16483), .ZN(
        n16491) );
  NOR2_X1 U19850 ( .A1(n16487), .A2(n16486), .ZN(n16490) );
  OAI21_X1 U19851 ( .B1(P1_FLUSH_REG_SCAN_IN), .B2(P1_MORE_REG_SCAN_IN), .A(
        n16488), .ZN(n16489) );
  OAI211_X1 U19852 ( .C1(n16491), .C2(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A(
        n16490), .B(n16489), .ZN(n16492) );
  NOR3_X1 U19853 ( .A1(n16494), .A2(n16493), .A3(n16492), .ZN(n16507) );
  INV_X1 U19854 ( .A(n16507), .ZN(n16497) );
  NAND2_X1 U19855 ( .A1(n16495), .A2(n21118), .ZN(n21289) );
  AOI21_X1 U19856 ( .B1(P1_STATE2_REG_0__SCAN_IN), .B2(
        P1_STATE2_REG_1__SCAN_IN), .A(n21113), .ZN(n21176) );
  NAND2_X1 U19857 ( .A1(n21287), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n16830) );
  OAI211_X1 U19858 ( .C1(n16496), .C2(n21289), .A(n21176), .B(n16830), .ZN(
        n16834) );
  AOI221_X1 U19859 ( .B1(n9954), .B2(n16839), .C1(n16497), .C2(n16839), .A(
        n16834), .ZN(n16840) );
  INV_X1 U19860 ( .A(n21291), .ZN(n16837) );
  NOR2_X1 U19861 ( .A1(n16837), .A2(n16498), .ZN(n16499) );
  NOR2_X1 U19862 ( .A1(n16840), .A2(n16499), .ZN(n16505) );
  INV_X1 U19863 ( .A(n16500), .ZN(n16501) );
  AOI211_X1 U19864 ( .C1(n21190), .C2(n21113), .A(n16502), .B(n16501), .ZN(
        n16503) );
  NAND2_X1 U19865 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n16503), .ZN(n16504) );
  OAI22_X1 U19866 ( .A1(n16505), .A2(P1_STATE2_REG_0__SCAN_IN), .B1(n16840), 
        .B2(n16504), .ZN(n16506) );
  OAI21_X1 U19867 ( .B1(n16507), .B2(n20767), .A(n16506), .ZN(P1_U3161) );
  INV_X1 U19868 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n17140) );
  INV_X1 U19869 ( .A(n19013), .ZN(n18866) );
  NOR2_X1 U19870 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16509), .ZN(
        n17115) );
  AOI22_X1 U19871 ( .A1(n18866), .A2(P3_REIP_REG_30__SCAN_IN), .B1(n17115), 
        .B2(n16510), .ZN(n16514) );
  AOI221_X1 U19872 ( .B1(n18931), .B2(n16511), .C1(n17138), .C2(n16511), .A(
        n18866), .ZN(n17143) );
  OAI21_X1 U19873 ( .B1(n17143), .B2(n16512), .A(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n16513) );
  OAI211_X1 U19874 ( .C1(n17119), .C2(n18877), .A(n16514), .B(n16513), .ZN(
        P3_U2832) );
  INV_X1 U19875 ( .A(HOLD), .ZN(n21186) );
  INV_X1 U19876 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n21197) );
  NAND2_X1 U19877 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(
        P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n21181) );
  OAI21_X1 U19878 ( .B1(n21186), .B2(n21180), .A(n21181), .ZN(n16515) );
  OAI21_X1 U19879 ( .B1(n21186), .B2(n21197), .A(n16515), .ZN(n16517) );
  NOR2_X1 U19880 ( .A1(n21180), .A2(n21287), .ZN(n21189) );
  INV_X1 U19881 ( .A(n21189), .ZN(n21179) );
  NAND3_X1 U19882 ( .A1(n16517), .A2(n16516), .A3(n21179), .ZN(P1_U3195) );
  INV_X1 U19883 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n17257) );
  NOR2_X1 U19884 ( .A1(n20864), .A2(n17257), .ZN(P1_U2905) );
  NOR3_X1 U19885 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(P2_STATEBS16_REG_SCAN_IN), .ZN(n16519) );
  NOR2_X1 U19886 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n16518) );
  NAND2_X1 U19887 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n20607), .ZN(n20610) );
  NOR2_X1 U19888 ( .A1(n20748), .A2(n20610), .ZN(n17079) );
  NOR4_X1 U19889 ( .A1(n16519), .A2(n16518), .A3(n17079), .A4(n17080), .ZN(
        P2_U3178) );
  INV_X1 U19890 ( .A(n17081), .ZN(n20736) );
  AOI221_X1 U19891 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(n17080), .C1(n20736), .C2(
        n17080), .A(n20512), .ZN(n20730) );
  INV_X1 U19892 ( .A(n20730), .ZN(n20731) );
  NOR2_X1 U19893 ( .A1(n16520), .A2(n20731), .ZN(P2_U3047) );
  NAND2_X1 U19894 ( .A1(n19068), .A2(n18049), .ZN(n18198) );
  INV_X1 U19895 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n18270) );
  INV_X1 U19896 ( .A(n18195), .ZN(n18197) );
  NAND2_X1 U19897 ( .A1(n19516), .A2(n18049), .ZN(n18192) );
  AOI22_X1 U19898 ( .A1(n18197), .A2(BUF2_REG_0__SCAN_IN), .B1(n18196), .B2(
        n18683), .ZN(n16525) );
  OAI221_X1 U19899 ( .B1(P3_EAX_REG_0__SCAN_IN), .B2(n18198), .C1(n18270), 
        .C2(n18049), .A(n16525), .ZN(P3_U2735) );
  AOI22_X1 U19900 ( .A1(n20850), .A2(P1_EBX_REG_25__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n20849), .ZN(n16531) );
  INV_X1 U19901 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n21241) );
  OAI22_X1 U19902 ( .A1(n16653), .A2(n20847), .B1(n21241), .B2(n16547), .ZN(
        n16526) );
  INV_X1 U19903 ( .A(n16526), .ZN(n16530) );
  AOI22_X1 U19904 ( .A1(n16650), .A2(n20808), .B1(n16745), .B2(n16609), .ZN(
        n16529) );
  OAI211_X1 U19905 ( .C1(P1_REIP_REG_24__SCAN_IN), .C2(P1_REIP_REG_25__SCAN_IN), .A(n16539), .B(n16527), .ZN(n16528) );
  NAND4_X1 U19906 ( .A1(n16531), .A2(n16530), .A3(n16529), .A4(n16528), .ZN(
        P1_U2815) );
  INV_X1 U19907 ( .A(n16547), .ZN(n16535) );
  AOI22_X1 U19908 ( .A1(n20849), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .B1(
        n16629), .B2(n16532), .ZN(n16533) );
  OAI21_X1 U19909 ( .B1(n16622), .B2(n15487), .A(n16533), .ZN(n16534) );
  AOI21_X1 U19910 ( .B1(n16535), .B2(P1_REIP_REG_24__SCAN_IN), .A(n16534), 
        .ZN(n16536) );
  OAI21_X1 U19911 ( .B1(n16537), .B2(n16617), .A(n16536), .ZN(n16538) );
  AOI21_X1 U19912 ( .B1(n16539), .B2(n21239), .A(n16538), .ZN(n16540) );
  OAI21_X1 U19913 ( .B1(n20860), .B2(n16541), .A(n16540), .ZN(P1_U2816) );
  AOI21_X1 U19914 ( .B1(P1_REIP_REG_22__SCAN_IN), .B2(n16548), .A(
        P1_REIP_REG_23__SCAN_IN), .ZN(n16546) );
  INV_X1 U19915 ( .A(n16660), .ZN(n16542) );
  AOI222_X1 U19916 ( .A1(n16542), .A2(n16629), .B1(n20849), .B2(
        P1_PHYADDRPOINTER_REG_23__SCAN_IN), .C1(n20850), .C2(
        P1_EBX_REG_23__SCAN_IN), .ZN(n16545) );
  NOR2_X1 U19917 ( .A1(n16753), .A2(n20860), .ZN(n16543) );
  AOI21_X1 U19918 ( .B1(n16657), .B2(n20808), .A(n16543), .ZN(n16544) );
  OAI211_X1 U19919 ( .C1(n16547), .C2(n16546), .A(n16545), .B(n16544), .ZN(
        P1_U2817) );
  AOI22_X1 U19920 ( .A1(n20850), .A2(P1_EBX_REG_22__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n20849), .ZN(n16555) );
  INV_X1 U19921 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n21236) );
  AOI22_X1 U19922 ( .A1(n16549), .A2(n16629), .B1(n16548), .B2(n21236), .ZN(
        n16554) );
  AOI22_X1 U19923 ( .A1(n16550), .A2(n20808), .B1(n16609), .B2(n16761), .ZN(
        n16553) );
  NOR2_X1 U19924 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(n16551), .ZN(n16558) );
  OAI21_X1 U19925 ( .B1(n16558), .B2(n16570), .A(P1_REIP_REG_22__SCAN_IN), 
        .ZN(n16552) );
  NAND4_X1 U19926 ( .A1(n16555), .A2(n16554), .A3(n16553), .A4(n16552), .ZN(
        P1_U2818) );
  AOI22_X1 U19927 ( .A1(n20850), .A2(P1_EBX_REG_21__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n20849), .ZN(n16562) );
  AOI22_X1 U19928 ( .A1(n16662), .A2(n16629), .B1(P1_REIP_REG_21__SCAN_IN), 
        .B2(n16570), .ZN(n16561) );
  OAI22_X1 U19929 ( .A1(n16665), .A2(n16617), .B1(n20860), .B2(n16556), .ZN(
        n16557) );
  INV_X1 U19930 ( .A(n16557), .ZN(n16560) );
  INV_X1 U19931 ( .A(n16558), .ZN(n16559) );
  NAND4_X1 U19932 ( .A1(n16562), .A2(n16561), .A3(n16560), .A4(n16559), .ZN(
        P1_U2819) );
  AOI22_X1 U19933 ( .A1(n20850), .A2(P1_EBX_REG_20__SCAN_IN), .B1(n16629), 
        .B2(n16563), .ZN(n16572) );
  INV_X1 U19934 ( .A(n16594), .ZN(n16564) );
  OAI21_X1 U19935 ( .B1(n16565), .B2(n16564), .A(n21232), .ZN(n16569) );
  OAI22_X1 U19936 ( .A1(n16567), .A2(n16617), .B1(n20860), .B2(n16566), .ZN(
        n16568) );
  AOI21_X1 U19937 ( .B1(n16570), .B2(n16569), .A(n16568), .ZN(n16571) );
  OAI211_X1 U19938 ( .C1(n16573), .C2(n20818), .A(n16572), .B(n16571), .ZN(
        P1_U2820) );
  OAI21_X1 U19939 ( .B1(P1_REIP_REG_18__SCAN_IN), .B2(n20813), .A(n16574), 
        .ZN(n16593) );
  OAI222_X1 U19940 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(P1_REIP_REG_18__SCAN_IN), .B1(P1_REIP_REG_19__SCAN_IN), .B2(n16594), .C1(n21229), .C2(n16593), .ZN(
        n16585) );
  NOR2_X1 U19941 ( .A1(n20847), .A2(n16681), .ZN(n16577) );
  INV_X1 U19942 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n16575) );
  OAI21_X1 U19943 ( .B1(n20818), .B2(n16575), .A(n20816), .ZN(n16576) );
  AOI211_X1 U19944 ( .C1(n20850), .C2(P1_EBX_REG_19__SCAN_IN), .A(n16577), .B(
        n16576), .ZN(n16584) );
  NOR2_X1 U19945 ( .A1(n16579), .A2(n16578), .ZN(n16580) );
  OR2_X1 U19946 ( .A1(n16581), .A2(n16580), .ZN(n16769) );
  OAI22_X1 U19947 ( .A1(n16677), .A2(n16617), .B1(n20860), .B2(n16769), .ZN(
        n16582) );
  INV_X1 U19948 ( .A(n16582), .ZN(n16583) );
  NAND3_X1 U19949 ( .A1(n16585), .A2(n16584), .A3(n16583), .ZN(P1_U2821) );
  NAND2_X1 U19950 ( .A1(n20849), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n16586) );
  NAND2_X1 U19951 ( .A1(n16586), .A2(n20816), .ZN(n16587) );
  AOI21_X1 U19952 ( .B1(n20850), .B2(P1_EBX_REG_18__SCAN_IN), .A(n16587), .ZN(
        n16590) );
  NAND2_X1 U19953 ( .A1(n16588), .A2(n16629), .ZN(n16589) );
  OAI211_X1 U19954 ( .C1(n16591), .C2(n16617), .A(n16590), .B(n16589), .ZN(
        n16592) );
  INV_X1 U19955 ( .A(n16592), .ZN(n16596) );
  OAI21_X1 U19956 ( .B1(P1_REIP_REG_18__SCAN_IN), .B2(n16594), .A(n16593), 
        .ZN(n16595) );
  OAI211_X1 U19957 ( .C1(n16597), .C2(n20860), .A(n16596), .B(n16595), .ZN(
        P1_U2822) );
  INV_X1 U19958 ( .A(n16598), .ZN(n16603) );
  NAND2_X1 U19959 ( .A1(n20849), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n16599) );
  OAI211_X1 U19960 ( .C1(n16622), .C2(n16600), .A(n16599), .B(n20816), .ZN(
        n16601) );
  AOI21_X1 U19961 ( .B1(n16694), .B2(n16629), .A(n16601), .ZN(n16602) );
  OAI21_X1 U19962 ( .B1(n16603), .B2(P1_REIP_REG_16__SCAN_IN), .A(n16602), 
        .ZN(n16604) );
  AOI21_X1 U19963 ( .B1(n16695), .B2(n20808), .A(n16604), .ZN(n16607) );
  NOR3_X1 U19964 ( .A1(P1_REIP_REG_15__SCAN_IN), .A2(n21222), .A3(n16605), 
        .ZN(n16614) );
  OAI21_X1 U19965 ( .B1(n16614), .B2(n16613), .A(P1_REIP_REG_16__SCAN_IN), 
        .ZN(n16606) );
  OAI211_X1 U19966 ( .C1(n16777), .C2(n20860), .A(n16607), .B(n16606), .ZN(
        P1_U2824) );
  AOI22_X1 U19967 ( .A1(n16698), .A2(n16629), .B1(n16609), .B2(n16608), .ZN(
        n16620) );
  NAND2_X1 U19968 ( .A1(n20849), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n16610) );
  OAI211_X1 U19969 ( .C1(n16622), .C2(n16611), .A(n20816), .B(n16610), .ZN(
        n16612) );
  AOI21_X1 U19970 ( .B1(P1_REIP_REG_15__SCAN_IN), .B2(n16613), .A(n16612), 
        .ZN(n16616) );
  INV_X1 U19971 ( .A(n16614), .ZN(n16615) );
  OAI211_X1 U19972 ( .C1(n16701), .C2(n16617), .A(n16616), .B(n16615), .ZN(
        n16618) );
  INV_X1 U19973 ( .A(n16618), .ZN(n16619) );
  NAND2_X1 U19974 ( .A1(n16620), .A2(n16619), .ZN(P1_U2825) );
  OAI22_X1 U19975 ( .A1(n16788), .A2(n20860), .B1(n16622), .B2(n16621), .ZN(
        n16623) );
  INV_X1 U19976 ( .A(n16623), .ZN(n16624) );
  OAI211_X1 U19977 ( .C1(n20818), .C2(n16625), .A(n16624), .B(n20816), .ZN(
        n16626) );
  AOI221_X1 U19978 ( .B1(n16628), .B2(P1_REIP_REG_13__SCAN_IN), .C1(n16627), 
        .C2(n21219), .A(n16626), .ZN(n16631) );
  AOI22_X1 U19979 ( .A1(n16711), .A2(n20808), .B1(n16629), .B2(n16710), .ZN(
        n16630) );
  NAND2_X1 U19980 ( .A1(n16631), .A2(n16630), .ZN(P1_U2827) );
  NOR2_X1 U19981 ( .A1(n21213), .A2(n16632), .ZN(n16633) );
  AOI22_X1 U19982 ( .A1(n20850), .A2(P1_EBX_REG_10__SCAN_IN), .B1(n21215), 
        .B2(n16633), .ZN(n16634) );
  OAI21_X1 U19983 ( .B1(n20860), .B2(n16635), .A(n16634), .ZN(n16636) );
  AOI211_X1 U19984 ( .C1(n20849), .C2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n20831), .B(n16636), .ZN(n16639) );
  AOI22_X1 U19985 ( .A1(n16723), .A2(n20808), .B1(n16637), .B2(
        P1_REIP_REG_10__SCAN_IN), .ZN(n16638) );
  OAI211_X1 U19986 ( .C1(n16720), .C2(n20847), .A(n16639), .B(n16638), .ZN(
        P1_U2830) );
  OAI22_X1 U19987 ( .A1(n16677), .A2(n16640), .B1(n15543), .B2(n16769), .ZN(
        n16641) );
  INV_X1 U19988 ( .A(n16641), .ZN(n16642) );
  OAI21_X1 U19989 ( .B1(n16644), .B2(n16643), .A(n16642), .ZN(P1_U2853) );
  AOI22_X1 U19990 ( .A1(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n16734), .B1(
        n16782), .B2(P1_REIP_REG_25__SCAN_IN), .ZN(n16652) );
  NAND3_X1 U19991 ( .A1(n16645), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n16647) );
  OAI21_X1 U19992 ( .B1(n16648), .B2(n16647), .A(n16646), .ZN(n16649) );
  XOR2_X1 U19993 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .B(n16649), .Z(
        n16746) );
  AOI22_X1 U19994 ( .A1(n16746), .A2(n16740), .B1(n16650), .B2(n16739), .ZN(
        n16651) );
  OAI211_X1 U19995 ( .C1(n16743), .C2(n16653), .A(n16652), .B(n16651), .ZN(
        P1_U2974) );
  AOI22_X1 U19996 ( .A1(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n16734), .B1(
        n16782), .B2(P1_REIP_REG_23__SCAN_IN), .ZN(n16659) );
  NOR2_X1 U19997 ( .A1(n16673), .A2(n9980), .ZN(n16655) );
  MUX2_X1 U19998 ( .A(n9980), .B(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .S(
        n16673), .Z(n16654) );
  MUX2_X1 U19999 ( .A(n16655), .B(n16654), .S(n15627), .Z(n16656) );
  AOI22_X1 U20000 ( .A1(n16740), .A2(n16755), .B1(n16657), .B2(n16739), .ZN(
        n16658) );
  OAI211_X1 U20001 ( .C1(n16743), .C2(n16660), .A(n16659), .B(n16658), .ZN(
        P1_U2976) );
  INV_X1 U20002 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n16669) );
  NAND2_X1 U20003 ( .A1(n16661), .A2(n16740), .ZN(n16664) );
  NAND2_X1 U20004 ( .A1(n16662), .A2(n16722), .ZN(n16663) );
  OAI211_X1 U20005 ( .C1(n16665), .C2(n16700), .A(n16664), .B(n16663), .ZN(
        n16666) );
  INV_X1 U20006 ( .A(n16666), .ZN(n16668) );
  NAND2_X1 U20007 ( .A1(n16782), .A2(P1_REIP_REG_21__SCAN_IN), .ZN(n16667) );
  OAI211_X1 U20008 ( .C1(n16670), .C2(n16669), .A(n16668), .B(n16667), .ZN(
        P1_U2978) );
  AOI22_X1 U20009 ( .A1(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n16734), .B1(
        n16782), .B2(P1_REIP_REG_19__SCAN_IN), .ZN(n16680) );
  NAND2_X1 U20010 ( .A1(n16672), .A2(n16671), .ZN(n16676) );
  MUX2_X1 U20011 ( .A(n16674), .B(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .S(
        n16673), .Z(n16675) );
  XNOR2_X1 U20012 ( .A(n16676), .B(n16675), .ZN(n16771) );
  INV_X1 U20013 ( .A(n16677), .ZN(n16678) );
  AOI22_X1 U20014 ( .A1(n16740), .A2(n16771), .B1(n16678), .B2(n16739), .ZN(
        n16679) );
  OAI211_X1 U20015 ( .C1(n16743), .C2(n16681), .A(n16680), .B(n16679), .ZN(
        P1_U2980) );
  AOI22_X1 U20016 ( .A1(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n16734), .B1(
        n16782), .B2(P1_REIP_REG_17__SCAN_IN), .ZN(n16685) );
  AOI22_X1 U20017 ( .A1(n16683), .A2(n16739), .B1(n16722), .B2(n16682), .ZN(
        n16684) );
  OAI211_X1 U20018 ( .C1(n20773), .C2(n16686), .A(n16685), .B(n16684), .ZN(
        P1_U2982) );
  NOR2_X1 U20019 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n16776) );
  NOR2_X1 U20020 ( .A1(n16688), .A2(n16687), .ZN(n16691) );
  NOR2_X1 U20021 ( .A1(n16776), .A2(n16691), .ZN(n16693) );
  INV_X1 U20022 ( .A(n16689), .ZN(n16690) );
  OAI22_X1 U20023 ( .A1(n16693), .A2(n16692), .B1(n16691), .B2(n16690), .ZN(
        n16778) );
  AOI22_X1 U20024 ( .A1(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n16734), .B1(
        n16782), .B2(P1_REIP_REG_16__SCAN_IN), .ZN(n16697) );
  AOI22_X1 U20025 ( .A1(n16695), .A2(n16739), .B1(n16694), .B2(n16722), .ZN(
        n16696) );
  OAI211_X1 U20026 ( .C1(n20773), .C2(n16778), .A(n16697), .B(n16696), .ZN(
        P1_U2983) );
  AOI22_X1 U20027 ( .A1(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n16734), .B1(
        n16782), .B2(P1_REIP_REG_15__SCAN_IN), .ZN(n16704) );
  INV_X1 U20028 ( .A(n16698), .ZN(n16699) );
  OAI22_X1 U20029 ( .A1(n16701), .A2(n16700), .B1(n16699), .B2(n16743), .ZN(
        n16702) );
  INV_X1 U20030 ( .A(n16702), .ZN(n16703) );
  OAI211_X1 U20031 ( .C1(n16705), .C2(n20773), .A(n16704), .B(n16703), .ZN(
        P1_U2984) );
  NOR2_X1 U20032 ( .A1(n16707), .A2(n16706), .ZN(n16708) );
  XOR2_X1 U20033 ( .A(n16709), .B(n16708), .Z(n16793) );
  AOI22_X1 U20034 ( .A1(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n16734), .B1(
        n16782), .B2(P1_REIP_REG_13__SCAN_IN), .ZN(n16713) );
  AOI22_X1 U20035 ( .A1(n16711), .A2(n16739), .B1(n16722), .B2(n16710), .ZN(
        n16712) );
  OAI211_X1 U20036 ( .C1(n20773), .C2(n16793), .A(n16713), .B(n16712), .ZN(
        P1_U2986) );
  AOI22_X1 U20037 ( .A1(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n16734), .B1(
        n16782), .B2(P1_REIP_REG_12__SCAN_IN), .ZN(n16718) );
  INV_X1 U20038 ( .A(n16714), .ZN(n16715) );
  AOI22_X1 U20039 ( .A1(n16716), .A2(n16739), .B1(n16715), .B2(n16722), .ZN(
        n16717) );
  OAI211_X1 U20040 ( .C1(n16719), .C2(n20773), .A(n16718), .B(n16717), .ZN(
        P1_U2987) );
  AOI22_X1 U20041 ( .A1(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n16734), .B1(
        n16782), .B2(P1_REIP_REG_10__SCAN_IN), .ZN(n16725) );
  INV_X1 U20042 ( .A(n16720), .ZN(n16721) );
  AOI22_X1 U20043 ( .A1(n16723), .A2(n16739), .B1(n16722), .B2(n16721), .ZN(
        n16724) );
  OAI211_X1 U20044 ( .C1(n20773), .C2(n16726), .A(n16725), .B(n16724), .ZN(
        P1_U2989) );
  AOI22_X1 U20045 ( .A1(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n16734), .B1(
        n16782), .B2(P1_REIP_REG_7__SCAN_IN), .ZN(n16733) );
  INV_X1 U20046 ( .A(n16728), .ZN(n16730) );
  NAND2_X1 U20047 ( .A1(n16730), .A2(n16729), .ZN(n16731) );
  XNOR2_X1 U20048 ( .A(n9732), .B(n16731), .ZN(n16818) );
  AOI22_X1 U20049 ( .A1(n16818), .A2(n16740), .B1(n16739), .B2(n20797), .ZN(
        n16732) );
  OAI211_X1 U20050 ( .C1(n16743), .C2(n20799), .A(n16733), .B(n16732), .ZN(
        P1_U2992) );
  AOI22_X1 U20051 ( .A1(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n16734), .B1(
        n16782), .B2(P1_REIP_REG_6__SCAN_IN), .ZN(n16742) );
  NAND2_X1 U20052 ( .A1(n16737), .A2(n16736), .ZN(n16738) );
  XNOR2_X1 U20053 ( .A(n16735), .B(n16738), .ZN(n16825) );
  AOI22_X1 U20054 ( .A1(n16825), .A2(n16740), .B1(n16739), .B2(n20809), .ZN(
        n16741) );
  OAI211_X1 U20055 ( .C1(n16743), .C2(n20812), .A(n16742), .B(n16741), .ZN(
        P1_U2993) );
  INV_X1 U20056 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n16749) );
  AOI21_X1 U20057 ( .B1(P1_REIP_REG_25__SCAN_IN), .B2(n16782), .A(n16744), 
        .ZN(n16748) );
  AOI22_X1 U20058 ( .A1(n16746), .A2(n20927), .B1(n16809), .B2(n16745), .ZN(
        n16747) );
  OAI211_X1 U20059 ( .C1(n16750), .C2(n16749), .A(n16748), .B(n16747), .ZN(
        P1_U3006) );
  INV_X1 U20060 ( .A(n16751), .ZN(n16752) );
  AOI22_X1 U20061 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n16752), .B1(
        n16782), .B2(P1_REIP_REG_23__SCAN_IN), .ZN(n16757) );
  INV_X1 U20062 ( .A(n16753), .ZN(n16754) );
  AOI22_X1 U20063 ( .A1(n16755), .A2(n20927), .B1(n16809), .B2(n16754), .ZN(
        n16756) );
  OAI211_X1 U20064 ( .C1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n16758), .A(
        n16757), .B(n16756), .ZN(P1_U3008) );
  AOI22_X1 U20065 ( .A1(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n16759), .B1(
        n16782), .B2(P1_REIP_REG_22__SCAN_IN), .ZN(n16767) );
  INV_X1 U20066 ( .A(n16760), .ZN(n16762) );
  AOI22_X1 U20067 ( .A1(n16762), .A2(n20927), .B1(n16809), .B2(n16761), .ZN(
        n16766) );
  OAI211_X1 U20068 ( .C1(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A(n16764), .B(n16763), .ZN(
        n16765) );
  NAND3_X1 U20069 ( .A1(n16767), .A2(n16766), .A3(n16765), .ZN(P1_U3009) );
  AOI22_X1 U20070 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n16768), .B1(
        n16782), .B2(P1_REIP_REG_19__SCAN_IN), .ZN(n16773) );
  INV_X1 U20071 ( .A(n16769), .ZN(n16770) );
  AOI22_X1 U20072 ( .A1(n16771), .A2(n20927), .B1(n16809), .B2(n16770), .ZN(
        n16772) );
  OAI211_X1 U20073 ( .C1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n16774), .A(
        n16773), .B(n16772), .ZN(P1_U3012) );
  NOR2_X1 U20074 ( .A1(n16776), .A2(n16775), .ZN(n16781) );
  OAI22_X1 U20075 ( .A1(n16778), .A2(n16792), .B1(n20925), .B2(n16777), .ZN(
        n16779) );
  AOI21_X1 U20076 ( .B1(n16781), .B2(n16780), .A(n16779), .ZN(n16784) );
  NAND2_X1 U20077 ( .A1(n16782), .A2(P1_REIP_REG_16__SCAN_IN), .ZN(n16783) );
  OAI211_X1 U20078 ( .C1(n16786), .C2(n16785), .A(n16784), .B(n16783), .ZN(
        P1_U3015) );
  INV_X1 U20079 ( .A(n16787), .ZN(n16790) );
  OAI22_X1 U20080 ( .A1(n16788), .A2(n20925), .B1(n21219), .B2(n16823), .ZN(
        n16789) );
  AOI21_X1 U20081 ( .B1(n16790), .B2(n16796), .A(n16789), .ZN(n16791) );
  OAI21_X1 U20082 ( .B1(n16793), .B2(n16792), .A(n16791), .ZN(n16794) );
  INV_X1 U20083 ( .A(n16794), .ZN(n16795) );
  OAI21_X1 U20084 ( .B1(n16797), .B2(n16796), .A(n16795), .ZN(P1_U3018) );
  INV_X1 U20085 ( .A(n16798), .ZN(n16800) );
  AOI21_X1 U20086 ( .B1(n16800), .B2(n16809), .A(n16799), .ZN(n16805) );
  NOR2_X1 U20087 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n16801), .ZN(
        n16802) );
  AOI22_X1 U20088 ( .A1(n16803), .A2(n20927), .B1(n16802), .B2(n16822), .ZN(
        n16804) );
  OAI211_X1 U20089 ( .C1(n16807), .C2(n16806), .A(n16805), .B(n16804), .ZN(
        P1_U3020) );
  AOI21_X1 U20090 ( .B1(n16810), .B2(n16809), .A(n16808), .ZN(n16814) );
  AOI22_X1 U20091 ( .A1(n16812), .A2(n20927), .B1(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n16811), .ZN(n16813) );
  OAI211_X1 U20092 ( .C1(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n16815), .A(
        n16814), .B(n16813), .ZN(P1_U3022) );
  OAI22_X1 U20093 ( .A1(n20795), .A2(n20925), .B1(n16823), .B2(n21208), .ZN(
        n16816) );
  INV_X1 U20094 ( .A(n16816), .ZN(n16820) );
  AOI22_X1 U20095 ( .A1(n16818), .A2(n20927), .B1(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n16817), .ZN(n16819) );
  OAI211_X1 U20096 ( .C1(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .C2(n16821), .A(
        n16820), .B(n16819), .ZN(P1_U3024) );
  INV_X1 U20097 ( .A(n16822), .ZN(n16829) );
  OAI22_X1 U20098 ( .A1(n20802), .A2(n20925), .B1(n21206), .B2(n16823), .ZN(
        n16824) );
  AOI21_X1 U20099 ( .B1(n16825), .B2(n20927), .A(n16824), .ZN(n16826) );
  OAI221_X1 U20100 ( .B1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n16829), .C1(
        n16828), .C2(n16827), .A(n16826), .ZN(P1_U3025) );
  INV_X1 U20101 ( .A(n16830), .ZN(n16831) );
  NAND3_X1 U20102 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n21113), .A3(n16831), 
        .ZN(n16832) );
  NAND2_X1 U20103 ( .A1(n16833), .A2(n16832), .ZN(n21175) );
  OAI21_X1 U20104 ( .B1(n16835), .B2(n21175), .A(n16834), .ZN(n16836) );
  OAI221_X1 U20105 ( .B1(n16837), .B2(n20953), .C1(n16837), .C2(n21287), .A(
        n16836), .ZN(n16838) );
  AOI221_X1 U20106 ( .B1(n16840), .B2(n16839), .C1(n9954), .C2(n16839), .A(
        n16838), .ZN(P1_U3162) );
  NOR2_X1 U20107 ( .A1(n16840), .A2(n9954), .ZN(n16842) );
  OAI22_X1 U20108 ( .A1(n20953), .A2(n16842), .B1(n16841), .B2(n9954), .ZN(
        P1_U3466) );
  AOI22_X1 U20109 ( .A1(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n19929), .B1(
        P2_REIP_REG_30__SCAN_IN), .B2(n19927), .ZN(n16853) );
  INV_X1 U20110 ( .A(n16843), .ZN(n16844) );
  AOI22_X1 U20111 ( .A1(n16844), .A2(n19877), .B1(P2_EBX_REG_30__SCAN_IN), 
        .B2(n19917), .ZN(n16852) );
  INV_X1 U20112 ( .A(n16845), .ZN(n16846) );
  AOI22_X1 U20113 ( .A1(n16846), .A2(n19922), .B1(n19915), .B2(n15144), .ZN(
        n16851) );
  OAI211_X1 U20114 ( .C1(n16849), .C2(n16848), .A(n19897), .B(n16847), .ZN(
        n16850) );
  NAND4_X1 U20115 ( .A1(n16853), .A2(n16852), .A3(n16851), .A4(n16850), .ZN(
        P2_U2825) );
  AOI22_X1 U20116 ( .A1(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n19929), .B1(
        P2_REIP_REG_29__SCAN_IN), .B2(n19927), .ZN(n16865) );
  INV_X1 U20117 ( .A(n16854), .ZN(n16855) );
  AOI22_X1 U20118 ( .A1(n16855), .A2(n19877), .B1(P2_EBX_REG_29__SCAN_IN), 
        .B2(n19917), .ZN(n16864) );
  INV_X1 U20119 ( .A(n16856), .ZN(n16858) );
  AOI22_X1 U20120 ( .A1(n16858), .A2(n19922), .B1(n19915), .B2(n16857), .ZN(
        n16863) );
  OAI211_X1 U20121 ( .C1(n16861), .C2(n16860), .A(n19897), .B(n16859), .ZN(
        n16862) );
  NAND4_X1 U20122 ( .A1(n16865), .A2(n16864), .A3(n16863), .A4(n16862), .ZN(
        P2_U2826) );
  AOI22_X1 U20123 ( .A1(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n19929), .B1(
        P2_REIP_REG_28__SCAN_IN), .B2(n19927), .ZN(n16876) );
  AOI22_X1 U20124 ( .A1(n16866), .A2(n19877), .B1(P2_EBX_REG_28__SCAN_IN), 
        .B2(n19917), .ZN(n16875) );
  INV_X1 U20125 ( .A(n16867), .ZN(n16868) );
  AOI22_X1 U20126 ( .A1(n16869), .A2(n19922), .B1(n16868), .B2(n19915), .ZN(
        n16874) );
  OAI211_X1 U20127 ( .C1(n16872), .C2(n16871), .A(n19897), .B(n16870), .ZN(
        n16873) );
  NAND4_X1 U20128 ( .A1(n16876), .A2(n16875), .A3(n16874), .A4(n16873), .ZN(
        P2_U2827) );
  NOR2_X1 U20129 ( .A1(n19888), .A2(n11011), .ZN(n16878) );
  OAI22_X1 U20130 ( .A1(n10080), .A2(n19815), .B1(n20675), .B2(n19887), .ZN(
        n16877) );
  NOR2_X1 U20131 ( .A1(n16878), .A2(n16877), .ZN(n16879) );
  OAI21_X1 U20132 ( .B1(n16880), .B2(n19919), .A(n16879), .ZN(n16881) );
  AOI21_X1 U20133 ( .B1(n16882), .B2(n19922), .A(n16881), .ZN(n16887) );
  OAI211_X1 U20134 ( .C1(n16885), .C2(n16884), .A(n19897), .B(n16883), .ZN(
        n16886) );
  OAI211_X1 U20135 ( .C1(n19914), .C2(n16888), .A(n16887), .B(n16886), .ZN(
        P2_U2828) );
  AOI22_X1 U20136 ( .A1(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n19929), .B1(
        P2_REIP_REG_26__SCAN_IN), .B2(n19927), .ZN(n16899) );
  AOI22_X1 U20137 ( .A1(n16889), .A2(n19877), .B1(P2_EBX_REG_26__SCAN_IN), 
        .B2(n19917), .ZN(n16898) );
  INV_X1 U20138 ( .A(n16890), .ZN(n16892) );
  AOI22_X1 U20139 ( .A1(n16892), .A2(n19922), .B1(n16891), .B2(n19915), .ZN(
        n16897) );
  OAI211_X1 U20140 ( .C1(n16895), .C2(n16894), .A(n19897), .B(n16893), .ZN(
        n16896) );
  NAND4_X1 U20141 ( .A1(n16899), .A2(n16898), .A3(n16897), .A4(n16896), .ZN(
        P2_U2829) );
  AOI22_X1 U20142 ( .A1(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n19929), .B1(
        P2_REIP_REG_23__SCAN_IN), .B2(n19927), .ZN(n16909) );
  AOI22_X1 U20143 ( .A1(n16900), .A2(n19877), .B1(P2_EBX_REG_23__SCAN_IN), 
        .B2(n19917), .ZN(n16908) );
  AOI22_X1 U20144 ( .A1(n16902), .A2(n19922), .B1(n16901), .B2(n19915), .ZN(
        n16907) );
  OAI211_X1 U20145 ( .C1(n16905), .C2(n16904), .A(n19897), .B(n16903), .ZN(
        n16906) );
  NAND4_X1 U20146 ( .A1(n16909), .A2(n16908), .A3(n16907), .A4(n16906), .ZN(
        P2_U2832) );
  AOI22_X1 U20147 ( .A1(n19969), .A2(n12092), .B1(n12107), .B2(n19947), .ZN(
        P2_U2856) );
  NOR2_X1 U20148 ( .A1(n16910), .A2(n20755), .ZN(n16911) );
  XNOR2_X1 U20149 ( .A(n16912), .B(n16911), .ZN(n16913) );
  XNOR2_X1 U20150 ( .A(n16914), .B(n16913), .ZN(n16937) );
  AOI22_X1 U20151 ( .A1(n16937), .A2(n16926), .B1(n19965), .B2(n16915), .ZN(
        n16916) );
  OAI21_X1 U20152 ( .B1(n19969), .B2(n10814), .A(n16916), .ZN(P2_U2863) );
  INV_X1 U20153 ( .A(n16917), .ZN(n16918) );
  AOI22_X1 U20154 ( .A1(n16918), .A2(n16926), .B1(P2_EBX_REG_21__SCAN_IN), 
        .B2(n19947), .ZN(n16919) );
  OAI21_X1 U20155 ( .B1(n19947), .B2(n16920), .A(n16919), .ZN(P2_U2866) );
  OAI22_X1 U20156 ( .A1(n16921), .A2(n19959), .B1(n19969), .B2(n10747), .ZN(
        n16922) );
  INV_X1 U20157 ( .A(n16922), .ZN(n16923) );
  OAI21_X1 U20158 ( .B1(n19947), .B2(n16924), .A(n16923), .ZN(P2_U2868) );
  INV_X1 U20159 ( .A(n16925), .ZN(n16927) );
  AOI22_X1 U20160 ( .A1(n16927), .A2(n16926), .B1(P2_EBX_REG_17__SCAN_IN), 
        .B2(n19947), .ZN(n16928) );
  OAI21_X1 U20161 ( .B1(n19947), .B2(n16929), .A(n16928), .ZN(P2_U2870) );
  INV_X1 U20162 ( .A(n16930), .ZN(n16931) );
  AOI22_X1 U20163 ( .A1(n16931), .A2(n19975), .B1(P2_EAX_REG_24__SCAN_IN), 
        .B2(n19974), .ZN(n16940) );
  AOI22_X1 U20164 ( .A1(n16933), .A2(BUF2_REG_24__SCAN_IN), .B1(n16932), .B2(
        BUF1_REG_24__SCAN_IN), .ZN(n16939) );
  AOI22_X1 U20165 ( .A1(n16937), .A2(n16936), .B1(n16935), .B2(n16934), .ZN(
        n16938) );
  NAND3_X1 U20166 ( .A1(n16940), .A2(n16939), .A3(n16938), .ZN(P2_U2895) );
  AOI22_X1 U20167 ( .A1(P2_REIP_REG_15__SCAN_IN), .A2(n20028), .B1(n17008), 
        .B2(n19822), .ZN(n16951) );
  NAND2_X1 U20168 ( .A1(n16942), .A2(n16941), .ZN(n16943) );
  XNOR2_X1 U20169 ( .A(n16944), .B(n16943), .ZN(n17023) );
  INV_X1 U20170 ( .A(n17023), .ZN(n16949) );
  NAND2_X1 U20171 ( .A1(n13714), .A2(n16945), .ZN(n16946) );
  NAND2_X1 U20172 ( .A1(n16947), .A2(n16946), .ZN(n19940) );
  INV_X1 U20173 ( .A(n19940), .ZN(n19823) );
  XNOR2_X1 U20174 ( .A(n16948), .B(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n17020) );
  AOI222_X1 U20175 ( .A1(n16949), .A2(n20046), .B1(n20051), .B2(n19823), .C1(
        n17010), .C2(n17020), .ZN(n16950) );
  OAI211_X1 U20176 ( .C1(n19816), .C2(n20055), .A(n16951), .B(n16950), .ZN(
        P2_U2999) );
  AOI22_X1 U20177 ( .A1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n20029), .B1(
        P2_REIP_REG_14__SCAN_IN), .B2(n19905), .ZN(n16956) );
  OAI22_X1 U20178 ( .A1(n16953), .A2(n16974), .B1(n20043), .B2(n16952), .ZN(
        n16954) );
  AOI21_X1 U20179 ( .B1(n20051), .B2(n19835), .A(n16954), .ZN(n16955) );
  OAI211_X1 U20180 ( .C1(n20045), .C2(n19829), .A(n16956), .B(n16955), .ZN(
        P2_U3000) );
  AOI22_X1 U20181 ( .A1(P2_REIP_REG_13__SCAN_IN), .A2(n20028), .B1(n17008), 
        .B2(n19844), .ZN(n16970) );
  NAND2_X1 U20182 ( .A1(n16959), .A2(n16958), .ZN(n16960) );
  XNOR2_X1 U20183 ( .A(n16957), .B(n16960), .ZN(n17031) );
  INV_X1 U20184 ( .A(n17031), .ZN(n16968) );
  OR2_X1 U20185 ( .A1(n16961), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n16962) );
  AND2_X1 U20186 ( .A1(n16965), .A2(n16964), .ZN(n16967) );
  OR2_X1 U20187 ( .A1(n16967), .A2(n16966), .ZN(n19948) );
  INV_X1 U20188 ( .A(n19948), .ZN(n19845) );
  AOI222_X1 U20189 ( .A1(n16968), .A2(n20046), .B1(n17028), .B2(n17010), .C1(
        n20051), .C2(n19845), .ZN(n16969) );
  OAI211_X1 U20190 ( .C1(n16971), .C2(n20055), .A(n16970), .B(n16969), .ZN(
        P2_U3001) );
  AOI22_X1 U20191 ( .A1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n20029), .B1(
        P2_REIP_REG_12__SCAN_IN), .B2(n19905), .ZN(n16978) );
  INV_X1 U20192 ( .A(n16972), .ZN(n16975) );
  OAI22_X1 U20193 ( .A1(n16975), .A2(n20043), .B1(n16974), .B2(n16973), .ZN(
        n16976) );
  AOI21_X1 U20194 ( .B1(n20051), .B2(n19856), .A(n16976), .ZN(n16977) );
  OAI211_X1 U20195 ( .C1(n20045), .C2(n19852), .A(n16978), .B(n16977), .ZN(
        P2_U3002) );
  AOI22_X1 U20196 ( .A1(P2_REIP_REG_11__SCAN_IN), .A2(n20028), .B1(n17008), 
        .B2(n19869), .ZN(n16985) );
  NAND2_X1 U20197 ( .A1(n16979), .A2(n20046), .ZN(n16981) );
  NAND2_X1 U20198 ( .A1(n20051), .A2(n19954), .ZN(n16980) );
  OAI211_X1 U20199 ( .C1(n16982), .C2(n20043), .A(n16981), .B(n16980), .ZN(
        n16983) );
  INV_X1 U20200 ( .A(n16983), .ZN(n16984) );
  OAI211_X1 U20201 ( .C1(n16986), .C2(n20055), .A(n16985), .B(n16984), .ZN(
        P2_U3003) );
  AOI22_X1 U20202 ( .A1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n20029), .B1(
        P2_REIP_REG_10__SCAN_IN), .B2(n19905), .ZN(n16998) );
  XOR2_X1 U20203 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .B(n16987), .Z(
        n17039) );
  INV_X1 U20204 ( .A(n17039), .ZN(n16994) );
  NAND2_X1 U20205 ( .A1(n16401), .A2(n16988), .ZN(n16993) );
  INV_X1 U20206 ( .A(n16989), .ZN(n16990) );
  NOR2_X1 U20207 ( .A1(n16991), .A2(n16990), .ZN(n16992) );
  XNOR2_X1 U20208 ( .A(n16993), .B(n16992), .ZN(n17041) );
  OAI22_X1 U20209 ( .A1(n16994), .A2(n20043), .B1(n17041), .B2(n16974), .ZN(
        n16995) );
  AOI21_X1 U20210 ( .B1(n20051), .B2(n16996), .A(n16995), .ZN(n16997) );
  OAI211_X1 U20211 ( .C1(n20045), .C2(n16999), .A(n16998), .B(n16997), .ZN(
        P2_U3004) );
  AOI22_X1 U20212 ( .A1(P2_REIP_REG_9__SCAN_IN), .A2(n20028), .B1(n17008), 
        .B2(n17000), .ZN(n17006) );
  INV_X1 U20213 ( .A(n17001), .ZN(n17004) );
  INV_X1 U20214 ( .A(n17002), .ZN(n19964) );
  AOI222_X1 U20215 ( .A1(n17004), .A2(n17010), .B1(n17003), .B2(n20046), .C1(
        n20051), .C2(n19964), .ZN(n17005) );
  OAI211_X1 U20216 ( .C1(n17007), .C2(n20055), .A(n17006), .B(n17005), .ZN(
        P2_U3005) );
  AOI22_X1 U20217 ( .A1(P2_REIP_REG_5__SCAN_IN), .A2(n20028), .B1(n17008), 
        .B2(n19908), .ZN(n17013) );
  AOI222_X1 U20218 ( .A1(n17011), .A2(n17010), .B1(n20051), .B2(n19909), .C1(
        n20046), .C2(n17009), .ZN(n17012) );
  OAI211_X1 U20219 ( .C1(n17014), .C2(n20055), .A(n17013), .B(n17012), .ZN(
        P2_U3009) );
  NOR2_X1 U20220 ( .A1(n10972), .A2(n12009), .ZN(n17018) );
  INV_X1 U20221 ( .A(n17015), .ZN(n17016) );
  OAI22_X1 U20222 ( .A1(n17048), .A2(n19827), .B1(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n17016), .ZN(n17017) );
  AOI211_X1 U20223 ( .C1(n17019), .C2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n17018), .B(n17017), .ZN(n17022) );
  AOI22_X1 U20224 ( .A1(n17020), .A2(n17052), .B1(n17074), .B2(n19823), .ZN(
        n17021) );
  OAI211_X1 U20225 ( .C1(n17023), .C2(n17071), .A(n17022), .B(n17021), .ZN(
        P2_U3031) );
  AOI21_X1 U20226 ( .B1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n17024), .A(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n17025) );
  OAI22_X1 U20227 ( .A1(n17026), .A2(n17025), .B1(n17048), .B2(n19849), .ZN(
        n17027) );
  AOI21_X1 U20228 ( .B1(P2_REIP_REG_13__SCAN_IN), .B2(n19905), .A(n17027), 
        .ZN(n17030) );
  AOI22_X1 U20229 ( .A1(n17028), .A2(n17052), .B1(n17074), .B2(n19845), .ZN(
        n17029) );
  OAI211_X1 U20230 ( .C1(n17071), .C2(n17031), .A(n17030), .B(n17029), .ZN(
        P2_U3033) );
  NAND2_X1 U20231 ( .A1(P2_REIP_REG_10__SCAN_IN), .A2(n19905), .ZN(n17032) );
  OAI221_X1 U20232 ( .B1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n17034), 
        .C1(n10722), .C2(n17033), .A(n17032), .ZN(n17038) );
  OAI22_X1 U20233 ( .A1(n20062), .A2(n17036), .B1(n17048), .B2(n17035), .ZN(
        n17037) );
  AOI211_X1 U20234 ( .C1(n17039), .C2(n17052), .A(n17038), .B(n17037), .ZN(
        n17040) );
  OAI21_X1 U20235 ( .B1(n17041), .B2(n17071), .A(n17040), .ZN(P2_U3036) );
  NOR2_X1 U20236 ( .A1(n17042), .A2(n20061), .ZN(n17046) );
  OR2_X1 U20237 ( .A1(n17044), .A2(n17043), .ZN(n17045) );
  MUX2_X1 U20238 ( .A(n17046), .B(n17045), .S(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .Z(n17050) );
  INV_X1 U20239 ( .A(n17047), .ZN(n19978) );
  OAI22_X1 U20240 ( .A1(n17048), .A2(n19978), .B1(n10945), .B2(n20073), .ZN(
        n17049) );
  NOR2_X1 U20241 ( .A1(n17050), .A2(n17049), .ZN(n17055) );
  AOI22_X1 U20242 ( .A1(n17053), .A2(n17052), .B1(n17074), .B2(n17051), .ZN(
        n17054) );
  OAI211_X1 U20243 ( .C1(n17056), .C2(n17071), .A(n17055), .B(n17054), .ZN(
        P2_U3038) );
  AOI21_X1 U20244 ( .B1(n20057), .B2(n20700), .A(n17057), .ZN(n17059) );
  OAI211_X1 U20245 ( .C1(n17060), .C2(n20068), .A(n17059), .B(n17058), .ZN(
        n17061) );
  AOI21_X1 U20246 ( .B1(n20059), .B2(n17062), .A(n17061), .ZN(n17063) );
  OAI221_X1 U20247 ( .B1(n17066), .B2(n17065), .C1(n17066), .C2(n17064), .A(
        n17063), .ZN(P2_U3043) );
  AOI22_X1 U20248 ( .A1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n17067), .B1(
        n20057), .B2(n19916), .ZN(n17076) );
  INV_X1 U20249 ( .A(n17068), .ZN(n17069) );
  OAI22_X1 U20250 ( .A1(n17071), .A2(n17070), .B1(n20068), .B2(n17069), .ZN(
        n17072) );
  AOI211_X1 U20251 ( .C1(n17074), .C2(n19923), .A(n17073), .B(n17072), .ZN(
        n17075) );
  OAI211_X1 U20252 ( .C1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(n17077), .A(
        n17076), .B(n17075), .ZN(P2_U3046) );
  AOI211_X1 U20253 ( .C1(n17081), .C2(n17080), .A(n17079), .B(n17078), .ZN(
        n17087) );
  MUX2_X1 U20254 ( .A(n20609), .B(n17082), .S(n20749), .Z(n17083) );
  NAND2_X1 U20255 ( .A1(n17083), .A2(n20753), .ZN(n17085) );
  INV_X1 U20256 ( .A(n20609), .ZN(n20612) );
  NAND3_X1 U20257 ( .A1(n20612), .A2(n20744), .A3(n20749), .ZN(n17084) );
  NAND2_X1 U20258 ( .A1(n17085), .A2(n17084), .ZN(n17086) );
  OAI211_X1 U20259 ( .C1(n17089), .C2(n17088), .A(n17087), .B(n17086), .ZN(
        P2_U3176) );
  NAND2_X1 U20260 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n12931), .ZN(
        n17095) );
  OAI221_X1 U20261 ( .B1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n17140), 
        .C1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .C2(n12931), .A(n17093), .ZN(
        n17091) );
  INV_X1 U20262 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n19661) );
  OAI22_X1 U20263 ( .A1(n17091), .A2(n17092), .B1(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n19661), .ZN(n17094) );
  INV_X1 U20264 ( .A(n19020), .ZN(n19693) );
  INV_X1 U20265 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n19637) );
  NOR2_X1 U20266 ( .A1(n19637), .A2(n19013), .ZN(n17142) );
  NOR2_X1 U20267 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n19712), .ZN(n18445) );
  NAND2_X1 U20268 ( .A1(n19388), .A2(n19116), .ZN(n19354) );
  OR2_X1 U20269 ( .A1(n17097), .A2(n18483), .ZN(n17110) );
  XOR2_X1 U20270 ( .A(n12659), .B(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .Z(
        n17099) );
  NOR2_X1 U20271 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n18430), .ZN(
        n17132) );
  INV_X1 U20272 ( .A(n18445), .ZN(n19560) );
  INV_X2 U20273 ( .A(n19354), .ZN(n19423) );
  NAND2_X1 U20274 ( .A1(n19423), .A2(n17097), .ZN(n17120) );
  OAI211_X1 U20275 ( .C1(n17098), .C2(n19560), .A(n18684), .B(n17120), .ZN(
        n17121) );
  NOR2_X1 U20276 ( .A1(n17132), .A2(n17121), .ZN(n17108) );
  OAI22_X1 U20277 ( .A1(n17110), .A2(n17099), .B1(n17108), .B2(n12659), .ZN(
        n17100) );
  AOI211_X1 U20278 ( .C1(n18547), .C2(n10033), .A(n17142), .B(n17100), .ZN(
        n17106) );
  NAND2_X1 U20279 ( .A1(n17126), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n17102) );
  XNOR2_X1 U20280 ( .A(n17102), .B(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n17145) );
  NAND2_X1 U20281 ( .A1(n17124), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n17104) );
  XNOR2_X1 U20282 ( .A(n17104), .B(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n17144) );
  AOI22_X1 U20283 ( .A1(n18674), .A2(n17145), .B1(n9716), .B2(n17144), .ZN(
        n17105) );
  OAI211_X1 U20284 ( .C1(n17148), .C2(n18540), .A(n17106), .B(n17105), .ZN(
        P3_U2799) );
  NAND2_X1 U20285 ( .A1(n18948), .A2(P3_REIP_REG_30__SCAN_IN), .ZN(n17107) );
  OAI221_X1 U20286 ( .B1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n17110), .C1(
        n17109), .C2(n17108), .A(n17107), .ZN(n17111) );
  AOI21_X1 U20287 ( .B1(n18547), .B2(n17289), .A(n17111), .ZN(n17118) );
  INV_X1 U20288 ( .A(n9716), .ZN(n18594) );
  OAI22_X1 U20289 ( .A1(n17126), .A2(n18689), .B1(n17124), .B2(n18594), .ZN(
        n17116) );
  INV_X1 U20290 ( .A(n17113), .ZN(n17114) );
  NOR3_X1 U20291 ( .A1(n18586), .A2(n17114), .A3(n18393), .ZN(n18349) );
  AOI22_X1 U20292 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n17116), .B1(
        n17115), .B2(n18349), .ZN(n17117) );
  OAI211_X1 U20293 ( .C1(n17119), .C2(n18540), .A(n17118), .B(n17117), .ZN(
        P3_U2800) );
  INV_X1 U20294 ( .A(n17120), .ZN(n17122) );
  AOI22_X1 U20295 ( .A1(n9848), .A2(n17122), .B1(
        P3_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n17121), .ZN(n17136) );
  NOR2_X1 U20296 ( .A1(n17152), .A2(n17123), .ZN(n17155) );
  INV_X1 U20297 ( .A(n17155), .ZN(n17125) );
  AOI211_X1 U20298 ( .C1(n17128), .C2(n17125), .A(n17124), .B(n18594), .ZN(
        n17130) );
  OR2_X1 U20299 ( .A1(n18327), .A2(n17152), .ZN(n17127) );
  AOI211_X1 U20300 ( .C1(n17128), .C2(n17127), .A(n17126), .B(n18689), .ZN(
        n17129) );
  OAI21_X1 U20301 ( .B1(n17132), .B2(n18547), .A(n17300), .ZN(n17133) );
  NAND4_X1 U20302 ( .A1(n17135), .A2(n17136), .A3(n17134), .A4(n17133), .ZN(
        P3_U2801) );
  NAND2_X1 U20303 ( .A1(n17138), .A2(n17137), .ZN(n17139) );
  OAI33_X1 U20304 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n19001), .A3(
        n19661), .B1(n17140), .B2(n17139), .B3(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n17141) );
  AOI211_X1 U20305 ( .C1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .C2(n17143), .A(
        n17142), .B(n17141), .ZN(n17147) );
  AOI22_X1 U20306 ( .A1(n17145), .A2(n18832), .B1(n17144), .B2(n18862), .ZN(
        n17146) );
  AOI22_X1 U20307 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n12931), .B1(
        n18509), .B2(n18328), .ZN(n18324) );
  AOI21_X1 U20308 ( .B1(n18509), .B2(n17159), .A(n17158), .ZN(n18325) );
  NOR2_X1 U20309 ( .A1(n18324), .A2(n18325), .ZN(n18326) );
  OR2_X1 U20310 ( .A1(n17149), .A2(n18171), .ZN(n17150) );
  NOR3_X1 U20311 ( .A1(n18326), .A2(n17151), .A3(n17150), .ZN(n17157) );
  INV_X1 U20312 ( .A(n19483), .ZN(n18891) );
  OAI21_X1 U20313 ( .B1(n18327), .B2(n17152), .A(n18891), .ZN(n17153) );
  OAI211_X1 U20314 ( .C1(n17155), .C2(n18871), .A(n17154), .B(n17153), .ZN(
        n17156) );
  OAI211_X1 U20315 ( .C1(n17157), .C2(n17156), .A(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B(n19013), .ZN(n17169) );
  NAND3_X1 U20316 ( .A1(n17158), .A2(n18926), .A3(n18324), .ZN(n17168) );
  INV_X1 U20317 ( .A(n17159), .ZN(n18342) );
  NAND3_X1 U20318 ( .A1(n18342), .A2(n19012), .A3(n17160), .ZN(n17167) );
  INV_X1 U20319 ( .A(n18871), .ZN(n18834) );
  AOI22_X1 U20320 ( .A1(n18891), .A2(n18512), .B1(n17112), .B2(n18834), .ZN(
        n18797) );
  INV_X1 U20321 ( .A(n18456), .ZN(n17163) );
  INV_X1 U20322 ( .A(n17161), .ZN(n17162) );
  OAI21_X1 U20323 ( .B1(n18797), .B2(n17163), .A(n17162), .ZN(n18704) );
  NAND2_X1 U20324 ( .A1(n17164), .A2(n18704), .ZN(n18743) );
  NOR2_X1 U20325 ( .A1(n17165), .A2(n18743), .ZN(n18700) );
  NOR2_X1 U20326 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n10095), .ZN(
        n18330) );
  AOI22_X1 U20327 ( .A1(n18866), .A2(P3_REIP_REG_28__SCAN_IN), .B1(n18700), 
        .B2(n18330), .ZN(n17166) );
  NAND4_X1 U20328 ( .A1(n17169), .A2(n17168), .A3(n17167), .A4(n17166), .ZN(
        P3_U2834) );
  NOR3_X1 U20329 ( .A1(P3_D_C_N_REG_SCAN_IN), .A2(P3_W_R_N_REG_SCAN_IN), .A3(
        P3_BE_N_REG_0__SCAN_IN), .ZN(n17171) );
  NOR4_X1 U20330 ( .A1(P3_BE_N_REG_1__SCAN_IN), .A2(P3_BE_N_REG_2__SCAN_IN), 
        .A3(P3_BE_N_REG_3__SCAN_IN), .A4(P3_ADS_N_REG_SCAN_IN), .ZN(n17170) );
  NAND4_X1 U20331 ( .A1(P3_M_IO_N_REG_SCAN_IN), .A2(n17171), .A3(n17170), .A4(
        U215), .ZN(U213) );
  INV_X1 U20332 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n19989) );
  NOR2_X2 U20333 ( .A1(n17216), .A2(n17172), .ZN(n17220) );
  INV_X1 U20334 ( .A(n17220), .ZN(n17218) );
  OAI222_X1 U20335 ( .A1(U212), .A2(n19989), .B1(n17218), .B2(n17173), .C1(
        U214), .C2(n17257), .ZN(U216) );
  INV_X1 U20336 ( .A(BUF1_REG_30__SCAN_IN), .ZN(n20112) );
  INV_X1 U20337 ( .A(U212), .ZN(n17215) );
  AOI22_X1 U20338 ( .A1(P1_DATAO_REG_30__SCAN_IN), .A2(n17216), .B1(
        P2_DATAO_REG_30__SCAN_IN), .B2(n17215), .ZN(n17174) );
  OAI21_X1 U20339 ( .B1(n20112), .B2(n17218), .A(n17174), .ZN(U217) );
  INV_X1 U20340 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n17176) );
  AOI22_X1 U20341 ( .A1(P1_DATAO_REG_29__SCAN_IN), .A2(n17216), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n17215), .ZN(n17175) );
  OAI21_X1 U20342 ( .B1(n17176), .B2(n17218), .A(n17175), .ZN(U218) );
  AOI22_X1 U20343 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(n17216), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(n17215), .ZN(n17177) );
  OAI21_X1 U20344 ( .B1(n20103), .B2(n17218), .A(n17177), .ZN(U219) );
  AOI222_X1 U20345 ( .A1(n17215), .A2(P2_DATAO_REG_27__SCAN_IN), .B1(n17220), 
        .B2(BUF1_REG_27__SCAN_IN), .C1(n17216), .C2(P1_DATAO_REG_27__SCAN_IN), 
        .ZN(n17178) );
  INV_X1 U20346 ( .A(n17178), .ZN(U220) );
  INV_X1 U20347 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n17180) );
  AOI22_X1 U20348 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(n17216), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n17215), .ZN(n17179) );
  OAI21_X1 U20349 ( .B1(n17180), .B2(n17218), .A(n17179), .ZN(U221) );
  INV_X1 U20350 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n17182) );
  AOI22_X1 U20351 ( .A1(P1_DATAO_REG_25__SCAN_IN), .A2(n17216), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(n17215), .ZN(n17181) );
  OAI21_X1 U20352 ( .B1(n17182), .B2(n17218), .A(n17181), .ZN(U222) );
  INV_X1 U20353 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n17184) );
  AOI22_X1 U20354 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n17216), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(n17215), .ZN(n17183) );
  OAI21_X1 U20355 ( .B1(n17184), .B2(n17218), .A(n17183), .ZN(U223) );
  INV_X1 U20356 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n17186) );
  AOI22_X1 U20357 ( .A1(P1_DATAO_REG_23__SCAN_IN), .A2(n17216), .B1(
        P2_DATAO_REG_23__SCAN_IN), .B2(n17215), .ZN(n17185) );
  OAI21_X1 U20358 ( .B1(n17186), .B2(n17218), .A(n17185), .ZN(U224) );
  INV_X1 U20359 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n17188) );
  AOI22_X1 U20360 ( .A1(P1_DATAO_REG_22__SCAN_IN), .A2(n17216), .B1(
        P2_DATAO_REG_22__SCAN_IN), .B2(n17215), .ZN(n17187) );
  OAI21_X1 U20361 ( .B1(n17188), .B2(n17218), .A(n17187), .ZN(U225) );
  INV_X1 U20362 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n17190) );
  AOI22_X1 U20363 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(n17216), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(n17215), .ZN(n17189) );
  OAI21_X1 U20364 ( .B1(n17190), .B2(n17218), .A(n17189), .ZN(U226) );
  AOI22_X1 U20365 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n17220), .B1(
        P1_DATAO_REG_20__SCAN_IN), .B2(n17216), .ZN(n17191) );
  OAI21_X1 U20366 ( .B1(n17243), .B2(U212), .A(n17191), .ZN(U227) );
  INV_X1 U20367 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n20097) );
  INV_X1 U20368 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n17192) );
  OAI222_X1 U20369 ( .A1(U212), .A2(n17242), .B1(n17218), .B2(n20097), .C1(
        U214), .C2(n17192), .ZN(U228) );
  INV_X1 U20370 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n17194) );
  AOI22_X1 U20371 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(n17216), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n17215), .ZN(n17193) );
  OAI21_X1 U20372 ( .B1(n17194), .B2(n17218), .A(n17193), .ZN(U229) );
  AOI22_X1 U20373 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n17220), .B1(
        P1_DATAO_REG_17__SCAN_IN), .B2(n17216), .ZN(n17195) );
  OAI21_X1 U20374 ( .B1(n17240), .B2(U212), .A(n17195), .ZN(U230) );
  INV_X1 U20375 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n17197) );
  AOI22_X1 U20376 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n17216), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n17215), .ZN(n17196) );
  OAI21_X1 U20377 ( .B1(n17197), .B2(n17218), .A(n17196), .ZN(U231) );
  INV_X1 U20378 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n17237) );
  AOI22_X1 U20379 ( .A1(BUF1_REG_15__SCAN_IN), .A2(n17220), .B1(
        P1_DATAO_REG_15__SCAN_IN), .B2(n17216), .ZN(n17198) );
  OAI21_X1 U20380 ( .B1(n17237), .B2(U212), .A(n17198), .ZN(U232) );
  AOI22_X1 U20381 ( .A1(P1_DATAO_REG_14__SCAN_IN), .A2(n17216), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n17215), .ZN(n17199) );
  OAI21_X1 U20382 ( .B1(n17200), .B2(n17218), .A(n17199), .ZN(U233) );
  INV_X1 U20383 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n17234) );
  AOI22_X1 U20384 ( .A1(BUF1_REG_13__SCAN_IN), .A2(n17220), .B1(
        P1_DATAO_REG_13__SCAN_IN), .B2(n17216), .ZN(n17201) );
  OAI21_X1 U20385 ( .B1(n17234), .B2(U212), .A(n17201), .ZN(U234) );
  INV_X1 U20386 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n17233) );
  AOI22_X1 U20387 ( .A1(BUF1_REG_12__SCAN_IN), .A2(n17220), .B1(
        P1_DATAO_REG_12__SCAN_IN), .B2(n17216), .ZN(n17202) );
  OAI21_X1 U20388 ( .B1(n17233), .B2(U212), .A(n17202), .ZN(U235) );
  INV_X1 U20389 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n17232) );
  AOI22_X1 U20390 ( .A1(BUF1_REG_11__SCAN_IN), .A2(n17220), .B1(
        P1_DATAO_REG_11__SCAN_IN), .B2(n17216), .ZN(n17203) );
  OAI21_X1 U20391 ( .B1(n17232), .B2(U212), .A(n17203), .ZN(U236) );
  INV_X1 U20392 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n17231) );
  AOI22_X1 U20393 ( .A1(BUF1_REG_10__SCAN_IN), .A2(n17220), .B1(
        P1_DATAO_REG_10__SCAN_IN), .B2(n17216), .ZN(n17204) );
  OAI21_X1 U20394 ( .B1(n17231), .B2(U212), .A(n17204), .ZN(U237) );
  INV_X1 U20395 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n17229) );
  AOI22_X1 U20396 ( .A1(BUF1_REG_9__SCAN_IN), .A2(n17220), .B1(
        P1_DATAO_REG_9__SCAN_IN), .B2(n17216), .ZN(n17205) );
  OAI21_X1 U20397 ( .B1(n17229), .B2(U212), .A(n17205), .ZN(U238) );
  AOI22_X1 U20398 ( .A1(P1_DATAO_REG_8__SCAN_IN), .A2(n17216), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n17215), .ZN(n17206) );
  OAI21_X1 U20399 ( .B1(n17207), .B2(n17218), .A(n17206), .ZN(U239) );
  INV_X1 U20400 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n20006) );
  AOI22_X1 U20401 ( .A1(BUF1_REG_7__SCAN_IN), .A2(n17220), .B1(
        P1_DATAO_REG_7__SCAN_IN), .B2(n17216), .ZN(n17208) );
  OAI21_X1 U20402 ( .B1(n20006), .B2(U212), .A(n17208), .ZN(U240) );
  INV_X1 U20403 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n17227) );
  AOI22_X1 U20404 ( .A1(BUF1_REG_6__SCAN_IN), .A2(n17220), .B1(
        P1_DATAO_REG_6__SCAN_IN), .B2(n17216), .ZN(n17209) );
  OAI21_X1 U20405 ( .B1(n17227), .B2(U212), .A(n17209), .ZN(U241) );
  INV_X1 U20406 ( .A(BUF1_REG_5__SCAN_IN), .ZN(n17211) );
  AOI22_X1 U20407 ( .A1(P1_DATAO_REG_5__SCAN_IN), .A2(n17216), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n17215), .ZN(n17210) );
  OAI21_X1 U20408 ( .B1(n17211), .B2(n17218), .A(n17210), .ZN(U242) );
  INV_X1 U20409 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n17225) );
  AOI22_X1 U20410 ( .A1(BUF1_REG_4__SCAN_IN), .A2(n17220), .B1(
        P1_DATAO_REG_4__SCAN_IN), .B2(n17216), .ZN(n17212) );
  OAI21_X1 U20411 ( .B1(n17225), .B2(U212), .A(n17212), .ZN(U243) );
  INV_X1 U20412 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n17224) );
  AOI22_X1 U20413 ( .A1(BUF1_REG_3__SCAN_IN), .A2(n17220), .B1(
        P1_DATAO_REG_3__SCAN_IN), .B2(n17216), .ZN(n17213) );
  OAI21_X1 U20414 ( .B1(n17224), .B2(U212), .A(n17213), .ZN(U244) );
  AOI22_X1 U20415 ( .A1(BUF1_REG_2__SCAN_IN), .A2(n17220), .B1(
        P1_DATAO_REG_2__SCAN_IN), .B2(n17216), .ZN(n17214) );
  OAI21_X1 U20416 ( .B1(n20019), .B2(U212), .A(n17214), .ZN(U245) );
  AOI22_X1 U20417 ( .A1(P1_DATAO_REG_1__SCAN_IN), .A2(n17216), .B1(
        P2_DATAO_REG_1__SCAN_IN), .B2(n17215), .ZN(n17217) );
  OAI21_X1 U20418 ( .B1(n17219), .B2(n17218), .A(n17217), .ZN(U246) );
  INV_X1 U20419 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n17222) );
  AOI22_X1 U20420 ( .A1(BUF1_REG_0__SCAN_IN), .A2(n17220), .B1(
        P1_DATAO_REG_0__SCAN_IN), .B2(n17216), .ZN(n17221) );
  OAI21_X1 U20421 ( .B1(n17222), .B2(U212), .A(n17221), .ZN(U247) );
  INV_X1 U20422 ( .A(BUF2_REG_0__SCAN_IN), .ZN(n19033) );
  AOI22_X1 U20423 ( .A1(n17253), .A2(n17222), .B1(n19033), .B2(U215), .ZN(U251) );
  INV_X1 U20424 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n17223) );
  INV_X1 U20425 ( .A(BUF2_REG_1__SCAN_IN), .ZN(n19039) );
  AOI22_X1 U20426 ( .A1(n17253), .A2(n17223), .B1(n19039), .B2(U215), .ZN(U252) );
  INV_X1 U20427 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n19043) );
  AOI22_X1 U20428 ( .A1(n17253), .A2(n20019), .B1(n19043), .B2(U215), .ZN(U253) );
  INV_X1 U20429 ( .A(BUF2_REG_3__SCAN_IN), .ZN(n19047) );
  AOI22_X1 U20430 ( .A1(n17253), .A2(n17224), .B1(n19047), .B2(U215), .ZN(U254) );
  INV_X1 U20431 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n19051) );
  AOI22_X1 U20432 ( .A1(n17253), .A2(n17225), .B1(n19051), .B2(U215), .ZN(U255) );
  INV_X1 U20433 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n17226) );
  INV_X1 U20434 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n19055) );
  AOI22_X1 U20435 ( .A1(n17255), .A2(n17226), .B1(n19055), .B2(U215), .ZN(U256) );
  INV_X1 U20436 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n19060) );
  AOI22_X1 U20437 ( .A1(n17255), .A2(n17227), .B1(n19060), .B2(U215), .ZN(U257) );
  INV_X1 U20438 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n19064) );
  AOI22_X1 U20439 ( .A1(n17253), .A2(n20006), .B1(n19064), .B2(U215), .ZN(U258) );
  INV_X1 U20440 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n17228) );
  AOI22_X1 U20441 ( .A1(n17255), .A2(n17228), .B1(n18301), .B2(U215), .ZN(U259) );
  INV_X1 U20442 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n18303) );
  AOI22_X1 U20443 ( .A1(n17253), .A2(n17229), .B1(n18303), .B2(U215), .ZN(U260) );
  INV_X1 U20444 ( .A(BUF2_REG_10__SCAN_IN), .ZN(n17230) );
  AOI22_X1 U20445 ( .A1(n17255), .A2(n17231), .B1(n17230), .B2(U215), .ZN(U261) );
  INV_X1 U20446 ( .A(BUF2_REG_11__SCAN_IN), .ZN(n18307) );
  AOI22_X1 U20447 ( .A1(n17253), .A2(n17232), .B1(n18307), .B2(U215), .ZN(U262) );
  INV_X1 U20448 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n18309) );
  AOI22_X1 U20449 ( .A1(n17255), .A2(n17233), .B1(n18309), .B2(U215), .ZN(U263) );
  INV_X1 U20450 ( .A(BUF2_REG_13__SCAN_IN), .ZN(n18313) );
  AOI22_X1 U20451 ( .A1(n17253), .A2(n17234), .B1(n18313), .B2(U215), .ZN(U264) );
  OAI22_X1 U20452 ( .A1(U215), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n17253), .ZN(n17235) );
  INV_X1 U20453 ( .A(n17235), .ZN(U265) );
  AOI22_X1 U20454 ( .A1(n17253), .A2(n17237), .B1(n17236), .B2(U215), .ZN(U266) );
  OAI22_X1 U20455 ( .A1(U215), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n17253), .ZN(n17238) );
  INV_X1 U20456 ( .A(n17238), .ZN(U267) );
  AOI22_X1 U20457 ( .A1(n17253), .A2(n17240), .B1(n17239), .B2(U215), .ZN(U268) );
  OAI22_X1 U20458 ( .A1(U215), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n17253), .ZN(n17241) );
  INV_X1 U20459 ( .A(n17241), .ZN(U269) );
  INV_X1 U20460 ( .A(BUF2_REG_19__SCAN_IN), .ZN(n20096) );
  AOI22_X1 U20461 ( .A1(n17255), .A2(n17242), .B1(n20096), .B2(U215), .ZN(U270) );
  AOI22_X1 U20462 ( .A1(n17253), .A2(n17243), .B1(n16014), .B2(U215), .ZN(U271) );
  OAI22_X1 U20463 ( .A1(U215), .A2(P2_DATAO_REG_21__SCAN_IN), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n17253), .ZN(n17244) );
  INV_X1 U20464 ( .A(n17244), .ZN(U272) );
  INV_X1 U20465 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n17245) );
  AOI22_X1 U20466 ( .A1(n17253), .A2(n17245), .B1(n19059), .B2(U215), .ZN(U273) );
  OAI22_X1 U20467 ( .A1(U215), .A2(P2_DATAO_REG_23__SCAN_IN), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n17253), .ZN(n17246) );
  INV_X1 U20468 ( .A(n17246), .ZN(U274) );
  OAI22_X1 U20469 ( .A1(U215), .A2(P2_DATAO_REG_24__SCAN_IN), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n17255), .ZN(n17247) );
  INV_X1 U20470 ( .A(n17247), .ZN(U275) );
  OAI22_X1 U20471 ( .A1(U215), .A2(P2_DATAO_REG_25__SCAN_IN), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n17255), .ZN(n17248) );
  INV_X1 U20472 ( .A(n17248), .ZN(U276) );
  OAI22_X1 U20473 ( .A1(U215), .A2(P2_DATAO_REG_26__SCAN_IN), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n17253), .ZN(n17249) );
  INV_X1 U20474 ( .A(n17249), .ZN(U277) );
  OAI22_X1 U20475 ( .A1(U215), .A2(P2_DATAO_REG_27__SCAN_IN), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n17253), .ZN(n17250) );
  INV_X1 U20476 ( .A(n17250), .ZN(U278) );
  INV_X1 U20477 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n17251) );
  INV_X1 U20478 ( .A(BUF2_REG_28__SCAN_IN), .ZN(n20102) );
  AOI22_X1 U20479 ( .A1(n17253), .A2(n17251), .B1(n20102), .B2(U215), .ZN(U279) );
  INV_X1 U20480 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n17252) );
  AOI22_X1 U20481 ( .A1(n17253), .A2(n17252), .B1(n15938), .B2(U215), .ZN(U280) );
  INV_X1 U20482 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n17254) );
  AOI22_X1 U20483 ( .A1(n17255), .A2(n17254), .B1(n20114), .B2(U215), .ZN(U281) );
  OAI22_X1 U20484 ( .A1(U215), .A2(P2_DATAO_REG_31__SCAN_IN), .B1(
        BUF2_REG_31__SCAN_IN), .B2(n17255), .ZN(n17256) );
  INV_X1 U20485 ( .A(n17256), .ZN(U282) );
  AOI222_X1 U20486 ( .A1(n19989), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(n17257), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .C1(n18206), .C2(
        P3_DATAO_REG_30__SCAN_IN), .ZN(n17258) );
  INV_X1 U20487 ( .A(n17260), .ZN(n17259) );
  INV_X1 U20488 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n19597) );
  INV_X1 U20489 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n20647) );
  AOI22_X1 U20490 ( .A1(n17259), .A2(n19597), .B1(n20647), .B2(n17260), .ZN(
        U347) );
  INV_X1 U20491 ( .A(n17260), .ZN(n17261) );
  INV_X1 U20492 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n19595) );
  INV_X1 U20493 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n20646) );
  AOI22_X1 U20494 ( .A1(n17261), .A2(n19595), .B1(n20646), .B2(n17260), .ZN(
        U348) );
  INV_X1 U20495 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n19592) );
  INV_X1 U20496 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n20645) );
  AOI22_X1 U20497 ( .A1(n17259), .A2(n19592), .B1(n20645), .B2(n17260), .ZN(
        U349) );
  INV_X1 U20498 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n19591) );
  INV_X1 U20499 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n20644) );
  AOI22_X1 U20500 ( .A1(n17259), .A2(n19591), .B1(n20644), .B2(n17260), .ZN(
        U350) );
  INV_X1 U20501 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n19589) );
  INV_X1 U20502 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n20643) );
  AOI22_X1 U20503 ( .A1(n17259), .A2(n19589), .B1(n20643), .B2(n17260), .ZN(
        U351) );
  INV_X1 U20504 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n19587) );
  INV_X1 U20505 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n20642) );
  AOI22_X1 U20506 ( .A1(n17259), .A2(n19587), .B1(n20642), .B2(n17260), .ZN(
        U352) );
  INV_X1 U20507 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n19585) );
  INV_X1 U20508 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n20640) );
  AOI22_X1 U20509 ( .A1(n17261), .A2(n19585), .B1(n20640), .B2(n17260), .ZN(
        U353) );
  INV_X1 U20510 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n19583) );
  AOI22_X1 U20511 ( .A1(n17259), .A2(n19583), .B1(n20639), .B2(n17260), .ZN(
        U354) );
  INV_X1 U20512 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n19638) );
  INV_X1 U20513 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n20682) );
  AOI22_X1 U20514 ( .A1(n17259), .A2(n19638), .B1(n20682), .B2(n17260), .ZN(
        U355) );
  INV_X1 U20515 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n19635) );
  INV_X1 U20516 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n20679) );
  AOI22_X1 U20517 ( .A1(n17259), .A2(n19635), .B1(n20679), .B2(n17260), .ZN(
        U356) );
  INV_X1 U20518 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n19632) );
  INV_X1 U20519 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n20677) );
  AOI22_X1 U20520 ( .A1(n17259), .A2(n19632), .B1(n20677), .B2(n17260), .ZN(
        U357) );
  INV_X1 U20521 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n19631) );
  INV_X1 U20522 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n20674) );
  AOI22_X1 U20523 ( .A1(n17259), .A2(n19631), .B1(n20674), .B2(n17260), .ZN(
        U358) );
  INV_X1 U20524 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n19629) );
  INV_X1 U20525 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n20673) );
  AOI22_X1 U20526 ( .A1(n17259), .A2(n19629), .B1(n20673), .B2(n17260), .ZN(
        U359) );
  INV_X1 U20527 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n19627) );
  INV_X1 U20528 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n20671) );
  AOI22_X1 U20529 ( .A1(n17259), .A2(n19627), .B1(n20671), .B2(n17260), .ZN(
        U360) );
  INV_X1 U20530 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n19625) );
  INV_X1 U20531 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n20669) );
  AOI22_X1 U20532 ( .A1(n17259), .A2(n19625), .B1(n20669), .B2(n17260), .ZN(
        U361) );
  INV_X1 U20533 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n20667) );
  AOI22_X1 U20534 ( .A1(n17259), .A2(n19622), .B1(n20667), .B2(n17260), .ZN(
        U362) );
  INV_X1 U20535 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n19621) );
  AOI22_X1 U20536 ( .A1(n17259), .A2(n19621), .B1(n20665), .B2(n17260), .ZN(
        U363) );
  INV_X1 U20537 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n19619) );
  INV_X1 U20538 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n20664) );
  AOI22_X1 U20539 ( .A1(n17259), .A2(n19619), .B1(n20664), .B2(n17260), .ZN(
        U364) );
  INV_X1 U20540 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n19581) );
  INV_X1 U20541 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n20638) );
  AOI22_X1 U20542 ( .A1(n17259), .A2(n19581), .B1(n20638), .B2(n17260), .ZN(
        U365) );
  INV_X1 U20543 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n19616) );
  INV_X1 U20544 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n20662) );
  AOI22_X1 U20545 ( .A1(n17259), .A2(n19616), .B1(n20662), .B2(n17260), .ZN(
        U366) );
  INV_X1 U20546 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n19615) );
  INV_X1 U20547 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n20661) );
  AOI22_X1 U20548 ( .A1(n17259), .A2(n19615), .B1(n20661), .B2(n17260), .ZN(
        U367) );
  INV_X1 U20549 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n19613) );
  AOI22_X1 U20550 ( .A1(n17259), .A2(n19613), .B1(n20659), .B2(n17260), .ZN(
        U368) );
  INV_X1 U20551 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n19610) );
  AOI22_X1 U20552 ( .A1(n17259), .A2(n19610), .B1(n20657), .B2(n17260), .ZN(
        U369) );
  INV_X1 U20553 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n19609) );
  INV_X1 U20554 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n20655) );
  AOI22_X1 U20555 ( .A1(n17259), .A2(n19609), .B1(n20655), .B2(n17260), .ZN(
        U370) );
  INV_X1 U20556 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n19607) );
  INV_X1 U20557 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n20653) );
  AOI22_X1 U20558 ( .A1(n17261), .A2(n19607), .B1(n20653), .B2(n17260), .ZN(
        U371) );
  INV_X1 U20559 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n19605) );
  INV_X1 U20560 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n20652) );
  AOI22_X1 U20561 ( .A1(n17261), .A2(n19605), .B1(n20652), .B2(n17260), .ZN(
        U372) );
  INV_X1 U20562 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n19603) );
  AOI22_X1 U20563 ( .A1(n17261), .A2(n19603), .B1(n20651), .B2(n17260), .ZN(
        U373) );
  INV_X1 U20564 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n19601) );
  INV_X1 U20565 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n20650) );
  AOI22_X1 U20566 ( .A1(n17261), .A2(n19601), .B1(n20650), .B2(n17260), .ZN(
        U374) );
  INV_X1 U20567 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n19599) );
  INV_X1 U20568 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n20649) );
  AOI22_X1 U20569 ( .A1(n17261), .A2(n19599), .B1(n20649), .B2(n17260), .ZN(
        U375) );
  INV_X1 U20570 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n19579) );
  INV_X1 U20571 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n20637) );
  AOI22_X1 U20572 ( .A1(n17261), .A2(n19579), .B1(n20637), .B2(n17260), .ZN(
        U376) );
  INV_X1 U20573 ( .A(P3_ADS_N_REG_SCAN_IN), .ZN(n17262) );
  INV_X1 U20574 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n19578) );
  NAND2_X1 U20575 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(n19578), .ZN(n19569) );
  AOI22_X1 U20576 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n19569), .B1(
        P3_STATE_REG_1__SCAN_IN), .B2(n19577), .ZN(n19648) );
  INV_X1 U20577 ( .A(n19648), .ZN(n19562) );
  OAI21_X1 U20578 ( .B1(n19577), .B2(n17262), .A(n19562), .ZN(P3_U2633) );
  NOR2_X1 U20579 ( .A1(n18272), .A2(n17263), .ZN(n17267) );
  OAI21_X1 U20580 ( .B1(n17267), .B2(n18204), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n17264) );
  OAI21_X1 U20581 ( .B1(n17265), .B2(n19549), .A(n17264), .ZN(P3_U2634) );
  AOI21_X1 U20582 ( .B1(n19577), .B2(n19578), .A(P3_D_C_N_REG_SCAN_IN), .ZN(
        n17266) );
  AOI22_X1 U20583 ( .A1(n19710), .A2(P3_CODEFETCH_REG_SCAN_IN), .B1(n17266), 
        .B2(n19708), .ZN(P3_U2635) );
  NOR2_X1 U20584 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(P3_STATE_REG_2__SCAN_IN), 
        .ZN(n19563) );
  OAI21_X1 U20585 ( .B1(n19563), .B2(BS16), .A(n19648), .ZN(n19646) );
  OAI21_X1 U20586 ( .B1(n19648), .B2(n19699), .A(n19646), .ZN(P3_U2636) );
  AOI211_X1 U20587 ( .C1(n17268), .C2(n19701), .A(n17267), .B(n19479), .ZN(
        n19485) );
  NOR2_X1 U20588 ( .A1(n19485), .A2(n19546), .ZN(n19691) );
  OAI21_X1 U20589 ( .B1(n19691), .B2(n17270), .A(n17269), .ZN(P3_U2637) );
  NOR4_X1 U20590 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_20__SCAN_IN), .A3(P3_DATAWIDTH_REG_21__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_22__SCAN_IN), .ZN(n17274) );
  NOR4_X1 U20591 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_16__SCAN_IN), .A3(P3_DATAWIDTH_REG_17__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_18__SCAN_IN), .ZN(n17273) );
  NOR4_X1 U20592 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_29__SCAN_IN), .A3(P3_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_31__SCAN_IN), .ZN(n17272) );
  NOR4_X1 U20593 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_25__SCAN_IN), .A3(P3_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_27__SCAN_IN), .ZN(n17271) );
  NAND4_X1 U20594 ( .A1(n17274), .A2(n17273), .A3(n17272), .A4(n17271), .ZN(
        n17280) );
  NOR4_X1 U20595 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_4__SCAN_IN), .A3(P3_DATAWIDTH_REG_5__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_6__SCAN_IN), .ZN(n17278) );
  AOI211_X1 U20596 ( .C1(P3_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A(P3_DATAWIDTH_REG_23__SCAN_IN), .B(
        P3_DATAWIDTH_REG_2__SCAN_IN), .ZN(n17277) );
  NOR4_X1 U20597 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_12__SCAN_IN), .A3(P3_DATAWIDTH_REG_13__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_14__SCAN_IN), .ZN(n17276) );
  NOR4_X1 U20598 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_8__SCAN_IN), .A3(P3_DATAWIDTH_REG_9__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_10__SCAN_IN), .ZN(n17275) );
  NAND4_X1 U20599 ( .A1(n17278), .A2(n17277), .A3(n17276), .A4(n17275), .ZN(
        n17279) );
  NOR2_X1 U20600 ( .A1(n17280), .A2(n17279), .ZN(n19685) );
  INV_X1 U20601 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n19643) );
  INV_X1 U20602 ( .A(n19685), .ZN(n19688) );
  INV_X1 U20603 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n19681) );
  NOR2_X1 U20604 ( .A1(P3_DATAWIDTH_REG_1__SCAN_IN), .A2(n19688), .ZN(n17282)
         );
  INV_X1 U20605 ( .A(P3_REIP_REG_0__SCAN_IN), .ZN(n19687) );
  INV_X1 U20606 ( .A(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(n17281) );
  NAND3_X1 U20607 ( .A1(n17282), .A2(n19687), .A3(n17281), .ZN(n17285) );
  OAI221_X1 U20608 ( .B1(n19685), .B2(n19643), .C1(n19688), .C2(n19681), .A(
        n17285), .ZN(P3_U2638) );
  OAI21_X1 U20609 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A(n19685), .ZN(n17283) );
  OAI21_X1 U20610 ( .B1(P3_BYTEENABLE_REG_3__SCAN_IN), .B2(n19685), .A(n17283), 
        .ZN(n17284) );
  NAND2_X1 U20611 ( .A1(n17285), .A2(n17284), .ZN(P3_U2639) );
  NOR3_X1 U20612 ( .A1(P3_REIP_REG_31__SCAN_IN), .A2(n19639), .A3(n17286), 
        .ZN(n17287) );
  AOI21_X1 U20613 ( .B1(n17581), .B2(P3_EBX_REG_31__SCAN_IN), .A(n17287), .ZN(
        n17297) );
  INV_X1 U20614 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n17294) );
  NOR4_X1 U20615 ( .A1(n17289), .A2(n17288), .A3(n17576), .A4(n19555), .ZN(
        n17293) );
  INV_X1 U20616 ( .A(n17290), .ZN(n17291) );
  AOI21_X1 U20617 ( .B1(n17301), .B2(n17291), .A(n19637), .ZN(n17292) );
  AOI211_X1 U20618 ( .C1(n17295), .C2(n17294), .A(n17293), .B(n17292), .ZN(
        n17296) );
  NOR2_X1 U20619 ( .A1(n17309), .A2(n17743), .ZN(n17307) );
  AOI211_X1 U20620 ( .C1(n17300), .C2(n17299), .A(n17298), .B(n19555), .ZN(
        n17303) );
  INV_X1 U20621 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n19634) );
  OAI22_X1 U20622 ( .A1(n17301), .A2(n19634), .B1(n10042), .B2(n17586), .ZN(
        n17302) );
  AOI211_X1 U20623 ( .C1(P3_EBX_REG_29__SCAN_IN), .C2(n17581), .A(n17303), .B(
        n17302), .ZN(n17305) );
  NAND4_X1 U20624 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .A3(n17308), .A4(n19634), .ZN(n17304) );
  OAI211_X1 U20625 ( .C1(n17307), .C2(n17306), .A(n17305), .B(n17304), .ZN(
        P3_U2642) );
  NAND2_X1 U20626 ( .A1(P3_REIP_REG_27__SCAN_IN), .A2(n17308), .ZN(n17317) );
  AOI22_X1 U20627 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n17606), .B1(
        n17581), .B2(P3_EBX_REG_28__SCAN_IN), .ZN(n17316) );
  INV_X1 U20628 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n19630) );
  NAND2_X1 U20629 ( .A1(n17308), .A2(n19630), .ZN(n17328) );
  NAND2_X1 U20630 ( .A1(n17321), .A2(n17328), .ZN(n17314) );
  AOI211_X1 U20631 ( .C1(P3_EBX_REG_28__SCAN_IN), .C2(n17324), .A(n17309), .B(
        n17618), .ZN(n17313) );
  AOI211_X1 U20632 ( .C1(n18323), .C2(n17311), .A(n17310), .B(n19555), .ZN(
        n17312) );
  AOI211_X1 U20633 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(n17314), .A(n17313), 
        .B(n17312), .ZN(n17315) );
  OAI211_X1 U20634 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(n17317), .A(n17316), 
        .B(n17315), .ZN(P3_U2643) );
  AOI211_X1 U20635 ( .C1(n17320), .C2(n17319), .A(n17318), .B(n19555), .ZN(
        n17323) );
  OAI22_X1 U20636 ( .A1(n18347), .A2(n17586), .B1(n19630), .B2(n17321), .ZN(
        n17322) );
  AOI211_X1 U20637 ( .C1(n17581), .C2(P3_EBX_REG_27__SCAN_IN), .A(n17323), .B(
        n17322), .ZN(n17329) );
  OAI211_X1 U20638 ( .C1(n17326), .C2(n17325), .A(n17583), .B(n17324), .ZN(
        n17327) );
  NAND3_X1 U20639 ( .A1(n17329), .A2(n17328), .A3(n17327), .ZN(P3_U2644) );
  INV_X1 U20640 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n19624) );
  OAI21_X1 U20641 ( .B1(n17341), .B2(n17609), .A(n17459), .ZN(n17356) );
  AOI21_X1 U20642 ( .B1(n17602), .B2(n19624), .A(n17356), .ZN(n17339) );
  AOI211_X1 U20643 ( .C1(n17331), .C2(n9815), .A(n17330), .B(n19555), .ZN(
        n17334) );
  INV_X1 U20644 ( .A(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n17332) );
  OAI22_X1 U20645 ( .A1(n17737), .A2(n17619), .B1(n17332), .B2(n17586), .ZN(
        n17333) );
  AOI211_X1 U20646 ( .C1(n17335), .C2(n19626), .A(n17334), .B(n17333), .ZN(
        n17338) );
  OAI211_X1 U20647 ( .C1(n17342), .C2(n17737), .A(n17583), .B(n17336), .ZN(
        n17337) );
  OAI211_X1 U20648 ( .C1(n17339), .C2(n19626), .A(n17338), .B(n17337), .ZN(
        P3_U2646) );
  NOR2_X1 U20649 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n17609), .ZN(n17340) );
  AOI22_X1 U20650 ( .A1(n17581), .A2(P3_EBX_REG_24__SCAN_IN), .B1(n17341), 
        .B2(n17340), .ZN(n17348) );
  AOI211_X1 U20651 ( .C1(P3_EBX_REG_24__SCAN_IN), .C2(n17357), .A(n17342), .B(
        n17618), .ZN(n17346) );
  AOI211_X1 U20652 ( .C1(n18378), .C2(n17344), .A(n17343), .B(n19555), .ZN(
        n17345) );
  AOI211_X1 U20653 ( .C1(P3_REIP_REG_24__SCAN_IN), .C2(n17356), .A(n17346), 
        .B(n17345), .ZN(n17347) );
  OAI211_X1 U20654 ( .C1(n18380), .C2(n17586), .A(n17348), .B(n17347), .ZN(
        P3_U2647) );
  OR2_X1 U20655 ( .A1(n17609), .A2(n17361), .ZN(n17377) );
  OAI21_X1 U20656 ( .B1(n17349), .B2(n17377), .A(n19623), .ZN(n17355) );
  AOI211_X1 U20657 ( .C1(n18395), .C2(n17351), .A(n17350), .B(n19555), .ZN(
        n17354) );
  INV_X1 U20658 ( .A(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n17352) );
  OAI22_X1 U20659 ( .A1(n17736), .A2(n17619), .B1(n17352), .B2(n17586), .ZN(
        n17353) );
  AOI211_X1 U20660 ( .C1(n17356), .C2(n17355), .A(n17354), .B(n17353), .ZN(
        n17359) );
  OAI211_X1 U20661 ( .C1(n17362), .C2(n17736), .A(n17583), .B(n17357), .ZN(
        n17358) );
  NAND2_X1 U20662 ( .A1(n17359), .A2(n17358), .ZN(P3_U2648) );
  NOR2_X1 U20663 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(n17377), .ZN(n17360) );
  AOI22_X1 U20664 ( .A1(n17581), .A2(P3_EBX_REG_22__SCAN_IN), .B1(
        P3_REIP_REG_21__SCAN_IN), .B2(n17360), .ZN(n17368) );
  AOI21_X1 U20665 ( .B1(n17602), .B2(n17361), .A(n17621), .ZN(n17385) );
  OAI21_X1 U20666 ( .B1(P3_REIP_REG_21__SCAN_IN), .B2(n17377), .A(n17385), 
        .ZN(n17366) );
  AOI211_X1 U20667 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n17374), .A(n17362), .B(
        n17618), .ZN(n17365) );
  AOI211_X1 U20668 ( .C1(n18412), .C2(n9831), .A(n17363), .B(n19555), .ZN(
        n17364) );
  AOI211_X1 U20669 ( .C1(P3_REIP_REG_22__SCAN_IN), .C2(n17366), .A(n17365), 
        .B(n17364), .ZN(n17367) );
  OAI211_X1 U20670 ( .C1(n18414), .C2(n17586), .A(n17368), .B(n17367), .ZN(
        P3_U2649) );
  INV_X1 U20671 ( .A(n17385), .ZN(n17373) );
  AOI211_X1 U20672 ( .C1(n18425), .C2(n17370), .A(n17369), .B(n19555), .ZN(
        n17372) );
  OAI22_X1 U20673 ( .A1(n18422), .A2(n17586), .B1(n17619), .B2(n17801), .ZN(
        n17371) );
  AOI211_X1 U20674 ( .C1(n17373), .C2(P3_REIP_REG_21__SCAN_IN), .A(n17372), 
        .B(n17371), .ZN(n17376) );
  OAI211_X1 U20675 ( .C1(n17380), .C2(n17801), .A(n17583), .B(n17374), .ZN(
        n17375) );
  OAI211_X1 U20676 ( .C1(P3_REIP_REG_21__SCAN_IN), .C2(n17377), .A(n17376), 
        .B(n17375), .ZN(P3_U2650) );
  NOR3_X1 U20677 ( .A1(n17609), .A2(n19611), .A3(n17408), .ZN(n17403) );
  NAND3_X1 U20678 ( .A1(P3_REIP_REG_19__SCAN_IN), .A2(P3_REIP_REG_18__SCAN_IN), 
        .A3(n17403), .ZN(n17386) );
  INV_X1 U20679 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n19617) );
  AOI211_X1 U20680 ( .C1(n18431), .C2(n17379), .A(n17378), .B(n19555), .ZN(
        n17383) );
  AOI211_X1 U20681 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n17390), .A(n17380), .B(
        n17618), .ZN(n17382) );
  INV_X1 U20682 ( .A(P3_EBX_REG_20__SCAN_IN), .ZN(n17786) );
  OAI22_X1 U20683 ( .A1(n18409), .A2(n17586), .B1(n17619), .B2(n17786), .ZN(
        n17381) );
  NOR3_X1 U20684 ( .A1(n17383), .A2(n17382), .A3(n17381), .ZN(n17384) );
  OAI221_X1 U20685 ( .B1(P3_REIP_REG_20__SCAN_IN), .B2(n17386), .C1(n19617), 
        .C2(n17385), .A(n17384), .ZN(P3_U2651) );
  NAND2_X1 U20686 ( .A1(P3_REIP_REG_18__SCAN_IN), .A2(n17403), .ZN(n17397) );
  INV_X1 U20687 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n19614) );
  INV_X1 U20688 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n19612) );
  OAI21_X1 U20689 ( .B1(n17387), .B2(n17609), .A(n17459), .ZN(n17409) );
  AOI21_X1 U20690 ( .B1(n17403), .B2(n19612), .A(n17409), .ZN(n17396) );
  AOI211_X1 U20691 ( .C1(n18449), .C2(n17389), .A(n17388), .B(n19555), .ZN(
        n17394) );
  OAI211_X1 U20692 ( .C1(n17398), .C2(n17392), .A(n17583), .B(n17390), .ZN(
        n17391) );
  OAI211_X1 U20693 ( .C1(n17619), .C2(n17392), .A(n19013), .B(n17391), .ZN(
        n17393) );
  AOI211_X1 U20694 ( .C1(n17606), .C2(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n17394), .B(n17393), .ZN(n17395) );
  OAI221_X1 U20695 ( .B1(P3_REIP_REG_19__SCAN_IN), .B2(n17397), .C1(n19614), 
        .C2(n17396), .A(n17395), .ZN(P3_U2652) );
  AOI211_X1 U20696 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n17411), .A(n17398), .B(
        n17618), .ZN(n17399) );
  AOI211_X1 U20697 ( .C1(n17581), .C2(P3_EBX_REG_18__SCAN_IN), .A(n18866), .B(
        n17399), .ZN(n17405) );
  AOI211_X1 U20698 ( .C1(n18462), .C2(n17401), .A(n17400), .B(n19555), .ZN(
        n17402) );
  AOI221_X1 U20699 ( .B1(n17403), .B2(n19612), .C1(n17409), .C2(
        P3_REIP_REG_18__SCAN_IN), .A(n17402), .ZN(n17404) );
  OAI211_X1 U20700 ( .C1(n18459), .C2(n17586), .A(n17405), .B(n17404), .ZN(
        P3_U2653) );
  OAI21_X1 U20701 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17420), .A(
        n10033), .ZN(n17407) );
  AOI21_X1 U20702 ( .B1(n17415), .B2(n17420), .A(n17406), .ZN(n18472) );
  XOR2_X1 U20703 ( .A(n17407), .B(n18472), .Z(n17418) );
  NOR2_X1 U20704 ( .A1(n17609), .A2(n17408), .ZN(n17410) );
  OAI21_X1 U20705 ( .B1(P3_REIP_REG_17__SCAN_IN), .B2(n17410), .A(n17409), 
        .ZN(n17414) );
  OAI211_X1 U20706 ( .C1(n17422), .C2(n17412), .A(n17583), .B(n17411), .ZN(
        n17413) );
  OAI211_X1 U20707 ( .C1(n17586), .C2(n17415), .A(n17414), .B(n17413), .ZN(
        n17416) );
  AOI211_X1 U20708 ( .C1(n17581), .C2(P3_EBX_REG_17__SCAN_IN), .A(n18866), .B(
        n17416), .ZN(n17417) );
  OAI21_X1 U20709 ( .B1(n17418), .B2(n19555), .A(n17417), .ZN(P3_U2654) );
  OR2_X1 U20710 ( .A1(n17419), .A2(n17576), .ZN(n17435) );
  INV_X1 U20711 ( .A(n17433), .ZN(n17421) );
  OAI21_X1 U20712 ( .B1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n17421), .A(
        n17420), .ZN(n18487) );
  XNOR2_X1 U20713 ( .A(n17435), .B(n18487), .ZN(n17429) );
  AOI211_X1 U20714 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n17436), .A(n17422), .B(
        n17618), .ZN(n17426) );
  INV_X1 U20715 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n19608) );
  NAND3_X1 U20716 ( .A1(n17602), .A2(n17423), .A3(n19608), .ZN(n17424) );
  OAI211_X1 U20717 ( .C1(n17627), .C2(n17619), .A(n19013), .B(n17424), .ZN(
        n17425) );
  AOI211_X1 U20718 ( .C1(n17606), .C2(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n17426), .B(n17425), .ZN(n17428) );
  NOR2_X1 U20719 ( .A1(n17621), .A2(n17430), .ZN(n17448) );
  NOR2_X1 U20720 ( .A1(n17617), .A2(n17448), .ZN(n17450) );
  NOR2_X1 U20721 ( .A1(P3_REIP_REG_15__SCAN_IN), .A2(n17609), .ZN(n17431) );
  OAI21_X1 U20722 ( .B1(n17450), .B2(n17431), .A(P3_REIP_REG_16__SCAN_IN), 
        .ZN(n17427) );
  OAI211_X1 U20723 ( .C1(n19555), .C2(n17429), .A(n17428), .B(n17427), .ZN(
        P3_U2655) );
  INV_X1 U20724 ( .A(n17430), .ZN(n17432) );
  AOI22_X1 U20725 ( .A1(n17581), .A2(P3_EBX_REG_15__SCAN_IN), .B1(n17432), 
        .B2(n17431), .ZN(n17442) );
  OAI21_X1 U20726 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n18481), .A(
        n17433), .ZN(n18493) );
  NAND2_X1 U20727 ( .A1(n17608), .A2(n17576), .ZN(n17598) );
  INV_X1 U20728 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n17620) );
  OAI221_X1 U20729 ( .B1(n18493), .B2(n18481), .C1(n18493), .C2(n17620), .A(
        n17608), .ZN(n17434) );
  AOI22_X1 U20730 ( .A1(n18493), .A2(n17435), .B1(n17598), .B2(n17434), .ZN(
        n17440) );
  INV_X1 U20731 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n18496) );
  OAI211_X1 U20732 ( .C1(n17444), .C2(n17437), .A(n17583), .B(n17436), .ZN(
        n17438) );
  OAI21_X1 U20733 ( .B1(n17586), .B2(n18496), .A(n17438), .ZN(n17439) );
  AOI211_X1 U20734 ( .C1(n17450), .C2(P3_REIP_REG_15__SCAN_IN), .A(n17440), 
        .B(n17439), .ZN(n17441) );
  NAND3_X1 U20735 ( .A1(n17442), .A2(n17441), .A3(n19013), .ZN(P3_U2656) );
  INV_X1 U20736 ( .A(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n17443) );
  NAND2_X1 U20737 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18526), .ZN(
        n17472) );
  INV_X1 U20738 ( .A(n17472), .ZN(n18525) );
  NAND2_X1 U20739 ( .A1(n18524), .A2(n18525), .ZN(n17457) );
  AOI21_X1 U20740 ( .B1(n17443), .B2(n17457), .A(n18481), .ZN(n18507) );
  OAI21_X1 U20741 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17457), .A(
        n9843), .ZN(n17456) );
  XOR2_X1 U20742 ( .A(n18507), .B(n17456), .Z(n17453) );
  AOI211_X1 U20743 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n17461), .A(n17444), .B(
        n17618), .ZN(n17445) );
  AOI21_X1 U20744 ( .B1(n17606), .B2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n17445), .ZN(n17452) );
  NAND2_X1 U20745 ( .A1(n17602), .A2(n17446), .ZN(n17447) );
  INV_X1 U20746 ( .A(P3_EBX_REG_14__SCAN_IN), .ZN(n17909) );
  OAI22_X1 U20747 ( .A1(n17448), .A2(n17447), .B1(n17619), .B2(n17909), .ZN(
        n17449) );
  AOI211_X1 U20748 ( .C1(P3_REIP_REG_14__SCAN_IN), .C2(n17450), .A(n18866), 
        .B(n17449), .ZN(n17451) );
  OAI211_X1 U20749 ( .C1(n19555), .C2(n17453), .A(n17452), .B(n17451), .ZN(
        P3_U2657) );
  NOR3_X1 U20750 ( .A1(P3_REIP_REG_13__SCAN_IN), .A2(n17609), .A3(n17454), 
        .ZN(n17455) );
  AOI211_X1 U20751 ( .C1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .C2(n17606), .A(
        n18866), .B(n17455), .ZN(n17466) );
  NOR2_X1 U20752 ( .A1(n17456), .A2(n19555), .ZN(n17458) );
  NOR2_X1 U20753 ( .A1(n18542), .A2(n17472), .ZN(n17471) );
  OAI21_X1 U20754 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n17471), .A(
        n17457), .ZN(n18528) );
  AOI22_X1 U20755 ( .A1(n17581), .A2(P3_EBX_REG_13__SCAN_IN), .B1(n17458), 
        .B2(n18528), .ZN(n17465) );
  OAI21_X1 U20756 ( .B1(n17470), .B2(n17609), .A(n17459), .ZN(n17488) );
  NOR2_X1 U20757 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n17609), .ZN(n17469) );
  NOR2_X1 U20758 ( .A1(n17576), .A2(n17620), .ZN(n17607) );
  OR2_X1 U20759 ( .A1(n19555), .A2(n17607), .ZN(n17616) );
  AOI211_X1 U20760 ( .C1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .C2(n10033), .A(
        n18528), .B(n17616), .ZN(n17460) );
  AOI221_X1 U20761 ( .B1(n17488), .B2(P3_REIP_REG_13__SCAN_IN), .C1(n17469), 
        .C2(P3_REIP_REG_13__SCAN_IN), .A(n17460), .ZN(n17464) );
  OAI211_X1 U20762 ( .C1(n17467), .C2(n17462), .A(n17583), .B(n17461), .ZN(
        n17463) );
  NAND4_X1 U20763 ( .A1(n17466), .A2(n17465), .A3(n17464), .A4(n17463), .ZN(
        P3_U2658) );
  AOI22_X1 U20764 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n17606), .B1(
        n17581), .B2(P3_EBX_REG_12__SCAN_IN), .ZN(n17477) );
  AOI211_X1 U20765 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n17482), .A(n17467), .B(
        n17618), .ZN(n17468) );
  AOI211_X1 U20766 ( .C1(n17470), .C2(n17469), .A(n18866), .B(n17468), .ZN(
        n17476) );
  AOI21_X1 U20767 ( .B1(n18542), .B2(n17472), .A(n17471), .ZN(n18546) );
  NOR2_X1 U20768 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n17615), .ZN(
        n17595) );
  AOI21_X1 U20769 ( .B1(n18526), .B2(n17595), .A(n17576), .ZN(n17473) );
  XOR2_X1 U20770 ( .A(n18546), .B(n17473), .Z(n17474) );
  AOI22_X1 U20771 ( .A1(n17608), .A2(n17474), .B1(P3_REIP_REG_12__SCAN_IN), 
        .B2(n17488), .ZN(n17475) );
  NAND3_X1 U20772 ( .A1(n17477), .A2(n17476), .A3(n17475), .ZN(P3_U2659) );
  NAND3_X1 U20773 ( .A1(n17602), .A2(P3_REIP_REG_8__SCAN_IN), .A3(n17521), 
        .ZN(n17499) );
  OAI21_X1 U20774 ( .B1(n17500), .B2(n17499), .A(n19598), .ZN(n17487) );
  INV_X1 U20775 ( .A(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n17485) );
  INV_X1 U20776 ( .A(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n18555) );
  INV_X1 U20777 ( .A(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n18587) );
  NOR3_X1 U20778 ( .A1(n17615), .A2(n18618), .A3(n18619), .ZN(n17539) );
  NAND2_X1 U20779 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n17539), .ZN(
        n17531) );
  NOR3_X1 U20780 ( .A1(n17478), .A2(n18587), .A3(n17531), .ZN(n17493) );
  INV_X1 U20781 ( .A(n17493), .ZN(n17504) );
  NOR2_X1 U20782 ( .A1(n18555), .A2(n17504), .ZN(n17492) );
  INV_X1 U20783 ( .A(n17492), .ZN(n17479) );
  AOI21_X1 U20784 ( .B1(n17485), .B2(n17479), .A(n18525), .ZN(n18559) );
  AOI21_X1 U20785 ( .B1(n17492), .B2(n17620), .A(n17576), .ZN(n17481) );
  AOI21_X1 U20786 ( .B1(n18559), .B2(n17481), .A(n19555), .ZN(n17480) );
  OAI21_X1 U20787 ( .B1(n18559), .B2(n17481), .A(n17480), .ZN(n17484) );
  OAI211_X1 U20788 ( .C1(n17495), .C2(n17490), .A(n17583), .B(n17482), .ZN(
        n17483) );
  OAI211_X1 U20789 ( .C1(n17586), .C2(n17485), .A(n17484), .B(n17483), .ZN(
        n17486) );
  AOI21_X1 U20790 ( .B1(n17488), .B2(n17487), .A(n17486), .ZN(n17489) );
  OAI211_X1 U20791 ( .C1(n17619), .C2(n17490), .A(n17489), .B(n19013), .ZN(
        P3_U2660) );
  INV_X1 U20792 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n19596) );
  AOI21_X1 U20793 ( .B1(n17602), .B2(n17491), .A(n17621), .ZN(n17503) );
  AOI21_X1 U20794 ( .B1(n18555), .B2(n17504), .A(n17492), .ZN(n18566) );
  AOI21_X1 U20795 ( .B1(n17493), .B2(n17620), .A(n17576), .ZN(n17508) );
  OAI21_X1 U20796 ( .B1(n18566), .B2(n17508), .A(n17608), .ZN(n17494) );
  AOI21_X1 U20797 ( .B1(n18566), .B2(n17508), .A(n17494), .ZN(n17498) );
  AOI211_X1 U20798 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n17510), .A(n17495), .B(
        n17618), .ZN(n17497) );
  OAI22_X1 U20799 ( .A1(n18555), .A2(n17586), .B1(n17619), .B2(n17962), .ZN(
        n17496) );
  NOR4_X1 U20800 ( .A1(n18948), .A2(n17498), .A3(n17497), .A4(n17496), .ZN(
        n17502) );
  INV_X1 U20801 ( .A(n17499), .ZN(n17506) );
  OAI211_X1 U20802 ( .C1(P3_REIP_REG_10__SCAN_IN), .C2(P3_REIP_REG_9__SCAN_IN), 
        .A(n17506), .B(n17500), .ZN(n17501) );
  OAI211_X1 U20803 ( .C1(n19596), .C2(n17503), .A(n17502), .B(n17501), .ZN(
        P3_U2661) );
  INV_X1 U20804 ( .A(n17503), .ZN(n17524) );
  AOI22_X1 U20805 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n17606), .B1(
        P3_REIP_REG_9__SCAN_IN), .B2(n17524), .ZN(n17515) );
  INV_X1 U20806 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n19594) );
  NOR2_X1 U20807 ( .A1(n18587), .A2(n17531), .ZN(n17516) );
  OAI21_X1 U20808 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n17516), .A(
        n17504), .ZN(n18579) );
  OAI22_X1 U20809 ( .A1(n17619), .A2(n17511), .B1(n18579), .B2(n17598), .ZN(
        n17505) );
  AOI211_X1 U20810 ( .C1(n17506), .C2(n19594), .A(n18866), .B(n17505), .ZN(
        n17514) );
  NAND3_X1 U20811 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n17507), .A3(
        n17595), .ZN(n17517) );
  NOR2_X1 U20812 ( .A1(n18587), .A2(n17517), .ZN(n17509) );
  OAI211_X1 U20813 ( .C1(n17509), .C2(n18579), .A(n17508), .B(n17608), .ZN(
        n17513) );
  OAI211_X1 U20814 ( .C1(n17519), .C2(n17511), .A(n17583), .B(n17510), .ZN(
        n17512) );
  NAND4_X1 U20815 ( .A1(n17515), .A2(n17514), .A3(n17513), .A4(n17512), .ZN(
        P3_U2662) );
  AOI21_X1 U20816 ( .B1(n18587), .B2(n17531), .A(n17516), .ZN(n18589) );
  NAND2_X1 U20817 ( .A1(n10033), .A2(n17517), .ZN(n17518) );
  XOR2_X1 U20818 ( .A(n18589), .B(n17518), .Z(n17527) );
  AOI211_X1 U20819 ( .C1(P3_EBX_REG_8__SCAN_IN), .C2(n17528), .A(n17519), .B(
        n17618), .ZN(n17520) );
  AOI21_X1 U20820 ( .B1(P3_EBX_REG_8__SCAN_IN), .B2(n17581), .A(n17520), .ZN(
        n17526) );
  NAND2_X1 U20821 ( .A1(n17602), .A2(n17521), .ZN(n17522) );
  OAI22_X1 U20822 ( .A1(P3_REIP_REG_8__SCAN_IN), .A2(n17522), .B1(n18587), 
        .B2(n17586), .ZN(n17523) );
  AOI211_X1 U20823 ( .C1(P3_REIP_REG_8__SCAN_IN), .C2(n17524), .A(n18866), .B(
        n17523), .ZN(n17525) );
  OAI211_X1 U20824 ( .C1(n19555), .C2(n17527), .A(n17526), .B(n17525), .ZN(
        P3_U2663) );
  AOI221_X1 U20825 ( .B1(n19588), .B2(n17602), .C1(n17537), .C2(n17602), .A(
        n17621), .ZN(n17536) );
  OAI211_X1 U20826 ( .C1(n17540), .C2(n18012), .A(n17583), .B(n17528), .ZN(
        n17529) );
  OAI211_X1 U20827 ( .C1(n17619), .C2(n18012), .A(n19013), .B(n17529), .ZN(
        n17530) );
  AOI21_X1 U20828 ( .B1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n17606), .A(
        n17530), .ZN(n17535) );
  OAI21_X1 U20829 ( .B1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n17539), .A(
        n17531), .ZN(n18608) );
  AOI21_X1 U20830 ( .B1(n17507), .B2(n17595), .A(n17576), .ZN(n17541) );
  XNOR2_X1 U20831 ( .A(n18608), .B(n17541), .ZN(n17533) );
  NOR4_X1 U20832 ( .A1(P3_REIP_REG_7__SCAN_IN), .A2(n17609), .A3(n19588), .A4(
        n17537), .ZN(n17532) );
  AOI21_X1 U20833 ( .B1(n17533), .B2(n17608), .A(n17532), .ZN(n17534) );
  OAI211_X1 U20834 ( .C1(n17536), .C2(n19590), .A(n17535), .B(n17534), .ZN(
        P3_U2664) );
  AOI21_X1 U20835 ( .B1(n17602), .B2(n17537), .A(n17621), .ZN(n17552) );
  NOR3_X1 U20836 ( .A1(P3_REIP_REG_6__SCAN_IN), .A2(n17609), .A3(n17537), .ZN(
        n17538) );
  AOI211_X1 U20837 ( .C1(n17581), .C2(P3_EBX_REG_6__SCAN_IN), .A(n18866), .B(
        n17538), .ZN(n17547) );
  AOI21_X1 U20838 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n10033), .A(
        n17616), .ZN(n17545) );
  OR2_X1 U20839 ( .A1(n17615), .A2(n18618), .ZN(n17550) );
  AOI21_X1 U20840 ( .B1(n18619), .B2(n17550), .A(n17539), .ZN(n18621) );
  AOI211_X1 U20841 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n17555), .A(n17540), .B(
        n17618), .ZN(n17544) );
  NAND2_X1 U20842 ( .A1(n17608), .A2(n17541), .ZN(n17542) );
  OAI22_X1 U20843 ( .A1(n18621), .A2(n17542), .B1(n18619), .B2(n17586), .ZN(
        n17543) );
  AOI211_X1 U20844 ( .C1(n17545), .C2(n18621), .A(n17544), .B(n17543), .ZN(
        n17546) );
  OAI211_X1 U20845 ( .C1(n19588), .C2(n17552), .A(n17547), .B(n17546), .ZN(
        P3_U2665) );
  INV_X1 U20846 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n17558) );
  INV_X1 U20847 ( .A(n17548), .ZN(n17574) );
  NOR2_X1 U20848 ( .A1(n17609), .A2(n17574), .ZN(n17560) );
  AOI21_X1 U20849 ( .B1(P3_REIP_REG_4__SCAN_IN), .B2(n17560), .A(
        P3_REIP_REG_5__SCAN_IN), .ZN(n17553) );
  INV_X1 U20850 ( .A(n18630), .ZN(n17549) );
  INV_X1 U20851 ( .A(n17595), .ZN(n17563) );
  OAI21_X1 U20852 ( .B1(n17549), .B2(n17563), .A(n10033), .ZN(n17564) );
  NOR2_X1 U20853 ( .A1(n17615), .A2(n17549), .ZN(n17559) );
  OAI21_X1 U20854 ( .B1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n17559), .A(
        n17550), .ZN(n18633) );
  XNOR2_X1 U20855 ( .A(n17564), .B(n18633), .ZN(n17551) );
  OAI22_X1 U20856 ( .A1(n17553), .A2(n17552), .B1(n19555), .B2(n17551), .ZN(
        n17554) );
  AOI211_X1 U20857 ( .C1(n17581), .C2(P3_EBX_REG_5__SCAN_IN), .A(n18948), .B(
        n17554), .ZN(n17557) );
  OAI211_X1 U20858 ( .C1(n17565), .C2(n18011), .A(n17583), .B(n17555), .ZN(
        n17556) );
  OAI211_X1 U20859 ( .C1(n17586), .C2(n17558), .A(n17557), .B(n17556), .ZN(
        P3_U2666) );
  AOI21_X1 U20860 ( .B1(n17602), .B2(n17574), .A(n17621), .ZN(n17590) );
  INV_X1 U20861 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n19584) );
  INV_X1 U20862 ( .A(n17598), .ZN(n17561) );
  INV_X1 U20863 ( .A(n18636), .ZN(n17562) );
  NAND2_X1 U20864 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17562), .ZN(
        n17573) );
  AOI21_X1 U20865 ( .B1(n18650), .B2(n17573), .A(n17559), .ZN(n18647) );
  AOI22_X1 U20866 ( .A1(n17561), .A2(n18647), .B1(n17560), .B2(n19584), .ZN(
        n17572) );
  NAND2_X1 U20867 ( .A1(n17562), .A2(n18650), .ZN(n18641) );
  OAI22_X1 U20868 ( .A1(n18647), .A2(n17564), .B1(n17563), .B2(n18641), .ZN(
        n17570) );
  AOI211_X1 U20869 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n17582), .A(n17565), .B(
        n17618), .ZN(n17569) );
  NAND2_X1 U20870 ( .A1(n9751), .A2(n19715), .ZN(n17626) );
  AOI21_X1 U20871 ( .B1(n17995), .B2(n19488), .A(n17626), .ZN(n17566) );
  AOI211_X1 U20872 ( .C1(n17581), .C2(P3_EBX_REG_4__SCAN_IN), .A(n18866), .B(
        n17566), .ZN(n17567) );
  OAI21_X1 U20873 ( .B1(n18650), .B2(n17586), .A(n17567), .ZN(n17568) );
  AOI211_X1 U20874 ( .C1(n17608), .C2(n17570), .A(n17569), .B(n17568), .ZN(
        n17571) );
  OAI211_X1 U20875 ( .C1(n17590), .C2(n19584), .A(n17572), .B(n17571), .ZN(
        P3_U2667) );
  NOR2_X1 U20876 ( .A1(n18671), .A2(n17615), .ZN(n17575) );
  AOI211_X1 U20877 ( .C1(n17575), .C2(n17620), .A(n19555), .B(n17576), .ZN(
        n17594) );
  OAI21_X1 U20878 ( .B1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n17575), .A(
        n17573), .ZN(n18656) );
  NAND2_X1 U20879 ( .A1(n17602), .A2(n17574), .ZN(n17579) );
  INV_X1 U20880 ( .A(n17575), .ZN(n17593) );
  NOR2_X1 U20881 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n17593), .ZN(
        n17577) );
  OAI21_X1 U20882 ( .B1(n17577), .B2(n17576), .A(n17608), .ZN(n17578) );
  OAI22_X1 U20883 ( .A1(n17601), .A2(n17579), .B1(n18656), .B2(n17578), .ZN(
        n17588) );
  INV_X1 U20884 ( .A(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n18660) );
  OAI21_X1 U20885 ( .B1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n19497), .A(
        n17995), .ZN(n17580) );
  INV_X1 U20886 ( .A(n17580), .ZN(n19652) );
  INV_X1 U20887 ( .A(n17626), .ZN(n19717) );
  AOI22_X1 U20888 ( .A1(n17581), .A2(P3_EBX_REG_3__SCAN_IN), .B1(n19652), .B2(
        n19717), .ZN(n17585) );
  OAI211_X1 U20889 ( .C1(n17591), .C2(n18026), .A(n17583), .B(n17582), .ZN(
        n17584) );
  OAI211_X1 U20890 ( .C1(n17586), .C2(n18660), .A(n17585), .B(n17584), .ZN(
        n17587) );
  AOI211_X1 U20891 ( .C1(n17594), .C2(n18656), .A(n17588), .B(n17587), .ZN(
        n17589) );
  OAI21_X1 U20892 ( .B1(n17590), .B2(n19582), .A(n17589), .ZN(P3_U2668) );
  INV_X1 U20893 ( .A(P3_EBX_REG_0__SCAN_IN), .ZN(n18047) );
  INV_X1 U20894 ( .A(P3_EBX_REG_1__SCAN_IN), .ZN(n18041) );
  NAND2_X1 U20895 ( .A1(n18047), .A2(n18041), .ZN(n17592) );
  AOI211_X1 U20896 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n17592), .A(n17591), .B(
        n17618), .ZN(n17600) );
  OAI21_X1 U20897 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A(n17593), .ZN(n18668) );
  AOI21_X1 U20898 ( .B1(n19666), .B2(n19506), .A(n19497), .ZN(n19663) );
  AOI22_X1 U20899 ( .A1(P3_REIP_REG_2__SCAN_IN), .A2(n17621), .B1(n19663), 
        .B2(n19717), .ZN(n17597) );
  OAI21_X1 U20900 ( .B1(n17595), .B2(n18668), .A(n17594), .ZN(n17596) );
  OAI211_X1 U20901 ( .C1(n17598), .C2(n18668), .A(n17597), .B(n17596), .ZN(
        n17599) );
  AOI211_X1 U20902 ( .C1(n17606), .C2(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A(
        n17600), .B(n17599), .ZN(n17604) );
  OAI211_X1 U20903 ( .C1(P3_REIP_REG_2__SCAN_IN), .C2(P3_REIP_REG_1__SCAN_IN), 
        .A(n17602), .B(n17601), .ZN(n17603) );
  OAI211_X1 U20904 ( .C1(n17605), .C2(n17619), .A(n17604), .B(n17603), .ZN(
        P3_U2669) );
  AOI21_X1 U20905 ( .B1(n17608), .B2(n17607), .A(n17606), .ZN(n17614) );
  OAI22_X1 U20906 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n17609), .B1(n17619), 
        .B2(n18041), .ZN(n17612) );
  OAI21_X1 U20907 ( .B1(P3_EBX_REG_0__SCAN_IN), .B2(P3_EBX_REG_1__SCAN_IN), 
        .A(n18034), .ZN(n18042) );
  NAND2_X1 U20908 ( .A1(n19506), .A2(n17610), .ZN(n19667) );
  OAI22_X1 U20909 ( .A1(n17618), .A2(n18042), .B1(n19667), .B2(n17626), .ZN(
        n17611) );
  AOI211_X1 U20910 ( .C1(P3_REIP_REG_1__SCAN_IN), .C2(n17621), .A(n17612), .B(
        n17611), .ZN(n17613) );
  OAI221_X1 U20911 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n17616), .C1(
        n17615), .C2(n17614), .A(n17613), .ZN(P3_U2670) );
  INV_X1 U20912 ( .A(n17617), .ZN(n17624) );
  AOI21_X1 U20913 ( .B1(n17619), .B2(n17618), .A(n18047), .ZN(n17623) );
  NOR3_X1 U20914 ( .A1(n19713), .A2(n17621), .A3(n17620), .ZN(n17622) );
  AOI211_X1 U20915 ( .C1(P3_REIP_REG_0__SCAN_IN), .C2(n17624), .A(n17623), .B(
        n17622), .ZN(n17625) );
  OAI21_X1 U20916 ( .B1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n17626), .A(
        n17625), .ZN(P3_U2671) );
  NAND2_X1 U20917 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(P3_EBX_REG_28__SCAN_IN), 
        .ZN(n17738) );
  NAND4_X1 U20918 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(P3_EBX_REG_24__SCAN_IN), 
        .A3(P3_EBX_REG_22__SCAN_IN), .A4(P3_EBX_REG_21__SCAN_IN), .ZN(n17628)
         );
  NOR4_X1 U20919 ( .A1(n17737), .A2(n17736), .A3(n17738), .A4(n17628), .ZN(
        n17741) );
  INV_X1 U20920 ( .A(n17741), .ZN(n17629) );
  NOR4_X1 U20921 ( .A1(n17743), .A2(n17786), .A3(n17830), .A4(n17629), .ZN(
        n17734) );
  NAND2_X1 U20922 ( .A1(P3_EBX_REG_30__SCAN_IN), .A2(n17734), .ZN(n17733) );
  INV_X1 U20923 ( .A(n17733), .ZN(n17630) );
  OAI33_X1 U20924 ( .A1(P3_EBX_REG_31__SCAN_IN), .A2(n9754), .A3(n17733), .B1(
        n17631), .B2(n18045), .B3(n17630), .ZN(P3_U2672) );
  AOI22_X1 U20925 ( .A1(n17972), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17979), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n17641) );
  INV_X1 U20926 ( .A(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n19184) );
  AOI22_X1 U20927 ( .A1(n12839), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n9714), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n17633) );
  AOI22_X1 U20928 ( .A1(n17992), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n17967), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n17632) );
  OAI211_X1 U20929 ( .C1(n17975), .C2(n19184), .A(n17633), .B(n17632), .ZN(
        n17639) );
  AOI22_X1 U20930 ( .A1(n17989), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17971), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17637) );
  AOI22_X1 U20931 ( .A1(n17970), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17948), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n17636) );
  AOI22_X1 U20932 ( .A1(n17991), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12899), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n17635) );
  NAND2_X1 U20933 ( .A1(n18002), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n17634) );
  NAND4_X1 U20934 ( .A1(n17637), .A2(n17636), .A3(n17635), .A4(n17634), .ZN(
        n17638) );
  AOI211_X1 U20935 ( .C1(n17864), .C2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A(
        n17639), .B(n17638), .ZN(n17640) );
  OAI211_X1 U20936 ( .C1(n12867), .C2(n17642), .A(n17641), .B(n17640), .ZN(
        n17739) );
  AOI22_X1 U20937 ( .A1(n17971), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n12899), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n17644) );
  OAI21_X1 U20938 ( .B1(n17811), .B2(n17643), .A(n17644), .ZN(n17654) );
  AOI22_X1 U20939 ( .A1(n17970), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n12846), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n17652) );
  OAI22_X1 U20940 ( .A1(n17918), .A2(n17958), .B1(n17946), .B2(n17645), .ZN(
        n17650) );
  AOI22_X1 U20941 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n9714), .B1(
        n17948), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n17648) );
  AOI22_X1 U20942 ( .A1(n12839), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17989), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n17647) );
  AOI22_X1 U20943 ( .A1(n17864), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12840), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n17646) );
  NAND3_X1 U20944 ( .A1(n17648), .A2(n17647), .A3(n17646), .ZN(n17649) );
  AOI211_X1 U20945 ( .C1(n17979), .C2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A(
        n17650), .B(n17649), .ZN(n17651) );
  OAI211_X1 U20946 ( .C1(n17983), .C2(n17915), .A(n17652), .B(n17651), .ZN(
        n17653) );
  AOI211_X1 U20947 ( .C1(n17991), .C2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A(
        n17654), .B(n17653), .ZN(n17748) );
  AOI22_X1 U20948 ( .A1(n12899), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n9714), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n17655) );
  OAI21_X1 U20949 ( .B1(n17983), .B2(n17957), .A(n17655), .ZN(n17665) );
  AOI22_X1 U20950 ( .A1(n17972), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n9740), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17663) );
  AOI22_X1 U20951 ( .A1(n12846), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12840), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n17656) );
  OAI21_X1 U20952 ( .B1(n17966), .B2(n17947), .A(n17656), .ZN(n17661) );
  AOI22_X1 U20953 ( .A1(n17989), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17991), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n17658) );
  AOI22_X1 U20954 ( .A1(n17970), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n17967), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n17657) );
  OAI211_X1 U20955 ( .C1(n10201), .C2(n17659), .A(n17658), .B(n17657), .ZN(
        n17660) );
  AOI211_X1 U20956 ( .C1(n17979), .C2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A(
        n17661), .B(n17660), .ZN(n17662) );
  OAI211_X1 U20957 ( .C1(n17958), .C2(n19081), .A(n17663), .B(n17662), .ZN(
        n17664) );
  AOI211_X1 U20958 ( .C1(n12839), .C2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A(
        n17665), .B(n17664), .ZN(n17757) );
  AOI22_X1 U20959 ( .A1(n17967), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12899), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n17666) );
  OAI21_X1 U20960 ( .B1(n17999), .B2(n17966), .A(n17666), .ZN(n17675) );
  AOI22_X1 U20961 ( .A1(n17992), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n12846), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n17673) );
  INV_X1 U20962 ( .A(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n19167) );
  OAI22_X1 U20963 ( .A1(n17958), .A2(n19075), .B1(n17975), .B2(n19167), .ZN(
        n17671) );
  AOI22_X1 U20964 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n9714), .B1(n9740), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n17669) );
  AOI22_X1 U20965 ( .A1(n17970), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17991), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n17668) );
  AOI22_X1 U20966 ( .A1(n17979), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17864), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n17667) );
  NAND3_X1 U20967 ( .A1(n17669), .A2(n17668), .A3(n17667), .ZN(n17670) );
  AOI211_X1 U20968 ( .C1(n12839), .C2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A(
        n17671), .B(n17670), .ZN(n17672) );
  OAI211_X1 U20969 ( .C1(n12726), .C2(n17990), .A(n17673), .B(n17672), .ZN(
        n17674) );
  AOI211_X1 U20970 ( .C1(n17972), .C2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A(
        n17675), .B(n17674), .ZN(n17767) );
  INV_X1 U20971 ( .A(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n17728) );
  AOI22_X1 U20972 ( .A1(n17970), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n12899), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n17676) );
  OAI21_X1 U20973 ( .B1(n17966), .B2(n17728), .A(n17676), .ZN(n17686) );
  INV_X1 U20974 ( .A(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n17684) );
  AOI22_X1 U20975 ( .A1(n17972), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n9714), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n17683) );
  AOI22_X1 U20976 ( .A1(n17991), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12840), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n17677) );
  OAI21_X1 U20977 ( .B1(n17958), .B2(n18014), .A(n17677), .ZN(n17681) );
  INV_X1 U20978 ( .A(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n17877) );
  AOI22_X1 U20979 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n17954), .B1(
        n17989), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n17679) );
  AOI22_X1 U20980 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n17971), .B1(
        n17967), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n17678) );
  OAI211_X1 U20981 ( .C1(n10201), .C2(n17877), .A(n17679), .B(n17678), .ZN(
        n17680) );
  AOI211_X1 U20982 ( .C1(n17979), .C2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A(
        n17681), .B(n17680), .ZN(n17682) );
  OAI211_X1 U20983 ( .C1(n12867), .C2(n17684), .A(n17683), .B(n17682), .ZN(
        n17685) );
  AOI211_X1 U20984 ( .C1(n12839), .C2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A(
        n17686), .B(n17685), .ZN(n17766) );
  NOR2_X1 U20985 ( .A1(n17767), .A2(n17766), .ZN(n17762) );
  AOI22_X1 U20986 ( .A1(n12839), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n12846), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n17696) );
  AOI22_X1 U20987 ( .A1(n17970), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n17972), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n17688) );
  AOI22_X1 U20988 ( .A1(n17992), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_10__1__SCAN_IN), .B2(n12899), .ZN(n17687) );
  OAI211_X1 U20989 ( .C1(n17982), .C2(n10201), .A(n17688), .B(n17687), .ZN(
        n17694) );
  AOI22_X1 U20990 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n17967), .B1(
        P3_INSTQUEUE_REG_0__1__SCAN_IN), .B2(n17971), .ZN(n17692) );
  AOI22_X1 U20991 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n17989), .B1(
        P3_INSTQUEUE_REG_6__1__SCAN_IN), .B2(n9714), .ZN(n17691) );
  AOI22_X1 U20992 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n17948), .B1(
        n18002), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n17690) );
  NAND2_X1 U20993 ( .A1(n17991), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n17689) );
  NAND4_X1 U20994 ( .A1(n17692), .A2(n17691), .A3(n17690), .A4(n17689), .ZN(
        n17693) );
  AOI211_X1 U20995 ( .C1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .C2(n12840), .A(
        n17694), .B(n17693), .ZN(n17695) );
  OAI211_X1 U20996 ( .C1(n17976), .C2(n17995), .A(n17696), .B(n17695), .ZN(
        n17761) );
  NAND2_X1 U20997 ( .A1(n17762), .A2(n17761), .ZN(n17760) );
  NOR2_X1 U20998 ( .A1(n17757), .A2(n17760), .ZN(n17753) );
  AOI22_X1 U20999 ( .A1(n17991), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n9714), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n17706) );
  AOI22_X1 U21000 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n17989), .B1(
        n17971), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17705) );
  AOI22_X1 U21001 ( .A1(n17864), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12840), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n17704) );
  OAI22_X1 U21002 ( .A1(n17930), .A2(n17643), .B1(n12867), .B2(n17819), .ZN(
        n17702) );
  AOI22_X1 U21003 ( .A1(n17992), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17948), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n17700) );
  AOI22_X1 U21004 ( .A1(n17970), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17967), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n17699) );
  AOI22_X1 U21005 ( .A1(n12839), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n12899), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n17698) );
  NAND2_X1 U21006 ( .A1(n18002), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n17697) );
  NAND4_X1 U21007 ( .A1(n17700), .A2(n17699), .A3(n17698), .A4(n17697), .ZN(
        n17701) );
  AOI211_X1 U21008 ( .C1(n17979), .C2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A(
        n17702), .B(n17701), .ZN(n17703) );
  NAND4_X1 U21009 ( .A1(n17706), .A2(n17705), .A3(n17704), .A4(n17703), .ZN(
        n17752) );
  NAND2_X1 U21010 ( .A1(n17753), .A2(n17752), .ZN(n17751) );
  NOR2_X1 U21011 ( .A1(n17748), .A2(n17751), .ZN(n18067) );
  AOI22_X1 U21012 ( .A1(n9748), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n18002), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n17717) );
  AOI22_X1 U21013 ( .A1(n17989), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17991), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n17707) );
  OAI21_X1 U21014 ( .B1(n18021), .B2(n12838), .A(n17707), .ZN(n17715) );
  OAI22_X1 U21015 ( .A1(n12867), .A2(n17708), .B1(n12705), .B2(n17789), .ZN(
        n17709) );
  AOI21_X1 U21016 ( .B1(n12840), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A(
        n17709), .ZN(n17713) );
  AOI22_X1 U21017 ( .A1(n17970), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n9714), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n17712) );
  AOI22_X1 U21018 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n12839), .B1(
        n17954), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n17711) );
  AOI22_X1 U21019 ( .A1(n17979), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n17864), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n17710) );
  NAND4_X1 U21020 ( .A1(n17713), .A2(n17712), .A3(n17711), .A4(n17710), .ZN(
        n17714) );
  AOI211_X1 U21021 ( .C1(n17972), .C2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A(
        n17715), .B(n17714), .ZN(n17716) );
  OAI211_X1 U21022 ( .C1(n17788), .C2(n17966), .A(n17717), .B(n17716), .ZN(
        n18066) );
  NAND2_X1 U21023 ( .A1(n18067), .A2(n18066), .ZN(n18065) );
  INV_X1 U21024 ( .A(n18065), .ZN(n17718) );
  NAND2_X1 U21025 ( .A1(n17739), .A2(n17718), .ZN(n17732) );
  AOI22_X1 U21026 ( .A1(n17970), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n17948), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n17719) );
  OAI21_X1 U21027 ( .B1(n12838), .B2(n18014), .A(n17719), .ZN(n17730) );
  AOI22_X1 U21028 ( .A1(n12846), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n17979), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n17727) );
  OAI22_X1 U21029 ( .A1(n17720), .A2(n17946), .B1(n17887), .B2(n17983), .ZN(
        n17725) );
  AOI22_X1 U21030 ( .A1(n17972), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17991), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n17723) );
  AOI22_X1 U21031 ( .A1(n17989), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12899), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n17722) );
  AOI22_X1 U21032 ( .A1(n17864), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12840), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n17721) );
  NAND3_X1 U21033 ( .A1(n17723), .A2(n17722), .A3(n17721), .ZN(n17724) );
  AOI211_X1 U21034 ( .C1(n18002), .C2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A(
        n17725), .B(n17724), .ZN(n17726) );
  OAI211_X1 U21035 ( .C1(n12829), .C2(n17728), .A(n17727), .B(n17726), .ZN(
        n17729) );
  AOI211_X1 U21036 ( .C1(n12839), .C2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A(
        n17730), .B(n17729), .ZN(n17731) );
  XNOR2_X1 U21037 ( .A(n17732), .B(n17731), .ZN(n18057) );
  OAI211_X1 U21038 ( .C1(P3_EBX_REG_30__SCAN_IN), .C2(n17734), .A(n17733), .B(
        n18039), .ZN(n17735) );
  OAI21_X1 U21039 ( .B1(n18057), .B2(n18039), .A(n17735), .ZN(P3_U2673) );
  NAND2_X1 U21040 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n17770), .ZN(n17765) );
  OAI21_X1 U21041 ( .B1(n17750), .B2(n17738), .A(n18039), .ZN(n17745) );
  XNOR2_X1 U21042 ( .A(n18065), .B(n17739), .ZN(n18061) );
  NOR2_X1 U21043 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n17802), .ZN(n17740) );
  AOI22_X1 U21044 ( .A1(n18045), .A2(n18061), .B1(n17741), .B2(n17740), .ZN(
        n17742) );
  OAI21_X1 U21045 ( .B1(n17743), .B2(n17745), .A(n17742), .ZN(P3_U2674) );
  INV_X1 U21046 ( .A(n17750), .ZN(n17755) );
  NAND2_X1 U21047 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(n17755), .ZN(n17747) );
  INV_X1 U21048 ( .A(P3_EBX_REG_28__SCAN_IN), .ZN(n17746) );
  OAI211_X1 U21049 ( .C1(n18067), .C2(n18066), .A(n18045), .B(n18065), .ZN(
        n17744) );
  OAI221_X1 U21050 ( .B1(P3_EBX_REG_28__SCAN_IN), .B2(n17747), .C1(n17746), 
        .C2(n17745), .A(n17744), .ZN(P3_U2675) );
  XNOR2_X1 U21051 ( .A(n17748), .B(n17751), .ZN(n18076) );
  NAND3_X1 U21052 ( .A1(n17750), .A2(P3_EBX_REG_27__SCAN_IN), .A3(n18039), 
        .ZN(n17749) );
  OAI221_X1 U21053 ( .B1(n17750), .B2(P3_EBX_REG_27__SCAN_IN), .C1(n18039), 
        .C2(n18076), .A(n17749), .ZN(P3_U2676) );
  AOI21_X1 U21054 ( .B1(P3_EBX_REG_26__SCAN_IN), .B2(n18039), .A(n17759), .ZN(
        n17754) );
  OAI21_X1 U21055 ( .B1(n17753), .B2(n17752), .A(n17751), .ZN(n18081) );
  OAI22_X1 U21056 ( .A1(n17755), .A2(n17754), .B1(n18039), .B2(n18081), .ZN(
        P3_U2677) );
  INV_X1 U21057 ( .A(n17756), .ZN(n17764) );
  AOI21_X1 U21058 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n18039), .A(n17764), .ZN(
        n17758) );
  XNOR2_X1 U21059 ( .A(n17757), .B(n17760), .ZN(n18086) );
  OAI22_X1 U21060 ( .A1(n17759), .A2(n17758), .B1(n18039), .B2(n18086), .ZN(
        P3_U2678) );
  AOI21_X1 U21061 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n18039), .A(n17769), .ZN(
        n17763) );
  OAI21_X1 U21062 ( .B1(n17762), .B2(n17761), .A(n17760), .ZN(n18091) );
  OAI22_X1 U21063 ( .A1(n17764), .A2(n17763), .B1(n18039), .B2(n18091), .ZN(
        P3_U2679) );
  INV_X1 U21064 ( .A(n17765), .ZN(n17785) );
  AOI21_X1 U21065 ( .B1(P3_EBX_REG_23__SCAN_IN), .B2(n18039), .A(n17785), .ZN(
        n17768) );
  XNOR2_X1 U21066 ( .A(n17767), .B(n17766), .ZN(n18096) );
  OAI22_X1 U21067 ( .A1(n17769), .A2(n17768), .B1(n18039), .B2(n18096), .ZN(
        P3_U2680) );
  AOI21_X1 U21068 ( .B1(P3_EBX_REG_22__SCAN_IN), .B2(n18039), .A(n17770), .ZN(
        n17784) );
  AOI22_X1 U21069 ( .A1(n17989), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n9748), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n17771) );
  OAI21_X1 U21070 ( .B1(n12829), .B2(n19184), .A(n17771), .ZN(n17783) );
  AOI22_X1 U21071 ( .A1(n17972), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12899), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n17780) );
  INV_X1 U21072 ( .A(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n17773) );
  AOI22_X1 U21073 ( .A1(n12846), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17991), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n17772) );
  OAI21_X1 U21074 ( .B1(n10201), .B2(n17773), .A(n17772), .ZN(n17778) );
  AOI22_X1 U21075 ( .A1(n12839), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n17948), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n17775) );
  AOI22_X1 U21076 ( .A1(n17970), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n9740), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n17774) );
  OAI211_X1 U21077 ( .C1(n17995), .C2(n17776), .A(n17775), .B(n17774), .ZN(
        n17777) );
  AOI211_X1 U21078 ( .C1(n12840), .C2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A(
        n17778), .B(n17777), .ZN(n17779) );
  OAI211_X1 U21079 ( .C1(n17958), .C2(n17781), .A(n17780), .B(n17779), .ZN(
        n17782) );
  AOI211_X1 U21080 ( .C1(n17954), .C2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A(
        n17783), .B(n17782), .ZN(n18099) );
  OAI22_X1 U21081 ( .A1(n17785), .A2(n17784), .B1(n18099), .B2(n18039), .ZN(
        P3_U2681) );
  OAI21_X1 U21082 ( .B1(n17786), .B2(n17830), .A(n18039), .ZN(n17815) );
  AOI22_X1 U21083 ( .A1(n12846), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n9748), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n17798) );
  AOI22_X1 U21084 ( .A1(n17991), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n9714), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n17787) );
  OAI21_X1 U21085 ( .B1(n17788), .B2(n17643), .A(n17787), .ZN(n17796) );
  OAI22_X1 U21086 ( .A1(n18021), .A2(n17958), .B1(n12726), .B2(n17789), .ZN(
        n17790) );
  AOI21_X1 U21087 ( .B1(n12839), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A(
        n17790), .ZN(n17794) );
  AOI22_X1 U21088 ( .A1(n17971), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12899), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n17793) );
  AOI22_X1 U21089 ( .A1(n17970), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n17948), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n17792) );
  AOI22_X1 U21090 ( .A1(n17864), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12840), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n17791) );
  NAND4_X1 U21091 ( .A1(n17794), .A2(n17793), .A3(n17792), .A4(n17791), .ZN(
        n17795) );
  AOI211_X1 U21092 ( .C1(n17954), .C2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A(
        n17796), .B(n17795), .ZN(n17797) );
  OAI211_X1 U21093 ( .C1(n17799), .C2(n17995), .A(n17798), .B(n17797), .ZN(
        n18105) );
  NAND2_X1 U21094 ( .A1(n18045), .A2(n18105), .ZN(n17800) );
  OAI221_X1 U21095 ( .B1(P3_EBX_REG_21__SCAN_IN), .B2(n17802), .C1(n17801), 
        .C2(n17815), .A(n17800), .ZN(P3_U2682) );
  AOI22_X1 U21096 ( .A1(n17991), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12899), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n17803) );
  OAI21_X1 U21097 ( .B1(n17918), .B2(n17879), .A(n17803), .ZN(n17813) );
  AOI22_X1 U21098 ( .A1(n17970), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17972), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n17810) );
  INV_X1 U21099 ( .A(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n17912) );
  INV_X1 U21100 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n18027) );
  OAI22_X1 U21101 ( .A1(n17995), .A2(n17912), .B1(n17958), .B2(n18027), .ZN(
        n17808) );
  AOI22_X1 U21102 ( .A1(n17971), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n9714), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n17806) );
  AOI22_X1 U21103 ( .A1(n17992), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n17989), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n17805) );
  AOI22_X1 U21104 ( .A1(n17864), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12840), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n17804) );
  NAND3_X1 U21105 ( .A1(n17806), .A2(n17805), .A3(n17804), .ZN(n17807) );
  AOI211_X1 U21106 ( .C1(n9748), .C2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A(
        n17808), .B(n17807), .ZN(n17809) );
  OAI211_X1 U21107 ( .C1(n17811), .C2(n12867), .A(n17810), .B(n17809), .ZN(
        n17812) );
  AOI211_X1 U21108 ( .C1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .C2(n17948), .A(
        n17813), .B(n17812), .ZN(n18113) );
  NOR2_X1 U21109 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n17814), .ZN(n17816) );
  OAI22_X1 U21110 ( .A1(n18113), .A2(n18039), .B1(n17816), .B2(n17815), .ZN(
        P3_U2683) );
  AOI22_X1 U21111 ( .A1(n17967), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17971), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n17817) );
  OAI21_X1 U21112 ( .B1(n17983), .B2(n17818), .A(n17817), .ZN(n17829) );
  AOI22_X1 U21113 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n12846), .B1(
        n9714), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n17826) );
  OAI22_X1 U21114 ( .A1(n17958), .A2(n18031), .B1(n12705), .B2(n17819), .ZN(
        n17824) );
  AOI22_X1 U21115 ( .A1(n17970), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17948), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n17822) );
  AOI22_X1 U21116 ( .A1(n17972), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17989), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n17821) );
  AOI22_X1 U21117 ( .A1(n17979), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17864), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n17820) );
  NAND3_X1 U21118 ( .A1(n17822), .A2(n17821), .A3(n17820), .ZN(n17823) );
  AOI211_X1 U21119 ( .C1(n12840), .C2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A(
        n17824), .B(n17823), .ZN(n17825) );
  OAI211_X1 U21120 ( .C1(n17933), .C2(n17827), .A(n17826), .B(n17825), .ZN(
        n17828) );
  AOI211_X1 U21121 ( .C1(n12839), .C2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A(
        n17829), .B(n17828), .ZN(n18119) );
  OAI21_X1 U21122 ( .B1(P3_EBX_REG_19__SCAN_IN), .B2(n17846), .A(n17830), .ZN(
        n17831) );
  AOI22_X1 U21123 ( .A1(n18045), .A2(n18119), .B1(n17831), .B2(n18039), .ZN(
        P3_U2684) );
  OAI21_X1 U21124 ( .B1(P3_EBX_REG_18__SCAN_IN), .B2(n17832), .A(n18039), .ZN(
        n17845) );
  AOI22_X1 U21125 ( .A1(n9748), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n9714), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n17833) );
  OAI21_X1 U21126 ( .B1(n12838), .B2(n17957), .A(n17833), .ZN(n17844) );
  AOI22_X1 U21127 ( .A1(n18002), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n12899), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n17841) );
  AOI22_X1 U21128 ( .A1(n12846), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17979), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n17834) );
  OAI21_X1 U21129 ( .B1(n17643), .B2(n17947), .A(n17834), .ZN(n17839) );
  AOI22_X1 U21130 ( .A1(n12839), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n17989), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n17836) );
  AOI22_X1 U21131 ( .A1(n17991), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17948), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n17835) );
  OAI211_X1 U21132 ( .C1(n17975), .C2(n17837), .A(n17836), .B(n17835), .ZN(
        n17838) );
  AOI211_X1 U21133 ( .C1(n17864), .C2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A(
        n17839), .B(n17838), .ZN(n17840) );
  OAI211_X1 U21134 ( .C1(n17913), .C2(n17842), .A(n17841), .B(n17840), .ZN(
        n17843) );
  AOI211_X1 U21135 ( .C1(n17954), .C2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A(
        n17844), .B(n17843), .ZN(n18124) );
  OAI22_X1 U21136 ( .A1(n17846), .A2(n17845), .B1(n18124), .B2(n18039), .ZN(
        P3_U2685) );
  OAI22_X1 U21137 ( .A1(n18040), .A2(n17958), .B1(n17946), .B2(n17982), .ZN(
        n17858) );
  AOI22_X1 U21138 ( .A1(n17972), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n17948), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n17856) );
  AOI22_X1 U21139 ( .A1(n12839), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_9__1__SCAN_IN), .B2(n12899), .ZN(n17855) );
  AOI22_X1 U21140 ( .A1(n17989), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n17864), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n17847) );
  OAI21_X1 U21141 ( .B1(n12867), .B2(n17848), .A(n17847), .ZN(n17853) );
  AOI22_X1 U21142 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n17991), .B1(
        n17954), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n17850) );
  AOI22_X1 U21143 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n17970), .B1(
        P3_INSTQUEUE_REG_5__1__SCAN_IN), .B2(n9714), .ZN(n17849) );
  OAI211_X1 U21144 ( .C1(n17995), .C2(n17851), .A(n17850), .B(n17849), .ZN(
        n17852) );
  AOI211_X1 U21145 ( .C1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .C2(n12840), .A(
        n17853), .B(n17852), .ZN(n17854) );
  NAND3_X1 U21146 ( .A1(n17856), .A2(n17855), .A3(n17854), .ZN(n17857) );
  AOI211_X1 U21147 ( .C1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .C2(n17971), .A(
        n17858), .B(n17857), .ZN(n18129) );
  OAI21_X1 U21148 ( .B1(P3_EBX_REG_17__SCAN_IN), .B2(n17875), .A(n17859), .ZN(
        n17860) );
  AOI22_X1 U21149 ( .A1(n18045), .A2(n18129), .B1(n17860), .B2(n18039), .ZN(
        P3_U2686) );
  INV_X1 U21150 ( .A(n17890), .ZN(n17861) );
  OAI21_X1 U21151 ( .B1(P3_EBX_REG_16__SCAN_IN), .B2(n17861), .A(n18039), .ZN(
        n17874) );
  AOI22_X1 U21152 ( .A1(n17989), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n9748), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n17862) );
  OAI21_X1 U21153 ( .B1(n17999), .B2(n17643), .A(n17862), .ZN(n17873) );
  AOI22_X1 U21154 ( .A1(n17992), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12846), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n17871) );
  OAI22_X1 U21155 ( .A1(n17958), .A2(n17863), .B1(n12829), .B2(n19167), .ZN(
        n17869) );
  AOI22_X1 U21156 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n17948), .B1(
        n12899), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n17867) );
  AOI22_X1 U21157 ( .A1(n17991), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n9740), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n17866) );
  AOI22_X1 U21158 ( .A1(n17979), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n17864), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n17865) );
  NAND3_X1 U21159 ( .A1(n17867), .A2(n17866), .A3(n17865), .ZN(n17868) );
  AOI211_X1 U21160 ( .C1(n12840), .C2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A(
        n17869), .B(n17868), .ZN(n17870) );
  OAI211_X1 U21161 ( .C1(n17879), .C2(n19075), .A(n17871), .B(n17870), .ZN(
        n17872) );
  AOI211_X1 U21162 ( .C1(n17970), .C2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A(
        n17873), .B(n17872), .ZN(n18136) );
  OAI22_X1 U21163 ( .A1(n17875), .A2(n17874), .B1(n18136), .B2(n18039), .ZN(
        P3_U2687) );
  AOI22_X1 U21164 ( .A1(n17989), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12899), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n17876) );
  OAI21_X1 U21165 ( .B1(n17946), .B2(n17877), .A(n17876), .ZN(n17889) );
  AOI22_X1 U21166 ( .A1(n17970), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n17948), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n17886) );
  INV_X1 U21167 ( .A(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n17878) );
  OAI22_X1 U21168 ( .A1(n17879), .A2(n18014), .B1(n10201), .B2(n17878), .ZN(
        n17884) );
  AOI22_X1 U21169 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n9740), .B1(
        n17972), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n17882) );
  AOI22_X1 U21170 ( .A1(n17991), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n9714), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n17881) );
  AOI22_X1 U21171 ( .A1(n17979), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n12840), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n17880) );
  NAND3_X1 U21172 ( .A1(n17882), .A2(n17881), .A3(n17880), .ZN(n17883) );
  AOI211_X1 U21173 ( .C1(n12846), .C2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A(
        n17884), .B(n17883), .ZN(n17885) );
  OAI211_X1 U21174 ( .C1(n17887), .C2(n17958), .A(n17886), .B(n17885), .ZN(
        n17888) );
  AOI211_X1 U21175 ( .C1(n17954), .C2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A(
        n17889), .B(n17888), .ZN(n18142) );
  OAI21_X1 U21176 ( .B1(P3_EBX_REG_15__SCAN_IN), .B2(n17891), .A(n17890), .ZN(
        n17892) );
  AOI22_X1 U21177 ( .A1(n18045), .A2(n18142), .B1(n17892), .B2(n18039), .ZN(
        P3_U2688) );
  AOI22_X1 U21178 ( .A1(n12839), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n17989), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n17904) );
  AOI22_X1 U21179 ( .A1(n17991), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17948), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n17903) );
  AOI22_X1 U21180 ( .A1(n17864), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12840), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n17902) );
  OAI22_X1 U21181 ( .A1(n17958), .A2(n17894), .B1(n12838), .B2(n17893), .ZN(
        n17900) );
  AOI22_X1 U21182 ( .A1(n17992), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12899), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n17898) );
  AOI22_X1 U21183 ( .A1(n17972), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n9748), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n17897) );
  AOI22_X1 U21184 ( .A1(n12846), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n9714), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n17896) );
  NAND2_X1 U21185 ( .A1(n17979), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n17895) );
  NAND4_X1 U21186 ( .A1(n17898), .A2(n17897), .A3(n17896), .A4(n17895), .ZN(
        n17899) );
  AOI211_X1 U21187 ( .C1(n17970), .C2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A(
        n17900), .B(n17899), .ZN(n17901) );
  NAND4_X1 U21188 ( .A1(n17904), .A2(n17903), .A3(n17902), .A4(n17901), .ZN(
        n18144) );
  NOR2_X1 U21189 ( .A1(n9754), .A2(n17905), .ZN(n17906) );
  AOI22_X1 U21190 ( .A1(n18045), .A2(n18144), .B1(n17906), .B2(n17909), .ZN(
        n17907) );
  OAI21_X1 U21191 ( .B1(n17909), .B2(n17908), .A(n17907), .ZN(P3_U2689) );
  OAI21_X1 U21192 ( .B1(P3_EBX_REG_12__SCAN_IN), .B2(n17910), .A(n18039), .ZN(
        n17926) );
  AOI22_X1 U21193 ( .A1(n17992), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n9714), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n17911) );
  OAI21_X1 U21194 ( .B1(n17913), .B2(n17912), .A(n17911), .ZN(n17925) );
  AOI22_X1 U21195 ( .A1(n12846), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n9740), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n17922) );
  AOI22_X1 U21196 ( .A1(n17989), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12840), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n17914) );
  OAI21_X1 U21197 ( .B1(n17958), .B2(n17915), .A(n17914), .ZN(n17920) );
  AOI22_X1 U21198 ( .A1(n17991), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n17948), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n17917) );
  AOI22_X1 U21199 ( .A1(n12839), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n9748), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n17916) );
  OAI211_X1 U21200 ( .C1(n17918), .C2(n17995), .A(n17917), .B(n17916), .ZN(
        n17919) );
  AOI211_X1 U21201 ( .C1(n17864), .C2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A(
        n17920), .B(n17919), .ZN(n17921) );
  OAI211_X1 U21202 ( .C1(n17923), .C2(n17643), .A(n17922), .B(n17921), .ZN(
        n17924) );
  AOI211_X1 U21203 ( .C1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .C2(n12899), .A(
        n17925), .B(n17924), .ZN(n18152) );
  OAI22_X1 U21204 ( .A1(n17927), .A2(n17926), .B1(n18152), .B2(n18039), .ZN(
        P3_U2691) );
  INV_X1 U21205 ( .A(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n19175) );
  AOI22_X1 U21206 ( .A1(n17972), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n9714), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n17928) );
  OAI21_X1 U21207 ( .B1(n17966), .B2(n19175), .A(n17928), .ZN(n17940) );
  INV_X1 U21208 ( .A(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n17938) );
  AOI22_X1 U21209 ( .A1(n9748), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17991), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n17937) );
  AOI22_X1 U21210 ( .A1(n18002), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12840), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n17929) );
  OAI21_X1 U21211 ( .B1(n17930), .B2(n12705), .A(n17929), .ZN(n17935) );
  AOI22_X1 U21212 ( .A1(n12839), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n17989), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n17932) );
  AOI22_X1 U21213 ( .A1(n17970), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n9740), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n17931) );
  OAI211_X1 U21214 ( .C1(n17933), .C2(n10201), .A(n17932), .B(n17931), .ZN(
        n17934) );
  AOI211_X1 U21215 ( .C1(n17979), .C2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A(
        n17935), .B(n17934), .ZN(n17936) );
  OAI211_X1 U21216 ( .C1(n12867), .C2(n17938), .A(n17937), .B(n17936), .ZN(
        n17939) );
  AOI211_X1 U21217 ( .C1(n17954), .C2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A(
        n17940), .B(n17939), .ZN(n18155) );
  OAI21_X1 U21218 ( .B1(P3_EBX_REG_11__SCAN_IN), .B2(n17942), .A(n17941), .ZN(
        n17943) );
  AOI22_X1 U21219 ( .A1(n18045), .A2(n18155), .B1(n17943), .B2(n18039), .ZN(
        P3_U2692) );
  AOI22_X1 U21220 ( .A1(n17970), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n9740), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n17944) );
  OAI21_X1 U21221 ( .B1(n17946), .B2(n17945), .A(n17944), .ZN(n17960) );
  AOI22_X1 U21222 ( .A1(n17972), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17989), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n17956) );
  OAI22_X1 U21223 ( .A1(n12867), .A2(n17947), .B1(n17995), .B2(n19081), .ZN(
        n17953) );
  AOI22_X1 U21224 ( .A1(n17948), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n9714), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n17951) );
  AOI22_X1 U21225 ( .A1(n17991), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12899), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n17950) );
  AOI22_X1 U21226 ( .A1(n17864), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12840), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n17949) );
  NAND3_X1 U21227 ( .A1(n17951), .A2(n17950), .A3(n17949), .ZN(n17952) );
  AOI211_X1 U21228 ( .C1(n17954), .C2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A(
        n17953), .B(n17952), .ZN(n17955) );
  OAI211_X1 U21229 ( .C1(n17958), .C2(n17957), .A(n17956), .B(n17955), .ZN(
        n17959) );
  AOI211_X1 U21230 ( .C1(n12839), .C2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A(
        n17960), .B(n17959), .ZN(n18161) );
  INV_X1 U21231 ( .A(n17986), .ZN(n17961) );
  OAI33_X1 U21232 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n9754), .A3(n17986), .B1(
        n17962), .B2(n18045), .B3(n17961), .ZN(n17963) );
  INV_X1 U21233 ( .A(n17963), .ZN(n17964) );
  OAI21_X1 U21234 ( .B1(n18161), .B2(n18039), .A(n17964), .ZN(P3_U2693) );
  AOI22_X1 U21235 ( .A1(n17989), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_10__1__SCAN_IN), .B2(n17991), .ZN(n17965) );
  OAI21_X1 U21236 ( .B1(n19170), .B2(n17966), .A(n17965), .ZN(n17985) );
  AOI22_X1 U21237 ( .A1(n12839), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n12846), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n17981) );
  AOI22_X1 U21238 ( .A1(n17967), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_15__1__SCAN_IN), .B2(n18002), .ZN(n17968) );
  OAI21_X1 U21239 ( .B1(n17969), .B2(n10201), .A(n17968), .ZN(n17978) );
  AOI22_X1 U21240 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n17971), .B1(
        n17970), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n17974) );
  AOI22_X1 U21241 ( .A1(n17972), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_8__1__SCAN_IN), .B2(n12899), .ZN(n17973) );
  OAI211_X1 U21242 ( .C1(n17976), .C2(n17975), .A(n17974), .B(n17973), .ZN(
        n17977) );
  AOI211_X1 U21243 ( .C1(n17979), .C2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A(
        n17978), .B(n17977), .ZN(n17980) );
  OAI211_X1 U21244 ( .C1(n17983), .C2(n17982), .A(n17981), .B(n17980), .ZN(
        n17984) );
  AOI211_X1 U21245 ( .C1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .C2(n9714), .A(
        n17985), .B(n17984), .ZN(n18163) );
  OAI211_X1 U21246 ( .C1(P3_EBX_REG_9__SCAN_IN), .C2(n17987), .A(n17986), .B(
        n18039), .ZN(n17988) );
  OAI21_X1 U21247 ( .B1(n18163), .B2(n18039), .A(n17988), .ZN(P3_U2694) );
  AOI22_X1 U21248 ( .A1(n12839), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n9714), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n18005) );
  AOI22_X1 U21249 ( .A1(n17989), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17971), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n18004) );
  OAI22_X1 U21250 ( .A1(n10201), .A2(n17990), .B1(n17966), .B2(n19167), .ZN(
        n18001) );
  AOI22_X1 U21251 ( .A1(n17970), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n17991), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n17998) );
  AOI22_X1 U21252 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n17972), .B1(
        n12899), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n17994) );
  AOI22_X1 U21253 ( .A1(n17992), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n9748), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n17993) );
  OAI211_X1 U21254 ( .C1(n17995), .C2(n19075), .A(n17994), .B(n17993), .ZN(
        n17996) );
  AOI21_X1 U21255 ( .B1(n12840), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A(
        n17996), .ZN(n17997) );
  OAI211_X1 U21256 ( .C1(n17999), .C2(n12867), .A(n17998), .B(n17997), .ZN(
        n18000) );
  AOI211_X1 U21257 ( .C1(n18002), .C2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A(
        n18001), .B(n18000), .ZN(n18003) );
  NAND3_X1 U21258 ( .A1(n18005), .A2(n18004), .A3(n18003), .ZN(n18166) );
  AOI22_X1 U21259 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n18010), .B1(n18045), .B2(
        n18166), .ZN(n18009) );
  NAND2_X1 U21260 ( .A1(n19068), .A2(n18048), .ZN(n18043) );
  INV_X1 U21261 ( .A(n18043), .ZN(n18044) );
  OAI211_X1 U21262 ( .C1(P3_EBX_REG_8__SCAN_IN), .C2(n18007), .A(n18044), .B(
        n18006), .ZN(n18008) );
  NAND2_X1 U21263 ( .A1(n18009), .A2(n18008), .ZN(P3_U2695) );
  NOR2_X1 U21264 ( .A1(n18010), .A2(n18024), .ZN(n18020) );
  NAND2_X1 U21265 ( .A1(P3_EBX_REG_5__SCAN_IN), .A2(n18020), .ZN(n18016) );
  OAI21_X1 U21266 ( .B1(n18019), .B2(n18016), .A(P3_EBX_REG_7__SCAN_IN), .ZN(
        n18015) );
  NOR3_X1 U21267 ( .A1(n18011), .A2(n18024), .A3(n18043), .ZN(n18017) );
  NAND3_X1 U21268 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n18017), .A3(n18012), .ZN(
        n18013) );
  OAI221_X1 U21269 ( .B1(n18045), .B2(n18015), .C1(n18039), .C2(n18014), .A(
        n18013), .ZN(P3_U2696) );
  NAND2_X1 U21270 ( .A1(n18039), .A2(n18016), .ZN(n18022) );
  AOI22_X1 U21271 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n18045), .B1(
        n18017), .B2(n18019), .ZN(n18018) );
  OAI21_X1 U21272 ( .B1(n18019), .B2(n18022), .A(n18018), .ZN(P3_U2697) );
  NOR2_X1 U21273 ( .A1(P3_EBX_REG_5__SCAN_IN), .A2(n18020), .ZN(n18023) );
  OAI22_X1 U21274 ( .A1(n18023), .A2(n18022), .B1(n18021), .B2(n18039), .ZN(
        P3_U2698) );
  NOR2_X1 U21275 ( .A1(n18024), .A2(n18043), .ZN(n18029) );
  NAND2_X1 U21276 ( .A1(n18025), .A2(n18044), .ZN(n18035) );
  NOR2_X1 U21277 ( .A1(n18026), .A2(n18035), .ZN(n18033) );
  AOI21_X1 U21278 ( .B1(P3_EBX_REG_4__SCAN_IN), .B2(n18039), .A(n18033), .ZN(
        n18028) );
  OAI22_X1 U21279 ( .A1(n18029), .A2(n18028), .B1(n18027), .B2(n18039), .ZN(
        P3_U2699) );
  INV_X1 U21280 ( .A(n18035), .ZN(n18030) );
  AOI21_X1 U21281 ( .B1(P3_EBX_REG_3__SCAN_IN), .B2(n18039), .A(n18030), .ZN(
        n18032) );
  OAI22_X1 U21282 ( .A1(n18033), .A2(n18032), .B1(n18031), .B2(n18039), .ZN(
        P3_U2700) );
  INV_X1 U21283 ( .A(n18034), .ZN(n18036) );
  OAI221_X1 U21284 ( .B1(P3_EBX_REG_2__SCAN_IN), .B2(n18048), .C1(
        P3_EBX_REG_2__SCAN_IN), .C2(n18036), .A(n18035), .ZN(n18037) );
  AOI22_X1 U21285 ( .A1(n18045), .A2(n18038), .B1(n18037), .B2(n18039), .ZN(
        P3_U2701) );
  OAI222_X1 U21286 ( .A1(n18043), .A2(n18042), .B1(n18041), .B2(n18048), .C1(
        n18040), .C2(n18039), .ZN(P3_U2702) );
  AOI22_X1 U21287 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n18045), .B1(
        n18044), .B2(n18047), .ZN(n18046) );
  OAI21_X1 U21288 ( .B1(n18048), .B2(n18047), .A(n18046), .ZN(P3_U2703) );
  INV_X1 U21289 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n18211) );
  INV_X1 U21290 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n18285) );
  NAND4_X1 U21291 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(P3_EAX_REG_4__SCAN_IN), 
        .A3(P3_EAX_REG_3__SCAN_IN), .A4(P3_EAX_REG_2__SCAN_IN), .ZN(n18050) );
  NAND4_X1 U21292 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(P3_EAX_REG_6__SCAN_IN), 
        .A3(P3_EAX_REG_0__SCAN_IN), .A4(n18051), .ZN(n18167) );
  INV_X1 U21293 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n18237) );
  NAND2_X1 U21294 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(P3_EAX_REG_18__SCAN_IN), 
        .ZN(n18097) );
  NAND4_X1 U21295 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(P3_EAX_REG_20__SCAN_IN), 
        .A3(P3_EAX_REG_22__SCAN_IN), .A4(P3_EAX_REG_17__SCAN_IN), .ZN(n18052)
         );
  NAND2_X1 U21296 ( .A1(P3_EAX_REG_23__SCAN_IN), .A2(n18093), .ZN(n18092) );
  INV_X1 U21297 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n18291) );
  OR2_X1 U21298 ( .A1(n18062), .A2(n18291), .ZN(n18056) );
  NAND2_X1 U21299 ( .A1(n18053), .A2(n18114), .ZN(n18098) );
  AOI22_X1 U21300 ( .A1(BUF2_REG_31__SCAN_IN), .A2(n18130), .B1(
        P3_EAX_REG_31__SCAN_IN), .B2(n18054), .ZN(n18055) );
  OAI21_X1 U21301 ( .B1(P3_EAX_REG_31__SCAN_IN), .B2(n18056), .A(n18055), .ZN(
        P3_U2704) );
  NAND2_X1 U21302 ( .A1(n19056), .A2(n18114), .ZN(n18104) );
  OAI22_X1 U21303 ( .A1(n18057), .A2(n18186), .B1(n20114), .B2(n18098), .ZN(
        n18058) );
  AOI21_X1 U21304 ( .B1(BUF2_REG_14__SCAN_IN), .B2(n18131), .A(n18058), .ZN(
        n18059) );
  OAI221_X1 U21305 ( .B1(P3_EAX_REG_30__SCAN_IN), .B2(n18062), .C1(n18291), 
        .C2(n18060), .A(n18059), .ZN(P3_U2705) );
  AOI22_X1 U21306 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n18131), .B1(n18061), .B2(
        n18196), .ZN(n18064) );
  OAI211_X1 U21307 ( .C1(n18068), .C2(P3_EAX_REG_29__SCAN_IN), .A(n18190), .B(
        n18062), .ZN(n18063) );
  OAI211_X1 U21308 ( .C1(n18098), .C2(n15938), .A(n18064), .B(n18063), .ZN(
        P3_U2706) );
  OAI21_X1 U21309 ( .B1(n18067), .B2(n18066), .A(n18065), .ZN(n18072) );
  AOI22_X1 U21310 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n18131), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n18130), .ZN(n18071) );
  AOI211_X1 U21311 ( .C1(n18211), .C2(n18073), .A(n18068), .B(n18114), .ZN(
        n18069) );
  INV_X1 U21312 ( .A(n18069), .ZN(n18070) );
  OAI211_X1 U21313 ( .C1(n18192), .C2(n18072), .A(n18071), .B(n18070), .ZN(
        P3_U2707) );
  AOI22_X1 U21314 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n18131), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n18130), .ZN(n18075) );
  OAI211_X1 U21315 ( .C1(n18077), .C2(P3_EAX_REG_27__SCAN_IN), .A(n18190), .B(
        n18073), .ZN(n18074) );
  OAI211_X1 U21316 ( .C1(n18186), .C2(n18076), .A(n18075), .B(n18074), .ZN(
        P3_U2708) );
  AOI22_X1 U21317 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n18131), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n18130), .ZN(n18080) );
  AOI211_X1 U21318 ( .C1(n18285), .C2(n18082), .A(n18077), .B(n18114), .ZN(
        n18078) );
  INV_X1 U21319 ( .A(n18078), .ZN(n18079) );
  OAI211_X1 U21320 ( .C1(n18192), .C2(n18081), .A(n18080), .B(n18079), .ZN(
        P3_U2709) );
  AOI22_X1 U21321 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n18131), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n18130), .ZN(n18085) );
  OAI211_X1 U21322 ( .C1(n18083), .C2(P3_EAX_REG_25__SCAN_IN), .A(n18190), .B(
        n18082), .ZN(n18084) );
  OAI211_X1 U21323 ( .C1(n18192), .C2(n18086), .A(n18085), .B(n18084), .ZN(
        P3_U2710) );
  AOI22_X1 U21324 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n18131), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n18130), .ZN(n18090) );
  OAI211_X1 U21325 ( .C1(n18088), .C2(P3_EAX_REG_24__SCAN_IN), .A(n18190), .B(
        n18087), .ZN(n18089) );
  OAI211_X1 U21326 ( .C1(n18091), .C2(n18186), .A(n18090), .B(n18089), .ZN(
        P3_U2711) );
  AOI22_X1 U21327 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n18131), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n18130), .ZN(n18095) );
  OAI211_X1 U21328 ( .C1(P3_EAX_REG_23__SCAN_IN), .C2(n18093), .A(n18190), .B(
        n18092), .ZN(n18094) );
  OAI211_X1 U21329 ( .C1(n18096), .C2(n18186), .A(n18095), .B(n18094), .ZN(
        P3_U2712) );
  NAND2_X1 U21330 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n18115), .ZN(n18110) );
  NAND2_X1 U21331 ( .A1(n18190), .A2(n18110), .ZN(n18106) );
  OAI21_X1 U21332 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n18198), .A(n18106), .ZN(
        n18101) );
  OAI22_X1 U21333 ( .A1(n18099), .A2(n18186), .B1(n19059), .B2(n18098), .ZN(
        n18100) );
  AOI21_X1 U21334 ( .B1(P3_EAX_REG_22__SCAN_IN), .B2(n18101), .A(n18100), .ZN(
        n18103) );
  INV_X1 U21335 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n18222) );
  NAND4_X1 U21336 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(P3_EAX_REG_21__SCAN_IN), 
        .A3(n18115), .A4(n18222), .ZN(n18102) );
  OAI211_X1 U21337 ( .C1(n18104), .C2(n19060), .A(n18103), .B(n18102), .ZN(
        P3_U2713) );
  AOI22_X1 U21338 ( .A1(BUF2_REG_21__SCAN_IN), .A2(n18130), .B1(n18196), .B2(
        n18105), .ZN(n18109) );
  INV_X1 U21339 ( .A(n18106), .ZN(n18107) );
  AOI22_X1 U21340 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n18131), .B1(
        P3_EAX_REG_21__SCAN_IN), .B2(n18107), .ZN(n18108) );
  OAI211_X1 U21341 ( .C1(P3_EAX_REG_21__SCAN_IN), .C2(n18110), .A(n18109), .B(
        n18108), .ZN(P3_U2714) );
  AOI22_X1 U21342 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n18131), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n18130), .ZN(n18112) );
  OAI211_X1 U21343 ( .C1(n18115), .C2(P3_EAX_REG_20__SCAN_IN), .A(n18190), .B(
        n18110), .ZN(n18111) );
  OAI211_X1 U21344 ( .C1(n18113), .C2(n18186), .A(n18112), .B(n18111), .ZN(
        P3_U2715) );
  AOI22_X1 U21345 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n18131), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n18130), .ZN(n18118) );
  INV_X1 U21346 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n18228) );
  INV_X1 U21347 ( .A(n18125), .ZN(n18121) );
  NAND2_X1 U21348 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n18121), .ZN(n18120) );
  AOI211_X1 U21349 ( .C1(n18228), .C2(n18120), .A(n18115), .B(n18114), .ZN(
        n18116) );
  INV_X1 U21350 ( .A(n18116), .ZN(n18117) );
  OAI211_X1 U21351 ( .C1(n18119), .C2(n18186), .A(n18118), .B(n18117), .ZN(
        P3_U2716) );
  AOI22_X1 U21352 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n18131), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n18130), .ZN(n18123) );
  OAI211_X1 U21353 ( .C1(n18121), .C2(P3_EAX_REG_18__SCAN_IN), .A(n18190), .B(
        n18120), .ZN(n18122) );
  OAI211_X1 U21354 ( .C1(n18124), .C2(n18186), .A(n18123), .B(n18122), .ZN(
        P3_U2717) );
  AOI22_X1 U21355 ( .A1(BUF2_REG_17__SCAN_IN), .A2(n18130), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n18131), .ZN(n18128) );
  OAI211_X1 U21356 ( .C1(n18126), .C2(P3_EAX_REG_17__SCAN_IN), .A(n18190), .B(
        n18125), .ZN(n18127) );
  OAI211_X1 U21357 ( .C1(n18129), .C2(n18186), .A(n18128), .B(n18127), .ZN(
        P3_U2718) );
  AOI22_X1 U21358 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n18131), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n18130), .ZN(n18135) );
  OAI211_X1 U21359 ( .C1(P3_EAX_REG_16__SCAN_IN), .C2(n18133), .A(n18190), .B(
        n18132), .ZN(n18134) );
  OAI211_X1 U21360 ( .C1(n18136), .C2(n18186), .A(n18135), .B(n18134), .ZN(
        P3_U2719) );
  NOR2_X1 U21361 ( .A1(n9754), .A2(n18137), .ZN(n18139) );
  NAND2_X1 U21362 ( .A1(n18190), .A2(n18137), .ZN(n18146) );
  INV_X1 U21363 ( .A(n18146), .ZN(n18138) );
  MUX2_X1 U21364 ( .A(n18139), .B(n18138), .S(P3_EAX_REG_15__SCAN_IN), .Z(
        n18140) );
  AOI21_X1 U21365 ( .B1(BUF2_REG_15__SCAN_IN), .B2(n18197), .A(n18140), .ZN(
        n18141) );
  OAI21_X1 U21366 ( .B1(n18142), .B2(n18186), .A(n18141), .ZN(P3_U2720) );
  INV_X1 U21367 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n18305) );
  NOR2_X1 U21368 ( .A1(n9754), .A2(n18167), .ZN(n18173) );
  NAND3_X1 U21369 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(P3_EAX_REG_8__SCAN_IN), 
        .A3(n18173), .ZN(n18162) );
  NAND2_X1 U21370 ( .A1(P3_EAX_REG_11__SCAN_IN), .A2(n18158), .ZN(n18151) );
  NOR2_X1 U21371 ( .A1(n18242), .A2(n18151), .ZN(n18154) );
  NAND2_X1 U21372 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n18154), .ZN(n18147) );
  INV_X1 U21373 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n18316) );
  AOI22_X1 U21374 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n18197), .B1(n18196), .B2(
        n18144), .ZN(n18145) );
  OAI221_X1 U21375 ( .B1(P3_EAX_REG_14__SCAN_IN), .B2(n18147), .C1(n18316), 
        .C2(n18146), .A(n18145), .ZN(P3_U2721) );
  INV_X1 U21376 ( .A(n18147), .ZN(n18150) );
  AOI21_X1 U21377 ( .B1(P3_EAX_REG_13__SCAN_IN), .B2(n18190), .A(n18154), .ZN(
        n18149) );
  OAI222_X1 U21378 ( .A1(n18195), .A2(n18313), .B1(n18150), .B2(n18149), .C1(
        n18192), .C2(n18148), .ZN(P3_U2722) );
  INV_X1 U21379 ( .A(n18151), .ZN(n18157) );
  AOI21_X1 U21380 ( .B1(P3_EAX_REG_12__SCAN_IN), .B2(n18190), .A(n18157), .ZN(
        n18153) );
  OAI222_X1 U21381 ( .A1(n18195), .A2(n18309), .B1(n18154), .B2(n18153), .C1(
        n18192), .C2(n18152), .ZN(P3_U2723) );
  AOI21_X1 U21382 ( .B1(P3_EAX_REG_11__SCAN_IN), .B2(n18190), .A(n18158), .ZN(
        n18156) );
  OAI222_X1 U21383 ( .A1(n18195), .A2(n18307), .B1(n18157), .B2(n18156), .C1(
        n18192), .C2(n18155), .ZN(P3_U2724) );
  AOI21_X1 U21384 ( .B1(n18305), .B2(n18162), .A(n18158), .ZN(n18159) );
  AOI22_X1 U21385 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n18197), .B1(n18159), .B2(
        n18190), .ZN(n18160) );
  OAI21_X1 U21386 ( .B1(n18161), .B2(n18186), .A(n18160), .ZN(P3_U2725) );
  INV_X1 U21387 ( .A(n18162), .ZN(n18165) );
  AOI22_X1 U21388 ( .A1(n18173), .A2(P3_EAX_REG_8__SCAN_IN), .B1(
        P3_EAX_REG_9__SCAN_IN), .B2(n18190), .ZN(n18164) );
  OAI222_X1 U21389 ( .A1(n18195), .A2(n18303), .B1(n18165), .B2(n18164), .C1(
        n18192), .C2(n18163), .ZN(P3_U2726) );
  INV_X1 U21390 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n18249) );
  AOI22_X1 U21391 ( .A1(n18196), .A2(n18166), .B1(n18173), .B2(n18249), .ZN(
        n18169) );
  NAND3_X1 U21392 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n18190), .A3(n18167), .ZN(
        n18168) );
  OAI211_X1 U21393 ( .C1(n18195), .C2(n18301), .A(n18169), .B(n18168), .ZN(
        P3_U2727) );
  INV_X1 U21394 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n18253) );
  INV_X1 U21395 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n18257) );
  INV_X1 U21396 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n18170) );
  NOR3_X1 U21397 ( .A1(n18170), .A2(n18270), .A3(n18198), .ZN(n18189) );
  NAND2_X1 U21398 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n18194), .ZN(n18181) );
  NOR2_X1 U21399 ( .A1(n18257), .A2(n18181), .ZN(n18184) );
  NAND2_X1 U21400 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n18184), .ZN(n18174) );
  NOR2_X1 U21401 ( .A1(n18253), .A2(n18174), .ZN(n18177) );
  AOI21_X1 U21402 ( .B1(P3_EAX_REG_7__SCAN_IN), .B2(n18190), .A(n18177), .ZN(
        n18172) );
  OAI222_X1 U21403 ( .A1(n19064), .A2(n18195), .B1(n18173), .B2(n18172), .C1(
        n18192), .C2(n18171), .ZN(P3_U2728) );
  INV_X1 U21404 ( .A(n18174), .ZN(n18180) );
  AOI21_X1 U21405 ( .B1(P3_EAX_REG_6__SCAN_IN), .B2(n18190), .A(n18180), .ZN(
        n18176) );
  OAI222_X1 U21406 ( .A1(n19060), .A2(n18195), .B1(n18177), .B2(n18176), .C1(
        n18192), .C2(n18175), .ZN(P3_U2729) );
  AOI21_X1 U21407 ( .B1(P3_EAX_REG_5__SCAN_IN), .B2(n18190), .A(n18184), .ZN(
        n18179) );
  OAI222_X1 U21408 ( .A1(n19055), .A2(n18195), .B1(n18180), .B2(n18179), .C1(
        n18192), .C2(n18178), .ZN(P3_U2730) );
  INV_X1 U21409 ( .A(n18181), .ZN(n18188) );
  AOI21_X1 U21410 ( .B1(P3_EAX_REG_4__SCAN_IN), .B2(n18190), .A(n18188), .ZN(
        n18183) );
  OAI222_X1 U21411 ( .A1(n19051), .A2(n18195), .B1(n18184), .B2(n18183), .C1(
        n18186), .C2(n18182), .ZN(P3_U2731) );
  AOI21_X1 U21412 ( .B1(P3_EAX_REG_3__SCAN_IN), .B2(n18190), .A(n18194), .ZN(
        n18187) );
  OAI222_X1 U21413 ( .A1(n19047), .A2(n18195), .B1(n18188), .B2(n18187), .C1(
        n18186), .C2(n18185), .ZN(P3_U2732) );
  AOI21_X1 U21414 ( .B1(P3_EAX_REG_2__SCAN_IN), .B2(n18190), .A(n18189), .ZN(
        n18193) );
  OAI222_X1 U21415 ( .A1(n19043), .A2(n18195), .B1(n18194), .B2(n18193), .C1(
        n18192), .C2(n18191), .ZN(P3_U2733) );
  AOI22_X1 U21416 ( .A1(n18197), .A2(BUF2_REG_1__SCAN_IN), .B1(n18196), .B2(
        n9895), .ZN(n18203) );
  NOR2_X1 U21417 ( .A1(n18270), .A2(n18198), .ZN(n18201) );
  NOR2_X1 U21418 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(n18198), .ZN(n18200) );
  OAI22_X1 U21419 ( .A1(P3_EAX_REG_1__SCAN_IN), .A2(n18201), .B1(n18200), .B2(
        n18199), .ZN(n18202) );
  NAND2_X1 U21420 ( .A1(n18203), .A2(n18202), .ZN(P3_U2734) );
  OR2_X1 U21421 ( .A1(n19660), .A2(n19560), .ZN(n19695) );
  INV_X1 U21423 ( .A(n18204), .ZN(n18271) );
  NOR2_X1 U21424 ( .A1(n18206), .A2(n18264), .ZN(P3_U2736) );
  NAND2_X1 U21425 ( .A1(n18262), .A2(n9752), .ZN(n18232) );
  AOI22_X1 U21426 ( .A1(n19548), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(n18266), 
        .B2(P3_DATAO_REG_30__SCAN_IN), .ZN(n18207) );
  OAI21_X1 U21427 ( .B1(n18291), .B2(n18232), .A(n18207), .ZN(P3_U2737) );
  INV_X1 U21428 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n18209) );
  AOI22_X1 U21429 ( .A1(n19548), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n18266), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n18208) );
  OAI21_X1 U21430 ( .B1(n18209), .B2(n18232), .A(n18208), .ZN(P3_U2738) );
  AOI22_X1 U21431 ( .A1(n19548), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n18266), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n18210) );
  OAI21_X1 U21432 ( .B1(n18211), .B2(n18232), .A(n18210), .ZN(P3_U2739) );
  INV_X1 U21433 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n18213) );
  AOI22_X1 U21435 ( .A1(n19548), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n18266), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n18212) );
  OAI21_X1 U21436 ( .B1(n18213), .B2(n18232), .A(n18212), .ZN(P3_U2740) );
  AOI22_X1 U21437 ( .A1(n19548), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n18266), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n18214) );
  OAI21_X1 U21438 ( .B1(n18285), .B2(n18232), .A(n18214), .ZN(P3_U2741) );
  INV_X1 U21439 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n18216) );
  AOI22_X1 U21440 ( .A1(n19548), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n18266), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n18215) );
  OAI21_X1 U21441 ( .B1(n18216), .B2(n18232), .A(n18215), .ZN(P3_U2742) );
  INV_X1 U21442 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n18218) );
  AOI22_X1 U21443 ( .A1(n19548), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n18266), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n18217) );
  OAI21_X1 U21444 ( .B1(n18218), .B2(n18232), .A(n18217), .ZN(P3_U2743) );
  INV_X1 U21445 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n18220) );
  AOI22_X1 U21446 ( .A1(n19548), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n18266), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n18219) );
  OAI21_X1 U21447 ( .B1(n18220), .B2(n18232), .A(n18219), .ZN(P3_U2744) );
  AOI22_X1 U21448 ( .A1(P3_UWORD_REG_6__SCAN_IN), .A2(n19548), .B1(n18266), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n18221) );
  OAI21_X1 U21449 ( .B1(n18222), .B2(n18232), .A(n18221), .ZN(P3_U2745) );
  INV_X1 U21450 ( .A(n18232), .ZN(n18233) );
  AOI22_X1 U21451 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(n18233), .B1(n18266), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n18223) );
  OAI21_X1 U21452 ( .B1(n18224), .B2(n19695), .A(n18223), .ZN(P3_U2746) );
  INV_X1 U21453 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n18226) );
  AOI22_X1 U21454 ( .A1(n19548), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n18266), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n18225) );
  OAI21_X1 U21455 ( .B1(n18226), .B2(n18232), .A(n18225), .ZN(P3_U2747) );
  AOI22_X1 U21456 ( .A1(n19548), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n18266), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n18227) );
  OAI21_X1 U21457 ( .B1(n18228), .B2(n18232), .A(n18227), .ZN(P3_U2748) );
  INV_X1 U21458 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n18230) );
  INV_X2 U21459 ( .A(n18264), .ZN(n18266) );
  AOI22_X1 U21460 ( .A1(n19548), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n18266), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n18229) );
  OAI21_X1 U21461 ( .B1(n18230), .B2(n18232), .A(n18229), .ZN(P3_U2749) );
  INV_X1 U21462 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n18275) );
  AOI22_X1 U21463 ( .A1(n19548), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n18266), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n18231) );
  OAI21_X1 U21464 ( .B1(n18275), .B2(n18232), .A(n18231), .ZN(P3_U2750) );
  AOI22_X1 U21465 ( .A1(P3_EAX_REG_16__SCAN_IN), .A2(n18233), .B1(n19548), 
        .B2(P3_UWORD_REG_0__SCAN_IN), .ZN(n18234) );
  OAI21_X1 U21466 ( .B1(n18235), .B2(n18264), .A(n18234), .ZN(P3_U2751) );
  AOI22_X1 U21467 ( .A1(n19548), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n18266), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n18236) );
  OAI21_X1 U21468 ( .B1(n18237), .B2(n18269), .A(n18236), .ZN(P3_U2752) );
  AOI22_X1 U21469 ( .A1(n19548), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n18266), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n18238) );
  OAI21_X1 U21470 ( .B1(n18316), .B2(n18269), .A(n18238), .ZN(P3_U2753) );
  AOI22_X1 U21471 ( .A1(n19548), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n18266), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n18239) );
  OAI21_X1 U21472 ( .B1(n18240), .B2(n18269), .A(n18239), .ZN(P3_U2754) );
  AOI22_X1 U21473 ( .A1(n19548), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n18266), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n18241) );
  OAI21_X1 U21474 ( .B1(n18242), .B2(n18269), .A(n18241), .ZN(P3_U2755) );
  INV_X1 U21475 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n18244) );
  AOI22_X1 U21476 ( .A1(n19548), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n18266), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n18243) );
  OAI21_X1 U21477 ( .B1(n18244), .B2(n18269), .A(n18243), .ZN(P3_U2756) );
  AOI22_X1 U21478 ( .A1(n19548), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n18266), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n18245) );
  OAI21_X1 U21479 ( .B1(n18305), .B2(n18269), .A(n18245), .ZN(P3_U2757) );
  INV_X1 U21480 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n18247) );
  AOI22_X1 U21481 ( .A1(n19548), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n18266), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n18246) );
  OAI21_X1 U21482 ( .B1(n18247), .B2(n18269), .A(n18246), .ZN(P3_U2758) );
  AOI22_X1 U21483 ( .A1(n19548), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n18266), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n18248) );
  OAI21_X1 U21484 ( .B1(n18249), .B2(n18269), .A(n18248), .ZN(P3_U2759) );
  INV_X1 U21485 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n18251) );
  AOI22_X1 U21486 ( .A1(n19548), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n18266), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n18250) );
  OAI21_X1 U21487 ( .B1(n18251), .B2(n18269), .A(n18250), .ZN(P3_U2760) );
  AOI22_X1 U21488 ( .A1(n19548), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n18266), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n18252) );
  OAI21_X1 U21489 ( .B1(n18253), .B2(n18269), .A(n18252), .ZN(P3_U2761) );
  INV_X1 U21490 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n18255) );
  AOI22_X1 U21491 ( .A1(n19548), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n18266), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n18254) );
  OAI21_X1 U21492 ( .B1(n18255), .B2(n18269), .A(n18254), .ZN(P3_U2762) );
  AOI22_X1 U21493 ( .A1(n19548), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n18266), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n18256) );
  OAI21_X1 U21494 ( .B1(n18257), .B2(n18269), .A(n18256), .ZN(P3_U2763) );
  INV_X1 U21495 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n18259) );
  AOI22_X1 U21496 ( .A1(n19548), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n18266), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n18258) );
  OAI21_X1 U21497 ( .B1(n18259), .B2(n18269), .A(n18258), .ZN(P3_U2764) );
  INV_X1 U21498 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n18261) );
  AOI22_X1 U21499 ( .A1(n19548), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n18266), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n18260) );
  OAI21_X1 U21500 ( .B1(n18261), .B2(n18269), .A(n18260), .ZN(P3_U2765) );
  AOI22_X1 U21501 ( .A1(P3_EAX_REG_1__SCAN_IN), .A2(n18262), .B1(n19548), .B2(
        P3_LWORD_REG_1__SCAN_IN), .ZN(n18263) );
  OAI21_X1 U21502 ( .B1(n18265), .B2(n18264), .A(n18263), .ZN(P3_U2766) );
  AOI22_X1 U21503 ( .A1(n19548), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n18266), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n18268) );
  OAI21_X1 U21504 ( .B1(n18270), .B2(n18269), .A(n18268), .ZN(P3_U2767) );
  OAI211_X1 U21505 ( .C1(n19701), .C2(n19040), .A(n18272), .B(n18271), .ZN(
        n18289) );
  NOR2_X1 U21506 ( .A1(n18318), .A2(n19040), .ZN(n18317) );
  NAND3_X1 U21507 ( .A1(n19040), .A2(n18272), .A3(n18271), .ZN(n18315) );
  AOI22_X1 U21508 ( .A1(P3_EAX_REG_16__SCAN_IN), .A2(n18310), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n18318), .ZN(n18273) );
  OAI21_X1 U21509 ( .B1(n19033), .B2(n18312), .A(n18273), .ZN(P3_U2768) );
  AOI22_X1 U21510 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n18317), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n18318), .ZN(n18274) );
  OAI21_X1 U21511 ( .B1(n18275), .B2(n18315), .A(n18274), .ZN(P3_U2769) );
  AOI22_X1 U21512 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n18310), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n18289), .ZN(n18276) );
  OAI21_X1 U21513 ( .B1(n19043), .B2(n18312), .A(n18276), .ZN(P3_U2770) );
  AOI22_X1 U21514 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(n18310), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n18289), .ZN(n18277) );
  OAI21_X1 U21515 ( .B1(n19047), .B2(n18312), .A(n18277), .ZN(P3_U2771) );
  AOI22_X1 U21516 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n18310), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n18289), .ZN(n18278) );
  OAI21_X1 U21517 ( .B1(n19051), .B2(n18312), .A(n18278), .ZN(P3_U2772) );
  AOI22_X1 U21518 ( .A1(P3_UWORD_REG_5__SCAN_IN), .A2(n18318), .B1(
        P3_EAX_REG_21__SCAN_IN), .B2(n18310), .ZN(n18279) );
  OAI21_X1 U21519 ( .B1(n19055), .B2(n18312), .A(n18279), .ZN(P3_U2773) );
  AOI22_X1 U21520 ( .A1(P3_UWORD_REG_6__SCAN_IN), .A2(n18318), .B1(
        P3_EAX_REG_22__SCAN_IN), .B2(n18310), .ZN(n18280) );
  OAI21_X1 U21521 ( .B1(n19060), .B2(n18312), .A(n18280), .ZN(P3_U2774) );
  AOI22_X1 U21522 ( .A1(P3_EAX_REG_23__SCAN_IN), .A2(n18310), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n18289), .ZN(n18281) );
  OAI21_X1 U21523 ( .B1(n19064), .B2(n18312), .A(n18281), .ZN(P3_U2775) );
  AOI22_X1 U21524 ( .A1(P3_EAX_REG_24__SCAN_IN), .A2(n18310), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n18289), .ZN(n18282) );
  OAI21_X1 U21525 ( .B1(n18301), .B2(n18312), .A(n18282), .ZN(P3_U2776) );
  AOI22_X1 U21526 ( .A1(P3_EAX_REG_25__SCAN_IN), .A2(n18310), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n18289), .ZN(n18283) );
  OAI21_X1 U21527 ( .B1(n18303), .B2(n18312), .A(n18283), .ZN(P3_U2777) );
  AOI22_X1 U21528 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n18317), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n18318), .ZN(n18284) );
  OAI21_X1 U21529 ( .B1(n18285), .B2(n18315), .A(n18284), .ZN(P3_U2778) );
  AOI22_X1 U21530 ( .A1(P3_EAX_REG_27__SCAN_IN), .A2(n18310), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n18289), .ZN(n18286) );
  OAI21_X1 U21531 ( .B1(n18307), .B2(n18312), .A(n18286), .ZN(P3_U2779) );
  AOI22_X1 U21532 ( .A1(P3_EAX_REG_28__SCAN_IN), .A2(n18310), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n18289), .ZN(n18287) );
  OAI21_X1 U21533 ( .B1(n18309), .B2(n18312), .A(n18287), .ZN(P3_U2780) );
  AOI22_X1 U21534 ( .A1(P3_EAX_REG_29__SCAN_IN), .A2(n18310), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n18289), .ZN(n18288) );
  OAI21_X1 U21535 ( .B1(n18313), .B2(n18312), .A(n18288), .ZN(P3_U2781) );
  AOI22_X1 U21536 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n18317), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n18289), .ZN(n18290) );
  OAI21_X1 U21537 ( .B1(n18291), .B2(n18315), .A(n18290), .ZN(P3_U2782) );
  AOI22_X1 U21538 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(n18310), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n18318), .ZN(n18292) );
  OAI21_X1 U21539 ( .B1(n19033), .B2(n18312), .A(n18292), .ZN(P3_U2783) );
  AOI22_X1 U21540 ( .A1(P3_EAX_REG_1__SCAN_IN), .A2(n18310), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n18318), .ZN(n18293) );
  OAI21_X1 U21541 ( .B1(n19039), .B2(n18312), .A(n18293), .ZN(P3_U2784) );
  AOI22_X1 U21542 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(n18310), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n18318), .ZN(n18294) );
  OAI21_X1 U21543 ( .B1(n19043), .B2(n18312), .A(n18294), .ZN(P3_U2785) );
  AOI22_X1 U21544 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n18310), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n18318), .ZN(n18295) );
  OAI21_X1 U21545 ( .B1(n19047), .B2(n18312), .A(n18295), .ZN(P3_U2786) );
  AOI22_X1 U21546 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(n18310), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n18318), .ZN(n18296) );
  OAI21_X1 U21547 ( .B1(n19051), .B2(n18312), .A(n18296), .ZN(P3_U2787) );
  AOI22_X1 U21548 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n18310), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n18318), .ZN(n18297) );
  OAI21_X1 U21549 ( .B1(n19055), .B2(n18312), .A(n18297), .ZN(P3_U2788) );
  AOI22_X1 U21550 ( .A1(P3_EAX_REG_6__SCAN_IN), .A2(n18310), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n18318), .ZN(n18298) );
  OAI21_X1 U21551 ( .B1(n19060), .B2(n18312), .A(n18298), .ZN(P3_U2789) );
  AOI22_X1 U21552 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(n18310), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n18318), .ZN(n18299) );
  OAI21_X1 U21553 ( .B1(n19064), .B2(n18312), .A(n18299), .ZN(P3_U2790) );
  AOI22_X1 U21554 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n18310), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n18318), .ZN(n18300) );
  OAI21_X1 U21555 ( .B1(n18301), .B2(n18312), .A(n18300), .ZN(P3_U2791) );
  AOI22_X1 U21556 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(n18310), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n18318), .ZN(n18302) );
  OAI21_X1 U21557 ( .B1(n18303), .B2(n18312), .A(n18302), .ZN(P3_U2792) );
  AOI22_X1 U21558 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n18317), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n18318), .ZN(n18304) );
  OAI21_X1 U21559 ( .B1(n18305), .B2(n18315), .A(n18304), .ZN(P3_U2793) );
  AOI22_X1 U21560 ( .A1(P3_EAX_REG_11__SCAN_IN), .A2(n18310), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n18318), .ZN(n18306) );
  OAI21_X1 U21561 ( .B1(n18307), .B2(n18312), .A(n18306), .ZN(P3_U2794) );
  AOI22_X1 U21562 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n18310), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n18318), .ZN(n18308) );
  OAI21_X1 U21563 ( .B1(n18309), .B2(n18312), .A(n18308), .ZN(P3_U2795) );
  AOI22_X1 U21564 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n18310), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n18318), .ZN(n18311) );
  OAI21_X1 U21565 ( .B1(n18313), .B2(n18312), .A(n18311), .ZN(P3_U2796) );
  AOI22_X1 U21566 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n18317), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n18318), .ZN(n18314) );
  OAI21_X1 U21567 ( .B1(n18316), .B2(n18315), .A(n18314), .ZN(P3_U2797) );
  AOI222_X1 U21568 ( .A1(n18310), .A2(P3_EAX_REG_15__SCAN_IN), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n18318), .C1(BUF2_REG_15__SCAN_IN), 
        .C2(n18317), .ZN(n18319) );
  INV_X1 U21569 ( .A(n18319), .ZN(P3_U2798) );
  INV_X1 U21570 ( .A(n18336), .ZN(n18320) );
  OAI21_X1 U21571 ( .B1(n18320), .B2(n19023), .A(n18684), .ZN(n18321) );
  AOI21_X1 U21572 ( .B1(n18445), .B2(n18322), .A(n18321), .ZN(n18360) );
  OAI21_X1 U21573 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n18430), .A(
        n18360), .ZN(n18346) );
  AOI22_X1 U21574 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n18346), .B1(
        n18547), .B2(n18323), .ZN(n18341) );
  AOI21_X1 U21575 ( .B1(n18325), .B2(n18324), .A(n18540), .ZN(n18335) );
  INV_X1 U21576 ( .A(n18326), .ZN(n18334) );
  NOR2_X1 U21577 ( .A1(n18674), .A2(n9716), .ZN(n18432) );
  INV_X1 U21578 ( .A(n18327), .ZN(n18695) );
  OAI22_X1 U21579 ( .A1(n18695), .A2(n18689), .B1(n18694), .B2(n18594), .ZN(
        n18362) );
  NOR2_X1 U21580 ( .A1(n10095), .A2(n18362), .ZN(n18329) );
  NOR3_X1 U21581 ( .A1(n18432), .A2(n18329), .A3(n18328), .ZN(n18332) );
  AND2_X1 U21582 ( .A1(n18349), .A2(n18330), .ZN(n18331) );
  NAND2_X1 U21583 ( .A1(n18948), .A2(P3_REIP_REG_28__SCAN_IN), .ZN(n18339) );
  NOR2_X1 U21584 ( .A1(n18483), .A2(n18336), .ZN(n18348) );
  OAI221_X1 U21585 ( .B1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_27__SCAN_IN), .C1(n18337), .C2(n18347), .A(
        n18348), .ZN(n18338) );
  NAND4_X1 U21586 ( .A1(n18341), .A2(n18340), .A3(n18339), .A4(n18338), .ZN(
        P3_U2802) );
  NOR2_X1 U21587 ( .A1(n18342), .A2(n17158), .ZN(n18343) );
  XNOR2_X1 U21588 ( .A(n18343), .B(n12931), .ZN(n18703) );
  OAI22_X1 U21589 ( .A1(n19013), .A2(n19630), .B1(n18529), .B2(n18344), .ZN(
        n18345) );
  AOI221_X1 U21590 ( .B1(n18348), .B2(n18347), .C1(n18346), .C2(
        P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A(n18345), .ZN(n18351) );
  AOI22_X1 U21591 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n18362), .B1(
        n18349), .B2(n10095), .ZN(n18350) );
  OAI211_X1 U21592 ( .C1(n18703), .C2(n18540), .A(n18351), .B(n18350), .ZN(
        P3_U2803) );
  INV_X1 U21593 ( .A(n18352), .ZN(n18353) );
  AOI21_X1 U21594 ( .B1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n9731), .A(
        n18353), .ZN(n18712) );
  AOI21_X1 U21595 ( .B1(n19423), .B2(n18355), .A(
        P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n18359) );
  INV_X1 U21596 ( .A(n18430), .ZN(n18357) );
  OAI21_X1 U21597 ( .B1(n18547), .B2(n18357), .A(n18356), .ZN(n18358) );
  NAND2_X1 U21598 ( .A1(n18948), .A2(P3_REIP_REG_26__SCAN_IN), .ZN(n18710) );
  OAI211_X1 U21599 ( .C1(n18360), .C2(n18359), .A(n18358), .B(n18710), .ZN(
        n18361) );
  AOI21_X1 U21600 ( .B1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n18362), .A(
        n18361), .ZN(n18364) );
  NOR2_X1 U21601 ( .A1(n18730), .A2(n18721), .ZN(n18706) );
  NAND4_X1 U21602 ( .A1(n18383), .A2(n18706), .A3(n18426), .A4(n12936), .ZN(
        n18363) );
  OAI211_X1 U21603 ( .C1(n18712), .C2(n18540), .A(n18364), .B(n18363), .ZN(
        P3_U2804) );
  XNOR2_X1 U21604 ( .A(n18365), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n18728) );
  OAI21_X1 U21605 ( .B1(n18366), .B2(n19560), .A(n18684), .ZN(n18367) );
  AOI21_X1 U21606 ( .B1(n19423), .B2(n9770), .A(n18367), .ZN(n18398) );
  OAI21_X1 U21607 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n18430), .A(
        n18398), .ZN(n18379) );
  NOR2_X1 U21608 ( .A1(n18483), .A2(n9770), .ZN(n18381) );
  OAI211_X1 U21609 ( .C1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A(n18381), .B(n18368), .ZN(n18369) );
  NAND2_X1 U21610 ( .A1(n18948), .A2(P3_REIP_REG_25__SCAN_IN), .ZN(n18720) );
  OAI211_X1 U21611 ( .C1(n18529), .C2(n18370), .A(n18369), .B(n18720), .ZN(
        n18371) );
  AOI21_X1 U21612 ( .B1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n18379), .A(
        n18371), .ZN(n18377) );
  NAND2_X1 U21613 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n18735), .ZN(
        n18372) );
  AOI22_X1 U21614 ( .A1(n18706), .A2(n18735), .B1(n18721), .B2(n18372), .ZN(
        n18725) );
  AOI21_X1 U21615 ( .B1(n18374), .B2(n12931), .A(n18373), .ZN(n18375) );
  XNOR2_X1 U21616 ( .A(n18375), .B(n18721), .ZN(n18724) );
  AOI22_X1 U21617 ( .A1(n9716), .A2(n18725), .B1(n18596), .B2(n18724), .ZN(
        n18376) );
  OAI211_X1 U21618 ( .C1(n18689), .C2(n18728), .A(n18377), .B(n18376), .ZN(
        P3_U2805) );
  NOR2_X1 U21619 ( .A1(n19013), .A2(n19624), .ZN(n18729) );
  AOI221_X1 U21620 ( .B1(n18381), .B2(n18380), .C1(n18379), .C2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A(n18729), .ZN(n18389) );
  INV_X1 U21621 ( .A(n18732), .ZN(n18382) );
  OAI22_X1 U21622 ( .A1(n18382), .A2(n18689), .B1(n18735), .B2(n18594), .ZN(
        n18400) );
  NAND2_X1 U21623 ( .A1(n18383), .A2(n18426), .ZN(n18386) );
  AOI21_X1 U21624 ( .B1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n18385), .A(
        n18384), .ZN(n18742) );
  OAI22_X1 U21625 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n18386), .B1(
        n18742), .B2(n18540), .ZN(n18387) );
  AOI21_X1 U21626 ( .B1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n18400), .A(
        n18387), .ZN(n18388) );
  OAI211_X1 U21627 ( .C1(n18529), .C2(n10028), .A(n18389), .B(n18388), .ZN(
        P3_U2806) );
  OAI21_X1 U21628 ( .B1(n18465), .B2(n18390), .A(n18405), .ZN(n18391) );
  OAI211_X1 U21629 ( .C1(n18509), .C2(n18758), .A(n18433), .B(n18391), .ZN(
        n18392) );
  XOR2_X1 U21630 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B(n18392), .Z(
        n18748) );
  NOR2_X1 U21631 ( .A1(n18586), .A2(n18393), .ZN(n18401) );
  INV_X1 U21632 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n18736) );
  AOI21_X1 U21633 ( .B1(n18394), .B2(n19423), .A(
        P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n18397) );
  OAI21_X1 U21634 ( .B1(n18547), .B2(n18357), .A(n18395), .ZN(n18396) );
  NAND2_X1 U21635 ( .A1(n18866), .A2(P3_REIP_REG_23__SCAN_IN), .ZN(n18747) );
  OAI211_X1 U21636 ( .C1(n18398), .C2(n18397), .A(n18396), .B(n18747), .ZN(
        n18399) );
  AOI221_X1 U21637 ( .B1(n18401), .B2(n18736), .C1(n18400), .C2(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A(n18399), .ZN(n18402) );
  OAI21_X1 U21638 ( .B1(n18540), .B2(n18748), .A(n18402), .ZN(P3_U2807) );
  NAND2_X1 U21639 ( .A1(n18800), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n18751) );
  NOR2_X1 U21640 ( .A1(n18759), .A2(n18751), .ZN(n18755) );
  INV_X1 U21641 ( .A(n18755), .ZN(n18404) );
  INV_X1 U21642 ( .A(n18433), .ZN(n18403) );
  AOI221_X1 U21643 ( .B1(n18833), .B2(n18405), .C1(n18404), .C2(n18405), .A(
        n18403), .ZN(n18406) );
  XNOR2_X1 U21644 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B(n18406), .ZN(
        n18765) );
  NOR2_X1 U21645 ( .A1(n18846), .A2(n18689), .ZN(n18502) );
  AOI21_X1 U21646 ( .B1(n9716), .B2(n18833), .A(n18502), .ZN(n18490) );
  OAI21_X1 U21647 ( .B1(n18432), .B2(n18755), .A(n18490), .ZN(n18427) );
  NAND2_X1 U21648 ( .A1(n18445), .A2(n18407), .ZN(n18408) );
  OAI211_X1 U21649 ( .C1(n9806), .C2(n19023), .A(n18684), .B(n18408), .ZN(
        n18436) );
  AOI21_X1 U21650 ( .B1(n18357), .B2(n18409), .A(n18436), .ZN(n18421) );
  NAND2_X1 U21651 ( .A1(n9806), .A2(n18523), .ZN(n18423) );
  AOI21_X1 U21652 ( .B1(n18422), .B2(n18414), .A(n18423), .ZN(n18411) );
  AOI22_X1 U21653 ( .A1(n18412), .A2(n18547), .B1(n18411), .B2(n18410), .ZN(
        n18413) );
  NAND2_X1 U21654 ( .A1(n18948), .A2(P3_REIP_REG_22__SCAN_IN), .ZN(n18763) );
  OAI211_X1 U21655 ( .C1(n18421), .C2(n18414), .A(n18413), .B(n18763), .ZN(
        n18415) );
  AOI21_X1 U21656 ( .B1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n18427), .A(
        n18415), .ZN(n18417) );
  NAND3_X1 U21657 ( .A1(n18426), .A2(n18755), .A3(n18758), .ZN(n18416) );
  OAI211_X1 U21658 ( .C1(n18540), .C2(n18765), .A(n18417), .B(n18416), .ZN(
        P3_U2808) );
  NOR3_X1 U21659 ( .A1(n18767), .A2(n12931), .A3(n18418), .ZN(n18442) );
  AOI22_X1 U21660 ( .A1(n18771), .A2(n18442), .B1(n18465), .B2(n18419), .ZN(
        n18420) );
  XNOR2_X1 U21661 ( .A(n18420), .B(n18768), .ZN(n18777) );
  NAND2_X1 U21662 ( .A1(n18866), .A2(P3_REIP_REG_21__SCAN_IN), .ZN(n18775) );
  OAI221_X1 U21663 ( .B1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n18423), .C1(
        n18422), .C2(n18421), .A(n18775), .ZN(n18424) );
  AOI21_X1 U21664 ( .B1(n18547), .B2(n18425), .A(n18424), .ZN(n18429) );
  AND2_X1 U21665 ( .A1(n18768), .A2(n18771), .ZN(n18774) );
  NOR2_X1 U21666 ( .A1(n18491), .A2(n18751), .ZN(n18454) );
  AOI22_X1 U21667 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n18427), .B1(
        n18774), .B2(n18454), .ZN(n18428) );
  OAI211_X1 U21668 ( .C1(n18777), .C2(n18540), .A(n18429), .B(n18428), .ZN(
        P3_U2809) );
  NAND2_X1 U21669 ( .A1(n18529), .A2(n18430), .ZN(n18646) );
  AOI22_X1 U21670 ( .A1(n18866), .A2(P3_REIP_REG_20__SCAN_IN), .B1(n18431), 
        .B2(n18646), .ZN(n18441) );
  NOR2_X1 U21671 ( .A1(n18787), .A2(n18751), .ZN(n18750) );
  OAI21_X1 U21672 ( .B1(n18432), .B2(n18750), .A(n18490), .ZN(n18453) );
  OAI221_X1 U21673 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n18463), 
        .C1(n18787), .C2(n18442), .A(n18433), .ZN(n18434) );
  XNOR2_X1 U21674 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .B(n18434), .ZN(
        n18779) );
  AOI22_X1 U21675 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n18453), .B1(
        n18596), .B2(n18779), .ZN(n18440) );
  NAND3_X1 U21676 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18454), .A3(
        n18435), .ZN(n18439) );
  OAI221_X1 U21677 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n19423), .C1(
        P3_PHYADDRPOINTER_REG_20__SCAN_IN), .C2(n18437), .A(n18436), .ZN(
        n18438) );
  NAND4_X1 U21678 ( .A1(n18441), .A2(n18440), .A3(n18439), .A4(n18438), .ZN(
        P3_U2810) );
  AOI21_X1 U21679 ( .B1(n18465), .B2(n18463), .A(n18442), .ZN(n18443) );
  XNOR2_X1 U21680 ( .A(n18443), .B(n18787), .ZN(n18792) );
  INV_X1 U21681 ( .A(n18446), .ZN(n18457) );
  OAI21_X1 U21682 ( .B1(n18457), .B2(n19023), .A(n18684), .ZN(n18471) );
  AOI21_X1 U21683 ( .B1(n18445), .B2(n18444), .A(n18471), .ZN(n18458) );
  AOI211_X1 U21684 ( .C1(n18459), .C2(n18451), .A(n18483), .B(n18446), .ZN(
        n18448) );
  AOI22_X1 U21685 ( .A1(n18449), .A2(n18547), .B1(n18448), .B2(n18447), .ZN(
        n18450) );
  NAND2_X1 U21686 ( .A1(n18866), .A2(P3_REIP_REG_19__SCAN_IN), .ZN(n18790) );
  OAI211_X1 U21687 ( .C1(n18458), .C2(n18451), .A(n18450), .B(n18790), .ZN(
        n18452) );
  AOI221_X1 U21688 ( .B1(n18454), .B2(n18787), .C1(n18453), .C2(
        P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A(n18452), .ZN(n18455) );
  OAI21_X1 U21689 ( .B1(n18792), .B2(n18540), .A(n18455), .ZN(P3_U2811) );
  NAND2_X1 U21690 ( .A1(n18456), .A2(n18767), .ZN(n18807) );
  NAND2_X1 U21691 ( .A1(n18457), .A2(n18523), .ZN(n18460) );
  NAND2_X1 U21692 ( .A1(n18948), .A2(P3_REIP_REG_18__SCAN_IN), .ZN(n18805) );
  OAI221_X1 U21693 ( .B1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n18460), .C1(
        n18459), .C2(n18458), .A(n18805), .ZN(n18461) );
  AOI21_X1 U21694 ( .B1(n18547), .B2(n18462), .A(n18461), .ZN(n18467) );
  OAI21_X1 U21695 ( .B1(n18800), .B2(n18491), .A(n18490), .ZN(n18476) );
  AOI21_X1 U21696 ( .B1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n18509), .A(
        n18463), .ZN(n18464) );
  XOR2_X1 U21697 ( .A(n18465), .B(n18464), .Z(n18803) );
  AOI22_X1 U21698 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n18476), .B1(
        n18596), .B2(n18803), .ZN(n18466) );
  OAI211_X1 U21699 ( .C1(n18586), .C2(n18807), .A(n18467), .B(n18466), .ZN(
        P3_U2812) );
  AOI21_X1 U21700 ( .B1(n18468), .B2(n19423), .A(
        P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n18469) );
  INV_X1 U21701 ( .A(n18469), .ZN(n18470) );
  AOI22_X1 U21702 ( .A1(n18472), .A2(n18646), .B1(n18471), .B2(n18470), .ZN(
        n18478) );
  AOI21_X1 U21703 ( .B1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n18474), .A(
        n18473), .ZN(n18815) );
  NAND2_X1 U21704 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n18808), .ZN(
        n18810) );
  OAI22_X1 U21705 ( .A1(n18815), .A2(n18540), .B1(n18491), .B2(n18810), .ZN(
        n18475) );
  AOI21_X1 U21706 ( .B1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n18476), .A(
        n18475), .ZN(n18477) );
  OAI211_X1 U21707 ( .C1(n19013), .C2(n19611), .A(n18478), .B(n18477), .ZN(
        P3_U2813) );
  OAI21_X1 U21708 ( .B1(n12931), .B2(n18757), .A(n18479), .ZN(n18480) );
  XNOR2_X1 U21709 ( .A(n18480), .B(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n18826) );
  INV_X1 U21710 ( .A(n18684), .ZN(n18637) );
  OAI21_X1 U21711 ( .B1(n18637), .B2(n18482), .A(n18677), .ZN(n18517) );
  OAI21_X1 U21712 ( .B1(n18481), .B2(n19560), .A(n18517), .ZN(n18495) );
  AOI22_X1 U21713 ( .A1(n18866), .A2(P3_REIP_REG_16__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n18495), .ZN(n18486) );
  NOR2_X1 U21714 ( .A1(n18483), .A2(n18482), .ZN(n18497) );
  OAI211_X1 U21715 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(n18497), .B(n18484), .ZN(n18485) );
  OAI211_X1 U21716 ( .C1(n18529), .C2(n18487), .A(n18486), .B(n18485), .ZN(
        n18488) );
  AOI21_X1 U21717 ( .B1(n18596), .B2(n18826), .A(n18488), .ZN(n18489) );
  OAI221_X1 U21718 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n18491), 
        .C1(n18829), .C2(n18490), .A(n18489), .ZN(P3_U2814) );
  AOI21_X1 U21719 ( .B1(n18492), .B2(n17112), .A(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n18840) );
  NAND2_X1 U21720 ( .A1(n9716), .A2(n18833), .ZN(n18505) );
  OAI22_X1 U21721 ( .A1(n19013), .A2(n19606), .B1(n18529), .B2(n18493), .ZN(
        n18494) );
  AOI221_X1 U21722 ( .B1(n18497), .B2(n18496), .C1(n18495), .C2(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A(n18494), .ZN(n18504) );
  INV_X1 U21723 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n18847) );
  NOR3_X1 U21724 ( .A1(n18879), .A2(n18847), .A3(n18855), .ZN(n18499) );
  AOI21_X1 U21725 ( .B1(n17112), .B2(n18499), .A(n18498), .ZN(n18500) );
  AOI221_X1 U21726 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n18880), 
        .C1(n12931), .C2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A(n18500), .ZN(
        n18501) );
  XNOR2_X1 U21727 ( .A(n18501), .B(n18819), .ZN(n18841) );
  NAND2_X1 U21728 ( .A1(n18513), .A2(n18819), .ZN(n18831) );
  AOI22_X1 U21729 ( .A1(n18596), .A2(n18841), .B1(n18502), .B2(n18831), .ZN(
        n18503) );
  OAI211_X1 U21730 ( .C1(n18840), .C2(n18505), .A(n18504), .B(n18503), .ZN(
        P3_U2815) );
  NOR3_X1 U21731 ( .A1(n19354), .A2(n18554), .A3(n18506), .ZN(n18557) );
  AOI21_X1 U21732 ( .B1(n18524), .B2(n18557), .A(
        P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n18518) );
  AOI22_X1 U21733 ( .A1(n18866), .A2(P3_REIP_REG_14__SCAN_IN), .B1(n18507), 
        .B2(n18646), .ZN(n18516) );
  NAND2_X1 U21734 ( .A1(n18872), .A2(n17112), .ZN(n18534) );
  INV_X1 U21735 ( .A(n17112), .ZN(n18591) );
  NOR2_X1 U21736 ( .A1(n18821), .A2(n18591), .ZN(n18508) );
  AOI221_X1 U21737 ( .B1(n18847), .B2(n18855), .C1(n18534), .C2(n18855), .A(
        n18508), .ZN(n18861) );
  NAND2_X1 U21738 ( .A1(n18509), .A2(n17112), .ZN(n18567) );
  NAND2_X1 U21739 ( .A1(n18872), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n18848) );
  OAI21_X1 U21740 ( .B1(n18567), .B2(n18848), .A(n18510), .ZN(n18511) );
  XNOR2_X1 U21741 ( .A(n18511), .B(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n18859) );
  INV_X1 U21742 ( .A(n18512), .ZN(n18890) );
  INV_X1 U21743 ( .A(n18872), .ZN(n18536) );
  NOR2_X1 U21744 ( .A1(n18890), .A2(n18536), .ZN(n18533) );
  OAI221_X1 U21745 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .C1(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n18533), .A(n18513), .ZN(
        n18858) );
  OAI22_X1 U21746 ( .A1(n18859), .A2(n18540), .B1(n18689), .B2(n18858), .ZN(
        n18514) );
  AOI21_X1 U21747 ( .B1(n9716), .B2(n18861), .A(n18514), .ZN(n18515) );
  OAI211_X1 U21748 ( .C1(n18518), .C2(n18517), .A(n18516), .B(n18515), .ZN(
        P3_U2816) );
  NAND2_X1 U21749 ( .A1(n18880), .A2(n12931), .ZN(n18521) );
  OR2_X1 U21750 ( .A1(n18519), .A2(n18520), .ZN(n18548) );
  AOI22_X1 U21751 ( .A1(n18521), .A2(n18534), .B1(n18548), .B2(n12931), .ZN(
        n18522) );
  XNOR2_X1 U21752 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B(n18522), .ZN(
        n18878) );
  NAND2_X1 U21753 ( .A1(n18526), .A2(n18523), .ZN(n18543) );
  AOI211_X1 U21754 ( .C1(n18542), .C2(n18530), .A(n18524), .B(n18543), .ZN(
        n18532) );
  OAI22_X1 U21755 ( .A1(n18526), .A2(n19023), .B1(n18525), .B2(n19560), .ZN(
        n18527) );
  NOR2_X1 U21756 ( .A1(n18637), .A2(n18527), .ZN(n18541) );
  OAI22_X1 U21757 ( .A1(n18541), .A2(n18530), .B1(n18529), .B2(n18528), .ZN(
        n18531) );
  AOI211_X1 U21758 ( .C1(P3_REIP_REG_13__SCAN_IN), .C2(n18948), .A(n18532), 
        .B(n18531), .ZN(n18539) );
  INV_X1 U21759 ( .A(n18533), .ZN(n18869) );
  AOI22_X1 U21760 ( .A1(n18869), .A2(n18674), .B1(n18534), .B2(n9716), .ZN(
        n18535) );
  INV_X1 U21761 ( .A(n18535), .ZN(n18550) );
  NOR2_X1 U21762 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n18536), .ZN(
        n18865) );
  INV_X1 U21763 ( .A(n18586), .ZN(n18537) );
  AOI22_X1 U21764 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n18550), .B1(
        n18865), .B2(n18537), .ZN(n18538) );
  OAI211_X1 U21765 ( .C1(n18540), .C2(n18878), .A(n18539), .B(n18538), .ZN(
        P3_U2817) );
  NOR3_X1 U21766 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n18586), .A3(
        n18879), .ZN(n18545) );
  NAND2_X1 U21767 ( .A1(n18866), .A2(P3_REIP_REG_12__SCAN_IN), .ZN(n18885) );
  OAI221_X1 U21768 ( .B1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n18543), .C1(
        n18542), .C2(n18541), .A(n18885), .ZN(n18544) );
  AOI211_X1 U21769 ( .C1(n18547), .C2(n18546), .A(n18545), .B(n18544), .ZN(
        n18552) );
  OAI21_X1 U21770 ( .B1(n18879), .B2(n18567), .A(n18548), .ZN(n18549) );
  XNOR2_X1 U21771 ( .A(n18549), .B(n18880), .ZN(n18884) );
  AOI22_X1 U21772 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n18550), .B1(
        n18596), .B2(n18884), .ZN(n18551) );
  NAND2_X1 U21773 ( .A1(n18552), .A2(n18551), .ZN(P3_U2818) );
  INV_X1 U21774 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n18553) );
  NAND2_X1 U21775 ( .A1(n18895), .A2(n18553), .ZN(n18900) );
  NOR2_X1 U21776 ( .A1(n19354), .A2(n18554), .ZN(n18588) );
  NAND3_X1 U21777 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A3(n18588), .ZN(n18565) );
  NOR2_X1 U21778 ( .A1(n18555), .A2(n18565), .ZN(n18574) );
  AOI21_X1 U21779 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n18677), .A(
        n18574), .ZN(n18556) );
  OAI22_X1 U21780 ( .A1(n18557), .A2(n18556), .B1(n19013), .B2(n19598), .ZN(
        n18558) );
  AOI21_X1 U21781 ( .B1(n18559), .B2(n18646), .A(n18558), .ZN(n18564) );
  AOI22_X1 U21782 ( .A1(n18674), .A2(n18890), .B1(n9716), .B2(n18591), .ZN(
        n18585) );
  OAI21_X1 U21783 ( .B1(n18895), .B2(n18586), .A(n18585), .ZN(n18570) );
  INV_X1 U21784 ( .A(n18567), .ZN(n18577) );
  NOR2_X1 U21785 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n18519), .ZN(
        n18561) );
  AOI21_X1 U21786 ( .B1(n18895), .B2(n18577), .A(n18561), .ZN(n18562) );
  XNOR2_X1 U21787 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n18562), .ZN(
        n18888) );
  AOI22_X1 U21788 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n18570), .B1(
        n18596), .B2(n18888), .ZN(n18563) );
  OAI211_X1 U21789 ( .C1(n18586), .C2(n18900), .A(n18564), .B(n18563), .ZN(
        P3_U2819) );
  INV_X1 U21790 ( .A(n18565), .ZN(n18581) );
  AOI21_X1 U21791 ( .B1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n18677), .A(
        n18581), .ZN(n18573) );
  AOI22_X1 U21792 ( .A1(n18866), .A2(P3_REIP_REG_10__SCAN_IN), .B1(n18566), 
        .B2(n18646), .ZN(n18572) );
  OAI21_X1 U21793 ( .B1(n18919), .B2(n18567), .A(n18519), .ZN(n18568) );
  XNOR2_X1 U21794 ( .A(n18568), .B(n18906), .ZN(n18901) );
  OAI21_X1 U21795 ( .B1(n18586), .B2(n18919), .A(n18906), .ZN(n18569) );
  AOI22_X1 U21796 ( .A1(n18596), .A2(n18901), .B1(n18570), .B2(n18569), .ZN(
        n18571) );
  OAI211_X1 U21797 ( .C1(n18574), .C2(n18573), .A(n18572), .B(n18571), .ZN(
        P3_U2820) );
  AND2_X1 U21798 ( .A1(n12931), .A2(n18575), .ZN(n18576) );
  NOR2_X1 U21799 ( .A1(n18577), .A2(n18576), .ZN(n18578) );
  XNOR2_X1 U21800 ( .A(n18578), .B(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n18916) );
  NOR2_X1 U21801 ( .A1(n19013), .A2(n19594), .ZN(n18583) );
  AOI22_X1 U21802 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n18677), .B1(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n18588), .ZN(n18580) );
  OAI22_X1 U21803 ( .A1(n18581), .A2(n18580), .B1(n18681), .B2(n18579), .ZN(
        n18582) );
  AOI211_X1 U21804 ( .C1(n18596), .C2(n18916), .A(n18583), .B(n18582), .ZN(
        n18584) );
  OAI221_X1 U21805 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18586), .C1(
        n18919), .C2(n18585), .A(n18584), .ZN(P3_U2821) );
  AOI22_X1 U21806 ( .A1(n18589), .A2(n18646), .B1(n18588), .B2(n18587), .ZN(
        n18599) );
  NAND2_X1 U21807 ( .A1(n18591), .A2(n18590), .ZN(n18921) );
  XNOR2_X1 U21808 ( .A(n12931), .B(n18921), .ZN(n18925) );
  OAI21_X1 U21809 ( .B1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n18593), .A(
        n18592), .ZN(n18923) );
  OAI22_X1 U21810 ( .A1(n18689), .A2(n18923), .B1(n18594), .B2(n18921), .ZN(
        n18595) );
  AOI21_X1 U21811 ( .B1(n18596), .B2(n18925), .A(n18595), .ZN(n18598) );
  NAND2_X1 U21812 ( .A1(n18948), .A2(P3_REIP_REG_8__SCAN_IN), .ZN(n18936) );
  NOR2_X1 U21813 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n19354), .ZN(
        n18600) );
  OAI21_X1 U21814 ( .B1(n17507), .B2(n19023), .A(n18684), .ZN(n18601) );
  OAI21_X1 U21815 ( .B1(n18600), .B2(n18601), .A(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n18597) );
  NAND4_X1 U21816 ( .A1(n18599), .A2(n18598), .A3(n18936), .A4(n18597), .ZN(
        P3_U2822) );
  AOI22_X1 U21817 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n18601), .B1(
        n17507), .B2(n18600), .ZN(n18611) );
  AOI21_X1 U21818 ( .B1(n18946), .B2(n18603), .A(n18602), .ZN(n18943) );
  OAI21_X1 U21819 ( .B1(n18606), .B2(n18605), .A(n18604), .ZN(n18607) );
  XNOR2_X1 U21820 ( .A(n18607), .B(n18946), .ZN(n18940) );
  OAI22_X1 U21821 ( .A1(n18681), .A2(n18608), .B1(n18689), .B2(n18940), .ZN(
        n18609) );
  AOI21_X1 U21822 ( .B1(n18678), .B2(n18943), .A(n18609), .ZN(n18610) );
  OAI211_X1 U21823 ( .C1(n19013), .C2(n19590), .A(n18611), .B(n18610), .ZN(
        P3_U2823) );
  AOI21_X1 U21824 ( .B1(n18614), .B2(n18613), .A(n18612), .ZN(n18952) );
  NOR2_X1 U21825 ( .A1(n19354), .A2(n18618), .ZN(n18615) );
  AOI22_X1 U21826 ( .A1(n18678), .A2(n18952), .B1(n18615), .B2(n18619), .ZN(
        n18623) );
  OAI21_X1 U21827 ( .B1(n18617), .B2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n18616), .ZN(n18955) );
  OAI21_X1 U21828 ( .B1(n18618), .B2(n19354), .A(n18677), .ZN(n18631) );
  OAI22_X1 U21829 ( .A1(n18689), .A2(n18955), .B1(n18619), .B2(n18631), .ZN(
        n18620) );
  AOI21_X1 U21830 ( .B1(n18621), .B2(n18646), .A(n18620), .ZN(n18622) );
  OAI211_X1 U21831 ( .C1(n19013), .C2(n19588), .A(n18623), .B(n18622), .ZN(
        P3_U2824) );
  OAI21_X1 U21832 ( .B1(n18626), .B2(n18625), .A(n18624), .ZN(n18962) );
  AOI21_X1 U21833 ( .B1(n18629), .B2(n18628), .A(n18627), .ZN(n18959) );
  AOI21_X1 U21834 ( .B1(n18630), .B2(n18684), .A(
        P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n18632) );
  OAI22_X1 U21835 ( .A1(n18681), .A2(n18633), .B1(n18632), .B2(n18631), .ZN(
        n18634) );
  AOI21_X1 U21836 ( .B1(n18678), .B2(n18959), .A(n18634), .ZN(n18635) );
  NAND2_X1 U21837 ( .A1(n18948), .A2(P3_REIP_REG_5__SCAN_IN), .ZN(n18960) );
  OAI211_X1 U21838 ( .C1(n18689), .C2(n18962), .A(n18635), .B(n18960), .ZN(
        P3_U2825) );
  OAI21_X1 U21839 ( .B1(n18637), .B2(n18636), .A(n18677), .ZN(n18661) );
  OAI21_X1 U21840 ( .B1(n18640), .B2(n18639), .A(n18638), .ZN(n18974) );
  OAI22_X1 U21841 ( .A1(n18689), .A2(n18974), .B1(n19354), .B2(n18641), .ZN(
        n18642) );
  AOI21_X1 U21842 ( .B1(n18948), .B2(P3_REIP_REG_4__SCAN_IN), .A(n18642), .ZN(
        n18649) );
  AOI21_X1 U21843 ( .B1(n18645), .B2(n18644), .A(n18643), .ZN(n18972) );
  AOI22_X1 U21844 ( .A1(n18678), .A2(n18972), .B1(n18647), .B2(n18646), .ZN(
        n18648) );
  OAI211_X1 U21845 ( .C1(n18650), .C2(n18661), .A(n18649), .B(n18648), .ZN(
        P3_U2826) );
  NAND2_X1 U21846 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n18684), .ZN(
        n18659) );
  AOI21_X1 U21847 ( .B1(n18976), .B2(n18652), .A(n18651), .ZN(n18979) );
  NOR2_X1 U21848 ( .A1(n19013), .A2(n19582), .ZN(n18978) );
  OAI21_X1 U21849 ( .B1(n18655), .B2(n18654), .A(n18653), .ZN(n18975) );
  OAI22_X1 U21850 ( .A1(n18681), .A2(n18656), .B1(n18689), .B2(n18975), .ZN(
        n18657) );
  AOI211_X1 U21851 ( .C1(n18678), .C2(n18979), .A(n18978), .B(n18657), .ZN(
        n18658) );
  OAI221_X1 U21852 ( .B1(n18661), .B2(n18660), .C1(n18661), .C2(n18659), .A(
        n18658), .ZN(P3_U2827) );
  AOI21_X1 U21853 ( .B1(n18664), .B2(n18663), .A(n18662), .ZN(n18993) );
  NOR2_X1 U21854 ( .A1(n19580), .A2(n19013), .ZN(n18996) );
  OAI21_X1 U21855 ( .B1(n18667), .B2(n18666), .A(n18665), .ZN(n18992) );
  OAI22_X1 U21856 ( .A1(n18681), .A2(n18668), .B1(n18689), .B2(n18992), .ZN(
        n18669) );
  AOI211_X1 U21857 ( .C1(n18678), .C2(n18993), .A(n18996), .B(n18669), .ZN(
        n18670) );
  OAI221_X1 U21858 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n19354), .C1(
        n18671), .C2(n18684), .A(n18670), .ZN(P3_U2828) );
  NOR2_X1 U21859 ( .A1(n18683), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n18672) );
  XOR2_X1 U21860 ( .A(n18676), .B(n18672), .Z(n19009) );
  INV_X1 U21861 ( .A(n19009), .ZN(n18673) );
  AOI22_X1 U21862 ( .A1(n18674), .A2(n18673), .B1(n18948), .B2(
        P3_REIP_REG_1__SCAN_IN), .ZN(n18680) );
  AOI21_X1 U21863 ( .B1(n18676), .B2(n18682), .A(n18675), .ZN(n19004) );
  AOI22_X1 U21864 ( .A1(n18678), .A2(n19004), .B1(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n18677), .ZN(n18679) );
  OAI211_X1 U21865 ( .C1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n18681), .A(
        n18680), .B(n18679), .ZN(P3_U2829) );
  OAI21_X1 U21866 ( .B1(n18683), .B2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n18682), .ZN(n18688) );
  INV_X1 U21867 ( .A(n18688), .ZN(n19018) );
  NAND3_X1 U21868 ( .A1(n19660), .A2(n19560), .A3(n18684), .ZN(n18685) );
  AOI22_X1 U21869 ( .A1(n18866), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n18685), .ZN(n18686) );
  OAI221_X1 U21870 ( .B1(n19018), .B2(n18689), .C1(n18688), .C2(n18687), .A(
        n18686), .ZN(P3_U2830) );
  AOI22_X1 U21871 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n19006), .B1(
        n18948), .B2(P3_REIP_REG_27__SCAN_IN), .ZN(n18702) );
  INV_X1 U21872 ( .A(n18716), .ZN(n18692) );
  NOR2_X1 U21873 ( .A1(n18914), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n18963) );
  INV_X1 U21874 ( .A(n18690), .ZN(n18691) );
  INV_X1 U21875 ( .A(n18928), .ZN(n18965) );
  OAI21_X1 U21876 ( .B1(n18963), .B2(n18691), .A(n18965), .ZN(n18733) );
  OAI21_X1 U21877 ( .B1(n18928), .B2(n18692), .A(n18733), .ZN(n18715) );
  OAI22_X1 U21878 ( .A1(n19517), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B1(
        n18914), .B2(n18693), .ZN(n18697) );
  OAI22_X1 U21879 ( .A1(n18695), .A2(n19483), .B1(n18694), .B2(n18871), .ZN(
        n18696) );
  OAI211_X1 U21880 ( .C1(n19517), .C2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B(n18708), .ZN(n18699) );
  OAI211_X1 U21881 ( .C1(n18700), .C2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n18995), .B(n18699), .ZN(n18701) );
  OAI211_X1 U21882 ( .C1(n18703), .C2(n18877), .A(n18702), .B(n18701), .ZN(
        P3_U2835) );
  NAND2_X1 U21883 ( .A1(n18995), .A2(n18704), .ZN(n18766) );
  NOR2_X1 U21884 ( .A1(n18705), .A2(n18766), .ZN(n18731) );
  AOI22_X1 U21885 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n18995), .B1(
        n18706), .B2(n18731), .ZN(n18707) );
  AOI21_X1 U21886 ( .B1(n18708), .B2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n18707), .ZN(n18709) );
  AOI21_X1 U21887 ( .B1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n19006), .A(
        n18709), .ZN(n18711) );
  OAI211_X1 U21888 ( .C1(n18712), .C2(n18877), .A(n18711), .B(n18710), .ZN(
        P3_U2836) );
  NOR2_X1 U21889 ( .A1(n18716), .A2(n18713), .ZN(n18719) );
  INV_X1 U21890 ( .A(n19509), .ZN(n19489) );
  INV_X1 U21891 ( .A(n18714), .ZN(n18737) );
  AOI221_X1 U21892 ( .B1(n18716), .B2(n19489), .C1(n18737), .C2(n19489), .A(
        n18715), .ZN(n18717) );
  INV_X1 U21893 ( .A(n18717), .ZN(n18718) );
  MUX2_X1 U21894 ( .A(n18719), .B(n18718), .S(
        P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Z(n18723) );
  INV_X1 U21895 ( .A(n19006), .ZN(n19000) );
  OAI21_X1 U21896 ( .B1(n19000), .B2(n18721), .A(n18720), .ZN(n18722) );
  AOI21_X1 U21897 ( .B1(n18995), .B2(n18723), .A(n18722), .ZN(n18727) );
  AOI22_X1 U21898 ( .A1(n18862), .A2(n18725), .B1(n18926), .B2(n18724), .ZN(
        n18726) );
  OAI211_X1 U21899 ( .C1(n19017), .C2(n18728), .A(n18727), .B(n18726), .ZN(
        P3_U2837) );
  AOI21_X1 U21900 ( .B1(n18731), .B2(n18730), .A(n18729), .ZN(n18741) );
  AOI21_X1 U21901 ( .B1(n18891), .B2(n18732), .A(n19006), .ZN(n18734) );
  OAI211_X1 U21902 ( .C1(n18735), .C2(n18871), .A(n18734), .B(n18733), .ZN(
        n18739) );
  AOI211_X1 U21903 ( .C1(n19489), .C2(n18737), .A(n18736), .B(n18739), .ZN(
        n18738) );
  NOR2_X1 U21904 ( .A1(n18948), .A2(n18738), .ZN(n18744) );
  OAI211_X1 U21905 ( .C1(n18824), .C2(n18739), .A(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B(n18744), .ZN(n18740) );
  OAI211_X1 U21906 ( .C1(n18742), .C2(n18877), .A(n18741), .B(n18740), .ZN(
        P3_U2838) );
  NOR2_X1 U21907 ( .A1(n19006), .A2(n18743), .ZN(n18745) );
  OAI21_X1 U21908 ( .B1(n18745), .B2(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n18744), .ZN(n18746) );
  OAI211_X1 U21909 ( .C1(n18748), .C2(n18877), .A(n18747), .B(n18746), .ZN(
        P3_U2839) );
  OAI22_X1 U21910 ( .A1(n18758), .A2(n19014), .B1(n18749), .B2(n18766), .ZN(
        n18762) );
  INV_X1 U21911 ( .A(n18750), .ZN(n18782) );
  NOR3_X1 U21912 ( .A1(n18811), .A2(n18849), .A3(n18782), .ZN(n18754) );
  OAI21_X1 U21913 ( .B1(n18767), .B2(n18802), .A(n19489), .ZN(n18753) );
  NOR2_X1 U21914 ( .A1(n19677), .A2(n18849), .ZN(n18913) );
  NAND2_X1 U21915 ( .A1(n18816), .A2(n18913), .ZN(n18818) );
  OAI21_X1 U21916 ( .B1(n18751), .B2(n18818), .A(n19515), .ZN(n18752) );
  OAI211_X1 U21917 ( .C1(n19517), .C2(n18754), .A(n18753), .B(n18752), .ZN(
        n18780) );
  NOR2_X1 U21918 ( .A1(n18891), .A2(n18834), .ZN(n18894) );
  OAI22_X1 U21919 ( .A1(n19517), .A2(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .B1(
        n18755), .B2(n18894), .ZN(n18756) );
  NOR2_X1 U21920 ( .A1(n18780), .A2(n18756), .ZN(n18770) );
  OAI22_X1 U21921 ( .A1(n18846), .A2(n19483), .B1(n18757), .B2(n18871), .ZN(
        n18769) );
  AOI211_X1 U21922 ( .C1(n18824), .C2(n18759), .A(n18758), .B(n18769), .ZN(
        n18760) );
  NAND2_X1 U21923 ( .A1(n18770), .A2(n18760), .ZN(n18761) );
  AOI22_X1 U21924 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n19006), .B1(
        n18762), .B2(n18761), .ZN(n18764) );
  OAI211_X1 U21925 ( .C1(n18765), .C2(n18877), .A(n18764), .B(n18763), .ZN(
        P3_U2840) );
  NOR2_X1 U21926 ( .A1(n18767), .A2(n18766), .ZN(n18788) );
  NOR2_X1 U21927 ( .A1(n18948), .A2(n18768), .ZN(n18773) );
  NOR2_X1 U21928 ( .A1(n19489), .A2(n19515), .ZN(n19005) );
  OAI211_X1 U21929 ( .C1(n18771), .C2(n19005), .A(n18817), .B(n18770), .ZN(
        n18772) );
  AOI22_X1 U21930 ( .A1(n18774), .A2(n18788), .B1(n18773), .B2(n18772), .ZN(
        n18776) );
  OAI211_X1 U21931 ( .C1(n18777), .C2(n18877), .A(n18776), .B(n18775), .ZN(
        P3_U2841) );
  NOR2_X1 U21932 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n18787), .ZN(
        n18778) );
  AOI22_X1 U21933 ( .A1(n18926), .A2(n18779), .B1(n18788), .B2(n18778), .ZN(
        n18786) );
  INV_X1 U21934 ( .A(n18894), .ZN(n18781) );
  AOI21_X1 U21935 ( .B1(n18782), .B2(n18781), .A(n18780), .ZN(n18783) );
  AOI21_X1 U21936 ( .B1(n18817), .B2(n18783), .A(n18948), .ZN(n18789) );
  NOR3_X1 U21937 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n19005), .A3(
        n19712), .ZN(n18784) );
  OAI21_X1 U21938 ( .B1(n18789), .B2(n18784), .A(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n18785) );
  OAI211_X1 U21939 ( .C1(n19617), .C2(n19013), .A(n18786), .B(n18785), .ZN(
        P3_U2842) );
  AOI22_X1 U21940 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18789), .B1(
        n18788), .B2(n18787), .ZN(n18791) );
  OAI211_X1 U21941 ( .C1(n18792), .C2(n18877), .A(n18791), .B(n18790), .ZN(
        P3_U2843) );
  AOI22_X1 U21942 ( .A1(n19489), .A2(n18986), .B1(n18793), .B2(n18989), .ZN(
        n18794) );
  INV_X1 U21943 ( .A(n18794), .ZN(n18981) );
  NAND2_X1 U21944 ( .A1(n18981), .A2(n18795), .ZN(n18949) );
  INV_X1 U21945 ( .A(n18949), .ZN(n18939) );
  NAND2_X1 U21946 ( .A1(n18796), .A2(n18939), .ZN(n18835) );
  NAND2_X1 U21947 ( .A1(n18797), .A2(n18835), .ZN(n18882) );
  NAND2_X1 U21948 ( .A1(n18995), .A2(n18882), .ZN(n18920) );
  NAND2_X1 U21949 ( .A1(n18816), .A2(n18820), .ZN(n18798) );
  OAI21_X1 U21950 ( .B1(n18829), .B2(n18798), .A(n18965), .ZN(n18799) );
  OAI211_X1 U21951 ( .C1(n18800), .C2(n18894), .A(n18817), .B(n18799), .ZN(
        n18801) );
  AOI211_X1 U21952 ( .C1(n19489), .C2(n18802), .A(n18963), .B(n18801), .ZN(
        n18809) );
  AOI221_X1 U21953 ( .B1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n9712), .C1(
        n18928), .C2(n9712), .A(n18866), .ZN(n18804) );
  AOI22_X1 U21954 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n18804), .B1(
        n18926), .B2(n18803), .ZN(n18806) );
  OAI211_X1 U21955 ( .C1(n18807), .C2(n18920), .A(n18806), .B(n18805), .ZN(
        P3_U2844) );
  NOR2_X1 U21956 ( .A1(n9712), .A2(n18808), .ZN(n18813) );
  NOR3_X1 U21957 ( .A1(n18811), .A2(n18920), .A3(n18810), .ZN(n18812) );
  AOI221_X1 U21958 ( .B1(P3_REIP_REG_17__SCAN_IN), .B2(n18948), .C1(n18813), 
        .C2(n19013), .A(n18812), .ZN(n18814) );
  OAI21_X1 U21959 ( .B1(n18815), .B2(n18877), .A(n18814), .ZN(P3_U2845) );
  INV_X1 U21960 ( .A(n18920), .ZN(n18907) );
  NAND2_X1 U21961 ( .A1(n18816), .A2(n18907), .ZN(n18830) );
  INV_X1 U21962 ( .A(n18817), .ZN(n18825) );
  OAI21_X1 U21963 ( .B1(n18819), .B2(n19515), .A(n18818), .ZN(n18823) );
  NOR2_X1 U21964 ( .A1(n19517), .A2(n18820), .ZN(n18902) );
  OAI21_X1 U21965 ( .B1(n18902), .B2(n18821), .A(n18873), .ZN(n18822) );
  OAI211_X1 U21966 ( .C1(n18867), .C2(n19509), .A(n18823), .B(n18822), .ZN(
        n18837) );
  OAI221_X1 U21967 ( .B1(n18825), .B2(n18824), .C1(n18825), .C2(n18837), .A(
        n19013), .ZN(n18828) );
  AOI22_X1 U21968 ( .A1(n18948), .A2(P3_REIP_REG_16__SCAN_IN), .B1(n18926), 
        .B2(n18826), .ZN(n18827) );
  OAI221_X1 U21969 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n18830), 
        .C1(n18829), .C2(n18828), .A(n18827), .ZN(P3_U2846) );
  NAND2_X1 U21970 ( .A1(n18832), .A2(n18831), .ZN(n18845) );
  AOI22_X1 U21971 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n19006), .B1(
        n18948), .B2(P3_REIP_REG_15__SCAN_IN), .ZN(n18844) );
  NAND2_X1 U21972 ( .A1(n18834), .A2(n18833), .ZN(n18839) );
  NOR2_X1 U21973 ( .A1(n18835), .A2(n18848), .ZN(n18857) );
  OAI211_X1 U21974 ( .C1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n18857), .A(
        n18837), .B(n18836), .ZN(n18838) );
  OAI21_X1 U21975 ( .B1(n18840), .B2(n18839), .A(n18838), .ZN(n18842) );
  AOI22_X1 U21976 ( .A1(n18995), .A2(n18842), .B1(n18926), .B2(n18841), .ZN(
        n18843) );
  OAI211_X1 U21977 ( .C1(n18846), .C2(n18845), .A(n18844), .B(n18843), .ZN(
        P3_U2847) );
  INV_X1 U21978 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n19604) );
  AOI21_X1 U21979 ( .B1(n18872), .B2(n18867), .A(n19509), .ZN(n18853) );
  AOI21_X1 U21980 ( .B1(n18872), .B2(n18913), .A(n18914), .ZN(n18868) );
  NOR2_X1 U21981 ( .A1(n18868), .A2(n18847), .ZN(n18851) );
  OAI21_X1 U21982 ( .B1(n18849), .B2(n18848), .A(n19499), .ZN(n18850) );
  OAI211_X1 U21983 ( .C1(n19005), .C2(n18851), .A(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B(n18850), .ZN(n18852) );
  OAI21_X1 U21984 ( .B1(n18853), .B2(n18852), .A(n18995), .ZN(n18854) );
  OAI21_X1 U21985 ( .B1(n19000), .B2(n18855), .A(n18854), .ZN(n18856) );
  OAI21_X1 U21986 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n18857), .A(
        n18856), .ZN(n18864) );
  OAI22_X1 U21987 ( .A1(n18859), .A2(n18877), .B1(n19017), .B2(n18858), .ZN(
        n18860) );
  AOI21_X1 U21988 ( .B1(n18862), .B2(n18861), .A(n18860), .ZN(n18863) );
  OAI211_X1 U21989 ( .C1(n19013), .C2(n19604), .A(n18864), .B(n18863), .ZN(
        P3_U2848) );
  AOI22_X1 U21990 ( .A1(n18866), .A2(P3_REIP_REG_13__SCAN_IN), .B1(n18907), 
        .B2(n18865), .ZN(n18876) );
  OAI22_X1 U21991 ( .A1(n17112), .A2(n18871), .B1(n18867), .B2(n19509), .ZN(
        n18889) );
  AOI211_X1 U21992 ( .C1(n18891), .C2(n18869), .A(n18868), .B(n18889), .ZN(
        n18870) );
  OAI21_X1 U21993 ( .B1(n18902), .B2(n18879), .A(n18873), .ZN(n18896) );
  OAI211_X1 U21994 ( .C1(n18872), .C2(n18871), .A(n18870), .B(n18896), .ZN(
        n18881) );
  INV_X1 U21995 ( .A(n18873), .ZN(n18903) );
  OAI21_X1 U21996 ( .B1(n18903), .B2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n18995), .ZN(n18874) );
  OAI211_X1 U21997 ( .C1(n18881), .C2(n18874), .A(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B(n19013), .ZN(n18875) );
  OAI211_X1 U21998 ( .C1(n18878), .C2(n18877), .A(n18876), .B(n18875), .ZN(
        P3_U2849) );
  INV_X1 U21999 ( .A(n18879), .ZN(n18883) );
  OAI222_X1 U22000 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n18883), 
        .B1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n18882), .C1(n18881), 
        .C2(n18880), .ZN(n18887) );
  AOI22_X1 U22001 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n19006), .B1(
        n18926), .B2(n18884), .ZN(n18886) );
  OAI211_X1 U22002 ( .C1(n19014), .C2(n18887), .A(n18886), .B(n18885), .ZN(
        P3_U2850) );
  AOI22_X1 U22003 ( .A1(n18948), .A2(P3_REIP_REG_11__SCAN_IN), .B1(n18926), 
        .B2(n18888), .ZN(n18899) );
  AOI21_X1 U22004 ( .B1(n18891), .B2(n18890), .A(n18889), .ZN(n18912) );
  AOI21_X1 U22005 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18913), .A(
        n18914), .ZN(n18892) );
  INV_X1 U22006 ( .A(n18892), .ZN(n18893) );
  OAI211_X1 U22007 ( .C1(n18895), .C2(n18894), .A(n18912), .B(n18893), .ZN(
        n18905) );
  OAI211_X1 U22008 ( .C1(n18914), .C2(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n18995), .B(n18896), .ZN(n18897) );
  OAI211_X1 U22009 ( .C1(n18905), .C2(n18897), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n19013), .ZN(n18898) );
  OAI211_X1 U22010 ( .C1(n18900), .C2(n18920), .A(n18899), .B(n18898), .ZN(
        P3_U2851) );
  AOI22_X1 U22011 ( .A1(n18948), .A2(P3_REIP_REG_10__SCAN_IN), .B1(n18926), 
        .B2(n18901), .ZN(n18910) );
  NOR2_X1 U22012 ( .A1(n18902), .A2(n19014), .ZN(n18911) );
  OAI21_X1 U22013 ( .B1(n18903), .B2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n18911), .ZN(n18904) );
  OAI211_X1 U22014 ( .C1(n18905), .C2(n18904), .A(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B(n19013), .ZN(n18909) );
  NAND3_X1 U22015 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n18907), .A3(
        n18906), .ZN(n18908) );
  NAND3_X1 U22016 ( .A1(n18910), .A2(n18909), .A3(n18908), .ZN(P3_U2852) );
  OAI211_X1 U22017 ( .C1(n18914), .C2(n18913), .A(n18912), .B(n18911), .ZN(
        n18915) );
  NAND2_X1 U22018 ( .A1(n19013), .A2(n18915), .ZN(n18918) );
  AOI22_X1 U22019 ( .A1(n18948), .A2(P3_REIP_REG_9__SCAN_IN), .B1(n18926), 
        .B2(n18916), .ZN(n18917) );
  OAI221_X1 U22020 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18920), .C1(
        n18919), .C2(n18918), .A(n18917), .ZN(P3_U2853) );
  OAI22_X1 U22021 ( .A1(n19017), .A2(n18923), .B1(n18922), .B2(n18921), .ZN(
        n18924) );
  AOI21_X1 U22022 ( .B1(n18926), .B2(n18925), .A(n18924), .ZN(n18937) );
  INV_X1 U22023 ( .A(n19001), .ZN(n18966) );
  NOR2_X1 U22024 ( .A1(n18928), .A2(n18927), .ZN(n18929) );
  AOI211_X1 U22025 ( .C1(n19489), .C2(n18930), .A(n18963), .B(n18929), .ZN(
        n18947) );
  OAI21_X1 U22026 ( .B1(n18931), .B2(n18933), .A(n18947), .ZN(n18938) );
  OAI221_X1 U22027 ( .B1(n19006), .B2(n18966), .C1(n19006), .C2(n18938), .A(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n18935) );
  NAND4_X1 U22028 ( .A1(n18995), .A2(n18933), .A3(n18939), .A4(n18932), .ZN(
        n18934) );
  NAND4_X1 U22029 ( .A1(n18937), .A2(n18936), .A3(n18935), .A4(n18934), .ZN(
        P3_U2854) );
  OAI221_X1 U22030 ( .B1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .C1(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .C2(n18939), .A(n18938), .ZN(
        n18941) );
  OAI22_X1 U22031 ( .A1(n19014), .A2(n18941), .B1(n19017), .B2(n18940), .ZN(
        n18942) );
  AOI21_X1 U22032 ( .B1(n19012), .B2(n18943), .A(n18942), .ZN(n18945) );
  NAND2_X1 U22033 ( .A1(n18948), .A2(P3_REIP_REG_7__SCAN_IN), .ZN(n18944) );
  OAI211_X1 U22034 ( .C1(n19000), .C2(n18946), .A(n18945), .B(n18944), .ZN(
        P3_U2855) );
  OAI21_X1 U22035 ( .B1(n18947), .B2(n19014), .A(n19000), .ZN(n18956) );
  AOI22_X1 U22036 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n18956), .B1(
        n18948), .B2(P3_REIP_REG_6__SCAN_IN), .ZN(n18954) );
  NOR2_X1 U22037 ( .A1(n19014), .A2(n18949), .ZN(n18951) );
  AOI22_X1 U22038 ( .A1(n18952), .A2(n19012), .B1(n18951), .B2(n18950), .ZN(
        n18953) );
  OAI211_X1 U22039 ( .C1(n19017), .C2(n18955), .A(n18954), .B(n18953), .ZN(
        P3_U2856) );
  NAND3_X1 U22040 ( .A1(n18995), .A2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        n18981), .ZN(n18968) );
  NOR2_X1 U22041 ( .A1(n18967), .A2(n18968), .ZN(n18957) );
  MUX2_X1 U22042 ( .A(n18957), .B(n18956), .S(
        P3_INSTADDRPOINTER_REG_5__SCAN_IN), .Z(n18958) );
  AOI21_X1 U22043 ( .B1(n19012), .B2(n18959), .A(n18958), .ZN(n18961) );
  OAI211_X1 U22044 ( .C1(n19017), .C2(n18962), .A(n18961), .B(n18960), .ZN(
        P3_U2857) );
  NOR2_X1 U22045 ( .A1(n19013), .A2(n19584), .ZN(n18971) );
  AOI21_X1 U22046 ( .B1(n18965), .B2(n18964), .A(n18963), .ZN(n18984) );
  OAI211_X1 U22047 ( .C1(n19509), .C2(n18986), .A(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B(n18984), .ZN(n18980) );
  AOI21_X1 U22048 ( .B1(n18966), .B2(n18980), .A(n19006), .ZN(n18969) );
  AOI22_X1 U22049 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n18969), .B1(
        n18968), .B2(n18967), .ZN(n18970) );
  AOI211_X1 U22050 ( .C1(n18972), .C2(n19012), .A(n18971), .B(n18970), .ZN(
        n18973) );
  OAI21_X1 U22051 ( .B1(n19017), .B2(n18974), .A(n18973), .ZN(P3_U2858) );
  OAI22_X1 U22052 ( .A1(n18976), .A2(n19000), .B1(n19017), .B2(n18975), .ZN(
        n18977) );
  AOI211_X1 U22053 ( .C1(n19012), .C2(n18979), .A(n18978), .B(n18977), .ZN(
        n18983) );
  OAI211_X1 U22054 ( .C1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .C2(n18981), .A(
        n18995), .B(n18980), .ZN(n18982) );
  NAND2_X1 U22055 ( .A1(n18983), .A2(n18982), .ZN(P3_U2859) );
  NAND2_X1 U22056 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18985) );
  OAI21_X1 U22057 ( .B1(n19509), .B2(n18985), .A(n18984), .ZN(n18988) );
  NOR2_X1 U22058 ( .A1(n19509), .A2(n18986), .ZN(n18987) );
  AOI21_X1 U22059 ( .B1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n18988), .A(
        n18987), .ZN(n18991) );
  NAND3_X1 U22060 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n18989), .A3(
        n18999), .ZN(n18990) );
  OAI211_X1 U22061 ( .C1(n18992), .C2(n19483), .A(n18991), .B(n18990), .ZN(
        n18994) );
  AOI22_X1 U22062 ( .A1(n18995), .A2(n18994), .B1(n19012), .B2(n18993), .ZN(
        n18998) );
  INV_X1 U22063 ( .A(n18996), .ZN(n18997) );
  OAI211_X1 U22064 ( .C1(n19000), .C2(n18999), .A(n18998), .B(n18997), .ZN(
        P3_U2860) );
  NOR2_X1 U22065 ( .A1(n19013), .A2(n19681), .ZN(n19003) );
  AOI211_X1 U22066 ( .C1(n19517), .C2(n19677), .A(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B(n19001), .ZN(n19002) );
  AOI211_X1 U22067 ( .C1(n19004), .C2(n19012), .A(n19003), .B(n19002), .ZN(
        n19008) );
  NOR3_X1 U22068 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n19005), .A3(
        n19014), .ZN(n19010) );
  OAI21_X1 U22069 ( .B1(n19006), .B2(n19010), .A(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n19007) );
  OAI211_X1 U22070 ( .C1(n19009), .C2(n19017), .A(n19008), .B(n19007), .ZN(
        P3_U2861) );
  NOR2_X1 U22071 ( .A1(n19013), .A2(n19687), .ZN(n19011) );
  AOI211_X1 U22072 ( .C1(n19012), .C2(n19018), .A(n19011), .B(n19010), .ZN(
        n19016) );
  OAI211_X1 U22073 ( .C1(n19499), .C2(n19014), .A(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B(n19013), .ZN(n19015) );
  OAI211_X1 U22074 ( .C1(n19018), .C2(n19017), .A(n19016), .B(n19015), .ZN(
        P3_U2862) );
  OAI211_X1 U22075 ( .C1(P3_FLUSH_REG_SCAN_IN), .C2(n19019), .A(
        P3_STATE2_REG_2__SCAN_IN), .B(P3_STATE2_REG_1__SCAN_IN), .ZN(n19541)
         );
  OAI21_X1 U22076 ( .B1(n19022), .B2(n19020), .A(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19021) );
  OAI221_X1 U22077 ( .B1(n19022), .B2(n19541), .C1(n19022), .C2(n19072), .A(
        n19021), .ZN(P3_U2863) );
  NAND2_X1 U22078 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19189) );
  INV_X1 U22079 ( .A(n19023), .ZN(n19024) );
  NOR2_X1 U22080 ( .A1(n19693), .A2(n19024), .ZN(n19026) );
  AOI221_X1 U22081 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n19189), .C1(n19026), 
        .C2(n19189), .A(n19025), .ZN(n19031) );
  NOR2_X1 U22082 ( .A1(n19027), .A2(n19522), .ZN(n19028) );
  OAI21_X1 U22083 ( .B1(n19028), .B2(n19116), .A(n19032), .ZN(n19029) );
  AOI22_X1 U22084 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n19031), .B1(
        n19029), .B2(n19527), .ZN(P3_U2865) );
  INV_X1 U22085 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19530) );
  NAND2_X1 U22086 ( .A1(n19527), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19304) );
  NOR2_X1 U22087 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19527), .ZN(
        n19213) );
  INV_X1 U22088 ( .A(n19213), .ZN(n19214) );
  AND2_X1 U22089 ( .A1(n19304), .A2(n19214), .ZN(n19030) );
  OAI22_X1 U22090 ( .A1(n19031), .A2(n19530), .B1(n19030), .B2(n19029), .ZN(
        P3_U2866) );
  NOR2_X1 U22091 ( .A1(n19531), .A2(n19032), .ZN(P3_U2867) );
  NOR2_X1 U22092 ( .A1(n19530), .A2(n19189), .ZN(n19421) );
  NAND2_X1 U22093 ( .A1(n19421), .A2(n19325), .ZN(n19086) );
  NAND2_X1 U22094 ( .A1(n19423), .A2(BUF2_REG_16__SCAN_IN), .ZN(n19427) );
  NAND2_X1 U22095 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19352) );
  NOR2_X1 U22096 ( .A1(n19352), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19422) );
  NAND2_X1 U22097 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19422), .ZN(
        n19441) );
  INV_X1 U22098 ( .A(n19441), .ZN(n19469) );
  NAND2_X1 U22099 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n19423), .ZN(n19358) );
  INV_X1 U22100 ( .A(n19358), .ZN(n19419) );
  NOR2_X2 U22101 ( .A1(n19065), .A2(n19033), .ZN(n19418) );
  INV_X1 U22102 ( .A(n19550), .ZN(n19417) );
  NAND2_X1 U22103 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19521) );
  NOR2_X2 U22104 ( .A1(n19521), .A2(n19352), .ZN(n19471) );
  NAND2_X1 U22105 ( .A1(n19522), .A2(n19325), .ZN(n19523) );
  NAND2_X1 U22106 ( .A1(n19527), .A2(n19530), .ZN(n19118) );
  NOR2_X2 U22107 ( .A1(n19523), .A2(n19118), .ZN(n19127) );
  NOR2_X1 U22108 ( .A1(n19471), .A2(n19127), .ZN(n19095) );
  NOR2_X1 U22109 ( .A1(n19417), .A2(n19095), .ZN(n19066) );
  AOI22_X1 U22110 ( .A1(n19469), .A2(n19419), .B1(n19418), .B2(n19066), .ZN(
        n19038) );
  NAND2_X1 U22111 ( .A1(n19441), .A2(n19086), .ZN(n19383) );
  AOI211_X1 U22112 ( .C1(P3_STATE2_REG_3__SCAN_IN), .C2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n19095), .B(n19065), .ZN(
        n19034) );
  AOI21_X1 U22113 ( .B1(n19423), .B2(n19383), .A(n19034), .ZN(n19069) );
  NAND2_X1 U22114 ( .A1(n19036), .A2(n19035), .ZN(n19067) );
  NOR2_X2 U22115 ( .A1(n9751), .A2(n19067), .ZN(n19424) );
  AOI22_X1 U22116 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n19069), .B1(
        n19127), .B2(n19424), .ZN(n19037) );
  OAI211_X1 U22117 ( .C1(n19086), .C2(n19427), .A(n19038), .B(n19037), .ZN(
        P3_U2868) );
  NAND2_X1 U22118 ( .A1(BUF2_REG_17__SCAN_IN), .A2(n19423), .ZN(n19433) );
  NAND2_X1 U22119 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n19423), .ZN(n19394) );
  INV_X1 U22120 ( .A(n19394), .ZN(n19429) );
  NOR2_X2 U22121 ( .A1(n19065), .A2(n19039), .ZN(n19428) );
  AOI22_X1 U22122 ( .A1(n19469), .A2(n19429), .B1(n19066), .B2(n19428), .ZN(
        n19042) );
  NOR2_X2 U22123 ( .A1(n19040), .A2(n19067), .ZN(n19430) );
  AOI22_X1 U22124 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n19069), .B1(
        n19127), .B2(n19430), .ZN(n19041) );
  OAI211_X1 U22125 ( .C1(n19086), .C2(n19433), .A(n19042), .B(n19041), .ZN(
        P3_U2869) );
  NAND2_X1 U22126 ( .A1(n19423), .A2(BUF2_REG_18__SCAN_IN), .ZN(n19440) );
  NAND2_X1 U22127 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n19423), .ZN(n19398) );
  INV_X1 U22128 ( .A(n19398), .ZN(n19436) );
  NOR2_X2 U22129 ( .A1(n19065), .A2(n19043), .ZN(n19434) );
  AOI22_X1 U22130 ( .A1(n19469), .A2(n19436), .B1(n19066), .B2(n19434), .ZN(
        n19046) );
  NOR2_X2 U22131 ( .A1(n19044), .A2(n19067), .ZN(n19437) );
  AOI22_X1 U22132 ( .A1(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n19069), .B1(
        n19127), .B2(n19437), .ZN(n19045) );
  OAI211_X1 U22133 ( .C1(n19086), .C2(n19440), .A(n19046), .B(n19045), .ZN(
        P3_U2870) );
  NAND2_X1 U22134 ( .A1(n19423), .A2(BUF2_REG_19__SCAN_IN), .ZN(n19337) );
  NAND2_X1 U22135 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n19423), .ZN(n19447) );
  INV_X1 U22136 ( .A(n19447), .ZN(n19334) );
  NOR2_X2 U22137 ( .A1(n19065), .A2(n19047), .ZN(n19442) );
  AOI22_X1 U22138 ( .A1(n19469), .A2(n19334), .B1(n19066), .B2(n19442), .ZN(
        n19050) );
  NOR2_X2 U22139 ( .A1(n19048), .A2(n19067), .ZN(n19444) );
  AOI22_X1 U22140 ( .A1(P3_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n19069), .B1(
        n19127), .B2(n19444), .ZN(n19049) );
  OAI211_X1 U22141 ( .C1(n19086), .C2(n19337), .A(n19050), .B(n19049), .ZN(
        P3_U2871) );
  NAND2_X1 U22142 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n19423), .ZN(n19453) );
  INV_X1 U22143 ( .A(n19086), .ZN(n19411) );
  NAND2_X1 U22144 ( .A1(n19423), .A2(BUF2_REG_20__SCAN_IN), .ZN(n19405) );
  INV_X1 U22145 ( .A(n19405), .ZN(n19449) );
  NOR2_X2 U22146 ( .A1(n19065), .A2(n19051), .ZN(n19448) );
  AOI22_X1 U22147 ( .A1(n19411), .A2(n19449), .B1(n19066), .B2(n19448), .ZN(
        n19054) );
  NOR2_X2 U22148 ( .A1(n19052), .A2(n19067), .ZN(n19450) );
  AOI22_X1 U22149 ( .A1(P3_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n19069), .B1(
        n19127), .B2(n19450), .ZN(n19053) );
  OAI211_X1 U22150 ( .C1(n19441), .C2(n19453), .A(n19054), .B(n19053), .ZN(
        P3_U2872) );
  NAND2_X1 U22151 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n19423), .ZN(n19459) );
  NAND2_X1 U22152 ( .A1(n19423), .A2(BUF2_REG_21__SCAN_IN), .ZN(n19371) );
  INV_X1 U22153 ( .A(n19371), .ZN(n19455) );
  NOR2_X2 U22154 ( .A1(n19065), .A2(n19055), .ZN(n19454) );
  AOI22_X1 U22155 ( .A1(n19411), .A2(n19455), .B1(n19066), .B2(n19454), .ZN(
        n19058) );
  NOR2_X2 U22156 ( .A1(n19056), .A2(n19067), .ZN(n19456) );
  AOI22_X1 U22157 ( .A1(P3_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n19069), .B1(
        n19127), .B2(n19456), .ZN(n19057) );
  OAI211_X1 U22158 ( .C1(n19441), .C2(n19459), .A(n19058), .B(n19057), .ZN(
        P3_U2873) );
  NAND2_X1 U22159 ( .A1(BUF2_REG_30__SCAN_IN), .A2(n19423), .ZN(n19465) );
  NOR2_X2 U22160 ( .A1(n19065), .A2(n19060), .ZN(n19460) );
  AOI22_X1 U22161 ( .A1(n19411), .A2(n19461), .B1(n19066), .B2(n19460), .ZN(
        n19063) );
  NOR2_X2 U22162 ( .A1(n19061), .A2(n19067), .ZN(n19462) );
  AOI22_X1 U22163 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n19069), .B1(
        n19127), .B2(n19462), .ZN(n19062) );
  OAI211_X1 U22164 ( .C1(n19441), .C2(n19465), .A(n19063), .B(n19062), .ZN(
        P3_U2874) );
  NAND2_X1 U22165 ( .A1(n19423), .A2(BUF2_REG_31__SCAN_IN), .ZN(n19476) );
  NAND2_X1 U22166 ( .A1(n19423), .A2(BUF2_REG_23__SCAN_IN), .ZN(n19382) );
  INV_X1 U22167 ( .A(n19382), .ZN(n19468) );
  NOR2_X2 U22168 ( .A1(n19065), .A2(n19064), .ZN(n19467) );
  AOI22_X1 U22169 ( .A1(n19411), .A2(n19468), .B1(n19066), .B2(n19467), .ZN(
        n19071) );
  NOR2_X2 U22170 ( .A1(n19068), .A2(n19067), .ZN(n19470) );
  AOI22_X1 U22171 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n19069), .B1(
        n19127), .B2(n19470), .ZN(n19070) );
  OAI211_X1 U22172 ( .C1(n19441), .C2(n19476), .A(n19071), .B(n19070), .ZN(
        P3_U2875) );
  INV_X1 U22173 ( .A(n19421), .ZN(n19416) );
  AND2_X1 U22174 ( .A1(n19072), .A2(n19388), .ZN(n19420) );
  NAND2_X1 U22175 ( .A1(n19420), .A2(n19522), .ZN(n19351) );
  OAI22_X1 U22176 ( .A1(n19354), .A2(n19416), .B1(n19118), .B2(n19351), .ZN(
        n19080) );
  INV_X1 U22177 ( .A(n19427), .ZN(n19350) );
  NAND2_X1 U22178 ( .A1(n19522), .A2(n19550), .ZN(n19257) );
  NOR2_X1 U22179 ( .A1(n19118), .A2(n19257), .ZN(n19091) );
  AOI22_X1 U22180 ( .A1(n19471), .A2(n19350), .B1(n19418), .B2(n19091), .ZN(
        n19074) );
  NAND2_X1 U22181 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19522), .ZN(
        n19259) );
  NOR2_X2 U22182 ( .A1(n19118), .A2(n19259), .ZN(n19149) );
  AOI22_X1 U22183 ( .A1(n19411), .A2(n19419), .B1(n19424), .B2(n19149), .ZN(
        n19073) );
  OAI211_X1 U22184 ( .C1(n19075), .C2(n19080), .A(n19074), .B(n19073), .ZN(
        P3_U2876) );
  INV_X1 U22185 ( .A(n19471), .ZN(n19115) );
  AOI22_X1 U22186 ( .A1(n19411), .A2(n19429), .B1(n19428), .B2(n19091), .ZN(
        n19077) );
  INV_X1 U22187 ( .A(n19080), .ZN(n19092) );
  AOI22_X1 U22188 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19092), .B1(
        n19430), .B2(n19149), .ZN(n19076) );
  OAI211_X1 U22189 ( .C1(n19115), .C2(n19433), .A(n19077), .B(n19076), .ZN(
        P3_U2877) );
  INV_X1 U22190 ( .A(n19440), .ZN(n19395) );
  AOI22_X1 U22191 ( .A1(n19471), .A2(n19395), .B1(n19434), .B2(n19091), .ZN(
        n19079) );
  AOI22_X1 U22192 ( .A1(n19411), .A2(n19436), .B1(n19437), .B2(n19149), .ZN(
        n19078) );
  OAI211_X1 U22193 ( .C1(n19081), .C2(n19080), .A(n19079), .B(n19078), .ZN(
        P3_U2878) );
  AOI22_X1 U22194 ( .A1(n19411), .A2(n19334), .B1(n19442), .B2(n19091), .ZN(
        n19083) );
  AOI22_X1 U22195 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19092), .B1(
        n19444), .B2(n19149), .ZN(n19082) );
  OAI211_X1 U22196 ( .C1(n19115), .C2(n19337), .A(n19083), .B(n19082), .ZN(
        P3_U2879) );
  AOI22_X1 U22197 ( .A1(n19471), .A2(n19449), .B1(n19448), .B2(n19091), .ZN(
        n19085) );
  AOI22_X1 U22198 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19092), .B1(
        n19450), .B2(n19149), .ZN(n19084) );
  OAI211_X1 U22199 ( .C1(n19086), .C2(n19453), .A(n19085), .B(n19084), .ZN(
        P3_U2880) );
  INV_X1 U22200 ( .A(n19459), .ZN(n19368) );
  AOI22_X1 U22201 ( .A1(n19411), .A2(n19368), .B1(n19454), .B2(n19091), .ZN(
        n19088) );
  AOI22_X1 U22202 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19092), .B1(
        n19456), .B2(n19149), .ZN(n19087) );
  OAI211_X1 U22203 ( .C1(n19115), .C2(n19371), .A(n19088), .B(n19087), .ZN(
        P3_U2881) );
  INV_X1 U22204 ( .A(n19461), .ZN(n19375) );
  INV_X1 U22205 ( .A(n19465), .ZN(n19372) );
  AOI22_X1 U22206 ( .A1(n19411), .A2(n19372), .B1(n19460), .B2(n19091), .ZN(
        n19090) );
  AOI22_X1 U22207 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19092), .B1(
        n19462), .B2(n19149), .ZN(n19089) );
  OAI211_X1 U22208 ( .C1(n19115), .C2(n19375), .A(n19090), .B(n19089), .ZN(
        P3_U2882) );
  INV_X1 U22209 ( .A(n19476), .ZN(n19378) );
  AOI22_X1 U22210 ( .A1(n19411), .A2(n19378), .B1(n19467), .B2(n19091), .ZN(
        n19094) );
  AOI22_X1 U22211 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19092), .B1(
        n19470), .B2(n19149), .ZN(n19093) );
  OAI211_X1 U22212 ( .C1(n19115), .C2(n19382), .A(n19094), .B(n19093), .ZN(
        P3_U2883) );
  INV_X1 U22213 ( .A(n19127), .ZN(n19138) );
  NOR3_X1 U22214 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19522), .A3(
        n19118), .ZN(n19158) );
  INV_X1 U22215 ( .A(n19158), .ZN(n19180) );
  INV_X1 U22216 ( .A(n19180), .ZN(n19154) );
  INV_X1 U22217 ( .A(n19116), .ZN(n19385) );
  NOR2_X1 U22218 ( .A1(n19149), .A2(n19154), .ZN(n19139) );
  OAI21_X1 U22219 ( .B1(n19095), .B2(n19385), .A(n19139), .ZN(n19096) );
  OAI211_X1 U22220 ( .C1(n19154), .C2(n19651), .A(n19388), .B(n19096), .ZN(
        n19112) );
  NOR2_X1 U22221 ( .A1(n19417), .A2(n19139), .ZN(n19111) );
  AOI22_X1 U22222 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19112), .B1(
        n19418), .B2(n19111), .ZN(n19098) );
  AOI22_X1 U22223 ( .A1(n19471), .A2(n19419), .B1(n19424), .B2(n19158), .ZN(
        n19097) );
  OAI211_X1 U22224 ( .C1(n19138), .C2(n19427), .A(n19098), .B(n19097), .ZN(
        P3_U2884) );
  AOI22_X1 U22225 ( .A1(n19471), .A2(n19429), .B1(n19428), .B2(n19111), .ZN(
        n19100) );
  AOI22_X1 U22226 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19112), .B1(
        n19430), .B2(n19154), .ZN(n19099) );
  OAI211_X1 U22227 ( .C1(n19138), .C2(n19433), .A(n19100), .B(n19099), .ZN(
        P3_U2885) );
  AOI22_X1 U22228 ( .A1(n19127), .A2(n19395), .B1(n19434), .B2(n19111), .ZN(
        n19102) );
  AOI22_X1 U22229 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19112), .B1(
        n19437), .B2(n19154), .ZN(n19101) );
  OAI211_X1 U22230 ( .C1(n19115), .C2(n19398), .A(n19102), .B(n19101), .ZN(
        P3_U2886) );
  INV_X1 U22231 ( .A(n19337), .ZN(n19443) );
  AOI22_X1 U22232 ( .A1(n19127), .A2(n19443), .B1(n19442), .B2(n19111), .ZN(
        n19104) );
  AOI22_X1 U22233 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19112), .B1(
        n19444), .B2(n19154), .ZN(n19103) );
  OAI211_X1 U22234 ( .C1(n19115), .C2(n19447), .A(n19104), .B(n19103), .ZN(
        P3_U2887) );
  AOI22_X1 U22235 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19112), .B1(
        n19448), .B2(n19111), .ZN(n19106) );
  AOI22_X1 U22236 ( .A1(n19127), .A2(n19449), .B1(n19450), .B2(n19154), .ZN(
        n19105) );
  OAI211_X1 U22237 ( .C1(n19115), .C2(n19453), .A(n19106), .B(n19105), .ZN(
        P3_U2888) );
  AOI22_X1 U22238 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19112), .B1(
        n19454), .B2(n19111), .ZN(n19108) );
  AOI22_X1 U22239 ( .A1(n19127), .A2(n19455), .B1(n19456), .B2(n19154), .ZN(
        n19107) );
  OAI211_X1 U22240 ( .C1(n19115), .C2(n19459), .A(n19108), .B(n19107), .ZN(
        P3_U2889) );
  AOI22_X1 U22241 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19112), .B1(
        n19460), .B2(n19111), .ZN(n19110) );
  AOI22_X1 U22242 ( .A1(n19127), .A2(n19461), .B1(n19462), .B2(n19154), .ZN(
        n19109) );
  OAI211_X1 U22243 ( .C1(n19115), .C2(n19465), .A(n19110), .B(n19109), .ZN(
        P3_U2890) );
  AOI22_X1 U22244 ( .A1(n19127), .A2(n19468), .B1(n19467), .B2(n19111), .ZN(
        n19114) );
  AOI22_X1 U22245 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19112), .B1(
        n19470), .B2(n19158), .ZN(n19113) );
  OAI211_X1 U22246 ( .C1(n19115), .C2(n19476), .A(n19114), .B(n19113), .ZN(
        P3_U2891) );
  INV_X1 U22247 ( .A(n19149), .ZN(n19162) );
  AOI22_X1 U22248 ( .A1(n19127), .A2(n19419), .B1(n19418), .B2(n19134), .ZN(
        n19120) );
  INV_X1 U22249 ( .A(n19118), .ZN(n19163) );
  OAI21_X1 U22250 ( .B1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n19116), .A(
        n19388), .ZN(n19117) );
  AOI21_X1 U22251 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n19521), .A(n19117), 
        .ZN(n19212) );
  NAND2_X1 U22252 ( .A1(n19163), .A2(n19212), .ZN(n19135) );
  NOR2_X2 U22253 ( .A1(n19521), .A2(n19118), .ZN(n19204) );
  AOI22_X1 U22254 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19135), .B1(
        n19424), .B2(n19204), .ZN(n19119) );
  OAI211_X1 U22255 ( .C1(n19427), .C2(n19162), .A(n19120), .B(n19119), .ZN(
        P3_U2892) );
  AOI22_X1 U22256 ( .A1(n19127), .A2(n19429), .B1(n19428), .B2(n19134), .ZN(
        n19122) );
  AOI22_X1 U22257 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19135), .B1(
        n19430), .B2(n19204), .ZN(n19121) );
  OAI211_X1 U22258 ( .C1(n19433), .C2(n19162), .A(n19122), .B(n19121), .ZN(
        P3_U2893) );
  AOI22_X1 U22259 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19135), .B1(
        n19434), .B2(n19134), .ZN(n19124) );
  AOI22_X1 U22260 ( .A1(n19395), .A2(n19149), .B1(n19437), .B2(n19204), .ZN(
        n19123) );
  OAI211_X1 U22261 ( .C1(n19138), .C2(n19398), .A(n19124), .B(n19123), .ZN(
        P3_U2894) );
  AOI22_X1 U22262 ( .A1(n19443), .A2(n19149), .B1(n19442), .B2(n19134), .ZN(
        n19126) );
  AOI22_X1 U22263 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19135), .B1(
        n19444), .B2(n19204), .ZN(n19125) );
  OAI211_X1 U22264 ( .C1(n19138), .C2(n19447), .A(n19126), .B(n19125), .ZN(
        P3_U2895) );
  INV_X1 U22265 ( .A(n19453), .ZN(n19402) );
  AOI22_X1 U22266 ( .A1(n19127), .A2(n19402), .B1(n19448), .B2(n19134), .ZN(
        n19129) );
  AOI22_X1 U22267 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19135), .B1(
        n19450), .B2(n19204), .ZN(n19128) );
  OAI211_X1 U22268 ( .C1(n19405), .C2(n19162), .A(n19129), .B(n19128), .ZN(
        P3_U2896) );
  AOI22_X1 U22269 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19135), .B1(
        n19454), .B2(n19134), .ZN(n19131) );
  AOI22_X1 U22270 ( .A1(n19456), .A2(n19204), .B1(n19455), .B2(n19149), .ZN(
        n19130) );
  OAI211_X1 U22271 ( .C1(n19138), .C2(n19459), .A(n19131), .B(n19130), .ZN(
        P3_U2897) );
  AOI22_X1 U22272 ( .A1(n19461), .A2(n19149), .B1(n19460), .B2(n19134), .ZN(
        n19133) );
  AOI22_X1 U22273 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19135), .B1(
        n19462), .B2(n19204), .ZN(n19132) );
  OAI211_X1 U22274 ( .C1(n19138), .C2(n19465), .A(n19133), .B(n19132), .ZN(
        P3_U2898) );
  AOI22_X1 U22275 ( .A1(n19468), .A2(n19149), .B1(n19467), .B2(n19134), .ZN(
        n19137) );
  AOI22_X1 U22276 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19135), .B1(
        n19470), .B2(n19204), .ZN(n19136) );
  OAI211_X1 U22277 ( .C1(n19138), .C2(n19476), .A(n19137), .B(n19136), .ZN(
        P3_U2899) );
  NOR2_X2 U22278 ( .A1(n19523), .A2(n19214), .ZN(n19221) );
  NOR2_X1 U22279 ( .A1(n19204), .A2(n19221), .ZN(n19190) );
  NOR2_X1 U22280 ( .A1(n19417), .A2(n19190), .ZN(n19157) );
  AOI22_X1 U22281 ( .A1(n19350), .A2(n19154), .B1(n19418), .B2(n19157), .ZN(
        n19142) );
  OAI21_X1 U22282 ( .B1(n19139), .B2(n19385), .A(n19190), .ZN(n19140) );
  OAI211_X1 U22283 ( .C1(n19221), .C2(n19651), .A(n19388), .B(n19140), .ZN(
        n19159) );
  AOI22_X1 U22284 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n19159), .B1(
        n19424), .B2(n19221), .ZN(n19141) );
  OAI211_X1 U22285 ( .C1(n19358), .C2(n19162), .A(n19142), .B(n19141), .ZN(
        P3_U2900) );
  INV_X1 U22286 ( .A(n19433), .ZN(n19391) );
  AOI22_X1 U22287 ( .A1(n19391), .A2(n19158), .B1(n19428), .B2(n19157), .ZN(
        n19144) );
  AOI22_X1 U22288 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19159), .B1(
        n19430), .B2(n19221), .ZN(n19143) );
  OAI211_X1 U22289 ( .C1(n19394), .C2(n19162), .A(n19144), .B(n19143), .ZN(
        P3_U2901) );
  AOI22_X1 U22290 ( .A1(n19436), .A2(n19149), .B1(n19434), .B2(n19157), .ZN(
        n19146) );
  AOI22_X1 U22291 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19159), .B1(
        n19437), .B2(n19221), .ZN(n19145) );
  OAI211_X1 U22292 ( .C1(n19440), .C2(n19180), .A(n19146), .B(n19145), .ZN(
        P3_U2902) );
  AOI22_X1 U22293 ( .A1(n19334), .A2(n19149), .B1(n19442), .B2(n19157), .ZN(
        n19148) );
  AOI22_X1 U22294 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19159), .B1(
        n19444), .B2(n19221), .ZN(n19147) );
  OAI211_X1 U22295 ( .C1(n19337), .C2(n19180), .A(n19148), .B(n19147), .ZN(
        P3_U2903) );
  AOI22_X1 U22296 ( .A1(n19402), .A2(n19149), .B1(n19448), .B2(n19157), .ZN(
        n19151) );
  AOI22_X1 U22297 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19159), .B1(
        n19450), .B2(n19221), .ZN(n19150) );
  OAI211_X1 U22298 ( .C1(n19405), .C2(n19180), .A(n19151), .B(n19150), .ZN(
        P3_U2904) );
  AOI22_X1 U22299 ( .A1(n19454), .A2(n19157), .B1(n19455), .B2(n19158), .ZN(
        n19153) );
  AOI22_X1 U22300 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19159), .B1(
        n19456), .B2(n19221), .ZN(n19152) );
  OAI211_X1 U22301 ( .C1(n19459), .C2(n19162), .A(n19153), .B(n19152), .ZN(
        P3_U2905) );
  AOI22_X1 U22302 ( .A1(n19461), .A2(n19154), .B1(n19460), .B2(n19157), .ZN(
        n19156) );
  AOI22_X1 U22303 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19159), .B1(
        n19462), .B2(n19221), .ZN(n19155) );
  OAI211_X1 U22304 ( .C1(n19465), .C2(n19162), .A(n19156), .B(n19155), .ZN(
        P3_U2906) );
  AOI22_X1 U22305 ( .A1(n19468), .A2(n19158), .B1(n19467), .B2(n19157), .ZN(
        n19161) );
  AOI22_X1 U22306 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19159), .B1(
        n19470), .B2(n19221), .ZN(n19160) );
  OAI211_X1 U22307 ( .C1(n19476), .C2(n19162), .A(n19161), .B(n19160), .ZN(
        P3_U2907) );
  NAND2_X1 U22308 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19163), .ZN(
        n19164) );
  OAI22_X1 U22309 ( .A1(n19354), .A2(n19164), .B1(n19214), .B2(n19351), .ZN(
        n19183) );
  NOR2_X1 U22310 ( .A1(n19214), .A2(n19257), .ZN(n19185) );
  AOI22_X1 U22311 ( .A1(n19419), .A2(n19154), .B1(n19418), .B2(n19185), .ZN(
        n19166) );
  NOR2_X2 U22312 ( .A1(n19214), .A2(n19259), .ZN(n19249) );
  AOI22_X1 U22313 ( .A1(n19350), .A2(n19204), .B1(n19424), .B2(n19249), .ZN(
        n19165) );
  OAI211_X1 U22314 ( .C1(n19167), .C2(n19183), .A(n19166), .B(n19165), .ZN(
        P3_U2908) );
  AOI22_X1 U22315 ( .A1(n19429), .A2(n19154), .B1(n19428), .B2(n19185), .ZN(
        n19169) );
  AOI22_X1 U22316 ( .A1(n19391), .A2(n19204), .B1(n19430), .B2(n19249), .ZN(
        n19168) );
  OAI211_X1 U22317 ( .C1(n19170), .C2(n19183), .A(n19169), .B(n19168), .ZN(
        P3_U2909) );
  AOI22_X1 U22318 ( .A1(n19395), .A2(n19204), .B1(n19434), .B2(n19185), .ZN(
        n19172) );
  INV_X1 U22319 ( .A(n19183), .ZN(n19186) );
  AOI22_X1 U22320 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19186), .B1(
        n19437), .B2(n19249), .ZN(n19171) );
  OAI211_X1 U22321 ( .C1(n19398), .C2(n19180), .A(n19172), .B(n19171), .ZN(
        P3_U2910) );
  AOI22_X1 U22322 ( .A1(n19443), .A2(n19204), .B1(n19442), .B2(n19185), .ZN(
        n19174) );
  AOI22_X1 U22323 ( .A1(n19444), .A2(n19249), .B1(n19334), .B2(n19154), .ZN(
        n19173) );
  OAI211_X1 U22324 ( .C1(n19175), .C2(n19183), .A(n19174), .B(n19173), .ZN(
        P3_U2911) );
  AOI22_X1 U22325 ( .A1(n19449), .A2(n19204), .B1(n19448), .B2(n19185), .ZN(
        n19177) );
  AOI22_X1 U22326 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19186), .B1(
        n19450), .B2(n19249), .ZN(n19176) );
  OAI211_X1 U22327 ( .C1(n19453), .C2(n19180), .A(n19177), .B(n19176), .ZN(
        P3_U2912) );
  AOI22_X1 U22328 ( .A1(n19454), .A2(n19185), .B1(n19455), .B2(n19204), .ZN(
        n19179) );
  AOI22_X1 U22329 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19186), .B1(
        n19456), .B2(n19249), .ZN(n19178) );
  OAI211_X1 U22330 ( .C1(n19459), .C2(n19180), .A(n19179), .B(n19178), .ZN(
        P3_U2913) );
  AOI22_X1 U22331 ( .A1(n19372), .A2(n19154), .B1(n19460), .B2(n19185), .ZN(
        n19182) );
  AOI22_X1 U22332 ( .A1(n19462), .A2(n19249), .B1(n19461), .B2(n19204), .ZN(
        n19181) );
  OAI211_X1 U22333 ( .C1(n19184), .C2(n19183), .A(n19182), .B(n19181), .ZN(
        P3_U2914) );
  INV_X1 U22334 ( .A(n19204), .ZN(n19211) );
  AOI22_X1 U22335 ( .A1(n19378), .A2(n19154), .B1(n19467), .B2(n19185), .ZN(
        n19188) );
  AOI22_X1 U22336 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19186), .B1(
        n19470), .B2(n19249), .ZN(n19187) );
  OAI211_X1 U22337 ( .C1(n19382), .C2(n19211), .A(n19188), .B(n19187), .ZN(
        P3_U2915) );
  INV_X1 U22338 ( .A(n19249), .ZN(n19256) );
  NOR2_X1 U22339 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19189), .ZN(
        n19258) );
  NAND2_X1 U22340 ( .A1(n19258), .A2(n19325), .ZN(n19274) );
  AOI21_X1 U22341 ( .B1(n19256), .B2(n19274), .A(n19417), .ZN(n19207) );
  AOI22_X1 U22342 ( .A1(n19350), .A2(n19221), .B1(n19418), .B2(n19207), .ZN(
        n19193) );
  INV_X1 U22343 ( .A(n19274), .ZN(n19276) );
  AOI221_X1 U22344 ( .B1(n19190), .B2(n19256), .C1(n19385), .C2(n19256), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n19191) );
  OAI21_X1 U22345 ( .B1(n19276), .B2(n19191), .A(n19388), .ZN(n19208) );
  AOI22_X1 U22346 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n19208), .B1(
        n19424), .B2(n19276), .ZN(n19192) );
  OAI211_X1 U22347 ( .C1(n19358), .C2(n19211), .A(n19193), .B(n19192), .ZN(
        P3_U2916) );
  INV_X1 U22348 ( .A(n19221), .ZN(n19234) );
  AOI22_X1 U22349 ( .A1(n19429), .A2(n19204), .B1(n19428), .B2(n19207), .ZN(
        n19195) );
  AOI22_X1 U22350 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19208), .B1(
        n19430), .B2(n19276), .ZN(n19194) );
  OAI211_X1 U22351 ( .C1(n19433), .C2(n19234), .A(n19195), .B(n19194), .ZN(
        P3_U2917) );
  AOI22_X1 U22352 ( .A1(n19395), .A2(n19221), .B1(n19434), .B2(n19207), .ZN(
        n19197) );
  AOI22_X1 U22353 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19208), .B1(
        n19437), .B2(n19276), .ZN(n19196) );
  OAI211_X1 U22354 ( .C1(n19398), .C2(n19211), .A(n19197), .B(n19196), .ZN(
        P3_U2918) );
  AOI22_X1 U22355 ( .A1(n19443), .A2(n19221), .B1(n19442), .B2(n19207), .ZN(
        n19199) );
  AOI22_X1 U22356 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19208), .B1(
        n19444), .B2(n19276), .ZN(n19198) );
  OAI211_X1 U22357 ( .C1(n19447), .C2(n19211), .A(n19199), .B(n19198), .ZN(
        P3_U2919) );
  AOI22_X1 U22358 ( .A1(n19402), .A2(n19204), .B1(n19448), .B2(n19207), .ZN(
        n19201) );
  AOI22_X1 U22359 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19208), .B1(
        n19450), .B2(n19276), .ZN(n19200) );
  OAI211_X1 U22360 ( .C1(n19405), .C2(n19234), .A(n19201), .B(n19200), .ZN(
        P3_U2920) );
  AOI22_X1 U22361 ( .A1(n19368), .A2(n19204), .B1(n19454), .B2(n19207), .ZN(
        n19203) );
  AOI22_X1 U22362 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19208), .B1(
        n19456), .B2(n19276), .ZN(n19202) );
  OAI211_X1 U22363 ( .C1(n19371), .C2(n19234), .A(n19203), .B(n19202), .ZN(
        P3_U2921) );
  AOI22_X1 U22364 ( .A1(n19372), .A2(n19204), .B1(n19460), .B2(n19207), .ZN(
        n19206) );
  AOI22_X1 U22365 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19208), .B1(
        n19462), .B2(n19276), .ZN(n19205) );
  OAI211_X1 U22366 ( .C1(n19375), .C2(n19234), .A(n19206), .B(n19205), .ZN(
        P3_U2922) );
  AOI22_X1 U22367 ( .A1(n19468), .A2(n19221), .B1(n19467), .B2(n19207), .ZN(
        n19210) );
  AOI22_X1 U22368 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19208), .B1(
        n19470), .B2(n19276), .ZN(n19209) );
  OAI211_X1 U22369 ( .C1(n19476), .C2(n19211), .A(n19210), .B(n19209), .ZN(
        P3_U2923) );
  AND2_X1 U22370 ( .A1(n19550), .A2(n19258), .ZN(n19230) );
  AOI22_X1 U22371 ( .A1(n19419), .A2(n19221), .B1(n19418), .B2(n19230), .ZN(
        n19216) );
  NAND2_X1 U22372 ( .A1(n19213), .A2(n19212), .ZN(n19231) );
  NOR2_X2 U22373 ( .A1(n19521), .A2(n19214), .ZN(n19298) );
  AOI22_X1 U22374 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19231), .B1(
        n19424), .B2(n19298), .ZN(n19215) );
  OAI211_X1 U22375 ( .C1(n19427), .C2(n19256), .A(n19216), .B(n19215), .ZN(
        P3_U2924) );
  AOI22_X1 U22376 ( .A1(n19429), .A2(n19221), .B1(n19428), .B2(n19230), .ZN(
        n19218) );
  AOI22_X1 U22377 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19231), .B1(
        n19430), .B2(n19298), .ZN(n19217) );
  OAI211_X1 U22378 ( .C1(n19433), .C2(n19256), .A(n19218), .B(n19217), .ZN(
        P3_U2925) );
  AOI22_X1 U22379 ( .A1(n19395), .A2(n19249), .B1(n19434), .B2(n19230), .ZN(
        n19220) );
  AOI22_X1 U22380 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19231), .B1(
        n19437), .B2(n19298), .ZN(n19219) );
  OAI211_X1 U22381 ( .C1(n19398), .C2(n19234), .A(n19220), .B(n19219), .ZN(
        P3_U2926) );
  AOI22_X1 U22382 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19231), .B1(
        n19442), .B2(n19230), .ZN(n19223) );
  AOI22_X1 U22383 ( .A1(n19444), .A2(n19298), .B1(n19334), .B2(n19221), .ZN(
        n19222) );
  OAI211_X1 U22384 ( .C1(n19337), .C2(n19256), .A(n19223), .B(n19222), .ZN(
        P3_U2927) );
  AOI22_X1 U22385 ( .A1(n19449), .A2(n19249), .B1(n19448), .B2(n19230), .ZN(
        n19225) );
  AOI22_X1 U22386 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19231), .B1(
        n19450), .B2(n19298), .ZN(n19224) );
  OAI211_X1 U22387 ( .C1(n19453), .C2(n19234), .A(n19225), .B(n19224), .ZN(
        P3_U2928) );
  AOI22_X1 U22388 ( .A1(n19454), .A2(n19230), .B1(n19455), .B2(n19249), .ZN(
        n19227) );
  AOI22_X1 U22389 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19231), .B1(
        n19456), .B2(n19298), .ZN(n19226) );
  OAI211_X1 U22390 ( .C1(n19459), .C2(n19234), .A(n19227), .B(n19226), .ZN(
        P3_U2929) );
  AOI22_X1 U22391 ( .A1(n19461), .A2(n19249), .B1(n19460), .B2(n19230), .ZN(
        n19229) );
  AOI22_X1 U22392 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19231), .B1(
        n19462), .B2(n19298), .ZN(n19228) );
  OAI211_X1 U22393 ( .C1(n19465), .C2(n19234), .A(n19229), .B(n19228), .ZN(
        P3_U2930) );
  AOI22_X1 U22394 ( .A1(n19468), .A2(n19249), .B1(n19467), .B2(n19230), .ZN(
        n19233) );
  AOI22_X1 U22395 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19231), .B1(
        n19470), .B2(n19298), .ZN(n19232) );
  OAI211_X1 U22396 ( .C1(n19476), .C2(n19234), .A(n19233), .B(n19232), .ZN(
        P3_U2931) );
  NOR2_X2 U22397 ( .A1(n19523), .A2(n19304), .ZN(n19321) );
  NOR2_X1 U22398 ( .A1(n19298), .A2(n19321), .ZN(n19280) );
  NOR2_X1 U22399 ( .A1(n19417), .A2(n19280), .ZN(n19252) );
  AOI22_X1 U22400 ( .A1(n19419), .A2(n19249), .B1(n19418), .B2(n19252), .ZN(
        n19238) );
  NOR2_X1 U22401 ( .A1(n19249), .A2(n19276), .ZN(n19235) );
  OAI21_X1 U22402 ( .B1(n19235), .B2(n19385), .A(n19280), .ZN(n19236) );
  OAI211_X1 U22403 ( .C1(n19321), .C2(n19651), .A(n19388), .B(n19236), .ZN(
        n19253) );
  AOI22_X1 U22404 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19253), .B1(
        n19424), .B2(n19321), .ZN(n19237) );
  OAI211_X1 U22405 ( .C1(n19427), .C2(n19274), .A(n19238), .B(n19237), .ZN(
        P3_U2932) );
  AOI22_X1 U22406 ( .A1(n19429), .A2(n19249), .B1(n19428), .B2(n19252), .ZN(
        n19240) );
  AOI22_X1 U22407 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19253), .B1(
        n19430), .B2(n19321), .ZN(n19239) );
  OAI211_X1 U22408 ( .C1(n19433), .C2(n19274), .A(n19240), .B(n19239), .ZN(
        P3_U2933) );
  AOI22_X1 U22409 ( .A1(n19436), .A2(n19249), .B1(n19434), .B2(n19252), .ZN(
        n19242) );
  AOI22_X1 U22410 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19253), .B1(
        n19437), .B2(n19321), .ZN(n19241) );
  OAI211_X1 U22411 ( .C1(n19440), .C2(n19274), .A(n19242), .B(n19241), .ZN(
        P3_U2934) );
  AOI22_X1 U22412 ( .A1(n19334), .A2(n19249), .B1(n19442), .B2(n19252), .ZN(
        n19244) );
  AOI22_X1 U22413 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19253), .B1(
        n19444), .B2(n19321), .ZN(n19243) );
  OAI211_X1 U22414 ( .C1(n19337), .C2(n19274), .A(n19244), .B(n19243), .ZN(
        P3_U2935) );
  AOI22_X1 U22415 ( .A1(n19449), .A2(n19276), .B1(n19448), .B2(n19252), .ZN(
        n19246) );
  AOI22_X1 U22416 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19253), .B1(
        n19450), .B2(n19321), .ZN(n19245) );
  OAI211_X1 U22417 ( .C1(n19453), .C2(n19256), .A(n19246), .B(n19245), .ZN(
        P3_U2936) );
  AOI22_X1 U22418 ( .A1(n19454), .A2(n19252), .B1(n19455), .B2(n19276), .ZN(
        n19248) );
  AOI22_X1 U22419 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19253), .B1(
        n19456), .B2(n19321), .ZN(n19247) );
  OAI211_X1 U22420 ( .C1(n19459), .C2(n19256), .A(n19248), .B(n19247), .ZN(
        P3_U2937) );
  AOI22_X1 U22421 ( .A1(n19372), .A2(n19249), .B1(n19460), .B2(n19252), .ZN(
        n19251) );
  AOI22_X1 U22422 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19253), .B1(
        n19462), .B2(n19321), .ZN(n19250) );
  OAI211_X1 U22423 ( .C1(n19375), .C2(n19274), .A(n19251), .B(n19250), .ZN(
        P3_U2938) );
  AOI22_X1 U22424 ( .A1(n19468), .A2(n19276), .B1(n19467), .B2(n19252), .ZN(
        n19255) );
  AOI22_X1 U22425 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19253), .B1(
        n19470), .B2(n19321), .ZN(n19254) );
  OAI211_X1 U22426 ( .C1(n19476), .C2(n19256), .A(n19255), .B(n19254), .ZN(
        P3_U2939) );
  INV_X1 U22427 ( .A(n19298), .ZN(n19296) );
  NOR2_X1 U22428 ( .A1(n19304), .A2(n19257), .ZN(n19275) );
  AOI22_X1 U22429 ( .A1(n19419), .A2(n19276), .B1(n19418), .B2(n19275), .ZN(
        n19261) );
  NOR2_X1 U22430 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19304), .ZN(
        n19303) );
  AOI22_X1 U22431 ( .A1(n19423), .A2(n19258), .B1(n19420), .B2(n19303), .ZN(
        n19277) );
  NOR2_X2 U22432 ( .A1(n19304), .A2(n19259), .ZN(n19346) );
  AOI22_X1 U22433 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n19277), .B1(
        n19424), .B2(n19346), .ZN(n19260) );
  OAI211_X1 U22434 ( .C1(n19427), .C2(n19296), .A(n19261), .B(n19260), .ZN(
        P3_U2940) );
  AOI22_X1 U22435 ( .A1(n19429), .A2(n19276), .B1(n19428), .B2(n19275), .ZN(
        n19263) );
  AOI22_X1 U22436 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19277), .B1(
        n19430), .B2(n19346), .ZN(n19262) );
  OAI211_X1 U22437 ( .C1(n19433), .C2(n19296), .A(n19263), .B(n19262), .ZN(
        P3_U2941) );
  AOI22_X1 U22438 ( .A1(n19395), .A2(n19298), .B1(n19434), .B2(n19275), .ZN(
        n19265) );
  AOI22_X1 U22439 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19277), .B1(
        n19437), .B2(n19346), .ZN(n19264) );
  OAI211_X1 U22440 ( .C1(n19398), .C2(n19274), .A(n19265), .B(n19264), .ZN(
        P3_U2942) );
  AOI22_X1 U22441 ( .A1(n19334), .A2(n19276), .B1(n19442), .B2(n19275), .ZN(
        n19267) );
  AOI22_X1 U22442 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19277), .B1(
        n19444), .B2(n19346), .ZN(n19266) );
  OAI211_X1 U22443 ( .C1(n19337), .C2(n19296), .A(n19267), .B(n19266), .ZN(
        P3_U2943) );
  AOI22_X1 U22444 ( .A1(n19402), .A2(n19276), .B1(n19448), .B2(n19275), .ZN(
        n19269) );
  AOI22_X1 U22445 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19277), .B1(
        n19450), .B2(n19346), .ZN(n19268) );
  OAI211_X1 U22446 ( .C1(n19405), .C2(n19296), .A(n19269), .B(n19268), .ZN(
        P3_U2944) );
  AOI22_X1 U22447 ( .A1(n19368), .A2(n19276), .B1(n19454), .B2(n19275), .ZN(
        n19271) );
  AOI22_X1 U22448 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19277), .B1(
        n19456), .B2(n19346), .ZN(n19270) );
  OAI211_X1 U22449 ( .C1(n19371), .C2(n19296), .A(n19271), .B(n19270), .ZN(
        P3_U2945) );
  AOI22_X1 U22450 ( .A1(n19461), .A2(n19298), .B1(n19460), .B2(n19275), .ZN(
        n19273) );
  AOI22_X1 U22451 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19277), .B1(
        n19462), .B2(n19346), .ZN(n19272) );
  OAI211_X1 U22452 ( .C1(n19465), .C2(n19274), .A(n19273), .B(n19272), .ZN(
        P3_U2946) );
  AOI22_X1 U22453 ( .A1(n19378), .A2(n19276), .B1(n19467), .B2(n19275), .ZN(
        n19279) );
  AOI22_X1 U22454 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19277), .B1(
        n19470), .B2(n19346), .ZN(n19278) );
  OAI211_X1 U22455 ( .C1(n19382), .C2(n19296), .A(n19279), .B(n19278), .ZN(
        P3_U2947) );
  NOR2_X1 U22456 ( .A1(n19522), .A2(n19304), .ZN(n19302) );
  INV_X1 U22457 ( .A(n19302), .ZN(n19353) );
  NOR2_X2 U22458 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19353), .ZN(
        n19377) );
  NOR2_X1 U22459 ( .A1(n19346), .A2(n19377), .ZN(n19326) );
  OAI21_X1 U22460 ( .B1(n19280), .B2(n19385), .A(n19326), .ZN(n19281) );
  OAI211_X1 U22461 ( .C1(n19377), .C2(n19651), .A(n19388), .B(n19281), .ZN(
        n19299) );
  NOR2_X1 U22462 ( .A1(n19417), .A2(n19326), .ZN(n19297) );
  AOI22_X1 U22463 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19299), .B1(
        n19418), .B2(n19297), .ZN(n19283) );
  AOI22_X1 U22464 ( .A1(n19350), .A2(n19321), .B1(n19424), .B2(n19377), .ZN(
        n19282) );
  OAI211_X1 U22465 ( .C1(n19358), .C2(n19296), .A(n19283), .B(n19282), .ZN(
        P3_U2948) );
  INV_X1 U22466 ( .A(n19321), .ZN(n19319) );
  AOI22_X1 U22467 ( .A1(n19429), .A2(n19298), .B1(n19428), .B2(n19297), .ZN(
        n19285) );
  AOI22_X1 U22468 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19299), .B1(
        n19430), .B2(n19377), .ZN(n19284) );
  OAI211_X1 U22469 ( .C1(n19433), .C2(n19319), .A(n19285), .B(n19284), .ZN(
        P3_U2949) );
  AOI22_X1 U22470 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19299), .B1(
        n19434), .B2(n19297), .ZN(n19287) );
  AOI22_X1 U22471 ( .A1(n19437), .A2(n19377), .B1(n19436), .B2(n19298), .ZN(
        n19286) );
  OAI211_X1 U22472 ( .C1(n19440), .C2(n19319), .A(n19287), .B(n19286), .ZN(
        P3_U2950) );
  AOI22_X1 U22473 ( .A1(n19334), .A2(n19298), .B1(n19442), .B2(n19297), .ZN(
        n19289) );
  AOI22_X1 U22474 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19299), .B1(
        n19444), .B2(n19377), .ZN(n19288) );
  OAI211_X1 U22475 ( .C1(n19337), .C2(n19319), .A(n19289), .B(n19288), .ZN(
        P3_U2951) );
  AOI22_X1 U22476 ( .A1(n19449), .A2(n19321), .B1(n19448), .B2(n19297), .ZN(
        n19291) );
  AOI22_X1 U22477 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19299), .B1(
        n19450), .B2(n19377), .ZN(n19290) );
  OAI211_X1 U22478 ( .C1(n19453), .C2(n19296), .A(n19291), .B(n19290), .ZN(
        P3_U2952) );
  AOI22_X1 U22479 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19299), .B1(
        n19454), .B2(n19297), .ZN(n19293) );
  AOI22_X1 U22480 ( .A1(n19368), .A2(n19298), .B1(n19456), .B2(n19377), .ZN(
        n19292) );
  OAI211_X1 U22481 ( .C1(n19371), .C2(n19319), .A(n19293), .B(n19292), .ZN(
        P3_U2953) );
  AOI22_X1 U22482 ( .A1(n19461), .A2(n19321), .B1(n19460), .B2(n19297), .ZN(
        n19295) );
  AOI22_X1 U22483 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19299), .B1(
        n19462), .B2(n19377), .ZN(n19294) );
  OAI211_X1 U22484 ( .C1(n19465), .C2(n19296), .A(n19295), .B(n19294), .ZN(
        P3_U2954) );
  AOI22_X1 U22485 ( .A1(n19378), .A2(n19298), .B1(n19467), .B2(n19297), .ZN(
        n19301) );
  AOI22_X1 U22486 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19299), .B1(
        n19470), .B2(n19377), .ZN(n19300) );
  OAI211_X1 U22487 ( .C1(n19382), .C2(n19319), .A(n19301), .B(n19300), .ZN(
        P3_U2955) );
  NOR2_X1 U22488 ( .A1(n19417), .A2(n19353), .ZN(n19320) );
  AOI22_X1 U22489 ( .A1(n19350), .A2(n19346), .B1(n19418), .B2(n19320), .ZN(
        n19306) );
  AOI22_X1 U22490 ( .A1(n19423), .A2(n19303), .B1(n19420), .B2(n19302), .ZN(
        n19322) );
  NOR2_X2 U22491 ( .A1(n19521), .A2(n19304), .ZN(n19401) );
  AOI22_X1 U22492 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19322), .B1(
        n19424), .B2(n19401), .ZN(n19305) );
  OAI211_X1 U22493 ( .C1(n19358), .C2(n19319), .A(n19306), .B(n19305), .ZN(
        P3_U2956) );
  INV_X1 U22494 ( .A(n19346), .ZN(n19344) );
  AOI22_X1 U22495 ( .A1(n19429), .A2(n19321), .B1(n19428), .B2(n19320), .ZN(
        n19308) );
  AOI22_X1 U22496 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19322), .B1(
        n19430), .B2(n19401), .ZN(n19307) );
  OAI211_X1 U22497 ( .C1(n19433), .C2(n19344), .A(n19308), .B(n19307), .ZN(
        P3_U2957) );
  AOI22_X1 U22498 ( .A1(n19436), .A2(n19321), .B1(n19434), .B2(n19320), .ZN(
        n19310) );
  AOI22_X1 U22499 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19322), .B1(
        n19437), .B2(n19401), .ZN(n19309) );
  OAI211_X1 U22500 ( .C1(n19440), .C2(n19344), .A(n19310), .B(n19309), .ZN(
        P3_U2958) );
  AOI22_X1 U22501 ( .A1(n19443), .A2(n19346), .B1(n19442), .B2(n19320), .ZN(
        n19312) );
  AOI22_X1 U22502 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19322), .B1(
        n19444), .B2(n19401), .ZN(n19311) );
  OAI211_X1 U22503 ( .C1(n19447), .C2(n19319), .A(n19312), .B(n19311), .ZN(
        P3_U2959) );
  AOI22_X1 U22504 ( .A1(n19449), .A2(n19346), .B1(n19448), .B2(n19320), .ZN(
        n19314) );
  AOI22_X1 U22505 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19322), .B1(
        n19450), .B2(n19401), .ZN(n19313) );
  OAI211_X1 U22506 ( .C1(n19453), .C2(n19319), .A(n19314), .B(n19313), .ZN(
        P3_U2960) );
  AOI22_X1 U22507 ( .A1(n19454), .A2(n19320), .B1(n19455), .B2(n19346), .ZN(
        n19316) );
  AOI22_X1 U22508 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19322), .B1(
        n19456), .B2(n19401), .ZN(n19315) );
  OAI211_X1 U22509 ( .C1(n19459), .C2(n19319), .A(n19316), .B(n19315), .ZN(
        P3_U2961) );
  AOI22_X1 U22510 ( .A1(n19461), .A2(n19346), .B1(n19460), .B2(n19320), .ZN(
        n19318) );
  AOI22_X1 U22511 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19322), .B1(
        n19462), .B2(n19401), .ZN(n19317) );
  OAI211_X1 U22512 ( .C1(n19465), .C2(n19319), .A(n19318), .B(n19317), .ZN(
        P3_U2962) );
  AOI22_X1 U22513 ( .A1(n19378), .A2(n19321), .B1(n19467), .B2(n19320), .ZN(
        n19324) );
  AOI22_X1 U22514 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19322), .B1(
        n19470), .B2(n19401), .ZN(n19323) );
  OAI211_X1 U22515 ( .C1(n19382), .C2(n19344), .A(n19324), .B(n19323), .ZN(
        P3_U2963) );
  NAND2_X1 U22516 ( .A1(n19325), .A2(n19422), .ZN(n19475) );
  INV_X1 U22517 ( .A(n19475), .ZN(n19435) );
  NOR2_X1 U22518 ( .A1(n19401), .A2(n19435), .ZN(n19386) );
  NOR2_X1 U22519 ( .A1(n19417), .A2(n19386), .ZN(n19345) );
  AOI22_X1 U22520 ( .A1(n19350), .A2(n19377), .B1(n19418), .B2(n19345), .ZN(
        n19329) );
  OAI21_X1 U22521 ( .B1(n19326), .B2(n19385), .A(n19386), .ZN(n19327) );
  OAI211_X1 U22522 ( .C1(n19435), .C2(n19651), .A(n19388), .B(n19327), .ZN(
        n19347) );
  AOI22_X1 U22523 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n19347), .B1(
        n19424), .B2(n19435), .ZN(n19328) );
  OAI211_X1 U22524 ( .C1(n19358), .C2(n19344), .A(n19329), .B(n19328), .ZN(
        P3_U2964) );
  INV_X1 U22525 ( .A(n19377), .ZN(n19365) );
  AOI22_X1 U22526 ( .A1(n19429), .A2(n19346), .B1(n19428), .B2(n19345), .ZN(
        n19331) );
  AOI22_X1 U22527 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n19347), .B1(
        n19430), .B2(n19435), .ZN(n19330) );
  OAI211_X1 U22528 ( .C1(n19433), .C2(n19365), .A(n19331), .B(n19330), .ZN(
        P3_U2965) );
  AOI22_X1 U22529 ( .A1(n19395), .A2(n19377), .B1(n19434), .B2(n19345), .ZN(
        n19333) );
  AOI22_X1 U22530 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n19347), .B1(
        n19437), .B2(n19435), .ZN(n19332) );
  OAI211_X1 U22531 ( .C1(n19398), .C2(n19344), .A(n19333), .B(n19332), .ZN(
        P3_U2966) );
  AOI22_X1 U22532 ( .A1(n19334), .A2(n19346), .B1(n19442), .B2(n19345), .ZN(
        n19336) );
  AOI22_X1 U22533 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19347), .B1(
        n19444), .B2(n19435), .ZN(n19335) );
  OAI211_X1 U22534 ( .C1(n19337), .C2(n19365), .A(n19336), .B(n19335), .ZN(
        P3_U2967) );
  AOI22_X1 U22535 ( .A1(n19449), .A2(n19377), .B1(n19448), .B2(n19345), .ZN(
        n19339) );
  AOI22_X1 U22536 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n19347), .B1(
        n19450), .B2(n19435), .ZN(n19338) );
  OAI211_X1 U22537 ( .C1(n19453), .C2(n19344), .A(n19339), .B(n19338), .ZN(
        P3_U2968) );
  AOI22_X1 U22538 ( .A1(n19454), .A2(n19345), .B1(n19455), .B2(n19377), .ZN(
        n19341) );
  AOI22_X1 U22539 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19347), .B1(
        n19456), .B2(n19435), .ZN(n19340) );
  OAI211_X1 U22540 ( .C1(n19459), .C2(n19344), .A(n19341), .B(n19340), .ZN(
        P3_U2969) );
  AOI22_X1 U22541 ( .A1(n19461), .A2(n19377), .B1(n19460), .B2(n19345), .ZN(
        n19343) );
  AOI22_X1 U22542 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19347), .B1(
        n19462), .B2(n19435), .ZN(n19342) );
  OAI211_X1 U22543 ( .C1(n19465), .C2(n19344), .A(n19343), .B(n19342), .ZN(
        P3_U2970) );
  AOI22_X1 U22544 ( .A1(n19378), .A2(n19346), .B1(n19467), .B2(n19345), .ZN(
        n19349) );
  AOI22_X1 U22545 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n19347), .B1(
        n19470), .B2(n19435), .ZN(n19348) );
  OAI211_X1 U22546 ( .C1(n19382), .C2(n19365), .A(n19349), .B(n19348), .ZN(
        P3_U2971) );
  AND2_X1 U22547 ( .A1(n19550), .A2(n19422), .ZN(n19376) );
  AOI22_X1 U22548 ( .A1(n19350), .A2(n19401), .B1(n19418), .B2(n19376), .ZN(
        n19357) );
  OAI22_X1 U22549 ( .A1(n19354), .A2(n19353), .B1(n19352), .B2(n19351), .ZN(
        n19355) );
  INV_X1 U22550 ( .A(n19355), .ZN(n19379) );
  AOI22_X1 U22551 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n19379), .B1(
        n19469), .B2(n19424), .ZN(n19356) );
  OAI211_X1 U22552 ( .C1(n19358), .C2(n19365), .A(n19357), .B(n19356), .ZN(
        P3_U2972) );
  AOI22_X1 U22553 ( .A1(n19391), .A2(n19401), .B1(n19428), .B2(n19376), .ZN(
        n19360) );
  AOI22_X1 U22554 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19379), .B1(
        n19469), .B2(n19430), .ZN(n19359) );
  OAI211_X1 U22555 ( .C1(n19394), .C2(n19365), .A(n19360), .B(n19359), .ZN(
        P3_U2973) );
  AOI22_X1 U22556 ( .A1(n19395), .A2(n19401), .B1(n19434), .B2(n19376), .ZN(
        n19362) );
  AOI22_X1 U22557 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19379), .B1(
        n19469), .B2(n19437), .ZN(n19361) );
  OAI211_X1 U22558 ( .C1(n19398), .C2(n19365), .A(n19362), .B(n19361), .ZN(
        P3_U2974) );
  AOI22_X1 U22559 ( .A1(n19443), .A2(n19401), .B1(n19442), .B2(n19376), .ZN(
        n19364) );
  AOI22_X1 U22560 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19379), .B1(
        n19469), .B2(n19444), .ZN(n19363) );
  OAI211_X1 U22561 ( .C1(n19447), .C2(n19365), .A(n19364), .B(n19363), .ZN(
        P3_U2975) );
  INV_X1 U22562 ( .A(n19401), .ZN(n19415) );
  AOI22_X1 U22563 ( .A1(n19402), .A2(n19377), .B1(n19448), .B2(n19376), .ZN(
        n19367) );
  AOI22_X1 U22564 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19379), .B1(
        n19469), .B2(n19450), .ZN(n19366) );
  OAI211_X1 U22565 ( .C1(n19405), .C2(n19415), .A(n19367), .B(n19366), .ZN(
        P3_U2976) );
  AOI22_X1 U22566 ( .A1(n19368), .A2(n19377), .B1(n19454), .B2(n19376), .ZN(
        n19370) );
  AOI22_X1 U22567 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19379), .B1(
        n19469), .B2(n19456), .ZN(n19369) );
  OAI211_X1 U22568 ( .C1(n19371), .C2(n19415), .A(n19370), .B(n19369), .ZN(
        P3_U2977) );
  AOI22_X1 U22569 ( .A1(n19372), .A2(n19377), .B1(n19460), .B2(n19376), .ZN(
        n19374) );
  AOI22_X1 U22570 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19379), .B1(
        n19469), .B2(n19462), .ZN(n19373) );
  OAI211_X1 U22571 ( .C1(n19375), .C2(n19415), .A(n19374), .B(n19373), .ZN(
        P3_U2978) );
  AOI22_X1 U22572 ( .A1(n19378), .A2(n19377), .B1(n19467), .B2(n19376), .ZN(
        n19381) );
  AOI22_X1 U22573 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19379), .B1(
        n19469), .B2(n19470), .ZN(n19380) );
  OAI211_X1 U22574 ( .C1(n19382), .C2(n19415), .A(n19381), .B(n19380), .ZN(
        P3_U2979) );
  INV_X1 U22575 ( .A(n19383), .ZN(n19384) );
  NOR2_X1 U22576 ( .A1(n19417), .A2(n19384), .ZN(n19410) );
  AOI22_X1 U22577 ( .A1(n19419), .A2(n19401), .B1(n19418), .B2(n19410), .ZN(
        n19390) );
  OAI21_X1 U22578 ( .B1(n19386), .B2(n19385), .A(n19384), .ZN(n19387) );
  OAI211_X1 U22579 ( .C1(n19411), .C2(n19651), .A(n19388), .B(n19387), .ZN(
        n19412) );
  AOI22_X1 U22580 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n19412), .B1(
        n19411), .B2(n19424), .ZN(n19389) );
  OAI211_X1 U22581 ( .C1(n19427), .C2(n19475), .A(n19390), .B(n19389), .ZN(
        P3_U2980) );
  AOI22_X1 U22582 ( .A1(n19391), .A2(n19435), .B1(n19428), .B2(n19410), .ZN(
        n19393) );
  AOI22_X1 U22583 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n19412), .B1(
        n19411), .B2(n19430), .ZN(n19392) );
  OAI211_X1 U22584 ( .C1(n19394), .C2(n19415), .A(n19393), .B(n19392), .ZN(
        P3_U2981) );
  AOI22_X1 U22585 ( .A1(n19395), .A2(n19435), .B1(n19434), .B2(n19410), .ZN(
        n19397) );
  AOI22_X1 U22586 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n19412), .B1(
        n19411), .B2(n19437), .ZN(n19396) );
  OAI211_X1 U22587 ( .C1(n19398), .C2(n19415), .A(n19397), .B(n19396), .ZN(
        P3_U2982) );
  AOI22_X1 U22588 ( .A1(n19443), .A2(n19435), .B1(n19442), .B2(n19410), .ZN(
        n19400) );
  AOI22_X1 U22589 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n19412), .B1(
        n19411), .B2(n19444), .ZN(n19399) );
  OAI211_X1 U22590 ( .C1(n19447), .C2(n19415), .A(n19400), .B(n19399), .ZN(
        P3_U2983) );
  AOI22_X1 U22591 ( .A1(n19402), .A2(n19401), .B1(n19448), .B2(n19410), .ZN(
        n19404) );
  AOI22_X1 U22592 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n19412), .B1(
        n19411), .B2(n19450), .ZN(n19403) );
  OAI211_X1 U22593 ( .C1(n19405), .C2(n19475), .A(n19404), .B(n19403), .ZN(
        P3_U2984) );
  AOI22_X1 U22594 ( .A1(n19454), .A2(n19410), .B1(n19455), .B2(n19435), .ZN(
        n19407) );
  AOI22_X1 U22595 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n19412), .B1(
        n19411), .B2(n19456), .ZN(n19406) );
  OAI211_X1 U22596 ( .C1(n19459), .C2(n19415), .A(n19407), .B(n19406), .ZN(
        P3_U2985) );
  AOI22_X1 U22597 ( .A1(n19461), .A2(n19435), .B1(n19460), .B2(n19410), .ZN(
        n19409) );
  AOI22_X1 U22598 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n19412), .B1(
        n19411), .B2(n19462), .ZN(n19408) );
  OAI211_X1 U22599 ( .C1(n19465), .C2(n19415), .A(n19409), .B(n19408), .ZN(
        P3_U2986) );
  AOI22_X1 U22600 ( .A1(n19468), .A2(n19435), .B1(n19467), .B2(n19410), .ZN(
        n19414) );
  AOI22_X1 U22601 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n19412), .B1(
        n19411), .B2(n19470), .ZN(n19413) );
  OAI211_X1 U22602 ( .C1(n19476), .C2(n19415), .A(n19414), .B(n19413), .ZN(
        P3_U2987) );
  NOR2_X1 U22603 ( .A1(n19417), .A2(n19416), .ZN(n19466) );
  AOI22_X1 U22604 ( .A1(n19419), .A2(n19435), .B1(n19418), .B2(n19466), .ZN(
        n19426) );
  AOI22_X1 U22605 ( .A1(n19423), .A2(n19422), .B1(n19421), .B2(n19420), .ZN(
        n19472) );
  AOI22_X1 U22606 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n19472), .B1(
        n19471), .B2(n19424), .ZN(n19425) );
  OAI211_X1 U22607 ( .C1(n19441), .C2(n19427), .A(n19426), .B(n19425), .ZN(
        P3_U2988) );
  AOI22_X1 U22608 ( .A1(n19429), .A2(n19435), .B1(n19428), .B2(n19466), .ZN(
        n19432) );
  AOI22_X1 U22609 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n19472), .B1(
        n19471), .B2(n19430), .ZN(n19431) );
  OAI211_X1 U22610 ( .C1(n19441), .C2(n19433), .A(n19432), .B(n19431), .ZN(
        P3_U2989) );
  AOI22_X1 U22611 ( .A1(n19436), .A2(n19435), .B1(n19434), .B2(n19466), .ZN(
        n19439) );
  AOI22_X1 U22612 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n19472), .B1(
        n19471), .B2(n19437), .ZN(n19438) );
  OAI211_X1 U22613 ( .C1(n19441), .C2(n19440), .A(n19439), .B(n19438), .ZN(
        P3_U2990) );
  AOI22_X1 U22614 ( .A1(n19469), .A2(n19443), .B1(n19442), .B2(n19466), .ZN(
        n19446) );
  AOI22_X1 U22615 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n19472), .B1(
        n19471), .B2(n19444), .ZN(n19445) );
  OAI211_X1 U22616 ( .C1(n19447), .C2(n19475), .A(n19446), .B(n19445), .ZN(
        P3_U2991) );
  AOI22_X1 U22617 ( .A1(n19469), .A2(n19449), .B1(n19448), .B2(n19466), .ZN(
        n19452) );
  AOI22_X1 U22618 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n19472), .B1(
        n19471), .B2(n19450), .ZN(n19451) );
  OAI211_X1 U22619 ( .C1(n19453), .C2(n19475), .A(n19452), .B(n19451), .ZN(
        P3_U2992) );
  AOI22_X1 U22620 ( .A1(n19469), .A2(n19455), .B1(n19454), .B2(n19466), .ZN(
        n19458) );
  AOI22_X1 U22621 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19472), .B1(
        n19471), .B2(n19456), .ZN(n19457) );
  OAI211_X1 U22622 ( .C1(n19459), .C2(n19475), .A(n19458), .B(n19457), .ZN(
        P3_U2993) );
  AOI22_X1 U22623 ( .A1(n19469), .A2(n19461), .B1(n19460), .B2(n19466), .ZN(
        n19464) );
  AOI22_X1 U22624 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19472), .B1(
        n19471), .B2(n19462), .ZN(n19463) );
  OAI211_X1 U22625 ( .C1(n19465), .C2(n19475), .A(n19464), .B(n19463), .ZN(
        P3_U2994) );
  AOI22_X1 U22626 ( .A1(n19469), .A2(n19468), .B1(n19467), .B2(n19466), .ZN(
        n19474) );
  AOI22_X1 U22627 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n19472), .B1(
        n19471), .B2(n19470), .ZN(n19473) );
  OAI211_X1 U22628 ( .C1(n19476), .C2(n19475), .A(n19474), .B(n19473), .ZN(
        P3_U2995) );
  NAND2_X1 U22629 ( .A1(n19477), .A2(n19501), .ZN(n19478) );
  AOI22_X1 U22630 ( .A1(n19481), .A2(n19480), .B1(n19479), .B2(n19478), .ZN(
        n19482) );
  OAI221_X1 U22631 ( .B1(n19484), .B2(n19509), .C1(n19484), .C2(n19483), .A(
        n19482), .ZN(n19692) );
  OAI21_X1 U22632 ( .B1(P3_MORE_REG_SCAN_IN), .B2(P3_FLUSH_REG_SCAN_IN), .A(
        n19485), .ZN(n19486) );
  OAI211_X1 U22633 ( .C1(n19514), .C2(n19488), .A(n19487), .B(n19486), .ZN(
        n19536) );
  INV_X1 U22634 ( .A(n19512), .ZN(n19490) );
  NAND2_X1 U22635 ( .A1(n19517), .A2(n12663), .ZN(n19518) );
  NAND2_X1 U22636 ( .A1(n19666), .A2(n19506), .ZN(n19495) );
  AOI22_X1 U22637 ( .A1(n19490), .A2(n19518), .B1(n19489), .B2(n19495), .ZN(
        n19491) );
  NOR2_X1 U22638 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n19491), .ZN(
        n19653) );
  OAI21_X1 U22639 ( .B1(n19494), .B2(n19493), .A(n19492), .ZN(n19504) );
  INV_X1 U22640 ( .A(n19504), .ZN(n19496) );
  OAI21_X1 U22641 ( .B1(n19497), .B2(n19496), .A(n19495), .ZN(n19498) );
  AOI21_X1 U22642 ( .B1(n19512), .B2(n19499), .A(n19498), .ZN(n19654) );
  NAND2_X1 U22643 ( .A1(n19514), .A2(n19654), .ZN(n19500) );
  AOI22_X1 U22644 ( .A1(n19514), .A2(n19653), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n19500), .ZN(n19534) );
  INV_X1 U22645 ( .A(n19514), .ZN(n19525) );
  AOI21_X1 U22646 ( .B1(n19666), .B2(n19674), .A(n19501), .ZN(n19513) );
  NAND2_X1 U22647 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n19515), .ZN(
        n19502) );
  AOI211_X1 U22648 ( .C1(n19503), .C2(n19502), .A(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n19674), .ZN(n19511) );
  AOI21_X1 U22649 ( .B1(n19674), .B2(n19505), .A(n19504), .ZN(n19508) );
  NAND2_X1 U22650 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n19506), .ZN(
        n19507) );
  OAI22_X1 U22651 ( .A1(n19663), .A2(n19509), .B1(n19508), .B2(n19507), .ZN(
        n19510) );
  AOI211_X1 U22652 ( .C1(n19513), .C2(n19512), .A(n19511), .B(n19510), .ZN(
        n19659) );
  AOI22_X1 U22653 ( .A1(n19525), .A2(n19666), .B1(n19659), .B2(n19514), .ZN(
        n19529) );
  NOR2_X1 U22654 ( .A1(n19516), .A2(n19515), .ZN(n19520) );
  AOI22_X1 U22655 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n19517), .B1(
        n19520), .B2(n12663), .ZN(n19676) );
  INV_X1 U22656 ( .A(n19518), .ZN(n19519) );
  OAI22_X1 U22657 ( .A1(n19520), .A2(n19667), .B1(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n19519), .ZN(n19672) );
  AOI222_X1 U22658 ( .A1(n19676), .A2(n19672), .B1(n19676), .B2(n19522), .C1(
        n19672), .C2(n19521), .ZN(n19524) );
  OAI21_X1 U22659 ( .B1(n19525), .B2(n19524), .A(n19523), .ZN(n19528) );
  AND2_X1 U22660 ( .A1(n19529), .A2(n19528), .ZN(n19526) );
  OAI221_X1 U22661 ( .B1(n19529), .B2(n19528), .C1(n19527), .C2(n19526), .A(
        n19531), .ZN(n19533) );
  AOI21_X1 U22662 ( .B1(n19531), .B2(n19530), .A(n19529), .ZN(n19532) );
  AOI222_X1 U22663 ( .A1(n19534), .A2(n19533), .B1(n19534), .B2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C1(n19533), .C2(n19532), .ZN(
        n19535) );
  NOR4_X1 U22664 ( .A1(n19537), .A2(n19692), .A3(n19536), .A4(n19535), .ZN(
        n19547) );
  OAI211_X1 U22665 ( .C1(n19539), .C2(n19538), .A(n19694), .B(n19547), .ZN(
        n19650) );
  INV_X1 U22666 ( .A(n19650), .ZN(n19540) );
  AOI21_X1 U22667 ( .B1(n19696), .B2(n19712), .A(n19540), .ZN(n19551) );
  OAI211_X1 U22668 ( .C1(P3_STATE2_REG_1__SCAN_IN), .C2(n19550), .A(n19551), 
        .B(n19541), .ZN(n19544) );
  AOI22_X1 U22669 ( .A1(n19675), .A2(n19703), .B1(n19696), .B2(n19548), .ZN(
        n19543) );
  AOI22_X1 U22670 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n19544), .B1(n19543), 
        .B2(n19542), .ZN(n19545) );
  OAI21_X1 U22671 ( .B1(n19547), .B2(n19546), .A(n19545), .ZN(P3_U2996) );
  NAND2_X1 U22672 ( .A1(n19696), .A2(n19548), .ZN(n19554) );
  NAND4_X1 U22673 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(
        P3_STATE2_REG_1__SCAN_IN), .A3(n19696), .A4(n19712), .ZN(n19557) );
  INV_X1 U22674 ( .A(n19549), .ZN(n19552) );
  NAND3_X1 U22675 ( .A1(n19552), .A2(n19551), .A3(n19550), .ZN(n19553) );
  NAND4_X1 U22676 ( .A1(n19555), .A2(n19554), .A3(n19557), .A4(n19553), .ZN(
        P3_U2997) );
  OAI21_X1 U22677 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(
        P3_STATEBS16_REG_SCAN_IN), .A(n19556), .ZN(n19559) );
  INV_X1 U22678 ( .A(n19557), .ZN(n19558) );
  AOI21_X1 U22679 ( .B1(n19560), .B2(n19559), .A(n19558), .ZN(P3_U2998) );
  AND2_X1 U22680 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n19562), .ZN(
        P3_U2999) );
  AND2_X1 U22681 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n19562), .ZN(
        P3_U3000) );
  AND2_X1 U22682 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n19562), .ZN(
        P3_U3001) );
  AND2_X1 U22683 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n19562), .ZN(
        P3_U3002) );
  AND2_X1 U22684 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n19562), .ZN(
        P3_U3003) );
  AND2_X1 U22685 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n19562), .ZN(
        P3_U3004) );
  AND2_X1 U22686 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n19562), .ZN(
        P3_U3005) );
  AND2_X1 U22687 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n19562), .ZN(
        P3_U3006) );
  NOR2_X1 U22688 ( .A1(n19561), .A2(n19648), .ZN(P3_U3007) );
  AND2_X1 U22689 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n19562), .ZN(
        P3_U3008) );
  AND2_X1 U22690 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n19562), .ZN(
        P3_U3009) );
  AND2_X1 U22691 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n19562), .ZN(
        P3_U3010) );
  AND2_X1 U22692 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n19562), .ZN(
        P3_U3011) );
  AND2_X1 U22693 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n19562), .ZN(
        P3_U3012) );
  AND2_X1 U22694 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n19562), .ZN(
        P3_U3013) );
  AND2_X1 U22695 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n19562), .ZN(
        P3_U3014) );
  AND2_X1 U22696 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n19562), .ZN(
        P3_U3015) );
  AND2_X1 U22697 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n19562), .ZN(
        P3_U3016) );
  AND2_X1 U22698 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n19562), .ZN(
        P3_U3017) );
  AND2_X1 U22699 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n19562), .ZN(
        P3_U3018) );
  AND2_X1 U22700 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n19562), .ZN(
        P3_U3019) );
  AND2_X1 U22701 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n19562), .ZN(
        P3_U3020) );
  AND2_X1 U22702 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n19562), .ZN(P3_U3021) );
  AND2_X1 U22703 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n19562), .ZN(P3_U3022) );
  AND2_X1 U22704 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n19562), .ZN(P3_U3023) );
  AND2_X1 U22705 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n19562), .ZN(P3_U3024) );
  AND2_X1 U22706 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n19562), .ZN(P3_U3025) );
  AND2_X1 U22707 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n19562), .ZN(P3_U3026) );
  AND2_X1 U22708 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n19562), .ZN(P3_U3027) );
  AND2_X1 U22709 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n19562), .ZN(P3_U3028) );
  OAI21_X1 U22710 ( .B1(n19563), .B2(n21186), .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n19564) );
  AOI22_X1 U22711 ( .A1(n19577), .A2(n19578), .B1(n19708), .B2(n19564), .ZN(
        n19566) );
  NAND3_X1 U22712 ( .A1(NA), .A2(n19577), .A3(n19565), .ZN(n19573) );
  OAI211_X1 U22713 ( .C1(n19701), .C2(n19569), .A(n19566), .B(n19573), .ZN(
        P3_U3029) );
  NOR2_X1 U22714 ( .A1(n19578), .A2(n21186), .ZN(n19572) );
  NOR2_X1 U22715 ( .A1(n19577), .A2(n19572), .ZN(n19567) );
  NAND2_X1 U22716 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(n19696), .ZN(n19570) );
  INV_X1 U22717 ( .A(n19570), .ZN(n19574) );
  AOI21_X1 U22718 ( .B1(n19567), .B2(P3_REQUESTPENDING_REG_SCAN_IN), .A(n19574), .ZN(n19568) );
  OAI211_X1 U22719 ( .C1(n21186), .C2(n19569), .A(n19568), .B(n19698), .ZN(
        P3_U3030) );
  OAI22_X1 U22720 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(
        P3_REQUESTPENDING_REG_SCAN_IN), .B1(NA), .B2(n19570), .ZN(n19571) );
  OAI22_X1 U22721 ( .A1(n19572), .A2(n19571), .B1(
        P3_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .ZN(n19576) );
  OAI211_X1 U22722 ( .C1(n19574), .C2(n19577), .A(n19573), .B(
        P3_STATE_REG_2__SCAN_IN), .ZN(n19575) );
  OAI21_X1 U22723 ( .B1(n19577), .B2(n19576), .A(n19575), .ZN(P3_U3031) );
  OAI222_X1 U22724 ( .A1(n19640), .A2(n19681), .B1(n19579), .B2(n19710), .C1(
        n19580), .C2(n19636), .ZN(P3_U3032) );
  OAI222_X1 U22725 ( .A1(n19636), .A2(n19582), .B1(n19581), .B2(n19710), .C1(
        n19580), .C2(n19640), .ZN(P3_U3033) );
  OAI222_X1 U22726 ( .A1(n19636), .A2(n19584), .B1(n19583), .B2(n19710), .C1(
        n19582), .C2(n19640), .ZN(P3_U3034) );
  INV_X1 U22727 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n19586) );
  OAI222_X1 U22728 ( .A1(n19636), .A2(n19586), .B1(n19585), .B2(n19710), .C1(
        n19584), .C2(n19640), .ZN(P3_U3035) );
  OAI222_X1 U22729 ( .A1(n19636), .A2(n19588), .B1(n19587), .B2(n19710), .C1(
        n19586), .C2(n19640), .ZN(P3_U3036) );
  OAI222_X1 U22730 ( .A1(n19636), .A2(n19590), .B1(n19589), .B2(n19710), .C1(
        n19588), .C2(n19640), .ZN(P3_U3037) );
  INV_X1 U22731 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n19593) );
  OAI222_X1 U22732 ( .A1(n19636), .A2(n19593), .B1(n19591), .B2(n19710), .C1(
        n19590), .C2(n19640), .ZN(P3_U3038) );
  OAI222_X1 U22733 ( .A1(n19593), .A2(n19640), .B1(n19592), .B2(n19710), .C1(
        n19594), .C2(n19636), .ZN(P3_U3039) );
  OAI222_X1 U22734 ( .A1(n19636), .A2(n19596), .B1(n19595), .B2(n19710), .C1(
        n19594), .C2(n19640), .ZN(P3_U3040) );
  OAI222_X1 U22735 ( .A1(n19636), .A2(n19598), .B1(n19597), .B2(n19710), .C1(
        n19596), .C2(n19640), .ZN(P3_U3041) );
  INV_X1 U22736 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n19600) );
  OAI222_X1 U22737 ( .A1(n19636), .A2(n19600), .B1(n19599), .B2(n19710), .C1(
        n19598), .C2(n19640), .ZN(P3_U3042) );
  OAI222_X1 U22738 ( .A1(n19636), .A2(n19602), .B1(n19601), .B2(n19710), .C1(
        n19600), .C2(n19640), .ZN(P3_U3043) );
  OAI222_X1 U22739 ( .A1(n19636), .A2(n19604), .B1(n19603), .B2(n19710), .C1(
        n19602), .C2(n19640), .ZN(P3_U3044) );
  OAI222_X1 U22740 ( .A1(n19636), .A2(n19606), .B1(n19605), .B2(n19710), .C1(
        n19604), .C2(n19640), .ZN(P3_U3045) );
  OAI222_X1 U22741 ( .A1(n19636), .A2(n19608), .B1(n19607), .B2(n19710), .C1(
        n19606), .C2(n19640), .ZN(P3_U3046) );
  OAI222_X1 U22742 ( .A1(n19636), .A2(n19611), .B1(n19609), .B2(n19710), .C1(
        n19608), .C2(n19640), .ZN(P3_U3047) );
  OAI222_X1 U22743 ( .A1(n19611), .A2(n19640), .B1(n19610), .B2(n19710), .C1(
        n19612), .C2(n19636), .ZN(P3_U3048) );
  OAI222_X1 U22744 ( .A1(n19636), .A2(n19614), .B1(n19613), .B2(n19710), .C1(
        n19612), .C2(n19640), .ZN(P3_U3049) );
  OAI222_X1 U22745 ( .A1(n19636), .A2(n19617), .B1(n19615), .B2(n19710), .C1(
        n19614), .C2(n19640), .ZN(P3_U3050) );
  INV_X1 U22746 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n19618) );
  OAI222_X1 U22747 ( .A1(n19617), .A2(n19640), .B1(n19616), .B2(n19710), .C1(
        n19618), .C2(n19636), .ZN(P3_U3051) );
  INV_X1 U22748 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n19620) );
  OAI222_X1 U22749 ( .A1(n19636), .A2(n19620), .B1(n19619), .B2(n19710), .C1(
        n19618), .C2(n19640), .ZN(P3_U3052) );
  OAI222_X1 U22750 ( .A1(n19636), .A2(n19623), .B1(n19621), .B2(n19710), .C1(
        n19620), .C2(n19640), .ZN(P3_U3053) );
  OAI222_X1 U22751 ( .A1(n19623), .A2(n19640), .B1(n19622), .B2(n19710), .C1(
        n19624), .C2(n19636), .ZN(P3_U3054) );
  OAI222_X1 U22752 ( .A1(n19636), .A2(n19626), .B1(n19625), .B2(n19710), .C1(
        n19624), .C2(n19640), .ZN(P3_U3055) );
  OAI222_X1 U22753 ( .A1(n19636), .A2(n19628), .B1(n19627), .B2(n19710), .C1(
        n19626), .C2(n19640), .ZN(P3_U3056) );
  OAI222_X1 U22754 ( .A1(n19636), .A2(n19630), .B1(n19629), .B2(n19710), .C1(
        n19628), .C2(n19640), .ZN(P3_U3057) );
  INV_X1 U22755 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n19633) );
  OAI222_X1 U22756 ( .A1(n19636), .A2(n19633), .B1(n19631), .B2(n19710), .C1(
        n19630), .C2(n19640), .ZN(P3_U3058) );
  OAI222_X1 U22757 ( .A1(n19633), .A2(n19640), .B1(n19632), .B2(n19710), .C1(
        n19634), .C2(n19636), .ZN(P3_U3059) );
  OAI222_X1 U22758 ( .A1(n19636), .A2(n19639), .B1(n19635), .B2(n19710), .C1(
        n19634), .C2(n19640), .ZN(P3_U3060) );
  OAI222_X1 U22759 ( .A1(n19640), .A2(n19639), .B1(n19638), .B2(n19710), .C1(
        n19637), .C2(n19636), .ZN(P3_U3061) );
  MUX2_X1 U22760 ( .A(P3_BE_N_REG_3__SCAN_IN), .B(P3_BYTEENABLE_REG_3__SCAN_IN), .S(n19710), .Z(P3_U3274) );
  INV_X1 U22761 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n19684) );
  INV_X1 U22762 ( .A(P3_BE_N_REG_2__SCAN_IN), .ZN(n19641) );
  AOI22_X1 U22763 ( .A1(n19710), .A2(n19684), .B1(n19641), .B2(n19708), .ZN(
        P3_U3275) );
  INV_X1 U22764 ( .A(P3_BE_N_REG_1__SCAN_IN), .ZN(n19642) );
  AOI22_X1 U22765 ( .A1(n19710), .A2(n19643), .B1(n19642), .B2(n19708), .ZN(
        P3_U3276) );
  INV_X1 U22766 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n19689) );
  INV_X1 U22767 ( .A(P3_BE_N_REG_0__SCAN_IN), .ZN(n19644) );
  AOI22_X1 U22768 ( .A1(n19710), .A2(n19689), .B1(n19644), .B2(n19708), .ZN(
        P3_U3277) );
  OAI21_X1 U22769 ( .B1(n19648), .B2(P3_DATAWIDTH_REG_0__SCAN_IN), .A(n19646), 
        .ZN(n19645) );
  INV_X1 U22770 ( .A(n19645), .ZN(P3_U3280) );
  INV_X1 U22771 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n19647) );
  OAI21_X1 U22772 ( .B1(n19648), .B2(n19647), .A(n19646), .ZN(P3_U3281) );
  OAI221_X1 U22773 ( .B1(n19651), .B2(P3_STATE2_REG_0__SCAN_IN), .C1(n19651), 
        .C2(n19650), .A(n19649), .ZN(P3_U3282) );
  AOI22_X1 U22774 ( .A1(n19713), .A2(n19653), .B1(n19675), .B2(n19652), .ZN(
        n19658) );
  INV_X1 U22775 ( .A(n19654), .ZN(n19655) );
  AOI21_X1 U22776 ( .B1(n19713), .B2(n19655), .A(n19680), .ZN(n19657) );
  OAI22_X1 U22777 ( .A1(n19680), .A2(n19658), .B1(n19657), .B2(n19656), .ZN(
        P3_U3285) );
  INV_X1 U22778 ( .A(n19659), .ZN(n19664) );
  NOR2_X1 U22779 ( .A1(n19660), .A2(n19677), .ZN(n19669) );
  AOI22_X1 U22780 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n19662), .B2(n19661), .ZN(
        n19668) );
  AOI222_X1 U22781 ( .A1(n19664), .A2(n19713), .B1(n19669), .B2(n19668), .C1(
        n19675), .C2(n19663), .ZN(n19665) );
  INV_X1 U22782 ( .A(n19680), .ZN(n19678) );
  AOI22_X1 U22783 ( .A1(n19680), .A2(n19666), .B1(n19665), .B2(n19678), .ZN(
        P3_U3288) );
  INV_X1 U22784 ( .A(n19667), .ZN(n19671) );
  INV_X1 U22785 ( .A(n19668), .ZN(n19670) );
  AOI222_X1 U22786 ( .A1(n19672), .A2(n19713), .B1(n19675), .B2(n19671), .C1(
        n19670), .C2(n19669), .ZN(n19673) );
  AOI22_X1 U22787 ( .A1(n19680), .A2(n19674), .B1(n19673), .B2(n19678), .ZN(
        P3_U3289) );
  AOI222_X1 U22788 ( .A1(n19677), .A2(P3_STATE2_REG_1__SCAN_IN), .B1(n19713), 
        .B2(n19676), .C1(n12663), .C2(n19675), .ZN(n19679) );
  AOI22_X1 U22789 ( .A1(n19680), .A2(n12663), .B1(n19679), .B2(n19678), .ZN(
        P3_U3290) );
  AOI21_X1 U22790 ( .B1(P3_DATAWIDTH_REG_0__SCAN_IN), .B2(
        P3_REIP_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n19682)
         );
  OAI221_X1 U22791 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n19682), .C1(n19681), 
        .C2(P3_REIP_REG_0__SCAN_IN), .A(n19685), .ZN(n19683) );
  OAI21_X1 U22792 ( .B1(n19685), .B2(n19684), .A(n19683), .ZN(P3_U3292) );
  NOR2_X1 U22793 ( .A1(n19688), .A2(P3_REIP_REG_1__SCAN_IN), .ZN(n19686) );
  AOI22_X1 U22794 ( .A1(n19689), .A2(n19688), .B1(n19687), .B2(n19686), .ZN(
        P3_U3293) );
  INV_X1 U22795 ( .A(P3_W_R_N_REG_SCAN_IN), .ZN(n19690) );
  AOI22_X1 U22796 ( .A1(n19710), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n19690), 
        .B2(n19708), .ZN(P3_U3294) );
  MUX2_X1 U22797 ( .A(P3_MORE_REG_SCAN_IN), .B(n19692), .S(n19691), .Z(
        P3_U3295) );
  OAI22_X1 U22798 ( .A1(n19696), .A2(n19695), .B1(n19694), .B2(n19693), .ZN(
        n19697) );
  NOR2_X1 U22799 ( .A1(n19715), .A2(n19697), .ZN(n19707) );
  AOI21_X1 U22800 ( .B1(n9752), .B2(n19699), .A(n19698), .ZN(n19702) );
  OAI211_X1 U22801 ( .C1(n19702), .C2(n19711), .A(P3_STATE2_REG_2__SCAN_IN), 
        .B(n19701), .ZN(n19704) );
  AOI21_X1 U22802 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n19704), .A(n19703), 
        .ZN(n19706) );
  NAND2_X1 U22803 ( .A1(n19707), .A2(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n19705) );
  OAI21_X1 U22804 ( .B1(n19707), .B2(n19706), .A(n19705), .ZN(P3_U3296) );
  INV_X1 U22805 ( .A(P3_MEMORYFETCH_REG_SCAN_IN), .ZN(n19718) );
  INV_X1 U22806 ( .A(P3_M_IO_N_REG_SCAN_IN), .ZN(n19709) );
  AOI22_X1 U22807 ( .A1(n19710), .A2(n19718), .B1(n19709), .B2(n19708), .ZN(
        P3_U3297) );
  INV_X1 U22808 ( .A(n19711), .ZN(n19716) );
  AOI21_X1 U22809 ( .B1(n19713), .B2(n19712), .A(n19715), .ZN(n19719) );
  INV_X1 U22810 ( .A(P3_READREQUEST_REG_SCAN_IN), .ZN(n19714) );
  AOI22_X1 U22811 ( .A1(n19716), .A2(n19715), .B1(n19719), .B2(n19714), .ZN(
        P3_U3298) );
  AOI21_X1 U22812 ( .B1(n19719), .B2(n19718), .A(n19717), .ZN(P3_U3299) );
  INV_X1 U22813 ( .A(P2_ADS_N_REG_SCAN_IN), .ZN(n19721) );
  NAND2_X1 U22814 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n20636), .ZN(n20629) );
  NAND2_X1 U22815 ( .A1(n20625), .A2(n19720), .ZN(n20626) );
  OAI21_X1 U22816 ( .B1(n20625), .B2(n20629), .A(n20626), .ZN(n20694) );
  INV_X1 U22817 ( .A(n20694), .ZN(n20619) );
  OAI21_X1 U22818 ( .B1(n20625), .B2(n19721), .A(n20619), .ZN(P2_U2815) );
  INV_X1 U22819 ( .A(P2_CODEFETCH_REG_SCAN_IN), .ZN(n19722) );
  OAI22_X1 U22820 ( .A1(n20745), .A2(n19722), .B1(n20696), .B2(n20610), .ZN(
        P2_U2816) );
  AOI21_X1 U22821 ( .B1(n20625), .B2(n20636), .A(P2_D_C_N_REG_SCAN_IN), .ZN(
        n19723) );
  AOI22_X1 U22822 ( .A1(n20765), .A2(P2_CODEFETCH_REG_SCAN_IN), .B1(n19723), 
        .B2(n20762), .ZN(P2_U2817) );
  INV_X1 U22823 ( .A(n20630), .ZN(n19724) );
  OAI21_X1 U22824 ( .B1(n19724), .B2(BS16), .A(n20694), .ZN(n20692) );
  OAI21_X1 U22825 ( .B1(n20694), .B2(n11033), .A(n20692), .ZN(P2_U2818) );
  NOR4_X1 U22826 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_13__SCAN_IN), .A3(P2_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_15__SCAN_IN), .ZN(n19734) );
  NOR4_X1 U22827 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_7__SCAN_IN), .A3(P2_DATAWIDTH_REG_9__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_10__SCAN_IN), .ZN(n19733) );
  AOI211_X1 U22828 ( .C1(P2_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_1__SCAN_IN), .A(P2_DATAWIDTH_REG_4__SCAN_IN), .B(
        P2_DATAWIDTH_REG_5__SCAN_IN), .ZN(n19725) );
  NAND3_X1 U22829 ( .A1(n19725), .A2(n20620), .A3(n20617), .ZN(n19731) );
  NOR4_X1 U22830 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_21__SCAN_IN), .A3(P2_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_23__SCAN_IN), .ZN(n19729) );
  NOR4_X1 U22831 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_17__SCAN_IN), .A3(P2_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_19__SCAN_IN), .ZN(n19728) );
  NOR4_X1 U22832 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_29__SCAN_IN), .A3(P2_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_31__SCAN_IN), .ZN(n19727) );
  NOR4_X1 U22833 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_25__SCAN_IN), .A3(P2_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_27__SCAN_IN), .ZN(n19726) );
  NAND4_X1 U22834 ( .A1(n19729), .A2(n19728), .A3(n19727), .A4(n19726), .ZN(
        n19730) );
  NOR4_X1 U22835 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_3__SCAN_IN), .A3(n19731), .A4(n19730), .ZN(n19732) );
  NAND3_X1 U22836 ( .A1(n19734), .A2(n19733), .A3(n19732), .ZN(n19741) );
  NOR2_X1 U22837 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n19741), .ZN(n19735) );
  INV_X1 U22838 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n20690) );
  AOI22_X1 U22839 ( .A1(n19735), .A2(n19736), .B1(n19741), .B2(n20690), .ZN(
        P2_U2820) );
  OR3_X1 U22840 ( .A1(P2_REIP_REG_0__SCAN_IN), .A2(P2_DATAWIDTH_REG_1__SCAN_IN), .A3(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n19740) );
  INV_X1 U22841 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n20688) );
  AOI22_X1 U22842 ( .A1(n19735), .A2(n19740), .B1(n19741), .B2(n20688), .ZN(
        P2_U2821) );
  INV_X1 U22843 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20693) );
  NAND2_X1 U22844 ( .A1(n19735), .A2(n20693), .ZN(n19739) );
  INV_X1 U22845 ( .A(n19741), .ZN(n19742) );
  OAI21_X1 U22846 ( .B1(n19736), .B2(n10371), .A(n19742), .ZN(n19737) );
  OAI21_X1 U22847 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n19742), .A(n19737), 
        .ZN(n19738) );
  OAI221_X1 U22848 ( .B1(n19739), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n19739), .C2(P2_REIP_REG_0__SCAN_IN), .A(n19738), .ZN(P2_U2822) );
  INV_X1 U22849 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n20686) );
  OAI221_X1 U22850 ( .B1(n19742), .B2(n20686), .C1(n19741), .C2(n19740), .A(
        n19739), .ZN(P2_U2823) );
  OAI22_X1 U22851 ( .A1(n10085), .A2(n19815), .B1(n20663), .B2(n19887), .ZN(
        n19744) );
  NOR2_X1 U22852 ( .A1(n19888), .A2(n10990), .ZN(n19743) );
  AOI211_X1 U22853 ( .C1(n19745), .C2(n19922), .A(n19744), .B(n19743), .ZN(
        n19746) );
  OAI21_X1 U22854 ( .B1(n19747), .B2(n19919), .A(n19746), .ZN(n19748) );
  INV_X1 U22855 ( .A(n19748), .ZN(n19753) );
  OAI211_X1 U22856 ( .C1(n19751), .C2(n19750), .A(n19897), .B(n19749), .ZN(
        n19752) );
  OAI211_X1 U22857 ( .C1(n19914), .C2(n19754), .A(n19753), .B(n19752), .ZN(
        P2_U2834) );
  INV_X1 U22858 ( .A(n19755), .ZN(n19756) );
  AOI21_X1 U22859 ( .B1(n19760), .B2(n19756), .A(n19932), .ZN(n19759) );
  AOI22_X1 U22860 ( .A1(n19759), .A2(n19758), .B1(n19877), .B2(n19757), .ZN(
        n19767) );
  AOI22_X1 U22861 ( .A1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n19929), .B1(
        P2_REIP_REG_20__SCAN_IN), .B2(n19927), .ZN(n19766) );
  AOI22_X1 U22862 ( .A1(P2_EBX_REG_20__SCAN_IN), .A2(n19917), .B1(n19760), 
        .B2(n19928), .ZN(n19765) );
  OAI22_X1 U22863 ( .A1(n19762), .A2(n19880), .B1(n19761), .B2(n19914), .ZN(
        n19763) );
  INV_X1 U22864 ( .A(n19763), .ZN(n19764) );
  NAND4_X1 U22865 ( .A1(n19767), .A2(n19766), .A3(n19765), .A4(n19764), .ZN(
        P2_U2835) );
  OAI21_X1 U22866 ( .B1(n20660), .B2(n19887), .A(n20073), .ZN(n19771) );
  OAI22_X1 U22867 ( .A1(n19769), .A2(n19919), .B1(n19768), .B2(n19815), .ZN(
        n19770) );
  AOI211_X1 U22868 ( .C1(P2_EBX_REG_19__SCAN_IN), .C2(n19917), .A(n19771), .B(
        n19770), .ZN(n19778) );
  NAND2_X1 U22869 ( .A1(n9718), .A2(n19772), .ZN(n19774) );
  XNOR2_X1 U22870 ( .A(n19774), .B(n19773), .ZN(n19776) );
  AOI22_X1 U22871 ( .A1(n19776), .A2(n19897), .B1(n19775), .B2(n19922), .ZN(
        n19777) );
  OAI211_X1 U22872 ( .C1(n19779), .C2(n19914), .A(n19778), .B(n19777), .ZN(
        P2_U2836) );
  NOR2_X1 U22873 ( .A1(n9766), .A2(n19792), .ZN(n19781) );
  XOR2_X1 U22874 ( .A(n19781), .B(n19780), .Z(n19791) );
  OAI21_X1 U22875 ( .B1(n20658), .B2(n19887), .A(n20073), .ZN(n19785) );
  INV_X1 U22876 ( .A(n19782), .ZN(n19783) );
  OAI22_X1 U22877 ( .A1(n19783), .A2(n19919), .B1(n19888), .B2(n10748), .ZN(
        n19784) );
  AOI211_X1 U22878 ( .C1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(n19929), .A(
        n19785), .B(n19784), .ZN(n19790) );
  OAI22_X1 U22879 ( .A1(n19787), .A2(n19880), .B1(n19786), .B2(n19914), .ZN(
        n19788) );
  INV_X1 U22880 ( .A(n19788), .ZN(n19789) );
  OAI211_X1 U22881 ( .C1(n20613), .C2(n19791), .A(n19790), .B(n19789), .ZN(
        P2_U2837) );
  AOI211_X1 U22882 ( .C1(n19798), .C2(n19793), .A(n19792), .B(n19932), .ZN(
        n19797) );
  AOI22_X1 U22883 ( .A1(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n19929), .B1(
        P2_REIP_REG_17__SCAN_IN), .B2(n19927), .ZN(n19794) );
  OAI211_X1 U22884 ( .C1(n19795), .C2(n19919), .A(n19794), .B(n20073), .ZN(
        n19796) );
  AOI211_X1 U22885 ( .C1(P2_EBX_REG_17__SCAN_IN), .C2(n19917), .A(n19797), .B(
        n19796), .ZN(n19801) );
  AOI22_X1 U22886 ( .A1(n19799), .A2(n19922), .B1(n19928), .B2(n19798), .ZN(
        n19800) );
  OAI211_X1 U22887 ( .C1(n19802), .C2(n19914), .A(n19801), .B(n19800), .ZN(
        P2_U2838) );
  NOR2_X1 U22888 ( .A1(n9766), .A2(n19803), .ZN(n19805) );
  XOR2_X1 U22889 ( .A(n19805), .B(n19804), .Z(n19814) );
  OAI21_X1 U22890 ( .B1(n20654), .B2(n19887), .A(n20073), .ZN(n19808) );
  OAI22_X1 U22891 ( .A1(n19806), .A2(n19919), .B1(n19888), .B2(n14256), .ZN(
        n19807) );
  AOI211_X1 U22892 ( .C1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .C2(n19929), .A(
        n19808), .B(n19807), .ZN(n19813) );
  OAI22_X1 U22893 ( .A1(n19810), .A2(n19880), .B1(n19809), .B2(n19914), .ZN(
        n19811) );
  INV_X1 U22894 ( .A(n19811), .ZN(n19812) );
  OAI211_X1 U22895 ( .C1(n20613), .C2(n19814), .A(n19813), .B(n19812), .ZN(
        P2_U2839) );
  OAI21_X1 U22896 ( .B1(n10972), .B2(n19887), .A(n20073), .ZN(n19819) );
  OAI22_X1 U22897 ( .A1(n19817), .A2(n19919), .B1(n19816), .B2(n19815), .ZN(
        n19818) );
  AOI211_X1 U22898 ( .C1(P2_EBX_REG_15__SCAN_IN), .C2(n19917), .A(n19819), .B(
        n19818), .ZN(n19826) );
  NAND2_X1 U22899 ( .A1(n9718), .A2(n19820), .ZN(n19821) );
  XNOR2_X1 U22900 ( .A(n19822), .B(n19821), .ZN(n19824) );
  AOI22_X1 U22901 ( .A1(n19824), .A2(n19897), .B1(n19823), .B2(n19922), .ZN(
        n19825) );
  OAI211_X1 U22902 ( .C1(n19827), .C2(n19914), .A(n19826), .B(n19825), .ZN(
        P2_U2840) );
  NOR2_X1 U22903 ( .A1(n9766), .A2(n19828), .ZN(n19830) );
  XOR2_X1 U22904 ( .A(n19830), .B(n19829), .Z(n19838) );
  OAI21_X1 U22905 ( .B1(n10967), .B2(n19887), .A(n20073), .ZN(n19833) );
  OAI22_X1 U22906 ( .A1(n19831), .A2(n19919), .B1(n19888), .B2(n10757), .ZN(
        n19832) );
  AOI211_X1 U22907 ( .C1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .C2(n19929), .A(
        n19833), .B(n19832), .ZN(n19837) );
  AOI22_X1 U22908 ( .A1(n19835), .A2(n19922), .B1(n19834), .B2(n19915), .ZN(
        n19836) );
  OAI211_X1 U22909 ( .C1(n20613), .C2(n19838), .A(n19837), .B(n19836), .ZN(
        P2_U2841) );
  AOI22_X1 U22910 ( .A1(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n19929), .B1(
        P2_EBX_REG_13__SCAN_IN), .B2(n19917), .ZN(n19839) );
  OAI21_X1 U22911 ( .B1(n19840), .B2(n19919), .A(n19839), .ZN(n19841) );
  AOI211_X1 U22912 ( .C1(P2_REIP_REG_13__SCAN_IN), .C2(n19927), .A(n19905), 
        .B(n19841), .ZN(n19848) );
  NAND2_X1 U22913 ( .A1(n9718), .A2(n19842), .ZN(n19843) );
  XNOR2_X1 U22914 ( .A(n19844), .B(n19843), .ZN(n19846) );
  AOI22_X1 U22915 ( .A1(n19846), .A2(n19910), .B1(n19845), .B2(n19922), .ZN(
        n19847) );
  OAI211_X1 U22916 ( .C1(n19849), .C2(n19914), .A(n19848), .B(n19847), .ZN(
        P2_U2842) );
  NOR2_X1 U22917 ( .A1(n9766), .A2(n19850), .ZN(n19851) );
  XOR2_X1 U22918 ( .A(n19852), .B(n19851), .Z(n19862) );
  INV_X1 U22919 ( .A(n19853), .ZN(n19854) );
  AOI22_X1 U22920 ( .A1(n19854), .A2(n19877), .B1(
        P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n19929), .ZN(n19855) );
  OAI211_X1 U22921 ( .C1(n10962), .C2(n19887), .A(n19855), .B(n20073), .ZN(
        n19860) );
  INV_X1 U22922 ( .A(n19856), .ZN(n19858) );
  OAI22_X1 U22923 ( .A1(n19858), .A2(n19880), .B1(n19857), .B2(n19914), .ZN(
        n19859) );
  AOI211_X1 U22924 ( .C1(P2_EBX_REG_12__SCAN_IN), .C2(n19917), .A(n19860), .B(
        n19859), .ZN(n19861) );
  OAI21_X1 U22925 ( .B1(n20613), .B2(n19862), .A(n19861), .ZN(P2_U2843) );
  INV_X1 U22926 ( .A(n19863), .ZN(n19865) );
  AOI22_X1 U22927 ( .A1(P2_EBX_REG_11__SCAN_IN), .A2(n19917), .B1(
        P2_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n19929), .ZN(n19864) );
  OAI21_X1 U22928 ( .B1(n19865), .B2(n19919), .A(n19864), .ZN(n19866) );
  AOI211_X1 U22929 ( .C1(P2_REIP_REG_11__SCAN_IN), .C2(n19927), .A(n20028), 
        .B(n19866), .ZN(n19872) );
  NAND2_X1 U22930 ( .A1(n9718), .A2(n19867), .ZN(n19868) );
  XNOR2_X1 U22931 ( .A(n19869), .B(n19868), .ZN(n19870) );
  AOI22_X1 U22932 ( .A1(n19870), .A2(n19897), .B1(n19954), .B2(n19922), .ZN(
        n19871) );
  OAI211_X1 U22933 ( .C1(n19873), .C2(n19914), .A(n19872), .B(n19871), .ZN(
        P2_U2844) );
  NAND2_X1 U22934 ( .A1(n9719), .A2(n19874), .ZN(n19876) );
  XOR2_X1 U22935 ( .A(n19876), .B(n19875), .Z(n19886) );
  AOI22_X1 U22936 ( .A1(n19878), .A2(n19877), .B1(P2_EBX_REG_7__SCAN_IN), .B2(
        n19917), .ZN(n19879) );
  OAI211_X1 U22937 ( .C1(n10940), .C2(n19887), .A(n19879), .B(n20073), .ZN(
        n19884) );
  OAI22_X1 U22938 ( .A1(n19882), .A2(n19914), .B1(n19881), .B2(n19880), .ZN(
        n19883) );
  AOI211_X1 U22939 ( .C1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .C2(n19929), .A(
        n19884), .B(n19883), .ZN(n19885) );
  OAI21_X1 U22940 ( .B1(n19886), .B2(n20613), .A(n19885), .ZN(P2_U2848) );
  OAI21_X1 U22941 ( .B1(n14389), .B2(n19887), .A(n20073), .ZN(n19891) );
  OAI22_X1 U22942 ( .A1(n19889), .A2(n19919), .B1(n19888), .B2(n10932), .ZN(
        n19890) );
  AOI211_X1 U22943 ( .C1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .C2(n19929), .A(
        n19891), .B(n19890), .ZN(n19900) );
  NOR2_X1 U22944 ( .A1(n9766), .A2(n19892), .ZN(n19894) );
  XNOR2_X1 U22945 ( .A(n19894), .B(n19893), .ZN(n19898) );
  INV_X1 U22946 ( .A(n19895), .ZN(n19896) );
  AOI22_X1 U22947 ( .A1(n19898), .A2(n19897), .B1(n19896), .B2(n19922), .ZN(
        n19899) );
  OAI211_X1 U22948 ( .C1(n19914), .C2(n19901), .A(n19900), .B(n19899), .ZN(
        P2_U2849) );
  AOI22_X1 U22949 ( .A1(P2_EBX_REG_5__SCAN_IN), .A2(n19917), .B1(
        P2_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n19929), .ZN(n19902) );
  OAI21_X1 U22950 ( .B1(n19903), .B2(n19919), .A(n19902), .ZN(n19904) );
  AOI211_X1 U22951 ( .C1(P2_REIP_REG_5__SCAN_IN), .C2(n19927), .A(n19905), .B(
        n19904), .ZN(n19913) );
  NAND2_X1 U22952 ( .A1(n9719), .A2(n19906), .ZN(n19907) );
  XNOR2_X1 U22953 ( .A(n19908), .B(n19907), .ZN(n19911) );
  AOI22_X1 U22954 ( .A1(n19911), .A2(n19910), .B1(n19909), .B2(n19922), .ZN(
        n19912) );
  OAI211_X1 U22955 ( .C1(n19914), .C2(n19987), .A(n19913), .B(n19912), .ZN(
        P2_U2850) );
  AOI22_X1 U22956 ( .A1(n19917), .A2(P2_EBX_REG_0__SCAN_IN), .B1(n19916), .B2(
        n19915), .ZN(n19918) );
  OAI21_X1 U22957 ( .B1(n19920), .B2(n19919), .A(n19918), .ZN(n19921) );
  AOI21_X1 U22958 ( .B1(n19923), .B2(n19922), .A(n19921), .ZN(n19924) );
  OAI21_X1 U22959 ( .B1(n20727), .B2(n19925), .A(n19924), .ZN(n19926) );
  AOI21_X1 U22960 ( .B1(n19927), .B2(P2_REIP_REG_0__SCAN_IN), .A(n19926), .ZN(
        n19931) );
  OAI21_X1 U22961 ( .B1(n19929), .B2(n19928), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n19930) );
  OAI211_X1 U22962 ( .C1(n19933), .C2(n19932), .A(n19931), .B(n19930), .ZN(
        P2_U2855) );
  OR2_X1 U22963 ( .A1(n19944), .A2(n19934), .ZN(n19936) );
  AOI211_X1 U22964 ( .C1(n19937), .C2(n19936), .A(n19959), .B(n19935), .ZN(
        n19938) );
  AOI21_X1 U22965 ( .B1(P2_EBX_REG_15__SCAN_IN), .B2(n19947), .A(n19938), .ZN(
        n19939) );
  OAI21_X1 U22966 ( .B1(n19940), .B2(n19947), .A(n19939), .ZN(P2_U2872) );
  OR2_X1 U22967 ( .A1(n19953), .A2(n19941), .ZN(n19943) );
  AOI21_X1 U22968 ( .B1(n19943), .B2(n19942), .A(n19959), .ZN(n19945) );
  AOI22_X1 U22969 ( .A1(n19945), .A2(n19944), .B1(P2_EBX_REG_13__SCAN_IN), 
        .B2(n19947), .ZN(n19946) );
  OAI21_X1 U22970 ( .B1(n19948), .B2(n19947), .A(n19946), .ZN(P2_U2874) );
  INV_X1 U22971 ( .A(n19949), .ZN(n19950) );
  NOR2_X1 U22972 ( .A1(n19950), .A2(n19959), .ZN(n19956) );
  OAI21_X1 U22973 ( .B1(n19953), .B2(n19952), .A(n19951), .ZN(n19955) );
  AOI22_X1 U22974 ( .A1(n19956), .A2(n19955), .B1(n19969), .B2(n19954), .ZN(
        n19957) );
  OAI21_X1 U22975 ( .B1(n19969), .B2(n19958), .A(n19957), .ZN(P2_U2876) );
  NOR2_X1 U22976 ( .A1(n19960), .A2(n19959), .ZN(n19967) );
  OAI21_X1 U22977 ( .B1(n19963), .B2(n19962), .A(n19961), .ZN(n19966) );
  AOI22_X1 U22978 ( .A1(n19967), .A2(n19966), .B1(n19965), .B2(n19964), .ZN(
        n19968) );
  OAI21_X1 U22979 ( .B1(n19969), .B2(n9947), .A(n19968), .ZN(P2_U2878) );
  OAI22_X1 U22980 ( .A1(n19980), .A2(n19970), .B1(n19979), .B2(n19993), .ZN(
        n19971) );
  INV_X1 U22981 ( .A(n19971), .ZN(n19972) );
  OAI21_X1 U22982 ( .B1(n19988), .B2(n19973), .A(n19972), .ZN(P2_U2905) );
  INV_X1 U22983 ( .A(n19980), .ZN(n19976) );
  AOI22_X1 U22984 ( .A1(n19976), .A2(n19975), .B1(P2_EAX_REG_8__SCAN_IN), .B2(
        n19974), .ZN(n19977) );
  OAI21_X1 U22985 ( .B1(n19988), .B2(n19978), .A(n19977), .ZN(P2_U2911) );
  INV_X1 U22986 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n20012) );
  OAI22_X1 U22987 ( .A1(n19980), .A2(n20108), .B1(n19979), .B2(n20012), .ZN(
        n19981) );
  INV_X1 U22988 ( .A(n19981), .ZN(n19986) );
  OR3_X1 U22989 ( .A1(n19984), .A2(n19983), .A3(n19982), .ZN(n19985) );
  OAI211_X1 U22990 ( .C1(n19988), .C2(n19987), .A(n19986), .B(n19985), .ZN(
        P2_U2914) );
  NOR2_X1 U22991 ( .A1(n20020), .A2(n19989), .ZN(P2_U2920) );
  AOI22_X1 U22992 ( .A1(n20025), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n20024), 
        .B2(P2_DATAO_REG_15__SCAN_IN), .ZN(n19990) );
  OAI21_X1 U22993 ( .B1(n19991), .B2(n20027), .A(n19990), .ZN(P2_U2936) );
  AOI22_X1 U22994 ( .A1(n20025), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n20024), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n19992) );
  OAI21_X1 U22995 ( .B1(n19993), .B2(n20027), .A(n19992), .ZN(P2_U2937) );
  AOI22_X1 U22996 ( .A1(n20021), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n20024), 
        .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n19994) );
  OAI21_X1 U22997 ( .B1(n19995), .B2(n20027), .A(n19994), .ZN(P2_U2938) );
  AOI22_X1 U22998 ( .A1(n20021), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(n20024), 
        .B2(P2_DATAO_REG_12__SCAN_IN), .ZN(n19996) );
  OAI21_X1 U22999 ( .B1(n19997), .B2(n20027), .A(n19996), .ZN(P2_U2939) );
  AOI22_X1 U23000 ( .A1(n20021), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n20024), 
        .B2(P2_DATAO_REG_11__SCAN_IN), .ZN(n19998) );
  OAI21_X1 U23001 ( .B1(n19999), .B2(n20027), .A(n19998), .ZN(P2_U2940) );
  AOI22_X1 U23002 ( .A1(n20021), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n20024), 
        .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n20000) );
  OAI21_X1 U23003 ( .B1(n20001), .B2(n20027), .A(n20000), .ZN(P2_U2941) );
  AOI22_X1 U23004 ( .A1(n20021), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n20024), 
        .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n20002) );
  OAI21_X1 U23005 ( .B1(n20003), .B2(n20027), .A(n20002), .ZN(P2_U2942) );
  AOI22_X1 U23006 ( .A1(n20021), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n20024), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n20004) );
  OAI21_X1 U23007 ( .B1(n20005), .B2(n20027), .A(n20004), .ZN(P2_U2943) );
  OAI222_X1 U23008 ( .A1(n20743), .A2(n20008), .B1(n20027), .B2(n20007), .C1(
        n20020), .C2(n20006), .ZN(P2_U2944) );
  AOI22_X1 U23009 ( .A1(n20021), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n20024), 
        .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n20009) );
  OAI21_X1 U23010 ( .B1(n20010), .B2(n20027), .A(n20009), .ZN(P2_U2945) );
  AOI22_X1 U23011 ( .A1(n20021), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n20024), 
        .B2(P2_DATAO_REG_5__SCAN_IN), .ZN(n20011) );
  OAI21_X1 U23012 ( .B1(n20012), .B2(n20027), .A(n20011), .ZN(P2_U2946) );
  INV_X1 U23013 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n20014) );
  AOI22_X1 U23014 ( .A1(n20021), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n20024), 
        .B2(P2_DATAO_REG_4__SCAN_IN), .ZN(n20013) );
  OAI21_X1 U23015 ( .B1(n20014), .B2(n20027), .A(n20013), .ZN(P2_U2947) );
  INV_X1 U23016 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n20016) );
  AOI22_X1 U23017 ( .A1(n20021), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n20024), 
        .B2(P2_DATAO_REG_3__SCAN_IN), .ZN(n20015) );
  OAI21_X1 U23018 ( .B1(n20016), .B2(n20027), .A(n20015), .ZN(P2_U2948) );
  INV_X1 U23019 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n20018) );
  INV_X1 U23020 ( .A(P2_LWORD_REG_2__SCAN_IN), .ZN(n20017) );
  OAI222_X1 U23021 ( .A1(n20020), .A2(n20019), .B1(n20027), .B2(n20018), .C1(
        n20743), .C2(n20017), .ZN(P2_U2949) );
  INV_X1 U23022 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n20023) );
  AOI22_X1 U23023 ( .A1(n20021), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n20024), 
        .B2(P2_DATAO_REG_1__SCAN_IN), .ZN(n20022) );
  OAI21_X1 U23024 ( .B1(n20023), .B2(n20027), .A(n20022), .ZN(P2_U2950) );
  AOI22_X1 U23025 ( .A1(n20025), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n20024), 
        .B2(P2_DATAO_REG_0__SCAN_IN), .ZN(n20026) );
  OAI21_X1 U23026 ( .B1(n11744), .B2(n20027), .A(n20026), .ZN(P2_U2951) );
  AOI22_X1 U23027 ( .A1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n20029), .B1(
        P2_REIP_REG_4__SCAN_IN), .B2(n20028), .ZN(n20040) );
  INV_X1 U23028 ( .A(n20030), .ZN(n20031) );
  XNOR2_X1 U23029 ( .A(n20032), .B(n20031), .ZN(n20060) );
  INV_X1 U23030 ( .A(n20060), .ZN(n20036) );
  XNOR2_X1 U23031 ( .A(n20033), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n20035) );
  XNOR2_X1 U23032 ( .A(n20035), .B(n20034), .ZN(n20069) );
  OAI22_X1 U23033 ( .A1(n20036), .A2(n16974), .B1(n20043), .B2(n20069), .ZN(
        n20037) );
  AOI21_X1 U23034 ( .B1(n20051), .B2(n20038), .A(n20037), .ZN(n20039) );
  OAI211_X1 U23035 ( .C1(n20045), .C2(n20041), .A(n20040), .B(n20039), .ZN(
        P2_U3010) );
  INV_X1 U23036 ( .A(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n20054) );
  OAI22_X1 U23037 ( .A1(n20045), .A2(n20044), .B1(n20043), .B2(n20042), .ZN(
        n20050) );
  AND3_X1 U23038 ( .A1(n20048), .A2(n20047), .A3(n20046), .ZN(n20049) );
  AOI211_X1 U23039 ( .C1(n20051), .C2(n10430), .A(n20050), .B(n20049), .ZN(
        n20053) );
  OAI211_X1 U23040 ( .C1(n20055), .C2(n20054), .A(n20053), .B(n20052), .ZN(
        P2_U3012) );
  AOI22_X1 U23041 ( .A1(n20058), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B1(
        n20057), .B2(n20056), .ZN(n20072) );
  NAND2_X1 U23042 ( .A1(n20060), .A2(n20059), .ZN(n20067) );
  NOR2_X1 U23043 ( .A1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n20061), .ZN(
        n20065) );
  NOR2_X1 U23044 ( .A1(n20063), .A2(n20062), .ZN(n20064) );
  NOR2_X1 U23045 ( .A1(n20065), .A2(n20064), .ZN(n20066) );
  OAI211_X1 U23046 ( .C1(n20069), .C2(n20068), .A(n20067), .B(n20066), .ZN(
        n20070) );
  INV_X1 U23047 ( .A(n20070), .ZN(n20071) );
  OAI211_X1 U23048 ( .C1(n10921), .C2(n20073), .A(n20072), .B(n20071), .ZN(
        P2_U3042) );
  NAND2_X1 U23049 ( .A1(n10567), .A2(n20710), .ZN(n20188) );
  OR2_X1 U23050 ( .A1(n20188), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n20134) );
  NOR2_X1 U23051 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20134), .ZN(
        n20122) );
  AOI22_X1 U23052 ( .A1(n20579), .A2(n20557), .B1(n20548), .B2(n20122), .ZN(
        n20086) );
  AOI21_X1 U23053 ( .B1(n20605), .B2(n20156), .A(n11033), .ZN(n20076) );
  NOR2_X1 U23054 ( .A1(n20076), .A2(n20509), .ZN(n20081) );
  INV_X1 U23055 ( .A(n20077), .ZN(n20082) );
  AOI21_X1 U23056 ( .B1(n20082), .B2(n20333), .A(n20699), .ZN(n20078) );
  AOI21_X1 U23057 ( .B1(n20081), .B2(n20080), .A(n20078), .ZN(n20079) );
  INV_X1 U23058 ( .A(n20080), .ZN(n20597) );
  OAI21_X1 U23059 ( .B1(n20597), .B2(n20122), .A(n20081), .ZN(n20084) );
  OAI21_X1 U23060 ( .B1(n20082), .B2(n20122), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20083) );
  NAND2_X1 U23061 ( .A1(n20084), .A2(n20083), .ZN(n20124) );
  AOI22_X1 U23062 ( .A1(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n20125), .B1(
        n13591), .B2(n20124), .ZN(n20085) );
  OAI211_X1 U23063 ( .C1(n20560), .C2(n20156), .A(n20086), .B(n20085), .ZN(
        P2_U3048) );
  AOI22_X1 U23064 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n20119), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n20118), .ZN(n20428) );
  AOI22_X1 U23065 ( .A1(n20561), .A2(n20579), .B1(n20087), .B2(n20122), .ZN(
        n20091) );
  AOI22_X1 U23066 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n20125), .B1(
        n20089), .B2(n20124), .ZN(n20090) );
  OAI211_X1 U23067 ( .C1(n20564), .C2(n20156), .A(n20091), .B(n20090), .ZN(
        P2_U3049) );
  AOI22_X1 U23068 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n20119), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n20118), .ZN(n20527) );
  AOI22_X1 U23069 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n20119), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n20118), .ZN(n20569) );
  NOR2_X2 U23070 ( .A1(n10325), .A2(n20120), .ZN(n20565) );
  AOI22_X1 U23071 ( .A1(n20524), .A2(n20579), .B1(n20565), .B2(n20122), .ZN(
        n20095) );
  AOI22_X1 U23072 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n20125), .B1(
        n20093), .B2(n20124), .ZN(n20094) );
  OAI211_X1 U23073 ( .C1(n20527), .C2(n20156), .A(n20095), .B(n20094), .ZN(
        P2_U3050) );
  INV_X1 U23074 ( .A(n20119), .ZN(n20111) );
  INV_X1 U23075 ( .A(n20118), .ZN(n20113) );
  OAI22_X1 U23076 ( .A1(n20097), .A2(n20111), .B1(n20096), .B2(n20113), .ZN(
        n20455) );
  AOI22_X1 U23077 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n20118), .B1(
        BUF1_REG_27__SCAN_IN), .B2(n20119), .ZN(n20433) );
  NOR2_X2 U23078 ( .A1(n20098), .A2(n20120), .ZN(n20570) );
  AOI22_X1 U23079 ( .A1(n20572), .A2(n20579), .B1(n20570), .B2(n20122), .ZN(
        n20101) );
  NOR2_X2 U23080 ( .A1(n20099), .A2(n20551), .ZN(n20571) );
  AOI22_X1 U23081 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n20125), .B1(
        n20571), .B2(n20124), .ZN(n20100) );
  OAI211_X1 U23082 ( .C1(n20575), .C2(n20156), .A(n20101), .B(n20100), .ZN(
        P2_U3051) );
  AOI22_X1 U23083 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n20119), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n20118), .ZN(n20495) );
  AOI22_X1 U23084 ( .A1(n20492), .A2(n20579), .B1(n20576), .B2(n20122), .ZN(
        n20107) );
  NOR2_X2 U23085 ( .A1(n20105), .A2(n20551), .ZN(n20577) );
  AOI22_X1 U23086 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n20125), .B1(
        n20577), .B2(n20124), .ZN(n20106) );
  OAI211_X1 U23087 ( .C1(n20495), .C2(n20156), .A(n20107), .B(n20106), .ZN(
        P2_U3052) );
  AOI22_X1 U23088 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n20119), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n20118), .ZN(n20589) );
  AOI22_X1 U23089 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n20118), .B1(
        BUF1_REG_29__SCAN_IN), .B2(n20119), .ZN(n20438) );
  NOR2_X2 U23090 ( .A1(n10838), .A2(n20120), .ZN(n20584) );
  AOI22_X1 U23091 ( .A1(n20586), .A2(n20579), .B1(n20584), .B2(n20122), .ZN(
        n20110) );
  NOR2_X2 U23092 ( .A1(n20108), .A2(n20551), .ZN(n20585) );
  AOI22_X1 U23093 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n20125), .B1(
        n20585), .B2(n20124), .ZN(n20109) );
  OAI211_X1 U23094 ( .C1(n20589), .C2(n20156), .A(n20110), .B(n20109), .ZN(
        P2_U3053) );
  AOI22_X1 U23095 ( .A1(BUF2_REG_22__SCAN_IN), .A2(n20118), .B1(
        BUF1_REG_22__SCAN_IN), .B2(n20119), .ZN(n20595) );
  OAI22_X1 U23096 ( .A1(n20114), .A2(n20113), .B1(n20112), .B2(n20111), .ZN(
        n20592) );
  AOI22_X1 U23097 ( .A1(n20592), .A2(n20579), .B1(n21297), .B2(n20122), .ZN(
        n20117) );
  NOR2_X2 U23098 ( .A1(n20115), .A2(n20551), .ZN(n20591) );
  AOI22_X1 U23099 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n20125), .B1(
        n20591), .B2(n20124), .ZN(n20116) );
  OAI211_X1 U23100 ( .C1(n20595), .C2(n20156), .A(n20117), .B(n20116), .ZN(
        P2_U3054) );
  AOI22_X1 U23101 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n20119), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n20118), .ZN(n20606) );
  AOI22_X1 U23102 ( .A1(BUF1_REG_31__SCAN_IN), .A2(n20119), .B1(
        BUF2_REG_31__SCAN_IN), .B2(n20118), .ZN(n20396) );
  AOI22_X1 U23103 ( .A1(n20600), .A2(n20579), .B1(n20596), .B2(n20122), .ZN(
        n20127) );
  NOR2_X2 U23104 ( .A1(n20123), .A2(n20551), .ZN(n20598) );
  AOI22_X1 U23105 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n20125), .B1(
        n20598), .B2(n20124), .ZN(n20126) );
  OAI211_X1 U23106 ( .C1(n20606), .C2(n20156), .A(n20127), .B(n20126), .ZN(
        P2_U3055) );
  INV_X1 U23107 ( .A(n20128), .ZN(n20306) );
  INV_X1 U23108 ( .A(n20129), .ZN(n20130) );
  NOR2_X1 U23109 ( .A1(n20364), .A2(n20188), .ZN(n20151) );
  NOR3_X1 U23110 ( .A1(n20130), .A2(n20151), .A3(n20607), .ZN(n20133) );
  AOI211_X2 U23111 ( .C1(n20134), .C2(n20607), .A(n20306), .B(n20133), .ZN(
        n20152) );
  AOI22_X1 U23112 ( .A1(n20152), .A2(n13591), .B1(n20548), .B2(n20151), .ZN(
        n20138) );
  NAND2_X1 U23113 ( .A1(n20131), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n20297) );
  INV_X1 U23114 ( .A(n20297), .ZN(n20132) );
  NAND2_X1 U23115 ( .A1(n20132), .A2(n20365), .ZN(n20135) );
  AOI21_X1 U23116 ( .B1(n20135), .B2(n20134), .A(n20133), .ZN(n20136) );
  OAI211_X1 U23117 ( .C1(n20151), .C2(n20333), .A(n20136), .B(n20512), .ZN(
        n20153) );
  AOI22_X1 U23118 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n20153), .B1(
        n20182), .B2(n20506), .ZN(n20137) );
  OAI211_X1 U23119 ( .C1(n20521), .C2(n20156), .A(n20138), .B(n20137), .ZN(
        P2_U3056) );
  AOI22_X1 U23120 ( .A1(n20152), .A2(n20089), .B1(n20087), .B2(n20151), .ZN(
        n20140) );
  INV_X1 U23121 ( .A(n20564), .ZN(n20450) );
  AOI22_X1 U23122 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n20153), .B1(
        n20182), .B2(n20450), .ZN(n20139) );
  OAI211_X1 U23123 ( .C1(n20428), .C2(n20156), .A(n20140), .B(n20139), .ZN(
        P2_U3057) );
  AOI22_X1 U23124 ( .A1(n20152), .A2(n20093), .B1(n20565), .B2(n20151), .ZN(
        n20142) );
  INV_X1 U23125 ( .A(n20527), .ZN(n20566) );
  AOI22_X1 U23126 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n20153), .B1(
        n20182), .B2(n20566), .ZN(n20141) );
  OAI211_X1 U23127 ( .C1(n20569), .C2(n20156), .A(n20142), .B(n20141), .ZN(
        P2_U3058) );
  AOI22_X1 U23128 ( .A1(n20152), .A2(n20571), .B1(n20570), .B2(n20151), .ZN(
        n20144) );
  AOI22_X1 U23129 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n20153), .B1(
        n20182), .B2(n20455), .ZN(n20143) );
  OAI211_X1 U23130 ( .C1(n20433), .C2(n20156), .A(n20144), .B(n20143), .ZN(
        P2_U3059) );
  INV_X1 U23131 ( .A(n20492), .ZN(n20583) );
  AOI22_X1 U23132 ( .A1(n20152), .A2(n20577), .B1(n20576), .B2(n20151), .ZN(
        n20146) );
  INV_X1 U23133 ( .A(n20495), .ZN(n20578) );
  AOI22_X1 U23134 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n20153), .B1(
        n20182), .B2(n20578), .ZN(n20145) );
  OAI211_X1 U23135 ( .C1(n20583), .C2(n20156), .A(n20146), .B(n20145), .ZN(
        P2_U3060) );
  AOI22_X1 U23136 ( .A1(n20152), .A2(n20585), .B1(n20584), .B2(n20151), .ZN(
        n20148) );
  INV_X1 U23137 ( .A(n20589), .ZN(n20460) );
  AOI22_X1 U23138 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n20153), .B1(
        n20182), .B2(n20460), .ZN(n20147) );
  OAI211_X1 U23139 ( .C1(n20438), .C2(n20156), .A(n20148), .B(n20147), .ZN(
        P2_U3061) );
  INV_X1 U23140 ( .A(n20592), .ZN(n20538) );
  AOI22_X1 U23141 ( .A1(n20152), .A2(n20591), .B1(n21297), .B2(n20151), .ZN(
        n20150) );
  INV_X1 U23142 ( .A(n20595), .ZN(n20534) );
  AOI22_X1 U23143 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n20153), .B1(
        n20182), .B2(n20534), .ZN(n20149) );
  OAI211_X1 U23144 ( .C1(n20538), .C2(n20156), .A(n20150), .B(n20149), .ZN(
        P2_U3062) );
  AOI22_X1 U23145 ( .A1(n20152), .A2(n20598), .B1(n20596), .B2(n20151), .ZN(
        n20155) );
  INV_X1 U23146 ( .A(n20606), .ZN(n20468) );
  AOI22_X1 U23147 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n20153), .B1(
        n20182), .B2(n20468), .ZN(n20154) );
  OAI211_X1 U23148 ( .C1(n20396), .C2(n20156), .A(n20155), .B(n20154), .ZN(
        P2_U3063) );
  NOR2_X1 U23149 ( .A1(n20397), .A2(n20188), .ZN(n20180) );
  OAI21_X1 U23150 ( .B1(n20162), .B2(n20180), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20158) );
  NOR2_X1 U23151 ( .A1(n20400), .A2(n20188), .ZN(n20160) );
  INV_X1 U23152 ( .A(n20160), .ZN(n20157) );
  NAND2_X1 U23153 ( .A1(n20158), .A2(n20157), .ZN(n20181) );
  AOI22_X1 U23154 ( .A1(n20181), .A2(n13591), .B1(n20548), .B2(n20180), .ZN(
        n20167) );
  INV_X1 U23155 ( .A(n20182), .ZN(n20159) );
  NAND2_X1 U23156 ( .A1(n20203), .A2(n20159), .ZN(n20161) );
  AOI21_X1 U23157 ( .B1(n20161), .B2(P2_STATEBS16_REG_SCAN_IN), .A(n20160), 
        .ZN(n20164) );
  AOI21_X1 U23158 ( .B1(n20162), .B2(n20333), .A(n20180), .ZN(n20163) );
  MUX2_X1 U23159 ( .A(n20164), .B(n20163), .S(n20509), .Z(n20165) );
  AOI22_X1 U23160 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n20183), .B1(
        n20182), .B2(n20557), .ZN(n20166) );
  OAI211_X1 U23161 ( .C1(n20560), .C2(n20203), .A(n20167), .B(n20166), .ZN(
        P2_U3064) );
  AOI22_X1 U23162 ( .A1(n20181), .A2(n20089), .B1(n20087), .B2(n20180), .ZN(
        n20169) );
  AOI22_X1 U23163 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n20183), .B1(
        n20182), .B2(n20561), .ZN(n20168) );
  OAI211_X1 U23164 ( .C1(n20564), .C2(n20203), .A(n20169), .B(n20168), .ZN(
        P2_U3065) );
  AOI22_X1 U23165 ( .A1(n20181), .A2(n20093), .B1(n20565), .B2(n20180), .ZN(
        n20171) );
  AOI22_X1 U23166 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n20183), .B1(
        n20182), .B2(n20524), .ZN(n20170) );
  OAI211_X1 U23167 ( .C1(n20527), .C2(n20203), .A(n20171), .B(n20170), .ZN(
        P2_U3066) );
  AOI22_X1 U23168 ( .A1(n20181), .A2(n20571), .B1(n20570), .B2(n20180), .ZN(
        n20173) );
  AOI22_X1 U23169 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n20183), .B1(
        n20182), .B2(n20572), .ZN(n20172) );
  OAI211_X1 U23170 ( .C1(n20575), .C2(n20203), .A(n20173), .B(n20172), .ZN(
        P2_U3067) );
  AOI22_X1 U23171 ( .A1(n20181), .A2(n20577), .B1(n20576), .B2(n20180), .ZN(
        n20175) );
  AOI22_X1 U23172 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n20183), .B1(
        n20182), .B2(n20492), .ZN(n20174) );
  OAI211_X1 U23173 ( .C1(n20495), .C2(n20203), .A(n20175), .B(n20174), .ZN(
        P2_U3068) );
  AOI22_X1 U23174 ( .A1(n20181), .A2(n20585), .B1(n20584), .B2(n20180), .ZN(
        n20177) );
  AOI22_X1 U23175 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n20183), .B1(
        n20182), .B2(n20586), .ZN(n20176) );
  OAI211_X1 U23176 ( .C1(n20589), .C2(n20203), .A(n20177), .B(n20176), .ZN(
        P2_U3069) );
  AOI22_X1 U23177 ( .A1(n20181), .A2(n20591), .B1(n21297), .B2(n20180), .ZN(
        n20179) );
  AOI22_X1 U23178 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n20183), .B1(
        n20182), .B2(n20592), .ZN(n20178) );
  OAI211_X1 U23179 ( .C1(n20595), .C2(n20203), .A(n20179), .B(n20178), .ZN(
        P2_U3070) );
  AOI22_X1 U23180 ( .A1(n20181), .A2(n20598), .B1(n20596), .B2(n20180), .ZN(
        n20185) );
  AOI22_X1 U23181 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n20183), .B1(
        n20182), .B2(n20600), .ZN(n20184) );
  OAI211_X1 U23182 ( .C1(n20606), .C2(n20203), .A(n20185), .B(n20184), .ZN(
        P2_U3071) );
  NOR2_X1 U23183 ( .A1(n20186), .A2(n20188), .ZN(n20212) );
  AOI22_X1 U23184 ( .A1(n20213), .A2(n20557), .B1(n20548), .B2(n20212), .ZN(
        n20198) );
  OAI21_X1 U23185 ( .B1(n20297), .B2(n20187), .A(n20699), .ZN(n20196) );
  NOR2_X1 U23186 ( .A1(n20721), .A2(n20188), .ZN(n20193) );
  OAI21_X1 U23187 ( .B1(n20189), .B2(n20607), .A(n20333), .ZN(n20191) );
  INV_X1 U23188 ( .A(n20212), .ZN(n20190) );
  AOI21_X1 U23189 ( .B1(n20191), .B2(n20190), .A(n20551), .ZN(n20192) );
  OAI21_X1 U23190 ( .B1(n20196), .B2(n20193), .A(n20192), .ZN(n20215) );
  INV_X1 U23191 ( .A(n20193), .ZN(n20195) );
  OAI21_X1 U23192 ( .B1(n20189), .B2(n20212), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20194) );
  OAI21_X1 U23193 ( .B1(n20196), .B2(n20195), .A(n20194), .ZN(n20214) );
  AOI22_X1 U23194 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n20215), .B1(
        n13591), .B2(n20214), .ZN(n20197) );
  OAI211_X1 U23195 ( .C1(n20560), .C2(n20223), .A(n20198), .B(n20197), .ZN(
        P2_U3072) );
  AOI22_X1 U23196 ( .A1(n20561), .A2(n20213), .B1(n20212), .B2(n20087), .ZN(
        n20200) );
  AOI22_X1 U23197 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n20215), .B1(
        n20089), .B2(n20214), .ZN(n20199) );
  OAI211_X1 U23198 ( .C1(n20564), .C2(n20223), .A(n20200), .B(n20199), .ZN(
        P2_U3073) );
  AOI22_X1 U23199 ( .A1(n20245), .A2(n20566), .B1(n20212), .B2(n20565), .ZN(
        n20202) );
  AOI22_X1 U23200 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n20215), .B1(
        n20093), .B2(n20214), .ZN(n20201) );
  OAI211_X1 U23201 ( .C1(n20569), .C2(n20203), .A(n20202), .B(n20201), .ZN(
        P2_U3074) );
  AOI22_X1 U23202 ( .A1(n20572), .A2(n20213), .B1(n20212), .B2(n20570), .ZN(
        n20205) );
  AOI22_X1 U23203 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20215), .B1(
        n20571), .B2(n20214), .ZN(n20204) );
  OAI211_X1 U23204 ( .C1(n20575), .C2(n20223), .A(n20205), .B(n20204), .ZN(
        P2_U3075) );
  AOI22_X1 U23205 ( .A1(n20492), .A2(n20213), .B1(n20212), .B2(n20576), .ZN(
        n20207) );
  AOI22_X1 U23206 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n20215), .B1(
        n20577), .B2(n20214), .ZN(n20206) );
  OAI211_X1 U23207 ( .C1(n20495), .C2(n20223), .A(n20207), .B(n20206), .ZN(
        P2_U3076) );
  AOI22_X1 U23208 ( .A1(n20586), .A2(n20213), .B1(n20212), .B2(n20584), .ZN(
        n20209) );
  AOI22_X1 U23209 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n20215), .B1(
        n20585), .B2(n20214), .ZN(n20208) );
  OAI211_X1 U23210 ( .C1(n20589), .C2(n20223), .A(n20209), .B(n20208), .ZN(
        P2_U3077) );
  AOI22_X1 U23211 ( .A1(n20592), .A2(n20213), .B1(n20212), .B2(n21297), .ZN(
        n20211) );
  AOI22_X1 U23212 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20215), .B1(
        n20591), .B2(n20214), .ZN(n20210) );
  OAI211_X1 U23213 ( .C1(n20595), .C2(n20223), .A(n20211), .B(n20210), .ZN(
        P2_U3078) );
  AOI22_X1 U23214 ( .A1(n20600), .A2(n20213), .B1(n20212), .B2(n20596), .ZN(
        n20217) );
  AOI22_X1 U23215 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n20215), .B1(
        n20598), .B2(n20214), .ZN(n20216) );
  OAI211_X1 U23216 ( .C1(n20606), .C2(n20223), .A(n20217), .B(n20216), .ZN(
        P2_U3079) );
  NAND2_X1 U23217 ( .A1(n20219), .A2(n10567), .ZN(n20222) );
  INV_X1 U23218 ( .A(n20220), .ZN(n20221) );
  NOR2_X1 U23219 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20254), .ZN(
        n20243) );
  NOR3_X1 U23220 ( .A1(n20221), .A2(n20243), .A3(n20607), .ZN(n20224) );
  AOI211_X2 U23221 ( .C1(n20222), .C2(n20607), .A(n20306), .B(n20224), .ZN(
        n20244) );
  AOI22_X1 U23222 ( .A1(n20244), .A2(n13591), .B1(n20548), .B2(n20243), .ZN(
        n20230) );
  INV_X1 U23223 ( .A(n20222), .ZN(n20228) );
  AOI21_X1 U23224 ( .B1(n20223), .B2(n20276), .A(n11033), .ZN(n20227) );
  INV_X1 U23225 ( .A(n20243), .ZN(n20225) );
  AOI211_X1 U23226 ( .C1(P2_STATE2_REG_3__SCAN_IN), .C2(n20225), .A(n20551), 
        .B(n20224), .ZN(n20226) );
  AOI22_X1 U23227 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n20246), .B1(
        n20245), .B2(n20557), .ZN(n20229) );
  OAI211_X1 U23228 ( .C1(n20560), .C2(n20276), .A(n20230), .B(n20229), .ZN(
        P2_U3080) );
  AOI22_X1 U23229 ( .A1(n20244), .A2(n20089), .B1(n20087), .B2(n20243), .ZN(
        n20232) );
  AOI22_X1 U23230 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n20246), .B1(
        n20245), .B2(n20561), .ZN(n20231) );
  OAI211_X1 U23231 ( .C1(n20564), .C2(n20276), .A(n20232), .B(n20231), .ZN(
        P2_U3081) );
  AOI22_X1 U23232 ( .A1(n20244), .A2(n20093), .B1(n20565), .B2(n20243), .ZN(
        n20234) );
  AOI22_X1 U23233 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n20246), .B1(
        n20245), .B2(n20524), .ZN(n20233) );
  OAI211_X1 U23234 ( .C1(n20527), .C2(n20276), .A(n20234), .B(n20233), .ZN(
        P2_U3082) );
  AOI22_X1 U23235 ( .A1(n20244), .A2(n20571), .B1(n20570), .B2(n20243), .ZN(
        n20236) );
  AOI22_X1 U23236 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n20246), .B1(
        n20245), .B2(n20572), .ZN(n20235) );
  OAI211_X1 U23237 ( .C1(n20575), .C2(n20276), .A(n20236), .B(n20235), .ZN(
        P2_U3083) );
  AOI22_X1 U23238 ( .A1(n20244), .A2(n20577), .B1(n20576), .B2(n20243), .ZN(
        n20238) );
  AOI22_X1 U23239 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n20246), .B1(
        n20245), .B2(n20492), .ZN(n20237) );
  OAI211_X1 U23240 ( .C1(n20495), .C2(n20276), .A(n20238), .B(n20237), .ZN(
        P2_U3084) );
  AOI22_X1 U23241 ( .A1(n20244), .A2(n20585), .B1(n20584), .B2(n20243), .ZN(
        n20240) );
  AOI22_X1 U23242 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n20246), .B1(
        n20245), .B2(n20586), .ZN(n20239) );
  OAI211_X1 U23243 ( .C1(n20589), .C2(n20276), .A(n20240), .B(n20239), .ZN(
        P2_U3085) );
  AOI22_X1 U23244 ( .A1(n20244), .A2(n20591), .B1(n21297), .B2(n20243), .ZN(
        n20242) );
  AOI22_X1 U23245 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n20246), .B1(
        n20245), .B2(n20592), .ZN(n20241) );
  OAI211_X1 U23246 ( .C1(n20595), .C2(n20276), .A(n20242), .B(n20241), .ZN(
        P2_U3086) );
  AOI22_X1 U23247 ( .A1(n20244), .A2(n20598), .B1(n20596), .B2(n20243), .ZN(
        n20248) );
  AOI22_X1 U23248 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n20246), .B1(
        n20245), .B2(n20600), .ZN(n20247) );
  OAI211_X1 U23249 ( .C1(n20606), .C2(n20276), .A(n20248), .B(n20247), .ZN(
        P2_U3087) );
  AOI22_X1 U23250 ( .A1(n20286), .A2(n20506), .B1(n20548), .B2(n20271), .ZN(
        n20257) );
  OAI21_X1 U23251 ( .B1(n20297), .B2(n20473), .A(n20699), .ZN(n20255) );
  INV_X1 U23252 ( .A(n20254), .ZN(n20251) );
  INV_X1 U23253 ( .A(n20271), .ZN(n20249) );
  OAI211_X1 U23254 ( .C1(n10611), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n20249), 
        .B(n20509), .ZN(n20250) );
  OAI211_X1 U23255 ( .C1(n20255), .C2(n20251), .A(n20512), .B(n20250), .ZN(
        n20273) );
  OAI21_X1 U23256 ( .B1(n20252), .B2(n20271), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20253) );
  OAI21_X1 U23257 ( .B1(n20255), .B2(n20254), .A(n20253), .ZN(n20272) );
  AOI22_X1 U23258 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n20273), .B1(
        n13591), .B2(n20272), .ZN(n20256) );
  OAI211_X1 U23259 ( .C1(n20521), .C2(n20276), .A(n20257), .B(n20256), .ZN(
        P2_U3088) );
  INV_X1 U23260 ( .A(n20276), .ZN(n20264) );
  AOI22_X1 U23261 ( .A1(n20561), .A2(n20264), .B1(n20087), .B2(n20271), .ZN(
        n20259) );
  AOI22_X1 U23262 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n20273), .B1(
        n20089), .B2(n20272), .ZN(n20258) );
  OAI211_X1 U23263 ( .C1(n20564), .C2(n20296), .A(n20259), .B(n20258), .ZN(
        P2_U3089) );
  AOI22_X1 U23264 ( .A1(n20524), .A2(n20264), .B1(n20565), .B2(n20271), .ZN(
        n20261) );
  AOI22_X1 U23265 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n20273), .B1(
        n20093), .B2(n20272), .ZN(n20260) );
  OAI211_X1 U23266 ( .C1(n20527), .C2(n20296), .A(n20261), .B(n20260), .ZN(
        P2_U3090) );
  AOI22_X1 U23267 ( .A1(n20455), .A2(n20286), .B1(n20271), .B2(n20570), .ZN(
        n20263) );
  AOI22_X1 U23268 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20273), .B1(
        n20571), .B2(n20272), .ZN(n20262) );
  OAI211_X1 U23269 ( .C1(n20433), .C2(n20276), .A(n20263), .B(n20262), .ZN(
        P2_U3091) );
  AOI22_X1 U23270 ( .A1(n20492), .A2(n20264), .B1(n20271), .B2(n20576), .ZN(
        n20266) );
  AOI22_X1 U23271 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n20273), .B1(
        n20577), .B2(n20272), .ZN(n20265) );
  OAI211_X1 U23272 ( .C1(n20495), .C2(n20296), .A(n20266), .B(n20265), .ZN(
        P2_U3092) );
  AOI22_X1 U23273 ( .A1(n20460), .A2(n20286), .B1(n20271), .B2(n20584), .ZN(
        n20268) );
  AOI22_X1 U23274 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20273), .B1(
        n20585), .B2(n20272), .ZN(n20267) );
  OAI211_X1 U23275 ( .C1(n20438), .C2(n20276), .A(n20268), .B(n20267), .ZN(
        P2_U3093) );
  AOI22_X1 U23276 ( .A1(n20286), .A2(n20534), .B1(n20271), .B2(n21297), .ZN(
        n20270) );
  AOI22_X1 U23277 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n20273), .B1(
        n20591), .B2(n20272), .ZN(n20269) );
  OAI211_X1 U23278 ( .C1(n20538), .C2(n20276), .A(n20270), .B(n20269), .ZN(
        P2_U3094) );
  AOI22_X1 U23279 ( .A1(n20286), .A2(n20468), .B1(n20271), .B2(n20596), .ZN(
        n20275) );
  AOI22_X1 U23280 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n20273), .B1(
        n20598), .B2(n20272), .ZN(n20274) );
  OAI211_X1 U23281 ( .C1(n20396), .C2(n20276), .A(n20275), .B(n20274), .ZN(
        P2_U3095) );
  AOI22_X1 U23282 ( .A1(n20292), .A2(n20089), .B1(n20087), .B2(n20291), .ZN(
        n20279) );
  INV_X1 U23283 ( .A(n20277), .ZN(n20293) );
  AOI22_X1 U23284 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n20293), .B1(
        n20286), .B2(n20561), .ZN(n20278) );
  OAI211_X1 U23285 ( .C1(n20564), .C2(n20325), .A(n20279), .B(n20278), .ZN(
        P2_U3097) );
  AOI22_X1 U23286 ( .A1(n20292), .A2(n20093), .B1(n20565), .B2(n20291), .ZN(
        n20281) );
  AOI22_X1 U23287 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n20293), .B1(
        n20327), .B2(n20566), .ZN(n20280) );
  OAI211_X1 U23288 ( .C1(n20569), .C2(n20296), .A(n20281), .B(n20280), .ZN(
        P2_U3098) );
  AOI22_X1 U23289 ( .A1(n20292), .A2(n20571), .B1(n20570), .B2(n20291), .ZN(
        n20283) );
  AOI22_X1 U23290 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n20293), .B1(
        n20327), .B2(n20455), .ZN(n20282) );
  OAI211_X1 U23291 ( .C1(n20433), .C2(n20296), .A(n20283), .B(n20282), .ZN(
        P2_U3099) );
  AOI22_X1 U23292 ( .A1(n20292), .A2(n20577), .B1(n20576), .B2(n20291), .ZN(
        n20285) );
  AOI22_X1 U23293 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n20293), .B1(
        n20327), .B2(n20578), .ZN(n20284) );
  OAI211_X1 U23294 ( .C1(n20583), .C2(n20296), .A(n20285), .B(n20284), .ZN(
        P2_U3100) );
  AOI22_X1 U23295 ( .A1(n20292), .A2(n20585), .B1(n20584), .B2(n20291), .ZN(
        n20288) );
  AOI22_X1 U23296 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n20293), .B1(
        n20286), .B2(n20586), .ZN(n20287) );
  OAI211_X1 U23297 ( .C1(n20589), .C2(n20325), .A(n20288), .B(n20287), .ZN(
        P2_U3101) );
  AOI22_X1 U23298 ( .A1(n20292), .A2(n20591), .B1(n21297), .B2(n20291), .ZN(
        n20290) );
  AOI22_X1 U23299 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n20293), .B1(
        n20327), .B2(n20534), .ZN(n20289) );
  OAI211_X1 U23300 ( .C1(n20538), .C2(n20296), .A(n20290), .B(n20289), .ZN(
        P2_U3102) );
  AOI22_X1 U23301 ( .A1(n20292), .A2(n20598), .B1(n20596), .B2(n20291), .ZN(
        n20295) );
  AOI22_X1 U23302 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n20293), .B1(
        n20327), .B2(n20468), .ZN(n20294) );
  OAI211_X1 U23303 ( .C1(n20396), .C2(n20296), .A(n20295), .B(n20294), .ZN(
        P2_U3103) );
  NOR2_X1 U23304 ( .A1(n20297), .A2(n20308), .ZN(n20698) );
  OAI21_X1 U23305 ( .B1(n20298), .B2(n20698), .A(n20512), .ZN(n20303) );
  NAND2_X1 U23306 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20298), .ZN(
        n20335) );
  AND2_X1 U23307 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n20335), .ZN(n20299) );
  NAND2_X1 U23308 ( .A1(n20300), .A2(n20299), .ZN(n20304) );
  NAND2_X1 U23309 ( .A1(n20335), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n20301) );
  NAND2_X1 U23310 ( .A1(n20304), .A2(n20301), .ZN(n20302) );
  INV_X1 U23311 ( .A(n20328), .ZN(n20318) );
  INV_X1 U23312 ( .A(n20304), .ZN(n20305) );
  AOI211_X2 U23313 ( .C1(n20307), .C2(n20607), .A(n20306), .B(n20305), .ZN(
        n20326) );
  INV_X1 U23314 ( .A(n20335), .ZN(n20338) );
  AOI22_X1 U23315 ( .A1(n20326), .A2(n13591), .B1(n20548), .B2(n20338), .ZN(
        n20311) );
  NOR2_X2 U23316 ( .A1(n20309), .A2(n20308), .ZN(n20354) );
  AOI22_X1 U23317 ( .A1(n20354), .A2(n20506), .B1(n20327), .B2(n20557), .ZN(
        n20310) );
  OAI211_X1 U23318 ( .C1(n20318), .C2(n11802), .A(n20311), .B(n20310), .ZN(
        P2_U3104) );
  AOI22_X1 U23319 ( .A1(n20326), .A2(n20089), .B1(n20087), .B2(n20338), .ZN(
        n20313) );
  AOI22_X1 U23320 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n20328), .B1(
        n20354), .B2(n20450), .ZN(n20312) );
  OAI211_X1 U23321 ( .C1(n20428), .C2(n20325), .A(n20313), .B(n20312), .ZN(
        P2_U3105) );
  AOI22_X1 U23322 ( .A1(n20326), .A2(n20093), .B1(n20565), .B2(n20338), .ZN(
        n20315) );
  AOI22_X1 U23323 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n20328), .B1(
        n20354), .B2(n20566), .ZN(n20314) );
  OAI211_X1 U23324 ( .C1(n20569), .C2(n20325), .A(n20315), .B(n20314), .ZN(
        P2_U3106) );
  AOI22_X1 U23325 ( .A1(n20326), .A2(n20571), .B1(n20570), .B2(n20338), .ZN(
        n20317) );
  AOI22_X1 U23326 ( .A1(n20354), .A2(n20455), .B1(n20327), .B2(n20572), .ZN(
        n20316) );
  OAI211_X1 U23327 ( .C1(n20318), .C2(n10452), .A(n20317), .B(n20316), .ZN(
        P2_U3107) );
  AOI22_X1 U23328 ( .A1(n20326), .A2(n20577), .B1(n20576), .B2(n20338), .ZN(
        n20320) );
  AOI22_X1 U23329 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n20328), .B1(
        n20354), .B2(n20578), .ZN(n20319) );
  OAI211_X1 U23330 ( .C1(n20583), .C2(n20325), .A(n20320), .B(n20319), .ZN(
        P2_U3108) );
  AOI22_X1 U23331 ( .A1(n20326), .A2(n20585), .B1(n20584), .B2(n20338), .ZN(
        n20322) );
  AOI22_X1 U23332 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n20328), .B1(
        n20327), .B2(n20586), .ZN(n20321) );
  OAI211_X1 U23333 ( .C1(n20589), .C2(n20362), .A(n20322), .B(n20321), .ZN(
        P2_U3109) );
  AOI22_X1 U23334 ( .A1(n20326), .A2(n20591), .B1(n21297), .B2(n20338), .ZN(
        n20324) );
  AOI22_X1 U23335 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n20328), .B1(
        n20354), .B2(n20534), .ZN(n20323) );
  OAI211_X1 U23336 ( .C1(n20538), .C2(n20325), .A(n20324), .B(n20323), .ZN(
        P2_U3110) );
  AOI22_X1 U23337 ( .A1(n20326), .A2(n20598), .B1(n20596), .B2(n20338), .ZN(
        n20330) );
  AOI22_X1 U23338 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n20328), .B1(
        n20327), .B2(n20600), .ZN(n20329) );
  OAI211_X1 U23339 ( .C1(n20606), .C2(n20362), .A(n20330), .B(n20329), .ZN(
        P2_U3111) );
  NAND2_X1 U23340 ( .A1(n20331), .A2(n20721), .ZN(n20373) );
  NOR2_X1 U23341 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20373), .ZN(
        n20357) );
  AOI22_X1 U23342 ( .A1(n20354), .A2(n20557), .B1(n20548), .B2(n20357), .ZN(
        n20343) );
  NAND2_X1 U23343 ( .A1(n20362), .A2(n20395), .ZN(n20332) );
  AOI21_X1 U23344 ( .B1(n20332), .B2(P2_STATEBS16_REG_SCAN_IN), .A(n20509), 
        .ZN(n20337) );
  INV_X1 U23345 ( .A(n10616), .ZN(n20339) );
  OAI21_X1 U23346 ( .B1(n20339), .B2(n20607), .A(n20333), .ZN(n20334) );
  AOI21_X1 U23347 ( .B1(n20337), .B2(n20335), .A(n20334), .ZN(n20336) );
  OAI21_X1 U23348 ( .B1(n20357), .B2(n20338), .A(n20337), .ZN(n20341) );
  OAI21_X1 U23349 ( .B1(n20339), .B2(n20357), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20340) );
  NAND2_X1 U23350 ( .A1(n20341), .A2(n20340), .ZN(n20358) );
  AOI22_X1 U23351 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n20359), .B1(
        n13591), .B2(n20358), .ZN(n20342) );
  OAI211_X1 U23352 ( .C1(n20560), .C2(n20395), .A(n20343), .B(n20342), .ZN(
        P2_U3112) );
  AOI22_X1 U23353 ( .A1(n20354), .A2(n20561), .B1(n20087), .B2(n20357), .ZN(
        n20345) );
  AOI22_X1 U23354 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n20359), .B1(
        n20358), .B2(n20089), .ZN(n20344) );
  OAI211_X1 U23355 ( .C1(n20564), .C2(n20395), .A(n20345), .B(n20344), .ZN(
        P2_U3113) );
  AOI22_X1 U23356 ( .A1(n20354), .A2(n20524), .B1(n20565), .B2(n20357), .ZN(
        n20347) );
  AOI22_X1 U23357 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n20359), .B1(
        n20358), .B2(n20093), .ZN(n20346) );
  OAI211_X1 U23358 ( .C1(n20527), .C2(n20395), .A(n20347), .B(n20346), .ZN(
        P2_U3114) );
  AOI22_X1 U23359 ( .A1(n20455), .A2(n20383), .B1(n20570), .B2(n20357), .ZN(
        n20349) );
  AOI22_X1 U23360 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n20359), .B1(
        n20358), .B2(n20571), .ZN(n20348) );
  OAI211_X1 U23361 ( .C1(n20433), .C2(n20362), .A(n20349), .B(n20348), .ZN(
        P2_U3115) );
  AOI22_X1 U23362 ( .A1(n20492), .A2(n20354), .B1(n20576), .B2(n20357), .ZN(
        n20351) );
  AOI22_X1 U23363 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n20359), .B1(
        n20358), .B2(n20577), .ZN(n20350) );
  OAI211_X1 U23364 ( .C1(n20495), .C2(n20395), .A(n20351), .B(n20350), .ZN(
        P2_U3116) );
  AOI22_X1 U23365 ( .A1(n20460), .A2(n20383), .B1(n20584), .B2(n20357), .ZN(
        n20353) );
  AOI22_X1 U23366 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n20359), .B1(
        n20358), .B2(n20585), .ZN(n20352) );
  OAI211_X1 U23367 ( .C1(n20438), .C2(n20362), .A(n20353), .B(n20352), .ZN(
        P2_U3117) );
  AOI22_X1 U23368 ( .A1(n20592), .A2(n20354), .B1(n21297), .B2(n20357), .ZN(
        n20356) );
  AOI22_X1 U23369 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n20359), .B1(
        n20358), .B2(n20591), .ZN(n20355) );
  OAI211_X1 U23370 ( .C1(n20595), .C2(n20395), .A(n20356), .B(n20355), .ZN(
        P2_U3118) );
  AOI22_X1 U23371 ( .A1(n20468), .A2(n20383), .B1(n20596), .B2(n20357), .ZN(
        n20361) );
  AOI22_X1 U23372 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n20359), .B1(
        n20358), .B2(n20598), .ZN(n20360) );
  OAI211_X1 U23373 ( .C1(n20396), .C2(n20362), .A(n20361), .B(n20360), .ZN(
        P2_U3119) );
  NOR2_X1 U23374 ( .A1(n20364), .A2(n20401), .ZN(n20402) );
  AOI22_X1 U23375 ( .A1(n20383), .A2(n20557), .B1(n20548), .B2(n20402), .ZN(
        n20376) );
  AOI21_X1 U23376 ( .B1(n20554), .B2(n20365), .A(n20509), .ZN(n20370) );
  INV_X1 U23377 ( .A(n20402), .ZN(n20366) );
  NAND2_X1 U23378 ( .A1(n20367), .A2(n20366), .ZN(n20371) );
  NOR2_X1 U23379 ( .A1(n20371), .A2(n20607), .ZN(n20368) );
  AOI21_X1 U23380 ( .B1(n20370), .B2(n20373), .A(n20368), .ZN(n20369) );
  OAI211_X1 U23381 ( .C1(n20402), .C2(n20333), .A(n20369), .B(n20512), .ZN(
        n20392) );
  INV_X1 U23382 ( .A(n20370), .ZN(n20374) );
  INV_X1 U23383 ( .A(n20371), .ZN(n20372) );
  OAI22_X1 U23384 ( .A1(n20374), .A2(n20373), .B1(n20372), .B2(n20607), .ZN(
        n20391) );
  AOI22_X1 U23385 ( .A1(P2_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n20392), .B1(
        n13591), .B2(n20391), .ZN(n20375) );
  OAI211_X1 U23386 ( .C1(n20560), .C2(n20386), .A(n20376), .B(n20375), .ZN(
        P2_U3120) );
  AOI22_X1 U23387 ( .A1(n20450), .A2(n20422), .B1(n20087), .B2(n20402), .ZN(
        n20378) );
  AOI22_X1 U23388 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n20392), .B1(
        n20089), .B2(n20391), .ZN(n20377) );
  OAI211_X1 U23389 ( .C1(n20428), .C2(n20395), .A(n20378), .B(n20377), .ZN(
        P2_U3121) );
  AOI22_X1 U23390 ( .A1(n20566), .A2(n20422), .B1(n20565), .B2(n20402), .ZN(
        n20380) );
  AOI22_X1 U23391 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n20392), .B1(
        n20093), .B2(n20391), .ZN(n20379) );
  OAI211_X1 U23392 ( .C1(n20569), .C2(n20395), .A(n20380), .B(n20379), .ZN(
        P2_U3122) );
  AOI22_X1 U23393 ( .A1(n20572), .A2(n20383), .B1(n20570), .B2(n20402), .ZN(
        n20382) );
  AOI22_X1 U23394 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n20392), .B1(
        n20571), .B2(n20391), .ZN(n20381) );
  OAI211_X1 U23395 ( .C1(n20575), .C2(n20386), .A(n20382), .B(n20381), .ZN(
        P2_U3123) );
  AOI22_X1 U23396 ( .A1(n20492), .A2(n20383), .B1(n20576), .B2(n20402), .ZN(
        n20385) );
  AOI22_X1 U23397 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n20392), .B1(
        n20577), .B2(n20391), .ZN(n20384) );
  OAI211_X1 U23398 ( .C1(n20495), .C2(n20386), .A(n20385), .B(n20384), .ZN(
        P2_U3124) );
  AOI22_X1 U23399 ( .A1(n20460), .A2(n20422), .B1(n20584), .B2(n20402), .ZN(
        n20388) );
  AOI22_X1 U23400 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n20392), .B1(
        n20585), .B2(n20391), .ZN(n20387) );
  OAI211_X1 U23401 ( .C1(n20438), .C2(n20395), .A(n20388), .B(n20387), .ZN(
        P2_U3125) );
  AOI22_X1 U23402 ( .A1(n20534), .A2(n20422), .B1(n21297), .B2(n20402), .ZN(
        n20390) );
  AOI22_X1 U23403 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n20392), .B1(
        n20591), .B2(n20391), .ZN(n20389) );
  OAI211_X1 U23404 ( .C1(n20538), .C2(n20395), .A(n20390), .B(n20389), .ZN(
        P2_U3126) );
  AOI22_X1 U23405 ( .A1(n20468), .A2(n20422), .B1(n20596), .B2(n20402), .ZN(
        n20394) );
  AOI22_X1 U23406 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n20392), .B1(
        n20598), .B2(n20391), .ZN(n20393) );
  OAI211_X1 U23407 ( .C1(n20396), .C2(n20395), .A(n20394), .B(n20393), .ZN(
        P2_U3127) );
  INV_X1 U23408 ( .A(n20404), .ZN(n20398) );
  NOR2_X1 U23409 ( .A1(n20397), .A2(n20401), .ZN(n20420) );
  OAI21_X1 U23410 ( .B1(n20398), .B2(n20420), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20399) );
  OAI21_X1 U23411 ( .B1(n20401), .B2(n20400), .A(n20399), .ZN(n20421) );
  AOI22_X1 U23412 ( .A1(n20421), .A2(n13591), .B1(n20548), .B2(n20420), .ZN(
        n20407) );
  AOI221_X1 U23413 ( .B1(n20445), .B2(P2_STATEBS16_REG_SCAN_IN), .C1(n20422), 
        .C2(P2_STATEBS16_REG_SCAN_IN), .A(n20402), .ZN(n20403) );
  AOI211_X1 U23414 ( .C1(n20404), .C2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .B(n20403), .ZN(n20405) );
  AOI22_X1 U23415 ( .A1(P2_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n20423), .B1(
        n20422), .B2(n20557), .ZN(n20406) );
  OAI211_X1 U23416 ( .C1(n20560), .C2(n20442), .A(n20407), .B(n20406), .ZN(
        P2_U3128) );
  AOI22_X1 U23417 ( .A1(n20421), .A2(n20089), .B1(n20087), .B2(n20420), .ZN(
        n20409) );
  AOI22_X1 U23418 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n20423), .B1(
        n20422), .B2(n20561), .ZN(n20408) );
  OAI211_X1 U23419 ( .C1(n20564), .C2(n20442), .A(n20409), .B(n20408), .ZN(
        P2_U3129) );
  AOI22_X1 U23420 ( .A1(n20421), .A2(n20093), .B1(n20565), .B2(n20420), .ZN(
        n20411) );
  AOI22_X1 U23421 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n20423), .B1(
        n20422), .B2(n20524), .ZN(n20410) );
  OAI211_X1 U23422 ( .C1(n20527), .C2(n20442), .A(n20411), .B(n20410), .ZN(
        P2_U3130) );
  AOI22_X1 U23423 ( .A1(n20421), .A2(n20571), .B1(n20570), .B2(n20420), .ZN(
        n20413) );
  AOI22_X1 U23424 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n20423), .B1(
        n20422), .B2(n20572), .ZN(n20412) );
  OAI211_X1 U23425 ( .C1(n20575), .C2(n20442), .A(n20413), .B(n20412), .ZN(
        P2_U3131) );
  AOI22_X1 U23426 ( .A1(n20421), .A2(n20577), .B1(n20576), .B2(n20420), .ZN(
        n20415) );
  AOI22_X1 U23427 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n20423), .B1(
        n20422), .B2(n20492), .ZN(n20414) );
  OAI211_X1 U23428 ( .C1(n20495), .C2(n20442), .A(n20415), .B(n20414), .ZN(
        P2_U3132) );
  AOI22_X1 U23429 ( .A1(n20421), .A2(n20585), .B1(n20584), .B2(n20420), .ZN(
        n20417) );
  AOI22_X1 U23430 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n20423), .B1(
        n20422), .B2(n20586), .ZN(n20416) );
  OAI211_X1 U23431 ( .C1(n20589), .C2(n20442), .A(n20417), .B(n20416), .ZN(
        P2_U3133) );
  AOI22_X1 U23432 ( .A1(n20421), .A2(n20591), .B1(n21297), .B2(n20420), .ZN(
        n20419) );
  AOI22_X1 U23433 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n20423), .B1(
        n20422), .B2(n20592), .ZN(n20418) );
  OAI211_X1 U23434 ( .C1(n20595), .C2(n20442), .A(n20419), .B(n20418), .ZN(
        P2_U3134) );
  AOI22_X1 U23435 ( .A1(n20421), .A2(n20598), .B1(n20596), .B2(n20420), .ZN(
        n20425) );
  AOI22_X1 U23436 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n20423), .B1(
        n20422), .B2(n20600), .ZN(n20424) );
  OAI211_X1 U23437 ( .C1(n20606), .C2(n20442), .A(n20425), .B(n20424), .ZN(
        P2_U3135) );
  AOI22_X1 U23438 ( .A1(n20444), .A2(n20089), .B1(n20443), .B2(n20087), .ZN(
        n20427) );
  AOI22_X1 U23439 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n20439), .B1(
        n20467), .B2(n20450), .ZN(n20426) );
  OAI211_X1 U23440 ( .C1(n20428), .C2(n20442), .A(n20427), .B(n20426), .ZN(
        P2_U3137) );
  AOI22_X1 U23441 ( .A1(n20444), .A2(n20093), .B1(n20443), .B2(n20565), .ZN(
        n20430) );
  AOI22_X1 U23442 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n20439), .B1(
        n20467), .B2(n20566), .ZN(n20429) );
  OAI211_X1 U23443 ( .C1(n20569), .C2(n20442), .A(n20430), .B(n20429), .ZN(
        P2_U3138) );
  AOI22_X1 U23444 ( .A1(n20444), .A2(n20571), .B1(n20443), .B2(n20570), .ZN(
        n20432) );
  AOI22_X1 U23445 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n20439), .B1(
        n20467), .B2(n20455), .ZN(n20431) );
  OAI211_X1 U23446 ( .C1(n20433), .C2(n20442), .A(n20432), .B(n20431), .ZN(
        P2_U3139) );
  AOI22_X1 U23447 ( .A1(n20444), .A2(n20577), .B1(n20443), .B2(n20576), .ZN(
        n20435) );
  AOI22_X1 U23448 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n20439), .B1(
        n20467), .B2(n20578), .ZN(n20434) );
  OAI211_X1 U23449 ( .C1(n20583), .C2(n20442), .A(n20435), .B(n20434), .ZN(
        P2_U3140) );
  AOI22_X1 U23450 ( .A1(n20444), .A2(n20585), .B1(n20443), .B2(n20584), .ZN(
        n20437) );
  AOI22_X1 U23451 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n20439), .B1(
        n20467), .B2(n20460), .ZN(n20436) );
  OAI211_X1 U23452 ( .C1(n20438), .C2(n20442), .A(n20437), .B(n20436), .ZN(
        P2_U3141) );
  AOI22_X1 U23453 ( .A1(n20444), .A2(n20591), .B1(n20443), .B2(n21297), .ZN(
        n20441) );
  AOI22_X1 U23454 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n20439), .B1(
        n20467), .B2(n20534), .ZN(n20440) );
  OAI211_X1 U23455 ( .C1(n20538), .C2(n20442), .A(n20441), .B(n20440), .ZN(
        P2_U3142) );
  AOI22_X1 U23456 ( .A1(n20444), .A2(n20598), .B1(n20443), .B2(n20596), .ZN(
        n20447) );
  AOI22_X1 U23457 ( .A1(n20467), .A2(n20468), .B1(n20445), .B2(n20600), .ZN(
        n20446) );
  OAI211_X1 U23458 ( .C1(n20449), .C2(n20448), .A(n20447), .B(n20446), .ZN(
        P2_U3143) );
  AOI22_X1 U23459 ( .A1(n20466), .A2(n20089), .B1(n20465), .B2(n20087), .ZN(
        n20452) );
  AOI22_X1 U23460 ( .A1(n20467), .A2(n20561), .B1(n20501), .B2(n20450), .ZN(
        n20451) );
  OAI211_X1 U23461 ( .C1(n20472), .C2(n10472), .A(n20452), .B(n20451), .ZN(
        P2_U3145) );
  AOI22_X1 U23462 ( .A1(n20466), .A2(n20093), .B1(n20465), .B2(n20565), .ZN(
        n20454) );
  AOI22_X1 U23463 ( .A1(n20467), .A2(n20524), .B1(n20501), .B2(n20566), .ZN(
        n20453) );
  OAI211_X1 U23464 ( .C1(n20472), .C2(n15015), .A(n20454), .B(n20453), .ZN(
        P2_U3146) );
  AOI22_X1 U23465 ( .A1(n20466), .A2(n20571), .B1(n20465), .B2(n20570), .ZN(
        n20457) );
  AOI22_X1 U23466 ( .A1(n20501), .A2(n20455), .B1(n20467), .B2(n20572), .ZN(
        n20456) );
  OAI211_X1 U23467 ( .C1(n20472), .C2(n15037), .A(n20457), .B(n20456), .ZN(
        P2_U3147) );
  AOI22_X1 U23468 ( .A1(n20466), .A2(n20577), .B1(n20465), .B2(n20576), .ZN(
        n20459) );
  AOI22_X1 U23469 ( .A1(n20467), .A2(n20492), .B1(n20501), .B2(n20578), .ZN(
        n20458) );
  OAI211_X1 U23470 ( .C1(n20472), .C2(n15065), .A(n20459), .B(n20458), .ZN(
        P2_U3148) );
  AOI22_X1 U23471 ( .A1(n20466), .A2(n20585), .B1(n20465), .B2(n20584), .ZN(
        n20462) );
  AOI22_X1 U23472 ( .A1(n20501), .A2(n20460), .B1(n20467), .B2(n20586), .ZN(
        n20461) );
  OAI211_X1 U23473 ( .C1(n20472), .C2(n15090), .A(n20462), .B(n20461), .ZN(
        P2_U3149) );
  AOI22_X1 U23474 ( .A1(n20466), .A2(n20591), .B1(n20465), .B2(n21297), .ZN(
        n20464) );
  AOI22_X1 U23475 ( .A1(n20467), .A2(n20592), .B1(n20501), .B2(n20534), .ZN(
        n20463) );
  OAI211_X1 U23476 ( .C1(n20472), .C2(n10669), .A(n20464), .B(n20463), .ZN(
        P2_U3150) );
  INV_X1 U23477 ( .A(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n20471) );
  AOI22_X1 U23478 ( .A1(n20466), .A2(n20598), .B1(n20465), .B2(n20596), .ZN(
        n20470) );
  AOI22_X1 U23479 ( .A1(n20501), .A2(n20468), .B1(n20467), .B2(n20600), .ZN(
        n20469) );
  OAI211_X1 U23480 ( .C1(n20472), .C2(n20471), .A(n20470), .B(n20469), .ZN(
        P2_U3151) );
  OR2_X1 U23481 ( .A1(n20475), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n20478) );
  INV_X1 U23482 ( .A(n20476), .ZN(n20477) );
  NAND2_X1 U23483 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20483), .ZN(
        n20480) );
  INV_X1 U23484 ( .A(n20480), .ZN(n20508) );
  NOR3_X1 U23485 ( .A1(n20477), .A2(n20508), .A3(n20607), .ZN(n20479) );
  AOI21_X1 U23486 ( .B1(n20607), .B2(n20478), .A(n20479), .ZN(n20500) );
  AOI22_X1 U23487 ( .A1(n20500), .A2(n13591), .B1(n20548), .B2(n20508), .ZN(
        n20485) );
  AOI211_X1 U23488 ( .C1(P2_STATE2_REG_3__SCAN_IN), .C2(n20480), .A(n20551), 
        .B(n20479), .ZN(n20481) );
  OAI221_X1 U23489 ( .B1(n20483), .B2(n20482), .C1(n20483), .C2(n20554), .A(
        n20481), .ZN(n20502) );
  AOI22_X1 U23490 ( .A1(P2_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n20502), .B1(
        n20501), .B2(n20557), .ZN(n20484) );
  OAI211_X1 U23491 ( .C1(n20560), .C2(n20537), .A(n20485), .B(n20484), .ZN(
        P2_U3152) );
  AOI22_X1 U23492 ( .A1(n20500), .A2(n20089), .B1(n20087), .B2(n20508), .ZN(
        n20487) );
  AOI22_X1 U23493 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n20502), .B1(
        n20501), .B2(n20561), .ZN(n20486) );
  OAI211_X1 U23494 ( .C1(n20564), .C2(n20537), .A(n20487), .B(n20486), .ZN(
        P2_U3153) );
  AOI22_X1 U23495 ( .A1(n20500), .A2(n20093), .B1(n20565), .B2(n20508), .ZN(
        n20489) );
  AOI22_X1 U23496 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n20502), .B1(
        n20501), .B2(n20524), .ZN(n20488) );
  OAI211_X1 U23497 ( .C1(n20527), .C2(n20537), .A(n20489), .B(n20488), .ZN(
        P2_U3154) );
  AOI22_X1 U23498 ( .A1(n20500), .A2(n20571), .B1(n20570), .B2(n20508), .ZN(
        n20491) );
  AOI22_X1 U23499 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n20502), .B1(
        n20501), .B2(n20572), .ZN(n20490) );
  OAI211_X1 U23500 ( .C1(n20575), .C2(n20537), .A(n20491), .B(n20490), .ZN(
        P2_U3155) );
  AOI22_X1 U23501 ( .A1(n20500), .A2(n20577), .B1(n20576), .B2(n20508), .ZN(
        n20494) );
  AOI22_X1 U23502 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n20502), .B1(
        n20501), .B2(n20492), .ZN(n20493) );
  OAI211_X1 U23503 ( .C1(n20495), .C2(n20537), .A(n20494), .B(n20493), .ZN(
        P2_U3156) );
  AOI22_X1 U23504 ( .A1(n20500), .A2(n20585), .B1(n20584), .B2(n20508), .ZN(
        n20497) );
  AOI22_X1 U23505 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n20502), .B1(
        n20501), .B2(n20586), .ZN(n20496) );
  OAI211_X1 U23506 ( .C1(n20589), .C2(n20537), .A(n20497), .B(n20496), .ZN(
        P2_U3157) );
  AOI22_X1 U23507 ( .A1(n20500), .A2(n20591), .B1(n21297), .B2(n20508), .ZN(
        n20499) );
  AOI22_X1 U23508 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n20502), .B1(
        n20501), .B2(n20592), .ZN(n20498) );
  OAI211_X1 U23509 ( .C1(n20595), .C2(n20537), .A(n20499), .B(n20498), .ZN(
        P2_U3158) );
  AOI22_X1 U23510 ( .A1(n20500), .A2(n20598), .B1(n20596), .B2(n20508), .ZN(
        n20504) );
  AOI22_X1 U23511 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n20502), .B1(
        n20501), .B2(n20600), .ZN(n20503) );
  OAI211_X1 U23512 ( .C1(n20606), .C2(n20537), .A(n20504), .B(n20503), .ZN(
        P2_U3159) );
  NOR3_X2 U23513 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n10567), .A3(
        n20545), .ZN(n20539) );
  AOI22_X1 U23514 ( .A1(n20506), .A2(n20601), .B1(n20548), .B2(n20539), .ZN(
        n20520) );
  OAI21_X1 U23515 ( .B1(n20601), .B2(n20540), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n20507) );
  NAND2_X1 U23516 ( .A1(n20507), .A2(n20699), .ZN(n20518) );
  NOR2_X1 U23517 ( .A1(n20539), .A2(n20508), .ZN(n20517) );
  INV_X1 U23518 ( .A(n20517), .ZN(n20513) );
  INV_X1 U23519 ( .A(n20539), .ZN(n20510) );
  OAI211_X1 U23520 ( .C1(n20514), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n20510), 
        .B(n20509), .ZN(n20511) );
  OAI211_X1 U23521 ( .C1(n20518), .C2(n20513), .A(n20512), .B(n20511), .ZN(
        n20542) );
  INV_X1 U23522 ( .A(n20514), .ZN(n20515) );
  OAI21_X1 U23523 ( .B1(n20515), .B2(n20539), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20516) );
  AOI22_X1 U23524 ( .A1(P2_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n20542), .B1(
        n13591), .B2(n20541), .ZN(n20519) );
  OAI211_X1 U23525 ( .C1(n20521), .C2(n20537), .A(n20520), .B(n20519), .ZN(
        P2_U3160) );
  AOI22_X1 U23526 ( .A1(n20561), .A2(n20540), .B1(n20087), .B2(n20539), .ZN(
        n20523) );
  AOI22_X1 U23527 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n20542), .B1(
        n20089), .B2(n20541), .ZN(n20522) );
  OAI211_X1 U23528 ( .C1(n20564), .C2(n20582), .A(n20523), .B(n20522), .ZN(
        P2_U3161) );
  AOI22_X1 U23529 ( .A1(n20524), .A2(n20540), .B1(n20565), .B2(n20539), .ZN(
        n20526) );
  AOI22_X1 U23530 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n20542), .B1(
        n20093), .B2(n20541), .ZN(n20525) );
  OAI211_X1 U23531 ( .C1(n20527), .C2(n20582), .A(n20526), .B(n20525), .ZN(
        P2_U3162) );
  AOI22_X1 U23532 ( .A1(n20572), .A2(n20540), .B1(n20570), .B2(n20539), .ZN(
        n20529) );
  AOI22_X1 U23533 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n20542), .B1(
        n20571), .B2(n20541), .ZN(n20528) );
  OAI211_X1 U23534 ( .C1(n20575), .C2(n20582), .A(n20529), .B(n20528), .ZN(
        P2_U3163) );
  AOI22_X1 U23535 ( .A1(n20578), .A2(n20601), .B1(n20576), .B2(n20539), .ZN(
        n20531) );
  AOI22_X1 U23536 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n20542), .B1(
        n20577), .B2(n20541), .ZN(n20530) );
  OAI211_X1 U23537 ( .C1(n20583), .C2(n20537), .A(n20531), .B(n20530), .ZN(
        P2_U3164) );
  AOI22_X1 U23538 ( .A1(n20586), .A2(n20540), .B1(n20584), .B2(n20539), .ZN(
        n20533) );
  AOI22_X1 U23539 ( .A1(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n20542), .B1(
        n20585), .B2(n20541), .ZN(n20532) );
  OAI211_X1 U23540 ( .C1(n20589), .C2(n20582), .A(n20533), .B(n20532), .ZN(
        P2_U3165) );
  AOI22_X1 U23541 ( .A1(n20534), .A2(n20601), .B1(n21297), .B2(n20539), .ZN(
        n20536) );
  AOI22_X1 U23542 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n20542), .B1(
        n20591), .B2(n20541), .ZN(n20535) );
  OAI211_X1 U23543 ( .C1(n20538), .C2(n20537), .A(n20536), .B(n20535), .ZN(
        P2_U3166) );
  AOI22_X1 U23544 ( .A1(n20600), .A2(n20540), .B1(n20596), .B2(n20539), .ZN(
        n20544) );
  AOI22_X1 U23545 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n20542), .B1(
        n20598), .B2(n20541), .ZN(n20543) );
  OAI211_X1 U23546 ( .C1(n20606), .C2(n20582), .A(n20544), .B(n20543), .ZN(
        P2_U3167) );
  NOR2_X1 U23547 ( .A1(n20597), .A2(n20607), .ZN(n20547) );
  NOR2_X1 U23548 ( .A1(n10567), .A2(n20545), .ZN(n20556) );
  AOI21_X1 U23549 ( .B1(n20556), .B2(n20333), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20546) );
  AOI21_X1 U23550 ( .B1(n20549), .B2(n20547), .A(n20546), .ZN(n20599) );
  AOI22_X1 U23551 ( .A1(n20599), .A2(n13591), .B1(n20597), .B2(n20548), .ZN(
        n20559) );
  INV_X1 U23552 ( .A(n20549), .ZN(n20550) );
  AOI211_X1 U23553 ( .C1(n20550), .C2(n20333), .A(n20597), .B(n20699), .ZN(
        n20552) );
  NOR2_X1 U23554 ( .A1(n20552), .A2(n20551), .ZN(n20553) );
  OAI221_X1 U23555 ( .B1(n20556), .B2(n20555), .C1(n20556), .C2(n20554), .A(
        n20553), .ZN(n20602) );
  AOI22_X1 U23556 ( .A1(P2_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n20602), .B1(
        n20601), .B2(n20557), .ZN(n20558) );
  OAI211_X1 U23557 ( .C1(n20560), .C2(n20605), .A(n20559), .B(n20558), .ZN(
        P2_U3168) );
  AOI22_X1 U23558 ( .A1(n20599), .A2(n20089), .B1(n20597), .B2(n20087), .ZN(
        n20563) );
  AOI22_X1 U23559 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n20602), .B1(
        n20601), .B2(n20561), .ZN(n20562) );
  OAI211_X1 U23560 ( .C1(n20564), .C2(n20605), .A(n20563), .B(n20562), .ZN(
        P2_U3169) );
  AOI22_X1 U23561 ( .A1(n20599), .A2(n20093), .B1(n20597), .B2(n20565), .ZN(
        n20568) );
  AOI22_X1 U23562 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n20602), .B1(
        n20579), .B2(n20566), .ZN(n20567) );
  OAI211_X1 U23563 ( .C1(n20569), .C2(n20582), .A(n20568), .B(n20567), .ZN(
        P2_U3170) );
  AOI22_X1 U23564 ( .A1(n20599), .A2(n20571), .B1(n20597), .B2(n20570), .ZN(
        n20574) );
  AOI22_X1 U23565 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n20602), .B1(
        n20601), .B2(n20572), .ZN(n20573) );
  OAI211_X1 U23566 ( .C1(n20575), .C2(n20605), .A(n20574), .B(n20573), .ZN(
        P2_U3171) );
  AOI22_X1 U23567 ( .A1(n20599), .A2(n20577), .B1(n20597), .B2(n20576), .ZN(
        n20581) );
  AOI22_X1 U23568 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n20602), .B1(
        n20579), .B2(n20578), .ZN(n20580) );
  OAI211_X1 U23569 ( .C1(n20583), .C2(n20582), .A(n20581), .B(n20580), .ZN(
        P2_U3172) );
  AOI22_X1 U23570 ( .A1(n20599), .A2(n20585), .B1(n20597), .B2(n20584), .ZN(
        n20588) );
  AOI22_X1 U23571 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n20602), .B1(
        n20601), .B2(n20586), .ZN(n20587) );
  OAI211_X1 U23572 ( .C1(n20589), .C2(n20605), .A(n20588), .B(n20587), .ZN(
        P2_U3173) );
  AOI22_X1 U23573 ( .A1(n20599), .A2(n20591), .B1(n20597), .B2(n21297), .ZN(
        n20594) );
  AOI22_X1 U23574 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n20602), .B1(
        n20601), .B2(n20592), .ZN(n20593) );
  OAI211_X1 U23575 ( .C1(n20595), .C2(n20605), .A(n20594), .B(n20593), .ZN(
        P2_U3174) );
  AOI22_X1 U23576 ( .A1(n20599), .A2(n20598), .B1(n20597), .B2(n20596), .ZN(
        n20604) );
  AOI22_X1 U23577 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n20602), .B1(
        n20601), .B2(n20600), .ZN(n20603) );
  OAI211_X1 U23578 ( .C1(n20606), .C2(n20605), .A(n20604), .B(n20603), .ZN(
        P2_U3175) );
  OAI21_X1 U23579 ( .B1(n20744), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n20607), 
        .ZN(n20608) );
  NAND2_X1 U23580 ( .A1(n20609), .A2(n20608), .ZN(n20615) );
  INV_X1 U23581 ( .A(n20610), .ZN(n20611) );
  OAI211_X1 U23582 ( .C1(n20612), .C2(n20611), .A(P2_STATE2_REG_1__SCAN_IN), 
        .B(n20744), .ZN(n20614) );
  OAI211_X1 U23583 ( .C1(n20616), .C2(n20615), .A(n20614), .B(n20613), .ZN(
        P2_U3177) );
  AND2_X1 U23584 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n20619), .ZN(
        P2_U3179) );
  AND2_X1 U23585 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n20619), .ZN(
        P2_U3180) );
  AND2_X1 U23586 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n20619), .ZN(
        P2_U3181) );
  AND2_X1 U23587 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n20619), .ZN(
        P2_U3182) );
  AND2_X1 U23588 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n20619), .ZN(
        P2_U3183) );
  AND2_X1 U23589 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n20619), .ZN(
        P2_U3184) );
  AND2_X1 U23590 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n20619), .ZN(
        P2_U3185) );
  AND2_X1 U23591 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n20619), .ZN(
        P2_U3186) );
  AND2_X1 U23592 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n20619), .ZN(
        P2_U3187) );
  AND2_X1 U23593 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n20619), .ZN(
        P2_U3188) );
  AND2_X1 U23594 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n20619), .ZN(
        P2_U3189) );
  AND2_X1 U23595 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n20619), .ZN(
        P2_U3190) );
  AND2_X1 U23596 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n20619), .ZN(
        P2_U3191) );
  AND2_X1 U23597 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n20619), .ZN(
        P2_U3192) );
  AND2_X1 U23598 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n20619), .ZN(
        P2_U3193) );
  AND2_X1 U23599 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n20619), .ZN(
        P2_U3194) );
  AND2_X1 U23600 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n20619), .ZN(
        P2_U3195) );
  AND2_X1 U23601 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n20619), .ZN(
        P2_U3196) );
  AND2_X1 U23602 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n20619), .ZN(
        P2_U3197) );
  AND2_X1 U23603 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n20619), .ZN(
        P2_U3198) );
  NOR2_X1 U23604 ( .A1(n20617), .A2(n20694), .ZN(P2_U3199) );
  AND2_X1 U23605 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n20619), .ZN(
        P2_U3200) );
  AND2_X1 U23606 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n20619), .ZN(P2_U3201) );
  NOR2_X1 U23607 ( .A1(n20618), .A2(n20694), .ZN(P2_U3202) );
  AND2_X1 U23608 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n20619), .ZN(P2_U3203) );
  AND2_X1 U23609 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n20619), .ZN(P2_U3204) );
  AND2_X1 U23610 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n20619), .ZN(P2_U3205) );
  AND2_X1 U23611 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n20619), .ZN(P2_U3206) );
  AND2_X1 U23612 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n20619), .ZN(P2_U3207) );
  NOR2_X1 U23613 ( .A1(n20620), .A2(n20694), .ZN(P2_U3208) );
  INV_X1 U23614 ( .A(NA), .ZN(n21192) );
  OAI21_X1 U23615 ( .B1(n21192), .B2(n20626), .A(P2_STATE_REG_2__SCAN_IN), 
        .ZN(n20635) );
  INV_X1 U23616 ( .A(n20635), .ZN(n20623) );
  NAND2_X1 U23617 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n20744), .ZN(n20633) );
  INV_X1 U23618 ( .A(n20633), .ZN(n20624) );
  INV_X1 U23619 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n20761) );
  NOR3_X1 U23620 ( .A1(n20624), .A2(n20761), .A3(n20625), .ZN(n20622) );
  OAI211_X1 U23621 ( .C1(HOLD), .C2(n20761), .A(n20762), .B(n20630), .ZN(
        n20621) );
  OAI21_X1 U23622 ( .B1(n20623), .B2(n20622), .A(n20621), .ZN(P2_U3209) );
  NOR2_X1 U23623 ( .A1(n20756), .A2(n20624), .ZN(n20628) );
  NOR2_X1 U23624 ( .A1(HOLD), .A2(n20625), .ZN(n20634) );
  OAI211_X1 U23625 ( .C1(n20634), .C2(n20636), .A(
        P2_REQUESTPENDING_REG_SCAN_IN), .B(n20626), .ZN(n20627) );
  OAI211_X1 U23626 ( .C1(n20629), .C2(n21186), .A(n20628), .B(n20627), .ZN(
        P2_U3210) );
  OAI22_X1 U23627 ( .A1(P2_REQUESTPENDING_REG_SCAN_IN), .A2(n20630), .B1(NA), 
        .B2(n20633), .ZN(n20631) );
  OAI211_X1 U23628 ( .C1(P2_REQUESTPENDING_REG_SCAN_IN), .C2(HOLD), .A(
        P2_STATE_REG_0__SCAN_IN), .B(n20631), .ZN(n20632) );
  OAI221_X1 U23629 ( .B1(n20635), .B2(n20634), .C1(n20635), .C2(n20633), .A(
        n20632), .ZN(P2_U3211) );
  NAND2_X1 U23630 ( .A1(n20765), .A2(n20636), .ZN(n20684) );
  CLKBUF_X1 U23631 ( .A(n20684), .Z(n20680) );
  OAI222_X1 U23632 ( .A1(n20681), .A2(n10371), .B1(n20637), .B2(n20765), .C1(
        n10380), .C2(n20680), .ZN(P2_U3212) );
  OAI222_X1 U23633 ( .A1(n20681), .A2(n10380), .B1(n20638), .B2(n20765), .C1(
        n14775), .C2(n20680), .ZN(P2_U3213) );
  OAI222_X1 U23634 ( .A1(n20681), .A2(n14775), .B1(n20639), .B2(n20765), .C1(
        n10921), .C2(n20680), .ZN(P2_U3214) );
  INV_X1 U23635 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n20641) );
  OAI222_X1 U23636 ( .A1(n20680), .A2(n20641), .B1(n20640), .B2(n20765), .C1(
        n10921), .C2(n20681), .ZN(P2_U3215) );
  OAI222_X1 U23637 ( .A1(n20684), .A2(n14389), .B1(n20642), .B2(n20765), .C1(
        n20641), .C2(n20681), .ZN(P2_U3216) );
  OAI222_X1 U23638 ( .A1(n20684), .A2(n10940), .B1(n20643), .B2(n20765), .C1(
        n14389), .C2(n20681), .ZN(P2_U3217) );
  OAI222_X1 U23639 ( .A1(n20684), .A2(n10945), .B1(n20644), .B2(n20765), .C1(
        n10940), .C2(n20681), .ZN(P2_U3218) );
  OAI222_X1 U23640 ( .A1(n20684), .A2(n14291), .B1(n20645), .B2(n20765), .C1(
        n10945), .C2(n20681), .ZN(P2_U3219) );
  OAI222_X1 U23641 ( .A1(n20684), .A2(n14248), .B1(n20646), .B2(n20765), .C1(
        n14291), .C2(n20681), .ZN(P2_U3220) );
  INV_X1 U23642 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n20648) );
  OAI222_X1 U23643 ( .A1(n20680), .A2(n20648), .B1(n20647), .B2(n20765), .C1(
        n14248), .C2(n20681), .ZN(P2_U3221) );
  OAI222_X1 U23644 ( .A1(n20680), .A2(n10962), .B1(n20649), .B2(n20765), .C1(
        n20648), .C2(n20681), .ZN(P2_U3222) );
  OAI222_X1 U23645 ( .A1(n20680), .A2(n11913), .B1(n20650), .B2(n20765), .C1(
        n10962), .C2(n20681), .ZN(P2_U3223) );
  OAI222_X1 U23646 ( .A1(n20680), .A2(n10967), .B1(n20651), .B2(n20765), .C1(
        n11913), .C2(n20681), .ZN(P2_U3224) );
  OAI222_X1 U23647 ( .A1(n20680), .A2(n10972), .B1(n20652), .B2(n20765), .C1(
        n10967), .C2(n20681), .ZN(P2_U3225) );
  OAI222_X1 U23648 ( .A1(n20680), .A2(n20654), .B1(n20653), .B2(n20765), .C1(
        n10972), .C2(n20681), .ZN(P2_U3226) );
  OAI222_X1 U23649 ( .A1(n20684), .A2(n20656), .B1(n20655), .B2(n20765), .C1(
        n20654), .C2(n20681), .ZN(P2_U3227) );
  OAI222_X1 U23650 ( .A1(n20684), .A2(n20658), .B1(n20657), .B2(n20765), .C1(
        n20656), .C2(n20681), .ZN(P2_U3228) );
  OAI222_X1 U23651 ( .A1(n20684), .A2(n20660), .B1(n20659), .B2(n20765), .C1(
        n20658), .C2(n20681), .ZN(P2_U3229) );
  OAI222_X1 U23652 ( .A1(n20684), .A2(n16124), .B1(n20661), .B2(n20765), .C1(
        n20660), .C2(n20681), .ZN(P2_U3230) );
  OAI222_X1 U23653 ( .A1(n20684), .A2(n20663), .B1(n20662), .B2(n20765), .C1(
        n16124), .C2(n20681), .ZN(P2_U3231) );
  OAI222_X1 U23654 ( .A1(n20684), .A2(n10995), .B1(n20664), .B2(n20765), .C1(
        n20663), .C2(n20681), .ZN(P2_U3232) );
  OAI222_X1 U23655 ( .A1(n20680), .A2(n20666), .B1(n20665), .B2(n20765), .C1(
        n10995), .C2(n20681), .ZN(P2_U3233) );
  OAI222_X1 U23656 ( .A1(n20680), .A2(n20668), .B1(n20667), .B2(n20765), .C1(
        n20666), .C2(n20681), .ZN(P2_U3234) );
  OAI222_X1 U23657 ( .A1(n20680), .A2(n20670), .B1(n20669), .B2(n20765), .C1(
        n20668), .C2(n20681), .ZN(P2_U3235) );
  OAI222_X1 U23658 ( .A1(n20680), .A2(n20672), .B1(n20671), .B2(n20765), .C1(
        n20670), .C2(n20681), .ZN(P2_U3236) );
  OAI222_X1 U23659 ( .A1(n20680), .A2(n20675), .B1(n20673), .B2(n20765), .C1(
        n20672), .C2(n20681), .ZN(P2_U3237) );
  OAI222_X1 U23660 ( .A1(n20681), .A2(n20675), .B1(n20674), .B2(n20765), .C1(
        n20676), .C2(n20680), .ZN(P2_U3238) );
  OAI222_X1 U23661 ( .A1(n20680), .A2(n20678), .B1(n20677), .B2(n20765), .C1(
        n20676), .C2(n20681), .ZN(P2_U3239) );
  OAI222_X1 U23662 ( .A1(n20680), .A2(n11022), .B1(n20679), .B2(n20765), .C1(
        n20678), .C2(n20681), .ZN(P2_U3240) );
  OAI222_X1 U23663 ( .A1(n20684), .A2(n20683), .B1(n20682), .B2(n20765), .C1(
        n11022), .C2(n20681), .ZN(P2_U3241) );
  INV_X1 U23664 ( .A(P2_BE_N_REG_3__SCAN_IN), .ZN(n20685) );
  AOI22_X1 U23665 ( .A1(n20765), .A2(n20686), .B1(n20685), .B2(n20762), .ZN(
        P2_U3585) );
  MUX2_X1 U23666 ( .A(P2_BE_N_REG_2__SCAN_IN), .B(P2_BYTEENABLE_REG_2__SCAN_IN), .S(n20765), .Z(P2_U3586) );
  INV_X1 U23667 ( .A(P2_BE_N_REG_1__SCAN_IN), .ZN(n20687) );
  AOI22_X1 U23668 ( .A1(n20765), .A2(n20688), .B1(n20687), .B2(n20762), .ZN(
        P2_U3587) );
  INV_X1 U23669 ( .A(P2_BE_N_REG_0__SCAN_IN), .ZN(n20689) );
  AOI22_X1 U23670 ( .A1(n20765), .A2(n20690), .B1(n20689), .B2(n20762), .ZN(
        P2_U3588) );
  OAI21_X1 U23671 ( .B1(n20694), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .A(n20692), 
        .ZN(n20691) );
  INV_X1 U23672 ( .A(n20691), .ZN(P2_U3591) );
  OAI21_X1 U23673 ( .B1(n20694), .B2(n20693), .A(n20692), .ZN(P2_U3592) );
  NAND2_X1 U23674 ( .A1(n20695), .A2(n20711), .ZN(n20704) );
  NAND3_X1 U23675 ( .A1(n20718), .A2(n20696), .A3(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n20697) );
  NAND2_X1 U23676 ( .A1(n20697), .A2(n20722), .ZN(n20705) );
  NAND2_X1 U23677 ( .A1(n20704), .A2(n20705), .ZN(n20702) );
  AOI222_X1 U23678 ( .A1(n20702), .A2(n20701), .B1(P2_STATE2_REG_3__SCAN_IN), 
        .B2(n20700), .C1(n20699), .C2(n20698), .ZN(n20703) );
  AOI22_X1 U23679 ( .A1(n20730), .A2(n10567), .B1(n20703), .B2(n20731), .ZN(
        P2_U3602) );
  OAI21_X1 U23680 ( .B1(n20706), .B2(n20705), .A(n20704), .ZN(n20707) );
  AOI21_X1 U23681 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n20708), .A(n20707), 
        .ZN(n20709) );
  AOI22_X1 U23682 ( .A1(n20730), .A2(n20710), .B1(n20709), .B2(n20731), .ZN(
        P2_U3603) );
  INV_X1 U23683 ( .A(n20711), .ZN(n20717) );
  NAND2_X1 U23684 ( .A1(n20712), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n20716) );
  INV_X1 U23685 ( .A(n20713), .ZN(n20714) );
  NAND3_X1 U23686 ( .A1(n20718), .A2(n20722), .A3(n20714), .ZN(n20715) );
  OAI211_X1 U23687 ( .C1(n20718), .C2(n20717), .A(n20716), .B(n20715), .ZN(
        n20719) );
  INV_X1 U23688 ( .A(n20719), .ZN(n20720) );
  AOI22_X1 U23689 ( .A1(n20730), .A2(n20721), .B1(n20720), .B2(n20731), .ZN(
        P2_U3604) );
  INV_X1 U23690 ( .A(n20722), .ZN(n20726) );
  INV_X1 U23691 ( .A(n20723), .ZN(n20725) );
  OAI22_X1 U23692 ( .A1(n20727), .A2(n20726), .B1(n20725), .B2(n20724), .ZN(
        n20728) );
  AOI21_X1 U23693 ( .B1(n20732), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n20728), 
        .ZN(n20729) );
  OAI22_X1 U23694 ( .A1(n20732), .A2(n20731), .B1(n20730), .B2(n20729), .ZN(
        P2_U3605) );
  INV_X1 U23695 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n20733) );
  AOI22_X1 U23696 ( .A1(n20765), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n20733), 
        .B2(n20762), .ZN(P2_U3608) );
  INV_X1 U23697 ( .A(n20734), .ZN(n20739) );
  NAND2_X1 U23698 ( .A1(n20736), .A2(n20735), .ZN(n20737) );
  OAI211_X1 U23699 ( .C1(n20740), .C2(n20739), .A(n20738), .B(n20737), .ZN(
        n20742) );
  MUX2_X1 U23700 ( .A(P2_MORE_REG_SCAN_IN), .B(n20742), .S(n20741), .Z(
        P2_U3609) );
  NOR2_X1 U23701 ( .A1(n20744), .A2(n20743), .ZN(n20746) );
  AOI211_X1 U23702 ( .C1(n20333), .C2(n20747), .A(n20746), .B(n20745), .ZN(
        n20760) );
  NAND2_X1 U23703 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n20748), .ZN(n20752) );
  NOR4_X1 U23704 ( .A1(n20756), .A2(n9759), .A3(n20750), .A4(n20749), .ZN(
        n20751) );
  AOI21_X1 U23705 ( .B1(n20753), .B2(n20752), .A(n20751), .ZN(n20759) );
  AOI211_X1 U23706 ( .C1(P2_STATEBS16_REG_SCAN_IN), .C2(n20756), .A(n20755), 
        .B(n20754), .ZN(n20757) );
  NOR2_X1 U23707 ( .A1(n20760), .A2(n20757), .ZN(n20758) );
  AOI22_X1 U23708 ( .A1(n20761), .A2(n20760), .B1(n20759), .B2(n20758), .ZN(
        P2_U3610) );
  INV_X1 U23709 ( .A(P2_M_IO_N_REG_SCAN_IN), .ZN(n20763) );
  AOI22_X1 U23710 ( .A1(n20765), .A2(n20764), .B1(n20763), .B2(n20762), .ZN(
        P2_U3611) );
  OAI21_X1 U23711 ( .B1(P1_STATE_REG_2__SCAN_IN), .B2(n21180), .A(
        P1_STATE_REG_0__SCAN_IN), .ZN(n21195) );
  OR2_X1 U23712 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n21180), .ZN(n21283) );
  OAI21_X1 U23713 ( .B1(n21195), .B2(P1_ADS_N_REG_SCAN_IN), .A(n21283), .ZN(
        n20766) );
  INV_X1 U23714 ( .A(n20766), .ZN(P1_U2802) );
  NAND2_X1 U23715 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n21270), .ZN(n20770) );
  OAI21_X1 U23716 ( .B1(n20768), .B2(n20767), .A(P1_CODEFETCH_REG_SCAN_IN), 
        .ZN(n20769) );
  OAI21_X1 U23717 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n20770), .A(n20769), 
        .ZN(P1_U2803) );
  NOR2_X1 U23718 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(P1_STATE_REG_0__SCAN_IN), 
        .ZN(n20772) );
  OAI21_X1 U23719 ( .B1(P1_D_C_N_REG_SCAN_IN), .B2(n20772), .A(n21283), .ZN(
        n20771) );
  OAI21_X1 U23720 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(n21283), .A(n20771), 
        .ZN(P1_U2804) );
  NAND2_X1 U23721 ( .A1(n21195), .A2(n21283), .ZN(n21263) );
  INV_X1 U23722 ( .A(n21263), .ZN(n21267) );
  OAI21_X1 U23723 ( .B1(BS16), .B2(n20772), .A(n21267), .ZN(n21265) );
  OAI21_X1 U23724 ( .B1(n21267), .B2(n21118), .A(n21265), .ZN(P1_U2805) );
  OAI21_X1 U23725 ( .B1(n20775), .B2(n20774), .A(n20773), .ZN(P1_U2806) );
  NOR4_X1 U23726 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_20__SCAN_IN), .A3(P1_DATAWIDTH_REG_21__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_22__SCAN_IN), .ZN(n20779) );
  NOR4_X1 U23727 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_16__SCAN_IN), .A3(P1_DATAWIDTH_REG_17__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_18__SCAN_IN), .ZN(n20778) );
  NOR4_X1 U23728 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_29__SCAN_IN), .A3(P1_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_31__SCAN_IN), .ZN(n20777) );
  NOR4_X1 U23729 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_24__SCAN_IN), .A3(P1_DATAWIDTH_REG_25__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_27__SCAN_IN), .ZN(n20776) );
  NAND4_X1 U23730 ( .A1(n20779), .A2(n20778), .A3(n20777), .A4(n20776), .ZN(
        n20785) );
  NOR4_X1 U23731 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_3__SCAN_IN), .A3(P1_DATAWIDTH_REG_4__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_5__SCAN_IN), .ZN(n20783) );
  AOI211_X1 U23732 ( .C1(P1_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_26__SCAN_IN), .B(
        P1_DATAWIDTH_REG_9__SCAN_IN), .ZN(n20782) );
  NOR4_X1 U23733 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_12__SCAN_IN), .A3(P1_DATAWIDTH_REG_13__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_14__SCAN_IN), .ZN(n20781) );
  NOR4_X1 U23734 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_7__SCAN_IN), .A3(P1_DATAWIDTH_REG_8__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_10__SCAN_IN), .ZN(n20780) );
  NAND4_X1 U23735 ( .A1(n20783), .A2(n20782), .A3(n20781), .A4(n20780), .ZN(
        n20784) );
  NOR2_X1 U23736 ( .A1(n20785), .A2(n20784), .ZN(n21282) );
  INV_X1 U23737 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n21260) );
  NOR3_X1 U23738 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A3(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n20787) );
  OAI21_X1 U23739 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n20787), .A(n21282), .ZN(
        n20786) );
  OAI21_X1 U23740 ( .B1(n21282), .B2(n21260), .A(n20786), .ZN(P1_U2807) );
  INV_X1 U23741 ( .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n21266) );
  AOI21_X1 U23742 ( .B1(n20846), .B2(n21266), .A(n20787), .ZN(n20788) );
  INV_X1 U23743 ( .A(n21282), .ZN(n21277) );
  AOI22_X1 U23744 ( .A1(n21282), .A2(n20788), .B1(n21257), .B2(n21277), .ZN(
        P1_U2808) );
  OAI21_X1 U23745 ( .B1(P1_REIP_REG_7__SCAN_IN), .B2(n20789), .A(n20816), .ZN(
        n20791) );
  NOR2_X1 U23746 ( .A1(n20818), .A2(n12147), .ZN(n20790) );
  AOI211_X1 U23747 ( .C1(P1_EBX_REG_7__SCAN_IN), .C2(n20850), .A(n20791), .B(
        n20790), .ZN(n20794) );
  OR2_X1 U23748 ( .A1(n20813), .A2(n20792), .ZN(n20804) );
  NAND2_X1 U23749 ( .A1(n20804), .A2(n20845), .ZN(n20800) );
  NAND2_X1 U23750 ( .A1(n20800), .A2(P1_REIP_REG_7__SCAN_IN), .ZN(n20793) );
  OAI211_X1 U23751 ( .C1(n20795), .C2(n20860), .A(n20794), .B(n20793), .ZN(
        n20796) );
  AOI21_X1 U23752 ( .B1(n20797), .B2(n20808), .A(n20796), .ZN(n20798) );
  OAI21_X1 U23753 ( .B1(n20799), .B2(n20847), .A(n20798), .ZN(P1_U2833) );
  AOI22_X1 U23754 ( .A1(n20800), .A2(P1_REIP_REG_6__SCAN_IN), .B1(n20850), 
        .B2(P1_EBX_REG_6__SCAN_IN), .ZN(n20801) );
  OAI21_X1 U23755 ( .B1(n20860), .B2(n20802), .A(n20801), .ZN(n20803) );
  AOI211_X1 U23756 ( .C1(n20849), .C2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n20831), .B(n20803), .ZN(n20811) );
  INV_X1 U23757 ( .A(n20804), .ZN(n20807) );
  AOI21_X1 U23758 ( .B1(n20857), .B2(n20827), .A(n20805), .ZN(n20830) );
  INV_X1 U23759 ( .A(n20830), .ZN(n20806) );
  NOR2_X1 U23760 ( .A1(n20806), .A2(n21205), .ZN(n20814) );
  AOI22_X1 U23761 ( .A1(n20809), .A2(n20808), .B1(n20807), .B2(n20814), .ZN(
        n20810) );
  OAI211_X1 U23762 ( .C1(n20812), .C2(n20847), .A(n20811), .B(n20810), .ZN(
        P1_U2834) );
  OR2_X1 U23763 ( .A1(n20813), .A2(n20827), .ZN(n20815) );
  AOI21_X1 U23764 ( .B1(n21205), .B2(n20815), .A(n20814), .ZN(n20823) );
  INV_X1 U23765 ( .A(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n20817) );
  OAI21_X1 U23766 ( .B1(n20818), .B2(n20817), .A(n20816), .ZN(n20819) );
  AOI21_X1 U23767 ( .B1(n20850), .B2(P1_EBX_REG_5__SCAN_IN), .A(n20819), .ZN(
        n20820) );
  OAI21_X1 U23768 ( .B1(n20821), .B2(n20860), .A(n20820), .ZN(n20822) );
  AOI211_X1 U23769 ( .C1(n20824), .C2(n20855), .A(n20823), .B(n20822), .ZN(
        n20825) );
  OAI21_X1 U23770 ( .B1(n20826), .B2(n20847), .A(n20825), .ZN(P1_U2835) );
  NAND2_X1 U23771 ( .A1(n20857), .A2(n20827), .ZN(n20829) );
  NAND3_X1 U23772 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_2__SCAN_IN), 
        .A3(P1_REIP_REG_3__SCAN_IN), .ZN(n20828) );
  OAI22_X1 U23773 ( .A1(n21202), .A2(n20830), .B1(n20829), .B2(n20828), .ZN(
        n20832) );
  AOI211_X1 U23774 ( .C1(n20849), .C2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n20832), .B(n20831), .ZN(n20834) );
  NAND2_X1 U23775 ( .A1(n20850), .A2(P1_EBX_REG_4__SCAN_IN), .ZN(n20833) );
  OAI211_X1 U23776 ( .C1(n20860), .C2(n20835), .A(n20834), .B(n20833), .ZN(
        n20836) );
  AOI21_X1 U23777 ( .B1(n20838), .B2(n20837), .A(n20836), .ZN(n20843) );
  INV_X1 U23778 ( .A(n20839), .ZN(n20840) );
  AOI22_X1 U23779 ( .A1(n20841), .A2(n20855), .B1(n20840), .B2(n16629), .ZN(
        n20842) );
  NAND2_X1 U23780 ( .A1(n20843), .A2(n20842), .ZN(P1_U2836) );
  INV_X1 U23781 ( .A(n20844), .ZN(n20856) );
  OAI22_X1 U23782 ( .A1(n20847), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B1(
        n20846), .B2(n20845), .ZN(n20848) );
  AOI21_X1 U23783 ( .B1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n20849), .A(
        n20848), .ZN(n20852) );
  NAND2_X1 U23784 ( .A1(n20850), .A2(P1_EBX_REG_1__SCAN_IN), .ZN(n20851) );
  OAI211_X1 U23785 ( .C1(n20853), .C2(n14001), .A(n20852), .B(n20851), .ZN(
        n20854) );
  AOI21_X1 U23786 ( .B1(n20856), .B2(n20855), .A(n20854), .ZN(n20859) );
  NAND2_X1 U23787 ( .A1(n20857), .A2(n20846), .ZN(n20858) );
  OAI211_X1 U23788 ( .C1(n20861), .C2(n20860), .A(n20859), .B(n20858), .ZN(
        P1_U2839) );
  INV_X1 U23789 ( .A(n20862), .ZN(n20866) );
  AOI22_X1 U23790 ( .A1(n20866), .A2(P1_EAX_REG_27__SCAN_IN), .B1(
        P1_UWORD_REG_11__SCAN_IN), .B2(n21288), .ZN(n20863) );
  OAI21_X1 U23791 ( .B1(n20865), .B2(n20864), .A(n20863), .ZN(P1_U2909) );
  AOI22_X1 U23792 ( .A1(n20866), .A2(P1_EAX_REG_22__SCAN_IN), .B1(
        P1_DATAO_REG_22__SCAN_IN), .B2(n20901), .ZN(n20867) );
  OAI21_X1 U23793 ( .B1(n20868), .B2(n20871), .A(n20867), .ZN(P1_U2914) );
  AOI22_X1 U23794 ( .A1(P1_EAX_REG_15__SCAN_IN), .A2(n20869), .B1(n20901), 
        .B2(P1_DATAO_REG_15__SCAN_IN), .ZN(n20870) );
  OAI21_X1 U23795 ( .B1(n20872), .B2(n20871), .A(n20870), .ZN(P1_U2921) );
  INV_X1 U23796 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n20874) );
  AOI22_X1 U23797 ( .A1(P1_LWORD_REG_14__SCAN_IN), .A2(n21288), .B1(n20901), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n20873) );
  OAI21_X1 U23798 ( .B1(n20874), .B2(n20903), .A(n20873), .ZN(P1_U2922) );
  INV_X1 U23799 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n20876) );
  AOI22_X1 U23800 ( .A1(P1_LWORD_REG_13__SCAN_IN), .A2(n21288), .B1(n20901), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n20875) );
  OAI21_X1 U23801 ( .B1(n20876), .B2(n20903), .A(n20875), .ZN(P1_U2923) );
  AOI22_X1 U23802 ( .A1(P1_LWORD_REG_12__SCAN_IN), .A2(n21288), .B1(n20894), 
        .B2(P1_DATAO_REG_12__SCAN_IN), .ZN(n20877) );
  OAI21_X1 U23803 ( .B1(n14687), .B2(n20903), .A(n20877), .ZN(P1_U2924) );
  AOI22_X1 U23804 ( .A1(P1_LWORD_REG_11__SCAN_IN), .A2(n21288), .B1(n20894), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n20878) );
  OAI21_X1 U23805 ( .B1(n20879), .B2(n20903), .A(n20878), .ZN(P1_U2925) );
  INV_X1 U23806 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n20881) );
  AOI22_X1 U23807 ( .A1(P1_LWORD_REG_10__SCAN_IN), .A2(n21288), .B1(n20894), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n20880) );
  OAI21_X1 U23808 ( .B1(n20881), .B2(n20903), .A(n20880), .ZN(P1_U2926) );
  INV_X1 U23809 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n20883) );
  AOI22_X1 U23810 ( .A1(P1_LWORD_REG_9__SCAN_IN), .A2(n21288), .B1(n20894), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n20882) );
  OAI21_X1 U23811 ( .B1(n20883), .B2(n20903), .A(n20882), .ZN(P1_U2927) );
  INV_X1 U23812 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n20885) );
  AOI22_X1 U23813 ( .A1(P1_LWORD_REG_8__SCAN_IN), .A2(n21288), .B1(n20894), 
        .B2(P1_DATAO_REG_8__SCAN_IN), .ZN(n20884) );
  OAI21_X1 U23814 ( .B1(n20885), .B2(n20903), .A(n20884), .ZN(P1_U2928) );
  AOI22_X1 U23815 ( .A1(P1_LWORD_REG_7__SCAN_IN), .A2(n21288), .B1(n20894), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n20886) );
  OAI21_X1 U23816 ( .B1(n20887), .B2(n20903), .A(n20886), .ZN(P1_U2929) );
  AOI22_X1 U23817 ( .A1(P1_LWORD_REG_6__SCAN_IN), .A2(n21288), .B1(n20894), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n20888) );
  OAI21_X1 U23818 ( .B1(n20889), .B2(n20903), .A(n20888), .ZN(P1_U2930) );
  AOI22_X1 U23819 ( .A1(P1_LWORD_REG_5__SCAN_IN), .A2(n21288), .B1(n20894), 
        .B2(P1_DATAO_REG_5__SCAN_IN), .ZN(n20890) );
  OAI21_X1 U23820 ( .B1(n20891), .B2(n20903), .A(n20890), .ZN(P1_U2931) );
  AOI22_X1 U23821 ( .A1(P1_LWORD_REG_4__SCAN_IN), .A2(n21288), .B1(n20894), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n20892) );
  OAI21_X1 U23822 ( .B1(n20893), .B2(n20903), .A(n20892), .ZN(P1_U2932) );
  AOI22_X1 U23823 ( .A1(P1_LWORD_REG_3__SCAN_IN), .A2(n21288), .B1(n20894), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n20895) );
  OAI21_X1 U23824 ( .B1(n20896), .B2(n20903), .A(n20895), .ZN(P1_U2933) );
  AOI22_X1 U23825 ( .A1(P1_LWORD_REG_2__SCAN_IN), .A2(n21288), .B1(n20901), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n20897) );
  OAI21_X1 U23826 ( .B1(n20898), .B2(n20903), .A(n20897), .ZN(P1_U2934) );
  AOI22_X1 U23827 ( .A1(P1_LWORD_REG_1__SCAN_IN), .A2(n21288), .B1(n20901), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n20899) );
  OAI21_X1 U23828 ( .B1(n20900), .B2(n20903), .A(n20899), .ZN(P1_U2935) );
  AOI22_X1 U23829 ( .A1(P1_LWORD_REG_0__SCAN_IN), .A2(n21288), .B1(n20901), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n20902) );
  OAI21_X1 U23830 ( .B1(n20904), .B2(n20903), .A(n20902), .ZN(P1_U2936) );
  AOI22_X1 U23831 ( .A1(n9717), .A2(P1_EAX_REG_24__SCAN_IN), .B1(
        P1_UWORD_REG_8__SCAN_IN), .B2(n20921), .ZN(n20906) );
  NAND2_X1 U23832 ( .A1(n13652), .A2(n20905), .ZN(n20911) );
  NAND2_X1 U23833 ( .A1(n20906), .A2(n20911), .ZN(P1_U2945) );
  AOI22_X1 U23834 ( .A1(n9717), .A2(P1_EAX_REG_26__SCAN_IN), .B1(
        P1_UWORD_REG_10__SCAN_IN), .B2(n20921), .ZN(n20908) );
  NAND2_X1 U23835 ( .A1(n13652), .A2(n20907), .ZN(n20915) );
  NAND2_X1 U23836 ( .A1(n20908), .A2(n20915), .ZN(P1_U2947) );
  AOI22_X1 U23837 ( .A1(n9717), .A2(P1_EAX_REG_28__SCAN_IN), .B1(
        P1_UWORD_REG_12__SCAN_IN), .B2(n20921), .ZN(n20910) );
  NAND2_X1 U23838 ( .A1(n13652), .A2(n20909), .ZN(n20917) );
  NAND2_X1 U23839 ( .A1(n20910), .A2(n20917), .ZN(P1_U2949) );
  AOI22_X1 U23840 ( .A1(n9717), .A2(P1_EAX_REG_8__SCAN_IN), .B1(
        P1_LWORD_REG_8__SCAN_IN), .B2(n20921), .ZN(n20912) );
  NAND2_X1 U23841 ( .A1(n20912), .A2(n20911), .ZN(P1_U2960) );
  AOI22_X1 U23842 ( .A1(n9717), .A2(P1_EAX_REG_9__SCAN_IN), .B1(
        P1_LWORD_REG_9__SCAN_IN), .B2(n20921), .ZN(n20914) );
  NAND2_X1 U23843 ( .A1(n20914), .A2(n20913), .ZN(P1_U2961) );
  AOI22_X1 U23844 ( .A1(n9717), .A2(P1_EAX_REG_10__SCAN_IN), .B1(
        P1_LWORD_REG_10__SCAN_IN), .B2(n20921), .ZN(n20916) );
  NAND2_X1 U23845 ( .A1(n20916), .A2(n20915), .ZN(P1_U2962) );
  AOI22_X1 U23846 ( .A1(n9717), .A2(P1_EAX_REG_12__SCAN_IN), .B1(
        P1_LWORD_REG_12__SCAN_IN), .B2(n20921), .ZN(n20918) );
  NAND2_X1 U23847 ( .A1(n20918), .A2(n20917), .ZN(P1_U2964) );
  AOI22_X1 U23848 ( .A1(n9717), .A2(P1_EAX_REG_13__SCAN_IN), .B1(
        P1_LWORD_REG_13__SCAN_IN), .B2(n20921), .ZN(n20920) );
  NAND2_X1 U23849 ( .A1(n20920), .A2(n20919), .ZN(P1_U2965) );
  AOI22_X1 U23850 ( .A1(n9717), .A2(P1_EAX_REG_14__SCAN_IN), .B1(
        P1_LWORD_REG_14__SCAN_IN), .B2(n20921), .ZN(n20923) );
  NAND2_X1 U23851 ( .A1(n20923), .A2(n20922), .ZN(P1_U2966) );
  NOR2_X1 U23852 ( .A1(n20925), .A2(n20924), .ZN(n20926) );
  AOI21_X1 U23853 ( .B1(n20928), .B2(n20927), .A(n20926), .ZN(n20937) );
  NAND2_X1 U23854 ( .A1(n20930), .A2(n20929), .ZN(n20933) );
  OAI22_X1 U23855 ( .A1(n20934), .A2(n20933), .B1(n20932), .B2(n20931), .ZN(
        n20935) );
  NAND3_X1 U23856 ( .A1(n20937), .A2(n20936), .A3(n20935), .ZN(P1_U3031) );
  NOR2_X1 U23857 ( .A1(n20939), .A2(n20938), .ZN(P1_U3032) );
  NAND3_X1 U23858 ( .A1(n21010), .A2(n20941), .A3(n21009), .ZN(n20980) );
  NOR2_X1 U23859 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20980), .ZN(
        n20973) );
  AOI22_X1 U23860 ( .A1(n20973), .A2(n21115), .B1(n20972), .B2(n21019), .ZN(
        n20959) );
  NOR2_X1 U23861 ( .A1(n20972), .A2(n21122), .ZN(n20944) );
  INV_X1 U23862 ( .A(n20942), .ZN(n20943) );
  AOI21_X1 U23863 ( .B1(n21005), .B2(n20944), .A(n20943), .ZN(n20957) );
  INV_X1 U23864 ( .A(n20957), .ZN(n20950) );
  OR2_X1 U23865 ( .A1(n20946), .A2(n20945), .ZN(n20956) );
  INV_X1 U23866 ( .A(n20947), .ZN(n20948) );
  NAND2_X1 U23867 ( .A1(n20949), .A2(n20948), .ZN(n21013) );
  AOI22_X1 U23868 ( .A1(n20950), .A2(n20956), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n21013), .ZN(n20951) );
  OAI211_X1 U23869 ( .C1(n20973), .C2(n20953), .A(n20952), .B(n20951), .ZN(
        n20975) );
  INV_X1 U23870 ( .A(n20954), .ZN(n20955) );
  OAI22_X1 U23871 ( .A1(n20957), .A2(n20956), .B1(n20955), .B2(n21013), .ZN(
        n20974) );
  AOI22_X1 U23872 ( .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n20975), .B1(
        n21114), .B2(n20974), .ZN(n20958) );
  OAI211_X1 U23873 ( .C1(n21022), .C2(n21005), .A(n20959), .B(n20958), .ZN(
        P1_U3033) );
  AOI22_X1 U23874 ( .A1(n20973), .A2(n21129), .B1(n20972), .B2(n21023), .ZN(
        n20961) );
  AOI22_X1 U23875 ( .A1(P1_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n20975), .B1(
        n21128), .B2(n20974), .ZN(n20960) );
  OAI211_X1 U23876 ( .C1(n21026), .C2(n21005), .A(n20961), .B(n20960), .ZN(
        P1_U3034) );
  AOI22_X1 U23877 ( .A1(n20973), .A2(n21135), .B1(n20972), .B2(n21027), .ZN(
        n20963) );
  AOI22_X1 U23878 ( .A1(P1_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n20975), .B1(
        n21134), .B2(n20974), .ZN(n20962) );
  OAI211_X1 U23879 ( .C1(n21030), .C2(n21005), .A(n20963), .B(n20962), .ZN(
        P1_U3035) );
  AOI22_X1 U23880 ( .A1(n20973), .A2(n21141), .B1(n20972), .B2(n21031), .ZN(
        n20965) );
  AOI22_X1 U23881 ( .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n20975), .B1(
        n21140), .B2(n20974), .ZN(n20964) );
  OAI211_X1 U23882 ( .C1(n21034), .C2(n21005), .A(n20965), .B(n20964), .ZN(
        P1_U3036) );
  AOI22_X1 U23883 ( .A1(n20973), .A2(n21147), .B1(n20972), .B2(n21035), .ZN(
        n20967) );
  AOI22_X1 U23884 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n20975), .B1(
        n21146), .B2(n20974), .ZN(n20966) );
  OAI211_X1 U23885 ( .C1(n21038), .C2(n21005), .A(n20967), .B(n20966), .ZN(
        P1_U3037) );
  AOI22_X1 U23886 ( .A1(n20973), .A2(n21153), .B1(n20972), .B2(n21039), .ZN(
        n20969) );
  AOI22_X1 U23887 ( .A1(P1_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n20975), .B1(
        n21152), .B2(n20974), .ZN(n20968) );
  OAI211_X1 U23888 ( .C1(n21042), .C2(n21005), .A(n20969), .B(n20968), .ZN(
        P1_U3038) );
  AOI22_X1 U23889 ( .A1(n20973), .A2(n21159), .B1(n20972), .B2(n21043), .ZN(
        n20971) );
  AOI22_X1 U23890 ( .A1(P1_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n20975), .B1(
        n21158), .B2(n20974), .ZN(n20970) );
  OAI211_X1 U23891 ( .C1(n21046), .C2(n21005), .A(n20971), .B(n20970), .ZN(
        P1_U3039) );
  AOI22_X1 U23892 ( .A1(n20973), .A2(n21167), .B1(n20972), .B2(n21049), .ZN(
        n20977) );
  AOI22_X1 U23893 ( .A1(P1_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n20975), .B1(
        n21165), .B2(n20974), .ZN(n20976) );
  OAI211_X1 U23894 ( .C1(n21054), .C2(n21005), .A(n20977), .B(n20976), .ZN(
        P1_U3040) );
  NOR2_X1 U23895 ( .A1(n21110), .A2(n20980), .ZN(n21000) );
  INV_X1 U23896 ( .A(n20978), .ZN(n21111) );
  AOI21_X1 U23897 ( .B1(n20979), .B2(n21111), .A(n21000), .ZN(n20981) );
  OAI22_X1 U23898 ( .A1(n20981), .A2(n21122), .B1(n20980), .B2(n21113), .ZN(
        n20999) );
  AOI22_X1 U23899 ( .A1(n21115), .A2(n21000), .B1(n21114), .B2(n20999), .ZN(
        n20986) );
  INV_X1 U23900 ( .A(n20980), .ZN(n20984) );
  OAI211_X1 U23901 ( .C1(n20982), .C2(n21118), .A(n21085), .B(n20981), .ZN(
        n20983) );
  OAI211_X1 U23902 ( .C1(n21085), .C2(n20984), .A(n21120), .B(n20983), .ZN(
        n21002) );
  AOI22_X1 U23903 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n21002), .B1(
        n21001), .B2(n21124), .ZN(n20985) );
  OAI211_X1 U23904 ( .C1(n21127), .C2(n21005), .A(n20986), .B(n20985), .ZN(
        P1_U3041) );
  AOI22_X1 U23905 ( .A1(n21129), .A2(n21000), .B1(n21128), .B2(n20999), .ZN(
        n20988) );
  AOI22_X1 U23906 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n21002), .B1(
        n21001), .B2(n21130), .ZN(n20987) );
  OAI211_X1 U23907 ( .C1(n21133), .C2(n21005), .A(n20988), .B(n20987), .ZN(
        P1_U3042) );
  AOI22_X1 U23908 ( .A1(n21135), .A2(n21000), .B1(n21134), .B2(n20999), .ZN(
        n20990) );
  AOI22_X1 U23909 ( .A1(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n21002), .B1(
        n21001), .B2(n21136), .ZN(n20989) );
  OAI211_X1 U23910 ( .C1(n21139), .C2(n21005), .A(n20990), .B(n20989), .ZN(
        P1_U3043) );
  AOI22_X1 U23911 ( .A1(n21141), .A2(n21000), .B1(n21140), .B2(n20999), .ZN(
        n20992) );
  AOI22_X1 U23912 ( .A1(P1_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n21002), .B1(
        n21001), .B2(n21142), .ZN(n20991) );
  OAI211_X1 U23913 ( .C1(n21145), .C2(n21005), .A(n20992), .B(n20991), .ZN(
        P1_U3044) );
  AOI22_X1 U23914 ( .A1(n21147), .A2(n21000), .B1(n21146), .B2(n20999), .ZN(
        n20994) );
  AOI22_X1 U23915 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n21002), .B1(
        n21001), .B2(n21148), .ZN(n20993) );
  OAI211_X1 U23916 ( .C1(n21151), .C2(n21005), .A(n20994), .B(n20993), .ZN(
        P1_U3045) );
  AOI22_X1 U23917 ( .A1(n21153), .A2(n21000), .B1(n21152), .B2(n20999), .ZN(
        n20996) );
  AOI22_X1 U23918 ( .A1(P1_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n21002), .B1(
        n21001), .B2(n21154), .ZN(n20995) );
  OAI211_X1 U23919 ( .C1(n21157), .C2(n21005), .A(n20996), .B(n20995), .ZN(
        P1_U3046) );
  AOI22_X1 U23920 ( .A1(n21159), .A2(n21000), .B1(n21158), .B2(n20999), .ZN(
        n20998) );
  AOI22_X1 U23921 ( .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n21002), .B1(
        n21001), .B2(n21160), .ZN(n20997) );
  OAI211_X1 U23922 ( .C1(n21163), .C2(n21005), .A(n20998), .B(n20997), .ZN(
        P1_U3047) );
  AOI22_X1 U23923 ( .A1(n21167), .A2(n21000), .B1(n21165), .B2(n20999), .ZN(
        n21004) );
  AOI22_X1 U23924 ( .A1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n21002), .B1(
        n21001), .B2(n21168), .ZN(n21003) );
  OAI211_X1 U23925 ( .C1(n21174), .C2(n21005), .A(n21004), .B(n21003), .ZN(
        P1_U3048) );
  INV_X1 U23926 ( .A(n21006), .ZN(n21007) );
  NAND3_X1 U23927 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n21010), .A3(
        n21009), .ZN(n21057) );
  NOR2_X1 U23928 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21057), .ZN(
        n21048) );
  NAND3_X1 U23929 ( .A1(n21055), .A2(n21085), .A3(n14001), .ZN(n21011) );
  OAI21_X1 U23930 ( .B1(n21013), .B2(n21012), .A(n21011), .ZN(n21047) );
  AOI22_X1 U23931 ( .A1(n21115), .A2(n21048), .B1(n21114), .B2(n21047), .ZN(
        n21021) );
  AOI21_X1 U23932 ( .B1(n21018), .B2(n21080), .A(n21118), .ZN(n21014) );
  AOI21_X1 U23933 ( .B1(n21055), .B2(n14001), .A(n21014), .ZN(n21015) );
  NOR2_X1 U23934 ( .A1(n21015), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n21017) );
  AOI22_X1 U23935 ( .A1(n21051), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n21050), .B2(n21019), .ZN(n21020) );
  OAI211_X1 U23936 ( .C1(n21022), .C2(n21080), .A(n21021), .B(n21020), .ZN(
        P1_U3065) );
  AOI22_X1 U23937 ( .A1(n21129), .A2(n21048), .B1(n21128), .B2(n21047), .ZN(
        n21025) );
  AOI22_X1 U23938 ( .A1(n21051), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n21050), .B2(n21023), .ZN(n21024) );
  OAI211_X1 U23939 ( .C1(n21026), .C2(n21080), .A(n21025), .B(n21024), .ZN(
        P1_U3066) );
  AOI22_X1 U23940 ( .A1(n21135), .A2(n21048), .B1(n21134), .B2(n21047), .ZN(
        n21029) );
  AOI22_X1 U23941 ( .A1(n21051), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n21050), .B2(n21027), .ZN(n21028) );
  OAI211_X1 U23942 ( .C1(n21030), .C2(n21080), .A(n21029), .B(n21028), .ZN(
        P1_U3067) );
  AOI22_X1 U23943 ( .A1(n21141), .A2(n21048), .B1(n21140), .B2(n21047), .ZN(
        n21033) );
  AOI22_X1 U23944 ( .A1(n21051), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n21050), .B2(n21031), .ZN(n21032) );
  OAI211_X1 U23945 ( .C1(n21034), .C2(n21080), .A(n21033), .B(n21032), .ZN(
        P1_U3068) );
  AOI22_X1 U23946 ( .A1(n21147), .A2(n21048), .B1(n21146), .B2(n21047), .ZN(
        n21037) );
  AOI22_X1 U23947 ( .A1(n21051), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n21050), .B2(n21035), .ZN(n21036) );
  OAI211_X1 U23948 ( .C1(n21038), .C2(n21080), .A(n21037), .B(n21036), .ZN(
        P1_U3069) );
  AOI22_X1 U23949 ( .A1(n21153), .A2(n21048), .B1(n21152), .B2(n21047), .ZN(
        n21041) );
  AOI22_X1 U23950 ( .A1(n21051), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n21050), .B2(n21039), .ZN(n21040) );
  OAI211_X1 U23951 ( .C1(n21042), .C2(n21080), .A(n21041), .B(n21040), .ZN(
        P1_U3070) );
  AOI22_X1 U23952 ( .A1(n21159), .A2(n21048), .B1(n21158), .B2(n21047), .ZN(
        n21045) );
  AOI22_X1 U23953 ( .A1(n21051), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n21050), .B2(n21043), .ZN(n21044) );
  OAI211_X1 U23954 ( .C1(n21046), .C2(n21080), .A(n21045), .B(n21044), .ZN(
        P1_U3071) );
  AOI22_X1 U23955 ( .A1(n21167), .A2(n21048), .B1(n21165), .B2(n21047), .ZN(
        n21053) );
  AOI22_X1 U23956 ( .A1(n21051), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n21050), .B2(n21049), .ZN(n21052) );
  OAI211_X1 U23957 ( .C1(n21054), .C2(n21080), .A(n21053), .B(n21052), .ZN(
        P1_U3072) );
  NOR2_X1 U23958 ( .A1(n21110), .A2(n21057), .ZN(n21075) );
  AOI21_X1 U23959 ( .B1(n21055), .B2(n21111), .A(n21075), .ZN(n21056) );
  OAI22_X1 U23960 ( .A1(n21056), .A2(n21122), .B1(n21057), .B2(n21113), .ZN(
        n21074) );
  AOI22_X1 U23961 ( .A1(n21115), .A2(n21075), .B1(n21114), .B2(n21074), .ZN(
        n21061) );
  INV_X1 U23962 ( .A(n21057), .ZN(n21059) );
  OAI21_X1 U23963 ( .B1(n21059), .B2(n21058), .A(n21120), .ZN(n21077) );
  AOI22_X1 U23964 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n21077), .B1(
        n21076), .B2(n21124), .ZN(n21060) );
  OAI211_X1 U23965 ( .C1(n21127), .C2(n21080), .A(n21061), .B(n21060), .ZN(
        P1_U3073) );
  AOI22_X1 U23966 ( .A1(n21129), .A2(n21075), .B1(n21128), .B2(n21074), .ZN(
        n21063) );
  AOI22_X1 U23967 ( .A1(P1_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n21077), .B1(
        n21076), .B2(n21130), .ZN(n21062) );
  OAI211_X1 U23968 ( .C1(n21133), .C2(n21080), .A(n21063), .B(n21062), .ZN(
        P1_U3074) );
  AOI22_X1 U23969 ( .A1(n21135), .A2(n21075), .B1(n21134), .B2(n21074), .ZN(
        n21065) );
  AOI22_X1 U23970 ( .A1(P1_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n21077), .B1(
        n21076), .B2(n21136), .ZN(n21064) );
  OAI211_X1 U23971 ( .C1(n21139), .C2(n21080), .A(n21065), .B(n21064), .ZN(
        P1_U3075) );
  AOI22_X1 U23972 ( .A1(n21141), .A2(n21075), .B1(n21140), .B2(n21074), .ZN(
        n21067) );
  AOI22_X1 U23973 ( .A1(P1_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n21077), .B1(
        n21076), .B2(n21142), .ZN(n21066) );
  OAI211_X1 U23974 ( .C1(n21145), .C2(n21080), .A(n21067), .B(n21066), .ZN(
        P1_U3076) );
  AOI22_X1 U23975 ( .A1(n21147), .A2(n21075), .B1(n21146), .B2(n21074), .ZN(
        n21069) );
  AOI22_X1 U23976 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n21077), .B1(
        n21076), .B2(n21148), .ZN(n21068) );
  OAI211_X1 U23977 ( .C1(n21151), .C2(n21080), .A(n21069), .B(n21068), .ZN(
        P1_U3077) );
  AOI22_X1 U23978 ( .A1(n21153), .A2(n21075), .B1(n21152), .B2(n21074), .ZN(
        n21071) );
  AOI22_X1 U23979 ( .A1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n21077), .B1(
        n21076), .B2(n21154), .ZN(n21070) );
  OAI211_X1 U23980 ( .C1(n21157), .C2(n21080), .A(n21071), .B(n21070), .ZN(
        P1_U3078) );
  AOI22_X1 U23981 ( .A1(n21159), .A2(n21075), .B1(n21158), .B2(n21074), .ZN(
        n21073) );
  AOI22_X1 U23982 ( .A1(P1_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n21077), .B1(
        n21076), .B2(n21160), .ZN(n21072) );
  OAI211_X1 U23983 ( .C1(n21163), .C2(n21080), .A(n21073), .B(n21072), .ZN(
        P1_U3079) );
  AOI22_X1 U23984 ( .A1(n21167), .A2(n21075), .B1(n21165), .B2(n21074), .ZN(
        n21079) );
  AOI22_X1 U23985 ( .A1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n21077), .B1(
        n21076), .B2(n21168), .ZN(n21078) );
  OAI211_X1 U23986 ( .C1(n21174), .C2(n21080), .A(n21079), .B(n21078), .ZN(
        P1_U3080) );
  NOR2_X1 U23987 ( .A1(n21110), .A2(n21083), .ZN(n21104) );
  INV_X1 U23988 ( .A(n21081), .ZN(n21082) );
  AOI21_X1 U23989 ( .B1(n21082), .B2(n21111), .A(n21104), .ZN(n21084) );
  OAI22_X1 U23990 ( .A1(n21084), .A2(n21122), .B1(n21083), .B2(n21113), .ZN(
        n21103) );
  AOI22_X1 U23991 ( .A1(n21115), .A2(n21104), .B1(n21114), .B2(n21103), .ZN(
        n21090) );
  INV_X1 U23992 ( .A(n21083), .ZN(n21088) );
  OAI211_X1 U23993 ( .C1(n21086), .C2(n21118), .A(n21085), .B(n21084), .ZN(
        n21087) );
  OAI211_X1 U23994 ( .C1(n21085), .C2(n21088), .A(n21120), .B(n21087), .ZN(
        n21106) );
  AOI22_X1 U23995 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n21106), .B1(
        n21105), .B2(n21124), .ZN(n21089) );
  OAI211_X1 U23996 ( .C1(n21127), .C2(n21109), .A(n21090), .B(n21089), .ZN(
        P1_U3105) );
  AOI22_X1 U23997 ( .A1(n21129), .A2(n21104), .B1(n21128), .B2(n21103), .ZN(
        n21092) );
  AOI22_X1 U23998 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n21106), .B1(
        n21105), .B2(n21130), .ZN(n21091) );
  OAI211_X1 U23999 ( .C1(n21133), .C2(n21109), .A(n21092), .B(n21091), .ZN(
        P1_U3106) );
  AOI22_X1 U24000 ( .A1(n21135), .A2(n21104), .B1(n21134), .B2(n21103), .ZN(
        n21094) );
  AOI22_X1 U24001 ( .A1(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n21106), .B1(
        n21105), .B2(n21136), .ZN(n21093) );
  OAI211_X1 U24002 ( .C1(n21139), .C2(n21109), .A(n21094), .B(n21093), .ZN(
        P1_U3107) );
  AOI22_X1 U24003 ( .A1(n21141), .A2(n21104), .B1(n21140), .B2(n21103), .ZN(
        n21096) );
  AOI22_X1 U24004 ( .A1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n21106), .B1(
        n21105), .B2(n21142), .ZN(n21095) );
  OAI211_X1 U24005 ( .C1(n21145), .C2(n21109), .A(n21096), .B(n21095), .ZN(
        P1_U3108) );
  AOI22_X1 U24006 ( .A1(n21147), .A2(n21104), .B1(n21146), .B2(n21103), .ZN(
        n21098) );
  AOI22_X1 U24007 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n21106), .B1(
        n21105), .B2(n21148), .ZN(n21097) );
  OAI211_X1 U24008 ( .C1(n21151), .C2(n21109), .A(n21098), .B(n21097), .ZN(
        P1_U3109) );
  AOI22_X1 U24009 ( .A1(n21153), .A2(n21104), .B1(n21152), .B2(n21103), .ZN(
        n21100) );
  AOI22_X1 U24010 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n21106), .B1(
        n21105), .B2(n21154), .ZN(n21099) );
  OAI211_X1 U24011 ( .C1(n21157), .C2(n21109), .A(n21100), .B(n21099), .ZN(
        P1_U3110) );
  AOI22_X1 U24012 ( .A1(n21159), .A2(n21104), .B1(n21158), .B2(n21103), .ZN(
        n21102) );
  AOI22_X1 U24013 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n21106), .B1(
        n21105), .B2(n21160), .ZN(n21101) );
  OAI211_X1 U24014 ( .C1(n21163), .C2(n21109), .A(n21102), .B(n21101), .ZN(
        P1_U3111) );
  AOI22_X1 U24015 ( .A1(n21167), .A2(n21104), .B1(n21165), .B2(n21103), .ZN(
        n21108) );
  AOI22_X1 U24016 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n21106), .B1(
        n21105), .B2(n21168), .ZN(n21107) );
  OAI211_X1 U24017 ( .C1(n21174), .C2(n21109), .A(n21108), .B(n21107), .ZN(
        P1_U3112) );
  NOR2_X1 U24018 ( .A1(n21110), .A2(n21116), .ZN(n21166) );
  AOI21_X1 U24019 ( .B1(n21112), .B2(n21111), .A(n21166), .ZN(n21117) );
  OAI22_X1 U24020 ( .A1(n21117), .A2(n21122), .B1(n21116), .B2(n21113), .ZN(
        n21164) );
  AOI22_X1 U24021 ( .A1(n21115), .A2(n21166), .B1(n21114), .B2(n21164), .ZN(
        n21126) );
  INV_X1 U24022 ( .A(n21116), .ZN(n21123) );
  OAI21_X1 U24023 ( .B1(n21119), .B2(n21118), .A(n21117), .ZN(n21121) );
  OAI221_X1 U24024 ( .B1(n21085), .B2(n21123), .C1(n21122), .C2(n21121), .A(
        n21120), .ZN(n21170) );
  AOI22_X1 U24025 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n21170), .B1(
        n21169), .B2(n21124), .ZN(n21125) );
  OAI211_X1 U24026 ( .C1(n21127), .C2(n21173), .A(n21126), .B(n21125), .ZN(
        P1_U3137) );
  AOI22_X1 U24027 ( .A1(n21129), .A2(n21166), .B1(n21128), .B2(n21164), .ZN(
        n21132) );
  AOI22_X1 U24028 ( .A1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n21170), .B1(
        n21169), .B2(n21130), .ZN(n21131) );
  OAI211_X1 U24029 ( .C1(n21133), .C2(n21173), .A(n21132), .B(n21131), .ZN(
        P1_U3138) );
  AOI22_X1 U24030 ( .A1(n21135), .A2(n21166), .B1(n21134), .B2(n21164), .ZN(
        n21138) );
  AOI22_X1 U24031 ( .A1(P1_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n21170), .B1(
        n21169), .B2(n21136), .ZN(n21137) );
  OAI211_X1 U24032 ( .C1(n21139), .C2(n21173), .A(n21138), .B(n21137), .ZN(
        P1_U3139) );
  AOI22_X1 U24033 ( .A1(n21141), .A2(n21166), .B1(n21140), .B2(n21164), .ZN(
        n21144) );
  AOI22_X1 U24034 ( .A1(P1_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n21170), .B1(
        n21169), .B2(n21142), .ZN(n21143) );
  OAI211_X1 U24035 ( .C1(n21145), .C2(n21173), .A(n21144), .B(n21143), .ZN(
        P1_U3140) );
  AOI22_X1 U24036 ( .A1(n21147), .A2(n21166), .B1(n21146), .B2(n21164), .ZN(
        n21150) );
  AOI22_X1 U24037 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n21170), .B1(
        n21169), .B2(n21148), .ZN(n21149) );
  OAI211_X1 U24038 ( .C1(n21151), .C2(n21173), .A(n21150), .B(n21149), .ZN(
        P1_U3141) );
  AOI22_X1 U24039 ( .A1(n21153), .A2(n21166), .B1(n21152), .B2(n21164), .ZN(
        n21156) );
  AOI22_X1 U24040 ( .A1(P1_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n21170), .B1(
        n21169), .B2(n21154), .ZN(n21155) );
  OAI211_X1 U24041 ( .C1(n21157), .C2(n21173), .A(n21156), .B(n21155), .ZN(
        P1_U3142) );
  AOI22_X1 U24042 ( .A1(n21159), .A2(n21166), .B1(n21158), .B2(n21164), .ZN(
        n21162) );
  AOI22_X1 U24043 ( .A1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n21170), .B1(
        n21169), .B2(n21160), .ZN(n21161) );
  OAI211_X1 U24044 ( .C1(n21163), .C2(n21173), .A(n21162), .B(n21161), .ZN(
        P1_U3143) );
  AOI22_X1 U24045 ( .A1(n21167), .A2(n21166), .B1(n21165), .B2(n21164), .ZN(
        n21172) );
  AOI22_X1 U24046 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n21170), .B1(
        n21169), .B2(n21168), .ZN(n21171) );
  OAI211_X1 U24047 ( .C1(n21174), .C2(n21173), .A(n21172), .B(n21171), .ZN(
        P1_U3144) );
  OR2_X1 U24048 ( .A1(n21176), .A2(n21175), .ZN(P1_U3163) );
  AND2_X1 U24049 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n21263), .ZN(
        P1_U3164) );
  AND2_X1 U24050 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n21263), .ZN(
        P1_U3165) );
  AND2_X1 U24051 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n21263), .ZN(
        P1_U3166) );
  AND2_X1 U24052 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n21263), .ZN(
        P1_U3167) );
  AND2_X1 U24053 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n21263), .ZN(
        P1_U3168) );
  NOR2_X1 U24054 ( .A1(n21267), .A2(n21177), .ZN(P1_U3169) );
  AND2_X1 U24055 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n21263), .ZN(
        P1_U3170) );
  AND2_X1 U24056 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n21263), .ZN(
        P1_U3171) );
  AND2_X1 U24057 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n21263), .ZN(
        P1_U3172) );
  AND2_X1 U24058 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n21263), .ZN(
        P1_U3173) );
  AND2_X1 U24059 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n21263), .ZN(
        P1_U3174) );
  AND2_X1 U24060 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n21263), .ZN(
        P1_U3175) );
  AND2_X1 U24061 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n21263), .ZN(
        P1_U3176) );
  AND2_X1 U24062 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n21263), .ZN(
        P1_U3177) );
  AND2_X1 U24063 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n21263), .ZN(
        P1_U3178) );
  AND2_X1 U24064 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n21263), .ZN(
        P1_U3179) );
  AND2_X1 U24065 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n21263), .ZN(
        P1_U3180) );
  AND2_X1 U24066 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n21263), .ZN(
        P1_U3181) );
  AND2_X1 U24067 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n21263), .ZN(
        P1_U3182) );
  AND2_X1 U24068 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n21263), .ZN(
        P1_U3183) );
  AND2_X1 U24069 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(n21263), .ZN(
        P1_U3184) );
  AND2_X1 U24070 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n21263), .ZN(
        P1_U3185) );
  NOR2_X1 U24071 ( .A1(n21267), .A2(n21178), .ZN(P1_U3186) );
  AND2_X1 U24072 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n21263), .ZN(P1_U3187) );
  AND2_X1 U24073 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n21263), .ZN(P1_U3188) );
  AND2_X1 U24074 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n21263), .ZN(P1_U3189) );
  AND2_X1 U24075 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n21263), .ZN(P1_U3190) );
  AND2_X1 U24076 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n21263), .ZN(P1_U3191) );
  AND2_X1 U24077 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n21263), .ZN(P1_U3192) );
  AND2_X1 U24078 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n21263), .ZN(P1_U3193) );
  NAND2_X1 U24079 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n21179), .ZN(n21191) );
  INV_X1 U24080 ( .A(n21191), .ZN(n21184) );
  INV_X2 U24081 ( .A(n21283), .ZN(n21296) );
  NAND2_X1 U24082 ( .A1(n21180), .A2(n21197), .ZN(n21182) );
  NAND2_X1 U24083 ( .A1(n21192), .A2(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n21185) );
  AOI22_X1 U24084 ( .A1(HOLD), .A2(n21182), .B1(n21185), .B2(n21181), .ZN(
        n21183) );
  OAI22_X1 U24085 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n21184), .B1(n21296), 
        .B2(n21183), .ZN(P1_U3194) );
  INV_X1 U24086 ( .A(n21185), .ZN(n21188) );
  AOI21_X1 U24087 ( .B1(P1_REQUESTPENDING_REG_SCAN_IN), .B2(n21197), .A(n21186), .ZN(n21187) );
  AOI21_X1 U24088 ( .B1(n21189), .B2(n21188), .A(n21187), .ZN(n21196) );
  NAND3_X1 U24089 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n21190), .A3(n21192), 
        .ZN(n21194) );
  OAI211_X1 U24090 ( .C1(P1_STATE_REG_1__SCAN_IN), .C2(n21192), .A(
        P1_STATE_REG_2__SCAN_IN), .B(n21191), .ZN(n21193) );
  OAI221_X1 U24091 ( .B1(n21196), .B2(n21195), .C1(n21196), .C2(n21194), .A(
        n21193), .ZN(P1_U3196) );
  NAND2_X1 U24092 ( .A1(n21296), .A2(n21197), .ZN(n21254) );
  INV_X1 U24093 ( .A(n21254), .ZN(n21248) );
  NAND2_X1 U24094 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n21296), .ZN(n21250) );
  INV_X1 U24095 ( .A(n21250), .ZN(n21252) );
  AOI222_X1 U24096 ( .A1(n21248), .A2(P1_REIP_REG_2__SCAN_IN), .B1(
        P1_ADDRESS_REG_0__SCAN_IN), .B2(n21283), .C1(P1_REIP_REG_1__SCAN_IN), 
        .C2(n21252), .ZN(n21198) );
  INV_X1 U24097 ( .A(n21198), .ZN(P1_U3197) );
  AOI222_X1 U24098 ( .A1(n21248), .A2(P1_REIP_REG_3__SCAN_IN), .B1(
        P1_ADDRESS_REG_1__SCAN_IN), .B2(n21283), .C1(P1_REIP_REG_2__SCAN_IN), 
        .C2(n21252), .ZN(n21199) );
  INV_X1 U24099 ( .A(n21199), .ZN(P1_U3198) );
  INV_X1 U24100 ( .A(P1_ADDRESS_REG_2__SCAN_IN), .ZN(n21201) );
  OAI222_X1 U24101 ( .A1(n21254), .A2(n21202), .B1(n21201), .B2(n21296), .C1(
        n21200), .C2(n21250), .ZN(P1_U3199) );
  INV_X1 U24102 ( .A(P1_ADDRESS_REG_3__SCAN_IN), .ZN(n21203) );
  OAI222_X1 U24103 ( .A1(n21254), .A2(n21205), .B1(n21203), .B2(n21296), .C1(
        n21202), .C2(n21250), .ZN(P1_U3200) );
  INV_X1 U24104 ( .A(P1_ADDRESS_REG_4__SCAN_IN), .ZN(n21204) );
  OAI222_X1 U24105 ( .A1(n21250), .A2(n21205), .B1(n21204), .B2(n21296), .C1(
        n21206), .C2(n21254), .ZN(P1_U3201) );
  OAI222_X1 U24106 ( .A1(n21254), .A2(n21208), .B1(n21207), .B2(n21296), .C1(
        n21206), .C2(n21250), .ZN(P1_U3202) );
  INV_X1 U24107 ( .A(P1_ADDRESS_REG_6__SCAN_IN), .ZN(n21209) );
  OAI222_X1 U24108 ( .A1(n21254), .A2(n21210), .B1(n21209), .B2(n21296), .C1(
        n21208), .C2(n21250), .ZN(P1_U3203) );
  INV_X1 U24109 ( .A(P1_ADDRESS_REG_7__SCAN_IN), .ZN(n21211) );
  OAI222_X1 U24110 ( .A1(n21254), .A2(n21213), .B1(n21211), .B2(n21296), .C1(
        n21210), .C2(n21250), .ZN(P1_U3204) );
  OAI222_X1 U24111 ( .A1(n21250), .A2(n21213), .B1(n21212), .B2(n21296), .C1(
        n21215), .C2(n21254), .ZN(P1_U3205) );
  AOI22_X1 U24112 ( .A1(P1_ADDRESS_REG_9__SCAN_IN), .A2(n21283), .B1(
        P1_REIP_REG_11__SCAN_IN), .B2(n21248), .ZN(n21214) );
  OAI21_X1 U24113 ( .B1(n21215), .B2(n21250), .A(n21214), .ZN(P1_U3206) );
  AOI22_X1 U24114 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(n21283), .B1(
        P1_REIP_REG_11__SCAN_IN), .B2(n21252), .ZN(n21216) );
  OAI21_X1 U24115 ( .B1(n21217), .B2(n21254), .A(n21216), .ZN(P1_U3207) );
  INV_X1 U24116 ( .A(P1_ADDRESS_REG_11__SCAN_IN), .ZN(n21218) );
  OAI222_X1 U24117 ( .A1(n21254), .A2(n21219), .B1(n21218), .B2(n21296), .C1(
        n21217), .C2(n21250), .ZN(P1_U3208) );
  INV_X1 U24118 ( .A(P1_ADDRESS_REG_12__SCAN_IN), .ZN(n21220) );
  OAI222_X1 U24119 ( .A1(n21254), .A2(n21222), .B1(n21220), .B2(n21296), .C1(
        n21219), .C2(n21250), .ZN(P1_U3209) );
  AOI22_X1 U24120 ( .A1(P1_ADDRESS_REG_13__SCAN_IN), .A2(n21283), .B1(
        P1_REIP_REG_15__SCAN_IN), .B2(n21248), .ZN(n21221) );
  OAI21_X1 U24121 ( .B1(n21222), .B2(n21250), .A(n21221), .ZN(P1_U3210) );
  INV_X1 U24122 ( .A(P1_REIP_REG_16__SCAN_IN), .ZN(n21225) );
  AOI22_X1 U24123 ( .A1(P1_ADDRESS_REG_14__SCAN_IN), .A2(n21283), .B1(
        P1_REIP_REG_15__SCAN_IN), .B2(n21252), .ZN(n21223) );
  OAI21_X1 U24124 ( .B1(n21225), .B2(n21254), .A(n21223), .ZN(P1_U3211) );
  INV_X1 U24125 ( .A(P1_ADDRESS_REG_15__SCAN_IN), .ZN(n21224) );
  OAI222_X1 U24126 ( .A1(n21250), .A2(n21225), .B1(n21224), .B2(n21296), .C1(
        n21227), .C2(n21254), .ZN(P1_U3212) );
  AOI22_X1 U24127 ( .A1(P1_ADDRESS_REG_16__SCAN_IN), .A2(n21283), .B1(
        P1_REIP_REG_18__SCAN_IN), .B2(n21248), .ZN(n21226) );
  OAI21_X1 U24128 ( .B1(n21227), .B2(n21250), .A(n21226), .ZN(P1_U3213) );
  AOI22_X1 U24129 ( .A1(P1_ADDRESS_REG_17__SCAN_IN), .A2(n21283), .B1(
        P1_REIP_REG_18__SCAN_IN), .B2(n21252), .ZN(n21228) );
  OAI21_X1 U24130 ( .B1(n21229), .B2(n21254), .A(n21228), .ZN(P1_U3214) );
  INV_X1 U24131 ( .A(P1_ADDRESS_REG_18__SCAN_IN), .ZN(n21230) );
  OAI222_X1 U24132 ( .A1(n21254), .A2(n21232), .B1(n21230), .B2(n21296), .C1(
        n21229), .C2(n21250), .ZN(P1_U3215) );
  INV_X1 U24133 ( .A(P1_ADDRESS_REG_19__SCAN_IN), .ZN(n21231) );
  OAI222_X1 U24134 ( .A1(n21250), .A2(n21232), .B1(n21231), .B2(n21296), .C1(
        n21234), .C2(n21254), .ZN(P1_U3216) );
  INV_X1 U24135 ( .A(P1_ADDRESS_REG_20__SCAN_IN), .ZN(n21233) );
  OAI222_X1 U24136 ( .A1(n21250), .A2(n21234), .B1(n21233), .B2(n21296), .C1(
        n21236), .C2(n21254), .ZN(P1_U3217) );
  AOI22_X1 U24137 ( .A1(P1_ADDRESS_REG_21__SCAN_IN), .A2(n21283), .B1(
        P1_REIP_REG_23__SCAN_IN), .B2(n21248), .ZN(n21235) );
  OAI21_X1 U24138 ( .B1(n21236), .B2(n21250), .A(n21235), .ZN(P1_U3218) );
  AOI22_X1 U24139 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(n21283), .B1(
        P1_REIP_REG_23__SCAN_IN), .B2(n21252), .ZN(n21237) );
  OAI21_X1 U24140 ( .B1(n21239), .B2(n21254), .A(n21237), .ZN(P1_U3219) );
  AOI22_X1 U24141 ( .A1(P1_ADDRESS_REG_23__SCAN_IN), .A2(n21283), .B1(
        P1_REIP_REG_25__SCAN_IN), .B2(n21248), .ZN(n21238) );
  OAI21_X1 U24142 ( .B1(n21239), .B2(n21250), .A(n21238), .ZN(P1_U3220) );
  OAI222_X1 U24143 ( .A1(n21250), .A2(n21241), .B1(n21240), .B2(n21296), .C1(
        n21242), .C2(n21254), .ZN(P1_U3221) );
  INV_X1 U24144 ( .A(P1_ADDRESS_REG_25__SCAN_IN), .ZN(n21243) );
  OAI222_X1 U24145 ( .A1(n21254), .A2(n21245), .B1(n21243), .B2(n21296), .C1(
        n21242), .C2(n21250), .ZN(P1_U3222) );
  INV_X1 U24146 ( .A(P1_ADDRESS_REG_26__SCAN_IN), .ZN(n21244) );
  OAI222_X1 U24147 ( .A1(n21250), .A2(n21245), .B1(n21244), .B2(n21296), .C1(
        n21247), .C2(n21254), .ZN(P1_U3223) );
  INV_X1 U24148 ( .A(P1_ADDRESS_REG_27__SCAN_IN), .ZN(n21246) );
  OAI222_X1 U24149 ( .A1(n21250), .A2(n21247), .B1(n21246), .B2(n21296), .C1(
        n21251), .C2(n21254), .ZN(P1_U3224) );
  AOI22_X1 U24150 ( .A1(P1_ADDRESS_REG_28__SCAN_IN), .A2(n21283), .B1(
        P1_REIP_REG_30__SCAN_IN), .B2(n21248), .ZN(n21249) );
  OAI21_X1 U24151 ( .B1(n21251), .B2(n21250), .A(n21249), .ZN(P1_U3225) );
  AOI22_X1 U24152 ( .A1(P1_ADDRESS_REG_29__SCAN_IN), .A2(n21283), .B1(
        P1_REIP_REG_30__SCAN_IN), .B2(n21252), .ZN(n21253) );
  OAI21_X1 U24153 ( .B1(n21255), .B2(n21254), .A(n21253), .ZN(P1_U3226) );
  AOI22_X1 U24154 ( .A1(n21296), .A2(n21257), .B1(n21256), .B2(n21283), .ZN(
        P1_U3458) );
  INV_X1 U24155 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n21278) );
  INV_X1 U24156 ( .A(P1_BE_N_REG_2__SCAN_IN), .ZN(n21258) );
  AOI22_X1 U24157 ( .A1(n21296), .A2(n21278), .B1(n21258), .B2(n21283), .ZN(
        P1_U3459) );
  INV_X1 U24158 ( .A(P1_BE_N_REG_1__SCAN_IN), .ZN(n21259) );
  AOI22_X1 U24159 ( .A1(n21296), .A2(n21260), .B1(n21259), .B2(n21283), .ZN(
        P1_U3460) );
  INV_X1 U24160 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n21281) );
  INV_X1 U24161 ( .A(P1_BE_N_REG_0__SCAN_IN), .ZN(n21261) );
  AOI22_X1 U24162 ( .A1(n21296), .A2(n21281), .B1(n21261), .B2(n21283), .ZN(
        P1_U3461) );
  INV_X1 U24163 ( .A(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(n21264) );
  INV_X1 U24164 ( .A(n21265), .ZN(n21262) );
  AOI21_X1 U24165 ( .B1(n21264), .B2(n21263), .A(n21262), .ZN(P1_U3464) );
  OAI21_X1 U24166 ( .B1(n21267), .B2(n21266), .A(n21265), .ZN(P1_U3465) );
  NAND2_X1 U24167 ( .A1(n21269), .A2(n21268), .ZN(n21274) );
  NAND2_X1 U24168 ( .A1(n21271), .A2(n21270), .ZN(n21272) );
  MUX2_X1 U24169 ( .A(n21272), .B(n11043), .S(n21275), .Z(n21273) );
  OAI21_X1 U24170 ( .B1(n21275), .B2(n21274), .A(n21273), .ZN(P1_U3469) );
  AOI21_X1 U24171 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n21276) );
  AOI22_X1 U24172 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_0__SCAN_IN), 
        .B1(n21276), .B2(n20846), .ZN(n21279) );
  AOI22_X1 U24173 ( .A1(n21282), .A2(n21279), .B1(n21278), .B2(n21277), .ZN(
        P1_U3481) );
  OAI21_X1 U24174 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(P1_REIP_REG_0__SCAN_IN), 
        .A(n21282), .ZN(n21280) );
  OAI21_X1 U24175 ( .B1(n21282), .B2(n21281), .A(n21280), .ZN(P1_U3482) );
  INV_X1 U24176 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n21284) );
  AOI22_X1 U24177 ( .A1(n21296), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n21284), 
        .B2(n21283), .ZN(P1_U3483) );
  AOI211_X1 U24178 ( .C1(n21288), .C2(n21287), .A(n21286), .B(n21285), .ZN(
        n21295) );
  NAND3_X1 U24179 ( .A1(n21290), .A2(P1_STATE2_REG_2__SCAN_IN), .A3(n21289), 
        .ZN(n21292) );
  AOI21_X1 U24180 ( .B1(P1_STATE2_REG_0__SCAN_IN), .B2(n21292), .A(n21291), 
        .ZN(n21294) );
  NAND2_X1 U24181 ( .A1(n21295), .A2(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n21293) );
  OAI21_X1 U24182 ( .B1(n21295), .B2(n21294), .A(n21293), .ZN(P1_U3485) );
  MUX2_X1 U24183 ( .A(P1_M_IO_N_REG_SCAN_IN), .B(P1_MEMORYFETCH_REG_SCAN_IN), 
        .S(n21296), .Z(P1_U3486) );
  NAND2_X1 U12231 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n19506) );
  INV_X1 U11593 ( .A(n12838), .ZN(n9740) );
  NAND2_X1 U12715 ( .A1(n10075), .A2(n10074), .ZN(n15978) );
  CLKBUF_X2 U11181 ( .A(n11159), .Z(n12607) );
  CLKBUF_X1 U11182 ( .A(n9756), .Z(n11217) );
  CLKBUF_X2 U11189 ( .A(n10430), .Z(n13420) );
  CLKBUF_X1 U11194 ( .A(n10920), .Z(n10944) );
  CLKBUF_X1 U11199 ( .A(n12833), .Z(n9748) );
  INV_X2 U11214 ( .A(n17995), .ZN(n17979) );
  CLKBUF_X1 U11219 ( .A(n9765), .Z(n9718) );
  NAND2_X1 U11227 ( .A1(n13141), .A2(n13592), .ZN(n11712) );
  CLKBUF_X1 U11232 ( .A(n18809), .Z(n9712) );
  CLKBUF_X1 U11253 ( .A(n10373), .Z(n11732) );
  CLKBUF_X1 U11264 ( .A(n19700), .Z(n9752) );
  INV_X2 U11466 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n14882) );
  CLKBUF_X1 U11573 ( .A(n18143), .Z(n9754) );
  NOR2_X2 U11605 ( .A1(n13350), .A2(n20120), .ZN(n21297) );
  INV_X2 U11629 ( .A(n19695), .ZN(n19548) );
endmodule

