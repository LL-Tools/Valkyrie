

module b22_C_AntiSAT_k_256_5 ( P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, 
        keyinput128, keyinput129, keyinput130, keyinput131, keyinput132, 
        keyinput133, keyinput134, keyinput135, keyinput136, keyinput137, 
        keyinput138, keyinput139, keyinput140, keyinput141, keyinput142, 
        keyinput143, keyinput144, keyinput145, keyinput146, keyinput147, 
        keyinput148, keyinput149, keyinput150, keyinput151, keyinput152, 
        keyinput153, keyinput154, keyinput155, keyinput156, keyinput157, 
        keyinput158, keyinput159, keyinput160, keyinput161, keyinput162, 
        keyinput163, keyinput164, keyinput165, keyinput166, keyinput167, 
        keyinput168, keyinput169, keyinput170, keyinput171, keyinput172, 
        keyinput173, keyinput174, keyinput175, keyinput176, keyinput177, 
        keyinput178, keyinput179, keyinput180, keyinput181, keyinput182, 
        keyinput183, keyinput184, keyinput185, keyinput186, keyinput187, 
        keyinput188, keyinput189, keyinput190, keyinput191, keyinput192, 
        keyinput193, keyinput194, keyinput195, keyinput196, keyinput197, 
        keyinput198, keyinput199, keyinput200, keyinput201, keyinput202, 
        keyinput203, keyinput204, keyinput205, keyinput206, keyinput207, 
        keyinput208, keyinput209, keyinput210, keyinput211, keyinput212, 
        keyinput213, keyinput214, keyinput215, keyinput216, keyinput217, 
        keyinput218, keyinput219, keyinput220, keyinput221, keyinput222, 
        keyinput223, keyinput224, keyinput225, keyinput226, keyinput227, 
        keyinput228, keyinput229, keyinput230, keyinput231, keyinput232, 
        keyinput233, keyinput234, keyinput235, keyinput236, keyinput237, 
        keyinput238, keyinput239, keyinput240, keyinput241, keyinput242, 
        keyinput243, keyinput244, keyinput245, keyinput246, keyinput247, 
        keyinput248, keyinput249, keyinput250, keyinput251, keyinput252, 
        keyinput253, keyinput254, keyinput255, SUB_1596_U4, SUB_1596_U62, 
        SUB_1596_U63, SUB_1596_U64, SUB_1596_U65, SUB_1596_U66, SUB_1596_U67, 
        SUB_1596_U68, SUB_1596_U69, SUB_1596_U70, SUB_1596_U54, SUB_1596_U55, 
        SUB_1596_U56, SUB_1596_U57, SUB_1596_U58, SUB_1596_U59, SUB_1596_U60, 
        SUB_1596_U61, SUB_1596_U5, SUB_1596_U53, U29, U28, P1_U3355, P1_U3354, 
        P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, P1_U3347, 
        P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, P1_U3340, 
        P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, P1_U3333, 
        P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, P1_U3326, 
        P1_U3325, P1_U3324, P1_U3445, P1_U3446, P1_U3323, P1_U3322, P1_U3321, 
        P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, P1_U3314, 
        P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, P1_U3307, 
        P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, P1_U3300, 
        P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, P1_U3459, 
        P1_U3462, P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, 
        P1_U3483, P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, 
        P1_U3504, P1_U3507, P1_U3510, P1_U3513, P1_U3515, P1_U3516, P1_U3517, 
        P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, P1_U3524, 
        P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, P1_U3531, 
        P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, P1_U3538, 
        P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, P1_U3545, 
        P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, P1_U3552, 
        P1_U3553, P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, 
        P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, P1_U3288, P1_U3287, 
        P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, P1_U3280, 
        P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, P1_U3273, 
        P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, P1_U3266, 
        P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, P1_U3261, P1_U3260, 
        P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, P1_U3253, 
        P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, P1_U3246, 
        P1_U3245, P1_U3244, P1_U3243, P1_U3560, P1_U3561, P1_U3562, P1_U3563, 
        P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, P1_U3570, 
        P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, P1_U3577, 
        P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, P1_U3584, 
        P1_U3585, P1_U3586, P1_U3587, P1_U3588, P1_U3589, P1_U3590, P1_U3591, 
        P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, P1_U3237, P1_U3236, 
        P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, P1_U3229, 
        P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, 
        P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, 
        P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U4016, P2_U3327, P2_U3326, 
        P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321, P2_U3320, P2_U3319, 
        P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314, P2_U3313, P2_U3312, 
        P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307, P2_U3306, P2_U3305, 
        P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300, P2_U3299, P2_U3298, 
        P2_U3297, P2_U3296, P2_U3416, P2_U3417, P2_U3295, P2_U3294, P2_U3293, 
        P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, 
        P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, 
        P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, 
        P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3430, 
        P2_U3433, P2_U3436, P2_U3439, P2_U3442, P2_U3445, P2_U3448, P2_U3451, 
        P2_U3454, P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, 
        P2_U3475, P2_U3478, P2_U3481, P2_U3484, P2_U3486, P2_U3487, P2_U3488, 
        P2_U3489, P2_U3490, P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, 
        P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, 
        P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, 
        P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, 
        P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, 
        P2_U3524, P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, 
        P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, 
        P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, 
        P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, 
        P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, 
        P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, 
        P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, 
        P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, 
        P2_U3216, P2_U3215, P2_U3214, P2_U3531, P2_U3532, P2_U3533, P2_U3534, 
        P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540, P2_U3541, 
        P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547, P2_U3548, 
        P2_U3549, P2_U3550, P2_U3551, P2_U3552, P2_U3553, P2_U3554, P2_U3555, 
        P2_U3556, P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, 
        P2_U3328, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3088, P2_U3087, P2_U3947, P3_U3295, P3_U3294, 
        P3_U3293, P3_U3292, P3_U3291, P3_U3290, P3_U3289, P3_U3288, P3_U3287, 
        P3_U3286, P3_U3285, P3_U3284, P3_U3283, P3_U3282, P3_U3281, P3_U3280, 
        P3_U3279, P3_U3278, P3_U3277, P3_U3276, P3_U3275, P3_U3274, P3_U3273, 
        P3_U3272, P3_U3271, P3_U3270, P3_U3269, P3_U3268, P3_U3267, P3_U3266, 
        P3_U3265, P3_U3264, P3_U3376, P3_U3377, P3_U3263, P3_U3262, P3_U3261, 
        P3_U3260, P3_U3259, P3_U3258, P3_U3257, P3_U3256, P3_U3255, P3_U3254, 
        P3_U3253, P3_U3252, P3_U3251, P3_U3250, P3_U3249, P3_U3248, P3_U3247, 
        P3_U3246, P3_U3245, P3_U3244, P3_U3243, P3_U3242, P3_U3241, P3_U3240, 
        P3_U3239, P3_U3238, P3_U3237, P3_U3236, P3_U3235, P3_U3234, P3_U3390, 
        P3_U3393, P3_U3396, P3_U3399, P3_U3402, P3_U3405, P3_U3408, P3_U3411, 
        P3_U3414, P3_U3417, P3_U3420, P3_U3423, P3_U3426, P3_U3429, P3_U3432, 
        P3_U3435, P3_U3438, P3_U3441, P3_U3444, P3_U3446, P3_U3447, P3_U3448, 
        P3_U3449, P3_U3450, P3_U3451, P3_U3452, P3_U3453, P3_U3454, P3_U3455, 
        P3_U3456, P3_U3457, P3_U3458, P3_U3459, P3_U3460, P3_U3461, P3_U3462, 
        P3_U3463, P3_U3464, P3_U3465, P3_U3466, P3_U3467, P3_U3468, P3_U3469, 
        P3_U3470, P3_U3471, P3_U3472, P3_U3473, P3_U3474, P3_U3475, P3_U3476, 
        P3_U3477, P3_U3478, P3_U3479, P3_U3480, P3_U3481, P3_U3482, P3_U3483, 
        P3_U3484, P3_U3485, P3_U3486, P3_U3487, P3_U3488, P3_U3489, P3_U3490, 
        P3_U3233, P3_U3232, P3_U3231, P3_U3230, P3_U3229, P3_U3228, P3_U3227, 
        P3_U3226, P3_U3225, P3_U3224, P3_U3223, P3_U3222, P3_U3221, P3_U3220, 
        P3_U3219, P3_U3218, P3_U3217, P3_U3216, P3_U3215, P3_U3214, P3_U3213, 
        P3_U3212, P3_U3211, P3_U3210, P3_U3209, P3_U3208, P3_U3207, P3_U3206, 
        P3_U3205, P3_U3204, P3_U3203, P3_U3202, P3_U3201, P3_U3200, P3_U3199, 
        P3_U3198, P3_U3197, P3_U3196, P3_U3195, P3_U3194, P3_U3193, P3_U3192, 
        P3_U3191, P3_U3190, P3_U3189, P3_U3188, P3_U3187, P3_U3186, P3_U3185, 
        P3_U3184, P3_U3183, P3_U3182, P3_U3491, P3_U3492, P3_U3493, P3_U3494, 
        P3_U3495, P3_U3496, P3_U3497, P3_U3498, P3_U3499, P3_U3500, P3_U3501, 
        P3_U3502, P3_U3503, P3_U3504, P3_U3505, P3_U3506, P3_U3507, P3_U3508, 
        P3_U3509, P3_U3510, P3_U3511, P3_U3512, P3_U3513, P3_U3514, P3_U3515, 
        P3_U3516, P3_U3517, P3_U3518, P3_U3519, P3_U3520, P3_U3521, P3_U3522, 
        P3_U3296, P3_U3181, P3_U3180, P3_U3179, P3_U3178, P3_U3177, P3_U3176, 
        P3_U3175, P3_U3174, P3_U3173, P3_U3172, P3_U3171, P3_U3170, P3_U3169, 
        P3_U3168, P3_U3167, P3_U3166, P3_U3165, P3_U3164, P3_U3163, P3_U3162, 
        P3_U3161, P3_U3160, P3_U3159, P3_U3158, P3_U3157, P3_U3156, P3_U3155, 
        P3_U3154, P3_U3153, P3_U3151, P3_U3150, P3_U3897 );
  input P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput0,
         keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6,
         keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12,
         keyinput13, keyinput14, keyinput15, keyinput16, keyinput17,
         keyinput18, keyinput19, keyinput20, keyinput21, keyinput22,
         keyinput23, keyinput24, keyinput25, keyinput26, keyinput27,
         keyinput28, keyinput29, keyinput30, keyinput31, keyinput32,
         keyinput33, keyinput34, keyinput35, keyinput36, keyinput37,
         keyinput38, keyinput39, keyinput40, keyinput41, keyinput42,
         keyinput43, keyinput44, keyinput45, keyinput46, keyinput47,
         keyinput48, keyinput49, keyinput50, keyinput51, keyinput52,
         keyinput53, keyinput54, keyinput55, keyinput56, keyinput57,
         keyinput58, keyinput59, keyinput60, keyinput61, keyinput62,
         keyinput63, keyinput64, keyinput65, keyinput66, keyinput67,
         keyinput68, keyinput69, keyinput70, keyinput71, keyinput72,
         keyinput73, keyinput74, keyinput75, keyinput76, keyinput77,
         keyinput78, keyinput79, keyinput80, keyinput81, keyinput82,
         keyinput83, keyinput84, keyinput85, keyinput86, keyinput87,
         keyinput88, keyinput89, keyinput90, keyinput91, keyinput92,
         keyinput93, keyinput94, keyinput95, keyinput96, keyinput97,
         keyinput98, keyinput99, keyinput100, keyinput101, keyinput102,
         keyinput103, keyinput104, keyinput105, keyinput106, keyinput107,
         keyinput108, keyinput109, keyinput110, keyinput111, keyinput112,
         keyinput113, keyinput114, keyinput115, keyinput116, keyinput117,
         keyinput118, keyinput119, keyinput120, keyinput121, keyinput122,
         keyinput123, keyinput124, keyinput125, keyinput126, keyinput127,
         keyinput128, keyinput129, keyinput130, keyinput131, keyinput132,
         keyinput133, keyinput134, keyinput135, keyinput136, keyinput137,
         keyinput138, keyinput139, keyinput140, keyinput141, keyinput142,
         keyinput143, keyinput144, keyinput145, keyinput146, keyinput147,
         keyinput148, keyinput149, keyinput150, keyinput151, keyinput152,
         keyinput153, keyinput154, keyinput155, keyinput156, keyinput157,
         keyinput158, keyinput159, keyinput160, keyinput161, keyinput162,
         keyinput163, keyinput164, keyinput165, keyinput166, keyinput167,
         keyinput168, keyinput169, keyinput170, keyinput171, keyinput172,
         keyinput173, keyinput174, keyinput175, keyinput176, keyinput177,
         keyinput178, keyinput179, keyinput180, keyinput181, keyinput182,
         keyinput183, keyinput184, keyinput185, keyinput186, keyinput187,
         keyinput188, keyinput189, keyinput190, keyinput191, keyinput192,
         keyinput193, keyinput194, keyinput195, keyinput196, keyinput197,
         keyinput198, keyinput199, keyinput200, keyinput201, keyinput202,
         keyinput203, keyinput204, keyinput205, keyinput206, keyinput207,
         keyinput208, keyinput209, keyinput210, keyinput211, keyinput212,
         keyinput213, keyinput214, keyinput215, keyinput216, keyinput217,
         keyinput218, keyinput219, keyinput220, keyinput221, keyinput222,
         keyinput223, keyinput224, keyinput225, keyinput226, keyinput227,
         keyinput228, keyinput229, keyinput230, keyinput231, keyinput232,
         keyinput233, keyinput234, keyinput235, keyinput236, keyinput237,
         keyinput238, keyinput239, keyinput240, keyinput241, keyinput242,
         keyinput243, keyinput244, keyinput245, keyinput246, keyinput247,
         keyinput248, keyinput249, keyinput250, keyinput251, keyinput252,
         keyinput253, keyinput254, keyinput255;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665,
         n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675,
         n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685,
         n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695,
         n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705,
         n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715,
         n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725,
         n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735,
         n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745,
         n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755,
         n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765,
         n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775,
         n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785,
         n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795,
         n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805,
         n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815,
         n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825,
         n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835,
         n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845,
         n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855,
         n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865,
         n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875,
         n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885,
         n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895,
         n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905,
         n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915,
         n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925,
         n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935,
         n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945,
         n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955,
         n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965,
         n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975,
         n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985,
         n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995,
         n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005,
         n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015,
         n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025,
         n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035,
         n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045,
         n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055,
         n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065,
         n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075,
         n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085,
         n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095,
         n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105,
         n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115,
         n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125,
         n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135,
         n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145,
         n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155,
         n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165,
         n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175,
         n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185,
         n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195,
         n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205,
         n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215,
         n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225,
         n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235,
         n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245,
         n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255,
         n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265,
         n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275,
         n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285,
         n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295,
         n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305,
         n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315,
         n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325,
         n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335,
         n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345,
         n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355,
         n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365,
         n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375,
         n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385,
         n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395,
         n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405,
         n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415,
         n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425,
         n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435,
         n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445,
         n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455,
         n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465,
         n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475,
         n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485,
         n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495,
         n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505,
         n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515,
         n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525,
         n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535,
         n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545,
         n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555,
         n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565,
         n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575,
         n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585,
         n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595,
         n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605,
         n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615,
         n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625,
         n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635,
         n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645,
         n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655,
         n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665,
         n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675,
         n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685,
         n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695,
         n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705,
         n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715,
         n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725,
         n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735,
         n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745,
         n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755,
         n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765,
         n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775,
         n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785,
         n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795,
         n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805,
         n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815,
         n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825,
         n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835,
         n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845,
         n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855,
         n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865,
         n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875,
         n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885,
         n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895,
         n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905,
         n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915,
         n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925,
         n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935,
         n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945,
         n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955,
         n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965,
         n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975,
         n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985,
         n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995,
         n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005,
         n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015,
         n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025,
         n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035,
         n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045,
         n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055,
         n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065,
         n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075,
         n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085,
         n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095,
         n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105,
         n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115,
         n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125,
         n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135,
         n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145,
         n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155,
         n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165,
         n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175,
         n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185,
         n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195,
         n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205,
         n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215,
         n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225,
         n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235,
         n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245,
         n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255,
         n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265,
         n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275,
         n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285,
         n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295,
         n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305,
         n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315,
         n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325,
         n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335,
         n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345,
         n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355,
         n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365,
         n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375,
         n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385,
         n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395,
         n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405,
         n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415,
         n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425,
         n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435,
         n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445,
         n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455,
         n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465,
         n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475,
         n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485,
         n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495,
         n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505,
         n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515,
         n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525,
         n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535,
         n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545,
         n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555,
         n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565,
         n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575,
         n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585,
         n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595,
         n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605,
         n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615,
         n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625,
         n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635,
         n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645,
         n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655,
         n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665,
         n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675,
         n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685,
         n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695,
         n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705,
         n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715,
         n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725,
         n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735,
         n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745,
         n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755,
         n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765,
         n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775,
         n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785,
         n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795,
         n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805,
         n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815,
         n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825,
         n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835,
         n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845,
         n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855,
         n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865,
         n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875,
         n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885,
         n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895,
         n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905,
         n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915,
         n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925,
         n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935,
         n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945,
         n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955,
         n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965,
         n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975,
         n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985,
         n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995,
         n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005,
         n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015,
         n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025,
         n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035,
         n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045,
         n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055,
         n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065,
         n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075,
         n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085,
         n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095,
         n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105,
         n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115,
         n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125,
         n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135,
         n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145,
         n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155,
         n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165,
         n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175,
         n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185,
         n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195,
         n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205,
         n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215,
         n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225,
         n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235,
         n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245,
         n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255,
         n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265,
         n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275,
         n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285,
         n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295,
         n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305,
         n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315,
         n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325,
         n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335,
         n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345,
         n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355,
         n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365,
         n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375,
         n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385,
         n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395,
         n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405,
         n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415,
         n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425,
         n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435,
         n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445,
         n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455,
         n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465,
         n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475,
         n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485,
         n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495,
         n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505,
         n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515,
         n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525,
         n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535,
         n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545,
         n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555,
         n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565,
         n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575,
         n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585,
         n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595,
         n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605,
         n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615,
         n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625,
         n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635,
         n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645,
         n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655,
         n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665,
         n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675,
         n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685,
         n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695,
         n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705,
         n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715,
         n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725,
         n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735,
         n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745,
         n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755,
         n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765,
         n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775,
         n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785,
         n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795,
         n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805,
         n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815,
         n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825,
         n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835,
         n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845,
         n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855,
         n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865,
         n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875,
         n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885,
         n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895,
         n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905,
         n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915,
         n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925,
         n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935,
         n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945,
         n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955,
         n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965,
         n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975,
         n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985,
         n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995,
         n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004,
         n10005, n10006, n10007, n10008, n10009, n10010, n10011, n10012,
         n10013, n10014, n10015, n10016, n10017, n10018, n10019, n10020,
         n10021, n10022, n10023, n10024, n10025, n10026, n10027, n10028,
         n10029, n10030, n10031, n10032, n10033, n10034, n10035, n10036,
         n10037, n10038, n10039, n10040, n10041, n10042, n10043, n10044,
         n10045, n10046, n10047, n10048, n10049, n10050, n10051, n10052,
         n10053, n10054, n10055, n10056, n10057, n10058, n10059, n10060,
         n10061, n10062, n10063, n10064, n10065, n10066, n10067, n10068,
         n10069, n10070, n10071, n10072, n10073, n10074, n10075, n10076,
         n10077, n10078, n10079, n10080, n10081, n10082, n10083, n10084,
         n10085, n10086, n10087, n10088, n10089, n10090, n10091, n10092,
         n10093, n10094, n10095, n10096, n10097, n10098, n10099, n10100,
         n10101, n10102, n10103, n10104, n10105, n10106, n10107, n10108,
         n10109, n10110, n10111, n10112, n10113, n10114, n10115, n10116,
         n10117, n10118, n10119, n10120, n10121, n10122, n10123, n10124,
         n10125, n10126, n10127, n10128, n10129, n10130, n10131, n10132,
         n10133, n10134, n10135, n10136, n10137, n10138, n10139, n10140,
         n10141, n10142, n10143, n10144, n10145, n10146, n10147, n10148,
         n10149, n10150, n10151, n10152, n10153, n10154, n10155, n10156,
         n10157, n10158, n10159, n10160, n10161, n10162, n10163, n10164,
         n10165, n10166, n10167, n10168, n10169, n10170, n10171, n10172,
         n10173, n10174, n10175, n10176, n10177, n10178, n10179, n10180,
         n10181, n10182, n10183, n10184, n10185, n10186, n10187, n10188,
         n10189, n10190, n10191, n10192, n10193, n10194, n10195, n10196,
         n10197, n10198, n10199, n10200, n10201, n10202, n10203, n10204,
         n10205, n10206, n10207, n10208, n10209, n10210, n10211, n10212,
         n10213, n10214, n10215, n10216, n10217, n10218, n10219, n10220,
         n10221, n10222, n10223, n10224, n10225, n10226, n10227, n10228,
         n10229, n10230, n10231, n10232, n10233, n10234, n10235, n10236,
         n10237, n10238, n10239, n10240, n10241, n10242, n10243, n10244,
         n10245, n10246, n10247, n10248, n10249, n10250, n10251, n10252,
         n10253, n10254, n10255, n10256, n10257, n10258, n10259, n10260,
         n10261, n10262, n10263, n10264, n10265, n10266, n10267, n10268,
         n10269, n10270, n10271, n10272, n10273, n10274, n10275, n10276,
         n10277, n10278, n10279, n10280, n10281, n10282, n10283, n10284,
         n10285, n10286, n10287, n10288, n10289, n10290, n10291, n10292,
         n10293, n10294, n10295, n10296, n10297, n10298, n10299, n10300,
         n10301, n10302, n10303, n10304, n10305, n10306, n10307, n10308,
         n10309, n10310, n10311, n10312, n10313, n10314, n10315, n10316,
         n10317, n10318, n10319, n10320, n10321, n10322, n10323, n10324,
         n10325, n10326, n10327, n10328, n10329, n10330, n10331, n10332,
         n10333, n10334, n10335, n10336, n10337, n10338, n10339, n10340,
         n10341, n10342, n10343, n10344, n10345, n10346, n10347, n10348,
         n10349, n10350, n10351, n10352, n10353, n10354, n10355, n10356,
         n10357, n10358, n10359, n10360, n10361, n10362, n10363, n10364,
         n10365, n10366, n10367, n10368, n10369, n10370, n10371, n10372,
         n10373, n10374, n10375, n10376, n10377, n10378, n10379, n10380,
         n10381, n10382, n10383, n10384, n10385, n10386, n10387, n10388,
         n10389, n10390, n10391, n10392, n10393, n10394, n10395, n10396,
         n10397, n10398, n10399, n10400, n10401, n10402, n10403, n10404,
         n10405, n10406, n10407, n10408, n10409, n10410, n10411, n10412,
         n10413, n10414, n10415, n10416, n10417, n10418, n10419, n10420,
         n10421, n10422, n10423, n10424, n10425, n10426, n10427, n10428,
         n10429, n10430, n10431, n10432, n10433, n10434, n10435, n10436,
         n10437, n10438, n10439, n10440, n10441, n10442, n10443, n10444,
         n10445, n10446, n10447, n10448, n10449, n10450, n10451, n10452,
         n10453, n10454, n10455, n10456, n10457, n10458, n10459, n10460,
         n10461, n10462, n10463, n10464, n10465, n10466, n10467, n10468,
         n10469, n10470, n10471, n10472, n10473, n10474, n10475, n10476,
         n10477, n10478, n10479, n10480, n10481, n10482, n10483, n10484,
         n10485, n10486, n10487, n10488, n10489, n10490, n10491, n10492,
         n10493, n10494, n10495, n10496, n10497, n10498, n10499, n10500,
         n10501, n10502, n10503, n10504, n10505, n10506, n10507, n10508,
         n10509, n10510, n10511, n10512, n10513, n10514, n10515, n10516,
         n10517, n10518, n10519, n10520, n10521, n10522, n10523, n10524,
         n10525, n10526, n10527, n10528, n10529, n10530, n10531, n10532,
         n10533, n10534, n10535, n10536, n10537, n10538, n10539, n10540,
         n10541, n10542, n10543, n10544, n10545, n10546, n10547, n10548,
         n10549, n10550, n10551, n10552, n10553, n10554, n10555, n10556,
         n10557, n10558, n10559, n10560, n10561, n10562, n10563, n10564,
         n10565, n10566, n10567, n10568, n10569, n10570, n10571, n10572,
         n10573, n10574, n10575, n10576, n10577, n10578, n10579, n10580,
         n10581, n10582, n10583, n10584, n10585, n10586, n10587, n10588,
         n10589, n10590, n10591, n10592, n10593, n10594, n10595, n10596,
         n10597, n10598, n10599, n10600, n10601, n10602, n10603, n10604,
         n10605, n10606, n10607, n10608, n10609, n10610, n10611, n10612,
         n10613, n10614, n10615, n10616, n10617, n10618, n10619, n10620,
         n10621, n10622, n10623, n10624, n10625, n10626, n10627, n10628,
         n10629, n10630, n10631, n10632, n10633, n10634, n10635, n10636,
         n10637, n10638, n10639, n10640, n10641, n10642, n10643, n10644,
         n10645, n10646, n10647, n10648, n10649, n10650, n10651, n10652,
         n10653, n10654, n10655, n10656, n10657, n10658, n10659, n10660,
         n10661, n10662, n10663, n10664, n10665, n10666, n10667, n10668,
         n10669, n10670, n10671, n10672, n10673, n10674, n10675, n10676,
         n10677, n10678, n10679, n10680, n10681, n10682, n10683, n10684,
         n10685, n10686, n10687, n10688, n10689, n10690, n10691, n10692,
         n10693, n10694, n10695, n10696, n10697, n10698, n10699, n10700,
         n10701, n10702, n10703, n10704, n10705, n10706, n10707, n10708,
         n10709, n10710, n10711, n10712, n10713, n10714, n10715, n10716,
         n10717, n10718, n10719, n10720, n10721, n10722, n10723, n10724,
         n10725, n10726, n10727, n10728, n10729, n10730, n10731, n10732,
         n10733, n10734, n10735, n10736, n10737, n10738, n10739, n10740,
         n10741, n10742, n10743, n10744, n10745, n10746, n10747, n10748,
         n10749, n10750, n10751, n10752, n10753, n10754, n10755, n10756,
         n10757, n10758, n10759, n10760, n10761, n10762, n10763, n10764,
         n10765, n10766, n10767, n10768, n10769, n10770, n10771, n10772,
         n10773, n10774, n10775, n10776, n10777, n10778, n10779, n10780,
         n10781, n10782, n10783, n10784, n10785, n10786, n10787, n10788,
         n10789, n10790, n10791, n10792, n10793, n10794, n10795, n10796,
         n10797, n10798, n10799, n10800, n10801, n10802, n10803, n10804,
         n10805, n10806, n10807, n10808, n10809, n10810, n10811, n10812,
         n10813, n10814, n10815, n10816, n10817, n10818, n10819, n10820,
         n10821, n10822, n10823, n10824, n10825, n10826, n10827, n10828,
         n10829, n10830, n10831, n10832, n10833, n10834, n10835, n10836,
         n10837, n10838, n10839, n10840, n10841, n10842, n10843, n10844,
         n10845, n10846, n10847, n10848, n10849, n10850, n10851, n10852,
         n10853, n10854, n10855, n10856, n10857, n10858, n10859, n10860,
         n10861, n10862, n10863, n10864, n10865, n10866, n10867, n10868,
         n10869, n10870, n10871, n10872, n10873, n10874, n10875, n10876,
         n10877, n10878, n10879, n10880, n10881, n10882, n10883, n10884,
         n10885, n10886, n10887, n10888, n10889, n10890, n10891, n10892,
         n10893, n10894, n10895, n10896, n10897, n10898, n10899, n10900,
         n10901, n10902, n10903, n10904, n10905, n10906, n10907, n10908,
         n10909, n10910, n10911, n10912, n10913, n10914, n10915, n10916,
         n10917, n10918, n10919, n10920, n10921, n10922, n10923, n10924,
         n10925, n10926, n10927, n10928, n10929, n10930, n10931, n10932,
         n10933, n10934, n10935, n10936, n10937, n10938, n10939, n10940,
         n10941, n10942, n10943, n10944, n10945, n10946, n10947, n10948,
         n10949, n10950, n10951, n10952, n10953, n10954, n10955, n10956,
         n10957, n10958, n10959, n10960, n10961, n10962, n10963, n10964,
         n10965, n10966, n10967, n10968, n10969, n10970, n10971, n10972,
         n10973, n10974, n10975, n10976, n10977, n10978, n10979, n10980,
         n10981, n10982, n10983, n10984, n10985, n10986, n10987, n10988,
         n10989, n10990, n10991, n10992, n10993, n10994, n10995, n10996,
         n10997, n10998, n10999, n11000, n11001, n11002, n11003, n11004,
         n11005, n11006, n11007, n11008, n11009, n11010, n11011, n11012,
         n11013, n11014, n11015, n11016, n11017, n11018, n11019, n11020,
         n11021, n11022, n11023, n11024, n11025, n11026, n11027, n11028,
         n11029, n11030, n11031, n11032, n11033, n11034, n11035, n11036,
         n11037, n11038, n11039, n11040, n11041, n11042, n11043, n11044,
         n11045, n11046, n11047, n11048, n11049, n11050, n11051, n11052,
         n11053, n11054, n11055, n11056, n11057, n11058, n11059, n11060,
         n11061, n11062, n11063, n11064, n11065, n11066, n11067, n11068,
         n11069, n11070, n11071, n11072, n11073, n11074, n11075, n11076,
         n11077, n11078, n11079, n11080, n11081, n11082, n11083, n11084,
         n11085, n11086, n11087, n11088, n11089, n11090, n11091, n11092,
         n11093, n11094, n11095, n11096, n11097, n11098, n11099, n11100,
         n11101, n11102, n11103, n11104, n11105, n11106, n11107, n11108,
         n11109, n11110, n11111, n11112, n11113, n11114, n11115, n11116,
         n11117, n11118, n11119, n11120, n11121, n11122, n11123, n11124,
         n11125, n11126, n11127, n11128, n11129, n11130, n11131, n11132,
         n11133, n11134, n11135, n11136, n11137, n11138, n11139, n11140,
         n11141, n11142, n11143, n11144, n11145, n11146, n11147, n11148,
         n11149, n11150, n11151, n11152, n11153, n11154, n11155, n11156,
         n11157, n11158, n11159, n11160, n11161, n11162, n11163, n11164,
         n11165, n11166, n11167, n11168, n11169, n11170, n11171, n11172,
         n11173, n11174, n11175, n11176, n11177, n11178, n11179, n11180,
         n11181, n11182, n11183, n11184, n11185, n11186, n11187, n11188,
         n11189, n11190, n11191, n11192, n11193, n11194, n11195, n11196,
         n11197, n11198, n11199, n11200, n11201, n11202, n11203, n11204,
         n11205, n11206, n11207, n11208, n11209, n11210, n11211, n11212,
         n11213, n11214, n11215, n11216, n11217, n11218, n11219, n11220,
         n11221, n11222, n11223, n11224, n11225, n11226, n11227, n11228,
         n11229, n11230, n11231, n11232, n11233, n11234, n11235, n11236,
         n11237, n11238, n11239, n11240, n11241, n11242, n11243, n11244,
         n11245, n11246, n11247, n11248, n11249, n11250, n11251, n11252,
         n11253, n11254, n11255, n11256, n11257, n11258, n11259, n11260,
         n11261, n11262, n11263, n11264, n11265, n11266, n11267, n11268,
         n11269, n11270, n11271, n11272, n11273, n11274, n11275, n11276,
         n11277, n11278, n11279, n11280, n11281, n11282, n11283, n11284,
         n11285, n11286, n11287, n11288, n11289, n11290, n11291, n11292,
         n11293, n11294, n11295, n11296, n11297, n11298, n11299, n11300,
         n11301, n11302, n11303, n11304, n11305, n11306, n11307, n11308,
         n11309, n11310, n11311, n11312, n11313, n11314, n11315, n11316,
         n11317, n11318, n11319, n11320, n11321, n11322, n11323, n11324,
         n11325, n11326, n11327, n11328, n11329, n11330, n11331, n11332,
         n11333, n11334, n11335, n11336, n11337, n11338, n11339, n11340,
         n11341, n11342, n11343, n11344, n11345, n11346, n11347, n11348,
         n11349, n11350, n11351, n11352, n11353, n11354, n11355, n11356,
         n11357, n11358, n11359, n11360, n11361, n11362, n11363, n11364,
         n11365, n11366, n11367, n11368, n11369, n11370, n11371, n11372,
         n11373, n11374, n11375, n11376, n11377, n11378, n11379, n11380,
         n11381, n11382, n11383, n11384, n11385, n11386, n11387, n11388,
         n11389, n11390, n11391, n11392, n11393, n11394, n11395, n11396,
         n11397, n11398, n11399, n11400, n11401, n11402, n11403, n11404,
         n11405, n11406, n11407, n11408, n11409, n11410, n11411, n11412,
         n11413, n11414, n11415, n11416, n11417, n11418, n11419, n11420,
         n11421, n11422, n11423, n11424, n11425, n11426, n11427, n11428,
         n11429, n11430, n11431, n11432, n11433, n11434, n11435, n11436,
         n11437, n11438, n11439, n11440, n11441, n11442, n11443, n11444,
         n11445, n11446, n11447, n11448, n11449, n11450, n11451, n11452,
         n11453, n11454, n11455, n11456, n11457, n11458, n11459, n11460,
         n11461, n11462, n11463, n11464, n11465, n11466, n11467, n11468,
         n11469, n11470, n11471, n11472, n11473, n11474, n11475, n11476,
         n11477, n11478, n11479, n11480, n11481, n11482, n11483, n11484,
         n11485, n11486, n11487, n11488, n11489, n11490, n11491, n11492,
         n11493, n11494, n11495, n11496, n11497, n11498, n11499, n11500,
         n11501, n11502, n11503, n11504, n11505, n11506, n11507, n11508,
         n11509, n11510, n11511, n11512, n11513, n11514, n11515, n11516,
         n11517, n11518, n11519, n11520, n11521, n11522, n11523, n11524,
         n11525, n11526, n11527, n11528, n11529, n11530, n11531, n11532,
         n11533, n11534, n11535, n11536, n11537, n11538, n11539, n11540,
         n11541, n11542, n11543, n11544, n11545, n11546, n11547, n11548,
         n11549, n11550, n11551, n11552, n11553, n11554, n11555, n11556,
         n11557, n11558, n11559, n11560, n11561, n11562, n11563, n11564,
         n11565, n11566, n11567, n11568, n11569, n11570, n11571, n11572,
         n11573, n11574, n11575, n11576, n11577, n11578, n11579, n11580,
         n11581, n11582, n11583, n11584, n11585, n11586, n11587, n11588,
         n11589, n11590, n11591, n11592, n11593, n11594, n11595, n11596,
         n11597, n11598, n11599, n11600, n11601, n11602, n11603, n11604,
         n11605, n11606, n11607, n11608, n11609, n11610, n11611, n11612,
         n11613, n11614, n11615, n11616, n11617, n11618, n11619, n11620,
         n11621, n11622, n11623, n11624, n11625, n11626, n11627, n11628,
         n11629, n11630, n11631, n11632, n11633, n11634, n11635, n11636,
         n11637, n11638, n11639, n11640, n11641, n11642, n11643, n11644,
         n11645, n11646, n11647, n11648, n11649, n11650, n11651, n11652,
         n11653, n11654, n11655, n11656, n11657, n11658, n11659, n11660,
         n11661, n11662, n11663, n11664, n11665, n11666, n11667, n11668,
         n11669, n11670, n11671, n11672, n11673, n11674, n11675, n11676,
         n11677, n11678, n11679, n11680, n11681, n11682, n11683, n11684,
         n11685, n11686, n11687, n11688, n11689, n11690, n11691, n11692,
         n11693, n11694, n11695, n11696, n11697, n11698, n11699, n11700,
         n11701, n11702, n11703, n11704, n11705, n11706, n11707, n11708,
         n11709, n11710, n11711, n11712, n11713, n11714, n11715, n11716,
         n11717, n11718, n11719, n11720, n11721, n11722, n11723, n11724,
         n11725, n11726, n11727, n11728, n11729, n11730, n11731, n11732,
         n11733, n11734, n11735, n11736, n11737, n11738, n11739, n11740,
         n11741, n11742, n11743, n11744, n11745, n11746, n11747, n11748,
         n11749, n11750, n11751, n11752, n11753, n11754, n11755, n11756,
         n11757, n11758, n11759, n11760, n11761, n11762, n11763, n11764,
         n11765, n11766, n11767, n11768, n11769, n11770, n11771, n11772,
         n11773, n11774, n11775, n11776, n11777, n11778, n11779, n11780,
         n11781, n11782, n11783, n11784, n11785, n11786, n11787, n11788,
         n11789, n11790, n11791, n11792, n11793, n11794, n11795, n11796,
         n11797, n11798, n11799, n11800, n11801, n11802, n11803, n11804,
         n11805, n11806, n11807, n11808, n11809, n11810, n11811, n11812,
         n11813, n11814, n11815, n11816, n11817, n11818, n11819, n11820,
         n11821, n11822, n11823, n11824, n11825, n11826, n11827, n11828,
         n11829, n11830, n11831, n11832, n11833, n11834, n11835, n11836,
         n11837, n11838, n11839, n11840, n11841, n11842, n11843, n11844,
         n11845, n11846, n11847, n11848, n11849, n11850, n11851, n11852,
         n11853, n11854, n11855, n11856, n11857, n11858, n11859, n11860,
         n11861, n11862, n11863, n11864, n11865, n11866, n11867, n11868,
         n11869, n11870, n11871, n11872, n11873, n11874, n11875, n11876,
         n11877, n11878, n11879, n11880, n11881, n11882, n11883, n11884,
         n11885, n11886, n11887, n11888, n11889, n11890, n11891, n11892,
         n11893, n11894, n11895, n11896, n11897, n11898, n11899, n11900,
         n11901, n11902, n11903, n11904, n11905, n11906, n11907, n11908,
         n11909, n11910, n11911, n11912, n11913, n11914, n11915, n11916,
         n11917, n11918, n11919, n11920, n11921, n11922, n11923, n11924,
         n11925, n11926, n11927, n11928, n11929, n11930, n11931, n11932,
         n11933, n11934, n11935, n11936, n11937, n11938, n11939, n11940,
         n11941, n11942, n11943, n11944, n11945, n11946, n11947, n11948,
         n11949, n11950, n11951, n11952, n11953, n11954, n11955, n11956,
         n11957, n11958, n11959, n11960, n11961, n11962, n11963, n11964,
         n11965, n11966, n11967, n11968, n11969, n11970, n11971, n11972,
         n11973, n11974, n11975, n11976, n11977, n11978, n11979, n11980,
         n11981, n11982, n11983, n11984, n11985, n11986, n11987, n11988,
         n11989, n11990, n11991, n11992, n11993, n11994, n11995, n11996,
         n11997, n11998, n11999, n12000, n12001, n12002, n12003, n12004,
         n12005, n12006, n12007, n12008, n12009, n12010, n12011, n12012,
         n12013, n12014, n12015, n12016, n12017, n12018, n12019, n12020,
         n12021, n12022, n12023, n12024, n12025, n12026, n12027, n12028,
         n12029, n12030, n12031, n12032, n12033, n12034, n12035, n12036,
         n12037, n12038, n12039, n12040, n12041, n12042, n12043, n12044,
         n12045, n12046, n12047, n12048, n12049, n12050, n12051, n12052,
         n12053, n12054, n12055, n12056, n12057, n12058, n12059, n12060,
         n12061, n12062, n12063, n12064, n12065, n12066, n12067, n12068,
         n12069, n12070, n12071, n12072, n12073, n12074, n12075, n12076,
         n12077, n12078, n12079, n12080, n12081, n12082, n12083, n12084,
         n12085, n12086, n12087, n12088, n12089, n12090, n12091, n12092,
         n12093, n12094, n12095, n12096, n12097, n12098, n12099, n12100,
         n12101, n12102, n12103, n12104, n12105, n12106, n12107, n12108,
         n12109, n12110, n12111, n12112, n12113, n12114, n12115, n12116,
         n12117, n12118, n12119, n12120, n12121, n12122, n12123, n12124,
         n12125, n12126, n12127, n12128, n12129, n12130, n12131, n12132,
         n12133, n12134, n12135, n12136, n12137, n12138, n12139, n12140,
         n12141, n12142, n12143, n12144, n12145, n12146, n12147, n12148,
         n12149, n12150, n12151, n12152, n12153, n12154, n12155, n12156,
         n12157, n12158, n12159, n12160, n12161, n12162, n12163, n12164,
         n12165, n12166, n12167, n12168, n12169, n12170, n12171, n12172,
         n12173, n12174, n12175, n12176, n12177, n12178, n12179, n12180,
         n12181, n12182, n12183, n12184, n12185, n12186, n12187, n12188,
         n12189, n12190, n12191, n12192, n12193, n12194, n12195, n12196,
         n12197, n12198, n12199, n12200, n12201, n12202, n12203, n12204,
         n12205, n12206, n12207, n12208, n12209, n12210, n12211, n12212,
         n12213, n12214, n12215, n12216, n12217, n12218, n12219, n12220,
         n12221, n12222, n12223, n12224, n12225, n12226, n12227, n12228,
         n12229, n12230, n12231, n12232, n12233, n12234, n12235, n12236,
         n12237, n12238, n12239, n12240, n12241, n12242, n12243, n12244,
         n12245, n12246, n12247, n12248, n12249, n12250, n12251, n12252,
         n12253, n12254, n12255, n12256, n12257, n12258, n12259, n12260,
         n12261, n12262, n12263, n12264, n12265, n12266, n12267, n12268,
         n12269, n12270, n12271, n12272, n12273, n12274, n12275, n12276,
         n12277, n12278, n12279, n12280, n12281, n12282, n12283, n12284,
         n12285, n12286, n12287, n12288, n12289, n12290, n12291, n12292,
         n12293, n12294, n12295, n12296, n12297, n12298, n12299, n12300,
         n12301, n12302, n12303, n12304, n12305, n12306, n12307, n12308,
         n12309, n12310, n12311, n12312, n12313, n12314, n12315, n12316,
         n12317, n12318, n12319, n12320, n12321, n12322, n12323, n12324,
         n12325, n12326, n12327, n12328, n12329, n12330, n12331, n12332,
         n12333, n12334, n12335, n12336, n12337, n12338, n12339, n12340,
         n12341, n12342, n12343, n12344, n12345, n12346, n12347, n12348,
         n12349, n12350, n12351, n12352, n12353, n12354, n12355, n12356,
         n12357, n12358, n12359, n12360, n12361, n12362, n12363, n12364,
         n12365, n12366, n12367, n12368, n12369, n12370, n12371, n12372,
         n12373, n12374, n12375, n12376, n12377, n12378, n12379, n12380,
         n12381, n12382, n12383, n12384, n12385, n12386, n12387, n12388,
         n12389, n12390, n12391, n12392, n12393, n12394, n12395, n12396,
         n12397, n12398, n12399, n12400, n12401, n12402, n12403, n12404,
         n12405, n12406, n12407, n12408, n12409, n12410, n12411, n12412,
         n12413, n12414, n12415, n12416, n12417, n12418, n12419, n12420,
         n12421, n12422, n12423, n12424, n12425, n12426, n12427, n12428,
         n12429, n12430, n12431, n12432, n12433, n12434, n12435, n12436,
         n12437, n12438, n12439, n12440, n12441, n12442, n12443, n12444,
         n12445, n12446, n12447, n12448, n12449, n12450, n12451, n12452,
         n12453, n12454, n12455, n12456, n12457, n12458, n12459, n12460,
         n12461, n12462, n12463, n12464, n12465, n12466, n12467, n12468,
         n12469, n12470, n12471, n12472, n12473, n12474, n12475, n12476,
         n12477, n12478, n12479, n12480, n12481, n12482, n12483, n12484,
         n12485, n12486, n12487, n12488, n12489, n12490, n12491, n12492,
         n12493, n12494, n12495, n12496, n12497, n12498, n12499, n12500,
         n12501, n12502, n12503, n12504, n12505, n12506, n12507, n12508,
         n12509, n12510, n12511, n12512, n12513, n12514, n12515, n12516,
         n12517, n12518, n12519, n12520, n12521, n12522, n12523, n12524,
         n12525, n12526, n12527, n12528, n12529, n12530, n12531, n12532,
         n12533, n12534, n12535, n12536, n12537, n12538, n12539, n12540,
         n12541, n12542, n12543, n12544, n12545, n12546, n12547, n12548,
         n12549, n12550, n12551, n12552, n12553, n12554, n12555, n12556,
         n12557, n12558, n12559, n12560, n12561, n12562, n12563, n12564,
         n12565, n12566, n12567, n12568, n12569, n12570, n12571, n12572,
         n12573, n12574, n12575, n12576, n12577, n12578, n12579, n12580,
         n12581, n12582, n12583, n12584, n12585, n12586, n12587, n12588,
         n12589, n12590, n12591, n12592, n12593, n12594, n12595, n12596,
         n12597, n12598, n12599, n12600, n12601, n12602, n12603, n12604,
         n12605, n12606, n12607, n12608, n12609, n12610, n12611, n12612,
         n12613, n12614, n12615, n12616, n12617, n12618, n12619, n12620,
         n12621, n12622, n12623, n12624, n12625, n12626, n12627, n12628,
         n12629, n12630, n12631, n12632, n12633, n12634, n12635, n12636,
         n12637, n12638, n12639, n12640, n12641, n12642, n12643, n12644,
         n12645, n12646, n12647, n12648, n12649, n12650, n12651, n12652,
         n12653, n12654, n12655, n12656, n12657, n12658, n12659, n12660,
         n12661, n12662, n12663, n12664, n12665, n12666, n12667, n12668,
         n12669, n12670, n12671, n12672, n12673, n12674, n12675, n12676,
         n12677, n12678, n12679, n12680, n12681, n12682, n12683, n12684,
         n12685, n12686, n12687, n12688, n12689, n12690, n12691, n12692,
         n12693, n12694, n12695, n12696, n12697, n12698, n12699, n12700,
         n12701, n12702, n12703, n12704, n12705, n12706, n12707, n12708,
         n12709, n12710, n12711, n12712, n12713, n12714, n12715, n12716,
         n12717, n12718, n12719, n12720, n12721, n12722, n12723, n12724,
         n12725, n12726, n12727, n12728, n12729, n12730, n12731, n12732,
         n12733, n12734, n12735, n12736, n12737, n12738, n12739, n12740,
         n12741, n12742, n12743, n12744, n12745, n12746, n12747, n12748,
         n12749, n12750, n12751, n12752, n12753, n12754, n12755, n12756,
         n12757, n12758, n12759, n12760, n12761, n12762, n12763, n12764,
         n12765, n12766, n12767, n12768, n12769, n12770, n12771, n12772,
         n12773, n12774, n12775, n12776, n12777, n12778, n12779, n12780,
         n12781, n12782, n12783, n12784, n12785, n12786, n12787, n12788,
         n12789, n12790, n12791, n12792, n12793, n12794, n12795, n12796,
         n12797, n12798, n12799, n12800, n12801, n12802, n12803, n12804,
         n12805, n12806, n12807, n12808, n12809, n12810, n12811, n12812,
         n12813, n12814, n12815, n12816, n12817, n12818, n12819, n12820,
         n12821, n12822, n12823, n12824, n12825, n12826, n12827, n12828,
         n12829, n12830, n12831, n12832, n12833, n12834, n12835, n12836,
         n12837, n12838, n12839, n12840, n12841, n12842, n12843, n12844,
         n12845, n12846, n12847, n12848, n12849, n12850, n12851, n12852,
         n12853, n12854, n12855, n12856, n12857, n12858, n12859, n12860,
         n12861, n12862, n12863, n12864, n12865, n12866, n12867, n12868,
         n12869, n12870, n12871, n12872, n12873, n12874, n12875, n12876,
         n12877, n12878, n12879, n12880, n12881, n12882, n12883, n12884,
         n12885, n12886, n12887, n12888, n12889, n12890, n12891, n12892,
         n12893, n12894, n12895, n12896, n12897, n12898, n12899, n12900,
         n12901, n12902, n12903, n12904, n12905, n12906, n12907, n12908,
         n12909, n12910, n12911, n12912, n12913, n12914, n12915, n12916,
         n12917, n12918, n12919, n12920, n12921, n12922, n12923, n12924,
         n12925, n12926, n12927, n12928, n12929, n12930, n12931, n12932,
         n12933, n12934, n12935, n12936, n12937, n12938, n12939, n12940,
         n12941, n12942, n12943, n12944, n12945, n12946, n12947, n12948,
         n12949, n12950, n12951, n12952, n12953, n12954, n12955, n12956,
         n12957, n12958, n12959, n12960, n12961, n12962, n12963, n12964,
         n12965, n12966, n12967, n12968, n12969, n12970, n12971, n12972,
         n12973, n12974, n12975, n12976, n12977, n12978, n12979, n12980,
         n12981, n12982, n12983, n12984, n12985, n12986, n12987, n12988,
         n12989, n12990, n12991, n12992, n12993, n12994, n12995, n12996,
         n12997, n12998, n12999, n13000, n13001, n13002, n13003, n13004,
         n13005, n13006, n13007, n13008, n13009, n13010, n13011, n13012,
         n13013, n13014, n13015, n13016, n13017, n13018, n13019, n13020,
         n13021, n13022, n13023, n13024, n13025, n13026, n13027, n13028,
         n13029, n13030, n13031, n13032, n13033, n13034, n13035, n13036,
         n13037, n13038, n13039, n13040, n13041, n13042, n13043, n13044,
         n13045, n13046, n13047, n13048, n13049, n13050, n13051, n13052,
         n13053, n13054, n13055, n13056, n13057, n13058, n13059, n13060,
         n13061, n13062, n13063, n13064, n13065, n13066, n13067, n13068,
         n13069, n13070, n13071, n13072, n13073, n13074, n13075, n13076,
         n13077, n13078, n13079, n13080, n13081, n13082, n13083, n13084,
         n13085, n13086, n13087, n13088, n13089, n13090, n13091, n13092,
         n13093, n13094, n13095, n13096, n13097, n13098, n13099, n13100,
         n13101, n13102, n13103, n13104, n13105, n13106, n13107, n13108,
         n13109, n13110, n13111, n13112, n13113, n13114, n13115, n13116,
         n13117, n13118, n13119, n13120, n13121, n13122, n13123, n13124,
         n13125, n13126, n13127, n13128, n13129, n13130, n13131, n13132,
         n13133, n13134, n13135, n13136, n13137, n13138, n13139, n13140,
         n13141, n13142, n13143, n13144, n13145, n13146, n13147, n13148,
         n13149, n13150, n13151, n13152, n13153, n13154, n13155, n13156,
         n13157, n13158, n13159, n13160, n13161, n13162, n13163, n13164,
         n13165, n13166, n13167, n13168, n13169, n13170, n13171, n13172,
         n13173, n13174, n13175, n13176, n13177, n13178, n13179, n13180,
         n13181, n13182, n13183, n13184, n13185, n13186, n13187, n13188,
         n13189, n13190, n13191, n13192, n13193, n13194, n13195, n13196,
         n13197, n13198, n13199, n13200, n13201, n13202, n13203, n13204,
         n13205, n13206, n13207, n13208, n13209, n13210, n13211, n13212,
         n13213, n13214, n13215, n13216, n13217, n13218, n13219, n13220,
         n13221, n13222, n13223, n13224, n13225, n13226, n13227, n13228,
         n13229, n13230, n13231, n13232, n13233, n13234, n13235, n13236,
         n13237, n13238, n13239, n13240, n13241, n13242, n13243, n13244,
         n13245, n13246, n13247, n13248, n13249, n13250, n13251, n13252,
         n13253, n13254, n13255, n13256, n13257, n13258, n13259, n13260,
         n13261, n13262, n13263, n13264, n13265, n13266, n13267, n13268,
         n13269, n13270, n13271, n13272, n13273, n13274, n13275, n13276,
         n13277, n13278, n13279, n13280, n13281, n13282, n13283, n13284,
         n13285, n13286, n13287, n13288, n13289, n13290, n13291, n13292,
         n13293, n13294, n13295, n13296, n13297, n13298, n13299, n13300,
         n13301, n13302, n13303, n13304, n13305, n13306, n13307, n13308,
         n13309, n13310, n13311, n13312, n13313, n13314, n13315, n13316,
         n13317, n13318, n13319, n13320, n13321, n13322, n13323, n13324,
         n13325, n13326, n13327, n13328, n13329, n13330, n13331, n13332,
         n13333, n13334, n13335, n13336, n13337, n13338, n13339, n13340,
         n13341, n13342, n13343, n13344, n13345, n13346, n13347, n13348,
         n13349, n13350, n13351, n13352, n13353, n13354, n13355, n13356,
         n13357, n13358, n13359, n13360, n13361, n13362, n13363, n13364,
         n13365, n13366, n13367, n13368, n13369, n13370, n13371, n13372,
         n13373, n13374, n13375, n13376, n13377, n13378, n13379, n13380,
         n13381, n13382, n13383, n13384, n13385, n13386, n13387, n13388,
         n13389, n13390, n13391, n13392, n13393, n13394, n13395, n13396,
         n13397, n13398, n13399, n13400, n13401, n13402, n13403, n13404,
         n13405, n13406, n13407, n13408, n13409, n13410, n13411, n13412,
         n13413, n13414, n13415, n13416, n13417, n13418, n13419, n13420,
         n13421, n13422, n13423, n13424, n13425, n13426, n13427, n13428,
         n13429, n13430, n13431, n13432, n13433, n13434, n13435, n13436,
         n13437, n13438, n13439, n13440, n13441, n13442, n13443, n13444,
         n13445, n13446, n13447, n13448, n13449, n13450, n13451, n13452,
         n13453, n13454, n13455, n13456, n13457, n13458, n13459, n13460,
         n13461, n13462, n13463, n13464, n13465, n13466, n13467, n13468,
         n13469, n13470, n13471, n13472, n13473, n13474, n13475, n13476,
         n13477, n13478, n13479, n13480, n13481, n13482, n13483, n13484,
         n13485, n13486, n13487, n13488, n13489, n13490, n13491, n13492,
         n13493, n13494, n13495, n13496, n13497, n13498, n13499, n13500,
         n13501, n13502, n13503, n13504, n13505, n13506, n13507, n13508,
         n13509, n13510, n13511, n13512, n13513, n13514, n13515, n13516,
         n13517, n13518, n13519, n13520, n13521, n13522, n13523, n13524,
         n13525, n13526, n13527, n13528, n13529, n13530, n13531, n13532,
         n13533, n13534, n13535, n13536, n13537, n13538, n13539, n13540,
         n13541, n13542, n13543, n13544, n13545, n13546, n13547, n13548,
         n13549, n13550, n13551, n13552, n13553, n13554, n13555, n13556,
         n13557, n13558, n13559, n13560, n13561, n13562, n13563, n13564,
         n13565, n13566, n13567, n13568, n13569, n13570, n13571, n13572,
         n13573, n13574, n13575, n13576, n13577, n13578, n13579, n13580,
         n13581, n13582, n13583, n13584, n13585, n13586, n13587, n13588,
         n13589, n13590, n13591, n13592, n13593, n13594, n13595, n13596,
         n13597, n13598, n13599, n13600, n13601, n13602, n13603, n13604,
         n13605, n13606, n13607, n13608, n13609, n13610, n13611, n13612,
         n13613, n13614, n13615, n13616, n13617, n13618, n13619, n13620,
         n13621, n13622, n13623, n13624, n13625, n13626, n13627, n13628,
         n13629, n13630, n13631, n13632, n13633, n13634, n13635, n13636,
         n13637, n13638, n13639, n13640, n13641, n13642, n13643, n13644,
         n13645, n13646, n13647, n13648, n13649, n13650, n13651, n13652,
         n13653, n13654, n13655, n13656, n13657, n13658, n13659, n13660,
         n13661, n13662, n13663, n13664, n13665, n13666, n13667, n13668,
         n13669, n13670, n13671, n13672, n13673, n13674, n13675, n13676,
         n13677, n13678, n13679, n13680, n13681, n13682, n13683, n13684,
         n13685, n13686, n13687, n13688, n13689, n13690, n13691, n13692,
         n13693, n13694, n13695, n13696, n13697, n13698, n13699, n13700,
         n13701, n13702, n13703, n13704, n13705, n13706, n13707, n13708,
         n13709, n13710, n13711, n13712, n13713, n13714, n13715, n13716,
         n13717, n13718, n13719, n13720, n13721, n13722, n13723, n13724,
         n13725, n13726, n13727, n13728, n13729, n13730, n13731, n13732,
         n13733, n13734, n13735, n13736, n13737, n13738, n13739, n13740,
         n13741, n13742, n13743, n13744, n13745, n13746, n13747, n13748,
         n13749, n13750, n13751, n13752, n13753, n13754, n13755, n13756,
         n13757, n13758, n13759, n13760, n13761, n13762, n13763, n13764,
         n13765, n13766, n13767, n13768, n13769, n13770, n13771, n13772,
         n13773, n13774, n13775, n13776, n13777, n13778, n13779, n13780,
         n13781, n13782, n13783, n13784, n13785, n13786, n13787, n13788,
         n13789, n13790, n13791, n13792, n13793, n13794, n13795, n13796,
         n13797, n13798, n13799, n13800, n13801, n13802, n13803, n13804,
         n13805, n13806, n13807, n13808, n13809, n13810, n13811, n13812,
         n13813, n13814, n13815, n13816, n13817, n13818, n13819, n13820,
         n13821, n13822, n13823, n13824, n13825, n13826, n13827, n13828,
         n13829, n13830, n13831, n13832, n13833, n13834, n13835, n13836,
         n13837, n13838, n13839, n13840, n13841, n13842, n13843, n13844,
         n13845, n13846, n13847, n13848, n13849, n13850, n13851, n13852,
         n13853, n13854, n13855, n13856, n13857, n13858, n13859, n13860,
         n13861, n13862, n13863, n13864, n13865, n13866, n13867, n13868,
         n13869, n13870, n13871, n13872, n13873, n13874, n13875, n13876,
         n13877, n13878, n13879, n13880, n13881, n13882, n13883, n13884,
         n13885, n13886, n13887, n13888, n13889, n13890, n13891, n13892,
         n13893, n13894, n13895, n13896, n13897, n13898, n13899, n13900,
         n13901, n13902, n13903, n13904, n13905, n13906, n13907, n13908,
         n13909, n13910, n13911, n13912, n13913, n13914, n13915, n13916,
         n13917, n13918, n13919, n13920, n13921, n13922, n13923, n13924,
         n13925, n13926, n13927, n13928, n13929, n13930, n13931, n13932,
         n13933, n13934, n13935, n13936, n13937, n13938, n13939, n13940,
         n13941, n13942, n13943, n13944, n13945, n13946, n13947, n13948,
         n13949, n13950, n13951, n13952, n13953, n13954, n13955, n13956,
         n13957, n13958, n13959, n13960, n13961, n13962, n13963, n13964,
         n13965, n13966, n13967, n13968, n13969, n13970, n13971, n13972,
         n13973, n13974, n13975, n13976, n13977, n13978, n13979, n13980,
         n13981, n13982, n13983, n13984, n13985, n13986, n13987, n13988,
         n13989, n13990, n13991, n13992, n13993, n13994, n13995, n13996,
         n13997, n13998, n13999, n14000, n14001, n14002, n14003, n14004,
         n14005, n14006, n14007, n14008, n14009, n14010, n14011, n14012,
         n14013, n14014, n14015, n14016, n14017, n14018, n14019, n14020,
         n14021, n14022, n14023, n14024, n14025, n14026, n14027, n14028,
         n14029, n14030, n14031, n14032, n14033, n14034, n14035, n14036,
         n14037, n14038, n14039, n14040, n14041, n14042, n14043, n14044,
         n14045, n14046, n14047, n14048, n14049, n14050, n14051, n14052,
         n14053, n14054, n14055, n14056, n14057, n14058, n14059, n14060,
         n14061, n14062, n14063, n14064, n14065, n14066, n14067, n14068,
         n14069, n14070, n14071, n14072, n14073, n14074, n14075, n14076,
         n14077, n14078, n14079, n14080, n14081, n14082, n14083, n14084,
         n14085, n14086, n14087, n14088, n14089, n14090, n14091, n14092,
         n14093, n14094, n14095, n14096, n14097, n14098, n14099, n14100,
         n14101, n14102, n14103, n14104, n14105, n14106, n14107, n14108,
         n14109, n14110, n14111, n14112, n14113, n14114, n14115, n14116,
         n14117, n14118, n14119, n14120, n14121, n14122, n14123, n14124,
         n14125, n14126, n14127, n14128, n14129, n14130, n14131, n14132,
         n14133, n14134, n14135, n14136, n14137, n14138, n14139, n14140,
         n14141, n14142, n14143, n14144, n14145, n14146, n14147, n14148,
         n14149, n14150, n14151, n14152, n14153, n14154, n14155, n14156,
         n14157, n14158, n14159, n14160, n14161, n14162, n14163, n14164,
         n14165, n14166, n14167, n14168, n14169, n14170, n14171, n14172,
         n14173, n14174, n14175, n14176, n14177, n14178, n14179, n14180,
         n14181, n14182, n14183, n14184, n14185, n14186, n14187, n14188,
         n14189, n14190, n14191, n14192, n14193, n14194, n14195, n14196,
         n14197, n14198, n14199, n14200, n14201, n14202, n14203, n14204,
         n14205, n14206, n14207, n14208, n14209, n14210, n14211, n14212,
         n14213, n14214, n14215, n14216, n14217, n14218, n14219, n14220,
         n14221, n14222, n14223, n14224, n14225, n14226, n14227, n14228,
         n14229, n14230, n14231, n14232, n14233, n14234, n14235, n14236,
         n14237, n14238, n14239, n14240, n14241, n14242, n14243, n14245,
         n14246, n14247, n14248, n14249, n14250, n14251, n14252, n14253,
         n14254, n14255, n14256, n14257, n14258, n14259, n14260, n14261,
         n14262, n14263, n14264, n14265, n14266, n14267, n14268, n14269,
         n14270, n14271, n14272, n14273, n14274, n14275, n14276, n14277,
         n14278, n14279, n14280, n14281, n14282, n14283, n14284, n14285,
         n14286, n14287, n14288, n14289, n14290, n14291, n14292, n14293,
         n14294, n14295, n14296, n14297, n14298, n14299, n14300, n14301,
         n14302, n14303, n14304, n14305, n14306, n14307, n14308, n14309,
         n14310, n14311, n14312, n14313, n14314, n14315, n14316, n14317,
         n14318, n14319, n14320, n14321, n14322, n14323, n14324, n14325,
         n14326, n14327, n14328, n14329, n14330, n14331, n14332, n14333,
         n14334, n14335, n14336, n14337, n14338, n14339, n14340, n14341,
         n14342, n14343, n14344, n14345, n14346, n14347, n14348, n14349,
         n14350, n14351, n14352, n14353, n14354, n14355, n14356, n14357,
         n14358, n14359, n14360, n14361, n14362, n14363, n14364, n14365,
         n14366, n14367, n14368, n14369, n14370, n14371, n14372, n14373,
         n14374, n14375, n14376, n14377, n14378, n14379, n14380, n14381,
         n14382, n14383, n14384, n14385, n14386, n14387, n14388, n14389,
         n14390, n14391, n14392, n14393, n14394, n14395, n14396, n14397,
         n14398, n14399, n14400, n14401, n14402, n14403, n14404, n14405,
         n14406, n14407, n14408, n14409, n14410, n14411, n14412, n14413,
         n14414, n14415, n14416, n14417, n14418, n14419, n14420, n14421,
         n14422, n14423, n14424, n14425, n14426, n14427, n14428, n14429,
         n14430, n14431, n14432, n14433, n14434, n14435, n14436, n14437,
         n14438, n14439, n14440, n14441, n14442, n14443, n14444, n14445,
         n14446, n14447, n14448, n14449, n14450, n14451, n14452, n14453,
         n14454, n14455, n14456, n14457, n14458, n14459, n14460, n14461,
         n14462, n14463, n14464, n14465, n14466, n14467, n14468, n14469,
         n14470, n14471, n14472, n14473, n14474, n14475, n14476, n14477,
         n14478, n14479, n14480, n14481, n14482, n14483, n14484, n14485,
         n14486, n14487, n14488, n14489, n14490, n14491, n14492, n14493,
         n14494, n14495, n14496, n14497, n14498, n14499, n14500, n14501,
         n14502, n14503, n14504, n14505, n14506, n14507, n14508, n14509,
         n14510, n14511, n14512, n14513, n14514, n14515, n14516, n14517,
         n14518, n14519, n14520, n14521, n14522, n14523, n14524, n14525,
         n14526, n14527, n14528, n14529, n14530, n14531, n14532, n14533,
         n14534, n14535, n14536, n14537, n14538, n14539, n14540, n14541,
         n14542, n14543, n14544, n14545, n14546, n14547, n14548, n14549,
         n14550, n14551, n14552, n14553, n14554, n14555, n14556, n14557,
         n14558, n14559, n14560, n14561, n14562, n14563, n14564, n14565,
         n14566, n14567, n14568, n14569, n14570, n14571, n14572, n14573,
         n14574, n14575, n14576, n14577, n14578, n14579, n14580, n14581,
         n14582, n14583, n14584, n14585, n14586, n14587, n14588, n14589,
         n14590, n14591, n14592, n14593, n14594, n14595, n14596, n14597,
         n14598, n14599, n14600, n14601, n14602, n14603, n14604, n14605,
         n14606, n14607, n14608, n14609, n14610, n14611, n14612, n14613,
         n14614, n14615, n14616, n14617, n14618, n14619, n14620, n14621,
         n14622, n14623, n14624, n14625, n14626, n14627, n14628, n14629,
         n14630, n14631, n14632, n14633, n14634, n14635, n14636, n14637,
         n14638, n14639, n14640, n14641, n14642, n14643, n14644, n14645,
         n14646, n14647, n14648, n14649, n14650, n14651, n14652, n14653,
         n14654, n14655, n14656, n14657, n14658, n14659, n14660, n14661,
         n14662, n14663, n14664, n14665, n14666, n14667, n14668, n14669,
         n14670, n14671, n14672, n14673, n14674, n14675, n14676, n14677,
         n14678, n14679, n14680, n14681, n14682, n14683, n14684, n14685,
         n14686, n14687, n14688, n14689, n14690, n14691, n14692, n14693,
         n14694, n14695, n14696, n14697, n14698, n14699, n14700, n14701,
         n14702, n14703, n14704, n14705, n14706, n14707, n14708, n14709,
         n14710, n14711, n14712, n14713, n14714, n14715, n14716, n14717,
         n14718, n14719, n14720, n14721, n14722, n14723, n14724, n14725,
         n14726, n14727, n14728, n14729, n14730, n14731, n14732, n14733,
         n14734, n14735, n14736, n14737, n14738, n14739, n14740, n14741,
         n14742, n14743, n14744, n14745, n14746, n14747, n14748, n14749,
         n14750, n14751, n14752, n14753, n14754, n14755, n14756, n14757,
         n14758, n14759, n14760, n14761, n14762, n14763, n14764, n14765,
         n14766, n14767, n14768, n14769, n14770, n14771, n14772, n14773,
         n14774, n14775, n14776, n14777, n14778, n14779, n14780, n14781,
         n14782, n14783, n14784, n14785, n14786, n14787, n14788, n14789,
         n14790, n14791, n14792, n14793, n14794, n14795, n14796, n14797,
         n14798, n14799, n14801, n14802, n14803, n14804, n14805, n14806,
         n14807, n14808, n14809, n14810, n14811, n14812, n14813, n14814,
         n14815, n14816, n14817, n14818, n14819, n14820, n14821, n14822,
         n14823, n14824, n14825, n14826, n14827, n14828, n14829, n14830,
         n14831, n14832, n14833, n14834, n14835, n14836, n14837, n14838,
         n14839, n14840, n14841, n14842, n14843, n14844, n14845, n14846,
         n14847, n14848, n14849, n14850, n14851, n14852, n14853, n14854,
         n14855, n14856, n14857, n14858, n14859, n14860, n14861, n14862,
         n14863, n14864, n14865, n14866, n14867, n14868, n14869, n14870,
         n14871, n14872, n14873, n14874, n14875, n14876, n14877, n14878,
         n14879, n14880, n14881, n14882, n14883, n14884, n14885, n14886,
         n14887, n14888, n14889, n14890, n14891, n14892, n14893, n14894,
         n14895, n14896, n14897, n14898, n14899, n14900, n14901, n14902,
         n14903, n14904, n14905, n14906, n14907, n14908, n14909, n14910,
         n14911, n14912, n14913, n14914, n14915, n14916, n14917, n14918,
         n14919, n14920, n14921, n14922, n14923, n14924, n14925, n14926,
         n14927, n14928, n14929, n14930, n14931, n14932, n14933, n14934,
         n14935, n14936, n14937, n14938, n14939, n14940, n14941, n14942,
         n14943, n14944, n14945, n14946, n14947, n14948, n14949, n14950,
         n14951, n14952, n14953, n14954, n14955, n14956, n14957, n14958,
         n14959, n14960, n14961, n14962, n14963, n14964, n14965, n14966,
         n14967, n14968, n14969, n14970, n14971, n14972, n14973, n14974,
         n14975, n14976, n14977, n14978, n14979, n14980, n14981, n14982,
         n14983, n14984, n14985, n14986, n14987, n14988, n14989, n14990,
         n14991, n14992, n14993, n14994, n14995, n14996, n14997, n14998,
         n14999, n15000, n15001, n15002, n15003, n15004, n15005, n15006,
         n15007, n15008, n15009, n15010, n15012, n15013, n15014, n15015,
         n15016, n15017, n15018, n15019, n15020, n15021, n15022, n15023,
         n15024, n15025, n15026, n15027, n15028, n15029, n15030, n15031,
         n15032, n15033, n15034, n15035, n15036, n15037, n15038, n15039,
         n15040, n15041, n15042, n15043, n15044, n15045, n15046, n15047,
         n15048, n15049, n15050, n15051, n15052, n15053, n15054, n15055,
         n15056, n15057, n15058, n15059, n15060, n15061, n15062, n15063,
         n15064, n15065, n15066, n15067, n15068, n15069, n15070, n15071,
         n15072, n15073, n15074, n15075, n15076, n15077, n15078, n15079,
         n15080, n15081, n15082, n15083, n15084, n15085, n15086, n15087,
         n15088, n15089, n15090, n15091, n15092, n15093, n15094, n15095,
         n15096, n15097, n15098, n15099, n15100, n15101, n15102, n15103,
         n15104, n15105, n15106, n15107, n15108, n15109, n15110, n15111,
         n15112, n15113, n15114, n15115, n15116, n15117, n15118, n15119,
         n15120, n15121, n15122, n15123, n15124, n15125, n15126, n15127,
         n15128, n15129, n15130, n15131, n15132, n15133, n15134, n15135,
         n15136, n15137, n15138, n15139, n15140, n15141, n15142, n15143,
         n15144, n15145, n15146, n15147, n15148, n15149, n15150, n15151,
         n15152, n15153, n15154, n15155, n15156, n15157, n15158, n15159,
         n15160, n15161, n15162, n15163, n15164, n15165, n15166, n15167,
         n15168, n15169, n15170, n15171, n15172, n15173, n15174, n15175,
         n15176, n15177, n15178, n15179, n15180, n15181, n15182, n15183,
         n15184, n15185, n15186, n15187, n15188, n15189, n15190, n15191,
         n15192, n15193, n15194, n15195, n15196, n15197, n15198, n15199,
         n15200, n15201, n15202, n15203, n15204, n15205, n15206, n15207,
         n15208, n15209, n15210, n15211, n15212, n15213, n15214, n15215,
         n15216, n15217, n15218, n15219, n15220, n15221, n15222, n15223,
         n15224, n15225, n15226, n15227, n15228, n15229, n15230, n15231,
         n15232, n15233, n15234, n15235, n15236, n15237, n15238, n15239,
         n15240, n15241, n15242, n15243, n15244, n15245, n15246, n15247,
         n15248, n15249, n15250, n15251, n15252, n15253, n15254, n15255,
         n15256, n15257, n15258, n15259, n15260, n15261, n15262, n15263,
         n15264, n15265, n15266, n15267, n15268, n15269, n15270, n15271,
         n15272, n15273, n15274, n15275, n15276, n15277, n15278, n15279,
         n15280, n15281, n15282, n15283, n15284, n15285, n15286, n15287,
         n15288, n15289, n15290, n15291, n15292, n15293, n15294, n15295,
         n15296, n15297, n15298, n15299, n15300, n15301, n15302, n15303,
         n15304, n15305, n15306, n15307, n15308, n15309, n15310, n15311,
         n15312, n15313, n15314, n15315, n15316, n15317, n15318, n15319,
         n15320, n15321, n15322, n15323, n15324, n15325, n15326, n15327,
         n15328, n15329, n15330, n15331, n15332, n15333, n15334, n15335,
         n15336, n15337, n15338, n15339, n15340, n15341, n15342, n15343,
         n15344, n15345, n15346, n15347, n15348, n15349, n15350, n15351,
         n15352, n15353, n15354, n15355, n15356, n15357, n15358, n15359,
         n15360, n15361, n15362, n15363, n15364, n15365, n15366, n15367,
         n15368, n15369, n15370, n15371, n15372, n15373, n15374, n15375,
         n15376, n15377, n15378, n15379, n15380, n15381, n15382, n15383,
         n15384, n15385, n15386, n15387, n15388, n15389, n15390, n15391,
         n15392, n15393, n15394, n15395, n15396, n15397, n15398, n15399,
         n15400, n15401, n15402, n15403, n15404, n15405, n15406, n15407,
         n15408, n15409, n15410, n15411, n15412, n15413, n15414, n15415,
         n15416, n15417, n15418, n15419, n15420, n15421, n15422, n15423,
         n15424, n15425, n15426, n15427, n15428, n15429, n15430, n15431,
         n15432, n15433, n15434, n15435, n15436, n15437, n15438, n15439,
         n15440, n15441, n15442, n15443, n15444, n15445, n15446, n15447,
         n15448, n15449, n15450, n15451, n15452, n15453, n15454, n15455,
         n15456, n15457, n15458, n15459, n15460, n15461, n15462, n15463,
         n15464, n15465, n15466, n15467, n15468, n15469, n15470, n15471,
         n15472, n15473, n15474, n15475, n15476, n15477, n15478, n15479,
         n15480, n15481, n15482, n15483, n15484, n15485, n15486, n15487,
         n15488, n15489, n15490, n15491, n15492, n15493, n15494, n15495,
         n15496, n15497, n15498, n15499, n15500, n15501, n15502, n15503,
         n15504, n15505, n15506, n15507, n15508, n15509, n15510, n15511,
         n15512, n15513, n15514, n15515, n15516, n15517, n15518, n15519,
         n15520, n15521, n15522, n15523, n15524, n15525, n15526, n15527,
         n15528, n15529, n15530, n15531, n15532, n15533, n15534, n15535,
         n15536, n15537, n15538, n15539, n15540, n15541, n15542, n15543,
         n15544, n15545, n15546, n15547, n15548, n15549, n15550, n15551,
         n15552, n15553, n15554, n15555, n15556, n15557, n15558, n15559,
         n15560, n15561, n15562, n15563, n15564, n15565, n15566, n15567,
         n15568, n15569, n15570, n15571, n15572, n15573, n15574, n15575,
         n15576, n15577, n15578, n15579, n15580, n15581, n15582, n15583,
         n15584, n15585, n15586, n15587, n15588, n15589, n15590, n15591,
         n15592, n15593, n15594, n15595, n15596, n15597, n15598, n15599,
         n15600, n15601, n15602, n15603, n15604, n15605, n15606, n15607,
         n15608, n15609, n15610, n15611, n15612, n15613, n15614, n15615,
         n15616, n15617, n15618, n15619, n15620, n15621, n15622, n15623,
         n15624, n15625, n15626, n15627, n15628, n15629, n15630, n15631,
         n15632, n15633, n15634, n15635, n15636, n15637, n15638, n15639,
         n15640, n15641, n15642, n15643, n15644, n15645, n15646, n15647,
         n15648, n15649, n15650, n15651, n15652, n15653, n15654, n15655,
         n15656, n15657, n15658, n15659, n15660, n15661, n15662, n15663,
         n15664, n15665, n15666, n15667, n15668, n15669, n15670, n15671,
         n15672, n15673, n15674, n15675, n15676, n15677, n15678, n15679,
         n15680, n15681, n15682, n15683, n15684, n15685, n15686, n15687,
         n15688, n15689, n15690, n15691, n15692, n15693, n15694, n15695,
         n15696, n15697, n15698, n15699, n15700, n15701, n15702, n15703,
         n15704, n15705, n15706, n15707, n15708, n15709, n15710, n15711,
         n15712, n15713, n15714, n15715, n15716, n15717, n15718, n15719,
         n15720, n15721, n15722, n15723, n15724, n15725, n15726, n15727,
         n15728, n15729, n15730, n15731, n15732, n15733, n15734, n15735,
         n15736, n15737, n15738, n15739, n15740, n15741, n15742, n15743,
         n15744, n15745, n15746, n15747, n15748, n15749, n15750, n15751,
         n15752, n15753, n15754, n15755, n15756, n15757, n15758, n15759,
         n15760, n15761, n15762, n15763, n15764, n15765, n15766, n15767,
         n15768, n15769, n15770, n15771, n15772, n15773, n15774, n15775,
         n15776, n15777, n15778, n15779, n15780, n15781, n15782, n15783,
         n15784, n15785, n15786, n15787, n15788, n15789, n15790, n15791,
         n15792, n15793, n15794, n15795, n15796, n15797, n15798, n15799,
         n15800, n15801, n15802, n15803, n15804, n15805;

  NOR2_X1 U7404 ( .A1(n12183), .A2(n12182), .ZN(n12184) );
  OAI21_X1 U7405 ( .B1(n9106), .B2(n6807), .A(n7727), .ZN(n9147) );
  INV_X1 U7406 ( .A(n12382), .ZN(n8337) );
  CLKBUF_X2 U7407 ( .A(n8751), .Z(n6661) );
  OR2_X1 U7408 ( .A1(n12141), .A2(n12140), .ZN(n11956) );
  INV_X2 U7409 ( .A(n12109), .ZN(n11286) );
  NAND2_X1 U7410 ( .A1(n12120), .A2(n7323), .ZN(n11959) );
  AND2_X1 U7411 ( .A1(n14804), .A2(n9619), .ZN(n11088) );
  INV_X4 U7412 ( .A(n6657), .ZN(n6662) );
  NAND2_X1 U7413 ( .A1(n9557), .A2(n14795), .ZN(n14804) );
  XNOR2_X1 U7414 ( .A(n7508), .B(n9461), .ZN(n9722) );
  INV_X2 U7415 ( .A(n11959), .ZN(n12117) );
  INV_X1 U7416 ( .A(n12593), .ZN(n12585) );
  INV_X1 U7417 ( .A(n12130), .ZN(n12140) );
  INV_X2 U7418 ( .A(n12270), .ZN(n12234) );
  INV_X1 U7420 ( .A(n8059), .ZN(n8429) );
  OAI22_X1 U7421 ( .A1(n14536), .A2(n14535), .B1(n14404), .B2(n14440), .ZN(
        n14519) );
  INV_X1 U7422 ( .A(n7483), .ZN(n14536) );
  INV_X1 U7423 ( .A(n11778), .ZN(n11830) );
  NAND2_X1 U7424 ( .A1(n7928), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7929) );
  NAND2_X1 U7425 ( .A1(n8524), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8526) );
  OR2_X1 U7426 ( .A1(n9167), .A2(n9166), .ZN(n9169) );
  INV_X1 U7427 ( .A(n8013), .ZN(n13058) );
  AND2_X1 U7428 ( .A1(n7673), .A2(n10759), .ZN(n6656) );
  INV_X1 U7429 ( .A(n11865), .ZN(n15144) );
  NAND2_X1 U7430 ( .A1(n12191), .A2(n7622), .ZN(n6657) );
  CLKBUF_X3 U7431 ( .A(n6658), .Z(n11808) );
  AND2_X2 U7432 ( .A1(n14801), .A2(n14804), .ZN(n6658) );
  NOR2_X2 U7433 ( .A1(n9458), .A2(P1_IR_REG_28__SCAN_IN), .ZN(n9556) );
  OR2_X2 U7434 ( .A1(n14869), .A2(P1_ADDR_REG_4__SCAN_IN), .ZN(n7268) );
  CLKBUF_X2 U7435 ( .A(n14228), .Z(n6659) );
  NAND4_X1 U7436 ( .A1(n9838), .A2(n9837), .A3(n9836), .A4(n9835), .ZN(n14228)
         );
  OAI21_X2 U7437 ( .B1(n14183), .B2(n7592), .A(n6871), .ZN(n14134) );
  OAI21_X2 U7438 ( .B1(n14606), .B2(n14400), .A(n14583), .ZN(n14568) );
  NAND2_X2 U7439 ( .A1(n9288), .A2(n14029), .ZN(n8535) );
  AND2_X4 U7440 ( .A1(n8507), .A2(n7622), .ZN(n9214) );
  INV_X1 U7441 ( .A(n14225), .ZN(n10456) );
  OAI21_X2 U7442 ( .B1(n13495), .B2(n7837), .A(n7833), .ZN(n13099) );
  INV_X4 U7443 ( .A(n9817), .ZN(n11657) );
  INV_X2 U7445 ( .A(n9619), .ZN(n14801) );
  INV_X2 U7446 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n14232) );
  NAND4_X2 U7447 ( .A1(n8379), .A2(n8378), .A3(n8377), .A4(n8376), .ZN(n12722)
         );
  AND2_X1 U7448 ( .A1(n8535), .A2(n9816), .ZN(n8751) );
  XNOR2_X2 U7449 ( .A(n10842), .B(n11995), .ZN(n12157) );
  INV_X1 U7450 ( .A(n14223), .ZN(n10842) );
  CLKBUF_X3 U7451 ( .A(n11959), .Z(n6663) );
  OAI21_X2 U7452 ( .B1(n14802), .B2(n12109), .A(n12111), .ZN(n14682) );
  XNOR2_X2 U7453 ( .A(n7929), .B(n7996), .ZN(n12440) );
  XNOR2_X2 U7454 ( .A(n14822), .B(n7269), .ZN(n14883) );
  AND2_X2 U7455 ( .A1(n7271), .A2(n7270), .ZN(n14822) );
  NOR2_X2 U7456 ( .A1(n14829), .A2(n14828), .ZN(n14892) );
  NAND2_X2 U7457 ( .A1(n9640), .A2(n10763), .ZN(n9794) );
  XNOR2_X2 U7458 ( .A(n6836), .B(n6835), .ZN(n14925) );
  XNOR2_X2 U7459 ( .A(n8502), .B(n8501), .ZN(n12191) );
  AND2_X1 U7460 ( .A1(n6841), .A2(n7795), .ZN(n14989) );
  NAND2_X1 U7461 ( .A1(n9210), .A2(n9209), .ZN(n13905) );
  NAND2_X1 U7462 ( .A1(n8205), .A2(n12516), .ZN(n12895) );
  OR2_X1 U7463 ( .A1(n15096), .A2(n12514), .ZN(n8205) );
  NAND2_X1 U7464 ( .A1(n9021), .A2(n9020), .ZN(n13947) );
  NAND2_X1 U7465 ( .A1(n7176), .A2(n9040), .ZN(n9061) );
  NOR2_X1 U7466 ( .A1(n14935), .A2(n14934), .ZN(n14933) );
  XNOR2_X1 U7467 ( .A(n14890), .B(n15448), .ZN(n14935) );
  NAND2_X1 U7468 ( .A1(n12453), .A2(n12455), .ZN(n12417) );
  XNOR2_X1 U7469 ( .A(n6659), .B(n11957), .ZN(n10132) );
  XNOR2_X1 U7470 ( .A(n14888), .B(n14887), .ZN(n15794) );
  CLKBUF_X2 U7471 ( .A(P3_U3897), .Z(n15577) );
  CLKBUF_X2 U7472 ( .A(P2_U3947), .Z(n6666) );
  INV_X1 U7473 ( .A(n10851), .ZN(n8394) );
  NAND2_X2 U7474 ( .A1(n12444), .A2(n12452), .ZN(n15692) );
  INV_X4 U7475 ( .A(n7915), .ZN(n6664) );
  INV_X1 U7476 ( .A(n9173), .ZN(n9642) );
  NAND2_X1 U7477 ( .A1(n9763), .A2(n7108), .ZN(n11951) );
  INV_X4 U7479 ( .A(n9170), .ZN(n7114) );
  BUF_X1 U7480 ( .A(n9174), .Z(n6670) );
  NOR2_X1 U7481 ( .A1(n14823), .A2(n14824), .ZN(n14825) );
  XNOR2_X1 U7482 ( .A(n8514), .B(n13365), .ZN(n9288) );
  AND2_X1 U7483 ( .A1(n8562), .A2(n6881), .ZN(n8492) );
  AND2_X1 U7484 ( .A1(n7023), .A2(n7022), .ZN(n7021) );
  AOI21_X1 U7485 ( .B1(n12124), .B2(n12123), .A(n12122), .ZN(n12125) );
  OR2_X1 U7486 ( .A1(n14464), .A2(n14463), .ZN(n14697) );
  NAND2_X1 U7487 ( .A1(n14464), .A2(n14463), .ZN(n14696) );
  OAI21_X1 U7488 ( .B1(n13704), .B2(n15573), .A(n7740), .ZN(n7183) );
  OR2_X1 U7489 ( .A1(n7848), .A2(n15771), .ZN(n7847) );
  OR3_X1 U7490 ( .A1(n13729), .A2(n7425), .A3(n7428), .ZN(n7424) );
  NAND2_X1 U7491 ( .A1(n11854), .A2(n7142), .ZN(n12925) );
  AND2_X1 U7492 ( .A1(n7107), .A2(n7106), .ZN(n12183) );
  NAND2_X1 U7493 ( .A1(n13898), .A2(n6924), .ZN(n14001) );
  AND2_X1 U7494 ( .A1(n7197), .A2(n7190), .ZN(n7649) );
  OR2_X1 U7495 ( .A1(n13717), .A2(n7425), .ZN(n7191) );
  NAND2_X1 U7496 ( .A1(n14753), .A2(n14436), .ZN(n14578) );
  CLKBUF_X1 U7497 ( .A(n11904), .Z(n11905) );
  AND2_X1 U7498 ( .A1(n13721), .A2(n13720), .ZN(n13904) );
  CLKBUF_X1 U7499 ( .A(n14429), .Z(n7126) );
  NAND2_X1 U7500 ( .A1(n9169), .A2(n9168), .ZN(n14802) );
  OR2_X1 U7501 ( .A1(n12747), .A2(n12241), .ZN(n12575) );
  NAND2_X1 U7502 ( .A1(n7742), .A2(n7741), .ZN(n13807) );
  OAI21_X1 U7503 ( .B1(n15252), .B2(n7793), .A(n7790), .ZN(n15255) );
  NAND2_X1 U7504 ( .A1(n7437), .A2(n7436), .ZN(n7742) );
  OR4_X1 U7505 ( .A1(n13737), .A2(n13753), .A3(n13749), .A4(n9264), .ZN(n9265)
         );
  NAND2_X1 U7506 ( .A1(n7273), .A2(n15247), .ZN(n15252) );
  NAND2_X1 U7507 ( .A1(n11822), .A2(n11821), .ZN(n14468) );
  NAND2_X1 U7508 ( .A1(n9152), .A2(n9151), .ZN(n9188) );
  OR4_X1 U7509 ( .A1(n13770), .A2(n13800), .A3(n13783), .A4(n9263), .ZN(n9264)
         );
  NAND2_X1 U7510 ( .A1(n15245), .A2(n14916), .ZN(n15248) );
  OAI22_X1 U7511 ( .A1(n7606), .A2(n6862), .B1(n6863), .B2(n7610), .ZN(n14111)
         );
  NAND2_X1 U7512 ( .A1(n11880), .A2(n11879), .ZN(n13503) );
  NAND2_X1 U7513 ( .A1(n7659), .A2(n7657), .ZN(n15205) );
  NAND2_X1 U7514 ( .A1(n15120), .A2(n11877), .ZN(n11880) );
  AND2_X1 U7515 ( .A1(n14561), .A2(n7667), .ZN(n7666) );
  NAND2_X1 U7516 ( .A1(n9086), .A2(n9085), .ZN(n9106) );
  NAND2_X1 U7517 ( .A1(n7353), .A2(n7352), .ZN(n15120) );
  NAND2_X1 U7518 ( .A1(n11733), .A2(n11732), .ZN(n14730) );
  NAND2_X1 U7519 ( .A1(n14911), .A2(n14910), .ZN(n15243) );
  NOR2_X1 U7520 ( .A1(n7438), .A2(n6706), .ZN(n7436) );
  AND2_X1 U7521 ( .A1(n7263), .A2(n15236), .ZN(n14911) );
  NAND2_X1 U7522 ( .A1(n11180), .A2(n11181), .ZN(n11190) );
  NAND2_X1 U7523 ( .A1(n7151), .A2(n13815), .ZN(n13810) );
  AOI21_X1 U7524 ( .B1(n10817), .B2(n6994), .A(n6993), .ZN(n11180) );
  NOR2_X1 U7525 ( .A1(n14759), .A2(n7514), .ZN(n7513) );
  NAND2_X1 U7526 ( .A1(n9061), .A2(n9060), .ZN(n7007) );
  NAND2_X1 U7527 ( .A1(n14952), .A2(n14907), .ZN(n15237) );
  XNOR2_X1 U7528 ( .A(n11544), .B(n11542), .ZN(n11541) );
  OR2_X1 U7529 ( .A1(n6919), .A2(n13965), .ZN(n13821) );
  INV_X1 U7530 ( .A(n7515), .ZN(n7514) );
  NAND2_X1 U7531 ( .A1(n11659), .A2(n11658), .ZN(n14759) );
  NAND2_X1 U7532 ( .A1(n11698), .A2(n11697), .ZN(n14743) );
  OR2_X1 U7533 ( .A1(n9019), .A2(n7719), .ZN(n7715) );
  OR2_X1 U7534 ( .A1(n13681), .A2(n13682), .ZN(n7741) );
  NAND2_X1 U7535 ( .A1(n11563), .A2(n11562), .ZN(n14762) );
  OR2_X1 U7536 ( .A1(n10846), .A2(n12156), .ZN(n15360) );
  NAND2_X1 U7537 ( .A1(n11639), .A2(n11638), .ZN(n14769) );
  NAND2_X1 U7538 ( .A1(n8998), .A2(n8997), .ZN(n9016) );
  XNOR2_X1 U7539 ( .A(n8996), .B(SI_20_), .ZN(n8995) );
  NAND2_X1 U7540 ( .A1(n11453), .A2(n11452), .ZN(n15203) );
  NAND2_X1 U7541 ( .A1(n10570), .A2(n10536), .ZN(n10792) );
  NAND2_X1 U7542 ( .A1(n7029), .A2(n7027), .ZN(n8996) );
  NAND2_X1 U7543 ( .A1(n8803), .A2(n8802), .ZN(n11491) );
  NAND2_X1 U7544 ( .A1(n7751), .A2(n7753), .ZN(n10570) );
  NAND2_X1 U7545 ( .A1(n7234), .A2(n6726), .ZN(n7753) );
  OAI21_X1 U7546 ( .B1(n8182), .B2(n6980), .A(n6975), .ZN(n8207) );
  NAND2_X1 U7547 ( .A1(n7801), .A2(n6731), .ZN(n7800) );
  NAND2_X1 U7548 ( .A1(n10574), .A2(n6920), .ZN(n10891) );
  NAND2_X2 U7549 ( .A1(n10658), .A2(n15711), .ZN(n15719) );
  NAND2_X1 U7550 ( .A1(n9645), .A2(n9644), .ZN(n9695) );
  NAND2_X1 U7551 ( .A1(n8705), .A2(n8704), .ZN(n15538) );
  OAI21_X1 U7552 ( .B1(n8770), .B2(n8769), .A(n8771), .ZN(n8796) );
  INV_X2 U7553 ( .A(n14969), .ZN(n6665) );
  NAND2_X2 U7554 ( .A1(n7570), .A2(n7568), .ZN(n12270) );
  XNOR2_X1 U7555 ( .A(n10242), .B(n10704), .ZN(n10239) );
  NAND2_X1 U7556 ( .A1(n15794), .A2(n15793), .ZN(n15792) );
  BUF_X1 U7557 ( .A(n8679), .Z(n7174) );
  OAI21_X1 U7558 ( .B1(n7180), .B2(n8654), .A(n7005), .ZN(n8679) );
  NAND2_X2 U7559 ( .A1(n8564), .A2(n7147), .ZN(n6989) );
  NAND4_X1 U7560 ( .A1(n8575), .A2(n8574), .A3(n8573), .A4(n8572), .ZN(n13575)
         );
  CLKBUF_X3 U7561 ( .A(n8553), .Z(n9191) );
  AND3_X1 U7562 ( .A1(n7244), .A2(n8582), .A3(n7243), .ZN(n10556) );
  AND2_X1 U7563 ( .A1(n7113), .A2(n8563), .ZN(n7147) );
  AND4_X1 U7564 ( .A1(n8065), .A2(n8064), .A3(n8063), .A4(n8062), .ZN(n10775)
         );
  AND2_X2 U7565 ( .A1(n11956), .A2(n11951), .ZN(n11778) );
  NAND4_X1 U7566 ( .A1(n8039), .A2(n8036), .A3(n8038), .A4(n8037), .ZN(n12637)
         );
  OAI211_X1 U7567 ( .C1(n12109), .C2(n9982), .A(n9981), .B(n9980), .ZN(n11957)
         );
  AND2_X1 U7568 ( .A1(n9176), .A2(n9174), .ZN(n7335) );
  BUF_X1 U7569 ( .A(n15498), .Z(n6672) );
  XNOR2_X1 U7570 ( .A(n9467), .B(n9466), .ZN(n12131) );
  NOR2_X1 U7571 ( .A1(n8014), .A2(n13058), .ZN(n8386) );
  NAND2_X4 U7572 ( .A1(n10021), .A2(n9616), .ZN(n8066) );
  NAND2_X1 U7573 ( .A1(n10021), .A2(n9816), .ZN(n8305) );
  AND2_X2 U7574 ( .A1(n8014), .A2(n13058), .ZN(n8059) );
  AND2_X2 U7575 ( .A1(n8015), .A2(n13058), .ZN(n12382) );
  NAND2_X1 U7576 ( .A1(n9465), .A2(n9464), .ZN(n12141) );
  AND2_X2 U7577 ( .A1(n8014), .A2(n8013), .ZN(n12381) );
  NAND2_X1 U7578 ( .A1(n9611), .A2(n9610), .ZN(n12130) );
  XNOR2_X1 U7579 ( .A(n14825), .B(n7806), .ZN(n14869) );
  XNOR2_X1 U7580 ( .A(n8007), .B(n8006), .ZN(n8014) );
  NAND2_X1 U7581 ( .A1(n9460), .A2(n9554), .ZN(n14807) );
  NAND2_X2 U7582 ( .A1(n8001), .A2(n8000), .ZN(n12694) );
  INV_X1 U7583 ( .A(n9722), .ZN(n6667) );
  MUX2_X1 U7584 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9609), .S(
        P1_IR_REG_20__SCAN_IN), .Z(n9611) );
  NAND2_X1 U7585 ( .A1(n8505), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8502) );
  MUX2_X1 U7586 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9459), .S(
        P1_IR_REG_28__SCAN_IN), .Z(n9460) );
  NAND2_X1 U7587 ( .A1(n6917), .A2(n6906), .ZN(n14029) );
  XNOR2_X1 U7588 ( .A(n9613), .B(P1_IR_REG_19__SCAN_IN), .ZN(n14612) );
  OR2_X1 U7589 ( .A1(n9612), .A2(n6779), .ZN(n9610) );
  NAND2_X2 U7590 ( .A1(n9816), .A2(P1_U3086), .ZN(n14815) );
  OR2_X1 U7591 ( .A1(n9816), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n7417) );
  AOI21_X1 U7592 ( .B1(n7004), .B2(n7003), .A(n7002), .ZN(n6906) );
  AND2_X1 U7593 ( .A1(n7394), .A2(n7393), .ZN(n8138) );
  NOR2_X1 U7594 ( .A1(n9616), .A2(P3_STATE_REG_SCAN_IN), .ZN(n14945) );
  NOR2_X1 U7595 ( .A1(n7039), .A2(n7038), .ZN(n7395) );
  AND2_X1 U7596 ( .A1(n8491), .A2(n8492), .ZN(n7361) );
  AND4_X1 U7597 ( .A1(n7503), .A2(n9310), .A3(n9312), .A4(n9313), .ZN(n7502)
         );
  NOR2_X1 U7598 ( .A1(n7396), .A2(P3_IR_REG_9__SCAN_IN), .ZN(n7394) );
  OAI21_X1 U7599 ( .B1(n14874), .B2(n14876), .A(n7804), .ZN(n7803) );
  NAND2_X1 U7600 ( .A1(n6698), .A2(n7682), .ZN(n7680) );
  AND2_X1 U7601 ( .A1(n6916), .A2(n8494), .ZN(n8495) );
  AND2_X1 U7602 ( .A1(n7909), .A2(n8500), .ZN(n7908) );
  NOR2_X1 U7603 ( .A1(n7998), .A2(P3_IR_REG_17__SCAN_IN), .ZN(n7860) );
  AND3_X1 U7604 ( .A1(n8562), .A2(n6878), .A3(n7869), .ZN(n6876) );
  AND3_X1 U7605 ( .A1(n7553), .A2(n7551), .A3(n7552), .ZN(n6826) );
  AND2_X1 U7606 ( .A1(n7040), .A2(n8466), .ZN(n7584) );
  AND3_X1 U7607 ( .A1(n8851), .A2(n8800), .A3(n8493), .ZN(n6916) );
  AND2_X1 U7608 ( .A1(n6878), .A2(n6877), .ZN(n8491) );
  AND2_X1 U7609 ( .A1(n7589), .A2(n7588), .ZN(n9307) );
  XNOR2_X1 U7610 ( .A(n14232), .B(P3_ADDR_REG_1__SCAN_IN), .ZN(n14874) );
  NOR2_X1 U7611 ( .A1(P3_IR_REG_10__SCAN_IN), .A2(P3_IR_REG_14__SCAN_IN), .ZN(
        n7553) );
  NOR2_X1 U7612 ( .A1(P3_IR_REG_12__SCAN_IN), .A2(P3_IR_REG_11__SCAN_IN), .ZN(
        n7552) );
  NOR2_X1 U7613 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), .ZN(
        n8517) );
  NOR2_X1 U7614 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n7589) );
  NOR2_X1 U7615 ( .A1(P3_IR_REG_13__SCAN_IN), .A2(P3_IR_REG_15__SCAN_IN), .ZN(
        n7551) );
  NOR2_X1 U7616 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_4__SCAN_IN), .ZN(
        n6878) );
  INV_X1 U7617 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n10047) );
  NOR2_X1 U7618 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n6880) );
  NOR2_X1 U7619 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_5__SCAN_IN), .ZN(
        n6879) );
  INV_X1 U7620 ( .A(P3_IR_REG_19__SCAN_IN), .ZN(n13367) );
  INV_X1 U7621 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n9311) );
  INV_X1 U7622 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n10048) );
  INV_X1 U7623 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n10049) );
  NOR2_X1 U7624 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n6877) );
  NOR2_X1 U7625 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n6881) );
  INV_X1 U7626 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n7869) );
  INV_X1 U7627 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n8040) );
  NOR2_X1 U7628 ( .A1(P2_IR_REG_14__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), .ZN(
        n8494) );
  INV_X4 U7629 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  INV_X4 U7630 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  BUF_X2 U7631 ( .A(n9722), .Z(n6668) );
  BUF_X2 U7632 ( .A(n9722), .Z(n6669) );
  XNOR2_X1 U7633 ( .A(n8598), .B(SI_3_), .ZN(n8596) );
  AOI21_X2 U7634 ( .B1(n12320), .B2(n6679), .A(n12319), .ZN(n12298) );
  XNOR2_X1 U7635 ( .A(n8516), .B(n9269), .ZN(n9174) );
  NOR2_X2 U7636 ( .A1(n14882), .A2(n14923), .ZN(n15801) );
  NAND2_X2 U7637 ( .A1(n15792), .A2(n14889), .ZN(n14890) );
  INV_X1 U7638 ( .A(n9170), .ZN(n6671) );
  AND2_X4 U7639 ( .A1(n12191), .A2(n14023), .ZN(n8571) );
  NAND2_X4 U7640 ( .A1(n10073), .A2(n6670), .ZN(n11865) );
  INV_X1 U7641 ( .A(n8386), .ZN(n8375) );
  NAND2_X1 U7642 ( .A1(n7584), .A2(n7248), .ZN(n7039) );
  MUX2_X1 U7643 ( .A(n12587), .B(n12586), .S(n12585), .Z(n12588) );
  NAND2_X1 U7644 ( .A1(n9016), .A2(n9015), .ZN(n9019) );
  NOR2_X1 U7645 ( .A1(n12578), .A2(n7844), .ZN(n7843) );
  INV_X1 U7646 ( .A(n8421), .ZN(n7844) );
  INV_X1 U7647 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n7867) );
  AND4_X1 U7648 ( .A1(n7861), .A2(n7860), .A3(n7394), .A4(n7868), .ZN(n7250)
         );
  AND2_X1 U7649 ( .A1(n8138), .A2(n13367), .ZN(n7292) );
  OR2_X1 U7650 ( .A1(n13905), .A2(n13666), .ZN(n13696) );
  INV_X1 U7651 ( .A(n11488), .ZN(n7220) );
  NAND2_X1 U7652 ( .A1(n9307), .A2(n9306), .ZN(n9339) );
  AND2_X1 U7653 ( .A1(n10048), .A2(n10049), .ZN(n7505) );
  AND4_X1 U7654 ( .A1(n8234), .A2(n8233), .A3(n8232), .A4(n8231), .ZN(n12362)
         );
  AOI21_X1 U7655 ( .B1(n7866), .B2(n7864), .A(n6746), .ZN(n7863) );
  INV_X1 U7656 ( .A(n7866), .ZN(n7865) );
  NAND2_X1 U7657 ( .A1(n8482), .A2(n12402), .ZN(n15695) );
  NAND2_X1 U7658 ( .A1(n9190), .A2(n9189), .ZN(n13901) );
  AND2_X1 U7659 ( .A1(n7430), .A2(n7702), .ZN(n7247) );
  NAND2_X1 U7660 ( .A1(n11490), .A2(n13565), .ZN(n7430) );
  AND2_X1 U7661 ( .A1(n7638), .A2(n8495), .ZN(n7840) );
  NAND2_X1 U7662 ( .A1(n11541), .A2(n11540), .ZN(n11546) );
  INV_X1 U7663 ( .A(n9610), .ZN(n9462) );
  AND2_X1 U7664 ( .A1(n8695), .A2(n8696), .ZN(n7889) );
  NAND2_X1 U7665 ( .A1(n7888), .A2(n7887), .ZN(n7886) );
  INV_X1 U7666 ( .A(n8696), .ZN(n7888) );
  INV_X1 U7667 ( .A(n8695), .ZN(n7887) );
  NAND2_X1 U7668 ( .A1(n8674), .A2(n8676), .ZN(n6904) );
  INV_X1 U7669 ( .A(n12065), .ZN(n7302) );
  NAND2_X1 U7670 ( .A1(n7301), .A2(n7302), .ZN(n7300) );
  MUX2_X1 U7671 ( .A(n14543), .B(n14559), .S(n12117), .Z(n12072) );
  NAND2_X1 U7672 ( .A1(n7102), .A2(n7101), .ZN(n12073) );
  NAND2_X1 U7673 ( .A1(n14569), .A2(n12117), .ZN(n7101) );
  NAND2_X1 U7674 ( .A1(n14160), .A2(n6663), .ZN(n7102) );
  MUX2_X1 U7675 ( .A(n14440), .B(n14730), .S(n6663), .Z(n12075) );
  AND2_X1 U7676 ( .A1(n6728), .A2(n7723), .ZN(n7722) );
  AND2_X1 U7677 ( .A1(n7903), .A2(n9123), .ZN(n7902) );
  NAND2_X1 U7678 ( .A1(n7905), .A2(n7904), .ZN(n7903) );
  OAI21_X1 U7679 ( .B1(n7375), .B2(n12463), .A(n12478), .ZN(n7371) );
  OAI21_X1 U7680 ( .B1(n13497), .B2(n9241), .A(n9076), .ZN(n9077) );
  NAND2_X1 U7681 ( .A1(n7898), .A2(n7900), .ZN(n7896) );
  INV_X1 U7682 ( .A(n7902), .ZN(n7900) );
  NAND2_X1 U7683 ( .A1(n9963), .A2(n7634), .ZN(n7633) );
  NOR2_X1 U7684 ( .A1(n7636), .A2(n7635), .ZN(n7634) );
  INV_X1 U7685 ( .A(n9962), .ZN(n7635) );
  NAND2_X1 U7686 ( .A1(n12118), .A2(n12130), .ZN(n12120) );
  AOI21_X1 U7687 ( .B1(n8929), .B2(n7725), .A(n7724), .ZN(n7723) );
  INV_X1 U7688 ( .A(n8874), .ZN(n7725) );
  INV_X1 U7689 ( .A(n8931), .ZN(n7724) );
  INV_X1 U7690 ( .A(n8929), .ZN(n7726) );
  NAND2_X1 U7691 ( .A1(n8876), .A2(n13439), .ZN(n8931) );
  OAI21_X1 U7692 ( .B1(n12214), .B2(n7285), .A(n7282), .ZN(n12222) );
  AOI21_X1 U7693 ( .B1(n7284), .B2(n7288), .A(n7283), .ZN(n7282) );
  INV_X1 U7694 ( .A(n12221), .ZN(n7283) );
  AND2_X1 U7695 ( .A1(n7858), .A2(n7294), .ZN(n7293) );
  INV_X1 U7696 ( .A(P3_IR_REG_18__SCAN_IN), .ZN(n7294) );
  NAND2_X1 U7697 ( .A1(n12741), .A2(n8420), .ZN(n7845) );
  NOR2_X1 U7698 ( .A1(n12769), .A2(n12770), .ZN(n12568) );
  INV_X1 U7699 ( .A(n8414), .ZN(n7057) );
  OR2_X1 U7700 ( .A1(n12954), .A2(n12216), .ZN(n12550) );
  NAND2_X1 U7701 ( .A1(n11945), .A2(n8019), .ZN(n12590) );
  NAND2_X1 U7702 ( .A1(n7404), .A2(n7402), .ZN(n12377) );
  INV_X1 U7703 ( .A(n7403), .ZN(n7402) );
  OAI21_X1 U7704 ( .B1(n12584), .B2(n12578), .A(n12586), .ZN(n7403) );
  INV_X1 U7705 ( .A(n12440), .ZN(n10656) );
  NAND2_X1 U7706 ( .A1(n6966), .A2(n7974), .ZN(n7975) );
  OAI21_X1 U7707 ( .B1(n8251), .B2(n7523), .A(n7522), .ZN(n6966) );
  INV_X1 U7708 ( .A(n7524), .ZN(n7523) );
  AOI21_X1 U7709 ( .B1(n7524), .B2(n7526), .A(n8279), .ZN(n7522) );
  INV_X1 U7710 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n7957) );
  INV_X1 U7711 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n7953) );
  INV_X1 U7712 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n8800) );
  AOI21_X1 U7713 ( .B1(n7229), .B2(n7228), .A(n13783), .ZN(n7227) );
  INV_X1 U7714 ( .A(n7230), .ZN(n7228) );
  AND2_X1 U7715 ( .A1(n10897), .A2(n10787), .ZN(n7647) );
  INV_X1 U7716 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n13365) );
  INV_X1 U7717 ( .A(n8499), .ZN(n7638) );
  NOR2_X1 U7718 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n7360) );
  OAI21_X1 U7719 ( .B1(n6701), .B2(n7678), .A(n14604), .ZN(n7677) );
  NOR2_X1 U7720 ( .A1(n14561), .A2(n7482), .ZN(n7481) );
  INV_X1 U7721 ( .A(n14402), .ZN(n7482) );
  NAND3_X1 U7722 ( .A1(n7715), .A2(n7718), .A3(n7714), .ZN(n7176) );
  NAND2_X1 U7723 ( .A1(n9019), .A2(n9018), .ZN(n9039) );
  AOI21_X1 U7724 ( .B1(n8796), .B2(n7012), .A(n7009), .ZN(n7008) );
  NAND2_X1 U7725 ( .A1(n7010), .A2(n7746), .ZN(n7009) );
  AOI21_X1 U7726 ( .B1(n8817), .B2(n7748), .A(n7747), .ZN(n7746) );
  AND2_X1 U7727 ( .A1(n8869), .A2(n8850), .ZN(n8867) );
  AOI21_X1 U7728 ( .B1(n7712), .B2(n6688), .A(n6755), .ZN(n7711) );
  NAND2_X1 U7729 ( .A1(n14232), .A2(P3_ADDR_REG_1__SCAN_IN), .ZN(n7804) );
  NOR2_X1 U7730 ( .A1(n14833), .A2(n14832), .ZN(n14898) );
  NAND3_X1 U7731 ( .A1(n7571), .A2(n8453), .A3(n7572), .ZN(n7570) );
  OR2_X1 U7732 ( .A1(n8281), .A2(n6729), .ZN(n8034) );
  INV_X1 U7733 ( .A(n7564), .ZN(n7562) );
  NAND2_X1 U7734 ( .A1(n12440), .A2(n8481), .ZN(n12604) );
  AND4_X1 U7735 ( .A1(n8195), .A2(n8194), .A3(n8193), .A4(n8192), .ZN(n12199)
         );
  AND4_X1 U7736 ( .A1(n8150), .A2(n8149), .A3(n8148), .A4(n8147), .ZN(n12498)
         );
  NAND2_X1 U7737 ( .A1(n8013), .A2(P3_REG3_REG_1__SCAN_IN), .ZN(n7041) );
  XNOR2_X1 U7738 ( .A(n7696), .B(n14928), .ZN(n15601) );
  NOR2_X1 U7739 ( .A1(n12654), .A2(n6801), .ZN(n12656) );
  NAND2_X1 U7740 ( .A1(n7324), .A2(n12689), .ZN(n7688) );
  NAND2_X1 U7741 ( .A1(n7688), .A2(n12691), .ZN(n12661) );
  MUX2_X1 U7742 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7999), .S(
        P3_IR_REG_27__SCAN_IN), .Z(n8001) );
  NAND2_X1 U7743 ( .A1(n8438), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7999) );
  NAND2_X1 U7744 ( .A1(n12318), .A2(n12224), .ZN(n12566) );
  NAND2_X1 U7745 ( .A1(n7059), .A2(n7058), .ZN(n12818) );
  INV_X1 U7746 ( .A(n12816), .ZN(n7059) );
  AND2_X1 U7747 ( .A1(n12854), .A2(n7065), .ZN(n7064) );
  NOR2_X1 U7748 ( .A1(n8408), .A2(n7074), .ZN(n7073) );
  INV_X1 U7749 ( .A(n8407), .ZN(n7074) );
  AND2_X1 U7750 ( .A1(n12478), .A2(n12471), .ZN(n12412) );
  NAND2_X1 U7751 ( .A1(n10852), .A2(n12457), .ZN(n10853) );
  NAND2_X1 U7752 ( .A1(n10851), .A2(n10660), .ZN(n12455) );
  XNOR2_X1 U7753 ( .A(n12377), .B(n6713), .ZN(n11942) );
  INV_X1 U7754 ( .A(n8066), .ZN(n8282) );
  INV_X1 U7755 ( .A(n8305), .ZN(n12394) );
  AND2_X1 U7756 ( .A1(n8465), .A2(n8448), .ZN(n9497) );
  AND4_X1 U7757 ( .A1(n7861), .A2(n7395), .A3(n7860), .A4(n7394), .ZN(n8440)
         );
  INV_X1 U7758 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n8005) );
  AND2_X1 U7759 ( .A1(n8138), .A2(n7582), .ZN(n7581) );
  AND2_X1 U7760 ( .A1(n7584), .A2(n13374), .ZN(n7582) );
  NAND2_X1 U7761 ( .A1(n7977), .A2(n6987), .ZN(n8304) );
  AND2_X1 U7762 ( .A1(n7976), .A2(n7095), .ZN(n6987) );
  INV_X1 U7763 ( .A(n8301), .ZN(n7095) );
  INV_X1 U7764 ( .A(n7531), .ZN(n7528) );
  AND2_X1 U7765 ( .A1(n6826), .A2(n7862), .ZN(n7861) );
  INV_X1 U7766 ( .A(P3_IR_REG_16__SCAN_IN), .ZN(n7862) );
  NAND2_X1 U7767 ( .A1(n8138), .A2(n7858), .ZN(n8263) );
  INV_X1 U7768 ( .A(n7964), .ZN(n7538) );
  OAI21_X1 U7769 ( .B1(n6971), .B2(n6968), .A(n6967), .ZN(n8180) );
  INV_X1 U7770 ( .A(n6969), .ZN(n6968) );
  AOI21_X1 U7771 ( .B1(n6969), .B2(n8152), .A(n6798), .ZN(n6967) );
  AND2_X1 U7772 ( .A1(n6972), .A2(n6800), .ZN(n6969) );
  AND2_X1 U7773 ( .A1(n9236), .A2(n9225), .ZN(n7168) );
  NAND2_X1 U7774 ( .A1(n9266), .A2(n7089), .ZN(n9275) );
  AND2_X1 U7775 ( .A1(n9248), .A2(n7175), .ZN(n7089) );
  AND2_X1 U7776 ( .A1(n9267), .A2(n7425), .ZN(n7175) );
  INV_X1 U7777 ( .A(n12191), .ZN(n8507) );
  NAND2_X1 U7778 ( .A1(n13729), .A2(n13692), .ZN(n13693) );
  INV_X1 U7779 ( .A(n7624), .ZN(n7623) );
  OAI21_X1 U7780 ( .B1(n7627), .B2(n7625), .A(n6739), .ZN(n7624) );
  INV_X1 U7781 ( .A(n13664), .ZN(n7625) );
  OR2_X1 U7782 ( .A1(n13935), .A2(n13497), .ZN(n9251) );
  AND2_X1 U7783 ( .A1(n7239), .A2(n7439), .ZN(n7238) );
  NAND2_X1 U7784 ( .A1(n7240), .A2(n6694), .ZN(n7239) );
  AOI21_X1 U7785 ( .B1(n7211), .B2(n7209), .A(n6745), .ZN(n7208) );
  INV_X1 U7786 ( .A(n13648), .ZN(n7209) );
  NOR2_X1 U7787 ( .A1(n13845), .A2(n13673), .ZN(n6918) );
  OR2_X1 U7788 ( .A1(n13861), .A2(n6694), .ZN(n7241) );
  AOI21_X1 U7789 ( .B1(n6678), .B2(n7218), .A(n6753), .ZN(n7217) );
  INV_X1 U7790 ( .A(n7222), .ZN(n7218) );
  NAND2_X1 U7791 ( .A1(n15133), .A2(n6711), .ZN(n7703) );
  INV_X2 U7792 ( .A(n8535), .ZN(n8958) );
  NOR2_X1 U7793 ( .A1(n10567), .A2(n7752), .ZN(n7751) );
  INV_X1 U7794 ( .A(n10534), .ZN(n7752) );
  OAI22_X1 U7795 ( .A1(n7423), .A2(n7420), .B1(n13697), .B2(n7426), .ZN(n7419)
         );
  NAND2_X1 U7796 ( .A1(n13729), .A2(n7422), .ZN(n7421) );
  INV_X1 U7797 ( .A(n9279), .ZN(n9285) );
  INV_X1 U7798 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n9276) );
  AND2_X1 U7799 ( .A1(n6881), .A2(n6877), .ZN(n6875) );
  OR2_X1 U7800 ( .A1(n8662), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n8681) );
  AND2_X1 U7801 ( .A1(n11611), .A2(n11601), .ZN(n7605) );
  NAND2_X1 U7802 ( .A1(n11546), .A2(n6687), .ZN(n7619) );
  NAND2_X1 U7803 ( .A1(n14804), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n7653) );
  NAND2_X1 U7804 ( .A1(n7487), .A2(n7484), .ZN(n14473) );
  AOI21_X1 U7805 ( .B1(n7486), .B2(n7490), .A(n7485), .ZN(n7484) );
  NOR2_X1 U7806 ( .A1(n14406), .A2(n14444), .ZN(n7485) );
  AOI21_X1 U7807 ( .B1(n7685), .B2(n7687), .A(n6719), .ZN(n7684) );
  XNOR2_X1 U7808 ( .A(n14499), .B(n12142), .ZN(n14491) );
  XNOR2_X1 U7809 ( .A(n14514), .B(n7177), .ZN(n14503) );
  NAND2_X1 U7810 ( .A1(n14971), .A2(n11449), .ZN(n11461) );
  AND2_X1 U7811 ( .A1(n12131), .A2(n12141), .ZN(n9996) );
  XNOR2_X1 U7812 ( .A(n9125), .B(n9108), .ZN(n14032) );
  OAI21_X1 U7813 ( .B1(n9106), .B2(n9105), .A(n9107), .ZN(n9125) );
  INV_X1 U7814 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n6874) );
  AOI21_X1 U7815 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(n14848), .A(n14847), .ZN(
        n14857) );
  NOR2_X1 U7816 ( .A1(n14859), .A2(n14858), .ZN(n14847) );
  NAND2_X1 U7817 ( .A1(n15252), .A2(n7789), .ZN(n7788) );
  INV_X1 U7818 ( .A(n12217), .ZN(n12622) );
  INV_X1 U7819 ( .A(n7696), .ZN(n11014) );
  NAND2_X1 U7820 ( .A1(n7138), .A2(n11855), .ZN(n6988) );
  NAND2_X1 U7821 ( .A1(n11856), .A2(n15695), .ZN(n7138) );
  NOR2_X1 U7822 ( .A1(n11867), .A2(n7355), .ZN(n7354) );
  INV_X1 U7823 ( .A(n11189), .ZN(n7355) );
  AOI21_X1 U7824 ( .B1(n7830), .B2(n7832), .A(n7827), .ZN(n7826) );
  OAI21_X1 U7825 ( .B1(n7828), .B2(n13101), .A(n13113), .ZN(n7827) );
  INV_X1 U7826 ( .A(n13561), .ZN(n15123) );
  AND2_X1 U7827 ( .A1(n9409), .A2(n14029), .ZN(n15467) );
  OR3_X1 U7828 ( .A1(n6926), .A2(n13636), .A3(n11865), .ZN(n13898) );
  NOR2_X1 U7829 ( .A1(n13637), .A2(n13899), .ZN(n6926) );
  INV_X1 U7830 ( .A(n14694), .ZN(n7133) );
  OR2_X1 U7831 ( .A1(n7794), .A2(n15256), .ZN(n7793) );
  NAND2_X1 U7832 ( .A1(n7796), .A2(n7791), .ZN(n7790) );
  NAND2_X1 U7833 ( .A1(n7169), .A2(n8530), .ZN(n8547) );
  OAI21_X1 U7834 ( .B1(n8531), .B2(n13578), .A(n8529), .ZN(n7170) );
  AOI21_X1 U7835 ( .B1(n11965), .B2(n11964), .A(n11963), .ZN(n11966) );
  MUX2_X1 U7836 ( .A(n11962), .B(n11961), .S(n11960), .Z(n11963) );
  NAND2_X1 U7837 ( .A1(n8570), .A2(n8569), .ZN(n7870) );
  NAND2_X1 U7838 ( .A1(n6888), .A2(n6886), .ZN(n7173) );
  INV_X1 U7839 ( .A(n8585), .ZN(n7149) );
  NAND2_X1 U7840 ( .A1(n7305), .A2(n7304), .ZN(n12001) );
  AOI21_X1 U7841 ( .B1(n6682), .B2(n7308), .A(n6756), .ZN(n7304) );
  NOR2_X1 U7842 ( .A1(n11992), .A2(n7307), .ZN(n7308) );
  NAND2_X1 U7843 ( .A1(n7885), .A2(n8719), .ZN(n7884) );
  NAND2_X1 U7844 ( .A1(n7889), .A2(n7886), .ZN(n7885) );
  OAI21_X1 U7845 ( .B1(n8697), .B2(n7889), .A(n7172), .ZN(n8721) );
  AND2_X1 U7846 ( .A1(n7886), .A2(n8720), .ZN(n7172) );
  INV_X1 U7847 ( .A(n8718), .ZN(n7146) );
  NOR2_X1 U7848 ( .A1(n12009), .A2(n7320), .ZN(n7319) );
  INV_X1 U7849 ( .A(n12009), .ZN(n7318) );
  NAND2_X1 U7850 ( .A1(n12021), .A2(n7772), .ZN(n7770) );
  INV_X1 U7851 ( .A(n12018), .ZN(n7772) );
  NAND2_X1 U7852 ( .A1(n6764), .A2(n12034), .ZN(n7313) );
  NAND2_X1 U7853 ( .A1(n7773), .A2(n12018), .ZN(n7771) );
  INV_X1 U7854 ( .A(n8794), .ZN(n7879) );
  NAND2_X1 U7855 ( .A1(n7297), .A2(n7295), .ZN(n7299) );
  NAND2_X1 U7856 ( .A1(n6708), .A2(n7296), .ZN(n7295) );
  NAND2_X1 U7857 ( .A1(n6891), .A2(n6890), .ZN(n6889) );
  NAND2_X1 U7858 ( .A1(n6893), .A2(n8814), .ZN(n6892) );
  INV_X1 U7859 ( .A(n8815), .ZN(n6890) );
  INV_X1 U7860 ( .A(n12072), .ZN(n7764) );
  INV_X1 U7861 ( .A(n12073), .ZN(n7760) );
  NOR2_X1 U7862 ( .A1(n12073), .A2(n12072), .ZN(n7758) );
  AND2_X1 U7863 ( .A1(n7763), .A2(n12076), .ZN(n7762) );
  NAND2_X1 U7864 ( .A1(n12090), .A2(n7163), .ZN(n7162) );
  INV_X1 U7865 ( .A(n12089), .ZN(n7163) );
  INV_X1 U7866 ( .A(n9013), .ZN(n7882) );
  NAND2_X1 U7867 ( .A1(n6899), .A2(n6896), .ZN(n8991) );
  INV_X1 U7868 ( .A(n8893), .ZN(n7032) );
  AND2_X1 U7869 ( .A1(n9056), .A2(n9057), .ZN(n7877) );
  INV_X1 U7870 ( .A(n9035), .ZN(n7081) );
  NAND2_X1 U7871 ( .A1(n7876), .A2(n7875), .ZN(n7874) );
  INV_X1 U7872 ( .A(n9056), .ZN(n7875) );
  INV_X1 U7873 ( .A(n9057), .ZN(n7876) );
  NOR2_X1 U7874 ( .A1(n7906), .A2(n6725), .ZN(n7905) );
  NAND2_X1 U7875 ( .A1(n12101), .A2(n12100), .ZN(n7785) );
  AND2_X1 U7876 ( .A1(n9107), .A2(SI_26_), .ZN(n7734) );
  NAND2_X1 U7877 ( .A1(n7901), .A2(n7905), .ZN(n7895) );
  AOI21_X1 U7878 ( .B1(n7902), .B2(n7899), .A(n9122), .ZN(n7898) );
  NOR2_X1 U7879 ( .A1(n9123), .A2(n7899), .ZN(n7901) );
  NAND2_X1 U7880 ( .A1(n11952), .A2(n12141), .ZN(n12118) );
  AOI21_X1 U7881 ( .B1(n9105), .B2(n7734), .A(n7733), .ZN(n7732) );
  INV_X1 U7882 ( .A(n9124), .ZN(n7733) );
  AOI21_X1 U7883 ( .B1(n9105), .B2(n9107), .A(SI_26_), .ZN(n7735) );
  INV_X1 U7884 ( .A(n9107), .ZN(n7731) );
  NAND2_X1 U7885 ( .A1(n7732), .A2(n7729), .ZN(n7728) );
  INV_X1 U7886 ( .A(n7734), .ZN(n7729) );
  INV_X1 U7887 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n9304) );
  INV_X1 U7888 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n9303) );
  INV_X1 U7889 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n9302) );
  NOR3_X1 U7890 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .A3(
        P1_IR_REG_16__SCAN_IN), .ZN(n9305) );
  AOI21_X1 U7891 ( .B1(n7030), .B2(n7033), .A(n7028), .ZN(n7027) );
  NAND2_X1 U7892 ( .A1(n8894), .A2(n7030), .ZN(n7029) );
  INV_X1 U7893 ( .A(n8979), .ZN(n7028) );
  AND2_X1 U7894 ( .A1(n7748), .A2(n7013), .ZN(n7012) );
  NAND2_X1 U7895 ( .A1(n7014), .A2(n8797), .ZN(n7013) );
  INV_X1 U7896 ( .A(n7913), .ZN(n7014) );
  NAND2_X1 U7897 ( .A1(n8821), .A2(n14937), .ZN(n8847) );
  INV_X1 U7898 ( .A(n8797), .ZN(n7015) );
  INV_X1 U7899 ( .A(P2_RD_REG_SCAN_IN), .ZN(n7442) );
  INV_X1 U7900 ( .A(n12279), .ZN(n7290) );
  XOR2_X1 U7901 ( .A(n10336), .B(n10337), .Z(n10267) );
  NOR2_X1 U7902 ( .A1(n10261), .A2(n6707), .ZN(n10332) );
  NAND2_X1 U7903 ( .A1(n7326), .A2(n6751), .ZN(n10598) );
  NAND2_X1 U7904 ( .A1(n7695), .A2(n6742), .ZN(n7326) );
  INV_X1 U7905 ( .A(n7693), .ZN(n7325) );
  OR2_X1 U7906 ( .A1(n12693), .A2(n15032), .ZN(n7253) );
  NAND2_X1 U7907 ( .A1(n15048), .A2(n12651), .ZN(n12652) );
  OR2_X1 U7908 ( .A1(n15061), .A2(n12701), .ZN(n7249) );
  INV_X1 U7909 ( .A(n12566), .ZN(n7369) );
  AOI21_X1 U7910 ( .B1(n7389), .B2(n7391), .A(n7387), .ZN(n7386) );
  INV_X1 U7911 ( .A(n12558), .ZN(n7387) );
  OR2_X1 U7912 ( .A1(n12338), .A2(n8324), .ZN(n12558) );
  NAND2_X1 U7913 ( .A1(n7067), .A2(n7069), .ZN(n7065) );
  NOR2_X1 U7914 ( .A1(n8410), .A2(n7071), .ZN(n7070) );
  INV_X1 U7915 ( .A(n8409), .ZN(n7071) );
  AND2_X1 U7916 ( .A1(n12884), .A2(n7411), .ZN(n7410) );
  OR2_X1 U7917 ( .A1(n12628), .A2(n13044), .ZN(n12510) );
  INV_X1 U7918 ( .A(n12489), .ZN(n7857) );
  XNOR2_X1 U7919 ( .A(n15756), .B(n12633), .ZN(n12477) );
  OR2_X1 U7920 ( .A1(n8429), .A2(n8046), .ZN(n8049) );
  OR2_X1 U7921 ( .A1(n12637), .A2(n15690), .ZN(n12444) );
  OR2_X1 U7922 ( .A1(n10318), .A2(n7129), .ZN(n10312) );
  NAND2_X1 U7923 ( .A1(n10318), .A2(n10316), .ZN(n12438) );
  INV_X1 U7924 ( .A(n7371), .ZN(n7370) );
  INV_X1 U7925 ( .A(n7375), .ZN(n7373) );
  NAND2_X1 U7926 ( .A1(n6978), .A2(n9707), .ZN(n6977) );
  INV_X1 U7927 ( .A(n7959), .ZN(n6978) );
  INV_X1 U7928 ( .A(P3_IR_REG_10__SCAN_IN), .ZN(n8165) );
  INV_X1 U7929 ( .A(P3_IR_REG_3__SCAN_IN), .ZN(n7918) );
  INV_X1 U7930 ( .A(P3_IR_REG_7__SCAN_IN), .ZN(n8109) );
  INV_X1 U7931 ( .A(n7943), .ZN(n7534) );
  INV_X1 U7932 ( .A(P3_ADDR_REG_8__SCAN_IN), .ZN(n14836) );
  INV_X1 U7933 ( .A(n13525), .ZN(n7346) );
  NOR2_X1 U7934 ( .A1(n7346), .A2(n13066), .ZN(n7000) );
  INV_X1 U7935 ( .A(n13504), .ZN(n7811) );
  NAND2_X1 U7936 ( .A1(n13062), .A2(n7808), .ZN(n7807) );
  INV_X1 U7937 ( .A(n13064), .ZN(n7808) );
  INV_X1 U7938 ( .A(n13117), .ZN(n7341) );
  INV_X1 U7939 ( .A(n10904), .ZN(n7359) );
  OR2_X1 U7940 ( .A1(n12191), .A2(n7622), .ZN(n7621) );
  INV_X1 U7941 ( .A(n13807), .ZN(n7094) );
  NOR2_X1 U7942 ( .A1(n7644), .A2(n6723), .ZN(n7643) );
  INV_X1 U7943 ( .A(n13649), .ZN(n7206) );
  NOR2_X1 U7944 ( .A1(n8730), .A2(n13266), .ZN(n8786) );
  INV_X1 U7945 ( .A(n7188), .ZN(n7187) );
  OAI21_X1 U7946 ( .B1(n10798), .B2(n7189), .A(n11224), .ZN(n7188) );
  INV_X1 U7947 ( .A(n10986), .ZN(n7189) );
  AND2_X1 U7948 ( .A1(n10993), .A2(n15549), .ZN(n11235) );
  INV_X1 U7949 ( .A(n7632), .ZN(n7631) );
  NOR2_X2 U7950 ( .A1(n15143), .A2(n11491), .ZN(n11499) );
  INV_X1 U7951 ( .A(n10897), .ZN(n10890) );
  INV_X1 U7952 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n8493) );
  INV_X1 U7953 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n6860) );
  AND2_X1 U7954 ( .A1(n7597), .A2(n11730), .ZN(n7593) );
  INV_X1 U7955 ( .A(n7590), .ZN(n6872) );
  AOI21_X1 U7956 ( .B1(n7593), .B2(n7599), .A(n7591), .ZN(n7590) );
  INV_X1 U7957 ( .A(n14049), .ZN(n7591) );
  INV_X1 U7958 ( .A(n14161), .ZN(n7604) );
  NOR2_X1 U7959 ( .A1(n7136), .A2(n7135), .ZN(n7134) );
  NOR2_X1 U7960 ( .A1(n14069), .A2(n11688), .ZN(n7135) );
  INV_X1 U7961 ( .A(n14141), .ZN(n7136) );
  INV_X1 U7962 ( .A(n14804), .ZN(n9620) );
  OR2_X1 U7963 ( .A1(n9920), .A2(n6965), .ZN(n6964) );
  AND2_X1 U7964 ( .A1(n11072), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n6965) );
  NAND2_X1 U7965 ( .A1(n14503), .A2(n14442), .ZN(n7686) );
  INV_X1 U7966 ( .A(n14403), .ZN(n7478) );
  INV_X1 U7967 ( .A(n14432), .ZN(n7678) );
  INV_X1 U7968 ( .A(n14622), .ZN(n7467) );
  NOR2_X1 U7969 ( .A1(n14630), .A2(n14426), .ZN(n7143) );
  AND2_X1 U7970 ( .A1(n6705), .A2(n6680), .ZN(n7472) );
  OAI21_X1 U7971 ( .B1(n14659), .B2(n7663), .A(n14423), .ZN(n7662) );
  INV_X1 U7972 ( .A(n14422), .ZN(n7663) );
  OR2_X1 U7973 ( .A1(n15203), .A2(n14211), .ZN(n14660) );
  NOR2_X1 U7974 ( .A1(n15285), .A2(n15286), .ZN(n7511) );
  NAND2_X1 U7975 ( .A1(n7140), .A2(n10127), .ZN(n10184) );
  NAND2_X1 U7976 ( .A1(n10126), .A2(n7141), .ZN(n7140) );
  AND2_X1 U7977 ( .A1(n14449), .A2(n12168), .ZN(n14463) );
  NAND2_X1 U7978 ( .A1(n15187), .A2(n14098), .ZN(n14974) );
  INV_X1 U7979 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n9316) );
  NAND2_X1 U7980 ( .A1(n9019), .A2(n6788), .ZN(n7718) );
  OAI21_X1 U7981 ( .B1(n8875), .B2(n7726), .A(n7723), .ZN(n8978) );
  INV_X1 U7982 ( .A(SI_18_), .ZN(n8973) );
  NAND2_X1 U7983 ( .A1(n8871), .A2(n13466), .ZN(n8874) );
  AND2_X1 U7984 ( .A1(n8931), .A2(n8878), .ZN(n8929) );
  NAND2_X1 U7985 ( .A1(n7016), .A2(n7018), .ZN(n8770) );
  AOI21_X1 U7986 ( .B1(n8742), .B2(n7019), .A(n6754), .ZN(n7018) );
  OR2_X1 U7987 ( .A1(n9388), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n9392) );
  NAND2_X1 U7988 ( .A1(n7131), .A2(n8600), .ZN(n8617) );
  OAI21_X1 U7989 ( .B1(n9158), .B2(P2_DATAO_REG_1__SCAN_IN), .A(n7148), .ZN(
        n8558) );
  OR2_X1 U7990 ( .A1(n8534), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n7148) );
  INV_X1 U7991 ( .A(P3_ADDR_REG_5__SCAN_IN), .ZN(n14826) );
  NAND2_X1 U7992 ( .A1(n7268), .A2(n6730), .ZN(n7267) );
  XNOR2_X1 U7993 ( .A(n7267), .B(n14826), .ZN(n14868) );
  OAI22_X1 U7994 ( .A1(n14892), .A2(n14830), .B1(P1_ADDR_REG_6__SCAN_IN), .B2(
        n10346), .ZN(n14831) );
  AOI21_X1 U7995 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(n14836), .A(n14835), .ZN(
        n14866) );
  NOR2_X1 U7996 ( .A1(n14898), .A2(n14897), .ZN(n14835) );
  OAI21_X1 U7997 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(n14844), .A(n14843), .ZN(
        n14913) );
  AOI21_X1 U7998 ( .B1(n12238), .B2(n12236), .A(n12269), .ZN(n7281) );
  OR2_X1 U7999 ( .A1(n12215), .A2(n12216), .ZN(n7291) );
  NAND2_X1 U8000 ( .A1(n7554), .A2(n11132), .ZN(n15584) );
  AND2_X1 U8001 ( .A1(n11131), .A2(n7555), .ZN(n7554) );
  INV_X1 U8002 ( .A(n11135), .ZN(n7555) );
  INV_X1 U8003 ( .A(n12345), .ZN(n6825) );
  AND2_X1 U8004 ( .A1(n7566), .A2(n6823), .ZN(n6822) );
  NOR2_X1 U8005 ( .A1(n12261), .A2(n7567), .ZN(n7566) );
  NAND3_X1 U8006 ( .A1(n7578), .A2(n8324), .A3(n7580), .ZN(n12333) );
  NAND2_X1 U8007 ( .A1(n10973), .A2(n10974), .ZN(n11124) );
  OR2_X1 U8008 ( .A1(n15014), .A2(n12199), .ZN(n7565) );
  NAND2_X1 U8009 ( .A1(n7093), .A2(n7091), .ZN(n12601) );
  OR2_X1 U8010 ( .A1(n12595), .A2(n12593), .ZN(n7093) );
  AND4_X1 U8011 ( .A1(n8313), .A2(n8312), .A3(n8311), .A4(n8310), .ZN(n12217)
         );
  AND4_X1 U8012 ( .A1(n8121), .A2(n8120), .A3(n8119), .A4(n8118), .ZN(n11136)
         );
  OAI21_X1 U8013 ( .B1(n10365), .B2(n10524), .A(n10025), .ZN(n10355) );
  OR2_X1 U8014 ( .A1(n10030), .A2(n10029), .ZN(n6936) );
  XNOR2_X1 U8015 ( .A(n10598), .B(n10599), .ZN(n10403) );
  NOR2_X1 U8016 ( .A1(n10403), .A2(n10402), .ZN(n10600) );
  NAND2_X1 U8017 ( .A1(n6938), .A2(n6937), .ZN(n7698) );
  INV_X1 U8018 ( .A(n10603), .ZN(n6937) );
  AOI21_X1 U8019 ( .B1(n15598), .B2(n15595), .A(n11029), .ZN(n11031) );
  NOR2_X1 U8020 ( .A1(n11031), .A2(n11030), .ZN(n12677) );
  XOR2_X1 U8021 ( .A(n12644), .B(n15622), .Z(n15618) );
  AND2_X1 U8022 ( .A1(n6929), .A2(n6928), .ZN(n12659) );
  NAND2_X1 U8023 ( .A1(n15640), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n6928) );
  INV_X1 U8024 ( .A(n15632), .ZN(n6929) );
  OR2_X1 U8025 ( .A1(n15650), .A2(n8190), .ZN(n6927) );
  NAND2_X1 U8026 ( .A1(n7253), .A2(n7252), .ZN(n15036) );
  NAND2_X1 U8027 ( .A1(n12693), .A2(n15032), .ZN(n7252) );
  NOR2_X1 U8028 ( .A1(n15036), .A2(n15037), .ZN(n15035) );
  NAND2_X1 U8029 ( .A1(n15049), .A2(n15050), .ZN(n15048) );
  NOR2_X1 U8030 ( .A1(n15054), .A2(n7690), .ZN(n12663) );
  NOR2_X1 U8031 ( .A1(n15042), .A2(n13407), .ZN(n7690) );
  NOR2_X1 U8032 ( .A1(n15063), .A2(n15062), .ZN(n15061) );
  AND2_X1 U8033 ( .A1(n12586), .A2(n8425), .ZN(n12728) );
  NAND2_X1 U8034 ( .A1(n12738), .A2(n12575), .ZN(n11853) );
  NOR2_X1 U8035 ( .A1(n11853), .A2(n8422), .ZN(n12727) );
  NAND2_X1 U8036 ( .A1(n12752), .A2(n8419), .ZN(n12741) );
  INV_X1 U8037 ( .A(n12753), .ZN(n12757) );
  OAI21_X1 U8038 ( .B1(n12779), .B2(n7369), .A(n7367), .ZN(n12735) );
  NAND2_X1 U8039 ( .A1(n12783), .A2(n7851), .ZN(n12764) );
  NOR2_X1 U8040 ( .A1(n7853), .A2(n7852), .ZN(n7851) );
  INV_X1 U8041 ( .A(n8417), .ZN(n7852) );
  NAND2_X1 U8042 ( .A1(n6986), .A2(n6985), .ZN(n6984) );
  NAND2_X1 U8043 ( .A1(n12779), .A2(n12568), .ZN(n12772) );
  AOI21_X1 U8044 ( .B1(n7053), .B2(n7056), .A(n6737), .ZN(n7051) );
  OR2_X1 U8045 ( .A1(n12781), .A2(n12782), .ZN(n12783) );
  AOI21_X1 U8046 ( .B1(n7055), .B2(n12825), .A(n7054), .ZN(n7053) );
  INV_X1 U8047 ( .A(n12409), .ZN(n7054) );
  INV_X1 U8048 ( .A(n7399), .ZN(n7397) );
  AOI21_X1 U8049 ( .B1(n8278), .B2(n7400), .A(n8291), .ZN(n7399) );
  NOR2_X1 U8050 ( .A1(n12547), .A2(n7401), .ZN(n7400) );
  INV_X1 U8051 ( .A(n12624), .ZN(n12845) );
  OR2_X1 U8052 ( .A1(n12842), .A2(n12846), .ZN(n12840) );
  AND2_X1 U8053 ( .A1(n12536), .A2(n12542), .ZN(n12846) );
  XNOR2_X1 U8054 ( .A(n13032), .B(n12870), .ZN(n12854) );
  AND2_X1 U8055 ( .A1(n12529), .A2(n12524), .ZN(n12884) );
  AOI21_X1 U8056 ( .B1(n6681), .B2(n7063), .A(n6750), .ZN(n7061) );
  NAND2_X1 U8057 ( .A1(n8404), .A2(n8403), .ZN(n12904) );
  AND2_X1 U8058 ( .A1(n8158), .A2(n8157), .ZN(n11416) );
  NAND2_X1 U8059 ( .A1(n11337), .A2(n11341), .ZN(n11411) );
  AOI21_X1 U8060 ( .B1(n7383), .B2(n12483), .A(n7382), .ZN(n7381) );
  INV_X1 U8061 ( .A(n12487), .ZN(n7382) );
  INV_X1 U8062 ( .A(n8115), .ZN(n7383) );
  NAND2_X1 U8063 ( .A1(n6811), .A2(n7384), .ZN(n11143) );
  INV_X1 U8064 ( .A(n12477), .ZN(n6821) );
  NAND2_X1 U8065 ( .A1(n11152), .A2(n6821), .ZN(n11151) );
  NAND2_X1 U8066 ( .A1(n8396), .A2(n10853), .ZN(n10726) );
  AND3_X1 U8067 ( .A1(n8058), .A2(n8057), .A3(n8056), .ZN(n10660) );
  INV_X1 U8068 ( .A(n15695), .ZN(n15708) );
  NAND2_X1 U8069 ( .A1(n8371), .A2(n8370), .ZN(n12582) );
  OR2_X1 U8070 ( .A1(n8066), .A2(n13471), .ZN(n8370) );
  OR2_X1 U8071 ( .A1(n8066), .A2(n11167), .ZN(n8334) );
  NAND2_X1 U8072 ( .A1(n8328), .A2(n8327), .ZN(n12563) );
  OR2_X1 U8073 ( .A1(n8066), .A2(n10969), .ZN(n8327) );
  NAND2_X1 U8074 ( .A1(n8284), .A2(n8283), .ZN(n12411) );
  AND3_X1 U8075 ( .A1(n8142), .A2(n8141), .A3(n8140), .ZN(n11120) );
  NAND2_X1 U8076 ( .A1(n8008), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8009) );
  NAND2_X1 U8077 ( .A1(n8440), .A2(n7077), .ZN(n8008) );
  OAI22_X1 U8078 ( .A1(n8369), .A2(n7989), .B1(P2_DATAO_REG_27__SCAN_IN), .B2(
        n14028), .ZN(n8382) );
  NAND2_X1 U8079 ( .A1(n8440), .A2(n6704), .ZN(n8000) );
  AND2_X1 U8080 ( .A1(n8439), .A2(n8438), .ZN(n8465) );
  MUX2_X1 U8081 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8437), .S(
        P3_IR_REG_26__SCAN_IN), .Z(n8439) );
  NAND2_X1 U8082 ( .A1(n7986), .A2(n7985), .ZN(n8358) );
  AND2_X1 U8083 ( .A1(n7861), .A2(n7860), .ZN(n7859) );
  OR2_X1 U8084 ( .A1(n7975), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n7976) );
  AND2_X1 U8085 ( .A1(n7923), .A2(n7928), .ZN(n8481) );
  XNOR2_X1 U8086 ( .A(n7975), .B(n11860), .ZN(n8292) );
  AOI21_X1 U8087 ( .B1(n7527), .B2(n7969), .A(n7525), .ZN(n7524) );
  INV_X1 U8088 ( .A(n7972), .ZN(n7525) );
  AND2_X1 U8089 ( .A1(n7972), .A2(n7970), .ZN(n8261) );
  NAND2_X1 U8090 ( .A1(P2_DATAO_REG_17__SCAN_IN), .A2(n7532), .ZN(n7531) );
  NAND2_X1 U8091 ( .A1(n7967), .A2(n7966), .ZN(n8237) );
  INV_X1 U8092 ( .A(n7962), .ZN(n7540) );
  NAND2_X1 U8093 ( .A1(n7542), .A2(n8206), .ZN(n7541) );
  INV_X1 U8094 ( .A(n8207), .ZN(n7542) );
  NAND2_X1 U8095 ( .A1(n8182), .A2(n7959), .ZN(n6974) );
  OR2_X1 U8096 ( .A1(n8180), .A2(n8179), .ZN(n8182) );
  AOI21_X1 U8097 ( .B1(n7956), .B2(n6973), .A(n6799), .ZN(n6972) );
  INV_X1 U8098 ( .A(n7954), .ZN(n6973) );
  INV_X1 U8099 ( .A(n7955), .ZN(n6971) );
  INV_X1 U8100 ( .A(n7392), .ZN(n7393) );
  XNOR2_X1 U8101 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .ZN(n8067) );
  INV_X1 U8102 ( .A(P3_IR_REG_1__SCAN_IN), .ZN(n7917) );
  XNOR2_X1 U8103 ( .A(n8040), .B(n7334), .ZN(n10092) );
  OAI21_X1 U8104 ( .B1(P3_IR_REG_0__SCAN_IN), .B2(P3_IR_REG_1__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n7334) );
  AND2_X1 U8105 ( .A1(n9934), .A2(n9694), .ZN(n7817) );
  INV_X1 U8106 ( .A(n13106), .ZN(n7832) );
  XNOR2_X1 U8107 ( .A(n13107), .B(n7362), .ZN(n9693) );
  INV_X1 U8108 ( .A(n10704), .ZN(n7705) );
  OR2_X1 U8109 ( .A1(n9943), .A2(n9944), .ZN(n10160) );
  AND2_X1 U8110 ( .A1(n13578), .A2(n10295), .ZN(n9790) );
  NAND2_X1 U8111 ( .A1(n8981), .A2(n8980), .ZN(n13681) );
  XNOR2_X1 U8112 ( .A(n13107), .B(n6989), .ZN(n9931) );
  INV_X1 U8113 ( .A(n10162), .ZN(n7819) );
  AND2_X1 U8114 ( .A1(n9240), .A2(n9239), .ZN(n7166) );
  INV_X1 U8115 ( .A(n9214), .ZN(n9198) );
  NOR2_X1 U8116 ( .A1(n7621), .A2(n9400), .ZN(n7620) );
  OAI21_X1 U8117 ( .B1(n9432), .B2(P2_REG2_REG_2__SCAN_IN), .A(n6848), .ZN(
        n9428) );
  NAND2_X1 U8118 ( .A1(n9432), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6848) );
  NAND2_X1 U8119 ( .A1(n13696), .A2(n9249), .ZN(n13718) );
  INV_X1 U8120 ( .A(n7628), .ZN(n7626) );
  INV_X1 U8121 ( .A(n13659), .ZN(n7200) );
  NAND2_X1 U8122 ( .A1(n13741), .A2(n13689), .ZN(n13691) );
  NAND2_X1 U8123 ( .A1(n6675), .A2(n13661), .ZN(n7628) );
  NAND2_X1 U8124 ( .A1(n7629), .A2(n6675), .ZN(n7627) );
  NAND2_X1 U8125 ( .A1(n6699), .A2(n13770), .ZN(n13769) );
  NOR2_X1 U8126 ( .A1(n13806), .A2(n6696), .ZN(n7231) );
  XNOR2_X1 U8127 ( .A(n13947), .B(n13685), .ZN(n13800) );
  INV_X1 U8128 ( .A(n7211), .ZN(n7210) );
  NOR2_X1 U8129 ( .A1(n6686), .A2(n7736), .ZN(n7240) );
  INV_X1 U8130 ( .A(n13647), .ZN(n7213) );
  AND2_X1 U8131 ( .A1(n13855), .A2(n7212), .ZN(n7211) );
  NAND2_X1 U8132 ( .A1(n7213), .A2(n13648), .ZN(n7212) );
  OAI21_X1 U8133 ( .B1(n7429), .B2(n6793), .A(n7737), .ZN(n13861) );
  OR2_X1 U8134 ( .A1(n13985), .A2(n13671), .ZN(n7737) );
  INV_X1 U8135 ( .A(n13875), .ZN(n7429) );
  NAND2_X1 U8136 ( .A1(n13881), .A2(n13646), .ZN(n13860) );
  AOI21_X1 U8137 ( .B1(n7217), .B2(n7219), .A(n7216), .ZN(n7215) );
  OR2_X1 U8138 ( .A1(n13879), .A2(n13880), .ZN(n13881) );
  NAND2_X1 U8139 ( .A1(n13669), .A2(n13668), .ZN(n13875) );
  OR2_X1 U8140 ( .A1(n13991), .A2(n13667), .ZN(n13668) );
  OR2_X1 U8141 ( .A1(n8830), .A2(n8829), .ZN(n8858) );
  INV_X1 U8142 ( .A(n6678), .ZN(n7219) );
  NAND2_X1 U8143 ( .A1(n7246), .A2(n7245), .ZN(n11529) );
  AND2_X1 U8144 ( .A1(n11493), .A2(n6715), .ZN(n7245) );
  NOR2_X1 U8145 ( .A1(n11486), .A2(n7223), .ZN(n7222) );
  INV_X1 U8146 ( .A(n11322), .ZN(n7223) );
  OR2_X1 U8147 ( .A1(n15140), .A2(n11327), .ZN(n7702) );
  NAND2_X1 U8148 ( .A1(n15142), .A2(n11321), .ZN(n7637) );
  AOI21_X1 U8149 ( .B1(n11326), .B2(n11325), .A(n6795), .ZN(n15133) );
  OR2_X1 U8150 ( .A1(n11227), .A2(n11325), .ZN(n11320) );
  NAND2_X1 U8151 ( .A1(n7646), .A2(n7645), .ZN(n10789) );
  AOI21_X1 U8152 ( .B1(n7647), .B2(n10785), .A(n6724), .ZN(n7645) );
  NAND2_X1 U8153 ( .A1(n10789), .A2(n10798), .ZN(n10987) );
  NOR2_X2 U8154 ( .A1(n10891), .A2(n15538), .ZN(n10993) );
  INV_X1 U8155 ( .A(n10788), .ZN(n10798) );
  INV_X1 U8156 ( .A(n10243), .ZN(n7754) );
  NAND2_X1 U8157 ( .A1(n10536), .A2(n7434), .ZN(n10567) );
  NAND2_X1 U8158 ( .A1(n7435), .A2(n13572), .ZN(n7434) );
  NAND2_X1 U8159 ( .A1(n10242), .A2(n7705), .ZN(n10237) );
  OR2_X1 U8160 ( .A1(n9965), .A2(n10704), .ZN(n10248) );
  NAND2_X1 U8161 ( .A1(n9964), .A2(n10239), .ZN(n10238) );
  NAND2_X1 U8162 ( .A1(n9909), .A2(n10556), .ZN(n9965) );
  XNOR2_X1 U8163 ( .A(n13575), .B(n10556), .ZN(n9956) );
  INV_X1 U8164 ( .A(n15522), .ZN(n15551) );
  NAND2_X1 U8165 ( .A1(n9279), .A2(n7908), .ZN(n8503) );
  NAND2_X1 U8166 ( .A1(n6917), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8514) );
  INV_X1 U8167 ( .A(n10920), .ZN(n6867) );
  NOR2_X1 U8168 ( .A1(n7607), .A2(n10929), .ZN(n6870) );
  NAND2_X1 U8169 ( .A1(n14807), .A2(n6712), .ZN(n7778) );
  OR2_X1 U8170 ( .A1(n14194), .A2(n11802), .ZN(n7587) );
  NAND2_X1 U8171 ( .A1(n11273), .A2(n11272), .ZN(n11355) );
  INV_X1 U8172 ( .A(n11275), .ZN(n11273) );
  AND2_X1 U8173 ( .A1(n9817), .A2(n9616), .ZN(n10128) );
  NAND2_X1 U8174 ( .A1(n11695), .A2(n11694), .ZN(n7603) );
  OAI21_X1 U8175 ( .B1(n7605), .B2(n6865), .A(n7612), .ZN(n6864) );
  NAND2_X1 U8176 ( .A1(n7614), .A2(n7613), .ZN(n7612) );
  INV_X1 U8177 ( .A(n14205), .ZN(n7613) );
  NAND2_X1 U8178 ( .A1(n14152), .A2(n14151), .ZN(n7606) );
  NAND2_X1 U8179 ( .A1(n14059), .A2(n10687), .ZN(n10924) );
  NAND2_X1 U8180 ( .A1(n6861), .A2(n7615), .ZN(n11544) );
  AOI21_X1 U8181 ( .B1(n7616), .B2(n11276), .A(n6744), .ZN(n7615) );
  NAND2_X1 U8182 ( .A1(n11275), .A2(n7616), .ZN(n6861) );
  NAND2_X1 U8183 ( .A1(n7598), .A2(n7604), .ZN(n7597) );
  INV_X1 U8184 ( .A(n7600), .ZN(n7598) );
  AOI21_X1 U8185 ( .B1(n7601), .B2(n7602), .A(n11713), .ZN(n7600) );
  INV_X1 U8186 ( .A(n11694), .ZN(n7601) );
  NAND2_X1 U8187 ( .A1(n14183), .A2(n7134), .ZN(n11695) );
  NAND2_X1 U8188 ( .A1(n7603), .A2(n7602), .ZN(n14163) );
  AND2_X1 U8189 ( .A1(n14174), .A2(n11577), .ZN(n7618) );
  NAND2_X1 U8190 ( .A1(n14122), .A2(n11655), .ZN(n14183) );
  NAND2_X1 U8191 ( .A1(n14679), .A2(n6663), .ZN(n7144) );
  INV_X1 U8192 ( .A(n12173), .ZN(n7106) );
  NAND2_X1 U8193 ( .A1(n6951), .A2(n6950), .ZN(n14254) );
  OR2_X1 U8194 ( .A1(n14258), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6950) );
  NAND2_X1 U8195 ( .A1(n14258), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6951) );
  NOR2_X1 U8196 ( .A1(n14255), .A2(n14254), .ZN(n14253) );
  NOR2_X1 U8197 ( .A1(n9339), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n9370) );
  OR2_X1 U8198 ( .A1(n9713), .A2(n6784), .ZN(n6960) );
  OR2_X1 U8199 ( .A1(n6960), .A2(n6959), .ZN(n14295) );
  INV_X1 U8200 ( .A(n14297), .ZN(n6959) );
  NOR2_X1 U8201 ( .A1(n11216), .A2(n11217), .ZN(n11219) );
  NAND2_X1 U8202 ( .A1(n11219), .A2(n11218), .ZN(n14352) );
  XNOR2_X1 U8203 ( .A(n14368), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n6946) );
  INV_X1 U8204 ( .A(n14463), .ZN(n14454) );
  NAND2_X1 U8205 ( .A1(n14488), .A2(n14491), .ZN(n7034) );
  INV_X1 U8206 ( .A(n7520), .ZN(n14489) );
  INV_X1 U8207 ( .A(n7686), .ZN(n7687) );
  NAND2_X1 U8208 ( .A1(n14732), .A2(n14441), .ZN(n14524) );
  INV_X1 U8209 ( .A(n7685), .ZN(n14441) );
  NOR2_X1 U8210 ( .A1(n14586), .A2(n14743), .ZN(n14556) );
  NAND2_X1 U8211 ( .A1(n14556), .A2(n14559), .ZN(n14555) );
  INV_X1 U8212 ( .A(n14397), .ZN(n7469) );
  INV_X1 U8213 ( .A(n14428), .ZN(n7679) );
  NAND2_X1 U8214 ( .A1(n14623), .A2(n14622), .ZN(n14621) );
  NAND2_X1 U8215 ( .A1(n15205), .A2(n14420), .ZN(n14656) );
  NAND2_X1 U8216 ( .A1(n7664), .A2(n14659), .ZN(n14658) );
  INV_X1 U8217 ( .A(n14656), .ZN(n7664) );
  NAND2_X1 U8218 ( .A1(n7476), .A2(n7475), .ZN(n7474) );
  INV_X1 U8219 ( .A(n14660), .ZN(n7475) );
  NAND2_X1 U8220 ( .A1(n14970), .A2(n12162), .ZN(n7659) );
  NAND2_X1 U8221 ( .A1(n7511), .A2(n7510), .ZN(n15186) );
  INV_X1 U8222 ( .A(n15380), .ZN(n7510) );
  AND2_X1 U8223 ( .A1(n11280), .A2(n11083), .ZN(n11099) );
  NAND2_X1 U8224 ( .A1(n15360), .A2(n7507), .ZN(n15273) );
  AND2_X1 U8225 ( .A1(n15276), .A2(n11097), .ZN(n7507) );
  OAI21_X1 U8226 ( .B1(n10740), .B2(n10739), .A(n10741), .ZN(n10845) );
  NOR2_X1 U8227 ( .A1(n10759), .A2(n10758), .ZN(n7674) );
  CLKBUF_X1 U8228 ( .A(n10584), .Z(n7139) );
  NAND2_X1 U8229 ( .A1(n10451), .A2(n10192), .ZN(n10592) );
  XNOR2_X1 U8230 ( .A(n14227), .B(n10194), .ZN(n11976) );
  NOR2_X1 U8231 ( .A1(n14230), .A2(n10225), .ZN(n11953) );
  OAI21_X1 U8232 ( .B1(n14519), .B2(n7491), .A(n7490), .ZN(n14492) );
  OR2_X2 U8233 ( .A1(n14540), .A2(n14539), .ZN(n14732) );
  NAND2_X1 U8234 ( .A1(n14567), .A2(n14402), .ZN(n14560) );
  INV_X1 U8235 ( .A(n15320), .ZN(n15288) );
  INV_X1 U8236 ( .A(n15379), .ZN(n15366) );
  XNOR2_X1 U8237 ( .A(n9161), .B(n9160), .ZN(n14017) );
  NAND2_X1 U8238 ( .A1(n9169), .A2(n9157), .ZN(n9161) );
  NAND2_X1 U8239 ( .A1(n14795), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9558) );
  NAND2_X1 U8240 ( .A1(n9317), .A2(n9316), .ZN(n9457) );
  INV_X1 U8241 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n9466) );
  INV_X1 U8242 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n7617) );
  NAND2_X1 U8243 ( .A1(n7020), .A2(n8726), .ZN(n8743) );
  NAND2_X1 U8244 ( .A1(n8724), .A2(n8723), .ZN(n7020) );
  XNOR2_X1 U8245 ( .A(n7184), .B(n6703), .ZN(n10828) );
  AOI21_X1 U8246 ( .B1(n7174), .B2(n8678), .A(n6688), .ZN(n7184) );
  NAND2_X1 U8247 ( .A1(n7418), .A2(n6695), .ZN(n7413) );
  INV_X1 U8248 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n7588) );
  INV_X1 U8249 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n6953) );
  INV_X1 U8250 ( .A(n7803), .ZN(n14872) );
  OR2_X1 U8251 ( .A1(n15803), .A2(n14879), .ZN(n6836) );
  NAND2_X1 U8252 ( .A1(n14885), .A2(n15789), .ZN(n14888) );
  NOR2_X1 U8253 ( .A1(n14933), .A2(n14894), .ZN(n14896) );
  INV_X1 U8254 ( .A(n14902), .ZN(n7262) );
  INV_X1 U8255 ( .A(n7800), .ZN(n14899) );
  AND2_X1 U8256 ( .A1(n14901), .A2(n7262), .ZN(n7258) );
  AOI21_X1 U8257 ( .B1(n14840), .B2(n14839), .A(n14838), .ZN(n14908) );
  OAI21_X1 U8258 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(n14850), .A(n14849), .ZN(
        n14917) );
  AND2_X1 U8259 ( .A1(n7792), .A2(n15256), .ZN(n7789) );
  NAND2_X1 U8260 ( .A1(n7265), .A2(n14988), .ZN(n14996) );
  OAI21_X1 U8261 ( .B1(n14989), .B2(n14990), .A(n7266), .ZN(n7265) );
  INV_X1 U8262 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n7266) );
  XNOR2_X1 U8263 ( .A(n6830), .B(n12238), .ZN(n12239) );
  NAND2_X1 U8264 ( .A1(n12353), .A2(n12237), .ZN(n6830) );
  NAND2_X1 U8265 ( .A1(n12354), .A2(n12355), .ZN(n12353) );
  NOR2_X1 U8266 ( .A1(n10465), .A2(n10319), .ZN(n10324) );
  NAND2_X1 U8267 ( .A1(n7576), .A2(n12204), .ZN(n15003) );
  NAND2_X1 U8268 ( .A1(n12202), .A2(n6781), .ZN(n7576) );
  AOI21_X1 U8269 ( .B1(n6674), .B2(n7574), .A(n6792), .ZN(n7573) );
  NAND2_X1 U8270 ( .A1(n12365), .A2(n6674), .ZN(n6831) );
  INV_X1 U8271 ( .A(n6781), .ZN(n7574) );
  NAND2_X1 U8272 ( .A1(n12292), .A2(n12197), .ZN(n15016) );
  NAND2_X1 U8273 ( .A1(n9875), .A2(n12610), .ZN(n15585) );
  AND2_X1 U8274 ( .A1(n9868), .A2(n9323), .ZN(n12610) );
  NAND2_X1 U8275 ( .A1(n11015), .A2(n6933), .ZN(n6932) );
  OR2_X1 U8276 ( .A1(n15601), .A2(n6931), .ZN(n6930) );
  INV_X1 U8277 ( .A(n11016), .ZN(n6933) );
  XNOR2_X1 U8278 ( .A(n12661), .B(n15032), .ZN(n15026) );
  INV_X1 U8279 ( .A(n12709), .ZN(n15679) );
  NAND2_X1 U8280 ( .A1(n15074), .A2(n7086), .ZN(n7085) );
  OR2_X1 U8281 ( .A1(n15073), .A2(n13425), .ZN(n7086) );
  XNOR2_X1 U8282 ( .A(n7257), .B(n12704), .ZN(n7256) );
  NAND2_X1 U8283 ( .A1(n15077), .A2(n12703), .ZN(n7257) );
  OR2_X1 U8284 ( .A1(n12705), .A2(n7255), .ZN(n7254) );
  AND2_X1 U8285 ( .A1(n15604), .A2(n12706), .ZN(n7255) );
  AOI21_X1 U8286 ( .B1(P3_REG2_REG_18__SCAN_IN), .B2(n14948), .A(n15084), .ZN(
        n12667) );
  AND2_X1 U8287 ( .A1(n10034), .A2(n10024), .ZN(n15082) );
  AND2_X1 U8288 ( .A1(n12820), .A2(n12819), .ZN(n12957) );
  NAND2_X1 U8289 ( .A1(n7374), .A2(n12463), .ZN(n11049) );
  NAND2_X1 U8290 ( .A1(n10724), .A2(n12462), .ZN(n7374) );
  AND2_X1 U8291 ( .A1(n11920), .A2(n12394), .ZN(n7544) );
  NAND2_X1 U8292 ( .A1(n7043), .A2(n15695), .ZN(n7849) );
  XNOR2_X1 U8293 ( .A(n7044), .B(n6713), .ZN(n7043) );
  NAND2_X1 U8294 ( .A1(n7046), .A2(n7045), .ZN(n7044) );
  NAND2_X1 U8295 ( .A1(n8426), .A2(n12245), .ZN(n7045) );
  AND2_X1 U8296 ( .A1(n7850), .A2(n8435), .ZN(n7848) );
  INV_X1 U8297 ( .A(n11942), .ZN(n7846) );
  INV_X1 U8298 ( .A(n12582), .ZN(n12996) );
  NAND2_X1 U8299 ( .A1(n12927), .A2(n12926), .ZN(n12994) );
  AND2_X1 U8300 ( .A1(n8307), .A2(n8306), .ZN(n13018) );
  NAND2_X1 U8301 ( .A1(n8228), .A2(n8227), .ZN(n13040) );
  INV_X1 U8302 ( .A(n11120), .ZN(n11403) );
  AND2_X1 U8303 ( .A1(n7077), .A2(n7076), .ZN(n7075) );
  INV_X1 U8304 ( .A(P3_IR_REG_29__SCAN_IN), .ZN(n7076) );
  NAND2_X1 U8305 ( .A1(n9649), .A2(n9287), .ZN(n9398) );
  NAND2_X1 U8306 ( .A1(n9128), .A2(n9127), .ZN(n13912) );
  AOI21_X1 U8307 ( .B1(n7836), .B2(n7835), .A(n7834), .ZN(n7833) );
  INV_X1 U8308 ( .A(n13078), .ZN(n7834) );
  INV_X1 U8309 ( .A(n13494), .ZN(n7835) );
  AND2_X1 U8310 ( .A1(n15122), .A2(n6716), .ZN(n7352) );
  NAND2_X1 U8311 ( .A1(n13679), .A2(n11865), .ZN(n6992) );
  AND2_X1 U8312 ( .A1(n7826), .A2(n7831), .ZN(n7822) );
  NAND2_X1 U8313 ( .A1(n7829), .A2(n13106), .ZN(n7828) );
  INV_X1 U8314 ( .A(n13114), .ZN(n7829) );
  INV_X1 U8315 ( .A(n13116), .ZN(n7824) );
  XNOR2_X1 U8316 ( .A(n9693), .B(n9692), .ZN(n9648) );
  NAND2_X1 U8317 ( .A1(n9065), .A2(n9064), .ZN(n13935) );
  NAND2_X1 U8318 ( .A1(n9790), .A2(n11865), .ZN(n9685) );
  NAND2_X1 U8319 ( .A1(n8935), .A2(n8934), .ZN(n13845) );
  OR2_X1 U8320 ( .A1(n9677), .A2(n9669), .ZN(n13561) );
  NAND2_X1 U8321 ( .A1(n9220), .A2(n9219), .ZN(n13702) );
  NAND2_X1 U8322 ( .A1(n6844), .A2(n9479), .ZN(n13582) );
  OR2_X1 U8323 ( .A1(n15441), .A2(n13579), .ZN(n6844) );
  XNOR2_X1 U8324 ( .A(n13613), .B(n13618), .ZN(n11197) );
  INV_X1 U8325 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n8003) );
  OAI21_X1 U8326 ( .B1(n13623), .B2(n15442), .A(n6855), .ZN(n6854) );
  AOI21_X1 U8327 ( .B1(n13624), .B2(n15467), .A(n15453), .ZN(n6855) );
  NAND2_X1 U8328 ( .A1(n8828), .A2(n8827), .ZN(n15127) );
  NOR2_X1 U8329 ( .A1(n7198), .A2(n6789), .ZN(n7197) );
  NOR2_X1 U8330 ( .A1(n7193), .A2(n13998), .ZN(n7192) );
  NAND2_X1 U8331 ( .A1(n15573), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n7740) );
  INV_X1 U8332 ( .A(n6925), .ZN(n6924) );
  NAND2_X1 U8333 ( .A1(n9279), .A2(n7639), .ZN(n8505) );
  AND2_X1 U8334 ( .A1(n7908), .A2(n7117), .ZN(n7639) );
  AND2_X1 U8335 ( .A1(n13366), .A2(n14018), .ZN(n7002) );
  NOR2_X1 U8336 ( .A1(n13366), .A2(n14018), .ZN(n7003) );
  NAND2_X1 U8337 ( .A1(n10678), .A2(n10677), .ZN(n14058) );
  NOR2_X1 U8338 ( .A1(n11684), .A2(n11683), .ZN(n14606) );
  INV_X1 U8339 ( .A(n14749), .ZN(n14400) );
  NAND2_X1 U8340 ( .A1(n11448), .A2(n11447), .ZN(n15216) );
  INV_X1 U8341 ( .A(n15167), .ZN(n14195) );
  NAND2_X1 U8342 ( .A1(n11616), .A2(n11615), .ZN(n14672) );
  OR2_X1 U8343 ( .A1(n12175), .A2(n12174), .ZN(n7119) );
  NOR2_X1 U8344 ( .A1(n9889), .A2(n9888), .ZN(n14313) );
  NOR2_X1 U8345 ( .A1(n9717), .A2(n9718), .ZN(n14329) );
  INV_X1 U8346 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n8002) );
  NAND2_X1 U8347 ( .A1(n6942), .A2(n14378), .ZN(n6941) );
  INV_X1 U8348 ( .A(n6946), .ZN(n6942) );
  AOI21_X1 U8349 ( .B1(n14376), .B2(n14377), .A(n14612), .ZN(n6940) );
  NAND2_X1 U8350 ( .A1(n6946), .A2(n14378), .ZN(n6945) );
  NOR2_X1 U8351 ( .A1(n14375), .A2(n7108), .ZN(n6944) );
  NAND2_X1 U8352 ( .A1(n11788), .A2(n11787), .ZN(n14499) );
  NAND2_X1 U8353 ( .A1(n11770), .A2(n11769), .ZN(n14514) );
  NAND2_X1 U8354 ( .A1(n14818), .A2(n9817), .ZN(n14559) );
  NAND2_X1 U8355 ( .A1(n14576), .A2(n14437), .ZN(n14554) );
  INV_X1 U8356 ( .A(n15297), .ZN(n15282) );
  NOR2_X1 U8357 ( .A1(n7026), .A2(n15219), .ZN(n7024) );
  AOI21_X1 U8358 ( .B1(n14691), .B2(n15403), .A(n6809), .ZN(n7022) );
  INV_X1 U8359 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n7125) );
  AND2_X1 U8360 ( .A1(n7456), .A2(n7460), .ZN(n7455) );
  INV_X1 U8361 ( .A(n7459), .ZN(n7457) );
  XNOR2_X1 U8362 ( .A(n14451), .B(n7463), .ZN(n14692) );
  NAND2_X1 U8363 ( .A1(n14696), .A2(n14449), .ZN(n14451) );
  INV_X1 U8364 ( .A(n14881), .ZN(n6835) );
  XNOR2_X1 U8365 ( .A(n14896), .B(n13585), .ZN(n15797) );
  OR2_X1 U8366 ( .A1(n15797), .A2(n15798), .ZN(n7801) );
  XNOR2_X1 U8367 ( .A(n7800), .B(n14900), .ZN(n14943) );
  NAND2_X1 U8368 ( .A1(n14943), .A2(n9484), .ZN(n14942) );
  OR2_X1 U8369 ( .A1(n15253), .A2(n7798), .ZN(n7792) );
  AND2_X1 U8370 ( .A1(n15253), .A2(n7798), .ZN(n7794) );
  OAI21_X1 U8371 ( .B1(n15248), .B2(n15249), .A(n7274), .ZN(n7273) );
  INV_X1 U8372 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n7274) );
  OAI21_X1 U8373 ( .B1(n14996), .B2(n14997), .A(n11198), .ZN(n6843) );
  NAND2_X1 U8374 ( .A1(n8565), .A2(n13576), .ZN(n6887) );
  INV_X1 U8375 ( .A(n8569), .ZN(n6886) );
  AOI22_X1 U8376 ( .A1(n9222), .A2(n10543), .B1(n13573), .B2(n9199), .ZN(n8627) );
  NAND2_X1 U8377 ( .A1(n7111), .A2(n7110), .ZN(n7109) );
  INV_X1 U8378 ( .A(n8586), .ZN(n7110) );
  INV_X1 U8379 ( .A(n8627), .ZN(n7893) );
  NAND2_X1 U8380 ( .A1(n11989), .A2(n11991), .ZN(n7769) );
  NAND2_X1 U8381 ( .A1(n11992), .A2(n7307), .ZN(n7306) );
  NAND2_X1 U8382 ( .A1(n12007), .A2(n7767), .ZN(n7766) );
  INV_X1 U8383 ( .A(n12010), .ZN(n7320) );
  AND2_X1 U8384 ( .A1(n8738), .A2(n8739), .ZN(n7907) );
  AND2_X1 U8385 ( .A1(n7313), .A2(n12035), .ZN(n7312) );
  NAND2_X1 U8386 ( .A1(n6895), .A2(n7878), .ZN(n6894) );
  NAND2_X1 U8387 ( .A1(n7880), .A2(n7879), .ZN(n7878) );
  INV_X1 U8388 ( .A(n8795), .ZN(n7880) );
  INV_X1 U8389 ( .A(n7300), .ZN(n7296) );
  AND2_X1 U8390 ( .A1(n14397), .A2(n12053), .ZN(n7303) );
  NAND2_X1 U8391 ( .A1(n6894), .A2(n8815), .ZN(n6893) );
  INV_X1 U8392 ( .A(n6894), .ZN(n6891) );
  MUX2_X1 U8393 ( .A(n14440), .B(n14730), .S(n12117), .Z(n12076) );
  AOI21_X1 U8394 ( .B1(n7757), .B2(n7759), .A(n6759), .ZN(n7321) );
  NOR2_X1 U8395 ( .A1(n7764), .A2(n7760), .ZN(n7759) );
  NAND2_X1 U8396 ( .A1(n6883), .A2(n6882), .ZN(n8947) );
  AOI21_X1 U8397 ( .B1(n8844), .B2(n6884), .A(n8928), .ZN(n6883) );
  NAND2_X1 U8398 ( .A1(n8841), .A2(n6733), .ZN(n6882) );
  INV_X1 U8399 ( .A(n8970), .ZN(n6900) );
  NAND2_X1 U8400 ( .A1(n12091), .A2(n12089), .ZN(n7756) );
  INV_X1 U8401 ( .A(n9012), .ZN(n7881) );
  INV_X1 U8402 ( .A(n9103), .ZN(n7906) );
  AND2_X1 U8403 ( .A1(n9080), .A2(n7872), .ZN(n7871) );
  INV_X1 U8404 ( .A(n10567), .ZN(n10535) );
  INV_X1 U8405 ( .A(n10237), .ZN(n7636) );
  AND2_X1 U8406 ( .A1(n7720), .A2(n7031), .ZN(n7030) );
  AND2_X1 U8407 ( .A1(n7721), .A2(n8977), .ZN(n7720) );
  NAND2_X1 U8408 ( .A1(n7722), .A2(n7032), .ZN(n7031) );
  INV_X1 U8409 ( .A(n7722), .ZN(n7033) );
  NAND2_X1 U8410 ( .A1(n10401), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n7693) );
  INV_X1 U8411 ( .A(n10400), .ZN(n7327) );
  INV_X1 U8412 ( .A(n12555), .ZN(n7391) );
  INV_X1 U8413 ( .A(n7390), .ZN(n7389) );
  OAI21_X1 U8414 ( .B1(n12554), .B2(n7391), .A(n12559), .ZN(n7390) );
  NAND2_X1 U8415 ( .A1(n8425), .A2(n12725), .ZN(n12584) );
  INV_X1 U8416 ( .A(n12584), .ZN(n7405) );
  OAI21_X1 U8417 ( .B1(n12462), .B2(n7376), .A(n12412), .ZN(n7375) );
  NOR2_X1 U8418 ( .A1(P3_IR_REG_25__SCAN_IN), .A2(P3_IR_REG_26__SCAN_IN), .ZN(
        n7868) );
  INV_X1 U8419 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n13360) );
  INV_X1 U8420 ( .A(n14491), .ZN(n7489) );
  NAND2_X1 U8421 ( .A1(n14514), .A2(n7177), .ZN(n7495) );
  NAND2_X1 U8422 ( .A1(n14579), .A2(n14437), .ZN(n7667) );
  AND2_X1 U8423 ( .A1(n7781), .A2(n9311), .ZN(n7503) );
  AND2_X1 U8424 ( .A1(n7716), .A2(n9038), .ZN(n7714) );
  INV_X1 U8425 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n7781) );
  INV_X1 U8426 ( .A(n8820), .ZN(n7749) );
  INV_X1 U8427 ( .A(n8847), .ZN(n7747) );
  NAND2_X1 U8428 ( .A1(n7012), .A2(n7015), .ZN(n7010) );
  NAND2_X1 U8429 ( .A1(n8848), .A2(n9561), .ZN(n8869) );
  NOR2_X1 U8430 ( .A1(n8741), .A2(n8722), .ZN(n7017) );
  INV_X1 U8431 ( .A(n8726), .ZN(n7019) );
  INV_X1 U8432 ( .A(n7713), .ZN(n7712) );
  OAI21_X1 U8433 ( .B1(n8678), .B2(n6688), .A(n6703), .ZN(n7713) );
  OAI21_X1 U8434 ( .B1(n9616), .B2(n7179), .A(n7178), .ZN(n8618) );
  NAND2_X1 U8435 ( .A1(n9616), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n7178) );
  NAND2_X1 U8436 ( .A1(n12333), .A2(n7580), .ZN(n6833) );
  INV_X1 U8437 ( .A(n12211), .ZN(n7567) );
  NAND2_X1 U8438 ( .A1(n12345), .A2(n6824), .ZN(n6823) );
  INV_X1 U8439 ( .A(n12208), .ZN(n6824) );
  INV_X1 U8440 ( .A(n8308), .ZN(n8318) );
  INV_X1 U8441 ( .A(n7092), .ZN(n7091) );
  OAI21_X1 U8442 ( .B1(n12594), .B2(n12585), .A(n12597), .ZN(n7092) );
  NAND2_X1 U8443 ( .A1(n6936), .A2(n10028), .ZN(n10094) );
  NAND2_X1 U8444 ( .A1(n10110), .A2(n10094), .ZN(n10095) );
  NAND2_X1 U8445 ( .A1(n10266), .A2(n10265), .ZN(n10336) );
  NAND2_X1 U8446 ( .A1(n12643), .A2(n12642), .ZN(n12644) );
  NAND2_X1 U8447 ( .A1(n12690), .A2(n15669), .ZN(n12649) );
  INV_X1 U8448 ( .A(n7053), .ZN(n7052) );
  AOI21_X1 U8449 ( .B1(n12846), .B2(n8413), .A(n6743), .ZN(n7866) );
  INV_X1 U8450 ( .A(n8413), .ZN(n7864) );
  INV_X1 U8451 ( .A(n12536), .ZN(n7401) );
  OR2_X1 U8452 ( .A1(n8403), .A2(n7063), .ZN(n7062) );
  INV_X1 U8453 ( .A(n8405), .ZN(n7063) );
  INV_X1 U8454 ( .A(n8400), .ZN(n7049) );
  INV_X1 U8455 ( .A(n12492), .ZN(n7380) );
  NAND2_X1 U8456 ( .A1(n8394), .A2(n15732), .ZN(n12453) );
  INV_X1 U8457 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n7040) );
  AND2_X1 U8458 ( .A1(n7861), .A2(n7919), .ZN(n7858) );
  OR2_X1 U8459 ( .A1(n8183), .A2(P3_IR_REG_11__SCAN_IN), .ZN(n8197) );
  INV_X1 U8460 ( .A(P3_IR_REG_8__SCAN_IN), .ZN(n7248) );
  NAND4_X1 U8461 ( .A1(n8040), .A2(n7917), .A3(n7036), .A4(n7035), .ZN(n7038)
         );
  INV_X1 U8462 ( .A(P3_IR_REG_6__SCAN_IN), .ZN(n7035) );
  OR2_X1 U8463 ( .A1(n8108), .A2(P3_IR_REG_6__SCAN_IN), .ZN(n8122) );
  NOR2_X1 U8464 ( .A1(n7339), .A2(n7342), .ZN(n7336) );
  AOI21_X1 U8466 ( .B1(n9104), .B2(n7897), .A(n7894), .ZN(n9206) );
  OR2_X1 U8467 ( .A1(n7898), .A2(n7901), .ZN(n7897) );
  NAND2_X1 U8468 ( .A1(n7896), .A2(n7895), .ZN(n7894) );
  INV_X1 U8469 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n8608) );
  NOR2_X1 U8470 ( .A1(n13730), .A2(n13905), .ZN(n7446) );
  INV_X1 U8471 ( .A(n13912), .ZN(n13695) );
  NOR3_X1 U8472 ( .A1(n13810), .A2(n13935), .A3(n6921), .ZN(n7450) );
  OR2_X1 U8473 ( .A1(n13942), .A2(n13947), .ZN(n6921) );
  NOR2_X1 U8474 ( .A1(n13821), .A2(n13681), .ZN(n7151) );
  NOR2_X1 U8475 ( .A1(n7744), .A2(n7440), .ZN(n7439) );
  INV_X1 U8476 ( .A(n13677), .ZN(n7440) );
  NOR2_X1 U8477 ( .A1(n7745), .A2(n13965), .ZN(n7744) );
  NOR2_X1 U8478 ( .A1(n8858), .A2(n8857), .ZN(n8882) );
  AND2_X1 U8479 ( .A1(n8786), .A2(n8785), .ZN(n8804) );
  NOR2_X1 U8480 ( .A1(n13697), .A2(n7423), .ZN(n7422) );
  AOI21_X1 U8481 ( .B1(n7699), .B2(n13737), .A(n7427), .ZN(n7426) );
  INV_X1 U8482 ( .A(n13696), .ZN(n7427) );
  INV_X1 U8483 ( .A(n7426), .ZN(n7423) );
  NOR2_X1 U8484 ( .A1(n7699), .A2(n13697), .ZN(n7420) );
  INV_X1 U8485 ( .A(n7446), .ZN(n13720) );
  INV_X1 U8486 ( .A(n13660), .ZN(n13497) );
  NAND2_X1 U8487 ( .A1(n7235), .A2(n10795), .ZN(n10898) );
  NAND2_X1 U8488 ( .A1(n10792), .A2(n10791), .ZN(n7235) );
  INV_X1 U8489 ( .A(n7335), .ZN(n9641) );
  NAND2_X1 U8490 ( .A1(n9173), .A2(n7335), .ZN(n9639) );
  INV_X1 U8491 ( .A(n11619), .ZN(n7614) );
  NAND2_X1 U8492 ( .A1(n11956), .A2(n9630), .ZN(n11722) );
  NAND2_X1 U8493 ( .A1(n12140), .A2(n11952), .ZN(n7323) );
  NAND2_X1 U8494 ( .A1(n12107), .A2(n12108), .ZN(n7099) );
  NAND2_X1 U8495 ( .A1(n14363), .A2(n6815), .ZN(n14366) );
  NOR2_X1 U8496 ( .A1(n14477), .A2(n14468), .ZN(n7518) );
  NOR2_X1 U8497 ( .A1(n14506), .A2(n14499), .ZN(n7520) );
  AND2_X1 U8498 ( .A1(n7490), .A2(n7489), .ZN(n7488) );
  AND2_X1 U8499 ( .A1(n7489), .A2(n7491), .ZN(n7486) );
  NAND2_X1 U8500 ( .A1(n14525), .A2(n14523), .ZN(n7685) );
  NOR2_X1 U8501 ( .A1(n14555), .A2(n14730), .ZN(n7512) );
  NOR2_X1 U8502 ( .A1(n14769), .A2(n14773), .ZN(n7517) );
  INV_X1 U8503 ( .A(n11956), .ZN(n10185) );
  NAND2_X1 U8504 ( .A1(n7492), .A2(n7495), .ZN(n7491) );
  INV_X1 U8505 ( .A(n14525), .ZN(n7492) );
  NAND2_X1 U8506 ( .A1(n7493), .A2(n7495), .ZN(n7490) );
  NAND2_X1 U8507 ( .A1(n14405), .A2(n7494), .ZN(n7493) );
  INV_X1 U8508 ( .A(n7496), .ZN(n7494) );
  INV_X1 U8509 ( .A(n14503), .ZN(n14405) );
  NOR2_X1 U8510 ( .A1(n14762), .A2(n7516), .ZN(n7515) );
  INV_X1 U8511 ( .A(n7517), .ZN(n7516) );
  AND2_X1 U8512 ( .A1(n9461), .A2(n7682), .ZN(n7681) );
  AND2_X1 U8513 ( .A1(n7730), .A2(n7728), .ZN(n7727) );
  NAND2_X1 U8514 ( .A1(n7735), .A2(n7731), .ZN(n7730) );
  NAND2_X1 U8515 ( .A1(n7709), .A2(SI_24_), .ZN(n7708) );
  INV_X1 U8516 ( .A(n9063), .ZN(n7709) );
  NAND2_X1 U8517 ( .A1(n7717), .A2(SI_22_), .ZN(n7716) );
  INV_X1 U8518 ( .A(n9018), .ZN(n7717) );
  OR2_X1 U8519 ( .A1(n8996), .A2(n10463), .ZN(n8997) );
  AND2_X1 U8520 ( .A1(n9305), .A2(n7781), .ZN(n7780) );
  OR2_X1 U8521 ( .A1(n9689), .A2(P1_IR_REG_11__SCAN_IN), .ZN(n10051) );
  NOR2_X1 U8522 ( .A1(n9392), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n9550) );
  OAI21_X1 U8523 ( .B1(n9616), .B2(P2_DATAO_REG_3__SCAN_IN), .A(n7417), .ZN(
        n8598) );
  INV_X1 U8524 ( .A(P1_RD_REG_SCAN_IN), .ZN(n7444) );
  NAND2_X1 U8525 ( .A1(n7803), .A2(n7272), .ZN(n7271) );
  OAI21_X1 U8526 ( .B1(n7803), .B2(n7272), .A(P3_ADDR_REG_2__SCAN_IN), .ZN(
        n7270) );
  INV_X1 U8527 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n7272) );
  OAI21_X1 U8528 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(n15614), .A(n14837), .ZN(
        n14864) );
  AOI21_X1 U8529 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(n14842), .A(n14841), .ZN(
        n14860) );
  NOR2_X1 U8530 ( .A1(n14908), .A2(n14909), .ZN(n14841) );
  NAND2_X1 U8531 ( .A1(n15014), .A2(n12199), .ZN(n7564) );
  XNOR2_X1 U8532 ( .A(n6833), .B(n6832), .ZN(n12254) );
  INV_X1 U8533 ( .A(n6785), .ZN(n6832) );
  AND2_X1 U8534 ( .A1(n8128), .A2(n8010), .ZN(n8145) );
  XNOR2_X1 U8535 ( .A(n10660), .B(n12234), .ZN(n10771) );
  NAND2_X1 U8536 ( .A1(n12214), .A2(n7287), .ZN(n7286) );
  OR2_X1 U8537 ( .A1(n8229), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n8243) );
  INV_X1 U8538 ( .A(n12204), .ZN(n7575) );
  NAND2_X1 U8539 ( .A1(n12254), .A2(n12562), .ZN(n12320) );
  NAND2_X1 U8540 ( .A1(n10773), .A2(n7556), .ZN(n10972) );
  NOR2_X1 U8541 ( .A1(n10777), .A2(n7557), .ZN(n7556) );
  INV_X1 U8542 ( .A(n10772), .ZN(n7557) );
  XNOR2_X1 U8543 ( .A(n12477), .B(n12234), .ZN(n11248) );
  NAND2_X1 U8544 ( .A1(n7577), .A2(n7579), .ZN(n7578) );
  INV_X1 U8545 ( .A(n12223), .ZN(n7579) );
  NAND2_X1 U8546 ( .A1(n12222), .A2(n12223), .ZN(n7580) );
  INV_X1 U8547 ( .A(n6828), .ZN(n6827) );
  OAI21_X1 U8548 ( .B1(n11377), .B2(n6829), .A(n11380), .ZN(n6828) );
  INV_X1 U8549 ( .A(n11382), .ZN(n6829) );
  OR2_X1 U8550 ( .A1(n8159), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n8173) );
  MUX2_X1 U8551 ( .A(n10315), .B(n10314), .S(n12270), .Z(n10465) );
  OR2_X1 U8552 ( .A1(n8350), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n8361) );
  AND4_X1 U8553 ( .A1(n8300), .A2(n8299), .A3(n8298), .A4(n8297), .ZN(n12216)
         );
  NOR2_X1 U8554 ( .A1(n10099), .A2(n10098), .ZN(n10261) );
  OR2_X1 U8555 ( .A1(n10332), .A2(n10333), .ZN(n7694) );
  NAND2_X1 U8556 ( .A1(n10397), .A2(n10396), .ZN(n10612) );
  OR2_X1 U8557 ( .A1(n10600), .A2(n10601), .ZN(n6938) );
  NAND2_X1 U8558 ( .A1(n11026), .A2(n11027), .ZN(n15598) );
  NAND2_X1 U8559 ( .A1(n7698), .A2(n7697), .ZN(n7696) );
  NAND2_X1 U8560 ( .A1(n11024), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n7697) );
  OR2_X1 U8561 ( .A1(n11016), .A2(n15600), .ZN(n6931) );
  NOR2_X1 U8562 ( .A1(n12677), .A2(n7251), .ZN(n15627) );
  AND2_X1 U8563 ( .A1(n12678), .A2(n12679), .ZN(n7251) );
  NAND2_X1 U8564 ( .A1(n6927), .A2(n6740), .ZN(n7324) );
  XOR2_X1 U8565 ( .A(n12649), .B(n15032), .Z(n15029) );
  INV_X1 U8566 ( .A(n7253), .ZN(n12695) );
  OAI21_X1 U8567 ( .B1(n15047), .B2(n15043), .A(n15045), .ZN(n15063) );
  NAND2_X1 U8568 ( .A1(n15059), .A2(n12653), .ZN(n15075) );
  XNOR2_X1 U8569 ( .A(n7249), .B(n15073), .ZN(n15079) );
  INV_X1 U8570 ( .A(n7249), .ZN(n12702) );
  NOR2_X1 U8571 ( .A1(n12717), .A2(n12728), .ZN(n12719) );
  NAND2_X1 U8572 ( .A1(n7845), .A2(n8421), .ZN(n11850) );
  NOR2_X1 U8573 ( .A1(P3_REG3_REG_26__SCAN_IN), .A2(n8361), .ZN(n8372) );
  NAND2_X1 U8574 ( .A1(n12764), .A2(n8418), .ZN(n12752) );
  NOR2_X1 U8575 ( .A1(n8309), .A2(P3_REG3_REG_21__SCAN_IN), .ZN(n8308) );
  NAND2_X1 U8576 ( .A1(n8295), .A2(n12328), .ZN(n8309) );
  INV_X1 U8577 ( .A(n7070), .ZN(n7069) );
  AOI21_X1 U8578 ( .B1(n7068), .B2(n7070), .A(n6720), .ZN(n7067) );
  INV_X1 U8579 ( .A(n7073), .ZN(n7068) );
  AOI21_X1 U8580 ( .B1(n7410), .B2(n7408), .A(n7407), .ZN(n7406) );
  INV_X1 U8581 ( .A(n7410), .ZN(n7409) );
  INV_X1 U8582 ( .A(n12529), .ZN(n7407) );
  OR2_X1 U8583 ( .A1(n8173), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n8188) );
  INV_X1 U8584 ( .A(n8403), .ZN(n12908) );
  NAND2_X1 U8585 ( .A1(n11416), .A2(n8172), .ZN(n11415) );
  OAI21_X1 U8586 ( .B1(n11151), .B2(n7856), .A(n7047), .ZN(n11337) );
  AND2_X1 U8587 ( .A1(n7854), .A2(n7048), .ZN(n7047) );
  NAND2_X1 U8588 ( .A1(n7855), .A2(n7049), .ZN(n7048) );
  AOI21_X1 U8589 ( .B1(n12483), .B2(n7855), .A(n6683), .ZN(n7854) );
  AND2_X1 U8590 ( .A1(n8156), .A2(n11410), .ZN(n11341) );
  NOR2_X1 U8591 ( .A1(n8102), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n8128) );
  OR2_X1 U8592 ( .A1(n8088), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n8102) );
  AND3_X1 U8593 ( .A1(n8101), .A2(n8100), .A3(n8099), .ZN(n11041) );
  INV_X1 U8594 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n8076) );
  NAND2_X1 U8595 ( .A1(n10645), .A2(n8395), .ZN(n10852) );
  AND4_X1 U8596 ( .A1(n8050), .A2(n8051), .A3(n8049), .A4(n8048), .ZN(n10851)
         );
  OR2_X1 U8597 ( .A1(n8375), .A2(P3_REG3_REG_3__SCAN_IN), .ZN(n8050) );
  NAND2_X1 U8598 ( .A1(n12444), .A2(n8045), .ZN(n10644) );
  INV_X1 U8599 ( .A(n12417), .ZN(n10643) );
  AOI21_X1 U8600 ( .B1(n15693), .B2(n15692), .A(n8393), .ZN(n10646) );
  NAND2_X1 U8601 ( .A1(n10646), .A2(n12417), .ZN(n10645) );
  INV_X1 U8602 ( .A(n15017), .ZN(n12869) );
  NAND2_X1 U8603 ( .A1(n12442), .A2(n12438), .ZN(n15705) );
  INV_X1 U8604 ( .A(n12719), .ZN(n7046) );
  NAND2_X1 U8605 ( .A1(n8348), .A2(n8347), .ZN(n12296) );
  NAND2_X1 U8606 ( .A1(n8317), .A2(n8316), .ZN(n12338) );
  OR2_X1 U8607 ( .A1(n8066), .A2(n7719), .ZN(n8316) );
  XNOR2_X1 U8608 ( .A(n11150), .B(n6821), .ZN(n15758) );
  NAND2_X1 U8609 ( .A1(n7572), .A2(n8453), .ZN(n10313) );
  AND2_X1 U8610 ( .A1(n6704), .A2(n8005), .ZN(n7077) );
  AOI21_X1 U8611 ( .B1(n7152), .B2(n6692), .A(n6820), .ZN(n7990) );
  OAI21_X1 U8612 ( .B1(n8358), .B2(n7987), .A(n7988), .ZN(n8369) );
  OAI21_X1 U8613 ( .B1(n8333), .B2(P2_DATAO_REG_24__SCAN_IN), .A(n7983), .ZN(
        n8346) );
  NAND2_X1 U8614 ( .A1(n6981), .A2(n7983), .ZN(n8333) );
  NAND2_X1 U8615 ( .A1(n6983), .A2(n6982), .ZN(n6981) );
  INV_X1 U8616 ( .A(n7982), .ZN(n6983) );
  XNOR2_X1 U8617 ( .A(n8467), .B(n8466), .ZN(n10019) );
  OR2_X1 U8618 ( .A1(n7926), .A2(P3_IR_REG_20__SCAN_IN), .ZN(n7928) );
  NOR2_X1 U8619 ( .A1(n9707), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n6980) );
  INV_X1 U8620 ( .A(n6976), .ZN(n6975) );
  OAI21_X1 U8621 ( .B1(n6782), .B2(n6979), .A(n6977), .ZN(n6976) );
  INV_X1 U8622 ( .A(P3_IR_REG_11__SCAN_IN), .ZN(n8166) );
  INV_X1 U8623 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n7916) );
  NAND2_X1 U8624 ( .A1(n7037), .A2(n7248), .ZN(n7392) );
  INV_X1 U8625 ( .A(n7038), .ZN(n7037) );
  XNOR2_X1 U8626 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .ZN(n8124) );
  NOR2_X1 U8627 ( .A1(n7944), .A2(n7534), .ZN(n7533) );
  XNOR2_X1 U8628 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .ZN(n8094) );
  XNOR2_X1 U8629 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .ZN(n8052) );
  NAND2_X1 U8630 ( .A1(n13434), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n8029) );
  OR2_X1 U8631 ( .A1(n8667), .A2(n8666), .ZN(n8709) );
  INV_X1 U8632 ( .A(n13074), .ZN(n7838) );
  NAND2_X1 U8633 ( .A1(n6990), .A2(n11898), .ZN(n11902) );
  OR2_X1 U8634 ( .A1(n8937), .A2(n8936), .ZN(n8963) );
  INV_X1 U8635 ( .A(n13107), .ZN(n10624) );
  NOR2_X1 U8636 ( .A1(n7358), .A2(n6996), .ZN(n6994) );
  OAI21_X1 U8637 ( .B1(n7356), .B2(n6996), .A(n6752), .ZN(n6993) );
  INV_X1 U8638 ( .A(n11178), .ZN(n6996) );
  NOR2_X1 U8639 ( .A1(n7346), .A2(n13084), .ZN(n7344) );
  NAND2_X1 U8640 ( .A1(n6997), .A2(n13070), .ZN(n7345) );
  NAND2_X1 U8641 ( .A1(n7348), .A2(n7000), .ZN(n6997) );
  AOI21_X1 U8642 ( .B1(n13503), .B2(n7812), .A(n7811), .ZN(n7810) );
  INV_X1 U8643 ( .A(n11882), .ZN(n7812) );
  OR2_X1 U8644 ( .A1(n9066), .A2(n13527), .ZN(n9094) );
  OR2_X1 U8645 ( .A1(n10817), .A2(n10818), .ZN(n10905) );
  OAI21_X1 U8646 ( .B1(n8535), .B2(P2_IR_REG_0__SCAN_IN), .A(n7127), .ZN(n9795) );
  NAND2_X1 U8647 ( .A1(n8535), .A2(n14039), .ZN(n7127) );
  NAND2_X1 U8648 ( .A1(n8961), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8982) );
  INV_X1 U8649 ( .A(n8963), .ZN(n8961) );
  AOI22_X1 U8650 ( .A1(n7345), .A2(n13494), .B1(n7351), .B2(n7343), .ZN(n7839)
         );
  AND2_X1 U8651 ( .A1(n7344), .A2(n13494), .ZN(n7343) );
  AOI21_X1 U8652 ( .B1(n15409), .B2(n9427), .A(n9428), .ZN(n9443) );
  AOI21_X1 U8653 ( .B1(n15422), .B2(n9404), .A(n9403), .ZN(n9477) );
  NOR2_X1 U8654 ( .A1(n9477), .A2(n6845), .ZN(n15444) );
  NOR2_X1 U8655 ( .A1(n6847), .A2(n6846), .ZN(n6845) );
  NAND2_X1 U8656 ( .A1(n13602), .A2(n9530), .ZN(n13600) );
  NOR2_X1 U8657 ( .A1(n9562), .A2(n6856), .ZN(n9576) );
  AND2_X1 U8658 ( .A1(n9567), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n6856) );
  NAND2_X1 U8659 ( .A1(n6857), .A2(n10867), .ZN(n10868) );
  OR2_X1 U8660 ( .A1(n10866), .A2(n6858), .ZN(n6857) );
  INV_X1 U8661 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n6858) );
  NAND2_X1 U8662 ( .A1(n11109), .A2(n11110), .ZN(n11115) );
  NAND2_X1 U8663 ( .A1(n11115), .A2(n11114), .ZN(n11195) );
  NAND2_X1 U8664 ( .A1(n11195), .A2(n11196), .ZN(n13613) );
  NAND2_X1 U8665 ( .A1(n9172), .A2(n9171), .ZN(n13635) );
  OR2_X1 U8666 ( .A1(n14802), .A2(n9170), .ZN(n9172) );
  NAND2_X1 U8667 ( .A1(n7446), .A2(n7445), .ZN(n13705) );
  INV_X1 U8668 ( .A(n13901), .ZN(n7445) );
  NAND2_X1 U8669 ( .A1(n7450), .A2(n7449), .ZN(n13760) );
  NAND2_X1 U8670 ( .A1(n13755), .A2(n6718), .ZN(n13741) );
  NAND2_X1 U8671 ( .A1(n7224), .A2(n6738), .ZN(n13773) );
  INV_X1 U8672 ( .A(n7450), .ZN(n13774) );
  AOI21_X1 U8673 ( .B1(n7643), .B2(n7641), .A(n6748), .ZN(n7640) );
  INV_X1 U8674 ( .A(n7643), .ZN(n7642) );
  INV_X1 U8675 ( .A(n13655), .ZN(n7641) );
  OR2_X1 U8676 ( .A1(n9001), .A2(n13119), .ZN(n9024) );
  OR2_X1 U8677 ( .A1(n8982), .A2(n13537), .ZN(n9001) );
  INV_X1 U8678 ( .A(n7151), .ZN(n13822) );
  AOI21_X1 U8679 ( .B1(n7208), .B2(n7210), .A(n7206), .ZN(n7205) );
  NAND2_X1 U8680 ( .A1(n7448), .A2(n13979), .ZN(n13863) );
  NAND2_X1 U8681 ( .A1(n11529), .A2(n11528), .ZN(n11530) );
  NAND2_X1 U8682 ( .A1(n11530), .A2(n7216), .ZN(n13669) );
  NAND2_X1 U8683 ( .A1(n11231), .A2(n6710), .ZN(n11326) );
  AOI21_X1 U8684 ( .B1(n7187), .B2(n7189), .A(n6714), .ZN(n7186) );
  INV_X1 U8685 ( .A(n11229), .ZN(n15549) );
  NOR2_X1 U8686 ( .A1(n15530), .A2(n10794), .ZN(n6920) );
  NAND2_X1 U8687 ( .A1(n10574), .A2(n15521), .ZN(n10893) );
  NAND2_X1 U8688 ( .A1(n9963), .A2(n9962), .ZN(n9964) );
  NAND2_X1 U8689 ( .A1(n9904), .A2(n9903), .ZN(n9958) );
  INV_X1 U8690 ( .A(n7194), .ZN(n7193) );
  INV_X1 U8691 ( .A(n13902), .ZN(n7198) );
  INV_X1 U8692 ( .A(n13496), .ZN(n13701) );
  NAND2_X1 U8693 ( .A1(n8898), .A2(n8897), .ZN(n13985) );
  NAND2_X1 U8694 ( .A1(n8753), .A2(n8752), .ZN(n11323) );
  AND2_X1 U8695 ( .A1(n9794), .A2(n15554), .ZN(n13998) );
  NAND2_X1 U8696 ( .A1(n7648), .A2(n10787), .ZN(n10889) );
  OR2_X1 U8697 ( .A1(n10786), .A2(n10785), .ZN(n7648) );
  NAND2_X1 U8698 ( .A1(n7234), .A2(n10243), .ZN(n10533) );
  OR2_X1 U8699 ( .A1(n10130), .A2(n9170), .ZN(n7243) );
  NAND2_X1 U8700 ( .A1(n6660), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n7244) );
  OR2_X1 U8701 ( .A1(n9673), .A2(n9247), .ZN(n15554) );
  AND2_X1 U8702 ( .A1(n13365), .A2(n13366), .ZN(n7909) );
  NOR2_X1 U8703 ( .A1(P2_IR_REG_26__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), .ZN(
        n7841) );
  AND2_X1 U8704 ( .A1(n8491), .A2(n8683), .ZN(n6915) );
  INV_X1 U8705 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n9268) );
  INV_X1 U8706 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n9269) );
  NAND2_X1 U8707 ( .A1(n9271), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8527) );
  OR2_X1 U8708 ( .A1(n8853), .A2(P2_IR_REG_15__SCAN_IN), .ZN(n8895) );
  OR2_X1 U8709 ( .A1(n8825), .A2(P2_IR_REG_14__SCAN_IN), .ZN(n8853) );
  OR2_X1 U8710 ( .A1(n8685), .A2(n8684), .ZN(n8701) );
  OR2_X1 U8711 ( .A1(n6772), .A2(P2_IR_REG_3__SCAN_IN), .ZN(n8620) );
  AND3_X1 U8712 ( .A1(n6772), .A2(n6851), .A3(n6849), .ZN(n9432) );
  NAND2_X1 U8713 ( .A1(n14018), .A2(n6850), .ZN(n6849) );
  NAND2_X1 U8714 ( .A1(n8561), .A2(P2_IR_REG_2__SCAN_IN), .ZN(n6851) );
  INV_X1 U8715 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n13434) );
  OR2_X1 U8716 ( .A1(n11455), .A2(n11454), .ZN(n11464) );
  INV_X1 U8717 ( .A(n11088), .ZN(n11680) );
  INV_X1 U8718 ( .A(n9986), .ZN(n10116) );
  NAND2_X1 U8719 ( .A1(n10921), .A2(n10920), .ZN(n10926) );
  AOI21_X1 U8720 ( .B1(n7593), .B2(n6873), .A(n6872), .ZN(n6871) );
  INV_X1 U8721 ( .A(n7134), .ZN(n6873) );
  NOR2_X1 U8722 ( .A1(n11678), .A2(n11677), .ZN(n11699) );
  INV_X1 U8723 ( .A(n11807), .ZN(n11824) );
  NOR2_X1 U8724 ( .A1(n14106), .A2(n11771), .ZN(n11789) );
  INV_X1 U8725 ( .A(n11680), .ZN(n12113) );
  INV_X2 U8726 ( .A(n10116), .ZN(n11837) );
  AND2_X1 U8727 ( .A1(n14801), .A2(n9620), .ZN(n9986) );
  CLKBUF_X1 U8728 ( .A(n9339), .Z(n9343) );
  INV_X1 U8729 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n9374) );
  OAI21_X1 U8730 ( .B1(n14329), .B2(n14327), .A(n14328), .ZN(n14326) );
  NAND2_X1 U8731 ( .A1(n14326), .A2(n6955), .ZN(n9922) );
  OR2_X1 U8732 ( .A1(n14339), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6955) );
  OR2_X1 U8733 ( .A1(n6964), .A2(n6963), .ZN(n6962) );
  INV_X1 U8734 ( .A(n9859), .ZN(n6963) );
  INV_X1 U8735 ( .A(n6964), .ZN(n9860) );
  AND2_X1 U8736 ( .A1(n6962), .A2(n6961), .ZN(n10063) );
  NAND2_X1 U8737 ( .A1(n10061), .A2(n15227), .ZN(n6961) );
  NOR2_X1 U8738 ( .A1(n10063), .A2(n10062), .ZN(n10495) );
  NAND2_X1 U8739 ( .A1(n14352), .A2(n6816), .ZN(n14355) );
  NAND2_X1 U8740 ( .A1(n14355), .A2(n14356), .ZN(n14363) );
  XNOR2_X1 U8741 ( .A(n14366), .B(n7164), .ZN(n15262) );
  NAND2_X1 U8742 ( .A1(n15262), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n15261) );
  NAND2_X1 U8743 ( .A1(n7518), .A2(n14690), .ZN(n14415) );
  INV_X1 U8744 ( .A(n7518), .ZN(n14461) );
  NAND2_X1 U8745 ( .A1(n7520), .A2(n7519), .ZN(n14477) );
  NAND2_X1 U8746 ( .A1(n7512), .A2(n14532), .ZN(n14527) );
  NOR2_X1 U8747 ( .A1(n12143), .A2(n14724), .ZN(n7496) );
  AND2_X1 U8748 ( .A1(n11734), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n11753) );
  XNOR2_X1 U8749 ( .A(n14724), .B(n12143), .ZN(n14525) );
  NOR2_X1 U8750 ( .A1(n14519), .A2(n14525), .ZN(n14518) );
  INV_X1 U8751 ( .A(n7512), .ZN(n14537) );
  OAI21_X1 U8752 ( .B1(n14568), .B2(n7480), .A(n7477), .ZN(n7483) );
  INV_X1 U8753 ( .A(n7481), .ZN(n7480) );
  AOI21_X1 U8754 ( .B1(n7481), .B2(n7479), .A(n7478), .ZN(n7477) );
  NAND2_X1 U8755 ( .A1(n7668), .A2(n7479), .ZN(n14576) );
  INV_X1 U8756 ( .A(n14578), .ZN(n7668) );
  NAND2_X1 U8757 ( .A1(n14568), .A2(n14579), .ZN(n14567) );
  INV_X1 U8758 ( .A(n7677), .ZN(n7676) );
  AOI21_X1 U8759 ( .B1(n7465), .B2(n7468), .A(n7464), .ZN(n14584) );
  INV_X1 U8760 ( .A(n7466), .ZN(n7464) );
  AOI21_X1 U8761 ( .B1(n7468), .B2(n7467), .A(n14399), .ZN(n7466) );
  NAND2_X1 U8762 ( .A1(n14670), .A2(n7517), .ZN(n14636) );
  NAND2_X1 U8763 ( .A1(n11640), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n11663) );
  NAND2_X1 U8764 ( .A1(n6763), .A2(n6680), .ZN(n7471) );
  INV_X1 U8765 ( .A(n7662), .ZN(n7661) );
  NAND2_X1 U8766 ( .A1(n14670), .A2(n14651), .ZN(n14647) );
  NAND2_X1 U8767 ( .A1(n11461), .A2(n12147), .ZN(n14661) );
  NOR2_X1 U8768 ( .A1(n11292), .A2(n11291), .ZN(n11299) );
  NAND2_X1 U8769 ( .A1(n11290), .A2(n11289), .ZN(n14955) );
  OR2_X1 U8770 ( .A1(n11076), .A2(n11075), .ZN(n11086) );
  OR2_X1 U8771 ( .A1(n11086), .A2(n11085), .ZN(n11292) );
  AND2_X1 U8772 ( .A1(n15360), .A2(n11097), .ZN(n15274) );
  INV_X1 U8773 ( .A(n7511), .ZN(n15287) );
  OAI21_X1 U8774 ( .B1(n10845), .B2(n10844), .A(n10843), .ZN(n10846) );
  NAND2_X1 U8775 ( .A1(n10458), .A2(n10457), .ZN(n10740) );
  NOR2_X1 U8776 ( .A1(n10422), .A2(n7655), .ZN(n7654) );
  INV_X1 U8777 ( .A(n10131), .ZN(n7655) );
  INV_X1 U8778 ( .A(n15319), .ZN(n11960) );
  NAND2_X1 U8779 ( .A1(n15288), .A2(n14612), .ZN(n9974) );
  NOR2_X1 U8780 ( .A1(n14450), .A2(n6677), .ZN(n7454) );
  NOR2_X1 U8781 ( .A1(n7463), .A2(n6700), .ZN(n7459) );
  NAND2_X1 U8782 ( .A1(n7459), .A2(n6677), .ZN(n7456) );
  NAND2_X1 U8783 ( .A1(n7463), .A2(n6700), .ZN(n7460) );
  INV_X1 U8784 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n9308) );
  OAI21_X1 U8785 ( .B1(n9465), .B2(P1_IR_REG_22__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n9309) );
  XNOR2_X1 U8786 ( .A(n9188), .B(n9187), .ZN(n14021) );
  INV_X1 U8787 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n7682) );
  INV_X1 U8788 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n9461) );
  XNOR2_X1 U8789 ( .A(n9321), .B(P1_IR_REG_26__SCAN_IN), .ZN(n9383) );
  XNOR2_X1 U8790 ( .A(n9106), .B(n9105), .ZN(n14035) );
  XNOR2_X1 U8791 ( .A(n9320), .B(P1_IR_REG_24__SCAN_IN), .ZN(n9380) );
  XNOR2_X1 U8792 ( .A(n9061), .B(n9041), .ZN(n11731) );
  NAND3_X1 U8793 ( .A1(n7718), .A2(n7716), .A3(n7715), .ZN(n11714) );
  XNOR2_X1 U8794 ( .A(n8957), .B(n8956), .ZN(n11656) );
  NAND2_X1 U8795 ( .A1(n8875), .A2(n8874), .ZN(n8930) );
  NAND2_X1 U8796 ( .A1(n7750), .A2(n8820), .ZN(n8846) );
  NAND2_X1 U8797 ( .A1(n7011), .A2(n8816), .ZN(n7750) );
  AND2_X1 U8798 ( .A1(n9811), .A2(n9705), .ZN(n11446) );
  NAND2_X1 U8799 ( .A1(n7180), .A2(n8633), .ZN(n8656) );
  NAND2_X1 U8800 ( .A1(n14877), .A2(P3_ADDR_REG_0__SCAN_IN), .ZN(n14876) );
  XNOR2_X1 U8801 ( .A(n14874), .B(n6837), .ZN(n14878) );
  INV_X1 U8802 ( .A(n14876), .ZN(n6837) );
  XNOR2_X1 U8803 ( .A(n14869), .B(n7805), .ZN(n14870) );
  INV_X1 U8804 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n7805) );
  INV_X1 U8805 ( .A(n7267), .ZN(n14827) );
  OAI21_X1 U8806 ( .B1(n15237), .B2(n15238), .A(n7264), .ZN(n7263) );
  INV_X1 U8807 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n7264) );
  OAI21_X1 U8808 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(n14846), .A(n14845), .ZN(
        n14859) );
  INV_X1 U8809 ( .A(n7792), .ZN(n7791) );
  INV_X1 U8810 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n7798) );
  INV_X1 U8811 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n7787) );
  NAND2_X1 U8812 ( .A1(n7563), .A2(n7564), .ZN(n12249) );
  NAND2_X1 U8813 ( .A1(n15016), .A2(n7565), .ZN(n7563) );
  NAND2_X1 U8814 ( .A1(n10470), .A2(n10479), .ZN(n10773) );
  AND2_X1 U8815 ( .A1(n7550), .A2(n10471), .ZN(n10470) );
  XNOR2_X1 U8816 ( .A(n10771), .B(n10851), .ZN(n7550) );
  NAND2_X1 U8817 ( .A1(n12344), .A2(n12211), .ZN(n12263) );
  INV_X1 U8818 ( .A(n7281), .ZN(n7277) );
  NAND2_X1 U8819 ( .A1(n7286), .A2(n7291), .ZN(n12278) );
  NAND2_X1 U8820 ( .A1(n10773), .A2(n10772), .ZN(n10778) );
  NAND2_X1 U8821 ( .A1(n12214), .A2(n12260), .ZN(n12327) );
  NAND2_X1 U8822 ( .A1(n7580), .A2(n7578), .ZN(n12335) );
  NAND2_X1 U8823 ( .A1(n12346), .A2(n12345), .ZN(n12344) );
  NAND2_X1 U8824 ( .A1(n12308), .A2(n12208), .ZN(n12346) );
  OAI21_X1 U8825 ( .B1(n15016), .B2(n7561), .A(n7558), .ZN(n12365) );
  AOI21_X1 U8826 ( .B1(n7560), .B2(n7559), .A(n6796), .ZN(n7558) );
  INV_X1 U8827 ( .A(n7565), .ZN(n7559) );
  AND2_X1 U8828 ( .A1(n8434), .A2(n12593), .ZN(n12867) );
  NAND2_X1 U8829 ( .A1(n12609), .A2(n12608), .ZN(n7548) );
  NOR4_X1 U8830 ( .A1(n12599), .A2(n12434), .A3(n12598), .A4(n12596), .ZN(
        n12435) );
  INV_X1 U8831 ( .A(n12615), .ZN(n7546) );
  INV_X1 U8832 ( .A(n10765), .ZN(n12613) );
  INV_X1 U8833 ( .A(n12362), .ZN(n12868) );
  INV_X1 U8834 ( .A(n12199), .ZN(n15013) );
  INV_X1 U8835 ( .A(n12498), .ZN(n12630) );
  NOR2_X1 U8836 ( .A1(n7042), .A2(n6747), .ZN(n7124) );
  NAND2_X1 U8837 ( .A1(n10361), .A2(n10521), .ZN(n10360) );
  NOR2_X1 U8838 ( .A1(n10518), .A2(n10519), .ZN(n10521) );
  INV_X1 U8839 ( .A(n6936), .ZN(n10093) );
  INV_X1 U8840 ( .A(n7695), .ZN(n10334) );
  XOR2_X1 U8841 ( .A(n10612), .B(n10613), .Z(n10398) );
  INV_X1 U8842 ( .A(n7698), .ZN(n11013) );
  INV_X1 U8843 ( .A(n6938), .ZN(n10604) );
  INV_X1 U8844 ( .A(P3_ADDR_REG_9__SCAN_IN), .ZN(n15614) );
  OAI21_X1 U8845 ( .B1(n15616), .B2(n7332), .A(n7331), .ZN(n15632) );
  NAND2_X1 U8846 ( .A1(n7333), .A2(P3_REG2_REG_11__SCAN_IN), .ZN(n7332) );
  XNOR2_X1 U8847 ( .A(n12659), .B(n12688), .ZN(n15650) );
  INV_X1 U8848 ( .A(n6927), .ZN(n15649) );
  INV_X1 U8849 ( .A(n7688), .ZN(n15666) );
  INV_X1 U8850 ( .A(n7324), .ZN(n15668) );
  NOR2_X1 U8851 ( .A1(n15026), .A2(n15027), .ZN(n15025) );
  OAI22_X1 U8852 ( .A1(n6935), .A2(n15053), .B1(n15026), .B2(n6934), .ZN(
        n15054) );
  NAND2_X1 U8853 ( .A1(n7691), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n6934) );
  INV_X1 U8854 ( .A(n12662), .ZN(n6935) );
  XNOR2_X1 U8855 ( .A(n12663), .B(n7689), .ZN(n15066) );
  NOR2_X1 U8856 ( .A1(n15066), .A2(n15067), .ZN(n15068) );
  OAI21_X1 U8857 ( .B1(n15066), .B2(n7329), .A(n7328), .ZN(n15084) );
  NAND2_X1 U8858 ( .A1(n7330), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n7329) );
  NAND2_X1 U8859 ( .A1(n12664), .A2(n7330), .ZN(n7328) );
  INV_X1 U8860 ( .A(n15083), .ZN(n7330) );
  INV_X1 U8861 ( .A(n12672), .ZN(n7084) );
  NAND2_X1 U8862 ( .A1(n11853), .A2(n8422), .ZN(n7142) );
  NAND2_X1 U8863 ( .A1(n8360), .A2(n8359), .ZN(n12747) );
  OR2_X1 U8864 ( .A1(n8066), .A2(n11425), .ZN(n8359) );
  NAND2_X1 U8865 ( .A1(n12772), .A2(n12566), .ZN(n12758) );
  NAND2_X1 U8866 ( .A1(n12783), .A2(n8417), .ZN(n12766) );
  NAND2_X1 U8867 ( .A1(n7050), .A2(n7053), .ZN(n12795) );
  NAND2_X1 U8868 ( .A1(n12816), .A2(n7055), .ZN(n7050) );
  NAND2_X1 U8869 ( .A1(n7388), .A2(n12555), .ZN(n12799) );
  NAND2_X1 U8870 ( .A1(n12809), .A2(n12554), .ZN(n7388) );
  NAND2_X1 U8871 ( .A1(n12818), .A2(n8414), .ZN(n12805) );
  NAND2_X1 U8872 ( .A1(n8294), .A2(n8293), .ZN(n12954) );
  OR2_X1 U8873 ( .A1(n8066), .A2(n10463), .ZN(n8293) );
  NAND2_X1 U8874 ( .A1(n12840), .A2(n8413), .ZN(n12830) );
  NAND2_X1 U8875 ( .A1(n7398), .A2(n12536), .ZN(n12834) );
  OR2_X1 U8876 ( .A1(n12847), .A2(n8278), .ZN(n7398) );
  NAND2_X1 U8877 ( .A1(n7072), .A2(n8409), .ZN(n12866) );
  NAND2_X1 U8878 ( .A1(n7079), .A2(n7073), .ZN(n7072) );
  NAND2_X1 U8879 ( .A1(n7079), .A2(n8407), .ZN(n12881) );
  NAND2_X1 U8880 ( .A1(n12904), .A2(n8405), .ZN(n15091) );
  NAND2_X1 U8881 ( .A1(n11143), .A2(n7855), .ZN(n11366) );
  NAND2_X1 U8882 ( .A1(n11143), .A2(n8401), .ZN(n11364) );
  OAI21_X1 U8883 ( .B1(n8116), .B2(n7384), .A(n7381), .ZN(n11363) );
  NAND2_X1 U8884 ( .A1(n8116), .A2(n8115), .ZN(n11142) );
  OAI211_X1 U8885 ( .C1(n11152), .C2(n6821), .A(n11151), .B(n15695), .ZN(
        n11153) );
  INV_X1 U8886 ( .A(n12827), .ZN(n15098) );
  NAND2_X1 U8887 ( .A1(n10726), .A2(n8397), .ZN(n11053) );
  AND3_X1 U8888 ( .A1(n8073), .A2(n8072), .A3(n8071), .ZN(n15736) );
  NAND2_X1 U8889 ( .A1(n12610), .A2(n9883), .ZN(n15711) );
  INV_X1 U8890 ( .A(n15711), .ZN(n12911) );
  INV_X2 U8891 ( .A(n15719), .ZN(n15703) );
  INV_X1 U8892 ( .A(n12404), .ZN(n12990) );
  INV_X1 U8893 ( .A(n12747), .ZN(n12999) );
  INV_X1 U8894 ( .A(n12296), .ZN(n13003) );
  AND2_X1 U8895 ( .A1(n12957), .A2(n12956), .ZN(n13020) );
  NAND2_X1 U8896 ( .A1(n8255), .A2(n8254), .ZN(n13032) );
  AND3_X1 U8897 ( .A1(n8187), .A2(n8186), .A3(n8185), .ZN(n13044) );
  AND2_X1 U8898 ( .A1(n8451), .A2(n8450), .ZN(n13050) );
  INV_X1 U8899 ( .A(n9323), .ZN(n13051) );
  INV_X1 U8900 ( .A(P3_IR_REG_30__SCAN_IN), .ZN(n8006) );
  NAND2_X1 U8901 ( .A1(n7078), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8007) );
  NAND2_X1 U8902 ( .A1(n8000), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n6834) );
  INV_X1 U8903 ( .A(SI_27_), .ZN(n13471) );
  INV_X1 U8904 ( .A(n10016), .ZN(n12696) );
  INV_X1 U8905 ( .A(n8465), .ZN(n11427) );
  NAND2_X1 U8906 ( .A1(n8446), .A2(n8445), .ZN(n11169) );
  MUX2_X1 U8907 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8444), .S(
        P3_IR_REG_24__SCAN_IN), .Z(n8446) );
  NAND2_X1 U8908 ( .A1(n7583), .A2(n7859), .ZN(n8443) );
  XNOR2_X1 U8909 ( .A(n8333), .B(n11510), .ZN(n11166) );
  XNOR2_X1 U8910 ( .A(n7921), .B(n7920), .ZN(n10765) );
  INV_X1 U8911 ( .A(P3_IR_REG_22__SCAN_IN), .ZN(n7920) );
  OAI21_X1 U8912 ( .B1(n7928), .B2(P3_IR_REG_21__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n7921) );
  NAND2_X1 U8913 ( .A1(n7977), .A2(n7976), .ZN(n8302) );
  INV_X1 U8914 ( .A(n8481), .ZN(n10462) );
  NAND2_X1 U8915 ( .A1(n7521), .A2(n7524), .ZN(n8280) );
  NAND2_X1 U8916 ( .A1(n8251), .A2(n7527), .ZN(n7521) );
  NAND2_X1 U8917 ( .A1(n7529), .A2(n7531), .ZN(n8262) );
  NAND2_X1 U8918 ( .A1(n7530), .A2(n8250), .ZN(n7529) );
  INV_X1 U8919 ( .A(n8251), .ZN(n7530) );
  INV_X1 U8920 ( .A(n7967), .ZN(n8236) );
  INV_X1 U8921 ( .A(SI_16_), .ZN(n13466) );
  INV_X1 U8922 ( .A(SI_15_), .ZN(n9561) );
  NAND2_X1 U8923 ( .A1(n7541), .A2(n7539), .ZN(n8223) );
  NAND2_X1 U8924 ( .A1(n7541), .A2(n7962), .ZN(n8221) );
  INV_X1 U8925 ( .A(SI_14_), .ZN(n14937) );
  NAND2_X1 U8926 ( .A1(n7549), .A2(n7960), .ZN(n8196) );
  NAND2_X1 U8927 ( .A1(n8182), .A2(n6782), .ZN(n7549) );
  NAND2_X1 U8928 ( .A1(n6974), .A2(n9707), .ZN(n7960) );
  INV_X1 U8929 ( .A(n12685), .ZN(n15640) );
  NAND2_X1 U8930 ( .A1(n6970), .A2(n6972), .ZN(n8169) );
  NAND2_X1 U8931 ( .A1(n6971), .A2(n7956), .ZN(n6970) );
  INV_X1 U8932 ( .A(n15622), .ZN(n12682) );
  NAND2_X1 U8933 ( .A1(n7955), .A2(n7954), .ZN(n8153) );
  INV_X1 U8934 ( .A(n10611), .ZN(n11024) );
  INV_X1 U8935 ( .A(n10393), .ZN(n10401) );
  NAND2_X1 U8936 ( .A1(n7535), .A2(n7943), .ZN(n8085) );
  NAND2_X1 U8937 ( .A1(n7842), .A2(n7917), .ZN(n8054) );
  AND2_X1 U8938 ( .A1(n10519), .A2(n8040), .ZN(n7842) );
  INV_X1 U8939 ( .A(n10092), .ZN(n10107) );
  NAND2_X1 U8940 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), .ZN(
        n7692) );
  NAND2_X1 U8941 ( .A1(n9274), .A2(n9281), .ZN(n9394) );
  NAND2_X1 U8942 ( .A1(n10905), .A2(n10904), .ZN(n11002) );
  NAND2_X1 U8943 ( .A1(n7816), .A2(n7814), .ZN(n13092) );
  NAND2_X1 U8944 ( .A1(n8535), .A2(n6913), .ZN(n6914) );
  OR2_X1 U8945 ( .A1(n8535), .A2(n8537), .ZN(n8538) );
  AND2_X1 U8946 ( .A1(n9816), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n6913) );
  INV_X1 U8947 ( .A(n11908), .ZN(n7337) );
  INV_X1 U8948 ( .A(n13535), .ZN(n7338) );
  NAND2_X1 U8949 ( .A1(n10160), .A2(n10159), .ZN(n10161) );
  NAND2_X1 U8950 ( .A1(n7348), .A2(n7001), .ZN(n7347) );
  NAND2_X1 U8951 ( .A1(n7351), .A2(n7350), .ZN(n7349) );
  INV_X1 U8952 ( .A(n9795), .ZN(n10295) );
  INV_X1 U8953 ( .A(n13681), .ZN(n13958) );
  AOI21_X1 U8954 ( .B1(n11905), .B2(n13533), .A(n13532), .ZN(n13535) );
  NAND2_X1 U8955 ( .A1(n11190), .A2(n11189), .ZN(n11866) );
  NAND2_X1 U8956 ( .A1(n13656), .A2(n11865), .ZN(n7809) );
  XNOR2_X1 U8957 ( .A(n13062), .B(n13064), .ZN(n11915) );
  NAND2_X1 U8958 ( .A1(n6995), .A2(n7356), .ZN(n11179) );
  NAND2_X1 U8959 ( .A1(n10817), .A2(n7357), .ZN(n6995) );
  NAND2_X1 U8960 ( .A1(n9695), .A2(n9694), .ZN(n9696) );
  NAND2_X1 U8961 ( .A1(n9696), .A2(n9697), .ZN(n9935) );
  NAND2_X1 U8962 ( .A1(n13516), .A2(n11892), .ZN(n13544) );
  NAND2_X1 U8963 ( .A1(n7839), .A2(n13074), .ZN(n13552) );
  NAND2_X1 U8964 ( .A1(n9110), .A2(n9109), .ZN(n13918) );
  NAND2_X1 U8965 ( .A1(n8856), .A2(n8855), .ZN(n13991) );
  NAND2_X1 U8966 ( .A1(n9246), .A2(n9245), .ZN(n6909) );
  NOR2_X1 U8967 ( .A1(n9275), .A2(n7087), .ZN(n9292) );
  OR2_X1 U8968 ( .A1(n9298), .A2(n7088), .ZN(n7087) );
  NAND2_X1 U8969 ( .A1(n10983), .A2(n10763), .ZN(n7088) );
  NAND2_X1 U8970 ( .A1(n9138), .A2(n9137), .ZN(n13694) );
  NAND2_X1 U8971 ( .A1(n9119), .A2(n9118), .ZN(n13663) );
  NOR2_X1 U8972 ( .A1(n6735), .A2(n7620), .ZN(n8539) );
  AOI21_X1 U8973 ( .B1(n8553), .B2(P2_REG2_REG_0__SCAN_IN), .A(n6757), .ZN(
        n8510) );
  NOR2_X1 U8974 ( .A1(n15444), .A2(n15443), .ZN(n15441) );
  NOR2_X1 U8975 ( .A1(n9533), .A2(n9532), .ZN(n9562) );
  NAND2_X1 U8976 ( .A1(n13600), .A2(n13601), .ZN(n9533) );
  XNOR2_X1 U8977 ( .A(n10868), .B(n15478), .ZN(n15475) );
  INV_X1 U8978 ( .A(n13635), .ZN(n13899) );
  NOR2_X1 U8979 ( .A1(n13697), .A2(n6702), .ZN(n7196) );
  NAND2_X1 U8980 ( .A1(n6702), .A2(n13697), .ZN(n7194) );
  INV_X1 U8981 ( .A(n13905), .ZN(n13725) );
  NAND2_X1 U8982 ( .A1(n13693), .A2(n7699), .ZN(n7236) );
  NAND2_X1 U8983 ( .A1(n13693), .A2(n7700), .ZN(n13714) );
  OAI211_X1 U8984 ( .C1(n13659), .C2(n6697), .A(n7202), .B(n7623), .ZN(n13913)
         );
  INV_X1 U8985 ( .A(n7203), .ZN(n7202) );
  OAI21_X1 U8986 ( .B1(n6697), .B2(n13658), .A(n13737), .ZN(n7203) );
  OAI21_X1 U8987 ( .B1(n7201), .B2(n7200), .A(n7199), .ZN(n13738) );
  NAND2_X1 U8988 ( .A1(n7623), .A2(n13658), .ZN(n7201) );
  NAND2_X1 U8989 ( .A1(n7623), .A2(n6697), .ZN(n7199) );
  OAI21_X1 U8990 ( .B1(n6699), .B2(n7628), .A(n7627), .ZN(n13750) );
  NAND2_X1 U8991 ( .A1(n13769), .A2(n13661), .ZN(n13754) );
  NAND2_X1 U8992 ( .A1(n7226), .A2(n7229), .ZN(n13784) );
  NAND2_X1 U8993 ( .A1(n13807), .A2(n7230), .ZN(n7226) );
  AOI21_X1 U8994 ( .B1(n13807), .B2(n13806), .A(n6696), .ZN(n13793) );
  AND2_X1 U8995 ( .A1(n7437), .A2(n7743), .ZN(n13820) );
  OAI21_X1 U8996 ( .B1(n13860), .B2(n7210), .A(n7208), .ZN(n13837) );
  NAND2_X1 U8997 ( .A1(n13678), .A2(n13677), .ZN(n13829) );
  NAND2_X1 U8998 ( .A1(n7241), .A2(n7240), .ZN(n13678) );
  OAI21_X1 U8999 ( .B1(n13860), .B2(n7213), .A(n13648), .ZN(n13856) );
  NAND2_X1 U9000 ( .A1(n7207), .A2(n7211), .ZN(n13854) );
  NAND2_X1 U9001 ( .A1(n13860), .A2(n13648), .ZN(n7207) );
  AND2_X1 U9002 ( .A1(n7241), .A2(n7242), .ZN(n13841) );
  OAI21_X1 U9003 ( .B1(n7637), .B2(n7219), .A(n7217), .ZN(n13642) );
  AND2_X1 U9004 ( .A1(n7246), .A2(n6715), .ZN(n11494) );
  NAND2_X1 U9005 ( .A1(n7221), .A2(n11488), .ZN(n11527) );
  NAND2_X1 U9006 ( .A1(n7637), .A2(n7222), .ZN(n7221) );
  NAND2_X1 U9007 ( .A1(n7703), .A2(n7702), .ZN(n11489) );
  NAND2_X1 U9008 ( .A1(n7637), .A2(n11322), .ZN(n11487) );
  NAND2_X1 U9009 ( .A1(n8781), .A2(n8780), .ZN(n15140) );
  NAND2_X1 U9010 ( .A1(n10987), .A2(n10986), .ZN(n11225) );
  INV_X1 U9011 ( .A(n13859), .ZN(n13872) );
  NAND2_X1 U9012 ( .A1(n7753), .A2(n10534), .ZN(n10568) );
  NAND2_X1 U9013 ( .A1(n10238), .A2(n10237), .ZN(n10545) );
  OR2_X1 U9014 ( .A1(n15151), .A2(n9175), .ZN(n13870) );
  OR2_X1 U9015 ( .A1(n15151), .A2(n10236), .ZN(n13874) );
  OR2_X1 U9016 ( .A1(n15151), .A2(n10250), .ZN(n13890) );
  NAND2_X1 U9017 ( .A1(n15491), .A2(n9678), .ZN(n13865) );
  INV_X1 U9018 ( .A(n13870), .ZN(n15147) );
  NAND2_X1 U9019 ( .A1(n10706), .A2(n7704), .ZN(n9967) );
  AOI21_X1 U9020 ( .B1(n10704), .B2(n15539), .A(n6813), .ZN(n7704) );
  AND2_X1 U9021 ( .A1(n9945), .A2(P2_STATE_REG_SCAN_IN), .ZN(n15491) );
  NAND2_X1 U9022 ( .A1(n7118), .A2(n7116), .ZN(n8506) );
  NAND2_X1 U9023 ( .A1(n7117), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7116) );
  XNOR2_X1 U9024 ( .A(n9286), .B(n8500), .ZN(n14033) );
  NAND2_X1 U9025 ( .A1(n9284), .A2(n9283), .ZN(n11511) );
  INV_X1 U9026 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n11860) );
  INV_X1 U9027 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n13423) );
  INV_X1 U9028 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n10735) );
  NAND2_X1 U9029 ( .A1(n8495), .A2(n8778), .ZN(n8932) );
  INV_X1 U9030 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n10153) );
  INV_X1 U9031 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n9971) );
  INV_X1 U9032 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n9594) );
  INV_X1 U9033 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n9548) );
  AND2_X1 U9034 ( .A1(n8663), .A2(n8681), .ZN(n13589) );
  INV_X1 U9035 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n13274) );
  INV_X1 U9036 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n9331) );
  NAND2_X1 U9037 ( .A1(n10921), .A2(n6866), .ZN(n6869) );
  NOR2_X1 U9038 ( .A1(n6868), .A2(n6867), .ZN(n6866) );
  OAI21_X1 U9039 ( .B1(n14193), .B2(n11802), .A(n6676), .ZN(n14041) );
  NAND2_X1 U9040 ( .A1(n7606), .A2(n7605), .ZN(n15169) );
  NAND2_X1 U9041 ( .A1(n11546), .A2(n11545), .ZN(n11572) );
  NAND2_X1 U9042 ( .A1(n10678), .A2(n7608), .ZN(n14059) );
  NOR2_X1 U9043 ( .A1(n14057), .A2(n7609), .ZN(n7608) );
  INV_X1 U9044 ( .A(n10677), .ZN(n7609) );
  NAND2_X1 U9045 ( .A1(n10129), .A2(n7777), .ZN(n14064) );
  INV_X1 U9046 ( .A(n7775), .ZN(n7777) );
  OAI21_X1 U9047 ( .B1(n10130), .B2(n12109), .A(n7778), .ZN(n7775) );
  AOI21_X1 U9048 ( .B1(n6676), .B2(n11802), .A(n11820), .ZN(n7586) );
  NAND2_X1 U9049 ( .A1(n11355), .A2(n7616), .ZN(n11519) );
  AND2_X1 U9050 ( .A1(n11355), .A2(n11354), .ZN(n11356) );
  AND2_X1 U9051 ( .A1(n7603), .A2(n6717), .ZN(n14080) );
  NAND2_X1 U9052 ( .A1(n11612), .A2(n7611), .ZN(n6862) );
  INV_X1 U9053 ( .A(n6864), .ZN(n6863) );
  NAND2_X1 U9054 ( .A1(n10926), .A2(n10925), .ZN(n10928) );
  AOI21_X1 U9055 ( .B1(n14134), .B2(n14133), .A(n14132), .ZN(n14136) );
  XNOR2_X1 U9056 ( .A(n10924), .B(n10922), .ZN(n10921) );
  NAND2_X1 U9057 ( .A1(n7594), .A2(n7597), .ZN(n14165) );
  NAND2_X1 U9058 ( .A1(n7596), .A2(n7595), .ZN(n7594) );
  INV_X1 U9059 ( .A(n11695), .ZN(n7596) );
  AND2_X1 U9060 ( .A1(n7619), .A2(n11577), .ZN(n14173) );
  NAND4_X1 U9061 ( .A1(n9972), .A2(n9975), .A3(n9772), .A4(n9628), .ZN(n15167)
         );
  XNOR2_X1 U9062 ( .A(n11618), .B(n11619), .ZN(n14206) );
  NAND2_X1 U9063 ( .A1(n15169), .A2(n11612), .ZN(n11618) );
  AND2_X1 U9064 ( .A1(n14159), .A2(n15379), .ZN(n15172) );
  AND2_X1 U9065 ( .A1(n7499), .A2(n7500), .ZN(n7498) );
  INV_X1 U9066 ( .A(n14269), .ZN(n6949) );
  INV_X1 U9067 ( .A(n14268), .ZN(n6948) );
  INV_X1 U9068 ( .A(n14253), .ZN(n14270) );
  INV_X1 U9069 ( .A(n6960), .ZN(n14296) );
  NAND2_X1 U9070 ( .A1(n14295), .A2(n6956), .ZN(n9889) );
  NAND2_X1 U9071 ( .A1(n6958), .A2(n6957), .ZN(n6956) );
  NAND2_X1 U9072 ( .A1(n14311), .A2(n6787), .ZN(n9717) );
  INV_X1 U9073 ( .A(n6962), .ZN(n10060) );
  NAND2_X1 U9074 ( .A1(n12129), .A2(n12128), .ZN(n14679) );
  OAI21_X1 U9075 ( .B1(n14460), .B2(n15351), .A(n14459), .ZN(n14695) );
  AOI21_X1 U9076 ( .B1(n14447), .B2(n15378), .A(n14458), .ZN(n14459) );
  XNOR2_X1 U9077 ( .A(n14455), .B(n14454), .ZN(n14460) );
  NAND2_X1 U9078 ( .A1(n7034), .A2(n14445), .ZN(n14483) );
  NAND2_X1 U9079 ( .A1(n14524), .A2(n7687), .ZN(n14502) );
  AND2_X1 U9080 ( .A1(n14524), .A2(n14442), .ZN(n14504) );
  AND2_X1 U9081 ( .A1(n11676), .A2(n11675), .ZN(n14749) );
  NAND2_X1 U9082 ( .A1(n14621), .A2(n14397), .ZN(n14603) );
  AND2_X1 U9083 ( .A1(n14621), .A2(n7468), .ZN(n14602) );
  NAND2_X1 U9084 ( .A1(n7675), .A2(n14432), .ZN(n14601) );
  NAND2_X1 U9085 ( .A1(n7126), .A2(n6701), .ZN(n7675) );
  AND2_X1 U9086 ( .A1(n14625), .A2(n14624), .ZN(n14765) );
  NAND2_X1 U9087 ( .A1(n7126), .A2(n14428), .ZN(n14617) );
  AND2_X1 U9088 ( .A1(n7473), .A2(n6684), .ZN(n14646) );
  NAND2_X1 U9089 ( .A1(n14658), .A2(n14422), .ZN(n14644) );
  NAND2_X1 U9090 ( .A1(n7473), .A2(n7474), .ZN(n14664) );
  NOR2_X1 U9091 ( .A1(n12147), .A2(n7658), .ZN(n7657) );
  INV_X1 U9092 ( .A(n11479), .ZN(n7658) );
  NAND2_X1 U9093 ( .A1(n7659), .A2(n11479), .ZN(n11481) );
  NAND2_X1 U9094 ( .A1(n11284), .A2(n11283), .ZN(n15183) );
  NAND2_X1 U9095 ( .A1(n11074), .A2(n11073), .ZN(n15380) );
  NAND2_X1 U9096 ( .A1(n15273), .A2(n7506), .ZN(n15374) );
  AND2_X1 U9097 ( .A1(n11099), .A2(n11098), .ZN(n7506) );
  AND2_X1 U9098 ( .A1(n15273), .A2(n11098), .ZN(n11100) );
  NAND2_X1 U9099 ( .A1(n11067), .A2(n11066), .ZN(n15286) );
  NAND2_X1 U9100 ( .A1(n10831), .A2(n10830), .ZN(n11998) );
  OAI21_X1 U9101 ( .B1(n7139), .B2(n7674), .A(n7672), .ZN(n10825) );
  NAND2_X1 U9102 ( .A1(n7139), .A2(n10428), .ZN(n10760) );
  NAND2_X1 U9103 ( .A1(n7656), .A2(n10131), .ZN(n10423) );
  OR2_X1 U9104 ( .A1(n6665), .A2(n9997), .ZN(n15297) );
  OR2_X1 U9105 ( .A1(n14409), .A2(n14612), .ZN(n14550) );
  INV_X1 U9106 ( .A(n14982), .ZN(n15191) );
  NAND2_X1 U9107 ( .A1(n15389), .A2(n15375), .ZN(n7458) );
  INV_X1 U9108 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n7462) );
  AND4_X1 U9109 ( .A1(n14712), .A2(n14711), .A3(n14710), .A4(n14709), .ZN(
        n14713) );
  AND4_X1 U9110 ( .A1(n14740), .A2(n14739), .A3(n14738), .A4(n14737), .ZN(
        n14741) );
  NAND2_X1 U9111 ( .A1(n7159), .A2(n7157), .ZN(n9557) );
  NAND2_X1 U9112 ( .A1(n7158), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7157) );
  INV_X1 U9113 ( .A(n9317), .ZN(n9314) );
  XNOR2_X1 U9114 ( .A(n11715), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n14818) );
  OR2_X1 U9115 ( .A1(n11714), .A2(n9616), .ZN(n11715) );
  NAND2_X1 U9116 ( .A1(n9610), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9463) );
  INV_X1 U9117 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n10721) );
  INV_X1 U9118 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n10234) );
  INV_X1 U9119 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n10054) );
  INV_X1 U9120 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n9691) );
  INV_X1 U9121 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n9553) );
  INV_X1 U9122 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n9391) );
  INV_X1 U9123 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n9376) );
  INV_X1 U9124 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n9373) );
  INV_X1 U9125 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n10427) );
  XNOR2_X1 U9126 ( .A(n8596), .B(n8597), .ZN(n10130) );
  NAND2_X1 U9127 ( .A1(n7412), .A2(n8579), .ZN(n8597) );
  NAND2_X1 U9128 ( .A1(n7413), .A2(n7414), .ZN(n7412) );
  INV_X1 U9129 ( .A(n8577), .ZN(n7414) );
  XNOR2_X1 U9130 ( .A(n8576), .B(n8577), .ZN(n9982) );
  NAND2_X1 U9131 ( .A1(n6954), .A2(n6952), .ZN(n9333) );
  NAND2_X1 U9132 ( .A1(n9336), .A2(n6953), .ZN(n6952) );
  OAI211_X1 U9133 ( .C1(P1_IR_REG_0__SCAN_IN), .C2(P1_IR_REG_1__SCAN_IN), .A(
        P1_IR_REG_2__SCAN_IN), .B(P1_IR_REG_31__SCAN_IN), .ZN(n6954) );
  XNOR2_X1 U9134 ( .A(n9360), .B(P1_IR_REG_1__SCAN_IN), .ZN(n14234) );
  INV_X1 U9135 ( .A(n6836), .ZN(n14880) );
  XNOR2_X1 U9136 ( .A(n14870), .B(P2_ADDR_REG_4__SCAN_IN), .ZN(n15791) );
  OAI211_X1 U9137 ( .C1(n14942), .C2(n7262), .A(n7260), .B(n7259), .ZN(n14950)
         );
  NAND2_X1 U9138 ( .A1(n7261), .A2(n14902), .ZN(n7260) );
  NAND2_X1 U9139 ( .A1(n14942), .A2(n7258), .ZN(n7259) );
  NAND2_X1 U9140 ( .A1(n14954), .A2(n14953), .ZN(n14952) );
  NAND2_X1 U9141 ( .A1(n15237), .A2(n15238), .ZN(n15236) );
  XNOR2_X1 U9142 ( .A(n14914), .B(n7799), .ZN(n15246) );
  INV_X1 U9143 ( .A(n14915), .ZN(n7799) );
  NAND2_X1 U9144 ( .A1(n15246), .A2(n15449), .ZN(n15245) );
  NAND2_X1 U9145 ( .A1(n7788), .A2(n7786), .ZN(n7795) );
  INV_X1 U9146 ( .A(n15255), .ZN(n6841) );
  AOI21_X1 U9147 ( .B1(n7789), .B2(n7794), .A(n7787), .ZN(n7786) );
  INV_X1 U9148 ( .A(n14996), .ZN(n7123) );
  NOR2_X1 U9149 ( .A1(n9868), .A2(n13051), .ZN(P3_U3897) );
  INV_X1 U9150 ( .A(n7104), .ZN(n7103) );
  OAI21_X1 U9151 ( .B1(n12996), .B2(n15581), .A(n12246), .ZN(n7104) );
  NAND2_X1 U9152 ( .A1(n11132), .A2(n11131), .ZN(n11134) );
  NOR2_X1 U9153 ( .A1(n6806), .A2(n11015), .ZN(n11017) );
  AOI21_X1 U9154 ( .B1(n7256), .B2(n15681), .A(n7254), .ZN(n12707) );
  XNOR2_X1 U9155 ( .A(n7085), .B(n7084), .ZN(n12710) );
  AND2_X1 U9156 ( .A1(n7849), .A2(n8435), .ZN(n11947) );
  AOI211_X1 U9157 ( .C1(n15097), .C2(n11945), .A(n11944), .B(n11943), .ZN(
        n11946) );
  AOI21_X1 U9158 ( .B1(n11945), .B2(n8475), .A(n8474), .ZN(n8476) );
  AOI21_X1 U9159 ( .B1(n8426), .B2(n8475), .A(n7154), .ZN(n7153) );
  NOR2_X1 U9160 ( .A1(n15788), .A2(n12924), .ZN(n7154) );
  OAI211_X1 U9161 ( .C1(n7849), .C2(n15771), .A(n7847), .B(n8490), .ZN(
        P3_U3456) );
  AND2_X1 U9162 ( .A1(n8488), .A2(n8487), .ZN(n8490) );
  AOI21_X1 U9163 ( .B1(n8426), .B2(n8485), .A(n7156), .ZN(n7155) );
  NOR2_X1 U9164 ( .A1(n15773), .A2(n12992), .ZN(n7156) );
  OR2_X1 U9165 ( .A1(n15773), .A2(P3_REG0_REG_27__SCAN_IN), .ZN(n7096) );
  AND2_X1 U9166 ( .A1(n7353), .A2(n6716), .ZN(n15121) );
  NOR2_X1 U9167 ( .A1(n6786), .A2(n7824), .ZN(n7823) );
  NAND2_X1 U9168 ( .A1(n7826), .A2(n7828), .ZN(n7825) );
  NAND2_X1 U9169 ( .A1(n9950), .A2(n6802), .ZN(n9951) );
  OAI21_X1 U9170 ( .B1(n13625), .B2(n9175), .A(n6852), .ZN(P2_U3233) );
  AOI21_X1 U9171 ( .B1(n6854), .B2(n9175), .A(n6853), .ZN(n6852) );
  OAI21_X1 U9172 ( .B1(n15450), .B2(n8003), .A(n13626), .ZN(n6853) );
  NAND2_X1 U9173 ( .A1(n7739), .A2(n15576), .ZN(n7738) );
  INV_X1 U9174 ( .A(n7183), .ZN(n7182) );
  NAND2_X1 U9175 ( .A1(n7649), .A2(n13703), .ZN(n7739) );
  INV_X1 U9176 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n6922) );
  NAND2_X1 U9177 ( .A1(n7432), .A2(n6814), .ZN(P2_U3496) );
  NAND2_X1 U9178 ( .A1(n7433), .A2(n15561), .ZN(n7432) );
  INV_X1 U9179 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n7431) );
  NAND2_X1 U9180 ( .A1(n6943), .A2(n6939), .ZN(n14380) );
  NAND2_X1 U9181 ( .A1(n6945), .A2(n6944), .ZN(n6943) );
  NAND2_X1 U9182 ( .A1(n6941), .A2(n6940), .ZN(n6939) );
  OR2_X1 U9183 ( .A1(n7132), .A2(n7026), .ZN(n7025) );
  NAND2_X1 U9184 ( .A1(n7133), .A2(n15375), .ZN(n7132) );
  OAI21_X1 U9185 ( .B1(n14693), .B2(n15387), .A(n7082), .ZN(P1_U3525) );
  INV_X1 U9186 ( .A(n7083), .ZN(n7082) );
  AOI21_X1 U9187 ( .B1(n14692), .B2(n15386), .A(n14691), .ZN(n14693) );
  OAI21_X1 U9188 ( .B1(n14694), .B2(n7458), .A(n7461), .ZN(n7083) );
  INV_X1 U9189 ( .A(n7801), .ZN(n15796) );
  NOR2_X1 U9190 ( .A1(n15252), .A2(n15253), .ZN(n15251) );
  INV_X1 U9191 ( .A(n7797), .ZN(n15257) );
  OAI21_X1 U9192 ( .B1(n15252), .B2(n7794), .A(n7792), .ZN(n7797) );
  XNOR2_X1 U9193 ( .A(n15000), .B(n14999), .ZN(n7802) );
  XNOR2_X1 U9194 ( .A(n7914), .B(P3_ADDR_REG_19__SCAN_IN), .ZN(n14999) );
  NAND3_X1 U9195 ( .A1(n7124), .A2(n8028), .A3(n8027), .ZN(n10318) );
  NAND2_X1 U9196 ( .A1(n7857), .A2(n8401), .ZN(n7856) );
  AND2_X1 U9197 ( .A1(n7233), .A2(n13656), .ZN(n6673) );
  NOR2_X1 U9198 ( .A1(n15004), .A2(n7575), .ZN(n6674) );
  NAND2_X1 U9199 ( .A1(n13927), .A2(n13688), .ZN(n6675) );
  BUF_X1 U9200 ( .A(n9241), .Z(n9034) );
  INV_X2 U9201 ( .A(n9241), .ZN(n8565) );
  NAND2_X1 U9202 ( .A1(n8237), .A2(n7968), .ZN(n8251) );
  AND2_X1 U9203 ( .A1(n7587), .A2(n14043), .ZN(n6676) );
  NAND2_X1 U9204 ( .A1(n7130), .A2(n7129), .ZN(n12442) );
  OR2_X1 U9205 ( .A1(n12408), .A2(n7057), .ZN(n7056) );
  AND2_X1 U9206 ( .A1(n14468), .A2(n14414), .ZN(n6677) );
  INV_X1 U9207 ( .A(n12463), .ZN(n7376) );
  NOR2_X1 U9208 ( .A1(n11526), .A2(n7220), .ZN(n6678) );
  INV_X1 U9209 ( .A(n7856), .ZN(n7855) );
  NAND2_X1 U9210 ( .A1(n6833), .A2(n6785), .ZN(n6679) );
  XNOR2_X1 U9211 ( .A(n8009), .B(P3_IR_REG_29__SCAN_IN), .ZN(n8013) );
  NAND2_X1 U9212 ( .A1(n14773), .A2(n14395), .ZN(n6680) );
  AND2_X1 U9213 ( .A1(n8406), .A2(n7062), .ZN(n6681) );
  AND2_X1 U9214 ( .A1(n6761), .A2(n7306), .ZN(n6682) );
  INV_X1 U9215 ( .A(n12224), .ZN(n6985) );
  AND2_X1 U9216 ( .A1(n12631), .A2(n11120), .ZN(n6683) );
  INV_X1 U9217 ( .A(n8534), .ZN(n9158) );
  AND2_X1 U9218 ( .A1(n7474), .A2(n14394), .ZN(n6684) );
  NOR2_X1 U9219 ( .A1(n9292), .A2(n9291), .ZN(n6685) );
  NOR2_X1 U9220 ( .A1(n13971), .A2(n13675), .ZN(n6686) );
  AND2_X1 U9221 ( .A1(n11545), .A2(n6791), .ZN(n6687) );
  NAND2_X1 U9222 ( .A1(n7906), .A2(n6725), .ZN(n7904) );
  INV_X1 U9223 ( .A(n7904), .ZN(n7899) );
  AND2_X1 U9224 ( .A1(n8680), .A2(SI_7_), .ZN(n6688) );
  INV_X1 U9225 ( .A(P3_IR_REG_25__SCAN_IN), .ZN(n13374) );
  AND2_X1 U9226 ( .A1(n11006), .A2(n11005), .ZN(n6689) );
  AND2_X1 U9227 ( .A1(n14804), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n6690) );
  INV_X1 U9228 ( .A(n14579), .ZN(n7479) );
  INV_X1 U9229 ( .A(n13679), .ZN(n7745) );
  INV_X1 U9230 ( .A(n13673), .ZN(n13979) );
  NAND2_X1 U9231 ( .A1(n6783), .A2(n11882), .ZN(n11924) );
  NAND2_X1 U9232 ( .A1(n11619), .A2(n14205), .ZN(n7611) );
  INV_X1 U9233 ( .A(n13947), .ZN(n7233) );
  INV_X1 U9234 ( .A(n12483), .ZN(n7384) );
  AND2_X1 U9235 ( .A1(n9060), .A2(SI_24_), .ZN(n6691) );
  INV_X1 U9236 ( .A(n15548), .ZN(n15539) );
  OR2_X1 U9237 ( .A1(n13246), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n6692) );
  INV_X1 U9238 ( .A(n9175), .ZN(n10763) );
  NOR2_X1 U9239 ( .A1(n12421), .A2(n12514), .ZN(n6693) );
  XNOR2_X1 U9240 ( .A(n8578), .B(SI_2_), .ZN(n8577) );
  AND2_X1 U9241 ( .A1(n13979), .A2(n13672), .ZN(n6694) );
  OR2_X1 U9242 ( .A1(n8558), .A2(n9326), .ZN(n6695) );
  INV_X1 U9243 ( .A(n10132), .ZN(n7141) );
  AND2_X1 U9244 ( .A1(n13815), .A2(n13684), .ZN(n6696) );
  XNOR2_X1 U9245 ( .A(n13901), .B(n13115), .ZN(n13697) );
  INV_X1 U9246 ( .A(n13697), .ZN(n7425) );
  NAND2_X1 U9247 ( .A1(n7626), .A2(n13664), .ZN(n6697) );
  AND2_X1 U9248 ( .A1(n9316), .A2(n7683), .ZN(n6698) );
  AND2_X1 U9249 ( .A1(n13659), .A2(n13658), .ZN(n6699) );
  NAND2_X1 U9250 ( .A1(n9163), .A2(n9162), .ZN(n13632) );
  NAND3_X1 U9251 ( .A1(n8510), .A2(n8509), .A3(n8508), .ZN(n13578) );
  NOR2_X1 U9252 ( .A1(n13800), .A2(n7231), .ZN(n7230) );
  OAI211_X1 U9253 ( .C1(n9170), .C2(n9818), .A(n8538), .B(n6914), .ZN(n15498)
         );
  INV_X1 U9254 ( .A(n15498), .ZN(n7362) );
  INV_X1 U9255 ( .A(n10128), .ZN(n10435) );
  NOR2_X1 U9256 ( .A1(n14468), .A2(n14414), .ZN(n6700) );
  NOR2_X1 U9257 ( .A1(n14431), .A2(n7679), .ZN(n6701) );
  INV_X1 U9258 ( .A(n13641), .ZN(n7216) );
  NOR2_X1 U9259 ( .A1(n13725), .A2(n13666), .ZN(n6702) );
  INV_X1 U9260 ( .A(n14659), .ZN(n7476) );
  INV_X1 U9261 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n9336) );
  XOR2_X1 U9262 ( .A(n8698), .B(SI_8_), .Z(n6703) );
  AND2_X1 U9263 ( .A1(n7868), .A2(n7867), .ZN(n6704) );
  AND2_X1 U9264 ( .A1(n7476), .A2(n12147), .ZN(n6705) );
  NOR2_X1 U9265 ( .A1(n13958), .A2(n13680), .ZN(n6706) );
  NAND2_X1 U9266 ( .A1(n7349), .A2(n7347), .ZN(n13524) );
  AND2_X1 U9267 ( .A1(n10264), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n6707) );
  OR2_X1 U9268 ( .A1(n12634), .A2(n11041), .ZN(n12478) );
  OR2_X1 U9269 ( .A1(n7301), .A2(n7302), .ZN(n6708) );
  NAND2_X1 U9270 ( .A1(n9091), .A2(n9090), .ZN(n13927) );
  INV_X1 U9271 ( .A(n13927), .ZN(n7449) );
  AND2_X1 U9272 ( .A1(n14226), .A2(n11982), .ZN(n6709) );
  XNOR2_X1 U9273 ( .A(n12582), .B(n12722), .ZN(n12578) );
  INV_X1 U9274 ( .A(n10935), .ZN(n6868) );
  NAND2_X1 U9275 ( .A1(n11752), .A2(n11751), .ZN(n14724) );
  OR2_X1 U9276 ( .A1(n15549), .A2(n13568), .ZN(n6710) );
  OR2_X1 U9277 ( .A1(n15154), .A2(n13566), .ZN(n6711) );
  AND2_X1 U9278 ( .A1(n6669), .A2(n14265), .ZN(n6712) );
  AND2_X1 U9279 ( .A1(n12591), .A2(n12590), .ZN(n6713) );
  INV_X1 U9280 ( .A(n14450), .ZN(n7463) );
  NOR2_X1 U9281 ( .A1(n7392), .A2(n7396), .ZN(n8136) );
  NAND2_X1 U9282 ( .A1(n15584), .A2(n11377), .ZN(n11379) );
  AND2_X1 U9283 ( .A1(n6880), .A2(n6879), .ZN(n8683) );
  AND2_X1 U9284 ( .A1(n11229), .A2(n13568), .ZN(n6714) );
  NAND2_X1 U9285 ( .A1(n9043), .A2(n9042), .ZN(n13942) );
  INV_X1 U9286 ( .A(n13942), .ZN(n7451) );
  NAND2_X1 U9287 ( .A1(n12566), .A2(n6984), .ZN(n12769) );
  INV_X1 U9288 ( .A(n12769), .ZN(n7853) );
  INV_X1 U9289 ( .A(n11994), .ZN(n7307) );
  INV_X1 U9290 ( .A(n12008), .ZN(n7767) );
  INV_X1 U9291 ( .A(n11997), .ZN(n7782) );
  NAND2_X1 U9292 ( .A1(n11491), .A2(n11495), .ZN(n6715) );
  NAND2_X1 U9293 ( .A1(n11871), .A2(n11870), .ZN(n6716) );
  NAND2_X1 U9294 ( .A1(n11692), .A2(n11693), .ZN(n6717) );
  NAND2_X1 U9295 ( .A1(n8535), .A2(n9616), .ZN(n9170) );
  OR2_X1 U9296 ( .A1(n7449), .A2(n13688), .ZN(n6718) );
  NAND2_X1 U9297 ( .A1(n8506), .A2(n8505), .ZN(n14023) );
  NAND2_X1 U9298 ( .A1(n11949), .A2(n11948), .ZN(n14419) );
  INV_X1 U9299 ( .A(n12066), .ZN(n7301) );
  NOR2_X1 U9300 ( .A1(n14604), .A2(n7469), .ZN(n7468) );
  AND2_X1 U9301 ( .A1(n14514), .A2(n14443), .ZN(n6719) );
  AND2_X1 U9302 ( .A1(n15005), .A2(n12626), .ZN(n6720) );
  NAND2_X1 U9303 ( .A1(n11623), .A2(n11622), .ZN(n14773) );
  NAND2_X1 U9304 ( .A1(n8960), .A2(n8959), .ZN(n13965) );
  AND2_X1 U9305 ( .A1(n7839), .A2(n7836), .ZN(n6721) );
  AND3_X1 U9306 ( .A1(n7300), .A2(n7303), .A3(n14600), .ZN(n6722) );
  INV_X1 U9307 ( .A(n7699), .ZN(n7428) );
  NOR2_X1 U9308 ( .A1(n13718), .A2(n7701), .ZN(n7699) );
  NOR2_X1 U9309 ( .A1(n8845), .A2(n7749), .ZN(n7748) );
  AND2_X1 U9310 ( .A1(n13654), .A2(n13655), .ZN(n6723) );
  AND2_X1 U9311 ( .A1(n15530), .A2(n13570), .ZN(n6724) );
  AND2_X1 U9312 ( .A1(n9102), .A2(n9101), .ZN(n6725) );
  NOR2_X1 U9313 ( .A1(n10532), .A2(n7754), .ZN(n6726) );
  AND4_X1 U9314 ( .A1(n10047), .A2(n9304), .A3(n9303), .A4(n9302), .ZN(n6727)
         );
  OR2_X1 U9315 ( .A1(n8972), .A2(SI_18_), .ZN(n6728) );
  NAND2_X1 U9316 ( .A1(n9816), .A2(n8031), .ZN(n6729) );
  OR2_X1 U9317 ( .A1(n14825), .A2(n7806), .ZN(n6730) );
  OR2_X1 U9318 ( .A1(n14896), .A2(n13585), .ZN(n6731) );
  AND2_X1 U9319 ( .A1(n14660), .A2(n12025), .ZN(n12147) );
  AND4_X1 U9320 ( .A1(n8492), .A2(n6916), .A3(n7869), .A4(n8494), .ZN(n6732)
         );
  AND2_X1 U9321 ( .A1(n6885), .A2(n8840), .ZN(n6733) );
  INV_X1 U9322 ( .A(n13661), .ZN(n7630) );
  AND2_X1 U9323 ( .A1(n8398), .A2(n8397), .ZN(n6734) );
  AND2_X1 U9324 ( .A1(n8571), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n6735) );
  AND2_X1 U9325 ( .A1(n14567), .A2(n7481), .ZN(n6736) );
  AND2_X1 U9326 ( .A1(n12338), .A2(n12621), .ZN(n6737) );
  OR2_X1 U9327 ( .A1(n7227), .A2(n7225), .ZN(n6738) );
  AND3_X1 U9328 ( .A1(n8035), .A2(n8034), .A3(n8033), .ZN(n10316) );
  INV_X1 U9329 ( .A(n10316), .ZN(n7129) );
  NAND2_X1 U9330 ( .A1(n10092), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n10028) );
  OR2_X1 U9331 ( .A1(n13918), .A2(n13663), .ZN(n6739) );
  INV_X1 U9332 ( .A(n7599), .ZN(n7595) );
  NAND2_X1 U9333 ( .A1(n7604), .A2(n7602), .ZN(n7599) );
  OR2_X1 U9334 ( .A1(n12688), .A2(n12659), .ZN(n6740) );
  NAND2_X1 U9335 ( .A1(n8881), .A2(n8880), .ZN(n13673) );
  NOR2_X1 U9336 ( .A1(n15068), .A2(n12664), .ZN(n6741) );
  INV_X1 U9337 ( .A(n7288), .ZN(n7287) );
  OR2_X1 U9338 ( .A1(n12326), .A2(n7289), .ZN(n7288) );
  AND2_X1 U9339 ( .A1(n7694), .A2(n7693), .ZN(n6742) );
  AND2_X1 U9340 ( .A1(n12411), .A2(n12624), .ZN(n6743) );
  AND2_X1 U9341 ( .A1(n14079), .A2(n6717), .ZN(n7602) );
  AND2_X1 U9342 ( .A1(n11357), .A2(n11354), .ZN(n7616) );
  AND2_X1 U9343 ( .A1(n11518), .A2(n11517), .ZN(n6744) );
  OR2_X1 U9344 ( .A1(n14672), .A2(n15163), .ZN(n14394) );
  NOR2_X1 U9345 ( .A1(n13845), .A2(n13675), .ZN(n6745) );
  NOR2_X1 U9346 ( .A1(n12411), .A2(n12624), .ZN(n6746) );
  AND2_X1 U9347 ( .A1(n12381), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n6747) );
  AND2_X1 U9348 ( .A1(n13947), .A2(n13656), .ZN(n6748) );
  INV_X1 U9349 ( .A(n7358), .ZN(n7357) );
  OR2_X1 U9350 ( .A1(n11001), .A2(n7359), .ZN(n7358) );
  INV_X1 U9351 ( .A(n7701), .ZN(n7700) );
  NOR2_X1 U9352 ( .A1(n13695), .A2(n13694), .ZN(n7701) );
  AND2_X1 U9353 ( .A1(n6698), .A2(n7681), .ZN(n6749) );
  AND2_X1 U9354 ( .A1(n15110), .A2(n15013), .ZN(n6750) );
  OR2_X1 U9355 ( .A1(n7327), .A2(n7325), .ZN(n6751) );
  AND2_X1 U9356 ( .A1(n12487), .A2(n12486), .ZN(n12483) );
  INV_X1 U9357 ( .A(n12021), .ZN(n7773) );
  NAND2_X1 U9358 ( .A1(n11177), .A2(n11176), .ZN(n6752) );
  NOR2_X1 U9359 ( .A1(n15127), .A2(n13564), .ZN(n6753) );
  AND2_X1 U9360 ( .A1(n8744), .A2(SI_10_), .ZN(n6754) );
  AND2_X1 U9361 ( .A1(n8698), .A2(SI_8_), .ZN(n6755) );
  AND2_X1 U9362 ( .A1(n11996), .A2(n7782), .ZN(n6756) );
  INV_X1 U9363 ( .A(P3_IR_REG_17__SCAN_IN), .ZN(n7919) );
  INV_X1 U9364 ( .A(P3_IR_REG_26__SCAN_IN), .ZN(n13368) );
  INV_X1 U9365 ( .A(n7736), .ZN(n7242) );
  AND2_X1 U9366 ( .A1(n13673), .A2(n13674), .ZN(n7736) );
  AND2_X1 U9367 ( .A1(n8571), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n6757) );
  AND2_X1 U9368 ( .A1(n11911), .A2(n11910), .ZN(n6758) );
  INV_X1 U9369 ( .A(n7285), .ZN(n7284) );
  NAND2_X1 U9370 ( .A1(n7290), .A2(n7291), .ZN(n7285) );
  INV_X1 U9371 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n13054) );
  INV_X1 U9372 ( .A(n7561), .ZN(n7560) );
  OR2_X1 U9373 ( .A1(n12200), .A2(n7562), .ZN(n7561) );
  INV_X1 U9374 ( .A(n7593), .ZN(n7592) );
  AND2_X1 U9375 ( .A1(n12075), .A2(n7761), .ZN(n6759) );
  INV_X1 U9376 ( .A(n7011), .ZN(n8818) );
  AOI21_X1 U9377 ( .B1(n8796), .B2(n7913), .A(n7015), .ZN(n7011) );
  OR2_X1 U9378 ( .A1(n13810), .A2(n6921), .ZN(n6760) );
  OR2_X1 U9379 ( .A1(n7782), .A2(n11996), .ZN(n6761) );
  NAND2_X1 U9380 ( .A1(n14224), .A2(n10428), .ZN(n6762) );
  OAI21_X1 U9381 ( .B1(n13770), .B2(n7630), .A(n13662), .ZN(n7629) );
  OR2_X1 U9382 ( .A1(n14559), .A2(n14569), .ZN(n14403) );
  NAND2_X1 U9383 ( .A1(n6684), .A2(n14645), .ZN(n6763) );
  NAND2_X1 U9384 ( .A1(n12024), .A2(n7771), .ZN(n6764) );
  NOR2_X1 U9385 ( .A1(n14518), .A2(n7496), .ZN(n6765) );
  INV_X1 U9386 ( .A(n15256), .ZN(n7796) );
  AND2_X1 U9387 ( .A1(n7381), .A2(n7380), .ZN(n6766) );
  OR2_X1 U9388 ( .A1(n9012), .A2(n7882), .ZN(n6767) );
  INV_X1 U9389 ( .A(P3_IR_REG_4__SCAN_IN), .ZN(n7036) );
  AND2_X1 U9390 ( .A1(n7338), .A2(n7337), .ZN(n6768) );
  AND2_X1 U9391 ( .A1(n12550), .A2(n12551), .ZN(n12825) );
  INV_X1 U9392 ( .A(n12825), .ZN(n7058) );
  NOR2_X1 U9393 ( .A1(n12178), .A2(n12176), .ZN(n6769) );
  NOR2_X1 U9394 ( .A1(n15025), .A2(n12662), .ZN(n6770) );
  AND2_X1 U9395 ( .A1(n8657), .A2(SI_6_), .ZN(n6771) );
  INV_X1 U9396 ( .A(n7831), .ZN(n7830) );
  OAI21_X1 U9397 ( .B1(n13101), .B2(n7832), .A(n13112), .ZN(n7831) );
  NAND2_X1 U9398 ( .A1(n8562), .A2(n6850), .ZN(n6772) );
  AND2_X1 U9399 ( .A1(n14446), .A2(n14445), .ZN(n6773) );
  AND2_X1 U9400 ( .A1(n11893), .A2(n11892), .ZN(n6774) );
  AND2_X1 U9401 ( .A1(n6909), .A2(n9297), .ZN(n6775) );
  NOR2_X1 U9402 ( .A1(n7336), .A2(n6758), .ZN(n6776) );
  OR2_X1 U9403 ( .A1(n11991), .A2(n11989), .ZN(n6777) );
  OR2_X1 U9404 ( .A1(n7767), .A2(n12007), .ZN(n6778) );
  INV_X1 U9405 ( .A(n7340), .ZN(n7339) );
  NOR2_X1 U9406 ( .A1(n7341), .A2(n11908), .ZN(n7340) );
  NAND2_X1 U9407 ( .A1(n9310), .A2(n7617), .ZN(n6779) );
  NAND2_X1 U9408 ( .A1(n8794), .A2(n8795), .ZN(n6780) );
  INV_X1 U9409 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n8466) );
  INV_X1 U9410 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n13366) );
  INV_X1 U9411 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n7117) );
  INV_X1 U9412 ( .A(n7232), .ZN(n7225) );
  NAND2_X1 U9413 ( .A1(n7451), .A2(n13686), .ZN(n7232) );
  INV_X1 U9414 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n7158) );
  INV_X1 U9415 ( .A(n7837), .ZN(n7836) );
  OR2_X1 U9416 ( .A1(n13553), .A2(n7838), .ZN(n7837) );
  INV_X1 U9417 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n7269) );
  INV_X1 U9418 ( .A(P3_IR_REG_5__SCAN_IN), .ZN(n8096) );
  INV_X1 U9419 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n6850) );
  NAND2_X1 U9420 ( .A1(n10185), .A2(n9630), .ZN(n7915) );
  AND3_X1 U9421 ( .A1(n8683), .A2(n6876), .A3(n6875), .ZN(n8778) );
  INV_X1 U9422 ( .A(n14443), .ZN(n7177) );
  INV_X1 U9423 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n8699) );
  NAND2_X1 U9424 ( .A1(n12363), .A2(n12868), .ZN(n6781) );
  INV_X1 U9425 ( .A(n10021), .ZN(n8281) );
  NAND2_X1 U9426 ( .A1(n11461), .A2(n6705), .ZN(n7473) );
  INV_X1 U9427 ( .A(n11945), .ZN(n8478) );
  NAND2_X1 U9428 ( .A1(n7543), .A2(n8004), .ZN(n11945) );
  NOR2_X1 U9429 ( .A1(n14111), .A2(n14112), .ZN(n14110) );
  NAND2_X1 U9430 ( .A1(n11806), .A2(n11805), .ZN(n14705) );
  INV_X1 U9431 ( .A(n14705), .ZN(n7519) );
  NAND2_X1 U9432 ( .A1(n8335), .A2(n8334), .ZN(n12318) );
  INV_X1 U9433 ( .A(n12318), .ZN(n6986) );
  AOI21_X1 U9434 ( .B1(n7230), .B2(n6696), .A(n6673), .ZN(n7229) );
  INV_X1 U9435 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n9707) );
  AND2_X1 U9436 ( .A1(n7959), .A2(P2_DATAO_REG_13__SCAN_IN), .ZN(n6782) );
  AOI21_X1 U9437 ( .B1(n13059), .B2(n12394), .A(n8383), .ZN(n12993) );
  INV_X1 U9438 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n6957) );
  AND2_X1 U9439 ( .A1(n11881), .A2(n13503), .ZN(n6783) );
  AND2_X1 U9440 ( .A1(n14284), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6784) );
  XOR2_X1 U9441 ( .A(n12563), .B(n12234), .Z(n6785) );
  INV_X1 U9442 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n6846) );
  NAND2_X1 U9443 ( .A1(n9000), .A2(n8999), .ZN(n13953) );
  AND2_X1 U9444 ( .A1(n13715), .A2(n15125), .ZN(n6786) );
  INV_X1 U9445 ( .A(n12520), .ZN(n7408) );
  NAND2_X1 U9446 ( .A1(n7606), .A2(n11601), .ZN(n15165) );
  OR2_X1 U9447 ( .A1(n9716), .A2(n15396), .ZN(n6787) );
  AND2_X1 U9448 ( .A1(n9018), .A2(n7719), .ZN(n6788) );
  AND2_X1 U9449 ( .A1(n13901), .A2(n15539), .ZN(n6789) );
  NAND2_X1 U9450 ( .A1(n7448), .A2(n6918), .ZN(n6919) );
  INV_X1 U9451 ( .A(n7452), .ZN(n13796) );
  NAND2_X1 U9452 ( .A1(n14670), .A2(n7515), .ZN(n6790) );
  INV_X1 U9453 ( .A(n7448), .ZN(n13885) );
  NOR2_X1 U9454 ( .A1(n13884), .A2(n13985), .ZN(n7448) );
  NAND2_X1 U9455 ( .A1(n11573), .A2(n11574), .ZN(n6791) );
  INV_X1 U9456 ( .A(P3_ADDR_REG_4__SCAN_IN), .ZN(n7806) );
  AND2_X1 U9457 ( .A1(n12206), .A2(n12626), .ZN(n6792) );
  NOR2_X1 U9458 ( .A1(n13891), .A2(n13670), .ZN(n6793) );
  INV_X1 U9459 ( .A(n7056), .ZN(n7055) );
  AND2_X1 U9460 ( .A1(n7286), .A2(n7284), .ZN(n6794) );
  AND2_X1 U9461 ( .A1(n11323), .A2(n11324), .ZN(n6795) );
  AND2_X1 U9462 ( .A1(n12201), .A2(n12627), .ZN(n6796) );
  INV_X1 U9463 ( .A(n7611), .ZN(n7610) );
  NAND2_X1 U9464 ( .A1(n7994), .A2(n11920), .ZN(n6797) );
  INV_X1 U9465 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n6859) );
  INV_X1 U9466 ( .A(n11612), .ZN(n6865) );
  AND2_X1 U9467 ( .A1(n9548), .A2(P2_DATAO_REG_11__SCAN_IN), .ZN(n6798) );
  AND2_X1 U9468 ( .A1(n7957), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n6799) );
  INV_X1 U9469 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n10414) );
  INV_X1 U9470 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n7532) );
  NOR2_X1 U9471 ( .A1(n8220), .A2(n7540), .ZN(n7539) );
  AOI21_X1 U9472 ( .B1(n7961), .B2(n7539), .A(n7538), .ZN(n7537) );
  NAND2_X1 U9473 ( .A1(n9553), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n6800) );
  INV_X1 U9474 ( .A(n7743), .ZN(n7438) );
  NAND2_X1 U9475 ( .A1(n13965), .A2(n7745), .ZN(n7743) );
  INV_X1 U9476 ( .A(n15403), .ZN(n7026) );
  NAND2_X1 U9477 ( .A1(n10072), .A2(n13865), .ZN(n13852) );
  INV_X1 U9478 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6979) );
  AND2_X1 U9479 ( .A1(n12655), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n6801) );
  OR2_X1 U9480 ( .A1(n8202), .A2(n8201), .ZN(n15655) );
  OR2_X1 U9481 ( .A1(n13542), .A2(n7705), .ZN(n6802) );
  XNOR2_X1 U9482 ( .A(n12656), .B(n12682), .ZN(n15616) );
  INV_X1 U9483 ( .A(n12260), .ZN(n7289) );
  NAND2_X1 U9484 ( .A1(n6932), .A2(n6930), .ZN(n12654) );
  NAND2_X1 U9485 ( .A1(n8138), .A2(n7861), .ZN(n6803) );
  NAND2_X1 U9486 ( .A1(n7859), .A2(n8138), .ZN(n6804) );
  NOR2_X1 U9487 ( .A1(n15615), .A2(n12657), .ZN(n6805) );
  NOR2_X1 U9488 ( .A1(n15601), .A2(n15600), .ZN(n6806) );
  INV_X1 U9489 ( .A(n7527), .ZN(n7526) );
  NOR2_X1 U9490 ( .A1(n7971), .A2(n7528), .ZN(n7527) );
  INV_X1 U9491 ( .A(n13656), .ZN(n13685) );
  INV_X1 U9492 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n8525) );
  NOR2_X1 U9493 ( .A1(n7735), .A2(n7732), .ZN(n6807) );
  INV_X1 U9494 ( .A(n13084), .ZN(n7350) );
  AND2_X1 U9495 ( .A1(n7648), .A2(n7647), .ZN(n6808) );
  NOR2_X1 U9496 ( .A1(n15403), .A2(n7125), .ZN(n6809) );
  AND2_X1 U9497 ( .A1(n8778), .A2(n7840), .ZN(n9279) );
  AND2_X1 U9498 ( .A1(n9063), .A2(n11167), .ZN(n6810) );
  AND2_X1 U9499 ( .A1(n11151), .A2(n8400), .ZN(n6811) );
  AND2_X1 U9500 ( .A1(n7708), .A2(n9083), .ZN(n6812) );
  AND2_X1 U9501 ( .A1(n9900), .A2(n9899), .ZN(n15576) );
  NAND2_X1 U9502 ( .A1(n8636), .A2(n8635), .ZN(n15513) );
  INV_X1 U9503 ( .A(n15513), .ZN(n7435) );
  AND2_X2 U9504 ( .A1(n10655), .A2(n8473), .ZN(n15788) );
  AND2_X2 U9505 ( .A1(n8484), .A2(n12610), .ZN(n15773) );
  OR2_X1 U9506 ( .A1(n10263), .A2(n10262), .ZN(n7695) );
  INV_X1 U9507 ( .A(n12699), .ZN(n7689) );
  AND2_X2 U9508 ( .A1(n12613), .A2(n10656), .ZN(n12593) );
  NAND2_X1 U9509 ( .A1(n9949), .A2(n9948), .ZN(n6813) );
  NAND2_X1 U9510 ( .A1(n8688), .A2(n8687), .ZN(n15530) );
  INV_X1 U9511 ( .A(n15530), .ZN(n7447) );
  OR2_X1 U9512 ( .A1(n15561), .A2(n7431), .ZN(n6814) );
  INV_X1 U9513 ( .A(n15053), .ZN(n7691) );
  INV_X1 U9514 ( .A(SI_22_), .ZN(n7719) );
  OR2_X1 U9515 ( .A1(n14364), .A2(n14365), .ZN(n6815) );
  OR2_X1 U9516 ( .A1(n14353), .A2(n14354), .ZN(n6816) );
  OR2_X1 U9517 ( .A1(n15561), .A2(n6922), .ZN(n6817) );
  AND2_X1 U9518 ( .A1(n7695), .A2(n7694), .ZN(n6818) );
  AND2_X1 U9519 ( .A1(n15766), .A2(n15765), .ZN(n15106) );
  INV_X1 U9520 ( .A(SI_26_), .ZN(n11425) );
  AND2_X1 U9521 ( .A1(n7981), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n6819) );
  INV_X1 U9522 ( .A(n9485), .ZN(n6847) );
  INV_X1 U9523 ( .A(n14299), .ZN(n6958) );
  INV_X1 U9524 ( .A(n14372), .ZN(n7164) );
  INV_X1 U9525 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n12670) );
  INV_X1 U9526 ( .A(n14612), .ZN(n7108) );
  AND2_X1 U9527 ( .A1(n9762), .A2(n9761), .ZN(n15351) );
  INV_X1 U9528 ( .A(n12706), .ZN(n12666) );
  AND2_X1 U9529 ( .A1(n7927), .A2(n7926), .ZN(n12706) );
  AND2_X1 U9530 ( .A1(n13246), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n6820) );
  INV_X1 U9531 ( .A(n6947), .ZN(n14283) );
  OAI21_X1 U9532 ( .B1(n14253), .B2(n6949), .A(n6948), .ZN(n6947) );
  NAND2_X1 U9533 ( .A1(n7075), .A2(n8440), .ZN(n7078) );
  INV_X1 U9534 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n14877) );
  INV_X1 U9535 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n7179) );
  INV_X1 U9536 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n6982) );
  INV_X1 U9537 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n7501) );
  OAI21_X2 U9538 ( .B1(n12308), .B2(n6825), .A(n6822), .ZN(n12214) );
  NAND2_X1 U9539 ( .A1(n8138), .A2(n6826), .ZN(n8239) );
  OAI21_X1 U9540 ( .B1(n15584), .B2(n6829), .A(n6827), .ZN(n12194) );
  NAND2_X1 U9541 ( .A1(n12297), .A2(n12233), .ZN(n12354) );
  INV_X1 U9542 ( .A(n12365), .ZN(n12202) );
  NAND2_X1 U9543 ( .A1(n6831), .A2(n7573), .ZN(n12310) );
  XNOR2_X2 U9544 ( .A(n6834), .B(n8005), .ZN(n8427) );
  NOR2_X1 U9545 ( .A1(n14925), .A2(n14924), .ZN(n14923) );
  NOR2_X1 U9546 ( .A1(n15804), .A2(n15805), .ZN(n15803) );
  NOR2_X1 U9547 ( .A1(n14949), .A2(n14904), .ZN(n14905) );
  OAI211_X1 U9548 ( .C1(n14949), .C2(n6840), .A(n6839), .B(n6838), .ZN(n14954)
         );
  NAND2_X1 U9549 ( .A1(n14949), .A2(n14906), .ZN(n6838) );
  NAND2_X1 U9550 ( .A1(n14904), .A2(n14906), .ZN(n6839) );
  OR2_X1 U9551 ( .A1(n14904), .A2(n14906), .ZN(n6840) );
  NAND2_X1 U9552 ( .A1(n15242), .A2(n15240), .ZN(n14914) );
  XNOR2_X1 U9553 ( .A(n6842), .B(n7802), .ZN(SUB_1596_U4) );
  NAND2_X1 U9554 ( .A1(n6843), .A2(n14998), .ZN(n6842) );
  NAND2_X1 U9555 ( .A1(n14996), .A2(n14997), .ZN(n14998) );
  AND2_X2 U9556 ( .A1(n6860), .A2(n6859), .ZN(n8562) );
  OAI211_X1 U9557 ( .C1(n6870), .C2(n6868), .A(n6869), .B(n11268), .ZN(n11271)
         );
  NAND2_X1 U9558 ( .A1(n10936), .A2(n10935), .ZN(n11269) );
  NAND2_X1 U9559 ( .A1(n6870), .A2(n10926), .ZN(n10936) );
  NAND3_X1 U9560 ( .A1(n7779), .A2(n7780), .A3(n10230), .ZN(n10719) );
  NAND4_X1 U9561 ( .A1(n7779), .A2(n7780), .A3(n10230), .A4(n6874), .ZN(n9612)
         );
  NAND2_X2 U9562 ( .A1(n9996), .A2(n12130), .ZN(n15320) );
  NOR2_X1 U9563 ( .A1(n8910), .A2(n8843), .ZN(n6884) );
  INV_X1 U9564 ( .A(n8910), .ZN(n6885) );
  NAND2_X1 U9565 ( .A1(n8568), .A2(n6887), .ZN(n8569) );
  INV_X1 U9566 ( .A(n8570), .ZN(n6888) );
  AND2_X1 U9567 ( .A1(n8566), .A2(n8567), .ZN(n8570) );
  NAND2_X1 U9568 ( .A1(n6892), .A2(n6889), .ZN(n8842) );
  NAND3_X1 U9569 ( .A1(n8768), .A2(n8767), .A3(n6780), .ZN(n6895) );
  NAND2_X1 U9570 ( .A1(n6898), .A2(n6897), .ZN(n6896) );
  INV_X1 U9571 ( .A(n8971), .ZN(n6897) );
  INV_X1 U9572 ( .A(n6902), .ZN(n6898) );
  NAND2_X1 U9573 ( .A1(n6901), .A2(n6900), .ZN(n6899) );
  NAND2_X1 U9574 ( .A1(n6902), .A2(n8971), .ZN(n6901) );
  NAND2_X1 U9575 ( .A1(n8949), .A2(n8948), .ZN(n6902) );
  NAND3_X1 U9576 ( .A1(n8653), .A2(n8652), .A3(n8676), .ZN(n6903) );
  NAND3_X1 U9577 ( .A1(n6905), .A2(n6904), .A3(n6903), .ZN(n8697) );
  NAND3_X1 U9578 ( .A1(n8653), .A2(n8652), .A3(n8674), .ZN(n6905) );
  OAI211_X1 U9579 ( .C1(n6775), .C2(n6908), .A(n6907), .B(n6685), .ZN(P2_U3328) );
  OAI21_X1 U9580 ( .B1(n6909), .B2(n9247), .A(n7911), .ZN(n6907) );
  OAI21_X1 U9581 ( .B1(n6909), .B2(n9295), .A(n11245), .ZN(n6908) );
  NAND2_X1 U9582 ( .A1(n9058), .A2(n7874), .ZN(n7873) );
  NAND2_X1 U9583 ( .A1(n6911), .A2(n6910), .ZN(n9058) );
  OR2_X1 U9584 ( .A1(n9037), .A2(n9036), .ZN(n6910) );
  NAND2_X1 U9585 ( .A1(n6912), .A2(n7081), .ZN(n6911) );
  NAND2_X1 U9586 ( .A1(n9037), .A2(n9036), .ZN(n6912) );
  OR2_X2 U9587 ( .A1(n10248), .A2(n10543), .ZN(n10575) );
  NOR2_X2 U9588 ( .A1(n10296), .A2(n6989), .ZN(n9909) );
  NAND4_X1 U9589 ( .A1(n6732), .A2(n6915), .A3(n7638), .A4(n7841), .ZN(n6917)
         );
  INV_X1 U9590 ( .A(n6919), .ZN(n13844) );
  NOR2_X1 U9591 ( .A1(n13810), .A2(n13947), .ZN(n7452) );
  NAND2_X1 U9592 ( .A1(n6923), .A2(n6817), .ZN(P2_U3497) );
  NAND2_X1 U9593 ( .A1(n14001), .A2(n15561), .ZN(n6923) );
  OAI21_X1 U9594 ( .B1(n13899), .B2(n15548), .A(n13897), .ZN(n6925) );
  NOR2_X1 U9595 ( .A1(n10026), .A2(n10027), .ZN(n10030) );
  AOI21_X1 U9596 ( .B1(n8326), .B2(n8325), .A(n6819), .ZN(n7982) );
  NAND2_X1 U9597 ( .A1(n8304), .A2(n7979), .ZN(n8315) );
  AOI21_X2 U9598 ( .B1(n15760), .B2(n12925), .A(n6988), .ZN(n12927) );
  NAND3_X1 U9599 ( .A1(n7366), .A2(n8367), .A3(n7365), .ZN(n12738) );
  INV_X1 U9600 ( .A(n6989), .ZN(n10668) );
  NAND2_X1 U9601 ( .A1(n6989), .A2(n8565), .ZN(n8566) );
  NAND2_X1 U9602 ( .A1(n6989), .A2(n9034), .ZN(n8568) );
  NAND2_X1 U9603 ( .A1(n9905), .A2(n6989), .ZN(n9903) );
  NAND2_X1 U9604 ( .A1(n10296), .A2(n6989), .ZN(n9796) );
  XNOR2_X1 U9605 ( .A(n6989), .B(n13576), .ZN(n9901) );
  INV_X1 U9606 ( .A(n11902), .ZN(n11900) );
  NAND2_X1 U9607 ( .A1(n13516), .A2(n6774), .ZN(n6990) );
  NAND2_X1 U9608 ( .A1(n13517), .A2(n13518), .ZN(n13516) );
  AND2_X2 U9609 ( .A1(n6991), .A2(n6776), .ZN(n13062) );
  NAND3_X1 U9610 ( .A1(n13533), .A2(n11905), .A3(n7340), .ZN(n6991) );
  NAND2_X2 U9611 ( .A1(n11935), .A2(n6992), .ZN(n13533) );
  AND2_X2 U9612 ( .A1(n11904), .A2(n11903), .ZN(n11935) );
  INV_X1 U9613 ( .A(n7345), .ZN(n6999) );
  NAND2_X1 U9614 ( .A1(n7351), .A2(n7344), .ZN(n6998) );
  XNOR2_X2 U9615 ( .A(n13065), .B(n7001), .ZN(n7351) );
  NAND2_X1 U9616 ( .A1(n6999), .A2(n6998), .ZN(n13495) );
  INV_X1 U9617 ( .A(n7351), .ZN(n13085) );
  INV_X1 U9618 ( .A(n13066), .ZN(n7001) );
  NAND3_X1 U9619 ( .A1(n8778), .A2(n7755), .A3(n8495), .ZN(n7004) );
  NAND2_X1 U9620 ( .A1(n8679), .A2(n7712), .ZN(n7710) );
  AOI21_X1 U9621 ( .B1(n8655), .B2(n7006), .A(n6771), .ZN(n7005) );
  INV_X1 U9622 ( .A(n8633), .ZN(n7006) );
  NAND2_X1 U9623 ( .A1(n9061), .A2(n6691), .ZN(n7707) );
  NAND2_X1 U9624 ( .A1(n7007), .A2(n6810), .ZN(n7706) );
  NAND2_X1 U9625 ( .A1(n7007), .A2(n9063), .ZN(n9084) );
  INV_X1 U9626 ( .A(n7008), .ZN(n8868) );
  NAND2_X1 U9627 ( .A1(n8724), .A2(n7017), .ZN(n7016) );
  NAND2_X1 U9628 ( .A1(n7025), .A2(n7021), .ZN(P1_U3557) );
  NAND2_X1 U9629 ( .A1(n14692), .A2(n7024), .ZN(n7023) );
  NAND2_X1 U9630 ( .A1(n8894), .A2(n8893), .ZN(n8875) );
  NAND2_X1 U9631 ( .A1(n7034), .A2(n6773), .ZN(n14481) );
  NOR2_X1 U9632 ( .A1(n8014), .A2(n7041), .ZN(n7042) );
  OAI21_X1 U9633 ( .B1(n12816), .B2(n7052), .A(n7051), .ZN(n8416) );
  NAND2_X1 U9634 ( .A1(n8404), .A2(n6681), .ZN(n7060) );
  NAND2_X1 U9635 ( .A1(n7060), .A2(n7061), .ZN(n12891) );
  OAI21_X1 U9636 ( .B1(n7079), .B2(n7069), .A(n7067), .ZN(n12853) );
  NAND2_X1 U9637 ( .A1(n7066), .A2(n7064), .ZN(n8412) );
  NAND2_X1 U9638 ( .A1(n7079), .A2(n7067), .ZN(n7066) );
  OAI21_X1 U9639 ( .B1(n12842), .B2(n7865), .A(n7863), .ZN(n12816) );
  NAND2_X1 U9640 ( .A1(n7845), .A2(n7843), .ZN(n11852) );
  NAND2_X1 U9641 ( .A1(n12891), .A2(n12894), .ZN(n7079) );
  NAND2_X1 U9642 ( .A1(n11051), .A2(n8399), .ZN(n11152) );
  NAND2_X1 U9643 ( .A1(n10726), .A2(n6734), .ZN(n11051) );
  NAND2_X1 U9644 ( .A1(n8392), .A2(n10312), .ZN(n15693) );
  INV_X2 U9645 ( .A(n7621), .ZN(n8553) );
  OAI21_X1 U9646 ( .B1(n8947), .B2(n8946), .A(n8945), .ZN(n8949) );
  NAND2_X1 U9647 ( .A1(n7112), .A2(n7109), .ZN(n8607) );
  INV_X1 U9648 ( .A(n7170), .ZN(n7169) );
  OAI21_X1 U9649 ( .B1(n7080), .B2(n7891), .A(n7890), .ZN(n8649) );
  OAI21_X1 U9650 ( .B1(n7883), .B2(n7146), .A(n8721), .ZN(n8740) );
  OAI22_X1 U9651 ( .A1(n8992), .A2(n7171), .B1(n7881), .B2(n9013), .ZN(n9037)
         );
  NAND2_X1 U9652 ( .A1(n7150), .A2(n7149), .ZN(n7112) );
  AOI21_X1 U9653 ( .B1(n8607), .B2(n8606), .A(n8605), .ZN(n7080) );
  NAND2_X1 U9654 ( .A1(n9979), .A2(n9978), .ZN(n10126) );
  AOI21_X1 U9655 ( .B1(n7656), .B2(n7654), .A(n6709), .ZN(n10585) );
  BUF_X8 U9656 ( .A(n10117), .Z(n11839) );
  NAND2_X1 U9657 ( .A1(n8068), .A2(n8067), .ZN(n7535) );
  INV_X1 U9658 ( .A(n8382), .ZN(n7152) );
  NAND2_X1 U9659 ( .A1(n7947), .A2(n7946), .ZN(n8112) );
  NAND2_X1 U9660 ( .A1(n7090), .A2(n7951), .ZN(n8135) );
  OAI21_X1 U9661 ( .B1(n8315), .B2(n8314), .A(n7980), .ZN(n8326) );
  NAND2_X1 U9662 ( .A1(n7544), .A2(n7994), .ZN(n7543) );
  NAND2_X1 U9663 ( .A1(n8125), .A2(n8124), .ZN(n7090) );
  NAND2_X1 U9664 ( .A1(n12607), .A2(n7548), .ZN(n7547) );
  NAND3_X1 U9665 ( .A1(n7094), .A2(n7229), .A3(n7232), .ZN(n7224) );
  OAI21_X1 U9666 ( .B1(n9147), .B2(n13471), .A(n9146), .ZN(n9149) );
  INV_X1 U9667 ( .A(n7368), .ZN(n7367) );
  NAND2_X1 U9668 ( .A1(n7137), .A2(n7537), .ZN(n7967) );
  NAND2_X1 U9669 ( .A1(n7097), .A2(n7096), .ZN(n12995) );
  OR2_X1 U9670 ( .A1(n12994), .A2(n15771), .ZN(n7097) );
  NAND2_X1 U9671 ( .A1(n7536), .A2(n7945), .ZN(n8095) );
  NAND2_X1 U9672 ( .A1(n7535), .A2(n7533), .ZN(n7536) );
  NAND2_X1 U9673 ( .A1(n7942), .A2(n7941), .ZN(n8068) );
  OAI21_X1 U9674 ( .B1(n12605), .B2(n7547), .A(n7546), .ZN(n7545) );
  NAND2_X1 U9675 ( .A1(n8292), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n7977) );
  NAND2_X1 U9676 ( .A1(n8207), .A2(n7539), .ZN(n7137) );
  NAND2_X1 U9677 ( .A1(n7940), .A2(n7939), .ZN(n8053) );
  OAI21_X1 U9678 ( .B1(n14679), .B2(n14386), .A(n7144), .ZN(n12139) );
  NAND2_X1 U9679 ( .A1(n8346), .A2(n7984), .ZN(n7986) );
  MUX2_X1 U9680 ( .A(n12181), .B(n12180), .S(n12179), .Z(n12182) );
  NAND2_X1 U9681 ( .A1(n7395), .A2(n7250), .ZN(n8438) );
  NAND2_X1 U9682 ( .A1(n11731), .A2(n11286), .ZN(n11733) );
  NAND2_X1 U9683 ( .A1(n7181), .A2(n8619), .ZN(n8631) );
  NAND2_X1 U9684 ( .A1(n7710), .A2(n7711), .ZN(n8724) );
  NAND2_X1 U9685 ( .A1(n7161), .A2(n7756), .ZN(n12094) );
  NAND2_X1 U9686 ( .A1(n7098), .A2(n7785), .ZN(n12105) );
  NAND2_X1 U9687 ( .A1(n12084), .A2(n12083), .ZN(n12086) );
  NAND2_X1 U9688 ( .A1(n7757), .A2(n12074), .ZN(n7322) );
  NAND2_X1 U9689 ( .A1(n12094), .A2(n12095), .ZN(n12093) );
  NAND3_X1 U9690 ( .A1(n12099), .A2(n7783), .A3(n12098), .ZN(n7098) );
  NAND3_X1 U9691 ( .A1(n7415), .A2(n7416), .A3(n8596), .ZN(n7131) );
  AND2_X2 U9692 ( .A1(n7100), .A2(n7099), .ZN(n12124) );
  INV_X1 U9693 ( .A(n12106), .ZN(n7100) );
  INV_X1 U9694 ( .A(n10318), .ZN(n7130) );
  NAND2_X1 U9695 ( .A1(n7105), .A2(n7103), .ZN(P3_U3154) );
  NAND2_X1 U9696 ( .A1(n12239), .A2(n15021), .ZN(n7105) );
  XNOR2_X1 U9697 ( .A(n12172), .B(n7108), .ZN(n7107) );
  INV_X1 U9698 ( .A(n9639), .ZN(n9293) );
  NAND2_X1 U9699 ( .A1(n8627), .A2(n8628), .ZN(n7145) );
  OAI22_X1 U9700 ( .A1(n8740), .A2(n7907), .B1(n8738), .B2(n8739), .ZN(n8763)
         );
  NAND4_X1 U9701 ( .A1(n8003), .A2(n8002), .A3(n7444), .A4(
        P3_ADDR_REG_19__SCAN_IN), .ZN(n7443) );
  INV_X1 U9702 ( .A(n8587), .ZN(n7111) );
  NAND2_X1 U9703 ( .A1(n7115), .A2(n6671), .ZN(n7113) );
  INV_X1 U9704 ( .A(n9982), .ZN(n7115) );
  NAND2_X1 U9705 ( .A1(n8504), .A2(P2_IR_REG_29__SCAN_IN), .ZN(n7118) );
  NOR2_X1 U9706 ( .A1(n12135), .A2(n7119), .ZN(n12185) );
  INV_X1 U9707 ( .A(n8628), .ZN(n7892) );
  NAND2_X1 U9708 ( .A1(n14435), .A2(n12164), .ZN(n14753) );
  NOR2_X1 U9709 ( .A1(n9922), .A2(n9921), .ZN(n9920) );
  NOR2_X1 U9710 ( .A1(n10495), .A2(n10494), .ZN(n10498) );
  AOI21_X1 U9711 ( .B1(n10954), .B2(n15210), .A(n10953), .ZN(n11215) );
  NOR3_X1 U9712 ( .A1(n14236), .A2(n9709), .A3(n14247), .ZN(n14235) );
  XNOR2_X1 U9713 ( .A(n7120), .B(P2_ADDR_REG_18__SCAN_IN), .ZN(SUB_1596_U62)
         );
  NAND2_X1 U9714 ( .A1(n14998), .A2(n7121), .ZN(n7120) );
  NAND2_X1 U9715 ( .A1(n7123), .A2(n7122), .ZN(n7121) );
  INV_X1 U9716 ( .A(n14997), .ZN(n7122) );
  NOR2_X2 U9717 ( .A1(n14911), .A2(n14910), .ZN(n15241) );
  NAND2_X1 U9718 ( .A1(n7738), .A2(n7182), .ZN(P2_U3528) );
  NAND2_X1 U9719 ( .A1(n10585), .A2(n10586), .ZN(n10584) );
  OAI21_X1 U9720 ( .B1(n8991), .B2(n8990), .A(n6767), .ZN(n7171) );
  NAND2_X2 U9721 ( .A1(n7443), .A2(n7441), .ZN(n8534) );
  INV_X1 U9722 ( .A(n12076), .ZN(n7761) );
  NAND2_X1 U9723 ( .A1(n8416), .A2(n8415), .ZN(n12781) );
  NOR2_X1 U9724 ( .A1(n7762), .A2(n7758), .ZN(n7757) );
  AOI21_X1 U9725 ( .B1(n12127), .B2(n12126), .A(n12125), .ZN(n12135) );
  NAND2_X1 U9726 ( .A1(n11478), .A2(n11477), .ZN(n14970) );
  INV_X1 U9727 ( .A(n10428), .ZN(n7673) );
  NAND2_X1 U9728 ( .A1(n9831), .A2(n9832), .ZN(n10008) );
  AND2_X1 U9729 ( .A1(n9830), .A2(n10007), .ZN(n9831) );
  NAND2_X1 U9730 ( .A1(n9824), .A2(n9825), .ZN(n9826) );
  INV_X4 U9731 ( .A(n11722), .ZN(n11832) );
  NAND2_X1 U9732 ( .A1(n14192), .A2(n11803), .ZN(n14042) );
  INV_X1 U9733 ( .A(n10925), .ZN(n7607) );
  NAND2_X1 U9734 ( .A1(n7367), .A2(n7369), .ZN(n7365) );
  OAI211_X4 U9735 ( .C1(n6667), .C2(n9460), .A(n7776), .B(n9816), .ZN(n12109)
         );
  OAI21_X1 U9736 ( .B1(n12568), .B2(n7369), .A(n12757), .ZN(n7368) );
  INV_X1 U9737 ( .A(n7143), .ZN(n14429) );
  NAND2_X1 U9738 ( .A1(n14425), .A2(n14424), .ZN(n14630) );
  OAI21_X2 U9739 ( .B1(n14732), .B2(n7686), .A(n7684), .ZN(n14488) );
  NAND2_X1 U9740 ( .A1(n9556), .A2(n7158), .ZN(n14795) );
  NAND2_X1 U9741 ( .A1(n11915), .A2(n7809), .ZN(n13063) );
  NAND2_X1 U9742 ( .A1(n13092), .A2(n13091), .ZN(n13090) );
  INV_X1 U9743 ( .A(n9648), .ZN(n9645) );
  OAI21_X1 U9744 ( .B1(n14429), .B2(n7678), .A(n7676), .ZN(n14434) );
  INV_X1 U9745 ( .A(n12157), .ZN(n7671) );
  NAND2_X1 U9746 ( .A1(n13773), .A2(n13772), .ZN(n13771) );
  INV_X4 U9747 ( .A(n8534), .ZN(n9616) );
  OAI21_X1 U9748 ( .B1(n8607), .B2(n8606), .A(n7145), .ZN(n7891) );
  INV_X1 U9749 ( .A(n7413), .ZN(n8576) );
  NAND2_X1 U9750 ( .A1(n7167), .A2(n7166), .ZN(n9246) );
  NOR2_X2 U9751 ( .A1(n13760), .A2(n13918), .ZN(n13744) );
  NAND2_X1 U9752 ( .A1(n8587), .A2(n8586), .ZN(n7150) );
  NAND2_X1 U9753 ( .A1(n12079), .A2(n12080), .ZN(n12078) );
  NAND2_X1 U9754 ( .A1(n7321), .A2(n7322), .ZN(n12079) );
  NAND3_X1 U9755 ( .A1(n7316), .A2(n7314), .A3(n7162), .ZN(n7161) );
  NAND2_X1 U9756 ( .A1(n7545), .A2(n12614), .ZN(P3_U3296) );
  OAI21_X1 U9757 ( .B1(n12991), .B2(n15786), .A(n7153), .ZN(P3_U3487) );
  OAI21_X1 U9758 ( .B1(n12991), .B2(n15771), .A(n7155), .ZN(P3_U3455) );
  INV_X1 U9759 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n7683) );
  AOI21_X1 U9760 ( .B1(n7672), .B2(n7674), .A(n7671), .ZN(n7670) );
  NAND2_X1 U9761 ( .A1(n9555), .A2(P1_IR_REG_29__SCAN_IN), .ZN(n7159) );
  NAND2_X1 U9762 ( .A1(n7813), .A2(n7810), .ZN(n13507) );
  NAND2_X1 U9763 ( .A1(n7315), .A2(n12088), .ZN(n7314) );
  INV_X1 U9764 ( .A(n12075), .ZN(n7763) );
  NAND2_X1 U9765 ( .A1(n7160), .A2(n12188), .ZN(P1_U3242) );
  OAI21_X1 U9766 ( .B1(n7309), .B2(n12185), .A(n11243), .ZN(n7160) );
  NAND2_X1 U9767 ( .A1(n7165), .A2(n7870), .ZN(n8587) );
  NAND3_X1 U9768 ( .A1(n7173), .A2(n8552), .A3(n8551), .ZN(n7165) );
  OAI21_X1 U9769 ( .B1(n9206), .B2(n9205), .A(n9141), .ZN(n9227) );
  AOI21_X1 U9770 ( .B1(n8697), .B2(n7886), .A(n7884), .ZN(n7883) );
  OAI21_X1 U9771 ( .B1(n9081), .B2(n9080), .A(n9079), .ZN(n9104) );
  BUF_X2 U9772 ( .A(n9241), .Z(n9199) );
  NAND3_X1 U9773 ( .A1(n9227), .A2(n9226), .A3(n7168), .ZN(n7167) );
  INV_X1 U9774 ( .A(n14023), .ZN(n7622) );
  NAND2_X1 U9775 ( .A1(n8870), .A2(n8869), .ZN(n8894) );
  NAND4_X1 U9776 ( .A1(n12670), .A2(n7442), .A3(P2_ADDR_REG_19__SCAN_IN), .A4(
        P1_ADDR_REG_19__SCAN_IN), .ZN(n7441) );
  NAND2_X1 U9777 ( .A1(n8868), .A2(n8867), .ZN(n8870) );
  NAND2_X1 U9778 ( .A1(n8631), .A2(n8630), .ZN(n7180) );
  NAND2_X1 U9779 ( .A1(n8617), .A2(n8616), .ZN(n7181) );
  NAND2_X1 U9780 ( .A1(n10789), .A2(n7187), .ZN(n7185) );
  NAND2_X1 U9781 ( .A1(n7185), .A2(n7186), .ZN(n11227) );
  NAND2_X1 U9782 ( .A1(n13717), .A2(n7196), .ZN(n7195) );
  NAND3_X1 U9783 ( .A1(n7191), .A2(n7195), .A3(n7192), .ZN(n7190) );
  NAND3_X1 U9784 ( .A1(n7195), .A2(n7194), .A3(n7191), .ZN(n13903) );
  NAND2_X1 U9785 ( .A1(n13860), .A2(n7208), .ZN(n7204) );
  NAND2_X1 U9786 ( .A1(n7204), .A2(n7205), .ZN(n13651) );
  NAND2_X1 U9787 ( .A1(n7637), .A2(n7217), .ZN(n7214) );
  NAND2_X1 U9788 ( .A1(n7214), .A2(n7215), .ZN(n13645) );
  MUX2_X1 U9789 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .S(n8534), .Z(n8578) );
  NAND2_X1 U9790 ( .A1(n10241), .A2(n10240), .ZN(n7234) );
  AOI21_X2 U9791 ( .B1(n10898), .B2(n10890), .A(n10797), .ZN(n10991) );
  AOI21_X2 U9792 ( .B1(n13716), .B2(n7236), .A(n13715), .ZN(n13907) );
  NAND2_X2 U9793 ( .A1(n13691), .A2(n13690), .ZN(n13729) );
  NAND2_X1 U9794 ( .A1(n13861), .A2(n7240), .ZN(n7237) );
  NAND2_X1 U9795 ( .A1(n7237), .A2(n7238), .ZN(n7437) );
  INV_X1 U9796 ( .A(n10556), .ZN(n13094) );
  NAND2_X1 U9797 ( .A1(n7703), .A2(n7247), .ZN(n7246) );
  MUX2_X1 U9798 ( .A(P3_REG1_REG_0__SCAN_IN), .B(P3_REG2_REG_0__SCAN_IN), .S(
        n10016), .Z(n10518) );
  NAND2_X1 U9799 ( .A1(n14942), .A2(n14901), .ZN(n14903) );
  NOR2_X2 U9800 ( .A1(n14950), .A2(n14951), .ZN(n14949) );
  INV_X1 U9801 ( .A(n14901), .ZN(n7261) );
  OAI211_X1 U9802 ( .C1(n12353), .C2(n7280), .A(n7278), .B(n7275), .ZN(n12277)
         );
  NAND2_X1 U9803 ( .A1(n12353), .A2(n7276), .ZN(n7275) );
  NOR2_X1 U9804 ( .A1(n12271), .A2(n7277), .ZN(n7276) );
  OAI21_X1 U9805 ( .B1(n12271), .B2(n7281), .A(n7279), .ZN(n7278) );
  OAI21_X1 U9806 ( .B1(n12271), .B2(n12238), .A(n7281), .ZN(n7279) );
  NAND2_X1 U9807 ( .A1(n12238), .A2(n12271), .ZN(n7280) );
  NAND2_X1 U9808 ( .A1(n7292), .A2(n7293), .ZN(n7926) );
  AND2_X1 U9809 ( .A1(n7293), .A2(n8138), .ZN(n8266) );
  NAND2_X1 U9810 ( .A1(n12054), .A2(n6722), .ZN(n7298) );
  NAND3_X1 U9811 ( .A1(n6708), .A2(n12064), .A3(n12063), .ZN(n7297) );
  AND2_X1 U9812 ( .A1(n7299), .A2(n7298), .ZN(n12070) );
  NAND2_X1 U9813 ( .A1(n11993), .A2(n6682), .ZN(n7305) );
  NAND2_X1 U9814 ( .A1(n7310), .A2(n12184), .ZN(n7309) );
  NAND2_X1 U9815 ( .A1(n12135), .A2(n6769), .ZN(n7310) );
  NAND2_X1 U9816 ( .A1(n7311), .A2(n7312), .ZN(n12042) );
  NAND4_X1 U9817 ( .A1(n12020), .A2(n12019), .A3(n7770), .A4(n12034), .ZN(
        n7311) );
  INV_X1 U9818 ( .A(n12086), .ZN(n7315) );
  NAND2_X1 U9819 ( .A1(n7317), .A2(n12085), .ZN(n7316) );
  NAND2_X1 U9820 ( .A1(n12086), .A2(n12087), .ZN(n7317) );
  OAI22_X1 U9821 ( .A1(n12011), .A2(n7319), .B1(n12010), .B2(n7318), .ZN(
        n12014) );
  NAND2_X1 U9822 ( .A1(n12014), .A2(n12015), .ZN(n12013) );
  NAND2_X1 U9823 ( .A1(n12657), .A2(n7333), .ZN(n7331) );
  NOR2_X1 U9824 ( .A1(n15616), .A2(n11420), .ZN(n15615) );
  INV_X1 U9825 ( .A(n15633), .ZN(n7333) );
  NAND2_X1 U9826 ( .A1(n9175), .A2(n7335), .ZN(n10235) );
  NAND3_X1 U9827 ( .A1(n9241), .A2(n7335), .A3(n10295), .ZN(n8529) );
  AOI22_X1 U9828 ( .A1(n10295), .A2(n9241), .B1(n7335), .B2(n9673), .ZN(n8531)
         );
  INV_X1 U9829 ( .A(n13532), .ZN(n7342) );
  INV_X1 U9830 ( .A(n13065), .ZN(n7348) );
  NAND2_X1 U9831 ( .A1(n11190), .A2(n7354), .ZN(n7353) );
  AOI21_X1 U9832 ( .B1(n7357), .B2(n10818), .A(n6689), .ZN(n7356) );
  NAND4_X1 U9833 ( .A1(n7361), .A2(n8683), .A3(n8495), .A4(n7360), .ZN(n9271)
         );
  OAI211_X1 U9834 ( .C1(n10644), .C2(n7364), .A(n7363), .B(n10856), .ZN(n8075)
         );
  NAND2_X1 U9835 ( .A1(n12417), .A2(n12455), .ZN(n7363) );
  INV_X1 U9836 ( .A(n12455), .ZN(n7364) );
  NAND2_X1 U9837 ( .A1(n10642), .A2(n12455), .ZN(n10850) );
  NAND2_X1 U9838 ( .A1(n10644), .A2(n10643), .ZN(n10642) );
  NAND2_X1 U9839 ( .A1(n12779), .A2(n7367), .ZN(n7366) );
  NAND2_X1 U9840 ( .A1(n7372), .A2(n7370), .ZN(n11150) );
  NAND2_X1 U9841 ( .A1(n10724), .A2(n7373), .ZN(n7372) );
  AOI21_X1 U9842 ( .B1(n8116), .B2(n6766), .A(n7378), .ZN(n7377) );
  INV_X1 U9843 ( .A(n7377), .ZN(n11342) );
  NAND2_X1 U9844 ( .A1(n7379), .A2(n12491), .ZN(n7378) );
  NAND3_X1 U9845 ( .A1(n7381), .A2(n7384), .A3(n7380), .ZN(n7379) );
  NAND2_X1 U9846 ( .A1(n12809), .A2(n7389), .ZN(n7385) );
  NAND2_X1 U9847 ( .A1(n7385), .A2(n7386), .ZN(n12780) );
  NAND4_X1 U9848 ( .A1(n8109), .A2(n7918), .A3(n8096), .A4(n7916), .ZN(n7396)
         );
  INV_X1 U9849 ( .A(n12694), .ZN(n10016) );
  NAND2_X4 U9850 ( .A1(n8427), .A2(n12694), .ZN(n10021) );
  AOI21_X1 U9851 ( .B1(n12847), .B2(n7400), .A(n7397), .ZN(n12826) );
  NAND2_X1 U9852 ( .A1(n11853), .A2(n7405), .ZN(n7404) );
  OAI21_X1 U9853 ( .B1(n12895), .B2(n7409), .A(n7406), .ZN(n12875) );
  OAI21_X1 U9854 ( .B1(n12895), .B2(n8219), .A(n12520), .ZN(n12885) );
  NAND2_X1 U9855 ( .A1(n8219), .A2(n12520), .ZN(n7411) );
  NAND2_X1 U9856 ( .A1(n8577), .A2(n8579), .ZN(n7416) );
  NAND3_X1 U9857 ( .A1(n7418), .A2(n8579), .A3(n6695), .ZN(n7415) );
  NAND2_X1 U9858 ( .A1(n8560), .A2(n8559), .ZN(n7418) );
  NAND3_X1 U9859 ( .A1(n7424), .A2(n7421), .A3(n7419), .ZN(n13698) );
  NAND3_X1 U9860 ( .A1(n13704), .A2(n7649), .A3(n13703), .ZN(n7433) );
  NOR2_X2 U9861 ( .A1(n13705), .A2(n13635), .ZN(n13636) );
  NOR2_X2 U9862 ( .A1(n10575), .A2(n15513), .ZN(n10574) );
  NAND2_X1 U9863 ( .A1(n14455), .A2(n7454), .ZN(n7453) );
  OAI211_X1 U9864 ( .C1(n14455), .C2(n7457), .A(n7455), .B(n7453), .ZN(n14694)
         );
  OR2_X1 U9865 ( .A1(n15389), .A2(n7462), .ZN(n7461) );
  INV_X1 U9866 ( .A(n14623), .ZN(n7465) );
  NAND2_X1 U9867 ( .A1(n11461), .A2(n7472), .ZN(n7470) );
  NAND2_X1 U9868 ( .A1(n7470), .A2(n7471), .ZN(n14633) );
  NAND2_X1 U9869 ( .A1(n14519), .A2(n7488), .ZN(n7487) );
  NAND3_X2 U9870 ( .A1(n9621), .A2(n7498), .A3(n7497), .ZN(n14230) );
  NAND2_X1 U9871 ( .A1(n6690), .A2(n14801), .ZN(n7497) );
  NAND3_X1 U9872 ( .A1(n14801), .A2(P1_REG1_REG_0__SCAN_IN), .A3(n9620), .ZN(
        n7499) );
  NAND3_X1 U9873 ( .A1(n9619), .A2(n14804), .A3(P1_REG2_REG_0__SCAN_IN), .ZN(
        n7500) );
  AND2_X1 U9874 ( .A1(n9305), .A2(n7502), .ZN(n7504) );
  NAND3_X1 U9875 ( .A1(n7504), .A2(n10230), .A3(n7779), .ZN(n9319) );
  NAND4_X1 U9876 ( .A1(n7504), .A2(n10230), .A3(n7779), .A4(n6749), .ZN(n9458)
         );
  AND4_X2 U9877 ( .A1(n6727), .A2(n7505), .A3(n9300), .A4(n9301), .ZN(n10230)
         );
  OAI21_X2 U9878 ( .B1(n9319), .B2(n7680), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n7508) );
  NOR2_X2 U9879 ( .A1(n10590), .A2(n15337), .ZN(n10743) );
  NAND2_X1 U9880 ( .A1(n7509), .A2(n15296), .ZN(n10590) );
  INV_X1 U9881 ( .A(n10592), .ZN(n7509) );
  NOR2_X2 U9882 ( .A1(n10193), .A2(n14064), .ZN(n10192) );
  NOR2_X2 U9883 ( .A1(n15186), .A2(n15183), .ZN(n15187) );
  AND2_X2 U9884 ( .A1(n14670), .A2(n7513), .ZN(n14609) );
  AOI21_X1 U9885 ( .B1(n10479), .B2(n10471), .A(n7550), .ZN(n10477) );
  NAND2_X1 U9886 ( .A1(n10972), .A2(n10971), .ZN(n10973) );
  INV_X1 U9887 ( .A(n12604), .ZN(n7571) );
  NAND2_X1 U9888 ( .A1(n7569), .A2(n10462), .ZN(n7568) );
  NAND2_X1 U9889 ( .A1(n12440), .A2(n12706), .ZN(n7569) );
  NAND2_X1 U9890 ( .A1(n9497), .A2(n8452), .ZN(n7572) );
  INV_X1 U9891 ( .A(n12222), .ZN(n7577) );
  NAND2_X1 U9892 ( .A1(n7859), .A2(n7581), .ZN(n8436) );
  AND2_X1 U9893 ( .A1(n8138), .A2(n8466), .ZN(n7583) );
  NAND2_X1 U9894 ( .A1(n10467), .A2(n10466), .ZN(n10480) );
  NAND2_X1 U9895 ( .A1(n7950), .A2(n7949), .ZN(n8125) );
  NAND2_X1 U9896 ( .A1(n7585), .A2(n7586), .ZN(n11836) );
  NAND2_X1 U9897 ( .A1(n14193), .A2(n6676), .ZN(n7585) );
  NAND2_X1 U9898 ( .A1(n14193), .A2(n14194), .ZN(n14192) );
  INV_X1 U9899 ( .A(n9307), .ZN(n9337) );
  NAND2_X1 U9900 ( .A1(n10008), .A2(n10007), .ZN(n10009) );
  NAND2_X1 U9901 ( .A1(n10009), .A2(n10010), .ZN(n10678) );
  OR2_X1 U9902 ( .A1(n9612), .A2(P1_IR_REG_19__SCAN_IN), .ZN(n9608) );
  NAND2_X1 U9903 ( .A1(n7619), .A2(n7618), .ZN(n14172) );
  OAI21_X1 U9904 ( .B1(n10239), .B2(n7636), .A(n10544), .ZN(n7632) );
  NAND2_X1 U9905 ( .A1(n7633), .A2(n7631), .ZN(n10548) );
  NAND4_X1 U9906 ( .A1(n8496), .A2(n8497), .A3(n8498), .A4(n8517), .ZN(n8499)
         );
  OAI21_X1 U9907 ( .B1(n13805), .B2(n7642), .A(n7640), .ZN(n13782) );
  OAI21_X1 U9908 ( .B1(n13805), .B2(n13654), .A(n13655), .ZN(n13801) );
  INV_X1 U9909 ( .A(n13800), .ZN(n7644) );
  NAND2_X1 U9910 ( .A1(n10786), .A2(n7647), .ZN(n7646) );
  NAND3_X2 U9911 ( .A1(n9634), .A2(n7650), .A3(n9635), .ZN(n14229) );
  INV_X1 U9912 ( .A(n7651), .ZN(n7650) );
  OAI21_X1 U9913 ( .B1(n9619), .B2(n7653), .A(n7652), .ZN(n7651) );
  NAND3_X1 U9914 ( .A1(n14804), .A2(n9619), .A3(P1_REG2_REG_1__SCAN_IN), .ZN(
        n7652) );
  NAND2_X1 U9915 ( .A1(n10184), .A2(n11976), .ZN(n7656) );
  NAND2_X1 U9916 ( .A1(n14656), .A2(n14422), .ZN(n7660) );
  NAND2_X1 U9917 ( .A1(n7660), .A2(n7661), .ZN(n14425) );
  NAND2_X1 U9918 ( .A1(n14578), .A2(n14437), .ZN(n7665) );
  NAND2_X1 U9919 ( .A1(n7665), .A2(n7666), .ZN(n14439) );
  NAND2_X1 U9920 ( .A1(n10584), .A2(n7672), .ZN(n7669) );
  NAND2_X1 U9921 ( .A1(n7669), .A2(n7670), .ZN(n10827) );
  AOI21_X2 U9922 ( .B1(n6762), .B2(n10758), .A(n6656), .ZN(n7672) );
  NOR2_X1 U9923 ( .A1(n9319), .A2(P1_IR_REG_24__SCAN_IN), .ZN(n9317) );
  XNOR2_X2 U9924 ( .A(n7692), .B(n8032), .ZN(n10365) );
  NAND3_X1 U9925 ( .A1(n7707), .A2(n6812), .A3(n7706), .ZN(n9086) );
  NAND3_X1 U9926 ( .A1(n7707), .A2(n7708), .A3(n7706), .ZN(n9082) );
  NAND3_X1 U9927 ( .A1(n7723), .A2(n6728), .A3(n7726), .ZN(n7721) );
  NAND2_X1 U9928 ( .A1(n13704), .A2(n13703), .ZN(n13900) );
  NOR2_X1 U9929 ( .A1(n8499), .A2(P2_IR_REG_26__SCAN_IN), .ZN(n7755) );
  NAND2_X1 U9930 ( .A1(n7765), .A2(n7766), .ZN(n12011) );
  NAND3_X1 U9931 ( .A1(n12006), .A2(n6778), .A3(n12005), .ZN(n7765) );
  NAND2_X1 U9932 ( .A1(n7768), .A2(n7769), .ZN(n11993) );
  NAND3_X1 U9933 ( .A1(n11987), .A2(n6777), .A3(n11986), .ZN(n7768) );
  INV_X1 U9934 ( .A(n9554), .ZN(n7774) );
  NAND2_X1 U9935 ( .A1(n7774), .A2(n6669), .ZN(n7776) );
  NAND2_X2 U9936 ( .A1(n14807), .A2(n6668), .ZN(n9817) );
  INV_X2 U9937 ( .A(n9339), .ZN(n7779) );
  NAND2_X1 U9938 ( .A1(n12102), .A2(n7784), .ZN(n7783) );
  INV_X1 U9939 ( .A(n12100), .ZN(n7784) );
  NAND2_X2 U9940 ( .A1(n13063), .A2(n7807), .ZN(n13065) );
  NAND2_X1 U9941 ( .A1(n11878), .A2(n13503), .ZN(n7813) );
  NAND2_X1 U9942 ( .A1(n9695), .A2(n7817), .ZN(n7816) );
  INV_X1 U9943 ( .A(n9934), .ZN(n7815) );
  OR2_X1 U9944 ( .A1(n9697), .A2(n7815), .ZN(n7814) );
  NAND2_X1 U9945 ( .A1(n9943), .A2(n10159), .ZN(n7820) );
  NAND2_X1 U9946 ( .A1(n7820), .A2(n7818), .ZN(n10376) );
  AOI21_X1 U9947 ( .B1(n9944), .B2(n10159), .A(n7819), .ZN(n7818) );
  OAI211_X1 U9948 ( .C1(n13102), .C2(n7825), .A(n7821), .B(n7823), .ZN(
        P2_U3192) );
  NAND2_X1 U9949 ( .A1(n13102), .A2(n7822), .ZN(n7821) );
  NAND4_X1 U9950 ( .A1(n10519), .A2(n7918), .A3(n7917), .A4(n8040), .ZN(n8069)
         );
  NAND2_X1 U9951 ( .A1(n7846), .A2(n15746), .ZN(n7850) );
  NAND2_X1 U9952 ( .A1(n7849), .A2(n7848), .ZN(n8489) );
  NAND3_X1 U9953 ( .A1(n8492), .A2(n8491), .A3(n8683), .ZN(n8775) );
  OAI21_X1 U9954 ( .B1(n9058), .B2(n7877), .A(n7874), .ZN(n9081) );
  NAND2_X1 U9955 ( .A1(n7873), .A2(n7871), .ZN(n9078) );
  NAND2_X1 U9956 ( .A1(n7877), .A2(n7874), .ZN(n7872) );
  NAND2_X1 U9957 ( .A1(n7893), .A2(n7892), .ZN(n7890) );
  NAND2_X1 U9958 ( .A1(n8763), .A2(n8764), .ZN(n8762) );
  INV_X1 U9959 ( .A(n12727), .ZN(n11854) );
  AND2_X1 U9960 ( .A1(n12739), .A2(n12738), .ZN(n12931) );
  XNOR2_X1 U9961 ( .A(n9147), .B(n9126), .ZN(n11804) );
  NAND2_X1 U9962 ( .A1(n9462), .A2(n9311), .ZN(n9465) );
  NAND2_X1 U9963 ( .A1(n8995), .A2(n8994), .ZN(n8998) );
  INV_X2 U9964 ( .A(n9158), .ZN(n9816) );
  INV_X1 U9965 ( .A(n14596), .ZN(n14435) );
  XNOR2_X1 U9966 ( .A(n14868), .B(P1_ADDR_REG_5__SCAN_IN), .ZN(n14886) );
  AND2_X1 U9967 ( .A1(n14867), .A2(n14868), .ZN(n14828) );
  NAND2_X1 U9968 ( .A1(n10298), .A2(n9785), .ZN(n9902) );
  INV_X1 U9969 ( .A(n12381), .ZN(n8349) );
  NAND2_X1 U9970 ( .A1(n8489), .A2(n15788), .ZN(n8477) );
  OR2_X1 U9971 ( .A1(P3_REG3_REG_16__SCAN_IN), .A2(n8243), .ZN(n7910) );
  AND4_X1 U9972 ( .A1(n9275), .A2(n9175), .A3(n11245), .A4(n10983), .ZN(n7911)
         );
  INV_X1 U9973 ( .A(n12546), .ZN(n8291) );
  NOR2_X1 U9974 ( .A1(n10748), .A2(n10832), .ZN(n7912) );
  INV_X1 U9975 ( .A(n12578), .ZN(n8422) );
  AND2_X1 U9976 ( .A1(n8797), .A2(n8774), .ZN(n7913) );
  INV_X1 U9977 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n8500) );
  XOR2_X1 U9978 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(P1_ADDR_REG_19__SCAN_IN), 
        .Z(n7914) );
  INV_X1 U9979 ( .A(n15378), .ZN(n15212) );
  INV_X1 U9980 ( .A(n12147), .ZN(n11480) );
  AND2_X1 U9981 ( .A1(n8565), .A2(n9795), .ZN(n8528) );
  NAND2_X1 U9982 ( .A1(n12013), .A2(n12012), .ZN(n12020) );
  AND2_X1 U9983 ( .A1(n12147), .A2(n12023), .ZN(n12024) );
  AND2_X1 U9984 ( .A1(n12033), .A2(n12032), .ZN(n12034) );
  NAND2_X1 U9985 ( .A1(n12082), .A2(n12081), .ZN(n12083) );
  INV_X1 U9986 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n7995) );
  CLKBUF_X3 U9987 ( .A(n8565), .Z(n9222) );
  INV_X1 U9988 ( .A(n12412), .ZN(n8398) );
  OR2_X1 U9989 ( .A1(n14743), .A2(n14401), .ZN(n14402) );
  INV_X1 U9990 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n9310) );
  NAND2_X1 U9991 ( .A1(n15704), .A2(n12438), .ZN(n10321) );
  INV_X1 U9992 ( .A(n9024), .ZN(n9022) );
  INV_X1 U9993 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n8857) );
  INV_X1 U9994 ( .A(n15554), .ZN(n9674) );
  INV_X1 U9995 ( .A(n11276), .ZN(n11272) );
  INV_X1 U9996 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n13404) );
  NAND2_X1 U9997 ( .A1(n10137), .A2(n11970), .ZN(n10453) );
  INV_X1 U9998 ( .A(SI_11_), .ZN(n8745) );
  INV_X1 U9999 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n9306) );
  INV_X1 U10000 ( .A(P3_REG3_REG_14__SCAN_IN), .ZN(n8212) );
  NOR2_X1 U10001 ( .A1(P3_REG3_REG_22__SCAN_IN), .A2(n8318), .ZN(n8338) );
  INV_X1 U10002 ( .A(n14928), .ZN(n15605) );
  NOR2_X1 U10003 ( .A1(P3_REG3_REG_17__SCAN_IN), .A2(n7910), .ZN(n8271) );
  INV_X1 U10004 ( .A(n12414), .ZN(n8172) );
  OR2_X1 U10005 ( .A1(n12611), .A2(n12585), .ZN(n9867) );
  INV_X1 U10006 ( .A(n9647), .ZN(n9644) );
  INV_X1 U10007 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n13119) );
  AND2_X1 U10008 ( .A1(n11907), .A2(n11906), .ZN(n11908) );
  AND2_X1 U10009 ( .A1(n8882), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8883) );
  OR2_X1 U10010 ( .A1(n9112), .A2(n9111), .ZN(n9131) );
  NAND2_X1 U10011 ( .A1(n9022), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n9046) );
  OR2_X1 U10012 ( .A1(n8709), .A2(n8706), .ZN(n8730) );
  AND2_X1 U10013 ( .A1(n9642), .A2(n9176), .ZN(n9672) );
  INV_X1 U10014 ( .A(n13630), .ZN(n13555) );
  INV_X1 U10015 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n8501) );
  OR2_X1 U10016 ( .A1(n9271), .A2(n9270), .ZN(n9273) );
  AND2_X1 U10017 ( .A1(n11624), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n11640) );
  NOR2_X1 U10018 ( .A1(n11464), .A2(n13404), .ZN(n11624) );
  INV_X1 U10019 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n11291) );
  INV_X2 U10020 ( .A(n10435), .ZN(n12110) );
  AND2_X1 U10021 ( .A1(n9468), .A2(n9763), .ZN(n12134) );
  AND2_X1 U10022 ( .A1(n14895), .A2(P1_ADDR_REG_7__SCAN_IN), .ZN(n14832) );
  INV_X1 U10023 ( .A(P3_ADDR_REG_12__SCAN_IN), .ZN(n14844) );
  INV_X1 U10024 ( .A(P3_REG3_REG_10__SCAN_IN), .ZN(n8144) );
  AND2_X1 U10025 ( .A1(n8285), .A2(n12264), .ZN(n8295) );
  AND2_X1 U10026 ( .A1(n12233), .A2(n12232), .ZN(n12299) );
  AND2_X1 U10027 ( .A1(n8271), .A2(n8270), .ZN(n8285) );
  NAND2_X1 U10028 ( .A1(n12606), .A2(n15712), .ZN(n12607) );
  AND4_X1 U10029 ( .A1(n8344), .A2(n8343), .A3(n8342), .A4(n8341), .ZN(n12224)
         );
  AND2_X1 U10030 ( .A1(n12532), .A2(n12530), .ZN(n12874) );
  AND2_X1 U10031 ( .A1(n10462), .A2(n12706), .ZN(n15712) );
  INV_X1 U10032 ( .A(n13050), .ZN(n8479) );
  INV_X1 U10033 ( .A(P3_REG0_REG_29__SCAN_IN), .ZN(n8486) );
  OR2_X1 U10034 ( .A1(n8066), .A2(n11391), .ZN(n8347) );
  AND2_X1 U10035 ( .A1(n7935), .A2(n8470), .ZN(n15766) );
  NAND2_X1 U10036 ( .A1(n10765), .A2(n12440), .ZN(n15744) );
  NAND2_X1 U10037 ( .A1(n8433), .A2(n12593), .ZN(n15017) );
  INV_X1 U10038 ( .A(SI_13_), .ZN(n14929) );
  NAND2_X1 U10039 ( .A1(n13067), .A2(n13069), .ZN(n13070) );
  NAND2_X1 U10040 ( .A1(n8883), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n8937) );
  INV_X1 U10041 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n13537) );
  INV_X1 U10042 ( .A(n9782), .ZN(n9678) );
  INV_X1 U10043 ( .A(n13643), .ZN(n13667) );
  INV_X1 U10044 ( .A(n9294), .ZN(n9295) );
  AND2_X1 U10045 ( .A1(n9131), .A2(n9113), .ZN(n13745) );
  INV_X1 U10046 ( .A(n13694), .ZN(n13665) );
  OR2_X1 U10047 ( .A1(n13845), .A2(n13676), .ZN(n13677) );
  NOR2_X1 U10048 ( .A1(n9173), .A2(n9675), .ZN(n9897) );
  AND2_X1 U10049 ( .A1(n9642), .A2(n9175), .ZN(n9787) );
  NOR2_X1 U10050 ( .A1(n9273), .A2(P2_IR_REG_23__SCAN_IN), .ZN(n9277) );
  INV_X1 U10051 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n8851) );
  OR2_X1 U10052 ( .A1(n11663), .A2(n11662), .ZN(n11678) );
  AND2_X1 U10053 ( .A1(n11786), .A2(n11785), .ZN(n14100) );
  INV_X1 U10054 ( .A(n11735), .ZN(n11734) );
  INV_X1 U10055 ( .A(n14115), .ZN(n14200) );
  INV_X1 U10056 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n14867) );
  INV_X1 U10057 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n14862) );
  OR2_X1 U10058 ( .A1(n9853), .A2(n9852), .ZN(n10056) );
  INV_X1 U10059 ( .A(n12151), .ZN(n10586) );
  XNOR2_X1 U10060 ( .A(n14705), .B(n14447), .ZN(n14484) );
  INV_X1 U10061 ( .A(n11099), .ZN(n12158) );
  OR2_X1 U10062 ( .A1(n9977), .A2(n14612), .ZN(n15318) );
  OAI21_X1 U10063 ( .B1(n9755), .B2(P1_D_REG_1__SCAN_IN), .A(n9595), .ZN(n9760) );
  NAND2_X1 U10064 ( .A1(n9155), .A2(n9154), .ZN(n9167) );
  AND2_X1 U10065 ( .A1(n8874), .A2(n8873), .ZN(n8893) );
  NOR2_X1 U10066 ( .A1(n8188), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n8213) );
  AND2_X1 U10067 ( .A1(n10472), .A2(P3_STATE_REG_SCAN_IN), .ZN(n15002) );
  INV_X1 U10068 ( .A(n15585), .ZN(n15021) );
  AND4_X1 U10069 ( .A1(n12386), .A2(n12385), .A3(n12384), .A4(n12383), .ZN(
        n12713) );
  AND4_X1 U10070 ( .A1(n8355), .A2(n8354), .A3(n8353), .A4(n8352), .ZN(n12229)
         );
  AND4_X1 U10071 ( .A1(n8277), .A2(n8276), .A3(n8275), .A4(n8274), .ZN(n12857)
         );
  INV_X1 U10072 ( .A(n15661), .ZN(n15681) );
  AND2_X1 U10073 ( .A1(n15719), .A2(n15700), .ZN(n15716) );
  NOR2_X1 U10074 ( .A1(n15788), .A2(n13479), .ZN(n8474) );
  AND2_X1 U10075 ( .A1(n8469), .A2(n8468), .ZN(n10655) );
  INV_X1 U10076 ( .A(n15106), .ZN(n15746) );
  AND2_X1 U10077 ( .A1(n10019), .A2(P3_STATE_REG_SCAN_IN), .ZN(n9323) );
  INV_X1 U10078 ( .A(P3_IR_REG_21__SCAN_IN), .ZN(n7996) );
  INV_X1 U10079 ( .A(n10337), .ZN(n10333) );
  AND2_X1 U10080 ( .A1(n13708), .A2(n9213), .ZN(n13722) );
  AND2_X1 U10081 ( .A1(n9671), .A2(n9670), .ZN(n15125) );
  INV_X1 U10082 ( .A(n15131), .ZN(n13556) );
  INV_X1 U10083 ( .A(n13542), .ZN(n15128) );
  INV_X1 U10084 ( .A(n6662), .ZN(n9195) );
  INV_X1 U10085 ( .A(n8571), .ZN(n9217) );
  INV_X1 U10086 ( .A(n15442), .ZN(n15474) );
  INV_X1 U10087 ( .A(n15479), .ZN(n15453) );
  XNOR2_X1 U10088 ( .A(n13912), .B(n13665), .ZN(n13737) );
  INV_X1 U10089 ( .A(n13683), .ZN(n13806) );
  INV_X1 U10090 ( .A(n13890), .ZN(n15139) );
  INV_X1 U10091 ( .A(n13874), .ZN(n15148) );
  INV_X1 U10092 ( .A(n9790), .ZN(n10294) );
  NAND2_X1 U10093 ( .A1(n10073), .A2(n9667), .ZN(n15548) );
  INV_X1 U10094 ( .A(n13998), .ZN(n15527) );
  AND2_X1 U10095 ( .A1(n9783), .A2(n15490), .ZN(n9899) );
  AND2_X1 U10096 ( .A1(n9398), .A2(n9394), .ZN(n9945) );
  AND2_X1 U10097 ( .A1(n9280), .A2(n9285), .ZN(n9649) );
  AND2_X1 U10098 ( .A1(n8826), .A2(n8853), .ZN(n10865) );
  NAND2_X1 U10099 ( .A1(n9322), .A2(n9383), .ZN(n9630) );
  AND2_X1 U10100 ( .A1(n9996), .A2(n9629), .ZN(n15379) );
  AND4_X1 U10101 ( .A1(n11721), .A2(n11720), .A3(n11719), .A4(n11718), .ZN(
        n14543) );
  INV_X1 U10102 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n14891) );
  INV_X1 U10103 ( .A(n15267), .ZN(n14340) );
  AND2_X1 U10104 ( .A1(n9809), .A2(n6669), .ZN(n14378) );
  OR2_X1 U10105 ( .A1(n9975), .A2(n11243), .ZN(n9721) );
  NAND2_X1 U10106 ( .A1(n9973), .A2(n9972), .ZN(n14409) );
  NAND2_X1 U10107 ( .A1(n14584), .A2(n14595), .ZN(n14583) );
  INV_X1 U10108 ( .A(n15351), .ZN(n15375) );
  INV_X1 U10109 ( .A(n14550), .ZN(n15299) );
  NAND2_X1 U10110 ( .A1(n14409), .A2(n14986), .ZN(n14969) );
  INV_X1 U10111 ( .A(n9626), .ZN(n9772) );
  AND2_X1 U10112 ( .A1(n10693), .A2(P1_STATE_REG_SCAN_IN), .ZN(n12186) );
  INV_X1 U10113 ( .A(n15386), .ZN(n15219) );
  NAND2_X1 U10114 ( .A1(n15318), .A2(n15341), .ZN(n15386) );
  AND2_X1 U10115 ( .A1(n9974), .A2(n9760), .ZN(n9773) );
  XNOR2_X1 U10116 ( .A(n9309), .B(n9308), .ZN(n9631) );
  INV_X1 U10117 ( .A(n12131), .ZN(n9763) );
  XNOR2_X1 U10118 ( .A(n9812), .B(P1_IR_REG_14__SCAN_IN), .ZN(n11451) );
  INV_X1 U10119 ( .A(n14886), .ZN(n14887) );
  NAND2_X1 U10120 ( .A1(n8465), .A2(n8464), .ZN(n9868) );
  AND4_X1 U10121 ( .A1(n12275), .A2(n12274), .A3(n12273), .A4(n12272), .ZN(
        n12276) );
  OR2_X1 U10122 ( .A1(n9878), .A2(n9877), .ZN(n15009) );
  INV_X1 U10123 ( .A(n15002), .ZN(n15593) );
  AND2_X1 U10124 ( .A1(n9884), .A2(n15711), .ZN(n15581) );
  INV_X1 U10125 ( .A(n12229), .ZN(n12619) );
  INV_X1 U10126 ( .A(n12857), .ZN(n12625) );
  NAND2_X1 U10127 ( .A1(n15577), .A2(n8427), .ZN(n15661) );
  INV_X1 U10128 ( .A(n15674), .ZN(n15613) );
  INV_X1 U10129 ( .A(n15082), .ZN(n15687) );
  INV_X1 U10130 ( .A(n15097), .ZN(n12898) );
  NAND2_X1 U10131 ( .A1(n15719), .A2(n10723), .ZN(n12827) );
  NAND2_X1 U10132 ( .A1(n15788), .A2(n15770), .ZN(n12986) );
  INV_X1 U10133 ( .A(n15788), .ZN(n15786) );
  INV_X1 U10134 ( .A(n15773), .ZN(n15771) );
  INV_X1 U10135 ( .A(SI_17_), .ZN(n13439) );
  INV_X1 U10136 ( .A(SI_12_), .ZN(n9367) );
  NAND2_X1 U10137 ( .A1(n9616), .A2(P3_U3151), .ZN(n14936) );
  NAND2_X1 U10138 ( .A1(n9947), .A2(P2_STATE_REG_SCAN_IN), .ZN(n15131) );
  INV_X1 U10139 ( .A(n15125), .ZN(n13558) );
  AND2_X1 U10140 ( .A1(n9679), .A2(n13865), .ZN(n13542) );
  NAND2_X1 U10141 ( .A1(n9100), .A2(n9099), .ZN(n13688) );
  OR2_X1 U10142 ( .A1(n15420), .A2(P2_U3088), .ZN(n15479) );
  OR2_X1 U10143 ( .A1(n9408), .A2(n14029), .ZN(n15442) );
  OR2_X1 U10144 ( .A1(n15151), .A2(n15522), .ZN(n13859) );
  INV_X1 U10145 ( .A(n15573), .ZN(n15158) );
  NAND2_X1 U10146 ( .A1(n10071), .A2(n9899), .ZN(n15559) );
  NOR2_X1 U10147 ( .A1(n15488), .A2(n15480), .ZN(n15484) );
  INV_X1 U10148 ( .A(n15484), .ZN(n15485) );
  INV_X1 U10149 ( .A(n9176), .ZN(n10983) );
  INV_X1 U10150 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n9815) );
  INV_X1 U10151 ( .A(n15172), .ZN(n14191) );
  INV_X1 U10152 ( .A(n14543), .ZN(n14569) );
  OR2_X1 U10153 ( .A1(n9727), .A2(n9726), .ZN(n15266) );
  INV_X1 U10154 ( .A(n14378), .ZN(n15264) );
  NAND2_X1 U10155 ( .A1(n9721), .A2(n9719), .ZN(n15271) );
  NAND2_X1 U10156 ( .A1(n9976), .A2(n9975), .ZN(n14986) );
  OR2_X1 U10157 ( .A1(n6665), .A2(n15351), .ZN(n14599) );
  OR2_X1 U10158 ( .A1(n6665), .A2(n9977), .ZN(n14982) );
  AND4_X1 U10159 ( .A1(n14962), .A2(n14961), .A3(n14960), .A4(n14959), .ZN(
        n14965) );
  INV_X1 U10160 ( .A(n15389), .ZN(n15387) );
  AND2_X2 U10161 ( .A1(n9973), .A2(n9773), .ZN(n15389) );
  INV_X1 U10162 ( .A(n15314), .ZN(n15313) );
  AND2_X1 U10163 ( .A1(n9631), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9386) );
  INV_X1 U10164 ( .A(n9380), .ZN(n11509) );
  INV_X1 U10165 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n10770) );
  INV_X1 U10166 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n9813) );
  NOR2_X1 U10167 ( .A1(n9398), .A2(n9299), .ZN(P2_U3947) );
  AND2_X2 U10168 ( .A1(n9386), .A2(n9623), .ZN(P1_U4016) );
  NAND2_X1 U10169 ( .A1(n7926), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7922) );
  MUX2_X1 U10170 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7922), .S(
        P3_IR_REG_20__SCAN_IN), .Z(n7923) );
  INV_X1 U10171 ( .A(n8266), .ZN(n7924) );
  NAND2_X1 U10172 ( .A1(n7924), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7925) );
  MUX2_X1 U10173 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7925), .S(
        P3_IR_REG_19__SCAN_IN), .Z(n7927) );
  OAI21_X1 U10174 ( .B1(n10765), .B2(n8481), .A(n12706), .ZN(n7930) );
  NAND2_X1 U10175 ( .A1(n7930), .A2(n12440), .ZN(n7932) );
  OAI21_X1 U10176 ( .B1(n8481), .B2(n10656), .A(n10765), .ZN(n7931) );
  NAND2_X1 U10177 ( .A1(n7932), .A2(n7931), .ZN(n9872) );
  NAND2_X1 U10178 ( .A1(n10462), .A2(n12666), .ZN(n12602) );
  INV_X1 U10179 ( .A(n12602), .ZN(n12611) );
  AND2_X1 U10180 ( .A1(n15744), .A2(n12611), .ZN(n7933) );
  NAND2_X1 U10181 ( .A1(n9872), .A2(n7933), .ZN(n7935) );
  NOR2_X1 U10182 ( .A1(n10462), .A2(n12706), .ZN(n7934) );
  NAND2_X1 U10183 ( .A1(n12613), .A2(n7934), .ZN(n8470) );
  NAND2_X1 U10184 ( .A1(n10765), .A2(n15712), .ZN(n15765) );
  INV_X1 U10185 ( .A(n8029), .ZN(n7936) );
  XNOR2_X1 U10186 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .ZN(n8030) );
  NAND2_X1 U10187 ( .A1(n7936), .A2(n8030), .ZN(n7938) );
  INV_X1 U10188 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n9359) );
  NAND2_X1 U10189 ( .A1(n9359), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n7937) );
  NAND2_X1 U10190 ( .A1(n7938), .A2(n7937), .ZN(n8042) );
  XNOR2_X1 U10191 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .ZN(n8041) );
  NAND2_X1 U10192 ( .A1(n8042), .A2(n8041), .ZN(n7940) );
  INV_X1 U10193 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n9330) );
  NAND2_X1 U10194 ( .A1(n9330), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n7939) );
  NAND2_X1 U10195 ( .A1(n8053), .A2(n8052), .ZN(n7942) );
  NAND2_X1 U10196 ( .A1(n9331), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n7941) );
  NAND2_X1 U10197 ( .A1(n13274), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n7943) );
  NOR2_X1 U10198 ( .A1(n10427), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n7944) );
  NAND2_X1 U10199 ( .A1(n10427), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n7945) );
  NAND2_X1 U10200 ( .A1(n8095), .A2(n8094), .ZN(n7947) );
  NAND2_X1 U10201 ( .A1(n9373), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n7946) );
  XNOR2_X1 U10202 ( .A(n9376), .B(P1_DATAO_REG_7__SCAN_IN), .ZN(n8111) );
  INV_X1 U10203 ( .A(n8111), .ZN(n7948) );
  NAND2_X1 U10204 ( .A1(n8112), .A2(n7948), .ZN(n7950) );
  NAND2_X1 U10205 ( .A1(n9376), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n7949) );
  NAND2_X1 U10206 ( .A1(n9391), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n7951) );
  XNOR2_X1 U10207 ( .A(n7953), .B(P1_DATAO_REG_9__SCAN_IN), .ZN(n8134) );
  INV_X1 U10208 ( .A(n8134), .ZN(n7952) );
  NAND2_X1 U10209 ( .A1(n8135), .A2(n7952), .ZN(n7955) );
  NAND2_X1 U10210 ( .A1(n7953), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n7954) );
  XNOR2_X1 U10211 ( .A(n7957), .B(P1_DATAO_REG_10__SCAN_IN), .ZN(n8152) );
  INV_X1 U10212 ( .A(n8152), .ZN(n7956) );
  NAND2_X1 U10213 ( .A1(n9691), .A2(P1_DATAO_REG_12__SCAN_IN), .ZN(n7959) );
  NAND2_X1 U10214 ( .A1(n9594), .A2(P2_DATAO_REG_12__SCAN_IN), .ZN(n7958) );
  NAND2_X1 U10215 ( .A1(n7959), .A2(n7958), .ZN(n8179) );
  XNOR2_X1 U10216 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .ZN(n8206) );
  INV_X1 U10217 ( .A(n8206), .ZN(n7961) );
  NAND2_X1 U10218 ( .A1(n9815), .A2(P2_DATAO_REG_14__SCAN_IN), .ZN(n7962) );
  NAND2_X1 U10219 ( .A1(n10054), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n7964) );
  NAND2_X1 U10220 ( .A1(n9971), .A2(P2_DATAO_REG_15__SCAN_IN), .ZN(n7963) );
  NAND2_X1 U10221 ( .A1(n7964), .A2(n7963), .ZN(n8220) );
  NAND2_X1 U10222 ( .A1(n10234), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n7968) );
  NAND2_X1 U10223 ( .A1(n10153), .A2(P2_DATAO_REG_16__SCAN_IN), .ZN(n7965) );
  NAND2_X1 U10224 ( .A1(n7968), .A2(n7965), .ZN(n8235) );
  INV_X1 U10225 ( .A(n8235), .ZN(n7966) );
  XNOR2_X1 U10226 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(P2_DATAO_REG_17__SCAN_IN), 
        .ZN(n8250) );
  INV_X1 U10227 ( .A(n8250), .ZN(n7969) );
  NAND2_X1 U10228 ( .A1(n10721), .A2(P1_DATAO_REG_18__SCAN_IN), .ZN(n7972) );
  NAND2_X1 U10229 ( .A1(n10735), .A2(P2_DATAO_REG_18__SCAN_IN), .ZN(n7970) );
  INV_X1 U10230 ( .A(n8261), .ZN(n7971) );
  NAND2_X1 U10231 ( .A1(n10770), .A2(P1_DATAO_REG_19__SCAN_IN), .ZN(n7974) );
  NAND2_X1 U10232 ( .A1(n13423), .A2(P2_DATAO_REG_19__SCAN_IN), .ZN(n7973) );
  NAND2_X1 U10233 ( .A1(n7974), .A2(n7973), .ZN(n8279) );
  INV_X1 U10234 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n10982) );
  NAND2_X1 U10235 ( .A1(n10982), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n7979) );
  INV_X1 U10236 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n10985) );
  NAND2_X1 U10237 ( .A1(n10985), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n7978) );
  NAND2_X1 U10238 ( .A1(n7979), .A2(n7978), .ZN(n8301) );
  INV_X1 U10239 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n11864) );
  XNOR2_X1 U10240 ( .A(n11864), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n8314) );
  NAND2_X1 U10241 ( .A1(n11864), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n7980) );
  XNOR2_X1 U10242 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(P2_DATAO_REG_23__SCAN_IN), 
        .ZN(n8325) );
  INV_X1 U10243 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n7981) );
  NAND2_X1 U10244 ( .A1(n7982), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n7983) );
  INV_X1 U10245 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n14037) );
  NAND2_X1 U10246 ( .A1(n14037), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n7984) );
  INV_X1 U10247 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n14816) );
  NAND2_X1 U10248 ( .A1(n14816), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n7985) );
  INV_X1 U10249 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n14034) );
  NOR2_X1 U10250 ( .A1(n14034), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n7987) );
  NAND2_X1 U10251 ( .A1(n14034), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n7988) );
  INV_X1 U10252 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n11560) );
  NOR2_X1 U10253 ( .A1(n11560), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n7989) );
  INV_X1 U10254 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n14028) );
  INV_X1 U10255 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n13246) );
  XNOR2_X1 U10256 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .ZN(n7991) );
  NAND2_X1 U10257 ( .A1(n7990), .A2(n7991), .ZN(n11920) );
  INV_X1 U10258 ( .A(n7990), .ZN(n7993) );
  INV_X1 U10259 ( .A(n7991), .ZN(n7992) );
  NAND2_X1 U10260 ( .A1(n7993), .A2(n7992), .ZN(n7994) );
  NOR2_X1 U10261 ( .A1(P3_IR_REG_22__SCAN_IN), .A2(P3_IR_REG_18__SCAN_IN), 
        .ZN(n7997) );
  NAND4_X1 U10262 ( .A1(n7997), .A2(n7996), .A3(n7995), .A4(n13367), .ZN(n7998) );
  INV_X1 U10263 ( .A(SI_29_), .ZN(n13329) );
  OR2_X1 U10264 ( .A1(n8066), .A2(n13329), .ZN(n8004) );
  INV_X1 U10265 ( .A(P3_REG3_REG_28__SCAN_IN), .ZN(n8012) );
  NOR2_X1 U10266 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n8077) );
  NAND2_X1 U10267 ( .A1(n8077), .A2(n8076), .ZN(n8088) );
  NOR2_X1 U10268 ( .A1(P3_REG3_REG_9__SCAN_IN), .A2(P3_REG3_REG_8__SCAN_IN), 
        .ZN(n8010) );
  NAND2_X1 U10269 ( .A1(n8145), .A2(n8144), .ZN(n8159) );
  NAND2_X1 U10270 ( .A1(n8213), .A2(n8212), .ZN(n8229) );
  INV_X1 U10271 ( .A(P3_REG3_REG_18__SCAN_IN), .ZN(n8270) );
  INV_X1 U10272 ( .A(P3_REG3_REG_19__SCAN_IN), .ZN(n12264) );
  INV_X1 U10273 ( .A(P3_REG3_REG_20__SCAN_IN), .ZN(n12328) );
  NOR2_X1 U10274 ( .A1(P3_REG3_REG_24__SCAN_IN), .A2(P3_REG3_REG_23__SCAN_IN), 
        .ZN(n8011) );
  NAND2_X1 U10275 ( .A1(n8338), .A2(n8011), .ZN(n8350) );
  INV_X1 U10276 ( .A(P3_REG3_REG_27__SCAN_IN), .ZN(n12240) );
  NAND2_X1 U10277 ( .A1(n8372), .A2(n12240), .ZN(n8384) );
  INV_X1 U10278 ( .A(n8384), .ZN(n8373) );
  NAND2_X1 U10279 ( .A1(n8012), .A2(n8373), .ZN(n11939) );
  OR2_X1 U10280 ( .A1(n8375), .A2(n11939), .ZN(n12386) );
  INV_X1 U10281 ( .A(P3_REG1_REG_29__SCAN_IN), .ZN(n13479) );
  OR2_X1 U10282 ( .A1(n8349), .A2(n13479), .ZN(n8018) );
  NAND2_X1 U10283 ( .A1(n8059), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n8017) );
  INV_X1 U10284 ( .A(n8014), .ZN(n8015) );
  NAND2_X1 U10285 ( .A1(n12382), .A2(P3_REG2_REG_29__SCAN_IN), .ZN(n8016) );
  NAND4_X1 U10286 ( .A1(n12386), .A2(n8018), .A3(n8017), .A4(n8016), .ZN(
        n12721) );
  NAND2_X1 U10287 ( .A1(n8478), .A2(n12721), .ZN(n12591) );
  INV_X1 U10288 ( .A(n12721), .ZN(n8019) );
  INV_X1 U10289 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n10519) );
  INV_X1 U10290 ( .A(SI_0_), .ZN(n9615) );
  OR2_X1 U10291 ( .A1(n8066), .A2(n9615), .ZN(n8022) );
  INV_X1 U10292 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n9614) );
  NAND2_X1 U10293 ( .A1(n9614), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n8020) );
  AND2_X1 U10294 ( .A1(n8029), .A2(n8020), .ZN(n9332) );
  OR2_X1 U10295 ( .A1(n8305), .A2(n9332), .ZN(n8021) );
  OAI211_X1 U10296 ( .C1(n10519), .C2(n10021), .A(n8022), .B(n8021), .ZN(
        n10716) );
  INV_X1 U10297 ( .A(n10716), .ZN(n9876) );
  NAND2_X1 U10298 ( .A1(n12381), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n8026) );
  NAND2_X1 U10299 ( .A1(n8386), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n8025) );
  NAND2_X1 U10300 ( .A1(n8059), .A2(P3_REG0_REG_0__SCAN_IN), .ZN(n8024) );
  NAND2_X1 U10301 ( .A1(n12382), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n8023) );
  NAND4_X1 U10302 ( .A1(n8026), .A2(n8025), .A3(n8024), .A4(n8023), .ZN(n12638) );
  NOR2_X1 U10303 ( .A1(n9876), .A2(n12638), .ZN(n15704) );
  NAND2_X1 U10304 ( .A1(n8059), .A2(P3_REG0_REG_1__SCAN_IN), .ZN(n8028) );
  NAND2_X1 U10305 ( .A1(n12382), .A2(P3_REG2_REG_1__SCAN_IN), .ZN(n8027) );
  INV_X1 U10306 ( .A(SI_1_), .ZN(n9326) );
  OR2_X1 U10307 ( .A1(n8066), .A2(n9326), .ZN(n8035) );
  XNOR2_X1 U10308 ( .A(n8030), .B(n8029), .ZN(n9327) );
  INV_X1 U10309 ( .A(n9327), .ZN(n8031) );
  INV_X1 U10310 ( .A(P3_IR_REG_1__SCAN_IN), .ZN(n8032) );
  OR2_X1 U10311 ( .A1(n10021), .A2(n10365), .ZN(n8033) );
  NAND2_X1 U10312 ( .A1(n10321), .A2(n12442), .ZN(n15689) );
  NAND2_X1 U10313 ( .A1(n12381), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n8039) );
  NAND2_X1 U10314 ( .A1(n8386), .A2(P3_REG3_REG_2__SCAN_IN), .ZN(n8038) );
  NAND2_X1 U10315 ( .A1(n8059), .A2(P3_REG0_REG_2__SCAN_IN), .ZN(n8037) );
  NAND2_X1 U10316 ( .A1(n12382), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n8036) );
  XNOR2_X1 U10317 ( .A(n8042), .B(n8041), .ZN(n9349) );
  OR2_X1 U10318 ( .A1(n8305), .A2(n9349), .ZN(n8044) );
  OR2_X1 U10319 ( .A1(n8066), .A2(SI_2_), .ZN(n8043) );
  OAI211_X1 U10320 ( .C1(n10107), .C2(n10021), .A(n8044), .B(n8043), .ZN(
        n15690) );
  NAND2_X1 U10321 ( .A1(n12637), .A2(n15690), .ZN(n12452) );
  INV_X1 U10322 ( .A(n15692), .ZN(n12448) );
  NAND2_X1 U10323 ( .A1(n15689), .A2(n12448), .ZN(n8045) );
  NAND2_X1 U10324 ( .A1(n12381), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n8051) );
  INV_X1 U10325 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n8046) );
  INV_X1 U10326 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n8047) );
  OR2_X1 U10327 ( .A1(n8337), .A2(n8047), .ZN(n8048) );
  OR2_X1 U10328 ( .A1(n8066), .A2(SI_3_), .ZN(n8058) );
  XNOR2_X1 U10329 ( .A(n8053), .B(n8052), .ZN(n9353) );
  OR2_X1 U10330 ( .A1(n8305), .A2(n9353), .ZN(n8057) );
  NAND2_X1 U10331 ( .A1(n8054), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8055) );
  XNOR2_X1 U10332 ( .A(n8055), .B(P3_IR_REG_3__SCAN_IN), .ZN(n10280) );
  OR2_X1 U10333 ( .A1(n10021), .A2(n10280), .ZN(n8056) );
  INV_X1 U10334 ( .A(n10660), .ZN(n15732) );
  NAND2_X1 U10335 ( .A1(n8059), .A2(P3_REG0_REG_4__SCAN_IN), .ZN(n8065) );
  INV_X1 U10336 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n10859) );
  OR2_X1 U10337 ( .A1(n8337), .A2(n10859), .ZN(n8064) );
  INV_X1 U10338 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n8060) );
  OR2_X1 U10339 ( .A1(n8349), .A2(n8060), .ZN(n8063) );
  AND2_X1 U10340 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(P3_REG3_REG_3__SCAN_IN), 
        .ZN(n8061) );
  NOR2_X1 U10341 ( .A1(n8077), .A2(n8061), .ZN(n10781) );
  OR2_X1 U10342 ( .A1(n8375), .A2(n10781), .ZN(n8062) );
  OR2_X1 U10343 ( .A1(n8066), .A2(SI_4_), .ZN(n8073) );
  XNOR2_X1 U10344 ( .A(n8068), .B(n8067), .ZN(n9351) );
  OR2_X1 U10345 ( .A1(n8305), .A2(n9351), .ZN(n8072) );
  NAND2_X1 U10346 ( .A1(n8069), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8070) );
  XNOR2_X1 U10347 ( .A(n8070), .B(n7036), .ZN(n10264) );
  INV_X1 U10348 ( .A(n10264), .ZN(n10258) );
  OR2_X1 U10349 ( .A1(n10021), .A2(n10258), .ZN(n8071) );
  NAND2_X1 U10350 ( .A1(n10775), .A2(n15736), .ZN(n12467) );
  INV_X1 U10351 ( .A(n10775), .ZN(n12636) );
  INV_X1 U10352 ( .A(n15736), .ZN(n8074) );
  NAND2_X1 U10353 ( .A1(n12636), .A2(n8074), .ZN(n12461) );
  NAND2_X1 U10354 ( .A1(n12467), .A2(n12461), .ZN(n12457) );
  INV_X1 U10355 ( .A(n12457), .ZN(n10856) );
  NAND2_X1 U10356 ( .A1(n8075), .A2(n12467), .ZN(n10724) );
  NAND2_X1 U10357 ( .A1(n12382), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n8082) );
  NAND2_X1 U10358 ( .A1(n12381), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n8081) );
  OR2_X1 U10359 ( .A1(n8077), .A2(n8076), .ZN(n8078) );
  NAND2_X1 U10360 ( .A1(n8088), .A2(n8078), .ZN(n10970) );
  NAND2_X1 U10361 ( .A1(n7128), .A2(n10970), .ZN(n8080) );
  NAND2_X1 U10362 ( .A1(n8059), .A2(P3_REG0_REG_5__SCAN_IN), .ZN(n8079) );
  NAND4_X1 U10363 ( .A1(n8082), .A2(n8081), .A3(n8080), .A4(n8079), .ZN(n12635) );
  NOR2_X1 U10364 ( .A1(n8069), .A2(P3_IR_REG_4__SCAN_IN), .ZN(n8097) );
  OR2_X1 U10365 ( .A1(n8097), .A2(n13054), .ZN(n8083) );
  XNOR2_X1 U10366 ( .A(n8083), .B(n8096), .ZN(n10337) );
  XNOR2_X1 U10367 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .ZN(n8084) );
  XNOR2_X1 U10368 ( .A(n8085), .B(n8084), .ZN(n9357) );
  OR2_X1 U10369 ( .A1(n8305), .A2(n9357), .ZN(n8087) );
  OR2_X1 U10370 ( .A1(n8066), .A2(SI_5_), .ZN(n8086) );
  OAI211_X1 U10371 ( .C1(n10333), .C2(n10021), .A(n8087), .B(n8086), .ZN(
        n15743) );
  OR2_X1 U10372 ( .A1(n12635), .A2(n15743), .ZN(n12463) );
  NAND2_X1 U10373 ( .A1(n12635), .A2(n15743), .ZN(n12470) );
  NAND2_X1 U10374 ( .A1(n12463), .A2(n12470), .ZN(n12468) );
  INV_X1 U10375 ( .A(n12468), .ZN(n12462) );
  NAND2_X1 U10376 ( .A1(n12382), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n8093) );
  NAND2_X1 U10377 ( .A1(n12381), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n8092) );
  NAND2_X1 U10378 ( .A1(n8088), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n8089) );
  NAND2_X1 U10379 ( .A1(n8102), .A2(n8089), .ZN(n11057) );
  NAND2_X1 U10380 ( .A1(n7128), .A2(n11057), .ZN(n8091) );
  NAND2_X1 U10381 ( .A1(n8059), .A2(P3_REG0_REG_6__SCAN_IN), .ZN(n8090) );
  NAND4_X1 U10382 ( .A1(n8093), .A2(n8092), .A3(n8091), .A4(n8090), .ZN(n12634) );
  INV_X1 U10383 ( .A(SI_6_), .ZN(n9328) );
  OR2_X1 U10384 ( .A1(n8066), .A2(n9328), .ZN(n8101) );
  XNOR2_X1 U10385 ( .A(n8095), .B(n8094), .ZN(n9329) );
  OR2_X1 U10386 ( .A1(n8305), .A2(n9329), .ZN(n8100) );
  NAND2_X1 U10387 ( .A1(n8097), .A2(n8096), .ZN(n8108) );
  NAND2_X1 U10388 ( .A1(n8108), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8098) );
  XNOR2_X1 U10389 ( .A(n8098), .B(P3_IR_REG_6__SCAN_IN), .ZN(n10393) );
  OR2_X1 U10390 ( .A1(n10021), .A2(n10401), .ZN(n8099) );
  NAND2_X1 U10391 ( .A1(n12634), .A2(n11041), .ZN(n12471) );
  AND2_X1 U10392 ( .A1(n8102), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n8103) );
  NOR2_X1 U10393 ( .A1(n8128), .A2(n8103), .ZN(n11165) );
  OR2_X1 U10394 ( .A1(n8375), .A2(n11165), .ZN(n8107) );
  NAND2_X1 U10395 ( .A1(n12382), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n8106) );
  NAND2_X1 U10396 ( .A1(n12381), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n8105) );
  NAND2_X1 U10397 ( .A1(n8059), .A2(P3_REG0_REG_7__SCAN_IN), .ZN(n8104) );
  NAND4_X1 U10398 ( .A1(n8107), .A2(n8106), .A3(n8105), .A4(n8104), .ZN(n12633) );
  NAND2_X1 U10399 ( .A1(n8122), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8110) );
  XNOR2_X1 U10400 ( .A(n8110), .B(n8109), .ZN(n10613) );
  INV_X1 U10401 ( .A(n10613), .ZN(n10599) );
  XNOR2_X1 U10402 ( .A(n8112), .B(n8111), .ZN(n9355) );
  OR2_X1 U10403 ( .A1(n8305), .A2(n9355), .ZN(n8114) );
  OR2_X1 U10404 ( .A1(n8066), .A2(SI_7_), .ZN(n8113) );
  OAI211_X1 U10405 ( .C1(n10599), .C2(n10021), .A(n8114), .B(n8113), .ZN(
        n12479) );
  NAND2_X1 U10406 ( .A1(n11150), .A2(n12477), .ZN(n8116) );
  INV_X1 U10407 ( .A(n12633), .ZN(n11144) );
  INV_X1 U10408 ( .A(n12479), .ZN(n15756) );
  NAND2_X1 U10409 ( .A1(n11144), .A2(n15756), .ZN(n8115) );
  NAND2_X1 U10410 ( .A1(n8059), .A2(P3_REG0_REG_8__SCAN_IN), .ZN(n8121) );
  INV_X1 U10411 ( .A(P3_REG2_REG_8__SCAN_IN), .ZN(n11146) );
  OR2_X1 U10412 ( .A1(n8337), .A2(n11146), .ZN(n8120) );
  INV_X1 U10413 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n8117) );
  OR2_X1 U10414 ( .A1(n8349), .A2(n8117), .ZN(n8119) );
  XNOR2_X1 U10415 ( .A(n8128), .B(P3_REG3_REG_8__SCAN_IN), .ZN(n11254) );
  OR2_X1 U10416 ( .A1(n8375), .A2(n11254), .ZN(n8118) );
  OAI21_X1 U10417 ( .B1(n8122), .B2(P3_IR_REG_7__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8123) );
  XNOR2_X1 U10418 ( .A(n8123), .B(P3_IR_REG_8__SCAN_IN), .ZN(n10611) );
  INV_X1 U10419 ( .A(SI_8_), .ZN(n9324) );
  OR2_X1 U10420 ( .A1(n8066), .A2(n9324), .ZN(n8127) );
  XNOR2_X1 U10421 ( .A(n8125), .B(n8124), .ZN(n9325) );
  OR2_X1 U10422 ( .A1(n8305), .A2(n9325), .ZN(n8126) );
  OAI211_X1 U10423 ( .C1(n10021), .C2(n11024), .A(n8127), .B(n8126), .ZN(
        n15769) );
  NAND2_X1 U10424 ( .A1(n11136), .A2(n15769), .ZN(n12487) );
  INV_X1 U10425 ( .A(n11136), .ZN(n12632) );
  INV_X1 U10426 ( .A(n15769), .ZN(n11253) );
  NAND2_X1 U10427 ( .A1(n12632), .A2(n11253), .ZN(n12486) );
  NAND2_X1 U10428 ( .A1(n12381), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n8133) );
  NAND2_X1 U10429 ( .A1(n8059), .A2(P3_REG0_REG_9__SCAN_IN), .ZN(n8132) );
  INV_X1 U10430 ( .A(P3_REG3_REG_8__SCAN_IN), .ZN(n13445) );
  INV_X1 U10431 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n13429) );
  AOI21_X1 U10432 ( .B1(n8128), .B2(n13445), .A(n13429), .ZN(n8129) );
  OR2_X1 U10433 ( .A1(n8145), .A2(n8129), .ZN(n11137) );
  NAND2_X1 U10434 ( .A1(n7128), .A2(n11137), .ZN(n8131) );
  NAND2_X1 U10435 ( .A1(n12382), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n8130) );
  NAND4_X1 U10436 ( .A1(n8133), .A2(n8132), .A3(n8131), .A4(n8130), .ZN(n12631) );
  XNOR2_X1 U10437 ( .A(n8135), .B(n8134), .ZN(n14926) );
  OR2_X1 U10438 ( .A1(n8305), .A2(n14926), .ZN(n8142) );
  OR2_X1 U10439 ( .A1(n8066), .A2(SI_9_), .ZN(n8141) );
  NOR2_X1 U10440 ( .A1(n8136), .A2(n13054), .ZN(n8137) );
  MUX2_X1 U10441 ( .A(n13054), .B(n8137), .S(P3_IR_REG_9__SCAN_IN), .Z(n8139)
         );
  OR2_X1 U10442 ( .A1(n8139), .A2(n8138), .ZN(n14928) );
  OR2_X1 U10443 ( .A1(n10021), .A2(n15605), .ZN(n8140) );
  NOR2_X1 U10444 ( .A1(n12631), .A2(n11403), .ZN(n12492) );
  NAND2_X1 U10445 ( .A1(n12631), .A2(n11403), .ZN(n12491) );
  NAND2_X1 U10446 ( .A1(n8059), .A2(P3_REG0_REG_10__SCAN_IN), .ZN(n8150) );
  INV_X1 U10447 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n8143) );
  OR2_X1 U10448 ( .A1(n8349), .A2(n8143), .ZN(n8149) );
  OR2_X1 U10449 ( .A1(n8145), .A2(n8144), .ZN(n8146) );
  AND2_X1 U10450 ( .A1(n8159), .A2(n8146), .ZN(n15594) );
  OR2_X1 U10451 ( .A1(n8375), .A2(n15594), .ZN(n8148) );
  INV_X1 U10452 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n11343) );
  OR2_X1 U10453 ( .A1(n8337), .A2(n11343), .ZN(n8147) );
  OR2_X1 U10454 ( .A1(n8138), .A2(n13054), .ZN(n8151) );
  XNOR2_X1 U10455 ( .A(n8151), .B(n8165), .ZN(n12655) );
  INV_X1 U10456 ( .A(n12655), .ZN(n12679) );
  OR2_X1 U10457 ( .A1(n8066), .A2(SI_10_), .ZN(n8155) );
  XNOR2_X1 U10458 ( .A(n8153), .B(n8152), .ZN(n9345) );
  OR2_X1 U10459 ( .A1(n8305), .A2(n9345), .ZN(n8154) );
  OAI211_X1 U10460 ( .C1(n12679), .C2(n10021), .A(n8155), .B(n8154), .ZN(
        n15580) );
  NAND2_X1 U10461 ( .A1(n12498), .A2(n15580), .ZN(n8156) );
  INV_X1 U10462 ( .A(n15580), .ZN(n12497) );
  NAND2_X1 U10463 ( .A1(n12630), .A2(n12497), .ZN(n11410) );
  INV_X1 U10464 ( .A(n11341), .ZN(n12503) );
  NAND2_X1 U10465 ( .A1(n11342), .A2(n12503), .ZN(n8158) );
  NAND2_X1 U10466 ( .A1(n12630), .A2(n15580), .ZN(n8157) );
  NAND2_X1 U10467 ( .A1(n12382), .A2(P3_REG2_REG_11__SCAN_IN), .ZN(n8164) );
  NAND2_X1 U10468 ( .A1(n12381), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n8163) );
  NAND2_X1 U10469 ( .A1(n8159), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n8160) );
  NAND2_X1 U10470 ( .A1(n8173), .A2(n8160), .ZN(n11417) );
  NAND2_X1 U10471 ( .A1(n7128), .A2(n11417), .ZN(n8162) );
  NAND2_X1 U10472 ( .A1(n8059), .A2(P3_REG0_REG_11__SCAN_IN), .ZN(n8161) );
  NAND4_X1 U10473 ( .A1(n8164), .A2(n8163), .A3(n8162), .A4(n8161), .ZN(n12629) );
  NAND2_X1 U10474 ( .A1(n8138), .A2(n8165), .ZN(n8183) );
  NAND2_X1 U10475 ( .A1(n8183), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8167) );
  XNOR2_X1 U10476 ( .A(n8167), .B(n8166), .ZN(n15622) );
  OR2_X1 U10477 ( .A1(n8066), .A2(SI_11_), .ZN(n8171) );
  XNOR2_X1 U10478 ( .A(n9553), .B(P1_DATAO_REG_11__SCAN_IN), .ZN(n8168) );
  XNOR2_X1 U10479 ( .A(n8169), .B(n8168), .ZN(n9347) );
  OR2_X1 U10480 ( .A1(n8305), .A2(n9347), .ZN(n8170) );
  OAI211_X1 U10481 ( .C1(n12682), .C2(n10021), .A(n8171), .B(n8170), .ZN(
        n13048) );
  OR2_X1 U10482 ( .A1(n12629), .A2(n13048), .ZN(n12505) );
  NAND2_X1 U10483 ( .A1(n12629), .A2(n13048), .ZN(n12506) );
  NAND2_X1 U10484 ( .A1(n12505), .A2(n12506), .ZN(n12414) );
  NAND2_X1 U10485 ( .A1(n11415), .A2(n12505), .ZN(n12909) );
  NAND2_X1 U10486 ( .A1(n12382), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n8178) );
  NAND2_X1 U10487 ( .A1(n12381), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n8177) );
  NAND2_X1 U10488 ( .A1(n8173), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n8174) );
  NAND2_X1 U10489 ( .A1(n8188), .A2(n8174), .ZN(n12910) );
  NAND2_X1 U10490 ( .A1(n7128), .A2(n12910), .ZN(n8176) );
  NAND2_X1 U10491 ( .A1(n8059), .A2(P3_REG0_REG_12__SCAN_IN), .ZN(n8175) );
  NAND4_X1 U10492 ( .A1(n8178), .A2(n8177), .A3(n8176), .A4(n8175), .ZN(n12628) );
  NAND2_X1 U10493 ( .A1(n8180), .A2(n8179), .ZN(n8181) );
  NAND2_X1 U10494 ( .A1(n8182), .A2(n8181), .ZN(n9366) );
  OR2_X1 U10495 ( .A1(n8305), .A2(n9366), .ZN(n8187) );
  OR2_X1 U10496 ( .A1(n8066), .A2(n9367), .ZN(n8186) );
  NAND2_X1 U10497 ( .A1(n8197), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8184) );
  XNOR2_X1 U10498 ( .A(n8184), .B(P3_IR_REG_12__SCAN_IN), .ZN(n12685) );
  OR2_X1 U10499 ( .A1(n10021), .A2(n15640), .ZN(n8185) );
  NAND2_X1 U10500 ( .A1(n12628), .A2(n13044), .ZN(n12509) );
  NAND2_X1 U10501 ( .A1(n12510), .A2(n12509), .ZN(n8403) );
  NAND2_X1 U10502 ( .A1(n12909), .A2(n12908), .ZN(n12907) );
  NAND2_X1 U10503 ( .A1(n12907), .A2(n12510), .ZN(n15096) );
  NAND2_X1 U10504 ( .A1(n8059), .A2(P3_REG0_REG_13__SCAN_IN), .ZN(n8195) );
  AND2_X1 U10505 ( .A1(n8188), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n8189) );
  NOR2_X1 U10506 ( .A1(n8213), .A2(n8189), .ZN(n15094) );
  OR2_X1 U10507 ( .A1(n8375), .A2(n15094), .ZN(n8194) );
  INV_X1 U10508 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n8190) );
  OR2_X1 U10509 ( .A1(n8337), .A2(n8190), .ZN(n8193) );
  INV_X1 U10510 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n8191) );
  OR2_X1 U10511 ( .A1(n8349), .A2(n8191), .ZN(n8192) );
  XNOR2_X1 U10512 ( .A(n8196), .B(n6979), .ZN(n14930) );
  NAND2_X1 U10513 ( .A1(n14930), .A2(n12394), .ZN(n8204) );
  NOR2_X1 U10514 ( .A1(n8197), .A2(P3_IR_REG_12__SCAN_IN), .ZN(n8200) );
  NOR2_X1 U10515 ( .A1(n8200), .A2(n13054), .ZN(n8198) );
  MUX2_X1 U10516 ( .A(n13054), .B(n8198), .S(P3_IR_REG_13__SCAN_IN), .Z(n8202)
         );
  INV_X1 U10517 ( .A(P3_IR_REG_13__SCAN_IN), .ZN(n8199) );
  NAND2_X1 U10518 ( .A1(n8200), .A2(n8199), .ZN(n8224) );
  INV_X1 U10519 ( .A(n8224), .ZN(n8201) );
  AOI22_X1 U10520 ( .A1(n8282), .A2(n14929), .B1(n8281), .B2(n15655), .ZN(
        n8203) );
  NAND2_X1 U10521 ( .A1(n8204), .A2(n8203), .ZN(n12198) );
  NOR2_X1 U10522 ( .A1(n15013), .A2(n12198), .ZN(n12514) );
  NAND2_X1 U10523 ( .A1(n15013), .A2(n12198), .ZN(n12516) );
  XNOR2_X1 U10524 ( .A(n8207), .B(n8206), .ZN(n14939) );
  NAND2_X1 U10525 ( .A1(n14939), .A2(n12394), .ZN(n8211) );
  NAND2_X1 U10526 ( .A1(n8224), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8209) );
  INV_X1 U10527 ( .A(P3_IR_REG_14__SCAN_IN), .ZN(n8208) );
  XNOR2_X1 U10528 ( .A(n8209), .B(n8208), .ZN(n15676) );
  AOI22_X1 U10529 ( .A1(n8282), .A2(n14937), .B1(n8281), .B2(n15676), .ZN(
        n8210) );
  NAND2_X1 U10530 ( .A1(n8211), .A2(n8210), .ZN(n15105) );
  NAND2_X1 U10531 ( .A1(n12381), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n8218) );
  NAND2_X1 U10532 ( .A1(n8059), .A2(P3_REG0_REG_14__SCAN_IN), .ZN(n8217) );
  OR2_X1 U10533 ( .A1(n8213), .A2(n8212), .ZN(n8214) );
  NAND2_X1 U10534 ( .A1(n8229), .A2(n8214), .ZN(n12896) );
  NAND2_X1 U10535 ( .A1(n7128), .A2(n12896), .ZN(n8216) );
  NAND2_X1 U10536 ( .A1(n12382), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n8215) );
  NAND4_X1 U10537 ( .A1(n8218), .A2(n8217), .A3(n8216), .A4(n8215), .ZN(n12627) );
  NAND2_X1 U10538 ( .A1(n15105), .A2(n12627), .ZN(n12523) );
  INV_X1 U10539 ( .A(n12523), .ZN(n8219) );
  OR2_X1 U10540 ( .A1(n15105), .A2(n12627), .ZN(n12520) );
  NAND2_X1 U10541 ( .A1(n8221), .A2(n8220), .ZN(n8222) );
  NAND2_X1 U10542 ( .A1(n8223), .A2(n8222), .ZN(n9560) );
  NAND2_X1 U10543 ( .A1(n9560), .A2(n12394), .ZN(n8228) );
  OAI21_X1 U10544 ( .B1(n8224), .B2(P3_IR_REG_14__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8226) );
  INV_X1 U10545 ( .A(P3_IR_REG_15__SCAN_IN), .ZN(n8225) );
  XNOR2_X1 U10546 ( .A(n8226), .B(n8225), .ZN(n15032) );
  AOI22_X1 U10547 ( .A1(n8282), .A2(n9561), .B1(n8281), .B2(n15032), .ZN(n8227) );
  INV_X1 U10548 ( .A(n13040), .ZN(n12373) );
  NAND2_X1 U10549 ( .A1(n8059), .A2(P3_REG0_REG_15__SCAN_IN), .ZN(n8234) );
  INV_X1 U10550 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n12976) );
  OR2_X1 U10551 ( .A1(n8349), .A2(n12976), .ZN(n8233) );
  NAND2_X1 U10552 ( .A1(n8229), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n8230) );
  AND2_X1 U10553 ( .A1(n8243), .A2(n8230), .ZN(n12368) );
  OR2_X1 U10554 ( .A1(n8375), .A2(n12368), .ZN(n8232) );
  INV_X1 U10555 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n15027) );
  OR2_X1 U10556 ( .A1(n8337), .A2(n15027), .ZN(n8231) );
  NAND2_X1 U10557 ( .A1(n12373), .A2(n12362), .ZN(n12529) );
  NAND2_X1 U10558 ( .A1(n13040), .A2(n12868), .ZN(n12524) );
  NAND2_X1 U10559 ( .A1(n8236), .A2(n8235), .ZN(n8238) );
  AND2_X1 U10560 ( .A1(n8237), .A2(n8238), .ZN(n9776) );
  NAND2_X1 U10561 ( .A1(n9776), .A2(n12394), .ZN(n8242) );
  NAND2_X1 U10562 ( .A1(n8239), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8240) );
  XNOR2_X1 U10563 ( .A(n8240), .B(P3_IR_REG_16__SCAN_IN), .ZN(n15042) );
  AOI22_X1 U10564 ( .A1(n8282), .A2(SI_16_), .B1(n8281), .B2(n15042), .ZN(
        n8241) );
  NAND2_X1 U10565 ( .A1(n8242), .A2(n8241), .ZN(n15005) );
  INV_X1 U10566 ( .A(n15005), .ZN(n13036) );
  INV_X1 U10567 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n12972) );
  OR2_X1 U10568 ( .A1(n8349), .A2(n12972), .ZN(n8248) );
  INV_X1 U10569 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n13407) );
  OR2_X1 U10570 ( .A1(n8337), .A2(n13407), .ZN(n8247) );
  NAND2_X1 U10571 ( .A1(n8243), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n8244) );
  NAND2_X1 U10572 ( .A1(n8244), .A2(n7910), .ZN(n15001) );
  NAND2_X1 U10573 ( .A1(n7128), .A2(n15001), .ZN(n8246) );
  NAND2_X1 U10574 ( .A1(n8059), .A2(P3_REG0_REG_16__SCAN_IN), .ZN(n8245) );
  NAND4_X1 U10575 ( .A1(n8248), .A2(n8247), .A3(n8246), .A4(n8245), .ZN(n12626) );
  NAND2_X1 U10576 ( .A1(n13036), .A2(n12626), .ZN(n12532) );
  INV_X1 U10577 ( .A(n12626), .ZN(n12856) );
  NAND2_X1 U10578 ( .A1(n15005), .A2(n12856), .ZN(n12530) );
  NAND2_X1 U10579 ( .A1(n12875), .A2(n12874), .ZN(n8249) );
  NAND2_X1 U10580 ( .A1(n8249), .A2(n12530), .ZN(n12860) );
  XNOR2_X1 U10581 ( .A(n8251), .B(n8250), .ZN(n9802) );
  NAND2_X1 U10582 ( .A1(n9802), .A2(n12394), .ZN(n8255) );
  NAND2_X1 U10583 ( .A1(n6803), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8252) );
  MUX2_X1 U10584 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8252), .S(
        P3_IR_REG_17__SCAN_IN), .Z(n8253) );
  NAND2_X1 U10585 ( .A1(n8253), .A2(n8263), .ZN(n12699) );
  AOI22_X1 U10586 ( .A1(n8282), .A2(n13439), .B1(n8281), .B2(n12699), .ZN(
        n8254) );
  AND2_X1 U10587 ( .A1(P3_REG3_REG_17__SCAN_IN), .A2(n7910), .ZN(n8256) );
  NOR2_X1 U10588 ( .A1(n8271), .A2(n8256), .ZN(n12861) );
  OR2_X1 U10589 ( .A1(n8375), .A2(n12861), .ZN(n8260) );
  INV_X1 U10590 ( .A(P3_REG0_REG_17__SCAN_IN), .ZN(n13421) );
  OR2_X1 U10591 ( .A1(n8429), .A2(n13421), .ZN(n8259) );
  NAND2_X1 U10592 ( .A1(n12381), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n8258) );
  NAND2_X1 U10593 ( .A1(n12382), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n8257) );
  NAND4_X1 U10594 ( .A1(n8260), .A2(n8259), .A3(n8258), .A4(n8257), .ZN(n12870) );
  INV_X1 U10595 ( .A(n12854), .ZN(n12859) );
  NAND2_X1 U10596 ( .A1(n12860), .A2(n12859), .ZN(n12858) );
  OR2_X1 U10597 ( .A1(n13032), .A2(n12870), .ZN(n12539) );
  NAND2_X1 U10598 ( .A1(n12858), .A2(n12539), .ZN(n12847) );
  XNOR2_X1 U10599 ( .A(n8262), .B(n8261), .ZN(n14946) );
  NAND2_X1 U10600 ( .A1(n14946), .A2(n12394), .ZN(n8269) );
  NAND2_X1 U10601 ( .A1(n8263), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8264) );
  MUX2_X1 U10602 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8264), .S(
        P3_IR_REG_18__SCAN_IN), .Z(n8265) );
  INV_X1 U10603 ( .A(n8265), .ZN(n8267) );
  NOR2_X1 U10604 ( .A1(n8267), .A2(n8266), .ZN(n15073) );
  AOI22_X1 U10605 ( .A1(n8282), .A2(SI_18_), .B1(n8281), .B2(n15073), .ZN(
        n8268) );
  NAND2_X1 U10606 ( .A1(n8269), .A2(n8268), .ZN(n12343) );
  NAND2_X1 U10607 ( .A1(n12382), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n8277) );
  INV_X1 U10608 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n13425) );
  OR2_X1 U10609 ( .A1(n8349), .A2(n13425), .ZN(n8276) );
  NOR2_X1 U10610 ( .A1(n8271), .A2(n8270), .ZN(n8272) );
  OR2_X1 U10611 ( .A1(n8285), .A2(n8272), .ZN(n12848) );
  INV_X1 U10612 ( .A(n12848), .ZN(n8273) );
  OR2_X1 U10613 ( .A1(n8375), .A2(n8273), .ZN(n8275) );
  INV_X1 U10614 ( .A(P3_REG0_REG_18__SCAN_IN), .ZN(n13027) );
  OR2_X1 U10615 ( .A1(n8429), .A2(n13027), .ZN(n8274) );
  OR2_X1 U10616 ( .A1(n12343), .A2(n12857), .ZN(n12536) );
  NAND2_X1 U10617 ( .A1(n12343), .A2(n12857), .ZN(n12542) );
  INV_X1 U10618 ( .A(n12846), .ZN(n8278) );
  XNOR2_X1 U10619 ( .A(n8280), .B(n8279), .ZN(n10081) );
  NAND2_X1 U10620 ( .A1(n10081), .A2(n12394), .ZN(n8284) );
  AOI22_X1 U10621 ( .A1(n8282), .A2(SI_19_), .B1(n12706), .B2(n8281), .ZN(
        n8283) );
  INV_X1 U10622 ( .A(P3_REG0_REG_19__SCAN_IN), .ZN(n13243) );
  OR2_X1 U10623 ( .A1(n8429), .A2(n13243), .ZN(n8290) );
  NAND2_X1 U10624 ( .A1(n12381), .A2(P3_REG1_REG_19__SCAN_IN), .ZN(n8289) );
  NAND2_X1 U10625 ( .A1(n12382), .A2(P3_REG2_REG_19__SCAN_IN), .ZN(n8288) );
  NOR2_X1 U10626 ( .A1(n8285), .A2(n12264), .ZN(n8286) );
  OR2_X1 U10627 ( .A1(n8295), .A2(n8286), .ZN(n12835) );
  NAND2_X1 U10628 ( .A1(n7128), .A2(n12835), .ZN(n8287) );
  NAND4_X1 U10629 ( .A1(n8290), .A2(n8289), .A3(n8288), .A4(n8287), .ZN(n12624) );
  NOR2_X1 U10630 ( .A1(n12411), .A2(n12845), .ZN(n12547) );
  NAND2_X1 U10631 ( .A1(n12411), .A2(n12845), .ZN(n12546) );
  XNOR2_X1 U10632 ( .A(n8292), .B(P2_DATAO_REG_20__SCAN_IN), .ZN(n10461) );
  NAND2_X1 U10633 ( .A1(n10461), .A2(n12394), .ZN(n8294) );
  INV_X1 U10634 ( .A(SI_20_), .ZN(n10463) );
  NAND2_X1 U10635 ( .A1(n12382), .A2(P3_REG2_REG_20__SCAN_IN), .ZN(n8300) );
  INV_X1 U10636 ( .A(P3_REG1_REG_20__SCAN_IN), .ZN(n13219) );
  OR2_X1 U10637 ( .A1(n8349), .A2(n13219), .ZN(n8299) );
  OR2_X1 U10638 ( .A1(n8295), .A2(n12328), .ZN(n8296) );
  AND2_X1 U10639 ( .A1(n8309), .A2(n8296), .ZN(n12821) );
  OR2_X1 U10640 ( .A1(n8375), .A2(n12821), .ZN(n8298) );
  INV_X1 U10641 ( .A(P3_REG0_REG_20__SCAN_IN), .ZN(n13019) );
  OR2_X1 U10642 ( .A1(n8429), .A2(n13019), .ZN(n8297) );
  NAND2_X1 U10643 ( .A1(n12954), .A2(n12216), .ZN(n12551) );
  NAND2_X1 U10644 ( .A1(n12826), .A2(n12825), .ZN(n12824) );
  NAND2_X1 U10645 ( .A1(n12824), .A2(n12550), .ZN(n12809) );
  NAND2_X1 U10646 ( .A1(n8302), .A2(n8301), .ZN(n8303) );
  NAND2_X1 U10647 ( .A1(n8304), .A2(n8303), .ZN(n10565) );
  OR2_X1 U10648 ( .A1(n10565), .A2(n8305), .ZN(n8307) );
  INV_X1 U10649 ( .A(SI_21_), .ZN(n10564) );
  OR2_X1 U10650 ( .A1(n8066), .A2(n10564), .ZN(n8306) );
  INV_X1 U10651 ( .A(n13018), .ZN(n12283) );
  NAND2_X1 U10652 ( .A1(n12381), .A2(P3_REG1_REG_21__SCAN_IN), .ZN(n8313) );
  INV_X1 U10653 ( .A(P3_REG2_REG_21__SCAN_IN), .ZN(n12811) );
  OR2_X1 U10654 ( .A1(n8337), .A2(n12811), .ZN(n8312) );
  AOI21_X1 U10655 ( .B1(n8309), .B2(P3_REG3_REG_21__SCAN_IN), .A(n8308), .ZN(
        n12810) );
  OR2_X1 U10656 ( .A1(n8375), .A2(n12810), .ZN(n8311) );
  INV_X1 U10657 ( .A(P3_REG0_REG_21__SCAN_IN), .ZN(n13016) );
  OR2_X1 U10658 ( .A1(n8429), .A2(n13016), .ZN(n8310) );
  NAND2_X1 U10659 ( .A1(n12283), .A2(n12217), .ZN(n12554) );
  NAND2_X1 U10660 ( .A1(n13018), .A2(n12622), .ZN(n12555) );
  XNOR2_X1 U10661 ( .A(n8315), .B(n8314), .ZN(n10767) );
  NAND2_X1 U10662 ( .A1(n10767), .A2(n12394), .ZN(n8317) );
  AND2_X1 U10663 ( .A1(P3_REG3_REG_22__SCAN_IN), .A2(n8318), .ZN(n8319) );
  NOR2_X1 U10664 ( .A1(n8338), .A2(n8319), .ZN(n12336) );
  OR2_X1 U10665 ( .A1(n8375), .A2(n12336), .ZN(n8323) );
  NAND2_X1 U10666 ( .A1(n12382), .A2(P3_REG2_REG_22__SCAN_IN), .ZN(n8322) );
  NAND2_X1 U10667 ( .A1(n12381), .A2(P3_REG1_REG_22__SCAN_IN), .ZN(n8321) );
  NAND2_X1 U10668 ( .A1(n8059), .A2(P3_REG0_REG_22__SCAN_IN), .ZN(n8320) );
  NAND4_X1 U10669 ( .A1(n8323), .A2(n8322), .A3(n8321), .A4(n8320), .ZN(n12621) );
  INV_X1 U10670 ( .A(n12621), .ZN(n8324) );
  NAND2_X1 U10671 ( .A1(n12338), .A2(n8324), .ZN(n12559) );
  XNOR2_X1 U10672 ( .A(n8326), .B(n8325), .ZN(n10967) );
  NAND2_X1 U10673 ( .A1(n10967), .A2(n12394), .ZN(n8328) );
  INV_X1 U10674 ( .A(SI_23_), .ZN(n10969) );
  XNOR2_X1 U10675 ( .A(n8338), .B(P3_REG3_REG_23__SCAN_IN), .ZN(n12256) );
  OR2_X1 U10676 ( .A1(n8375), .A2(n12256), .ZN(n8332) );
  NAND2_X1 U10677 ( .A1(n12382), .A2(P3_REG2_REG_23__SCAN_IN), .ZN(n8331) );
  NAND2_X1 U10678 ( .A1(n12381), .A2(P3_REG1_REG_23__SCAN_IN), .ZN(n8330) );
  NAND2_X1 U10679 ( .A1(n8059), .A2(P3_REG0_REG_23__SCAN_IN), .ZN(n8329) );
  NAND4_X1 U10680 ( .A1(n8332), .A2(n8331), .A3(n8330), .A4(n8329), .ZN(n12620) );
  XNOR2_X1 U10681 ( .A(n12563), .B(n12620), .ZN(n12782) );
  NAND2_X1 U10682 ( .A1(n12780), .A2(n12782), .ZN(n12779) );
  INV_X1 U10683 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n11510) );
  NAND2_X1 U10684 ( .A1(n11166), .A2(n12394), .ZN(n8335) );
  INV_X1 U10685 ( .A(SI_24_), .ZN(n11167) );
  NAND2_X1 U10686 ( .A1(n12381), .A2(P3_REG1_REG_24__SCAN_IN), .ZN(n8344) );
  INV_X1 U10687 ( .A(P3_REG2_REG_24__SCAN_IN), .ZN(n8336) );
  OR2_X1 U10688 ( .A1(n8337), .A2(n8336), .ZN(n8343) );
  INV_X1 U10689 ( .A(P3_REG3_REG_23__SCAN_IN), .ZN(n13426) );
  NAND2_X1 U10690 ( .A1(n8338), .A2(n13426), .ZN(n8339) );
  NAND2_X1 U10691 ( .A1(n8339), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n8340) );
  AND2_X1 U10692 ( .A1(n8340), .A2(n8350), .ZN(n12322) );
  OR2_X1 U10693 ( .A1(n8375), .A2(n12322), .ZN(n8342) );
  INV_X1 U10694 ( .A(P3_REG0_REG_24__SCAN_IN), .ZN(n13005) );
  OR2_X1 U10695 ( .A1(n8429), .A2(n13005), .ZN(n8341) );
  INV_X1 U10696 ( .A(n12620), .ZN(n12562) );
  NOR2_X1 U10697 ( .A1(n12563), .A2(n12562), .ZN(n12770) );
  AOI22_X1 U10698 ( .A1(P2_DATAO_REG_25__SCAN_IN), .A2(
        P1_DATAO_REG_25__SCAN_IN), .B1(n14037), .B2(n14816), .ZN(n8345) );
  XNOR2_X1 U10699 ( .A(n8346), .B(n8345), .ZN(n11389) );
  NAND2_X1 U10700 ( .A1(n11389), .A2(n12394), .ZN(n8348) );
  INV_X1 U10701 ( .A(SI_25_), .ZN(n11391) );
  NAND2_X1 U10702 ( .A1(n12382), .A2(P3_REG2_REG_25__SCAN_IN), .ZN(n8355) );
  INV_X1 U10703 ( .A(P3_REG1_REG_25__SCAN_IN), .ZN(n13229) );
  OR2_X1 U10704 ( .A1(n8349), .A2(n13229), .ZN(n8354) );
  NAND2_X1 U10705 ( .A1(n8350), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n8351) );
  AND2_X1 U10706 ( .A1(n8361), .A2(n8351), .ZN(n12303) );
  OR2_X1 U10707 ( .A1(n8375), .A2(n12303), .ZN(n8353) );
  INV_X1 U10708 ( .A(P3_REG0_REG_25__SCAN_IN), .ZN(n13000) );
  OR2_X1 U10709 ( .A1(n8429), .A2(n13000), .ZN(n8352) );
  OR2_X1 U10710 ( .A1(n12296), .A2(n12229), .ZN(n12571) );
  NAND2_X1 U10711 ( .A1(n12296), .A2(n12229), .ZN(n12736) );
  NAND2_X1 U10712 ( .A1(n12571), .A2(n12736), .ZN(n12753) );
  INV_X1 U10713 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n14810) );
  AOI22_X1 U10714 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(n14034), .B1(
        P1_DATAO_REG_26__SCAN_IN), .B2(n14810), .ZN(n8356) );
  INV_X1 U10715 ( .A(n8356), .ZN(n8357) );
  XNOR2_X1 U10716 ( .A(n8358), .B(n8357), .ZN(n11424) );
  NAND2_X1 U10717 ( .A1(n11424), .A2(n12394), .ZN(n8360) );
  AOI21_X1 U10718 ( .B1(n8361), .B2(P3_REG3_REG_26__SCAN_IN), .A(n8372), .ZN(
        n12744) );
  OR2_X1 U10719 ( .A1(n8375), .A2(n12744), .ZN(n8365) );
  INV_X1 U10720 ( .A(P3_REG0_REG_26__SCAN_IN), .ZN(n13428) );
  OR2_X1 U10721 ( .A1(n8429), .A2(n13428), .ZN(n8364) );
  NAND2_X1 U10722 ( .A1(n12381), .A2(P3_REG1_REG_26__SCAN_IN), .ZN(n8363) );
  NAND2_X1 U10723 ( .A1(n12382), .A2(P3_REG2_REG_26__SCAN_IN), .ZN(n8362) );
  NAND4_X1 U10724 ( .A1(n8365), .A2(n8364), .A3(n8363), .A4(n8362), .ZN(n12618) );
  INV_X1 U10725 ( .A(n12618), .ZN(n12241) );
  NAND2_X1 U10726 ( .A1(n12747), .A2(n12241), .ZN(n12576) );
  NAND2_X1 U10727 ( .A1(n12575), .A2(n12576), .ZN(n12740) );
  INV_X1 U10728 ( .A(n12736), .ZN(n8366) );
  NOR2_X1 U10729 ( .A1(n12740), .A2(n8366), .ZN(n8367) );
  AOI22_X1 U10730 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(n14028), .B1(
        P1_DATAO_REG_27__SCAN_IN), .B2(n11560), .ZN(n8368) );
  XNOR2_X1 U10731 ( .A(n8369), .B(n8368), .ZN(n11507) );
  NAND2_X1 U10732 ( .A1(n11507), .A2(n12394), .ZN(n8371) );
  INV_X1 U10733 ( .A(n8372), .ZN(n8374) );
  AOI21_X1 U10734 ( .B1(P3_REG3_REG_27__SCAN_IN), .B2(n8374), .A(n8373), .ZN(
        n12242) );
  OR2_X1 U10735 ( .A1(n8375), .A2(n12242), .ZN(n8379) );
  NAND2_X1 U10736 ( .A1(n12382), .A2(P3_REG2_REG_27__SCAN_IN), .ZN(n8378) );
  NAND2_X1 U10737 ( .A1(n12381), .A2(P3_REG1_REG_27__SCAN_IN), .ZN(n8377) );
  NAND2_X1 U10738 ( .A1(n8059), .A2(P3_REG0_REG_27__SCAN_IN), .ZN(n8376) );
  INV_X1 U10739 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n14809) );
  AOI22_X1 U10740 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(n14809), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(n13246), .ZN(n8380) );
  INV_X1 U10741 ( .A(n8380), .ZN(n8381) );
  XNOR2_X1 U10742 ( .A(n8382), .B(n8381), .ZN(n13059) );
  INV_X1 U10743 ( .A(SI_28_), .ZN(n13061) );
  NOR2_X1 U10744 ( .A1(n8066), .A2(n13061), .ZN(n8383) );
  INV_X1 U10745 ( .A(n12993), .ZN(n8426) );
  NAND2_X1 U10746 ( .A1(n12381), .A2(P3_REG1_REG_28__SCAN_IN), .ZN(n8390) );
  NAND2_X1 U10747 ( .A1(n12382), .A2(P3_REG2_REG_28__SCAN_IN), .ZN(n8389) );
  NAND2_X1 U10748 ( .A1(P3_REG3_REG_28__SCAN_IN), .A2(n8384), .ZN(n8385) );
  NAND2_X1 U10749 ( .A1(n11939), .A2(n8385), .ZN(n12730) );
  NAND2_X1 U10750 ( .A1(n7128), .A2(n12730), .ZN(n8388) );
  NAND2_X1 U10751 ( .A1(n8059), .A2(P3_REG0_REG_28__SCAN_IN), .ZN(n8387) );
  NAND4_X1 U10752 ( .A1(n8390), .A2(n8389), .A3(n8388), .A4(n8387), .ZN(n12245) );
  INV_X1 U10753 ( .A(n12245), .ZN(n8391) );
  NAND2_X1 U10754 ( .A1(n8426), .A2(n8391), .ZN(n8425) );
  INV_X1 U10755 ( .A(n12722), .ZN(n8423) );
  NAND2_X1 U10756 ( .A1(n12582), .A2(n8423), .ZN(n12725) );
  NAND2_X1 U10757 ( .A1(n12993), .A2(n12245), .ZN(n12586) );
  NAND2_X1 U10758 ( .A1(n12638), .A2(n10716), .ZN(n15706) );
  NAND2_X1 U10759 ( .A1(n15705), .A2(n15706), .ZN(n8392) );
  INV_X1 U10760 ( .A(n15690), .ZN(n10483) );
  NOR2_X1 U10761 ( .A1(n12637), .A2(n10483), .ZN(n8393) );
  NAND2_X1 U10762 ( .A1(n8394), .A2(n10660), .ZN(n8395) );
  NAND2_X1 U10763 ( .A1(n12636), .A2(n15736), .ZN(n10725) );
  AND2_X1 U10764 ( .A1(n12468), .A2(n10725), .ZN(n8396) );
  INV_X1 U10765 ( .A(n12635), .ZN(n11050) );
  NAND2_X1 U10766 ( .A1(n11050), .A2(n15743), .ZN(n8397) );
  INV_X1 U10767 ( .A(n11041), .ZN(n15749) );
  NAND2_X1 U10768 ( .A1(n12634), .A2(n15749), .ZN(n8399) );
  NAND2_X1 U10769 ( .A1(n12633), .A2(n15756), .ZN(n8400) );
  NAND2_X1 U10770 ( .A1(n11136), .A2(n11253), .ZN(n8401) );
  XNOR2_X1 U10771 ( .A(n12631), .B(n11120), .ZN(n12489) );
  NAND2_X1 U10772 ( .A1(n11411), .A2(n11410), .ZN(n8402) );
  NAND2_X1 U10773 ( .A1(n8402), .A2(n12414), .ZN(n11409) );
  INV_X1 U10774 ( .A(n13048), .ZN(n11418) );
  NAND2_X1 U10775 ( .A1(n12629), .A2(n11418), .ZN(n12902) );
  NAND2_X1 U10776 ( .A1(n11409), .A2(n12902), .ZN(n8404) );
  INV_X1 U10777 ( .A(n13044), .ZN(n12912) );
  NAND2_X1 U10778 ( .A1(n12628), .A2(n12912), .ZN(n8405) );
  NAND2_X1 U10779 ( .A1(n12199), .A2(n12198), .ZN(n8406) );
  INV_X1 U10780 ( .A(n12198), .ZN(n15110) );
  NAND2_X1 U10781 ( .A1(n12520), .A2(n12523), .ZN(n12894) );
  INV_X1 U10782 ( .A(n12627), .ZN(n15018) );
  OR2_X1 U10783 ( .A1(n15018), .A2(n15105), .ZN(n8407) );
  NOR2_X1 U10784 ( .A1(n13040), .A2(n12362), .ZN(n8408) );
  NAND2_X1 U10785 ( .A1(n13040), .A2(n12362), .ZN(n8409) );
  NOR2_X1 U10786 ( .A1(n15005), .A2(n12626), .ZN(n8410) );
  INV_X1 U10787 ( .A(n12870), .ZN(n12844) );
  OR2_X1 U10788 ( .A1(n13032), .A2(n12844), .ZN(n8411) );
  NAND2_X1 U10789 ( .A1(n8412), .A2(n8411), .ZN(n12842) );
  OR2_X1 U10790 ( .A1(n12343), .A2(n12625), .ZN(n8413) );
  INV_X1 U10791 ( .A(n12216), .ZN(n12623) );
  NAND2_X1 U10792 ( .A1(n12954), .A2(n12623), .ZN(n8414) );
  AND2_X1 U10793 ( .A1(n12283), .A2(n12622), .ZN(n12408) );
  NAND2_X1 U10794 ( .A1(n13018), .A2(n12217), .ZN(n12409) );
  OR2_X1 U10795 ( .A1(n12338), .A2(n12621), .ZN(n8415) );
  NAND2_X1 U10796 ( .A1(n12563), .A2(n12620), .ZN(n8417) );
  OR2_X1 U10797 ( .A1(n12318), .A2(n6985), .ZN(n12751) );
  AND2_X1 U10798 ( .A1(n12751), .A2(n12753), .ZN(n8418) );
  NAND2_X1 U10799 ( .A1(n12296), .A2(n12619), .ZN(n8419) );
  OR2_X1 U10800 ( .A1(n12618), .A2(n12747), .ZN(n8420) );
  NAND2_X1 U10801 ( .A1(n12747), .A2(n12618), .ZN(n8421) );
  NAND2_X1 U10802 ( .A1(n12996), .A2(n8423), .ZN(n8424) );
  NAND2_X1 U10803 ( .A1(n11852), .A2(n8424), .ZN(n12717) );
  NAND2_X1 U10804 ( .A1(n12613), .A2(n12706), .ZN(n8482) );
  NAND2_X1 U10805 ( .A1(n10656), .A2(n8481), .ZN(n12402) );
  INV_X1 U10806 ( .A(n8427), .ZN(n10022) );
  NAND2_X1 U10807 ( .A1(n10022), .A2(n10016), .ZN(n10023) );
  NAND2_X1 U10808 ( .A1(n10021), .A2(n10023), .ZN(n8433) );
  AND2_X1 U10809 ( .A1(n10022), .A2(P3_B_REG_SCAN_IN), .ZN(n8428) );
  NOR2_X1 U10810 ( .A1(n15017), .A2(n8428), .ZN(n12711) );
  INV_X1 U10811 ( .A(P3_REG0_REG_30__SCAN_IN), .ZN(n15114) );
  OR2_X1 U10812 ( .A1(n8429), .A2(n15114), .ZN(n8432) );
  NAND2_X1 U10813 ( .A1(n12382), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n8431) );
  NAND2_X1 U10814 ( .A1(n12381), .A2(P3_REG1_REG_30__SCAN_IN), .ZN(n8430) );
  NAND4_X1 U10815 ( .A1(n12386), .A2(n8432), .A3(n8431), .A4(n8430), .ZN(
        n12617) );
  INV_X1 U10816 ( .A(n8433), .ZN(n8434) );
  AOI22_X1 U10817 ( .A1(n12711), .A2(n12617), .B1(n12245), .B2(n12867), .ZN(
        n8435) );
  NAND2_X1 U10818 ( .A1(n8436), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8437) );
  INV_X1 U10819 ( .A(n8440), .ZN(n8445) );
  NAND2_X1 U10820 ( .A1(n8445), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8441) );
  MUX2_X1 U10821 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8441), .S(
        P3_IR_REG_25__SCAN_IN), .Z(n8442) );
  NAND2_X1 U10822 ( .A1(n8442), .A2(n8436), .ZN(n11392) );
  NAND2_X1 U10823 ( .A1(n8443), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8444) );
  XNOR2_X1 U10824 ( .A(n11169), .B(P3_B_REG_SCAN_IN), .ZN(n8447) );
  NAND2_X1 U10825 ( .A1(n11392), .A2(n8447), .ZN(n8448) );
  INV_X1 U10826 ( .A(P3_D_REG_1__SCAN_IN), .ZN(n8449) );
  NAND2_X1 U10827 ( .A1(n9497), .A2(n8449), .ZN(n8451) );
  NAND2_X1 U10828 ( .A1(n11427), .A2(n11392), .ZN(n8450) );
  INV_X1 U10829 ( .A(P3_D_REG_0__SCAN_IN), .ZN(n8452) );
  NAND2_X1 U10830 ( .A1(n11427), .A2(n11169), .ZN(n8453) );
  XNOR2_X1 U10831 ( .A(n13050), .B(n10313), .ZN(n8469) );
  NOR2_X1 U10832 ( .A1(P3_D_REG_6__SCAN_IN), .A2(P3_D_REG_14__SCAN_IN), .ZN(
        n8457) );
  NOR4_X1 U10833 ( .A1(P3_D_REG_7__SCAN_IN), .A2(P3_D_REG_8__SCAN_IN), .A3(
        P3_D_REG_2__SCAN_IN), .A4(P3_D_REG_9__SCAN_IN), .ZN(n8456) );
  NOR4_X1 U10834 ( .A1(P3_D_REG_20__SCAN_IN), .A2(P3_D_REG_19__SCAN_IN), .A3(
        P3_D_REG_18__SCAN_IN), .A4(P3_D_REG_27__SCAN_IN), .ZN(n8455) );
  NOR4_X1 U10835 ( .A1(P3_D_REG_30__SCAN_IN), .A2(P3_D_REG_17__SCAN_IN), .A3(
        P3_D_REG_22__SCAN_IN), .A4(P3_D_REG_25__SCAN_IN), .ZN(n8454) );
  NAND4_X1 U10836 ( .A1(n8457), .A2(n8456), .A3(n8455), .A4(n8454), .ZN(n8463)
         );
  NOR4_X1 U10837 ( .A1(P3_D_REG_21__SCAN_IN), .A2(P3_D_REG_12__SCAN_IN), .A3(
        P3_D_REG_11__SCAN_IN), .A4(P3_D_REG_26__SCAN_IN), .ZN(n8461) );
  NOR4_X1 U10838 ( .A1(P3_D_REG_24__SCAN_IN), .A2(P3_D_REG_29__SCAN_IN), .A3(
        P3_D_REG_10__SCAN_IN), .A4(P3_D_REG_31__SCAN_IN), .ZN(n8460) );
  NOR4_X1 U10839 ( .A1(P3_D_REG_23__SCAN_IN), .A2(P3_D_REG_3__SCAN_IN), .A3(
        P3_D_REG_5__SCAN_IN), .A4(P3_D_REG_4__SCAN_IN), .ZN(n8459) );
  NOR4_X1 U10840 ( .A1(P3_D_REG_16__SCAN_IN), .A2(P3_D_REG_15__SCAN_IN), .A3(
        P3_D_REG_13__SCAN_IN), .A4(P3_D_REG_28__SCAN_IN), .ZN(n8458) );
  NAND4_X1 U10841 ( .A1(n8461), .A2(n8460), .A3(n8459), .A4(n8458), .ZN(n8462)
         );
  OAI21_X1 U10842 ( .B1(n8463), .B2(n8462), .A(n9497), .ZN(n8480) );
  NOR2_X1 U10843 ( .A1(n11392), .A2(n11169), .ZN(n8464) );
  NAND2_X1 U10844 ( .A1(n6804), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8467) );
  AND2_X1 U10845 ( .A1(n8480), .A2(n12610), .ZN(n8468) );
  NAND2_X1 U10846 ( .A1(n12585), .A2(n8470), .ZN(n10650) );
  AND2_X1 U10847 ( .A1(n9867), .A2(n10650), .ZN(n10652) );
  OAI22_X1 U10848 ( .A1(n15744), .A2(n8481), .B1(n12706), .B2(n10765), .ZN(
        n8471) );
  AOI21_X1 U10849 ( .B1(n8471), .B2(n12602), .A(n12593), .ZN(n8472) );
  MUX2_X1 U10850 ( .A(n10652), .B(n8472), .S(n8479), .Z(n8473) );
  INV_X1 U10851 ( .A(n15744), .ZN(n15770) );
  INV_X1 U10852 ( .A(n12986), .ZN(n8475) );
  NAND2_X1 U10853 ( .A1(n8477), .A2(n8476), .ZN(P3_U3488) );
  NAND3_X1 U10854 ( .A1(n8479), .A2(n10313), .A3(n8480), .ZN(n9878) );
  INV_X1 U10855 ( .A(n9872), .ZN(n8483) );
  INV_X1 U10856 ( .A(n10313), .ZN(n13052) );
  NAND3_X1 U10857 ( .A1(n13052), .A2(n13050), .A3(n8480), .ZN(n9879) );
  NAND2_X1 U10858 ( .A1(n12593), .A2(n12611), .ZN(n10307) );
  OR2_X1 U10859 ( .A1(n12604), .A2(n8482), .ZN(n9874) );
  AND2_X1 U10860 ( .A1(n10307), .A2(n9874), .ZN(n9865) );
  OAI22_X1 U10861 ( .A1(n9878), .A2(n8483), .B1(n9879), .B2(n9865), .ZN(n8484)
         );
  NAND2_X1 U10862 ( .A1(n15773), .A2(n15770), .ZN(n13049) );
  INV_X1 U10863 ( .A(n13049), .ZN(n8485) );
  NAND2_X1 U10864 ( .A1(n11945), .A2(n8485), .ZN(n8488) );
  OR2_X1 U10865 ( .A1(n15773), .A2(n8486), .ZN(n8487) );
  NOR2_X1 U10866 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), 
        .ZN(n8498) );
  NOR2_X1 U10867 ( .A1(P2_IR_REG_23__SCAN_IN), .A2(P2_IR_REG_22__SCAN_IN), 
        .ZN(n8497) );
  NOR2_X1 U10868 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), 
        .ZN(n8496) );
  NAND2_X1 U10869 ( .A1(n8503), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8504) );
  NAND2_X1 U10870 ( .A1(n9214), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n8509) );
  NAND2_X1 U10871 ( .A1(n6662), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n8508) );
  NAND2_X1 U10872 ( .A1(n9616), .A2(SI_0_), .ZN(n8511) );
  NAND2_X1 U10873 ( .A1(n8511), .A2(n13434), .ZN(n8513) );
  AND2_X1 U10874 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n8512) );
  NAND2_X1 U10875 ( .A1(n9158), .A2(n8512), .ZN(n8533) );
  NAND2_X1 U10876 ( .A1(n8513), .A2(n8533), .ZN(n14039) );
  NAND2_X1 U10877 ( .A1(n8527), .A2(n9268), .ZN(n8515) );
  NAND2_X1 U10878 ( .A1(n8515), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8516) );
  INV_X1 U10879 ( .A(n8517), .ZN(n8518) );
  NAND2_X1 U10880 ( .A1(n8518), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8519) );
  NAND2_X1 U10881 ( .A1(n8527), .A2(n8519), .ZN(n8522) );
  INV_X1 U10882 ( .A(n8522), .ZN(n8521) );
  INV_X1 U10883 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n8520) );
  NAND2_X1 U10884 ( .A1(n8521), .A2(n8520), .ZN(n8524) );
  NAND2_X1 U10885 ( .A1(n8522), .A2(P2_IR_REG_21__SCAN_IN), .ZN(n8523) );
  AND2_X2 U10886 ( .A1(n8524), .A2(n8523), .ZN(n9176) );
  XNOR2_X2 U10887 ( .A(n8526), .B(n8525), .ZN(n9173) );
  XNOR2_X1 U10888 ( .A(n8527), .B(P2_IR_REG_19__SCAN_IN), .ZN(n9175) );
  NAND2_X2 U10889 ( .A1(n9293), .A2(n9175), .ZN(n9241) );
  NAND2_X1 U10890 ( .A1(n9173), .A2(n9175), .ZN(n9673) );
  NAND2_X1 U10891 ( .A1(n13578), .A2(n8528), .ZN(n8530) );
  INV_X1 U10892 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n9362) );
  XNOR2_X1 U10893 ( .A(n8558), .B(SI_1_), .ZN(n8560) );
  AND2_X1 U10894 ( .A1(P2_DATAO_REG_0__SCAN_IN), .A2(SI_0_), .ZN(n8532) );
  NAND2_X1 U10895 ( .A1(n9816), .A2(n8532), .ZN(n9618) );
  NAND2_X1 U10896 ( .A1(n9618), .A2(n8533), .ZN(n8559) );
  XNOR2_X1 U10897 ( .A(n8560), .B(n8559), .ZN(n9818) );
  NAND2_X1 U10898 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), 
        .ZN(n8536) );
  XNOR2_X1 U10899 ( .A(n8536), .B(P2_IR_REG_1__SCAN_IN), .ZN(n9412) );
  INV_X1 U10900 ( .A(n9412), .ZN(n8537) );
  NAND2_X1 U10901 ( .A1(n6672), .A2(n9034), .ZN(n8543) );
  NAND2_X1 U10902 ( .A1(n6662), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n8541) );
  NAND2_X1 U10903 ( .A1(n9214), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n8540) );
  NAND3_X2 U10904 ( .A1(n8541), .A2(n8540), .A3(n8539), .ZN(n13577) );
  NAND2_X1 U10905 ( .A1(n13577), .A2(n8565), .ZN(n8542) );
  NAND2_X1 U10906 ( .A1(n8543), .A2(n8542), .ZN(n8548) );
  NAND2_X1 U10907 ( .A1(n8547), .A2(n8548), .ZN(n8546) );
  AOI22_X1 U10908 ( .A1(n13577), .A2(n9199), .B1(n8565), .B2(n6672), .ZN(n8544) );
  INV_X1 U10909 ( .A(n8544), .ZN(n8545) );
  NAND2_X1 U10910 ( .A1(n8546), .A2(n8545), .ZN(n8552) );
  INV_X1 U10911 ( .A(n8547), .ZN(n8550) );
  INV_X1 U10912 ( .A(n8548), .ZN(n8549) );
  NAND2_X1 U10913 ( .A1(n8550), .A2(n8549), .ZN(n8551) );
  NAND2_X1 U10914 ( .A1(n9214), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n8557) );
  NAND2_X1 U10915 ( .A1(n6662), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n8556) );
  NAND2_X1 U10916 ( .A1(n8571), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n8555) );
  NAND2_X1 U10917 ( .A1(n8553), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n8554) );
  NAND4_X1 U10918 ( .A1(n8557), .A2(n8556), .A3(n8555), .A4(n8554), .ZN(n13576) );
  NAND2_X1 U10919 ( .A1(n13576), .A2(n9034), .ZN(n8567) );
  NAND2_X1 U10920 ( .A1(n8751), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n8564) );
  NOR2_X1 U10921 ( .A1(n8562), .A2(n14018), .ZN(n8561) );
  NAND2_X1 U10922 ( .A1(n8958), .A2(n9432), .ZN(n8563) );
  INV_X1 U10923 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n13095) );
  NAND2_X1 U10924 ( .A1(n9214), .A2(n13095), .ZN(n8575) );
  NAND2_X1 U10925 ( .A1(n6662), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n8574) );
  NAND2_X1 U10926 ( .A1(n8571), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n8573) );
  NAND2_X1 U10927 ( .A1(n8553), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n8572) );
  NAND2_X1 U10928 ( .A1(n13575), .A2(n8565), .ZN(n8584) );
  NAND2_X1 U10929 ( .A1(n8578), .A2(SI_2_), .ZN(n8579) );
  INV_X1 U10930 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n9341) );
  NAND2_X1 U10931 ( .A1(n6772), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8580) );
  MUX2_X1 U10932 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8580), .S(
        P2_IR_REG_3__SCAN_IN), .Z(n8581) );
  AND2_X1 U10933 ( .A1(n8581), .A2(n8620), .ZN(n9448) );
  NAND2_X1 U10934 ( .A1(n8958), .A2(n9448), .ZN(n8582) );
  NAND2_X1 U10935 ( .A1(n13094), .A2(n9034), .ZN(n8583) );
  NAND2_X1 U10936 ( .A1(n8584), .A2(n8583), .ZN(n8586) );
  AOI22_X1 U10937 ( .A1(n13575), .A2(n9199), .B1(n8565), .B2(n13094), .ZN(
        n8585) );
  NAND2_X1 U10938 ( .A1(n8553), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n8593) );
  INV_X1 U10939 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n8588) );
  NAND2_X1 U10940 ( .A1(n13095), .A2(n8588), .ZN(n8589) );
  NAND2_X1 U10941 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n8609) );
  AND2_X1 U10942 ( .A1(n8589), .A2(n8609), .ZN(n10703) );
  NAND2_X1 U10943 ( .A1(n9214), .A2(n10703), .ZN(n8592) );
  NAND2_X1 U10944 ( .A1(n6662), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n8591) );
  NAND2_X1 U10945 ( .A1(n8571), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n8590) );
  NAND4_X1 U10946 ( .A1(n8593), .A2(n8592), .A3(n8591), .A4(n8590), .ZN(n13574) );
  NAND2_X1 U10947 ( .A1(n13574), .A2(n9034), .ZN(n8604) );
  NAND2_X1 U10948 ( .A1(n8620), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8595) );
  INV_X1 U10949 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n8594) );
  XNOR2_X1 U10950 ( .A(n8595), .B(n8594), .ZN(n15419) );
  INV_X1 U10951 ( .A(n8598), .ZN(n8599) );
  NAND2_X1 U10952 ( .A1(n8599), .A2(SI_3_), .ZN(n8600) );
  XNOR2_X1 U10953 ( .A(n8618), .B(SI_4_), .ZN(n8615) );
  XNOR2_X1 U10954 ( .A(n8617), .B(n8615), .ZN(n9342) );
  NAND2_X1 U10955 ( .A1(n9342), .A2(n7114), .ZN(n8602) );
  NAND2_X1 U10956 ( .A1(n8751), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n8601) );
  OAI211_X1 U10957 ( .C1(n8535), .C2(n15419), .A(n8602), .B(n8601), .ZN(n10704) );
  NAND2_X1 U10958 ( .A1(n10704), .A2(n8565), .ZN(n8603) );
  NAND2_X1 U10959 ( .A1(n8604), .A2(n8603), .ZN(n8606) );
  AOI22_X1 U10960 ( .A1(n13574), .A2(n9222), .B1(n9199), .B2(n10704), .ZN(
        n8605) );
  NAND2_X1 U10961 ( .A1(n9191), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n8614) );
  NOR2_X1 U10962 ( .A1(n8609), .A2(n8608), .ZN(n8637) );
  INV_X1 U10963 ( .A(n8637), .ZN(n8639) );
  NAND2_X1 U10964 ( .A1(n8609), .A2(n8608), .ZN(n8610) );
  AND2_X1 U10965 ( .A1(n8639), .A2(n8610), .ZN(n10154) );
  NAND2_X1 U10966 ( .A1(n9214), .A2(n10154), .ZN(n8613) );
  NAND2_X1 U10967 ( .A1(n6662), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n8612) );
  NAND2_X1 U10968 ( .A1(n8571), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n8611) );
  NAND4_X1 U10969 ( .A1(n8614), .A2(n8613), .A3(n8612), .A4(n8611), .ZN(n13573) );
  NAND2_X1 U10970 ( .A1(n13573), .A2(n8565), .ZN(n8626) );
  INV_X1 U10971 ( .A(n8615), .ZN(n8616) );
  NAND2_X1 U10972 ( .A1(n8618), .A2(SI_4_), .ZN(n8619) );
  MUX2_X1 U10973 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(P1_DATAO_REG_5__SCAN_IN), 
        .S(n9616), .Z(n8632) );
  XNOR2_X1 U10974 ( .A(n8632), .B(SI_5_), .ZN(n8629) );
  XNOR2_X1 U10975 ( .A(n8631), .B(n8629), .ZN(n10424) );
  NAND2_X1 U10976 ( .A1(n10424), .A2(n7114), .ZN(n8624) );
  INV_X1 U10977 ( .A(n8620), .ZN(n8621) );
  NAND2_X1 U10978 ( .A1(n8621), .A2(n8594), .ZN(n8685) );
  NAND2_X1 U10979 ( .A1(n8685), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8622) );
  XNOR2_X1 U10980 ( .A(n8622), .B(P2_IR_REG_5__SCAN_IN), .ZN(n9485) );
  AOI22_X1 U10981 ( .A1(n6661), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n8958), .B2(
        n9485), .ZN(n8623) );
  NAND2_X1 U10982 ( .A1(n8624), .A2(n8623), .ZN(n10543) );
  NAND2_X1 U10983 ( .A1(n10543), .A2(n9199), .ZN(n8625) );
  NAND2_X1 U10984 ( .A1(n8626), .A2(n8625), .ZN(n8628) );
  INV_X1 U10985 ( .A(n8629), .ZN(n8630) );
  NAND2_X1 U10986 ( .A1(n8632), .A2(SI_5_), .ZN(n8633) );
  MUX2_X1 U10987 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(P1_DATAO_REG_6__SCAN_IN), 
        .S(n9616), .Z(n8657) );
  XNOR2_X1 U10988 ( .A(n8657), .B(SI_6_), .ZN(n8654) );
  XNOR2_X1 U10989 ( .A(n8656), .B(n8654), .ZN(n10437) );
  NAND2_X1 U10990 ( .A1(n10437), .A2(n7114), .ZN(n8636) );
  OR2_X1 U10991 ( .A1(n8685), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n8658) );
  NAND2_X1 U10992 ( .A1(n8658), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8634) );
  XNOR2_X1 U10993 ( .A(n8634), .B(P2_IR_REG_6__SCAN_IN), .ZN(n9486) );
  AOI22_X1 U10994 ( .A1(n6661), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n8958), .B2(
        n9486), .ZN(n8635) );
  NAND2_X1 U10995 ( .A1(n8553), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n8644) );
  NAND2_X1 U10996 ( .A1(n8637), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n8667) );
  INV_X1 U10997 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n8638) );
  NAND2_X1 U10998 ( .A1(n8639), .A2(n8638), .ZN(n8640) );
  AND2_X1 U10999 ( .A1(n8667), .A2(n8640), .ZN(n10576) );
  NAND2_X1 U11000 ( .A1(n9214), .A2(n10576), .ZN(n8643) );
  NAND2_X1 U11001 ( .A1(n6662), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n8642) );
  NAND2_X1 U11002 ( .A1(n8571), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n8641) );
  NAND4_X1 U11003 ( .A1(n8644), .A2(n8643), .A3(n8642), .A4(n8641), .ZN(n13572) );
  AOI22_X1 U11004 ( .A1(n15513), .A2(n9222), .B1(n9199), .B2(n13572), .ZN(
        n8650) );
  INV_X1 U11005 ( .A(n8650), .ZN(n8645) );
  NAND2_X1 U11006 ( .A1(n8649), .A2(n8645), .ZN(n8648) );
  INV_X1 U11007 ( .A(n13572), .ZN(n9255) );
  NAND2_X1 U11008 ( .A1(n15513), .A2(n9034), .ZN(n8646) );
  OAI21_X1 U11009 ( .B1(n9255), .B2(n9241), .A(n8646), .ZN(n8647) );
  NAND2_X1 U11010 ( .A1(n8648), .A2(n8647), .ZN(n8653) );
  INV_X1 U11011 ( .A(n8649), .ZN(n8651) );
  NAND2_X1 U11012 ( .A1(n8651), .A2(n8650), .ZN(n8652) );
  INV_X1 U11013 ( .A(n8654), .ZN(n8655) );
  MUX2_X1 U11014 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(P1_DATAO_REG_7__SCAN_IN), 
        .S(n9616), .Z(n8680) );
  XNOR2_X1 U11015 ( .A(n8680), .B(SI_7_), .ZN(n8677) );
  XNOR2_X1 U11016 ( .A(n7174), .B(n8677), .ZN(n10736) );
  NAND2_X1 U11017 ( .A1(n10736), .A2(n7114), .ZN(n8665) );
  INV_X1 U11018 ( .A(n8658), .ZN(n8660) );
  INV_X1 U11019 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n8659) );
  NAND2_X1 U11020 ( .A1(n8660), .A2(n8659), .ZN(n8662) );
  NAND2_X1 U11021 ( .A1(n8662), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8661) );
  MUX2_X1 U11022 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8661), .S(
        P2_IR_REG_7__SCAN_IN), .Z(n8663) );
  AOI22_X1 U11023 ( .A1(n6661), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n8958), .B2(
        n13589), .ZN(n8664) );
  NAND2_X1 U11024 ( .A1(n8665), .A2(n8664), .ZN(n10794) );
  NAND2_X1 U11025 ( .A1(n9191), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n8672) );
  INV_X1 U11026 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n8666) );
  NAND2_X1 U11027 ( .A1(n8667), .A2(n8666), .ZN(n8668) );
  AND2_X1 U11028 ( .A1(n8709), .A2(n8668), .ZN(n10537) );
  NAND2_X1 U11029 ( .A1(n9214), .A2(n10537), .ZN(n8671) );
  NAND2_X1 U11030 ( .A1(n6662), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n8670) );
  NAND2_X1 U11031 ( .A1(n8571), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n8669) );
  NAND4_X1 U11032 ( .A1(n8672), .A2(n8671), .A3(n8670), .A4(n8669), .ZN(n13571) );
  AND2_X1 U11033 ( .A1(n13571), .A2(n8565), .ZN(n8673) );
  AOI21_X1 U11034 ( .B1(n10794), .B2(n9199), .A(n8673), .ZN(n8674) );
  INV_X1 U11035 ( .A(n13571), .ZN(n10793) );
  NAND2_X1 U11036 ( .A1(n10794), .A2(n8565), .ZN(n8675) );
  OAI21_X1 U11037 ( .B1(n9222), .B2(n10793), .A(n8675), .ZN(n8676) );
  INV_X1 U11038 ( .A(n8677), .ZN(n8678) );
  MUX2_X1 U11039 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(P1_DATAO_REG_8__SCAN_IN), 
        .S(n9616), .Z(n8698) );
  NAND2_X1 U11040 ( .A1(n10828), .A2(n7114), .ZN(n8688) );
  NAND2_X1 U11041 ( .A1(n8681), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8682) );
  MUX2_X1 U11042 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8682), .S(
        P2_IR_REG_8__SCAN_IN), .Z(n8686) );
  INV_X1 U11043 ( .A(n8683), .ZN(n8684) );
  NAND2_X1 U11044 ( .A1(n8686), .A2(n8701), .ZN(n9489) );
  INV_X1 U11045 ( .A(n9489), .ZN(n9535) );
  AOI22_X1 U11046 ( .A1(n6661), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n8958), .B2(
        n9535), .ZN(n8687) );
  NAND2_X1 U11047 ( .A1(n15530), .A2(n8565), .ZN(n8694) );
  NAND2_X1 U11048 ( .A1(n9191), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n8692) );
  XNOR2_X1 U11049 ( .A(n8709), .B(P2_REG3_REG_8__SCAN_IN), .ZN(n10894) );
  NAND2_X1 U11050 ( .A1(n9214), .A2(n10894), .ZN(n8691) );
  NAND2_X1 U11051 ( .A1(n6662), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n8690) );
  NAND2_X1 U11052 ( .A1(n8571), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n8689) );
  NAND4_X1 U11053 ( .A1(n8692), .A2(n8691), .A3(n8690), .A4(n8689), .ZN(n13570) );
  NAND2_X1 U11054 ( .A1(n13570), .A2(n9034), .ZN(n8693) );
  NAND2_X1 U11055 ( .A1(n8694), .A2(n8693), .ZN(n8696) );
  AOI22_X1 U11056 ( .A1(n15530), .A2(n9034), .B1(n9222), .B2(n13570), .ZN(
        n8695) );
  MUX2_X1 U11057 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(P1_DATAO_REG_9__SCAN_IN), 
        .S(n9616), .Z(n8725) );
  XNOR2_X1 U11058 ( .A(n8725), .B(SI_9_), .ZN(n8722) );
  XNOR2_X1 U11059 ( .A(n8724), .B(n8722), .ZN(n11065) );
  NAND2_X1 U11060 ( .A1(n11065), .A2(n7114), .ZN(n8705) );
  NAND2_X1 U11061 ( .A1(n8701), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8700) );
  MUX2_X1 U11062 ( .A(n8700), .B(P2_IR_REG_31__SCAN_IN), .S(n8699), .Z(n8703)
         );
  INV_X1 U11063 ( .A(n8701), .ZN(n8702) );
  NAND2_X1 U11064 ( .A1(n8702), .A2(n8699), .ZN(n8749) );
  NAND2_X1 U11065 ( .A1(n8703), .A2(n8749), .ZN(n9537) );
  INV_X1 U11066 ( .A(n9537), .ZN(n13605) );
  AOI22_X1 U11067 ( .A1(n6661), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n8958), .B2(
        n13605), .ZN(n8704) );
  NAND2_X1 U11068 ( .A1(n15538), .A2(n9034), .ZN(n8716) );
  NAND2_X1 U11069 ( .A1(n6662), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n8714) );
  NAND2_X1 U11070 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_REG3_REG_8__SCAN_IN), 
        .ZN(n8706) );
  INV_X1 U11071 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n8708) );
  INV_X1 U11072 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n8707) );
  OAI21_X1 U11073 ( .B1(n8709), .B2(n8708), .A(n8707), .ZN(n8710) );
  AND2_X1 U11074 ( .A1(n8730), .A2(n8710), .ZN(n10819) );
  NAND2_X1 U11075 ( .A1(n9214), .A2(n10819), .ZN(n8713) );
  NAND2_X1 U11076 ( .A1(n9191), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n8712) );
  NAND2_X1 U11077 ( .A1(n8571), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n8711) );
  NAND4_X1 U11078 ( .A1(n8714), .A2(n8713), .A3(n8712), .A4(n8711), .ZN(n13569) );
  NAND2_X1 U11079 ( .A1(n13569), .A2(n8565), .ZN(n8715) );
  NAND2_X1 U11080 ( .A1(n8716), .A2(n8715), .ZN(n8719) );
  INV_X1 U11081 ( .A(n13569), .ZN(n10988) );
  NAND2_X1 U11082 ( .A1(n15538), .A2(n8565), .ZN(n8717) );
  OAI21_X1 U11083 ( .B1(n9222), .B2(n10988), .A(n8717), .ZN(n8718) );
  INV_X1 U11084 ( .A(n8719), .ZN(n8720) );
  INV_X1 U11085 ( .A(n8722), .ZN(n8723) );
  NAND2_X1 U11086 ( .A1(n8725), .A2(SI_9_), .ZN(n8726) );
  MUX2_X1 U11087 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(P1_DATAO_REG_10__SCAN_IN), 
        .S(n9616), .Z(n8744) );
  XNOR2_X1 U11088 ( .A(n8744), .B(SI_10_), .ZN(n8741) );
  XNOR2_X1 U11089 ( .A(n8743), .B(n8741), .ZN(n11071) );
  NAND2_X1 U11090 ( .A1(n11071), .A2(n7114), .ZN(n8729) );
  NAND2_X1 U11091 ( .A1(n8749), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8727) );
  XNOR2_X1 U11092 ( .A(n8727), .B(P2_IR_REG_10__SCAN_IN), .ZN(n9567) );
  AOI22_X1 U11093 ( .A1(n6660), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n8958), 
        .B2(n9567), .ZN(n8728) );
  NAND2_X2 U11094 ( .A1(n8729), .A2(n8728), .ZN(n11229) );
  NAND2_X1 U11095 ( .A1(n11229), .A2(n8565), .ZN(n8737) );
  NAND2_X1 U11096 ( .A1(n6662), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n8735) );
  INV_X1 U11097 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n13266) );
  INV_X1 U11098 ( .A(n8786), .ZN(n8784) );
  NAND2_X1 U11099 ( .A1(n8730), .A2(n13266), .ZN(n8731) );
  AND2_X1 U11100 ( .A1(n8784), .A2(n8731), .ZN(n10994) );
  NAND2_X1 U11101 ( .A1(n9214), .A2(n10994), .ZN(n8734) );
  NAND2_X1 U11102 ( .A1(n9191), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n8733) );
  NAND2_X1 U11103 ( .A1(n8571), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n8732) );
  NAND4_X1 U11104 ( .A1(n8735), .A2(n8734), .A3(n8733), .A4(n8732), .ZN(n13568) );
  NAND2_X1 U11105 ( .A1(n13568), .A2(n9199), .ZN(n8736) );
  NAND2_X1 U11106 ( .A1(n8737), .A2(n8736), .ZN(n8739) );
  AOI22_X1 U11107 ( .A1(n11229), .A2(n9034), .B1(n9222), .B2(n13568), .ZN(
        n8738) );
  INV_X1 U11108 ( .A(n8741), .ZN(n8742) );
  MUX2_X1 U11109 ( .A(n9553), .B(n9548), .S(n9616), .Z(n8746) );
  NAND2_X1 U11110 ( .A1(n8746), .A2(n8745), .ZN(n8771) );
  INV_X1 U11111 ( .A(n8746), .ZN(n8747) );
  NAND2_X1 U11112 ( .A1(n8747), .A2(SI_11_), .ZN(n8748) );
  NAND2_X1 U11113 ( .A1(n8771), .A2(n8748), .ZN(n8769) );
  XNOR2_X1 U11114 ( .A(n8770), .B(n8769), .ZN(n11281) );
  NAND2_X1 U11115 ( .A1(n11281), .A2(n7114), .ZN(n8753) );
  OAI21_X1 U11116 ( .B1(n8749), .B2(P2_IR_REG_10__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8750) );
  XNOR2_X1 U11117 ( .A(n8750), .B(P2_IR_REG_11__SCAN_IN), .ZN(n9568) );
  AOI22_X1 U11118 ( .A1(n6661), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n8958), 
        .B2(n9568), .ZN(n8752) );
  NAND2_X1 U11119 ( .A1(n11323), .A2(n9199), .ZN(n8759) );
  NAND2_X1 U11120 ( .A1(n6662), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n8757) );
  XNOR2_X1 U11121 ( .A(n8784), .B(P2_REG3_REG_11__SCAN_IN), .ZN(n11393) );
  NAND2_X1 U11122 ( .A1(n9214), .A2(n11393), .ZN(n8756) );
  NAND2_X1 U11123 ( .A1(n8571), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n8755) );
  NAND2_X1 U11124 ( .A1(n9191), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n8754) );
  NAND4_X1 U11125 ( .A1(n8757), .A2(n8756), .A3(n8755), .A4(n8754), .ZN(n13567) );
  NAND2_X1 U11126 ( .A1(n13567), .A2(n9222), .ZN(n8758) );
  NAND2_X1 U11127 ( .A1(n8759), .A2(n8758), .ZN(n8764) );
  INV_X1 U11128 ( .A(n13567), .ZN(n11324) );
  NAND2_X1 U11129 ( .A1(n11323), .A2(n9222), .ZN(n8760) );
  OAI21_X1 U11130 ( .B1(n8565), .B2(n11324), .A(n8760), .ZN(n8761) );
  NAND2_X1 U11131 ( .A1(n8762), .A2(n8761), .ZN(n8768) );
  INV_X1 U11132 ( .A(n8763), .ZN(n8766) );
  INV_X1 U11133 ( .A(n8764), .ZN(n8765) );
  NAND2_X1 U11134 ( .A1(n8766), .A2(n8765), .ZN(n8767) );
  MUX2_X1 U11135 ( .A(n9691), .B(n9594), .S(n9616), .Z(n8772) );
  NAND2_X1 U11136 ( .A1(n8772), .A2(n9367), .ZN(n8797) );
  INV_X1 U11137 ( .A(n8772), .ZN(n8773) );
  NAND2_X1 U11138 ( .A1(n8773), .A2(SI_12_), .ZN(n8774) );
  XNOR2_X1 U11139 ( .A(n8796), .B(n7913), .ZN(n11287) );
  NAND2_X1 U11140 ( .A1(n11287), .A2(n7114), .ZN(n8781) );
  NAND2_X1 U11141 ( .A1(n8775), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8776) );
  MUX2_X1 U11142 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8776), .S(
        P2_IR_REG_12__SCAN_IN), .Z(n8777) );
  INV_X1 U11143 ( .A(n8777), .ZN(n8779) );
  NOR2_X1 U11144 ( .A1(n8779), .A2(n8778), .ZN(n10178) );
  AOI22_X1 U11145 ( .A1(n6660), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n8958), 
        .B2(n10178), .ZN(n8780) );
  NAND2_X1 U11146 ( .A1(n15140), .A2(n9222), .ZN(n8793) );
  NAND2_X1 U11147 ( .A1(n8553), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n8791) );
  INV_X1 U11148 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n8783) );
  INV_X1 U11149 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n8782) );
  OAI21_X1 U11150 ( .B1(n8784), .B2(n8783), .A(n8782), .ZN(n8787) );
  AND2_X1 U11151 ( .A1(P2_REG3_REG_11__SCAN_IN), .A2(P2_REG3_REG_12__SCAN_IN), 
        .ZN(n8785) );
  INV_X1 U11152 ( .A(n8804), .ZN(n8805) );
  AND2_X1 U11153 ( .A1(n8787), .A2(n8805), .ZN(n15138) );
  NAND2_X1 U11154 ( .A1(n9214), .A2(n15138), .ZN(n8790) );
  NAND2_X1 U11155 ( .A1(n6662), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n8789) );
  NAND2_X1 U11156 ( .A1(n8571), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n8788) );
  NAND4_X1 U11157 ( .A1(n8791), .A2(n8790), .A3(n8789), .A4(n8788), .ZN(n13566) );
  NAND2_X1 U11158 ( .A1(n13566), .A2(n9199), .ZN(n8792) );
  NAND2_X1 U11159 ( .A1(n8793), .A2(n8792), .ZN(n8795) );
  AOI22_X1 U11160 ( .A1(n15140), .A2(n9034), .B1(n9222), .B2(n13566), .ZN(
        n8794) );
  MUX2_X1 U11161 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(P1_DATAO_REG_13__SCAN_IN), 
        .S(n9616), .Z(n8819) );
  XNOR2_X1 U11162 ( .A(n8819), .B(n14929), .ZN(n8816) );
  XNOR2_X1 U11163 ( .A(n8818), .B(n8816), .ZN(n11445) );
  NAND2_X1 U11164 ( .A1(n11445), .A2(n7114), .ZN(n8803) );
  INV_X1 U11165 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n14018) );
  NOR2_X1 U11166 ( .A1(n8778), .A2(n14018), .ZN(n8798) );
  MUX2_X1 U11167 ( .A(n14018), .B(n8798), .S(P2_IR_REG_13__SCAN_IN), .Z(n8799)
         );
  INV_X1 U11168 ( .A(n8799), .ZN(n8801) );
  NAND2_X1 U11169 ( .A1(n8778), .A2(n8800), .ZN(n8825) );
  AND2_X1 U11170 ( .A1(n8801), .A2(n8825), .ZN(n15454) );
  AOI22_X1 U11171 ( .A1(n6661), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n8958), 
        .B2(n15454), .ZN(n8802) );
  NAND2_X1 U11172 ( .A1(n11491), .A2(n9199), .ZN(n8812) );
  NAND2_X1 U11173 ( .A1(n9191), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n8810) );
  NAND2_X1 U11174 ( .A1(n8804), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n8830) );
  INV_X1 U11175 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n15451) );
  NAND2_X1 U11176 ( .A1(n8805), .A2(n15451), .ZN(n8806) );
  AND2_X1 U11177 ( .A1(n8830), .A2(n8806), .ZN(n11330) );
  NAND2_X1 U11178 ( .A1(n9214), .A2(n11330), .ZN(n8809) );
  NAND2_X1 U11179 ( .A1(n6662), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n8808) );
  NAND2_X1 U11180 ( .A1(n8571), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n8807) );
  NAND4_X1 U11181 ( .A1(n8810), .A2(n8809), .A3(n8808), .A4(n8807), .ZN(n13565) );
  NAND2_X1 U11182 ( .A1(n13565), .A2(n9222), .ZN(n8811) );
  NAND2_X1 U11183 ( .A1(n8812), .A2(n8811), .ZN(n8815) );
  INV_X1 U11184 ( .A(n13565), .ZN(n11495) );
  NAND2_X1 U11185 ( .A1(n11491), .A2(n9222), .ZN(n8813) );
  OAI21_X1 U11186 ( .B1(n9222), .B2(n11495), .A(n8813), .ZN(n8814) );
  INV_X1 U11187 ( .A(n8816), .ZN(n8817) );
  NAND2_X1 U11188 ( .A1(n8819), .A2(SI_13_), .ZN(n8820) );
  MUX2_X1 U11189 ( .A(n9813), .B(n9815), .S(n9616), .Z(n8821) );
  INV_X1 U11190 ( .A(n8821), .ZN(n8822) );
  NAND2_X1 U11191 ( .A1(n8822), .A2(SI_14_), .ZN(n8823) );
  NAND2_X1 U11192 ( .A1(n8847), .A2(n8823), .ZN(n8845) );
  XNOR2_X1 U11193 ( .A(n8846), .B(n8845), .ZN(n11450) );
  NAND2_X1 U11194 ( .A1(n11450), .A2(n7114), .ZN(n8828) );
  NAND2_X1 U11195 ( .A1(n8825), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8824) );
  MUX2_X1 U11196 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8824), .S(
        P2_IR_REG_14__SCAN_IN), .Z(n8826) );
  AOI22_X1 U11197 ( .A1(n6661), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n8958), 
        .B2(n10865), .ZN(n8827) );
  NAND2_X1 U11198 ( .A1(n15127), .A2(n9222), .ZN(n8838) );
  NAND2_X1 U11199 ( .A1(n6662), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n8836) );
  INV_X1 U11200 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n8829) );
  NAND2_X1 U11201 ( .A1(n8830), .A2(n8829), .ZN(n8831) );
  NAND2_X1 U11202 ( .A1(n8858), .A2(n8831), .ZN(n15132) );
  INV_X1 U11203 ( .A(n15132), .ZN(n8832) );
  NAND2_X1 U11204 ( .A1(n9214), .A2(n8832), .ZN(n8835) );
  NAND2_X1 U11205 ( .A1(n8571), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n8834) );
  NAND2_X1 U11206 ( .A1(n9191), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n8833) );
  NAND4_X1 U11207 ( .A1(n8836), .A2(n8835), .A3(n8834), .A4(n8833), .ZN(n13564) );
  NAND2_X1 U11208 ( .A1(n13564), .A2(n9199), .ZN(n8837) );
  NAND2_X1 U11209 ( .A1(n8838), .A2(n8837), .ZN(n8843) );
  NAND2_X1 U11210 ( .A1(n8842), .A2(n8843), .ZN(n8841) );
  INV_X1 U11211 ( .A(n13564), .ZN(n9252) );
  NAND2_X1 U11212 ( .A1(n15127), .A2(n9199), .ZN(n8839) );
  OAI21_X1 U11213 ( .B1(n9252), .B2(n9241), .A(n8839), .ZN(n8840) );
  INV_X1 U11214 ( .A(n8842), .ZN(n8844) );
  MUX2_X1 U11215 ( .A(n10054), .B(n9971), .S(n9616), .Z(n8848) );
  INV_X1 U11216 ( .A(n8848), .ZN(n8849) );
  NAND2_X1 U11217 ( .A1(n8849), .A2(SI_15_), .ZN(n8850) );
  XNOR2_X1 U11218 ( .A(n8868), .B(n8867), .ZN(n11613) );
  NAND2_X1 U11219 ( .A1(n11613), .A2(n7114), .ZN(n8856) );
  NAND2_X1 U11220 ( .A1(n8853), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8852) );
  MUX2_X1 U11221 ( .A(n8852), .B(P2_IR_REG_31__SCAN_IN), .S(n8851), .Z(n8854)
         );
  NAND2_X1 U11222 ( .A1(n8854), .A2(n8895), .ZN(n15478) );
  INV_X1 U11223 ( .A(n15478), .ZN(n10879) );
  AOI22_X1 U11224 ( .A1(n6661), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n8958), 
        .B2(n10879), .ZN(n8855) );
  INV_X1 U11225 ( .A(n8882), .ZN(n8900) );
  NAND2_X1 U11226 ( .A1(n8858), .A2(n8857), .ZN(n8859) );
  AND2_X1 U11227 ( .A1(n8900), .A2(n8859), .ZN(n11925) );
  NAND2_X1 U11228 ( .A1(n9214), .A2(n11925), .ZN(n8863) );
  NAND2_X1 U11229 ( .A1(n6662), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n8862) );
  NAND2_X1 U11230 ( .A1(n8571), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n8861) );
  NAND2_X1 U11231 ( .A1(n9191), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n8860) );
  NAND4_X1 U11232 ( .A1(n8863), .A2(n8862), .A3(n8861), .A4(n8860), .ZN(n13643) );
  AND2_X1 U11233 ( .A1(n13643), .A2(n9199), .ZN(n8864) );
  AOI21_X1 U11234 ( .B1(n13991), .B2(n9222), .A(n8864), .ZN(n8917) );
  NAND2_X1 U11235 ( .A1(n13991), .A2(n9199), .ZN(n8866) );
  NAND2_X1 U11236 ( .A1(n13643), .A2(n9222), .ZN(n8865) );
  NAND2_X1 U11237 ( .A1(n8866), .A2(n8865), .ZN(n8916) );
  MUX2_X1 U11238 ( .A(n10234), .B(n10153), .S(n9616), .Z(n8871) );
  INV_X1 U11239 ( .A(n8871), .ZN(n8872) );
  NAND2_X1 U11240 ( .A1(n8872), .A2(SI_16_), .ZN(n8873) );
  MUX2_X1 U11241 ( .A(n10414), .B(n7532), .S(n9616), .Z(n8876) );
  INV_X1 U11242 ( .A(n8876), .ZN(n8877) );
  NAND2_X1 U11243 ( .A1(n8877), .A2(SI_17_), .ZN(n8878) );
  XNOR2_X1 U11244 ( .A(n8930), .B(n8929), .ZN(n11637) );
  NAND2_X1 U11245 ( .A1(n11637), .A2(n7114), .ZN(n8881) );
  OAI21_X1 U11246 ( .B1(n8895), .B2(P2_IR_REG_16__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8879) );
  XNOR2_X1 U11247 ( .A(n8879), .B(P2_IR_REG_17__SCAN_IN), .ZN(n11111) );
  AOI22_X1 U11248 ( .A1(n6660), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n8958), 
        .B2(n11111), .ZN(n8880) );
  NAND2_X1 U11249 ( .A1(n6662), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n8889) );
  INV_X1 U11250 ( .A(n8883), .ZN(n8902) );
  INV_X1 U11251 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n8884) );
  NAND2_X1 U11252 ( .A1(n8902), .A2(n8884), .ZN(n8885) );
  AND2_X1 U11253 ( .A1(n8937), .A2(n8885), .ZN(n13864) );
  NAND2_X1 U11254 ( .A1(n9214), .A2(n13864), .ZN(n8888) );
  NAND2_X1 U11255 ( .A1(n9191), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n8887) );
  NAND2_X1 U11256 ( .A1(n8571), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n8886) );
  NAND4_X1 U11257 ( .A1(n8889), .A2(n8888), .A3(n8887), .A4(n8886), .ZN(n13672) );
  AND2_X1 U11258 ( .A1(n13672), .A2(n8565), .ZN(n8890) );
  AOI21_X1 U11259 ( .B1(n13673), .B2(n9199), .A(n8890), .ZN(n8927) );
  NAND2_X1 U11260 ( .A1(n13673), .A2(n9222), .ZN(n8892) );
  NAND2_X1 U11261 ( .A1(n13672), .A2(n9199), .ZN(n8891) );
  NAND2_X1 U11262 ( .A1(n8892), .A2(n8891), .ZN(n8921) );
  XNOR2_X1 U11263 ( .A(n8894), .B(n8893), .ZN(n11620) );
  NAND2_X1 U11264 ( .A1(n11620), .A2(n7114), .ZN(n8898) );
  NAND2_X1 U11265 ( .A1(n8895), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8896) );
  XNOR2_X1 U11266 ( .A(n8896), .B(P2_IR_REG_16__SCAN_IN), .ZN(n10870) );
  AOI22_X1 U11267 ( .A1(n6661), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n8958), 
        .B2(n10870), .ZN(n8897) );
  NAND2_X1 U11268 ( .A1(n6662), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n8906) );
  INV_X1 U11269 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n8899) );
  NAND2_X1 U11270 ( .A1(n8900), .A2(n8899), .ZN(n8901) );
  AND2_X1 U11271 ( .A1(n8902), .A2(n8901), .ZN(n13887) );
  NAND2_X1 U11272 ( .A1(n9214), .A2(n13887), .ZN(n8905) );
  NAND2_X1 U11273 ( .A1(n8571), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n8904) );
  NAND2_X1 U11274 ( .A1(n8553), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n8903) );
  NAND4_X1 U11275 ( .A1(n8906), .A2(n8905), .A3(n8904), .A4(n8903), .ZN(n13670) );
  AND2_X1 U11276 ( .A1(n13670), .A2(n8565), .ZN(n8907) );
  AOI21_X1 U11277 ( .B1(n13985), .B2(n9199), .A(n8907), .ZN(n8912) );
  NAND2_X1 U11278 ( .A1(n13985), .A2(n9222), .ZN(n8909) );
  NAND2_X1 U11279 ( .A1(n13670), .A2(n9199), .ZN(n8908) );
  NAND2_X1 U11280 ( .A1(n8909), .A2(n8908), .ZN(n8911) );
  AOI22_X1 U11281 ( .A1(n8927), .A2(n8921), .B1(n8912), .B2(n8911), .ZN(n8915)
         );
  OAI21_X1 U11282 ( .B1(n8917), .B2(n8916), .A(n8915), .ZN(n8910) );
  INV_X1 U11283 ( .A(n8911), .ZN(n8914) );
  INV_X1 U11284 ( .A(n8912), .ZN(n8913) );
  AND2_X1 U11285 ( .A1(n8914), .A2(n8913), .ZN(n8923) );
  INV_X1 U11286 ( .A(n8923), .ZN(n8926) );
  INV_X1 U11287 ( .A(n8915), .ZN(n8920) );
  INV_X1 U11288 ( .A(n8916), .ZN(n8919) );
  INV_X1 U11289 ( .A(n8917), .ZN(n8918) );
  OR3_X1 U11290 ( .A1(n8920), .A2(n8919), .A3(n8918), .ZN(n8925) );
  OR2_X1 U11291 ( .A1(n13673), .A2(n13672), .ZN(n13648) );
  INV_X1 U11292 ( .A(n8921), .ZN(n8922) );
  OAI21_X1 U11293 ( .B1(n8923), .B2(n13648), .A(n8922), .ZN(n8924) );
  OAI211_X1 U11294 ( .C1(n8927), .C2(n8926), .A(n8925), .B(n8924), .ZN(n8928)
         );
  XNOR2_X1 U11295 ( .A(n8978), .B(SI_18_), .ZN(n8950) );
  MUX2_X1 U11296 ( .A(n10721), .B(n10735), .S(n9616), .Z(n8974) );
  XNOR2_X1 U11297 ( .A(n8950), .B(n8974), .ZN(n11561) );
  NAND2_X1 U11298 ( .A1(n11561), .A2(n7114), .ZN(n8935) );
  NAND2_X1 U11299 ( .A1(n8932), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8933) );
  XNOR2_X1 U11300 ( .A(n8933), .B(P2_IR_REG_18__SCAN_IN), .ZN(n13618) );
  AOI22_X1 U11301 ( .A1(n6661), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n8958), 
        .B2(n13618), .ZN(n8934) );
  INV_X1 U11302 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n8936) );
  NAND2_X1 U11303 ( .A1(n8937), .A2(n8936), .ZN(n8938) );
  AND2_X1 U11304 ( .A1(n8963), .A2(n8938), .ZN(n13846) );
  NAND2_X1 U11305 ( .A1(n13846), .A2(n9214), .ZN(n8942) );
  NAND2_X1 U11306 ( .A1(n9191), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n8941) );
  NAND2_X1 U11307 ( .A1(n6662), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n8940) );
  NAND2_X1 U11308 ( .A1(n8571), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n8939) );
  NAND4_X1 U11309 ( .A1(n8942), .A2(n8941), .A3(n8940), .A4(n8939), .ZN(n13675) );
  AND2_X1 U11310 ( .A1(n13675), .A2(n9199), .ZN(n8943) );
  AOI21_X1 U11311 ( .B1(n13845), .B2(n9222), .A(n8943), .ZN(n8946) );
  INV_X1 U11312 ( .A(n13675), .ZN(n13676) );
  NAND2_X1 U11313 ( .A1(n13845), .A2(n9199), .ZN(n8944) );
  OAI21_X1 U11314 ( .B1(n13676), .B2(n9241), .A(n8944), .ZN(n8945) );
  NAND2_X1 U11315 ( .A1(n8947), .A2(n8946), .ZN(n8948) );
  NAND2_X1 U11316 ( .A1(n8950), .A2(n8974), .ZN(n8952) );
  NAND2_X1 U11317 ( .A1(n8978), .A2(n8973), .ZN(n8951) );
  NAND2_X1 U11318 ( .A1(n8952), .A2(n8951), .ZN(n8957) );
  MUX2_X1 U11319 ( .A(n10770), .B(n13423), .S(n9616), .Z(n8953) );
  INV_X1 U11320 ( .A(SI_19_), .ZN(n10082) );
  NAND2_X1 U11321 ( .A1(n8953), .A2(n10082), .ZN(n8979) );
  INV_X1 U11322 ( .A(n8953), .ZN(n8954) );
  NAND2_X1 U11323 ( .A1(n8954), .A2(SI_19_), .ZN(n8955) );
  NAND2_X1 U11324 ( .A1(n8979), .A2(n8955), .ZN(n8976) );
  INV_X1 U11325 ( .A(n8976), .ZN(n8956) );
  NAND2_X1 U11326 ( .A1(n11656), .A2(n7114), .ZN(n8960) );
  AOI22_X1 U11327 ( .A1(n6661), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n9175), 
        .B2(n8958), .ZN(n8959) );
  NAND2_X1 U11328 ( .A1(n13965), .A2(n9199), .ZN(n8969) );
  INV_X1 U11329 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n8967) );
  INV_X1 U11330 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n8962) );
  NAND2_X1 U11331 ( .A1(n8963), .A2(n8962), .ZN(n8964) );
  NAND2_X1 U11332 ( .A1(n8982), .A2(n8964), .ZN(n13831) );
  OR2_X1 U11333 ( .A1(n13831), .A2(n9198), .ZN(n8966) );
  AOI22_X1 U11334 ( .A1(n6662), .A2(P2_REG1_REG_19__SCAN_IN), .B1(n9191), .B2(
        P2_REG2_REG_19__SCAN_IN), .ZN(n8965) );
  OAI211_X1 U11335 ( .C1(n9217), .C2(n8967), .A(n8966), .B(n8965), .ZN(n13679)
         );
  NAND2_X1 U11336 ( .A1(n13679), .A2(n9222), .ZN(n8968) );
  NAND2_X1 U11337 ( .A1(n8969), .A2(n8968), .ZN(n8971) );
  AOI22_X1 U11338 ( .A1(n13965), .A2(n8565), .B1(n9199), .B2(n13679), .ZN(
        n8970) );
  INV_X1 U11339 ( .A(n8974), .ZN(n8972) );
  NOR2_X1 U11340 ( .A1(n8974), .A2(n8973), .ZN(n8975) );
  NOR2_X1 U11341 ( .A1(n8976), .A2(n8975), .ZN(n8977) );
  INV_X1 U11342 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n10888) );
  MUX2_X1 U11343 ( .A(n10888), .B(n11860), .S(n9616), .Z(n8993) );
  XNOR2_X1 U11344 ( .A(n8995), .B(n8993), .ZN(n11674) );
  NAND2_X1 U11345 ( .A1(n11674), .A2(n7114), .ZN(n8981) );
  NAND2_X1 U11346 ( .A1(n6661), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n8980) );
  NAND2_X1 U11347 ( .A1(n13681), .A2(n9222), .ZN(n8988) );
  INV_X1 U11348 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n8986) );
  NAND2_X1 U11349 ( .A1(n8982), .A2(n13537), .ZN(n8983) );
  NAND2_X1 U11350 ( .A1(n9001), .A2(n8983), .ZN(n13823) );
  OR2_X1 U11351 ( .A1(n13823), .A2(n9198), .ZN(n8985) );
  AOI22_X1 U11352 ( .A1(n6662), .A2(P2_REG1_REG_20__SCAN_IN), .B1(n9191), .B2(
        P2_REG2_REG_20__SCAN_IN), .ZN(n8984) );
  OAI211_X1 U11353 ( .C1(n9217), .C2(n8986), .A(n8985), .B(n8984), .ZN(n13680)
         );
  NAND2_X1 U11354 ( .A1(n13680), .A2(n9199), .ZN(n8987) );
  NAND2_X1 U11355 ( .A1(n8988), .A2(n8987), .ZN(n8990) );
  AOI22_X1 U11356 ( .A1(n13681), .A2(n9199), .B1(n9222), .B2(n13680), .ZN(
        n8989) );
  AOI21_X1 U11357 ( .B1(n8991), .B2(n8990), .A(n8989), .ZN(n8992) );
  INV_X1 U11358 ( .A(n8993), .ZN(n8994) );
  MUX2_X1 U11359 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(P1_DATAO_REG_21__SCAN_IN), 
        .S(n9616), .Z(n9017) );
  XNOR2_X1 U11360 ( .A(n9017), .B(SI_21_), .ZN(n9014) );
  XNOR2_X1 U11361 ( .A(n9016), .B(n9014), .ZN(n11696) );
  NAND2_X1 U11362 ( .A1(n11696), .A2(n7114), .ZN(n9000) );
  NAND2_X1 U11363 ( .A1(n6660), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n8999) );
  NAND2_X1 U11364 ( .A1(n13953), .A2(n9034), .ZN(n9010) );
  NAND2_X1 U11365 ( .A1(n9001), .A2(n13119), .ZN(n9002) );
  AND2_X1 U11366 ( .A1(n9024), .A2(n9002), .ZN(n13812) );
  NAND2_X1 U11367 ( .A1(n13812), .A2(n9214), .ZN(n9008) );
  INV_X1 U11368 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n9005) );
  NAND2_X1 U11369 ( .A1(n8571), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n9004) );
  NAND2_X1 U11370 ( .A1(n9191), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n9003) );
  OAI211_X1 U11371 ( .C1(n9195), .C2(n9005), .A(n9004), .B(n9003), .ZN(n9006)
         );
  INV_X1 U11372 ( .A(n9006), .ZN(n9007) );
  NAND2_X1 U11373 ( .A1(n9008), .A2(n9007), .ZN(n13684) );
  NAND2_X1 U11374 ( .A1(n13684), .A2(n9222), .ZN(n9009) );
  NAND2_X1 U11375 ( .A1(n9010), .A2(n9009), .ZN(n9013) );
  INV_X1 U11376 ( .A(n13684), .ZN(n11912) );
  NAND2_X1 U11377 ( .A1(n13953), .A2(n9222), .ZN(n9011) );
  OAI21_X1 U11378 ( .B1(n9222), .B2(n11912), .A(n9011), .ZN(n9012) );
  INV_X1 U11379 ( .A(n9014), .ZN(n9015) );
  NAND2_X1 U11380 ( .A1(n9017), .A2(SI_21_), .ZN(n9018) );
  MUX2_X1 U11381 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(P1_DATAO_REG_22__SCAN_IN), 
        .S(n9616), .Z(n9038) );
  XNOR2_X1 U11382 ( .A(n11714), .B(n9038), .ZN(n11862) );
  NAND2_X1 U11383 ( .A1(n11862), .A2(n7114), .ZN(n9021) );
  NAND2_X1 U11384 ( .A1(n6661), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n9020) );
  NAND2_X1 U11385 ( .A1(n13947), .A2(n9222), .ZN(n9033) );
  INV_X1 U11386 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n9023) );
  NAND2_X1 U11387 ( .A1(n9024), .A2(n9023), .ZN(n9025) );
  NAND2_X1 U11388 ( .A1(n9046), .A2(n9025), .ZN(n13797) );
  OR2_X1 U11389 ( .A1(n13797), .A2(n9198), .ZN(n9031) );
  INV_X1 U11390 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n9028) );
  NAND2_X1 U11391 ( .A1(n8553), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n9027) );
  NAND2_X1 U11392 ( .A1(n8571), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n9026) );
  OAI211_X1 U11393 ( .C1(n9195), .C2(n9028), .A(n9027), .B(n9026), .ZN(n9029)
         );
  INV_X1 U11394 ( .A(n9029), .ZN(n9030) );
  NAND2_X1 U11395 ( .A1(n9031), .A2(n9030), .ZN(n13656) );
  NAND2_X1 U11396 ( .A1(n13656), .A2(n9034), .ZN(n9032) );
  NAND2_X1 U11397 ( .A1(n9033), .A2(n9032), .ZN(n9036) );
  AOI22_X1 U11398 ( .A1(n13947), .A2(n9034), .B1(n9222), .B2(n13656), .ZN(
        n9035) );
  NAND2_X1 U11399 ( .A1(n9039), .A2(SI_22_), .ZN(n9040) );
  MUX2_X1 U11400 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(P1_DATAO_REG_23__SCAN_IN), 
        .S(n9616), .Z(n9062) );
  XNOR2_X1 U11401 ( .A(n9062), .B(SI_23_), .ZN(n9041) );
  NAND2_X1 U11402 ( .A1(n11731), .A2(n7114), .ZN(n9043) );
  NAND2_X1 U11403 ( .A1(n6661), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n9042) );
  NAND2_X1 U11404 ( .A1(n13942), .A2(n9199), .ZN(n9055) );
  INV_X1 U11405 ( .A(n9046), .ZN(n9044) );
  NAND2_X1 U11406 ( .A1(n9044), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n9066) );
  INV_X1 U11407 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n9045) );
  NAND2_X1 U11408 ( .A1(n9046), .A2(n9045), .ZN(n9047) );
  NAND2_X1 U11409 ( .A1(n9066), .A2(n9047), .ZN(n13786) );
  OR2_X1 U11410 ( .A1(n13786), .A2(n9198), .ZN(n9053) );
  INV_X1 U11411 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n9050) );
  NAND2_X1 U11412 ( .A1(n9191), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n9049) );
  NAND2_X1 U11413 ( .A1(n8571), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n9048) );
  OAI211_X1 U11414 ( .C1(n9195), .C2(n9050), .A(n9049), .B(n9048), .ZN(n9051)
         );
  INV_X1 U11415 ( .A(n9051), .ZN(n9052) );
  NAND2_X1 U11416 ( .A1(n9053), .A2(n9052), .ZN(n13686) );
  NAND2_X1 U11417 ( .A1(n13686), .A2(n9222), .ZN(n9054) );
  NAND2_X1 U11418 ( .A1(n9055), .A2(n9054), .ZN(n9057) );
  AOI22_X1 U11419 ( .A1(n13942), .A2(n9222), .B1(n9199), .B2(n13686), .ZN(
        n9056) );
  INV_X1 U11420 ( .A(n9062), .ZN(n9059) );
  NAND2_X1 U11421 ( .A1(n9059), .A2(n10969), .ZN(n9060) );
  NAND2_X1 U11422 ( .A1(n9062), .A2(SI_23_), .ZN(n9063) );
  MUX2_X1 U11423 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(P1_DATAO_REG_24__SCAN_IN), 
        .S(n9616), .Z(n9083) );
  XNOR2_X1 U11424 ( .A(n9082), .B(n9083), .ZN(n11750) );
  NAND2_X1 U11425 ( .A1(n11750), .A2(n7114), .ZN(n9065) );
  NAND2_X1 U11426 ( .A1(n6660), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n9064) );
  NAND2_X1 U11427 ( .A1(n13935), .A2(n9222), .ZN(n9075) );
  INV_X1 U11428 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n13527) );
  NAND2_X1 U11429 ( .A1(n9066), .A2(n13527), .ZN(n9067) );
  AND2_X1 U11430 ( .A1(n9094), .A2(n9067), .ZN(n13776) );
  NAND2_X1 U11431 ( .A1(n13776), .A2(n9214), .ZN(n9073) );
  INV_X1 U11432 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n9070) );
  NAND2_X1 U11433 ( .A1(n8571), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n9069) );
  NAND2_X1 U11434 ( .A1(n9191), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n9068) );
  OAI211_X1 U11435 ( .C1(n9195), .C2(n9070), .A(n9069), .B(n9068), .ZN(n9071)
         );
  INV_X1 U11436 ( .A(n9071), .ZN(n9072) );
  NAND2_X1 U11437 ( .A1(n9073), .A2(n9072), .ZN(n13660) );
  NAND2_X1 U11438 ( .A1(n13660), .A2(n9034), .ZN(n9074) );
  NAND2_X1 U11439 ( .A1(n9075), .A2(n9074), .ZN(n9080) );
  NAND2_X1 U11440 ( .A1(n13935), .A2(n9199), .ZN(n9076) );
  NAND2_X1 U11441 ( .A1(n9078), .A2(n9077), .ZN(n9079) );
  NAND2_X1 U11442 ( .A1(n9084), .A2(SI_24_), .ZN(n9085) );
  MUX2_X1 U11443 ( .A(n14816), .B(n14037), .S(n9616), .Z(n9087) );
  NAND2_X1 U11444 ( .A1(n9087), .A2(n11391), .ZN(n9107) );
  INV_X1 U11445 ( .A(n9087), .ZN(n9088) );
  NAND2_X1 U11446 ( .A1(n9088), .A2(SI_25_), .ZN(n9089) );
  NAND2_X1 U11447 ( .A1(n9107), .A2(n9089), .ZN(n9105) );
  NAND2_X1 U11448 ( .A1(n14035), .A2(n7114), .ZN(n9091) );
  NAND2_X1 U11449 ( .A1(n6661), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n9090) );
  NAND2_X1 U11450 ( .A1(n13927), .A2(n9034), .ZN(n9102) );
  INV_X1 U11451 ( .A(n9094), .ZN(n9092) );
  NAND2_X1 U11452 ( .A1(n9092), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n9112) );
  INV_X1 U11453 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n9093) );
  NAND2_X1 U11454 ( .A1(n9094), .A2(n9093), .ZN(n9095) );
  NAND2_X1 U11455 ( .A1(n9112), .A2(n9095), .ZN(n13762) );
  OR2_X1 U11456 ( .A1(n13762), .A2(n9198), .ZN(n9100) );
  INV_X1 U11457 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n13315) );
  NAND2_X1 U11458 ( .A1(n6662), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n9097) );
  NAND2_X1 U11459 ( .A1(n9191), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n9096) );
  OAI211_X1 U11460 ( .C1(n13315), .C2(n9217), .A(n9097), .B(n9096), .ZN(n9098)
         );
  INV_X1 U11461 ( .A(n9098), .ZN(n9099) );
  NAND2_X1 U11462 ( .A1(n13688), .A2(n9222), .ZN(n9101) );
  AOI22_X1 U11463 ( .A1(n13927), .A2(n9222), .B1(n9199), .B2(n13688), .ZN(
        n9103) );
  MUX2_X1 U11464 ( .A(n14810), .B(n14034), .S(n9616), .Z(n9124) );
  XNOR2_X1 U11465 ( .A(n9124), .B(SI_26_), .ZN(n9108) );
  NAND2_X1 U11466 ( .A1(n14032), .A2(n7114), .ZN(n9110) );
  NAND2_X1 U11467 ( .A1(n6661), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n9109) );
  NAND2_X1 U11468 ( .A1(n13918), .A2(n9222), .ZN(n9121) );
  INV_X1 U11469 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n9111) );
  NAND2_X1 U11470 ( .A1(n9112), .A2(n9111), .ZN(n9113) );
  NAND2_X1 U11471 ( .A1(n13745), .A2(n9214), .ZN(n9119) );
  INV_X1 U11472 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n9116) );
  NAND2_X1 U11473 ( .A1(n9191), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n9115) );
  NAND2_X1 U11474 ( .A1(n8571), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n9114) );
  OAI211_X1 U11475 ( .C1(n9195), .C2(n9116), .A(n9115), .B(n9114), .ZN(n9117)
         );
  INV_X1 U11476 ( .A(n9117), .ZN(n9118) );
  NAND2_X1 U11477 ( .A1(n13663), .A2(n9199), .ZN(n9120) );
  NAND2_X1 U11478 ( .A1(n9121), .A2(n9120), .ZN(n9123) );
  AOI22_X1 U11479 ( .A1(n13918), .A2(n9199), .B1(n8565), .B2(n13663), .ZN(
        n9122) );
  MUX2_X1 U11480 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(P1_DATAO_REG_27__SCAN_IN), 
        .S(n9616), .Z(n9145) );
  XNOR2_X1 U11481 ( .A(n9145), .B(n13471), .ZN(n9126) );
  NAND2_X1 U11482 ( .A1(n11804), .A2(n7114), .ZN(n9128) );
  NAND2_X1 U11483 ( .A1(n6661), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n9127) );
  INV_X1 U11484 ( .A(n9131), .ZN(n9129) );
  NAND2_X1 U11485 ( .A1(n9129), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n9212) );
  INV_X1 U11486 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n9130) );
  NAND2_X1 U11487 ( .A1(n9131), .A2(n9130), .ZN(n9132) );
  NAND2_X1 U11488 ( .A1(n9212), .A2(n9132), .ZN(n13079) );
  OR2_X1 U11489 ( .A1(n13079), .A2(n9198), .ZN(n9138) );
  INV_X1 U11490 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n9135) );
  NAND2_X1 U11491 ( .A1(n8571), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n9134) );
  NAND2_X1 U11492 ( .A1(n9191), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n9133) );
  OAI211_X1 U11493 ( .C1(n9195), .C2(n9135), .A(n9134), .B(n9133), .ZN(n9136)
         );
  INV_X1 U11494 ( .A(n9136), .ZN(n9137) );
  AND2_X1 U11495 ( .A1(n13694), .A2(n8565), .ZN(n9139) );
  AOI21_X1 U11496 ( .B1(n13912), .B2(n9199), .A(n9139), .ZN(n9205) );
  NAND2_X1 U11497 ( .A1(n13912), .A2(n9222), .ZN(n9140) );
  OAI21_X1 U11498 ( .B1(n9222), .B2(n13665), .A(n9140), .ZN(n9141) );
  INV_X1 U11499 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n9144) );
  NAND2_X1 U11500 ( .A1(n9191), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n9143) );
  NAND2_X1 U11501 ( .A1(n8571), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n9142) );
  OAI211_X1 U11502 ( .C1(n9195), .C2(n9144), .A(n9143), .B(n9142), .ZN(n13631)
         );
  INV_X1 U11503 ( .A(n9145), .ZN(n9146) );
  NAND2_X1 U11504 ( .A1(n9147), .A2(n13471), .ZN(n9148) );
  NAND2_X1 U11505 ( .A1(n9149), .A2(n9148), .ZN(n9208) );
  MUX2_X1 U11506 ( .A(n14809), .B(n13246), .S(n9616), .Z(n9150) );
  XNOR2_X1 U11507 ( .A(n9150), .B(SI_28_), .ZN(n9207) );
  NAND2_X1 U11508 ( .A1(n9208), .A2(n9207), .ZN(n9152) );
  NAND2_X1 U11509 ( .A1(n9150), .A2(n13061), .ZN(n9151) );
  INV_X1 U11510 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n14806) );
  INV_X1 U11511 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n14022) );
  MUX2_X1 U11512 ( .A(n14806), .B(n14022), .S(n9616), .Z(n9153) );
  XNOR2_X1 U11513 ( .A(n9153), .B(SI_29_), .ZN(n9187) );
  NAND2_X1 U11514 ( .A1(n9188), .A2(n9187), .ZN(n9155) );
  NAND2_X1 U11515 ( .A1(n9153), .A2(n13329), .ZN(n9154) );
  MUX2_X1 U11516 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n9616), .Z(n9156) );
  NAND2_X1 U11517 ( .A1(n9156), .A2(SI_30_), .ZN(n9157) );
  OAI21_X1 U11518 ( .B1(n9156), .B2(SI_30_), .A(n9157), .ZN(n9166) );
  MUX2_X1 U11519 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n9616), .Z(n9159) );
  XNOR2_X1 U11520 ( .A(n9159), .B(SI_31_), .ZN(n9160) );
  NAND2_X1 U11521 ( .A1(n14017), .A2(n7114), .ZN(n9163) );
  NAND2_X1 U11522 ( .A1(n6661), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n9162) );
  MUX2_X1 U11523 ( .A(n13631), .B(n8565), .S(n13632), .Z(n9165) );
  NAND2_X1 U11524 ( .A1(n13631), .A2(n9222), .ZN(n9164) );
  NAND2_X1 U11525 ( .A1(n9165), .A2(n9164), .ZN(n9204) );
  NAND2_X1 U11526 ( .A1(n9167), .A2(n9166), .ZN(n9168) );
  NAND2_X1 U11527 ( .A1(n6661), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n9171) );
  NAND2_X1 U11528 ( .A1(n6670), .A2(n10763), .ZN(n9667) );
  NAND2_X1 U11529 ( .A1(n9667), .A2(n9176), .ZN(n9675) );
  AOI21_X1 U11530 ( .B1(n9787), .B2(n6670), .A(n9675), .ZN(n9177) );
  INV_X1 U11531 ( .A(n9177), .ZN(n9178) );
  AOI21_X1 U11532 ( .B1(n13631), .B2(n9199), .A(n9178), .ZN(n9182) );
  NAND2_X1 U11533 ( .A1(n6662), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n9181) );
  NAND2_X1 U11534 ( .A1(n9191), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n9180) );
  NAND2_X1 U11535 ( .A1(n8571), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n9179) );
  AND3_X1 U11536 ( .A1(n9181), .A2(n9180), .A3(n9179), .ZN(n9184) );
  NOR2_X1 U11537 ( .A1(n9182), .A2(n9184), .ZN(n9183) );
  AOI21_X1 U11538 ( .B1(n13635), .B2(n9222), .A(n9183), .ZN(n9238) );
  NAND2_X1 U11539 ( .A1(n13635), .A2(n9199), .ZN(n9186) );
  INV_X1 U11540 ( .A(n9184), .ZN(n13699) );
  NAND2_X1 U11541 ( .A1(n13699), .A2(n9222), .ZN(n9185) );
  NAND2_X1 U11542 ( .A1(n9186), .A2(n9185), .ZN(n9237) );
  NAND2_X1 U11543 ( .A1(n14021), .A2(n7114), .ZN(n9190) );
  NAND2_X1 U11544 ( .A1(n6661), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n9189) );
  INV_X1 U11545 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n9211) );
  OR2_X1 U11546 ( .A1(n9212), .A2(n9211), .ZN(n13708) );
  INV_X1 U11547 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n9194) );
  NAND2_X1 U11548 ( .A1(n9191), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n9193) );
  NAND2_X1 U11549 ( .A1(n8571), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n9192) );
  OAI211_X1 U11550 ( .C1(n9195), .C2(n9194), .A(n9193), .B(n9192), .ZN(n9196)
         );
  INV_X1 U11551 ( .A(n9196), .ZN(n9197) );
  OAI21_X1 U11552 ( .B1(n13708), .B2(n9198), .A(n9197), .ZN(n13563) );
  AND2_X1 U11553 ( .A1(n13563), .A2(n9199), .ZN(n9200) );
  AOI21_X1 U11554 ( .B1(n13901), .B2(n9222), .A(n9200), .ZN(n9233) );
  NAND2_X1 U11555 ( .A1(n13901), .A2(n9199), .ZN(n9202) );
  NAND2_X1 U11556 ( .A1(n13563), .A2(n9222), .ZN(n9201) );
  NAND2_X1 U11557 ( .A1(n9202), .A2(n9201), .ZN(n9232) );
  OAI22_X1 U11558 ( .A1(n9238), .A2(n9237), .B1(n9233), .B2(n9232), .ZN(n9203)
         );
  NAND2_X1 U11559 ( .A1(n9204), .A2(n9203), .ZN(n9236) );
  NAND2_X1 U11560 ( .A1(n9206), .A2(n9205), .ZN(n9226) );
  XNOR2_X1 U11561 ( .A(n9208), .B(n9207), .ZN(n14024) );
  NAND2_X1 U11562 ( .A1(n14024), .A2(n7114), .ZN(n9210) );
  NAND2_X1 U11563 ( .A1(n6660), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n9209) );
  NAND2_X1 U11564 ( .A1(n9212), .A2(n9211), .ZN(n9213) );
  NAND2_X1 U11565 ( .A1(n13722), .A2(n9214), .ZN(n9220) );
  INV_X1 U11566 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n13317) );
  NAND2_X1 U11567 ( .A1(n6662), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n9216) );
  NAND2_X1 U11568 ( .A1(n8553), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n9215) );
  OAI211_X1 U11569 ( .C1(n13317), .C2(n9217), .A(n9216), .B(n9215), .ZN(n9218)
         );
  INV_X1 U11570 ( .A(n9218), .ZN(n9219) );
  AND2_X1 U11571 ( .A1(n13702), .A2(n8565), .ZN(n9221) );
  AOI21_X1 U11572 ( .B1(n13905), .B2(n9199), .A(n9221), .ZN(n9229) );
  NAND2_X1 U11573 ( .A1(n13905), .A2(n9222), .ZN(n9224) );
  NAND2_X1 U11574 ( .A1(n13702), .A2(n9034), .ZN(n9223) );
  NAND2_X1 U11575 ( .A1(n9224), .A2(n9223), .ZN(n9228) );
  NAND2_X1 U11576 ( .A1(n9229), .A2(n9228), .ZN(n9225) );
  XNOR2_X1 U11577 ( .A(n13632), .B(n13631), .ZN(n9248) );
  INV_X1 U11578 ( .A(n9228), .ZN(n9231) );
  INV_X1 U11579 ( .A(n9229), .ZN(n9230) );
  AOI22_X1 U11580 ( .A1(n9233), .A2(n9232), .B1(n9231), .B2(n9230), .ZN(n9234)
         );
  NAND2_X1 U11581 ( .A1(n9248), .A2(n9234), .ZN(n9235) );
  NAND2_X1 U11582 ( .A1(n9236), .A2(n9235), .ZN(n9240) );
  NAND2_X1 U11583 ( .A1(n9238), .A2(n9237), .ZN(n9239) );
  INV_X1 U11584 ( .A(n13631), .ZN(n9242) );
  OR3_X1 U11585 ( .A1(n13632), .A2(n9242), .A3(n9034), .ZN(n9244) );
  NAND3_X1 U11586 ( .A1(n13632), .A2(n9242), .A3(n9241), .ZN(n9243) );
  AND2_X1 U11587 ( .A1(n9244), .A2(n9243), .ZN(n9245) );
  INV_X1 U11588 ( .A(n6670), .ZN(n9247) );
  INV_X1 U11589 ( .A(n13563), .ZN(n13115) );
  XNOR2_X1 U11590 ( .A(n13635), .B(n13699), .ZN(n9267) );
  INV_X1 U11591 ( .A(n13702), .ZN(n13666) );
  NAND2_X1 U11592 ( .A1(n13905), .A2(n13666), .ZN(n9249) );
  INV_X1 U11593 ( .A(n13688), .ZN(n9250) );
  XNOR2_X1 U11594 ( .A(n13927), .B(n9250), .ZN(n13753) );
  INV_X1 U11595 ( .A(n13663), .ZN(n13498) );
  OR2_X1 U11596 ( .A1(n13918), .A2(n13498), .ZN(n13689) );
  NAND2_X1 U11597 ( .A1(n13918), .A2(n13498), .ZN(n13690) );
  NAND2_X1 U11598 ( .A1(n13689), .A2(n13690), .ZN(n13749) );
  NAND2_X1 U11599 ( .A1(n13935), .A2(n13497), .ZN(n13687) );
  NAND2_X1 U11600 ( .A1(n13687), .A2(n9251), .ZN(n13770) );
  INV_X1 U11601 ( .A(n13686), .ZN(n11913) );
  XNOR2_X1 U11602 ( .A(n13942), .B(n11913), .ZN(n13783) );
  XNOR2_X1 U11603 ( .A(n13953), .B(n11912), .ZN(n13683) );
  INV_X1 U11604 ( .A(n13680), .ZN(n13682) );
  XNOR2_X1 U11605 ( .A(n13681), .B(n13682), .ZN(n13819) );
  XNOR2_X1 U11606 ( .A(n13845), .B(n13676), .ZN(n13855) );
  OR2_X1 U11607 ( .A1(n13965), .A2(n13679), .ZN(n13650) );
  NAND2_X1 U11608 ( .A1(n13965), .A2(n13679), .ZN(n13649) );
  NAND2_X1 U11609 ( .A1(n13650), .A2(n13649), .ZN(n13838) );
  XNOR2_X1 U11610 ( .A(n13991), .B(n13667), .ZN(n13641) );
  OR2_X1 U11611 ( .A1(n15127), .A2(n9252), .ZN(n11528) );
  NAND2_X1 U11612 ( .A1(n15127), .A2(n9252), .ZN(n9253) );
  NAND2_X1 U11613 ( .A1(n11528), .A2(n9253), .ZN(n11492) );
  XNOR2_X1 U11614 ( .A(n11491), .B(n11495), .ZN(n11328) );
  INV_X1 U11615 ( .A(n13566), .ZN(n11327) );
  XNOR2_X1 U11616 ( .A(n15140), .B(n11327), .ZN(n15141) );
  XNOR2_X1 U11617 ( .A(n11323), .B(n13567), .ZN(n11325) );
  INV_X1 U11618 ( .A(n13570), .ZN(n10796) );
  XNOR2_X1 U11619 ( .A(n15530), .B(n10796), .ZN(n10897) );
  XNOR2_X2 U11620 ( .A(n13577), .B(n6672), .ZN(n10299) );
  OAI21_X1 U11621 ( .B1(n13578), .B2(n10295), .A(n10294), .ZN(n15494) );
  NAND4_X1 U11622 ( .A1(n10299), .A2(n9901), .A3(n15494), .A4(n9247), .ZN(
        n9254) );
  NOR3_X1 U11623 ( .A1(n9254), .A2(n10239), .A3(n9956), .ZN(n9256) );
  XNOR2_X1 U11624 ( .A(n10794), .B(n13571), .ZN(n10552) );
  NAND2_X1 U11625 ( .A1(n15513), .A2(n9255), .ZN(n10536) );
  XNOR2_X1 U11626 ( .A(n13573), .B(n10543), .ZN(n10244) );
  NAND4_X1 U11627 ( .A1(n9256), .A2(n10552), .A3(n10535), .A4(n10244), .ZN(
        n9257) );
  NOR2_X1 U11628 ( .A1(n10897), .A2(n9257), .ZN(n9258) );
  XNOR2_X1 U11629 ( .A(n11229), .B(n13568), .ZN(n10992) );
  XNOR2_X1 U11630 ( .A(n15538), .B(n13569), .ZN(n10788) );
  NAND4_X1 U11631 ( .A1(n11325), .A2(n9258), .A3(n10992), .A4(n10788), .ZN(
        n9259) );
  OR4_X1 U11632 ( .A1(n11492), .A2(n11328), .A3(n15141), .A4(n9259), .ZN(n9260) );
  NOR2_X1 U11633 ( .A1(n13641), .A2(n9260), .ZN(n9261) );
  XNOR2_X1 U11634 ( .A(n13985), .B(n13670), .ZN(n13880) );
  NAND2_X1 U11635 ( .A1(n13673), .A2(n13672), .ZN(n13647) );
  NAND2_X1 U11636 ( .A1(n13648), .A2(n13647), .ZN(n13862) );
  NAND4_X1 U11637 ( .A1(n13838), .A2(n9261), .A3(n13880), .A4(n13862), .ZN(
        n9262) );
  OR4_X1 U11638 ( .A1(n13683), .A2(n13819), .A3(n13855), .A4(n9262), .ZN(n9263) );
  NOR2_X1 U11639 ( .A1(n13718), .A2(n9265), .ZN(n9266) );
  NAND4_X1 U11640 ( .A1(n8520), .A2(n9269), .A3(n9268), .A4(n8525), .ZN(n9270)
         );
  NAND2_X1 U11641 ( .A1(n9273), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9272) );
  MUX2_X1 U11642 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9272), .S(
        P2_IR_REG_23__SCAN_IN), .Z(n9274) );
  INV_X1 U11643 ( .A(n9277), .ZN(n9281) );
  NOR2_X1 U11644 ( .A1(n9394), .A2(P2_U3088), .ZN(n11245) );
  INV_X1 U11645 ( .A(n11245), .ZN(n9298) );
  INV_X1 U11646 ( .A(P2_B_REG_SCAN_IN), .ZN(n13628) );
  NAND2_X1 U11647 ( .A1(n9277), .A2(n9276), .ZN(n9283) );
  NAND2_X1 U11648 ( .A1(n9283), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9278) );
  MUX2_X1 U11649 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9278), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n9280) );
  NAND2_X1 U11650 ( .A1(n9281), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9282) );
  MUX2_X1 U11651 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9282), .S(
        P2_IR_REG_24__SCAN_IN), .Z(n9284) );
  NAND2_X1 U11652 ( .A1(n9285), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9286) );
  NOR2_X1 U11653 ( .A1(n11511), .A2(n14033), .ZN(n9287) );
  INV_X1 U11654 ( .A(n15491), .ZN(n15488) );
  INV_X1 U11655 ( .A(n9288), .ZN(n9289) );
  NAND2_X1 U11656 ( .A1(n9672), .A2(n9289), .ZN(n13496) );
  NOR4_X1 U11657 ( .A1(n15488), .A2(n9667), .A3(n14029), .A4(n13496), .ZN(
        n9290) );
  AOI211_X1 U11658 ( .C1(n11245), .C2(n9173), .A(n13628), .B(n9290), .ZN(n9291) );
  INV_X1 U11659 ( .A(n9667), .ZN(n9670) );
  AOI211_X1 U11660 ( .C1(n9176), .C2(n10763), .A(n9670), .B(n9293), .ZN(n9294)
         );
  MUX2_X1 U11661 ( .A(n9642), .B(n9176), .S(n9247), .Z(n9296) );
  NAND2_X1 U11662 ( .A1(n9296), .A2(n9175), .ZN(n9297) );
  NAND2_X1 U11663 ( .A1(n9394), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9299) );
  NOR2_X1 U11664 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n9301) );
  NOR2_X1 U11665 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n9300) );
  NOR2_X1 U11666 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), 
        .ZN(n9313) );
  NOR2_X1 U11667 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), 
        .ZN(n9312) );
  NAND2_X1 U11668 ( .A1(n9314), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9315) );
  MUX2_X1 U11669 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9315), .S(
        P1_IR_REG_25__SCAN_IN), .Z(n9318) );
  NAND2_X1 U11670 ( .A1(n9318), .A2(n9457), .ZN(n14813) );
  NAND2_X1 U11671 ( .A1(n9319), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9320) );
  NOR2_X1 U11672 ( .A1(n14813), .A2(n11509), .ZN(n9322) );
  NAND2_X1 U11673 ( .A1(n9457), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9321) );
  INV_X1 U11674 ( .A(n9630), .ZN(n9623) );
  INV_X2 U11675 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  INV_X1 U11676 ( .A(n14945), .ZN(n14938) );
  OAI222_X1 U11677 ( .A1(n14938), .A2(n9325), .B1(n14936), .B2(n9324), .C1(
        P3_U3151), .C2(n11024), .ZN(P3_U3287) );
  OAI222_X1 U11678 ( .A1(n14938), .A2(n9327), .B1(n14936), .B2(n9326), .C1(
        P3_U3151), .C2(n10365), .ZN(P3_U3294) );
  OAI222_X1 U11679 ( .A1(n14938), .A2(n9329), .B1(n14936), .B2(n9328), .C1(
        P3_U3151), .C2(n10401), .ZN(P3_U3289) );
  NOR2_X1 U11680 ( .A1(n9616), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14026) );
  INV_X2 U11681 ( .A(n14026), .ZN(n14038) );
  NAND2_X2 U11682 ( .A1(n9616), .A2(P2_U3088), .ZN(n14031) );
  INV_X1 U11683 ( .A(n9432), .ZN(n9438) );
  OAI222_X1 U11684 ( .A1(n14038), .A2(n9330), .B1(n14031), .B2(n9982), .C1(
        P2_U3088), .C2(n9438), .ZN(P2_U3325) );
  INV_X1 U11685 ( .A(n9448), .ZN(n9456) );
  OAI222_X1 U11686 ( .A1(n14038), .A2(n9331), .B1(n14031), .B2(n10130), .C1(
        P2_U3088), .C2(n9456), .ZN(P2_U3324) );
  OAI222_X1 U11687 ( .A1(P3_U3151), .A2(n10519), .B1(n14938), .B2(n9332), .C1(
        n9615), .C2(n14936), .ZN(P3_U3295) );
  NAND2_X2 U11688 ( .A1(n9616), .A2(P1_U3086), .ZN(n14817) );
  INV_X1 U11689 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n9335) );
  NOR2_X1 U11690 ( .A1(n9333), .A2(n9307), .ZN(n14258) );
  INV_X1 U11691 ( .A(n14258), .ZN(n9334) );
  OAI222_X1 U11692 ( .A1(n14817), .A2(n9335), .B1(n14815), .B2(n9982), .C1(
        P1_U3086), .C2(n9334), .ZN(P1_U3353) );
  NAND2_X1 U11693 ( .A1(n9337), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9338) );
  MUX2_X1 U11694 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9338), .S(
        P1_IR_REG_3__SCAN_IN), .Z(n9340) );
  AND2_X1 U11695 ( .A1(n9340), .A2(n9343), .ZN(n14265) );
  INV_X1 U11696 ( .A(n14265), .ZN(n9710) );
  OAI222_X1 U11697 ( .A1(n14817), .A2(n9341), .B1(n14815), .B2(n10130), .C1(
        P1_U3086), .C2(n9710), .ZN(P1_U3352) );
  INV_X1 U11698 ( .A(n9342), .ZN(n10125) );
  OAI222_X1 U11699 ( .A1(n14038), .A2(n13274), .B1(n14031), .B2(n10125), .C1(
        P2_U3088), .C2(n15419), .ZN(P2_U3323) );
  NAND2_X1 U11700 ( .A1(n9343), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9344) );
  XNOR2_X1 U11701 ( .A(n9344), .B(P1_IR_REG_4__SCAN_IN), .ZN(n14284) );
  INV_X1 U11702 ( .A(n14284), .ZN(n14275) );
  OAI222_X1 U11703 ( .A1(n14817), .A2(n7179), .B1(n14815), .B2(n10125), .C1(
        P1_U3086), .C2(n14275), .ZN(P1_U3351) );
  INV_X1 U11704 ( .A(n14936), .ZN(n14944) );
  AOI222_X1 U11705 ( .A1(n9345), .A2(n14945), .B1(SI_10_), .B2(n14944), .C1(
        n12679), .C2(P3_STATE_REG_SCAN_IN), .ZN(n9346) );
  INV_X1 U11706 ( .A(n9346), .ZN(P3_U3285) );
  AOI222_X1 U11707 ( .A1(n9347), .A2(n14945), .B1(SI_11_), .B2(n14944), .C1(
        n12682), .C2(P3_STATE_REG_SCAN_IN), .ZN(n9348) );
  INV_X1 U11708 ( .A(n9348), .ZN(P3_U3284) );
  AOI222_X1 U11709 ( .A1(n9349), .A2(n14945), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n10107), .C1(SI_2_), .C2(n14944), .ZN(n9350) );
  INV_X1 U11710 ( .A(n9350), .ZN(P3_U3293) );
  AOI222_X1 U11711 ( .A1(n9351), .A2(n14945), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n10258), .C1(SI_4_), .C2(n14944), .ZN(n9352) );
  INV_X1 U11712 ( .A(n9352), .ZN(P3_U3291) );
  AOI222_X1 U11713 ( .A1(n9353), .A2(n14945), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n10280), .C1(SI_3_), .C2(n14944), .ZN(n9354) );
  INV_X1 U11714 ( .A(n9354), .ZN(P3_U3292) );
  AOI222_X1 U11715 ( .A1(n9355), .A2(n14945), .B1(n10599), .B2(
        P3_STATE_REG_SCAN_IN), .C1(SI_7_), .C2(n14944), .ZN(n9356) );
  INV_X1 U11716 ( .A(n9356), .ZN(P3_U3288) );
  AOI222_X1 U11717 ( .A1(n9357), .A2(n14945), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n10333), .C1(SI_5_), .C2(n14944), .ZN(n9358) );
  INV_X1 U11718 ( .A(n9358), .ZN(P3_U3290) );
  OAI222_X1 U11719 ( .A1(n14038), .A2(n9359), .B1(n14031), .B2(n9818), .C1(
        P2_U3088), .C2(n8537), .ZN(P2_U3326) );
  NAND2_X1 U11720 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n9360) );
  INV_X1 U11721 ( .A(n14234), .ZN(n9361) );
  OAI222_X1 U11722 ( .A1(n14817), .A2(n9362), .B1(n14815), .B2(n9818), .C1(
        P1_U3086), .C2(n9361), .ZN(P1_U3354) );
  INV_X1 U11723 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n9363) );
  INV_X1 U11724 ( .A(n10424), .ZN(n9365) );
  OAI222_X1 U11725 ( .A1(n14038), .A2(n9363), .B1(n14031), .B2(n9365), .C1(
        P2_U3088), .C2(n6847), .ZN(P2_U3322) );
  OR2_X1 U11726 ( .A1(n9370), .A2(n9336), .ZN(n9364) );
  XNOR2_X1 U11727 ( .A(n9364), .B(P1_IR_REG_5__SCAN_IN), .ZN(n14299) );
  OAI222_X1 U11728 ( .A1(n14817), .A2(n10427), .B1(n14815), .B2(n9365), .C1(
        P1_U3086), .C2(n6958), .ZN(P1_U3350) );
  OAI222_X1 U11729 ( .A1(P3_U3151), .A2(n15640), .B1(n14936), .B2(n9367), .C1(
        n14938), .C2(n9366), .ZN(P3_U3283) );
  INV_X1 U11730 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n9368) );
  INV_X1 U11731 ( .A(n10437), .ZN(n9372) );
  INV_X1 U11732 ( .A(n9486), .ZN(n15439) );
  OAI222_X1 U11733 ( .A1(n14038), .A2(n9368), .B1(n14031), .B2(n9372), .C1(
        P2_U3088), .C2(n15439), .ZN(P2_U3321) );
  INV_X1 U11734 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n9369) );
  AND2_X1 U11735 ( .A1(n9370), .A2(n9369), .ZN(n10231) );
  OR2_X1 U11736 ( .A1(n10231), .A2(n9336), .ZN(n9371) );
  XNOR2_X1 U11737 ( .A(n9371), .B(P1_IR_REG_6__SCAN_IN), .ZN(n10436) );
  INV_X1 U11738 ( .A(n10436), .ZN(n9714) );
  OAI222_X1 U11739 ( .A1(n14817), .A2(n9373), .B1(n14815), .B2(n9372), .C1(
        P1_U3086), .C2(n9714), .ZN(P1_U3349) );
  INV_X1 U11740 ( .A(n10736), .ZN(n9378) );
  NAND2_X1 U11741 ( .A1(n10231), .A2(n9374), .ZN(n9388) );
  NAND2_X1 U11742 ( .A1(n9388), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9375) );
  XNOR2_X1 U11743 ( .A(n9375), .B(P1_IR_REG_7__SCAN_IN), .ZN(n14317) );
  INV_X1 U11744 ( .A(n14317), .ZN(n9716) );
  OAI222_X1 U11745 ( .A1(n14817), .A2(n9376), .B1(n14815), .B2(n9378), .C1(
        P1_U3086), .C2(n9716), .ZN(P1_U3348) );
  INV_X1 U11746 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n9379) );
  INV_X1 U11747 ( .A(n13589), .ZN(n9377) );
  OAI222_X1 U11748 ( .A1(n14038), .A2(n9379), .B1(n14031), .B2(n9378), .C1(
        P2_U3088), .C2(n9377), .ZN(P2_U3320) );
  AND2_X1 U11749 ( .A1(n9386), .A2(n9630), .ZN(n9975) );
  NAND2_X1 U11750 ( .A1(n14813), .A2(P1_B_REG_SCAN_IN), .ZN(n9381) );
  MUX2_X1 U11751 ( .A(n9381), .B(P1_B_REG_SCAN_IN), .S(n9380), .Z(n9382) );
  NAND2_X1 U11752 ( .A1(n9382), .A2(n9383), .ZN(n9755) );
  NAND2_X1 U11753 ( .A1(n9975), .A2(n9755), .ZN(n15314) );
  INV_X1 U11754 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n9385) );
  INV_X1 U11755 ( .A(n9383), .ZN(n14812) );
  NAND2_X1 U11756 ( .A1(n14812), .A2(n14813), .ZN(n9595) );
  INV_X1 U11757 ( .A(n9595), .ZN(n9384) );
  AOI22_X1 U11758 ( .A1(n15314), .A2(n9385), .B1(n9384), .B2(n9386), .ZN(
        P1_U3446) );
  INV_X1 U11759 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n9606) );
  NAND2_X1 U11760 ( .A1(n14812), .A2(n11509), .ZN(n9754) );
  INV_X1 U11761 ( .A(n9754), .ZN(n9387) );
  AOI22_X1 U11762 ( .A1(n15314), .A2(n9606), .B1(n9387), .B2(n9386), .ZN(
        P1_U3445) );
  INV_X1 U11763 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n13209) );
  INV_X1 U11764 ( .A(n10828), .ZN(n9390) );
  OAI222_X1 U11765 ( .A1(n14038), .A2(n13209), .B1(n14031), .B2(n9390), .C1(
        P2_U3088), .C2(n9489), .ZN(P2_U3319) );
  NAND2_X1 U11766 ( .A1(n9392), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9389) );
  XNOR2_X1 U11767 ( .A(n9389), .B(P1_IR_REG_8__SCAN_IN), .ZN(n10829) );
  INV_X1 U11768 ( .A(n10829), .ZN(n9723) );
  OAI222_X1 U11769 ( .A1(n14817), .A2(n9391), .B1(n14815), .B2(n9390), .C1(
        P1_U3086), .C2(n9723), .ZN(P1_U3347) );
  INV_X1 U11770 ( .A(n11065), .ZN(n9470) );
  OR2_X1 U11771 ( .A1(n9550), .A2(n9336), .ZN(n9473) );
  XNOR2_X1 U11772 ( .A(n9473), .B(P1_IR_REG_9__SCAN_IN), .ZN(n14339) );
  INV_X1 U11773 ( .A(n14817), .ZN(n14797) );
  AOI22_X1 U11774 ( .A1(n14339), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n14797), .ZN(n9393) );
  OAI21_X1 U11775 ( .B1(n9470), .B2(n14815), .A(n9393), .ZN(P1_U3346) );
  INV_X1 U11776 ( .A(n9394), .ZN(n9397) );
  NAND2_X1 U11777 ( .A1(n9672), .A2(n9394), .ZN(n9395) );
  NAND2_X1 U11778 ( .A1(n9395), .A2(n8535), .ZN(n9396) );
  OAI21_X1 U11779 ( .B1(n9398), .B2(n9397), .A(n9396), .ZN(n9399) );
  NAND2_X1 U11780 ( .A1(n9399), .A2(n9288), .ZN(n15420) );
  OR2_X1 U11781 ( .A1(n9399), .A2(P2_U3088), .ZN(n15450) );
  INV_X1 U11782 ( .A(n15450), .ZN(n15472) );
  NAND2_X1 U11783 ( .A1(P2_U3088), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n10166) );
  INV_X1 U11784 ( .A(n10166), .ZN(n9407) );
  NOR2_X1 U11785 ( .A1(n9288), .A2(P2_U3088), .ZN(n14025) );
  NAND2_X1 U11786 ( .A1(n9399), .A2(n14025), .ZN(n9408) );
  INV_X1 U11787 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n9401) );
  INV_X1 U11788 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n9400) );
  MUX2_X1 U11789 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n9400), .S(n9412), .Z(n15410) );
  NAND3_X1 U11790 ( .A1(n15410), .A2(P2_IR_REG_0__SCAN_IN), .A3(
        P2_REG2_REG_0__SCAN_IN), .ZN(n15409) );
  NAND2_X1 U11791 ( .A1(n9412), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n9427) );
  INV_X1 U11792 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n10666) );
  NOR2_X1 U11793 ( .A1(n9438), .A2(n10666), .ZN(n9442) );
  MUX2_X1 U11794 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n9401), .S(n9448), .Z(n9441)
         );
  OAI21_X1 U11795 ( .B1(n9443), .B2(n9442), .A(n9441), .ZN(n9440) );
  OAI21_X1 U11796 ( .B1(n9401), .B2(n9456), .A(n9440), .ZN(n15424) );
  INV_X1 U11797 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n9402) );
  MUX2_X1 U11798 ( .A(n9402), .B(P2_REG2_REG_4__SCAN_IN), .S(n15419), .Z(
        n15423) );
  NAND2_X1 U11799 ( .A1(n15424), .A2(n15423), .ZN(n15422) );
  OR2_X1 U11800 ( .A1(n15419), .A2(n9402), .ZN(n9404) );
  MUX2_X1 U11801 ( .A(n6846), .B(P2_REG2_REG_5__SCAN_IN), .S(n9485), .Z(n9403)
         );
  AND3_X1 U11802 ( .A1(n15422), .A2(n9404), .A3(n9403), .ZN(n9405) );
  NOR3_X1 U11803 ( .A1(n15442), .A2(n9477), .A3(n9405), .ZN(n9406) );
  AOI211_X1 U11804 ( .C1(n15472), .C2(P2_ADDR_REG_5__SCAN_IN), .A(n9407), .B(
        n9406), .ZN(n9426) );
  INV_X1 U11805 ( .A(n9408), .ZN(n9409) );
  INV_X1 U11806 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n9410) );
  MUX2_X1 U11807 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n9410), .S(n9432), .Z(n9414)
         );
  INV_X1 U11808 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n9411) );
  MUX2_X1 U11809 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n9411), .S(n9412), .Z(n15413) );
  AND2_X1 U11810 ( .A1(P2_REG1_REG_0__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), 
        .ZN(n15414) );
  NAND2_X1 U11811 ( .A1(n15413), .A2(n15414), .ZN(n15412) );
  NAND2_X1 U11812 ( .A1(n9412), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n9433) );
  NAND2_X1 U11813 ( .A1(n15412), .A2(n9433), .ZN(n9413) );
  NAND2_X1 U11814 ( .A1(n9414), .A2(n9413), .ZN(n9451) );
  NAND2_X1 U11815 ( .A1(n9432), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n9450) );
  NAND2_X1 U11816 ( .A1(n9451), .A2(n9450), .ZN(n9416) );
  MUX2_X1 U11817 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n9916), .S(n9448), .Z(n9415)
         );
  NAND2_X1 U11818 ( .A1(n9416), .A2(n9415), .ZN(n9453) );
  NAND2_X1 U11819 ( .A1(n9448), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n9417) );
  NAND2_X1 U11820 ( .A1(n9453), .A2(n9417), .ZN(n15427) );
  INV_X1 U11821 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n9418) );
  MUX2_X1 U11822 ( .A(n9418), .B(P2_REG1_REG_4__SCAN_IN), .S(n15419), .Z(
        n15426) );
  NAND2_X1 U11823 ( .A1(n15427), .A2(n15426), .ZN(n15425) );
  OR2_X1 U11824 ( .A1(n15419), .A2(n9418), .ZN(n9423) );
  NAND2_X1 U11825 ( .A1(n15425), .A2(n9423), .ZN(n9421) );
  INV_X1 U11826 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n9419) );
  MUX2_X1 U11827 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n9419), .S(n9485), .Z(n9420)
         );
  NAND2_X1 U11828 ( .A1(n9421), .A2(n9420), .ZN(n15434) );
  MUX2_X1 U11829 ( .A(n9419), .B(P2_REG1_REG_5__SCAN_IN), .S(n9485), .Z(n9422)
         );
  NAND3_X1 U11830 ( .A1(n15425), .A2(n9423), .A3(n9422), .ZN(n9424) );
  NAND3_X1 U11831 ( .A1(n15467), .A2(n15434), .A3(n9424), .ZN(n9425) );
  OAI211_X1 U11832 ( .C1(n15479), .C2(n6847), .A(n9426), .B(n9425), .ZN(
        P2_U3219) );
  AND2_X1 U11833 ( .A1(P2_U3088), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n9431) );
  AND3_X1 U11834 ( .A1(n9428), .A2(n15409), .A3(n9427), .ZN(n9429) );
  NOR3_X1 U11835 ( .A1(n15442), .A2(n9443), .A3(n9429), .ZN(n9430) );
  AOI211_X1 U11836 ( .C1(n15472), .C2(P2_ADDR_REG_2__SCAN_IN), .A(n9431), .B(
        n9430), .ZN(n9437) );
  MUX2_X1 U11837 ( .A(n9410), .B(P2_REG1_REG_2__SCAN_IN), .S(n9432), .Z(n9434)
         );
  NAND3_X1 U11838 ( .A1(n9434), .A2(n15412), .A3(n9433), .ZN(n9435) );
  NAND3_X1 U11839 ( .A1(n15467), .A2(n9451), .A3(n9435), .ZN(n9436) );
  OAI211_X1 U11840 ( .C1(n15479), .C2(n9438), .A(n9437), .B(n9436), .ZN(
        P2_U3216) );
  INV_X1 U11841 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n9439) );
  NOR2_X1 U11842 ( .A1(n15450), .A2(n9439), .ZN(n9447) );
  INV_X1 U11843 ( .A(n9440), .ZN(n9445) );
  NOR3_X1 U11844 ( .A1(n9443), .A2(n9442), .A3(n9441), .ZN(n9444) );
  NOR3_X1 U11845 ( .A1(n15442), .A2(n9445), .A3(n9444), .ZN(n9446) );
  AOI211_X1 U11846 ( .C1(P2_REG3_REG_3__SCAN_IN), .C2(P2_U3088), .A(n9447), 
        .B(n9446), .ZN(n9455) );
  INV_X1 U11847 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n9916) );
  MUX2_X1 U11848 ( .A(n9916), .B(P2_REG1_REG_3__SCAN_IN), .S(n9448), .Z(n9449)
         );
  NAND3_X1 U11849 ( .A1(n9451), .A2(n9450), .A3(n9449), .ZN(n9452) );
  NAND3_X1 U11850 ( .A1(n15467), .A2(n9453), .A3(n9452), .ZN(n9454) );
  OAI211_X1 U11851 ( .C1(n15479), .C2(n9456), .A(n9455), .B(n9454), .ZN(
        P2_U3217) );
  OR2_X1 U11852 ( .A1(n9631), .A2(P1_U3086), .ZN(n12189) );
  INV_X1 U11853 ( .A(n12189), .ZN(n11243) );
  INV_X1 U11854 ( .A(n9556), .ZN(n9554) );
  NAND2_X1 U11855 ( .A1(n9458), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9459) );
  MUX2_X1 U11856 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9463), .S(
        P1_IR_REG_21__SCAN_IN), .Z(n9464) );
  INV_X1 U11857 ( .A(n12141), .ZN(n9468) );
  NAND2_X1 U11858 ( .A1(n9465), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9467) );
  NAND2_X1 U11859 ( .A1(n12134), .A2(n9631), .ZN(n9469) );
  NAND2_X1 U11860 ( .A1(n9817), .A2(n9469), .ZN(n9719) );
  INV_X1 U11861 ( .A(n15271), .ZN(n14360) );
  NOR2_X1 U11862 ( .A1(n14360), .A2(P1_U4016), .ZN(P1_U3085) );
  INV_X1 U11863 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n9471) );
  OAI222_X1 U11864 ( .A1(n14038), .A2(n9471), .B1(n14031), .B2(n9470), .C1(
        P2_U3088), .C2(n9537), .ZN(P2_U3318) );
  INV_X1 U11865 ( .A(n11071), .ZN(n9527) );
  INV_X1 U11866 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n9472) );
  NAND2_X1 U11867 ( .A1(n9473), .A2(n9472), .ZN(n9474) );
  NAND2_X1 U11868 ( .A1(n9474), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9475) );
  XNOR2_X1 U11869 ( .A(n9475), .B(P1_IR_REG_10__SCAN_IN), .ZN(n11072) );
  AOI22_X1 U11870 ( .A1(n11072), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n14797), .ZN(n9476) );
  OAI21_X1 U11871 ( .B1(n9527), .B2(n14815), .A(n9476), .ZN(P1_U3345) );
  INV_X1 U11872 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n9478) );
  MUX2_X1 U11873 ( .A(n9478), .B(P2_REG2_REG_6__SCAN_IN), .S(n9486), .Z(n15443) );
  NOR2_X1 U11874 ( .A1(n15439), .A2(n9478), .ZN(n13579) );
  INV_X1 U11875 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n10538) );
  MUX2_X1 U11876 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n10538), .S(n13589), .Z(
        n9479) );
  NAND2_X1 U11877 ( .A1(n13589), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n9482) );
  INV_X1 U11878 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n9480) );
  MUX2_X1 U11879 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n9480), .S(n9489), .Z(n9481)
         );
  AOI21_X1 U11880 ( .B1(n13582), .B2(n9482), .A(n9481), .ZN(n9529) );
  NAND3_X1 U11881 ( .A1(n13582), .A2(n9482), .A3(n9481), .ZN(n9483) );
  NAND2_X1 U11882 ( .A1(n9483), .A2(n15474), .ZN(n9496) );
  INV_X1 U11883 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n9484) );
  NAND2_X1 U11884 ( .A1(P2_U3088), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n10637) );
  OAI21_X1 U11885 ( .B1(n15450), .B2(n9484), .A(n10637), .ZN(n9494) );
  INV_X1 U11886 ( .A(n15467), .ZN(n15459) );
  NAND2_X1 U11887 ( .A1(n9485), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n15433) );
  INV_X1 U11888 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n15566) );
  MUX2_X1 U11889 ( .A(n15566), .B(P2_REG1_REG_6__SCAN_IN), .S(n9486), .Z(
        n15432) );
  AOI21_X1 U11890 ( .B1(n15434), .B2(n15433), .A(n15432), .ZN(n13587) );
  NOR2_X1 U11891 ( .A1(n15439), .A2(n15566), .ZN(n13588) );
  INV_X1 U11892 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n9487) );
  MUX2_X1 U11893 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n9487), .S(n13589), .Z(n9488) );
  OAI21_X1 U11894 ( .B1(n13587), .B2(n13588), .A(n9488), .ZN(n13593) );
  NAND2_X1 U11895 ( .A1(n13589), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n9491) );
  INV_X1 U11896 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n15569) );
  MUX2_X1 U11897 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n15569), .S(n9489), .Z(n9490) );
  AOI21_X1 U11898 ( .B1(n13593), .B2(n9491), .A(n9490), .ZN(n9534) );
  AND3_X1 U11899 ( .A1(n13593), .A2(n9491), .A3(n9490), .ZN(n9492) );
  NOR3_X1 U11900 ( .A1(n15459), .A2(n9534), .A3(n9492), .ZN(n9493) );
  AOI211_X1 U11901 ( .C1(n15453), .C2(n9535), .A(n9494), .B(n9493), .ZN(n9495)
         );
  OAI21_X1 U11902 ( .B1(n9529), .B2(n9496), .A(n9495), .ZN(P2_U3222) );
  NOR2_X1 U11903 ( .A1(n9497), .A2(n13051), .ZN(n9499) );
  CLKBUF_X1 U11904 ( .A(n9499), .Z(n9525) );
  INV_X1 U11905 ( .A(P3_D_REG_15__SCAN_IN), .ZN(n9498) );
  NOR2_X1 U11906 ( .A1(n9525), .A2(n9498), .ZN(P3_U3250) );
  INV_X1 U11907 ( .A(P3_D_REG_20__SCAN_IN), .ZN(n9500) );
  NOR2_X1 U11908 ( .A1(n9525), .A2(n9500), .ZN(P3_U3245) );
  INV_X1 U11909 ( .A(P3_D_REG_27__SCAN_IN), .ZN(n9501) );
  NOR2_X1 U11910 ( .A1(n9499), .A2(n9501), .ZN(P3_U3238) );
  INV_X1 U11911 ( .A(P3_D_REG_14__SCAN_IN), .ZN(n9502) );
  NOR2_X1 U11912 ( .A1(n9525), .A2(n9502), .ZN(P3_U3251) );
  INV_X1 U11913 ( .A(P3_D_REG_29__SCAN_IN), .ZN(n9503) );
  NOR2_X1 U11914 ( .A1(n9499), .A2(n9503), .ZN(P3_U3236) );
  INV_X1 U11915 ( .A(P3_D_REG_24__SCAN_IN), .ZN(n9504) );
  NOR2_X1 U11916 ( .A1(n9499), .A2(n9504), .ZN(P3_U3241) );
  INV_X1 U11917 ( .A(P3_D_REG_13__SCAN_IN), .ZN(n9505) );
  NOR2_X1 U11918 ( .A1(n9525), .A2(n9505), .ZN(P3_U3252) );
  INV_X1 U11919 ( .A(P3_D_REG_19__SCAN_IN), .ZN(n9506) );
  NOR2_X1 U11920 ( .A1(n9525), .A2(n9506), .ZN(P3_U3246) );
  INV_X1 U11921 ( .A(P3_D_REG_3__SCAN_IN), .ZN(n9507) );
  NOR2_X1 U11922 ( .A1(n9499), .A2(n9507), .ZN(P3_U3262) );
  INV_X1 U11923 ( .A(P3_D_REG_28__SCAN_IN), .ZN(n9508) );
  NOR2_X1 U11924 ( .A1(n9499), .A2(n9508), .ZN(P3_U3237) );
  INV_X1 U11925 ( .A(P3_D_REG_5__SCAN_IN), .ZN(n9509) );
  NOR2_X1 U11926 ( .A1(n9499), .A2(n9509), .ZN(P3_U3260) );
  INV_X1 U11927 ( .A(P3_D_REG_21__SCAN_IN), .ZN(n9510) );
  NOR2_X1 U11928 ( .A1(n9499), .A2(n9510), .ZN(P3_U3244) );
  INV_X1 U11929 ( .A(P3_D_REG_18__SCAN_IN), .ZN(n9511) );
  NOR2_X1 U11930 ( .A1(n9525), .A2(n9511), .ZN(P3_U3247) );
  INV_X1 U11931 ( .A(P3_D_REG_8__SCAN_IN), .ZN(n9512) );
  NOR2_X1 U11932 ( .A1(n9525), .A2(n9512), .ZN(P3_U3257) );
  INV_X1 U11933 ( .A(P3_D_REG_9__SCAN_IN), .ZN(n13311) );
  NOR2_X1 U11934 ( .A1(n9525), .A2(n13311), .ZN(P3_U3256) );
  INV_X1 U11935 ( .A(P3_D_REG_10__SCAN_IN), .ZN(n9513) );
  NOR2_X1 U11936 ( .A1(n9525), .A2(n9513), .ZN(P3_U3255) );
  INV_X1 U11937 ( .A(P3_D_REG_26__SCAN_IN), .ZN(n9514) );
  NOR2_X1 U11938 ( .A1(n9499), .A2(n9514), .ZN(P3_U3239) );
  INV_X1 U11939 ( .A(P3_D_REG_12__SCAN_IN), .ZN(n9515) );
  NOR2_X1 U11940 ( .A1(n9525), .A2(n9515), .ZN(P3_U3253) );
  INV_X1 U11941 ( .A(P3_D_REG_25__SCAN_IN), .ZN(n9516) );
  NOR2_X1 U11942 ( .A1(n9499), .A2(n9516), .ZN(P3_U3240) );
  INV_X1 U11943 ( .A(P3_D_REG_11__SCAN_IN), .ZN(n9517) );
  NOR2_X1 U11944 ( .A1(n9525), .A2(n9517), .ZN(P3_U3254) );
  INV_X1 U11945 ( .A(P3_D_REG_30__SCAN_IN), .ZN(n13318) );
  NOR2_X1 U11946 ( .A1(n9499), .A2(n13318), .ZN(P3_U3235) );
  INV_X1 U11947 ( .A(P3_D_REG_16__SCAN_IN), .ZN(n9518) );
  NOR2_X1 U11948 ( .A1(n9525), .A2(n9518), .ZN(P3_U3249) );
  INV_X1 U11949 ( .A(P3_D_REG_2__SCAN_IN), .ZN(n9519) );
  NOR2_X1 U11950 ( .A1(n9525), .A2(n9519), .ZN(P3_U3263) );
  INV_X1 U11951 ( .A(P3_D_REG_17__SCAN_IN), .ZN(n9520) );
  NOR2_X1 U11952 ( .A1(n9525), .A2(n9520), .ZN(P3_U3248) );
  INV_X1 U11953 ( .A(P3_D_REG_4__SCAN_IN), .ZN(n9521) );
  NOR2_X1 U11954 ( .A1(n9525), .A2(n9521), .ZN(P3_U3261) );
  INV_X1 U11955 ( .A(P3_D_REG_31__SCAN_IN), .ZN(n9522) );
  NOR2_X1 U11956 ( .A1(n9499), .A2(n9522), .ZN(P3_U3234) );
  INV_X1 U11957 ( .A(P3_D_REG_7__SCAN_IN), .ZN(n9523) );
  NOR2_X1 U11958 ( .A1(n9525), .A2(n9523), .ZN(P3_U3258) );
  INV_X1 U11959 ( .A(P3_D_REG_22__SCAN_IN), .ZN(n9524) );
  NOR2_X1 U11960 ( .A1(n9525), .A2(n9524), .ZN(P3_U3243) );
  INV_X1 U11961 ( .A(P3_D_REG_6__SCAN_IN), .ZN(n13277) );
  NOR2_X1 U11962 ( .A1(n9525), .A2(n13277), .ZN(P3_U3259) );
  INV_X1 U11963 ( .A(P3_D_REG_23__SCAN_IN), .ZN(n9526) );
  NOR2_X1 U11964 ( .A1(n9525), .A2(n9526), .ZN(P3_U3242) );
  INV_X1 U11965 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n9528) );
  INV_X1 U11966 ( .A(n9567), .ZN(n9544) );
  OAI222_X1 U11967 ( .A1(n14038), .A2(n9528), .B1(n14031), .B2(n9527), .C1(
        P2_U3088), .C2(n9544), .ZN(P2_U3317) );
  AOI21_X1 U11968 ( .B1(n9535), .B2(P2_REG2_REG_8__SCAN_IN), .A(n9529), .ZN(
        n13602) );
  INV_X1 U11969 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n13597) );
  MUX2_X1 U11970 ( .A(n13597), .B(P2_REG2_REG_9__SCAN_IN), .S(n9537), .Z(n9530) );
  NAND2_X1 U11971 ( .A1(n9537), .A2(n13597), .ZN(n13601) );
  INV_X1 U11972 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n9531) );
  MUX2_X1 U11973 ( .A(n9531), .B(P2_REG2_REG_10__SCAN_IN), .S(n9567), .Z(n9532) );
  AOI211_X1 U11974 ( .C1(n9533), .C2(n9532), .A(n15442), .B(n9562), .ZN(n9547)
         );
  INV_X1 U11975 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n15571) );
  AOI21_X1 U11976 ( .B1(n9535), .B2(P2_REG1_REG_8__SCAN_IN), .A(n9534), .ZN(
        n13606) );
  MUX2_X1 U11977 ( .A(n15571), .B(P2_REG1_REG_9__SCAN_IN), .S(n9537), .Z(n9536) );
  AND2_X1 U11978 ( .A1(n13606), .A2(n9536), .ZN(n13607) );
  AOI21_X1 U11979 ( .B1(n15571), .B2(n9537), .A(n13607), .ZN(n9539) );
  INV_X1 U11980 ( .A(n9539), .ZN(n9542) );
  INV_X1 U11981 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n15574) );
  MUX2_X1 U11982 ( .A(n15574), .B(P2_REG1_REG_10__SCAN_IN), .S(n9567), .Z(
        n9541) );
  MUX2_X1 U11983 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n15574), .S(n9567), .Z(
        n9538) );
  NAND2_X1 U11984 ( .A1(n9539), .A2(n9538), .ZN(n9588) );
  INV_X1 U11985 ( .A(n9588), .ZN(n9540) );
  AOI211_X1 U11986 ( .C1(n9542), .C2(n9541), .A(n15459), .B(n9540), .ZN(n9546)
         );
  NAND2_X1 U11987 ( .A1(P2_U3088), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n10906)
         );
  NAND2_X1 U11988 ( .A1(n15472), .A2(P2_ADDR_REG_10__SCAN_IN), .ZN(n9543) );
  OAI211_X1 U11989 ( .C1(n15479), .C2(n9544), .A(n10906), .B(n9543), .ZN(n9545) );
  OR3_X1 U11990 ( .A1(n9547), .A2(n9546), .A3(n9545), .ZN(P2_U3224) );
  INV_X1 U11991 ( .A(n11281), .ZN(n9552) );
  INV_X1 U11992 ( .A(n9568), .ZN(n9582) );
  OAI222_X1 U11993 ( .A1(n14038), .A2(n9548), .B1(n14031), .B2(n9552), .C1(
        P2_U3088), .C2(n9582), .ZN(P2_U3316) );
  NOR2_X1 U11994 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n9549) );
  NAND2_X1 U11995 ( .A1(n9550), .A2(n9549), .ZN(n9689) );
  NAND2_X1 U11996 ( .A1(n9689), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9551) );
  XNOR2_X1 U11997 ( .A(n9551), .B(P1_IR_REG_11__SCAN_IN), .ZN(n11282) );
  INV_X1 U11998 ( .A(n11282), .ZN(n10061) );
  OAI222_X1 U11999 ( .A1(n14817), .A2(n9553), .B1(n14815), .B2(n9552), .C1(
        P1_U3086), .C2(n10061), .ZN(P1_U3344) );
  NAND2_X1 U12000 ( .A1(n9554), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9555) );
  XNOR2_X2 U12001 ( .A(n9558), .B(P1_IR_REG_30__SCAN_IN), .ZN(n9619) );
  INV_X2 U12002 ( .A(n10116), .ZN(n12112) );
  AOI222_X1 U12003 ( .A1(n12112), .A2(P1_REG1_REG_30__SCAN_IN), .B1(n12113), 
        .B2(P1_REG2_REG_30__SCAN_IN), .C1(n11808), .C2(P1_REG0_REG_30__SCAN_IN), .ZN(n14408) );
  INV_X1 U12004 ( .A(P1_U4016), .ZN(n14215) );
  NAND2_X1 U12005 ( .A1(n14215), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n9559) );
  OAI21_X1 U12006 ( .B1(n14408), .B2(n14215), .A(n9559), .ZN(P1_U3590) );
  OAI222_X1 U12007 ( .A1(P3_U3151), .A2(n15032), .B1(n14936), .B2(n9561), .C1(
        n14938), .C2(n9560), .ZN(P3_U3280) );
  INV_X1 U12008 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n9563) );
  MUX2_X1 U12009 ( .A(P2_REG2_REG_11__SCAN_IN), .B(n9563), .S(n9568), .Z(n9577) );
  NAND2_X1 U12010 ( .A1(n9576), .A2(n9577), .ZN(n9578) );
  NAND2_X1 U12011 ( .A1(n9582), .A2(n9563), .ZN(n9564) );
  INV_X1 U12012 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n10172) );
  MUX2_X1 U12013 ( .A(n10172), .B(P2_REG2_REG_12__SCAN_IN), .S(n10178), .Z(
        n9565) );
  AOI21_X1 U12014 ( .B1(n9578), .B2(n9564), .A(n9565), .ZN(n10170) );
  AND3_X1 U12015 ( .A1(n9578), .A2(n9565), .A3(n9564), .ZN(n9566) );
  OAI21_X1 U12016 ( .B1(n10170), .B2(n9566), .A(n15474), .ZN(n9575) );
  NAND2_X1 U12017 ( .A1(n9567), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n9587) );
  INV_X1 U12018 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n11239) );
  MUX2_X1 U12019 ( .A(n11239), .B(P2_REG1_REG_11__SCAN_IN), .S(n9568), .Z(
        n9586) );
  AOI21_X1 U12020 ( .B1(n9588), .B2(n9587), .A(n9586), .ZN(n9585) );
  AOI21_X1 U12021 ( .B1(n9568), .B2(P2_REG1_REG_11__SCAN_IN), .A(n9585), .ZN(
        n9570) );
  INV_X1 U12022 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n15157) );
  MUX2_X1 U12023 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n15157), .S(n10178), .Z(
        n9569) );
  NAND2_X1 U12024 ( .A1(n9570), .A2(n9569), .ZN(n10177) );
  OAI21_X1 U12025 ( .B1(n9570), .B2(n9569), .A(n10177), .ZN(n9573) );
  INV_X1 U12026 ( .A(n10178), .ZN(n10171) );
  NAND2_X1 U12027 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3088), .ZN(n11185)
         );
  NAND2_X1 U12028 ( .A1(n15472), .A2(P2_ADDR_REG_12__SCAN_IN), .ZN(n9571) );
  OAI211_X1 U12029 ( .C1(n15479), .C2(n10171), .A(n11185), .B(n9571), .ZN(
        n9572) );
  AOI21_X1 U12030 ( .B1(n9573), .B2(n15467), .A(n9572), .ZN(n9574) );
  NAND2_X1 U12031 ( .A1(n9575), .A2(n9574), .ZN(P2_U3226) );
  INV_X1 U12032 ( .A(n9576), .ZN(n9581) );
  INV_X1 U12033 ( .A(n9577), .ZN(n9580) );
  INV_X1 U12034 ( .A(n9578), .ZN(n9579) );
  AOI21_X1 U12035 ( .B1(n9581), .B2(n9580), .A(n9579), .ZN(n9593) );
  NOR2_X1 U12036 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8783), .ZN(n9584) );
  NOR2_X1 U12037 ( .A1(n15479), .A2(n9582), .ZN(n9583) );
  AOI211_X1 U12038 ( .C1(n15472), .C2(P2_ADDR_REG_11__SCAN_IN), .A(n9584), .B(
        n9583), .ZN(n9592) );
  INV_X1 U12039 ( .A(n9585), .ZN(n9590) );
  NAND3_X1 U12040 ( .A1(n9588), .A2(n9587), .A3(n9586), .ZN(n9589) );
  NAND3_X1 U12041 ( .A1(n9590), .A2(n15467), .A3(n9589), .ZN(n9591) );
  OAI211_X1 U12042 ( .C1(n9593), .C2(n15442), .A(n9592), .B(n9591), .ZN(
        P2_U3225) );
  INV_X1 U12043 ( .A(n11287), .ZN(n9690) );
  OAI222_X1 U12044 ( .A1(n14031), .A2(n9690), .B1(n10171), .B2(P2_U3088), .C1(
        n9594), .C2(n14038), .ZN(P2_U3315) );
  NOR4_X1 U12045 ( .A1(P1_D_REG_14__SCAN_IN), .A2(P1_D_REG_15__SCAN_IN), .A3(
        P1_D_REG_16__SCAN_IN), .A4(P1_D_REG_18__SCAN_IN), .ZN(n9599) );
  NOR4_X1 U12046 ( .A1(P1_D_REG_12__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_9__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n9598) );
  NOR4_X1 U12047 ( .A1(P1_D_REG_24__SCAN_IN), .A2(P1_D_REG_25__SCAN_IN), .A3(
        P1_D_REG_26__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n9597) );
  NOR4_X1 U12048 ( .A1(P1_D_REG_19__SCAN_IN), .A2(P1_D_REG_21__SCAN_IN), .A3(
        P1_D_REG_22__SCAN_IN), .A4(P1_D_REG_23__SCAN_IN), .ZN(n9596) );
  AND4_X1 U12049 ( .A1(n9599), .A2(n9598), .A3(n9597), .A4(n9596), .ZN(n9605)
         );
  NOR2_X1 U12050 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_17__SCAN_IN), .ZN(
        n9603) );
  NOR4_X1 U12051 ( .A1(P1_D_REG_27__SCAN_IN), .A2(P1_D_REG_28__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_11__SCAN_IN), .ZN(n9602) );
  NOR4_X1 U12052 ( .A1(P1_D_REG_3__SCAN_IN), .A2(P1_D_REG_4__SCAN_IN), .A3(
        P1_D_REG_5__SCAN_IN), .A4(P1_D_REG_6__SCAN_IN), .ZN(n9601) );
  NOR4_X1 U12053 ( .A1(P1_D_REG_30__SCAN_IN), .A2(P1_D_REG_29__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_2__SCAN_IN), .ZN(n9600) );
  AND4_X1 U12054 ( .A1(n9603), .A2(n9602), .A3(n9601), .A4(n9600), .ZN(n9604)
         );
  NAND2_X1 U12055 ( .A1(n9605), .A2(n9604), .ZN(n9756) );
  NOR2_X1 U12056 ( .A1(n9756), .A2(n9606), .ZN(n9607) );
  OAI21_X1 U12057 ( .B1(n9755), .B2(n9607), .A(n9754), .ZN(n9626) );
  NAND2_X1 U12058 ( .A1(n9608), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9609) );
  NAND2_X1 U12059 ( .A1(n9612), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9613) );
  OAI21_X1 U12060 ( .B1(n9760), .B2(n9626), .A(n9974), .ZN(n10694) );
  AND2_X1 U12061 ( .A1(n10694), .A2(n9975), .ZN(n14159) );
  NAND2_X1 U12062 ( .A1(n12130), .A2(n7108), .ZN(n9629) );
  INV_X1 U12063 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n14247) );
  OAI21_X1 U12064 ( .B1(n9616), .B2(n9615), .A(n9614), .ZN(n9617) );
  NAND2_X1 U12065 ( .A1(n9618), .A2(n9617), .ZN(n14819) );
  MUX2_X1 U12066 ( .A(n14247), .B(n14819), .S(n9817), .Z(n10225) );
  NAND2_X1 U12067 ( .A1(n11839), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n9621) );
  AND2_X2 U12068 ( .A1(n11832), .A2(n15320), .ZN(n10688) );
  OAI22_X1 U12069 ( .A1(n10225), .A2(n7915), .B1(n14247), .B2(n9630), .ZN(
        n9622) );
  AOI21_X1 U12070 ( .B1(n14230), .B2(n10688), .A(n9622), .ZN(n9823) );
  NAND2_X1 U12071 ( .A1(n14230), .A2(n6664), .ZN(n9625) );
  INV_X1 U12072 ( .A(n10225), .ZN(n10203) );
  AOI22_X1 U12073 ( .A1(n10203), .A2(n11832), .B1(P1_REG1_REG_0__SCAN_IN), 
        .B2(n9623), .ZN(n9624) );
  NAND2_X1 U12074 ( .A1(n9625), .A2(n9624), .ZN(n9822) );
  XNOR2_X1 U12075 ( .A(n9823), .B(n9822), .ZN(n14246) );
  INV_X1 U12076 ( .A(n9760), .ZN(n9972) );
  INV_X1 U12077 ( .A(n12134), .ZN(n9627) );
  AND2_X1 U12078 ( .A1(n15366), .A2(n9627), .ZN(n9628) );
  NAND2_X1 U12079 ( .A1(n14246), .A2(n14195), .ZN(n9637) );
  NAND2_X1 U12080 ( .A1(n12134), .A2(n9629), .ZN(n9633) );
  AND2_X1 U12081 ( .A1(n9631), .A2(n9630), .ZN(n9632) );
  AND2_X1 U12082 ( .A1(n9633), .A2(n9632), .ZN(n10693) );
  AND3_X1 U12083 ( .A1(n12186), .A2(n9972), .A3(n9772), .ZN(n14115) );
  NAND2_X1 U12084 ( .A1(n12134), .A2(n14807), .ZN(n14607) );
  NOR2_X1 U12085 ( .A1(n14200), .A2(n14607), .ZN(n14207) );
  NAND2_X1 U12086 ( .A1(n10117), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n9635) );
  NAND2_X1 U12087 ( .A1(n9986), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n9634) );
  NAND2_X1 U12088 ( .A1(n10694), .A2(n12186), .ZN(n10012) );
  AOI22_X1 U12089 ( .A1(n14207), .A2(n14229), .B1(P1_REG3_REG_0__SCAN_IN), 
        .B2(n10012), .ZN(n9636) );
  OAI211_X1 U12090 ( .C1(n14191), .C2(n10225), .A(n9637), .B(n9636), .ZN(
        P1_U3232) );
  NAND2_X1 U12091 ( .A1(n9641), .A2(n9642), .ZN(n9638) );
  NAND2_X1 U12092 ( .A1(n9639), .A2(n9638), .ZN(n9640) );
  NAND2_X4 U12093 ( .A1(n9794), .A2(n9641), .ZN(n13107) );
  NOR2_X2 U12094 ( .A1(n9642), .A2(n9176), .ZN(n10073) );
  NAND2_X1 U12095 ( .A1(n13577), .A2(n11865), .ZN(n9692) );
  NAND2_X1 U12096 ( .A1(n10624), .A2(n9795), .ZN(n9643) );
  NAND2_X1 U12097 ( .A1(n9685), .A2(n9643), .ZN(n9647) );
  INV_X1 U12098 ( .A(n9695), .ZN(n9646) );
  AOI21_X1 U12099 ( .B1(n9648), .B2(n9647), .A(n9646), .ZN(n9682) );
  INV_X1 U12100 ( .A(n9649), .ZN(n14036) );
  XNOR2_X1 U12101 ( .A(n11511), .B(P2_B_REG_SCAN_IN), .ZN(n9650) );
  NAND2_X1 U12102 ( .A1(n14036), .A2(n9650), .ZN(n9652) );
  INV_X1 U12103 ( .A(n14033), .ZN(n9651) );
  AND2_X1 U12104 ( .A1(n9652), .A2(n9651), .ZN(n15480) );
  INV_X1 U12105 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n15487) );
  AND2_X1 U12106 ( .A1(n11511), .A2(n14033), .ZN(n9653) );
  AOI21_X1 U12107 ( .B1(n15480), .B2(n15487), .A(n9653), .ZN(n9778) );
  NOR4_X1 U12108 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_21__SCAN_IN), .ZN(n9657) );
  NOR4_X1 U12109 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_13__SCAN_IN), .A3(
        P2_D_REG_14__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n9656) );
  NOR4_X1 U12110 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_29__SCAN_IN), .ZN(n9655) );
  NOR4_X1 U12111 ( .A1(P2_D_REG_22__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n9654) );
  NAND4_X1 U12112 ( .A1(n9657), .A2(n9656), .A3(n9655), .A4(n9654), .ZN(n9663)
         );
  NOR2_X1 U12113 ( .A1(P2_D_REG_8__SCAN_IN), .A2(P2_D_REG_17__SCAN_IN), .ZN(
        n9661) );
  NOR4_X1 U12114 ( .A1(P2_D_REG_31__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_7__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n9660) );
  NOR4_X1 U12115 ( .A1(P2_D_REG_9__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_11__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n9659) );
  NOR4_X1 U12116 ( .A1(P2_D_REG_3__SCAN_IN), .A2(P2_D_REG_4__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_6__SCAN_IN), .ZN(n9658) );
  NAND4_X1 U12117 ( .A1(n9661), .A2(n9660), .A3(n9659), .A4(n9658), .ZN(n9662)
         );
  OAI21_X1 U12118 ( .B1(n9663), .B2(n9662), .A(n15480), .ZN(n9780) );
  NAND2_X1 U12119 ( .A1(n9778), .A2(n9780), .ZN(n9898) );
  INV_X1 U12120 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n15489) );
  NAND2_X1 U12121 ( .A1(n15480), .A2(n15489), .ZN(n9665) );
  NAND2_X1 U12122 ( .A1(n14036), .A2(n14033), .ZN(n9664) );
  NAND2_X1 U12123 ( .A1(n9665), .A2(n9664), .ZN(n15490) );
  OR2_X1 U12124 ( .A1(n9898), .A2(n15490), .ZN(n9676) );
  INV_X1 U12125 ( .A(n9676), .ZN(n9666) );
  NAND2_X1 U12126 ( .A1(n9666), .A2(n15491), .ZN(n9677) );
  INV_X1 U12127 ( .A(n9672), .ZN(n9668) );
  NAND2_X1 U12128 ( .A1(n15548), .A2(n9668), .ZN(n9669) );
  INV_X1 U12129 ( .A(n9677), .ZN(n9671) );
  INV_X1 U12130 ( .A(n13578), .ZN(n9683) );
  INV_X1 U12131 ( .A(n13576), .ZN(n9905) );
  NAND2_X1 U12132 ( .A1(n9672), .A2(n9288), .ZN(n13630) );
  OAI22_X1 U12133 ( .A1(n9683), .A2(n13496), .B1(n9905), .B2(n13630), .ZN(
        n10301) );
  NAND2_X1 U12134 ( .A1(n9674), .A2(n10983), .ZN(n9782) );
  AOI21_X1 U12135 ( .B1(n9676), .B2(n9782), .A(n9897), .ZN(n9946) );
  NAND2_X1 U12136 ( .A1(n9946), .A2(n15491), .ZN(n9699) );
  AOI22_X1 U12137 ( .A1(n15125), .A2(n10301), .B1(n9699), .B2(
        P2_REG3_REG_1__SCAN_IN), .ZN(n9681) );
  NAND2_X1 U12138 ( .A1(n10073), .A2(n9247), .ZN(n10250) );
  OR2_X1 U12139 ( .A1(n9677), .A2(n10250), .ZN(n9679) );
  NAND2_X1 U12140 ( .A1(n15128), .A2(n6672), .ZN(n9680) );
  OAI211_X1 U12141 ( .C1(n9682), .C2(n13561), .A(n9681), .B(n9680), .ZN(
        P2_U3194) );
  INV_X1 U12142 ( .A(n13577), .ZN(n9784) );
  NOR2_X1 U12143 ( .A1(n9784), .A2(n13630), .ZN(n10074) );
  INV_X1 U12144 ( .A(n10074), .ZN(n9688) );
  AOI22_X1 U12145 ( .A1(n15128), .A2(n10295), .B1(P2_REG3_REG_0__SCAN_IN), 
        .B2(n9699), .ZN(n9687) );
  OAI21_X1 U12146 ( .B1(n9683), .B2(n15144), .A(n9795), .ZN(n9684) );
  NAND3_X1 U12147 ( .A1(n15123), .A2(n9685), .A3(n9684), .ZN(n9686) );
  OAI211_X1 U12148 ( .C1(n9688), .C2(n13558), .A(n9687), .B(n9686), .ZN(
        P2_U3204) );
  NAND2_X1 U12149 ( .A1(n10051), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9702) );
  XNOR2_X1 U12150 ( .A(n9702), .B(P1_IR_REG_12__SCAN_IN), .ZN(n11288) );
  INV_X1 U12151 ( .A(n11288), .ZN(n10065) );
  OAI222_X1 U12152 ( .A1(n14817), .A2(n9691), .B1(n14815), .B2(n9690), .C1(
        n10065), .C2(P1_U3086), .ZN(P1_U3343) );
  INV_X1 U12153 ( .A(n11445), .ZN(n9706) );
  INV_X1 U12154 ( .A(n15454), .ZN(n10174) );
  OAI222_X1 U12155 ( .A1(n14031), .A2(n9706), .B1(n10174), .B2(P2_U3088), .C1(
        n6979), .C2(n14038), .ZN(P2_U3314) );
  NAND2_X1 U12156 ( .A1(n13576), .A2(n11865), .ZN(n9932) );
  XNOR2_X1 U12157 ( .A(n9931), .B(n9932), .ZN(n9697) );
  NAND2_X1 U12158 ( .A1(n9693), .A2(n9692), .ZN(n9694) );
  OAI21_X1 U12159 ( .B1(n9697), .B2(n9696), .A(n9935), .ZN(n9698) );
  NAND2_X1 U12160 ( .A1(n9698), .A2(n15123), .ZN(n9701) );
  INV_X1 U12161 ( .A(n13575), .ZN(n9961) );
  OAI22_X1 U12162 ( .A1(n9961), .A2(n13630), .B1(n9784), .B2(n13496), .ZN(
        n9788) );
  AOI22_X1 U12163 ( .A1(n15125), .A2(n9788), .B1(n9699), .B2(
        P2_REG3_REG_2__SCAN_IN), .ZN(n9700) );
  OAI211_X1 U12164 ( .C1(n10668), .C2(n13542), .A(n9701), .B(n9700), .ZN(
        P2_U3209) );
  NAND2_X1 U12165 ( .A1(n9702), .A2(n10048), .ZN(n9703) );
  NAND2_X1 U12166 ( .A1(n9703), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9704) );
  NAND2_X1 U12167 ( .A1(n9704), .A2(n10049), .ZN(n9811) );
  OR2_X1 U12168 ( .A1(n9704), .A2(n10049), .ZN(n9705) );
  INV_X1 U12169 ( .A(n11446), .ZN(n10504) );
  OAI222_X1 U12170 ( .A1(n14817), .A2(n9707), .B1(n14815), .B2(n9706), .C1(
        n10504), .C2(P1_U3086), .ZN(P1_U3342) );
  INV_X1 U12171 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n9708) );
  MUX2_X1 U12172 ( .A(n9708), .B(P1_REG1_REG_8__SCAN_IN), .S(n10829), .Z(n9718) );
  INV_X1 U12173 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n15396) );
  INV_X1 U12174 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n15390) );
  MUX2_X1 U12175 ( .A(n15390), .B(P1_REG1_REG_1__SCAN_IN), .S(n14234), .Z(
        n14236) );
  INV_X1 U12176 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n9709) );
  AOI21_X1 U12177 ( .B1(n14234), .B2(P1_REG1_REG_1__SCAN_IN), .A(n14235), .ZN(
        n14255) );
  INV_X1 U12178 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n15392) );
  NAND2_X1 U12179 ( .A1(n14258), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n14269) );
  INV_X1 U12180 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n10222) );
  MUX2_X1 U12181 ( .A(n10222), .B(P1_REG1_REG_3__SCAN_IN), .S(n14265), .Z(
        n14268) );
  NOR2_X1 U12182 ( .A1(n9710), .A2(n10222), .ZN(n14278) );
  INV_X1 U12183 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n9711) );
  MUX2_X1 U12184 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n9711), .S(n14284), .Z(n9712) );
  OAI21_X1 U12185 ( .B1(n14283), .B2(n14278), .A(n9712), .ZN(n14281) );
  INV_X1 U12186 ( .A(n14281), .ZN(n9713) );
  MUX2_X1 U12187 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n6957), .S(n14299), .Z(
        n14297) );
  INV_X1 U12188 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n15394) );
  MUX2_X1 U12189 ( .A(n15394), .B(P1_REG1_REG_6__SCAN_IN), .S(n10436), .Z(
        n9888) );
  NOR2_X1 U12190 ( .A1(n9714), .A2(n15394), .ZN(n14308) );
  MUX2_X1 U12191 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n15396), .S(n14317), .Z(
        n9715) );
  OAI21_X1 U12192 ( .B1(n14313), .B2(n14308), .A(n9715), .ZN(n14311) );
  AOI21_X1 U12193 ( .B1(n9718), .B2(n9717), .A(n14329), .ZN(n9753) );
  INV_X1 U12194 ( .A(n9719), .ZN(n9720) );
  NAND2_X1 U12195 ( .A1(n9721), .A2(n9720), .ZN(n9727) );
  INV_X1 U12196 ( .A(n9727), .ZN(n9809) );
  AND2_X1 U12197 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n9725) );
  INV_X1 U12198 ( .A(n14807), .ZN(n9834) );
  OR2_X1 U12199 ( .A1(n9727), .A2(n9834), .ZN(n15267) );
  NOR2_X1 U12200 ( .A1(n15267), .A2(n9723), .ZN(n9724) );
  AOI211_X1 U12201 ( .C1(n14360), .C2(P1_ADDR_REG_8__SCAN_IN), .A(n9725), .B(
        n9724), .ZN(n9752) );
  NAND2_X1 U12203 ( .A1(n9834), .A2(n6667), .ZN(n9726) );
  INV_X1 U12204 ( .A(n15266), .ZN(n14377) );
  XNOR2_X1 U12205 ( .A(n14258), .B(P1_REG2_REG_2__SCAN_IN), .ZN(n14252) );
  INV_X1 U12206 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n9728) );
  MUX2_X1 U12207 ( .A(P1_REG2_REG_1__SCAN_IN), .B(n9728), .S(n14234), .Z(
        n14240) );
  AND2_X1 U12208 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n9729) );
  NAND2_X1 U12209 ( .A1(n14240), .A2(n9729), .ZN(n14239) );
  NAND2_X1 U12210 ( .A1(n14234), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n9730) );
  NAND2_X1 U12211 ( .A1(n14239), .A2(n9730), .ZN(n14251) );
  INV_X1 U12212 ( .A(n14251), .ZN(n9731) );
  OR2_X1 U12213 ( .A1(n14252), .A2(n9731), .ZN(n9733) );
  NAND2_X1 U12214 ( .A1(n14258), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n9732) );
  NAND2_X1 U12215 ( .A1(n9733), .A2(n9732), .ZN(n14266) );
  INV_X1 U12216 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n10191) );
  MUX2_X1 U12217 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n10191), .S(n14265), .Z(
        n14267) );
  NAND2_X1 U12218 ( .A1(n14266), .A2(n14267), .ZN(n14287) );
  NAND2_X1 U12219 ( .A1(n14265), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n14286) );
  NAND2_X1 U12220 ( .A1(n14287), .A2(n14286), .ZN(n9736) );
  INV_X1 U12221 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n9734) );
  MUX2_X1 U12222 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n9734), .S(n14284), .Z(n9735) );
  NAND2_X1 U12223 ( .A1(n9736), .A2(n9735), .ZN(n14302) );
  NAND2_X1 U12224 ( .A1(n14284), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n14301) );
  NAND2_X1 U12225 ( .A1(n14302), .A2(n14301), .ZN(n9739) );
  INV_X1 U12226 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n9737) );
  MUX2_X1 U12227 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n9737), .S(n14299), .Z(n9738) );
  NAND2_X1 U12228 ( .A1(n9739), .A2(n9738), .ZN(n14304) );
  NAND2_X1 U12229 ( .A1(n14299), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n9891) );
  NAND2_X1 U12230 ( .A1(n14304), .A2(n9891), .ZN(n9741) );
  INV_X1 U12231 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n10446) );
  MUX2_X1 U12232 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n10446), .S(n10436), .Z(
        n9740) );
  NAND2_X1 U12233 ( .A1(n9741), .A2(n9740), .ZN(n14320) );
  NAND2_X1 U12234 ( .A1(n10436), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n14319) );
  NAND2_X1 U12235 ( .A1(n14320), .A2(n14319), .ZN(n9744) );
  INV_X1 U12236 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n9742) );
  MUX2_X1 U12237 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n9742), .S(n14317), .Z(n9743) );
  NAND2_X1 U12238 ( .A1(n9744), .A2(n9743), .ZN(n14322) );
  NAND2_X1 U12239 ( .A1(n14317), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n9749) );
  NAND2_X1 U12240 ( .A1(n14322), .A2(n9749), .ZN(n9747) );
  INV_X1 U12241 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n9745) );
  MUX2_X1 U12242 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n9745), .S(n10829), .Z(n9746) );
  NAND2_X1 U12243 ( .A1(n9747), .A2(n9746), .ZN(n14336) );
  MUX2_X1 U12244 ( .A(n9745), .B(P1_REG2_REG_8__SCAN_IN), .S(n10829), .Z(n9748) );
  NAND3_X1 U12245 ( .A1(n14322), .A2(n9749), .A3(n9748), .ZN(n9750) );
  NAND3_X1 U12246 ( .A1(n14377), .A2(n14336), .A3(n9750), .ZN(n9751) );
  OAI211_X1 U12247 ( .C1(n9753), .C2(n15264), .A(n9752), .B(n9751), .ZN(
        P1_U3251) );
  OAI21_X1 U12248 ( .B1(n9755), .B2(P1_D_REG_0__SCAN_IN), .A(n9754), .ZN(n9759) );
  INV_X1 U12249 ( .A(n9755), .ZN(n9757) );
  NAND2_X1 U12250 ( .A1(n9757), .A2(n9756), .ZN(n9758) );
  AND3_X1 U12251 ( .A1(n12186), .A2(n9759), .A3(n9758), .ZN(n9973) );
  INV_X1 U12252 ( .A(n9996), .ZN(n9770) );
  OR2_X1 U12253 ( .A1(n12131), .A2(n7108), .ZN(n9762) );
  OR2_X1 U12254 ( .A1(n12141), .A2(n12130), .ZN(n9761) );
  INV_X1 U12255 ( .A(n11951), .ZN(n9764) );
  NAND2_X1 U12256 ( .A1(n9764), .A2(n10185), .ZN(n9765) );
  NAND2_X1 U12257 ( .A1(n11830), .A2(n9765), .ZN(n9977) );
  AND2_X1 U12258 ( .A1(n12130), .A2(n14612), .ZN(n9766) );
  NAND2_X1 U12259 ( .A1(n12131), .A2(n9766), .ZN(n15341) );
  INV_X1 U12260 ( .A(n11953), .ZN(n9768) );
  NAND2_X1 U12261 ( .A1(n14230), .A2(n10225), .ZN(n9767) );
  NAND2_X1 U12262 ( .A1(n9768), .A2(n9767), .ZN(n12148) );
  OAI21_X1 U12263 ( .B1(n15375), .B2(n15386), .A(n12148), .ZN(n9769) );
  INV_X2 U12264 ( .A(n14607), .ZN(n14966) );
  NAND2_X1 U12265 ( .A1(n14229), .A2(n14966), .ZN(n10224) );
  OAI211_X1 U12266 ( .C1(n9770), .C2(n10225), .A(n9769), .B(n10224), .ZN(n9774) );
  NAND2_X1 U12267 ( .A1(n9774), .A2(n15389), .ZN(n9771) );
  OAI21_X1 U12268 ( .B1(n15389), .B2(n7501), .A(n9771), .ZN(P1_U3459) );
  AND3_X2 U12269 ( .A1(n9773), .A2(n12186), .A3(n9772), .ZN(n15403) );
  NAND2_X1 U12270 ( .A1(n9774), .A2(n15403), .ZN(n9775) );
  OAI21_X1 U12271 ( .B1(n15403), .B2(n9709), .A(n9775), .ZN(P1_U3528) );
  INV_X1 U12272 ( .A(n15042), .ZN(n12674) );
  INV_X1 U12273 ( .A(n9776), .ZN(n9777) );
  OAI222_X1 U12274 ( .A1(P3_U3151), .A2(n12674), .B1(n14936), .B2(n13466), 
        .C1(n14938), .C2(n9777), .ZN(P3_U3279) );
  NOR2_X1 U12275 ( .A1(n9778), .A2(n15488), .ZN(n15486) );
  INV_X1 U12276 ( .A(n9897), .ZN(n9779) );
  AND2_X1 U12277 ( .A1(n9780), .A2(n9779), .ZN(n9781) );
  AND2_X1 U12278 ( .A1(n15486), .A2(n9781), .ZN(n10071) );
  AND2_X1 U12279 ( .A1(n15491), .A2(n9782), .ZN(n9783) );
  INV_X2 U12280 ( .A(n15559), .ZN(n15561) );
  INV_X1 U12281 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n9801) );
  NOR2_X1 U12282 ( .A1(n13578), .A2(n9795), .ZN(n10300) );
  NAND2_X1 U12283 ( .A1(n10299), .A2(n10300), .ZN(n10298) );
  NAND2_X1 U12284 ( .A1(n9784), .A2(n6672), .ZN(n9785) );
  XNOR2_X1 U12285 ( .A(n9902), .B(n9901), .ZN(n9789) );
  NOR2_X1 U12286 ( .A1(n10983), .A2(n6670), .ZN(n9786) );
  NOR2_X2 U12287 ( .A1(n9787), .A2(n9786), .ZN(n15522) );
  AOI21_X1 U12288 ( .B1(n9789), .B2(n15551), .A(n9788), .ZN(n10673) );
  OAI22_X1 U12289 ( .A1(n10299), .A2(n9790), .B1(n6672), .B2(n13577), .ZN(
        n9792) );
  INV_X1 U12290 ( .A(n9901), .ZN(n9791) );
  NAND2_X1 U12291 ( .A1(n9792), .A2(n9791), .ZN(n9907) );
  OR2_X1 U12292 ( .A1(n9792), .A2(n9791), .ZN(n9793) );
  NAND2_X1 U12293 ( .A1(n9907), .A2(n9793), .ZN(n10671) );
  NAND2_X1 U12294 ( .A1(n7362), .A2(n9795), .ZN(n10296) );
  NAND2_X1 U12295 ( .A1(n9796), .A2(n15144), .ZN(n9797) );
  OR2_X1 U12296 ( .A1(n9909), .A2(n9797), .ZN(n10665) );
  OAI21_X1 U12297 ( .B1(n10668), .B2(n15548), .A(n10665), .ZN(n9798) );
  AOI21_X1 U12298 ( .B1(n10671), .B2(n15527), .A(n9798), .ZN(n9799) );
  NAND2_X1 U12299 ( .A1(n10673), .A2(n9799), .ZN(n9954) );
  NAND2_X1 U12300 ( .A1(n9954), .A2(n15561), .ZN(n9800) );
  OAI21_X1 U12301 ( .B1(n15561), .B2(n9801), .A(n9800), .ZN(P2_U3436) );
  OAI222_X1 U12302 ( .A1(P3_U3151), .A2(n12699), .B1(n14936), .B2(n13439), 
        .C1(n14938), .C2(n9802), .ZN(P3_U3278) );
  INV_X1 U12303 ( .A(P3_DATAO_REG_3__SCAN_IN), .ZN(n13310) );
  NAND2_X1 U12304 ( .A1(n8394), .A2(n15577), .ZN(n9803) );
  OAI21_X1 U12305 ( .B1(n15577), .B2(n13310), .A(n9803), .ZN(P3_U3494) );
  INV_X1 U12306 ( .A(P3_DATAO_REG_1__SCAN_IN), .ZN(n13405) );
  NAND2_X1 U12307 ( .A1(n10318), .A2(n15577), .ZN(n9804) );
  OAI21_X1 U12308 ( .B1(n15577), .B2(n13405), .A(n9804), .ZN(P3_U3492) );
  OAI21_X1 U12309 ( .B1(P1_REG2_REG_0__SCAN_IN), .B2(n6668), .A(n9834), .ZN(
        n14248) );
  AOI21_X1 U12310 ( .B1(n9709), .B2(n6669), .A(n14248), .ZN(n9805) );
  MUX2_X1 U12311 ( .A(n14248), .B(n9805), .S(n14247), .Z(n9808) );
  INV_X1 U12312 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n10223) );
  OAI22_X1 U12313 ( .A1(n15271), .A2(n14877), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10223), .ZN(n9807) );
  NOR3_X1 U12314 ( .A1(n15264), .A2(n14247), .A3(P1_REG1_REG_0__SCAN_IN), .ZN(
        n9806) );
  AOI211_X1 U12315 ( .C1(n9809), .C2(n9808), .A(n9807), .B(n9806), .ZN(n9810)
         );
  INV_X1 U12316 ( .A(n9810), .ZN(P1_U3243) );
  INV_X1 U12317 ( .A(n11450), .ZN(n9814) );
  NAND2_X1 U12318 ( .A1(n9811), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9812) );
  INV_X1 U12319 ( .A(n11451), .ZN(n10954) );
  OAI222_X1 U12320 ( .A1(n14817), .A2(n9813), .B1(n14815), .B2(n9814), .C1(
        P1_U3086), .C2(n10954), .ZN(P1_U3341) );
  INV_X1 U12321 ( .A(n10865), .ZN(n10875) );
  OAI222_X1 U12322 ( .A1(n14038), .A2(n9815), .B1(n14031), .B2(n9814), .C1(
        P2_U3088), .C2(n10875), .ZN(P2_U3313) );
  NAND2_X1 U12323 ( .A1(n11657), .A2(n14234), .ZN(n9821) );
  NAND2_X1 U12324 ( .A1(n10128), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n9820) );
  OR2_X1 U12325 ( .A1(n12109), .A2(n9818), .ZN(n9819) );
  AND3_X2 U12326 ( .A1(n9821), .A2(n9820), .A3(n9819), .ZN(n15319) );
  MUX2_X1 U12327 ( .A(n11830), .B(n9823), .S(n9822), .Z(n9832) );
  NAND2_X1 U12328 ( .A1(n14229), .A2(n6664), .ZN(n9825) );
  NAND2_X1 U12329 ( .A1(n11960), .A2(n11832), .ZN(n9824) );
  XNOR2_X1 U12330 ( .A(n9826), .B(n11778), .ZN(n9829) );
  AND2_X1 U12331 ( .A1(n11960), .A2(n6664), .ZN(n9827) );
  AOI21_X1 U12332 ( .B1(n14229), .B2(n10688), .A(n9827), .ZN(n9828) );
  NAND2_X1 U12333 ( .A1(n9829), .A2(n9828), .ZN(n10007) );
  OR2_X1 U12334 ( .A1(n9829), .A2(n9828), .ZN(n9830) );
  OAI21_X1 U12335 ( .B1(n9832), .B2(n9831), .A(n10008), .ZN(n9833) );
  NAND2_X1 U12336 ( .A1(n9833), .A2(n14195), .ZN(n9842) );
  AND2_X2 U12337 ( .A1(n9834), .A2(n12134), .ZN(n15378) );
  NAND2_X1 U12338 ( .A1(n14115), .A2(n15378), .ZN(n15161) );
  INV_X1 U12339 ( .A(n15161), .ZN(n14063) );
  INV_X1 U12340 ( .A(n14207), .ZN(n15164) );
  NAND2_X1 U12341 ( .A1(n9986), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n9838) );
  NAND2_X1 U12342 ( .A1(n10117), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n9837) );
  NAND2_X1 U12343 ( .A1(n11088), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n9836) );
  NAND2_X1 U12344 ( .A1(n6658), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n9835) );
  INV_X1 U12345 ( .A(n6659), .ZN(n10201) );
  INV_X1 U12346 ( .A(n10012), .ZN(n9839) );
  INV_X1 U12347 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n14231) );
  OAI22_X1 U12348 ( .A1(n15164), .A2(n10201), .B1(n9839), .B2(n14231), .ZN(
        n9840) );
  AOI21_X1 U12349 ( .B1(n14063), .B2(n14230), .A(n9840), .ZN(n9841) );
  OAI211_X1 U12350 ( .C1(n15319), .C2(n14191), .A(n9842), .B(n9841), .ZN(
        P1_U3222) );
  NOR2_X1 U12351 ( .A1(n10829), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n14327) );
  INV_X1 U12352 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n15399) );
  MUX2_X1 U12353 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n15399), .S(n14339), .Z(
        n14328) );
  INV_X1 U12354 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n15401) );
  MUX2_X1 U12355 ( .A(n15401), .B(P1_REG1_REG_10__SCAN_IN), .S(n11072), .Z(
        n9921) );
  INV_X1 U12356 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n15227) );
  NOR3_X1 U12357 ( .A1(n9860), .A2(n15227), .A3(n15264), .ZN(n9851) );
  NAND2_X1 U12358 ( .A1(n10829), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n14335) );
  NAND2_X1 U12359 ( .A1(n14336), .A2(n14335), .ZN(n9845) );
  INV_X1 U12360 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n9843) );
  MUX2_X1 U12361 ( .A(P1_REG2_REG_9__SCAN_IN), .B(n9843), .S(n14339), .Z(n9844) );
  NAND2_X1 U12362 ( .A1(n9845), .A2(n9844), .ZN(n14338) );
  NAND2_X1 U12363 ( .A1(n14339), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n9846) );
  NAND2_X1 U12364 ( .A1(n14338), .A2(n9846), .ZN(n9926) );
  INV_X1 U12365 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n9847) );
  MUX2_X1 U12366 ( .A(P1_REG2_REG_10__SCAN_IN), .B(n9847), .S(n11072), .Z(
        n9925) );
  NAND2_X1 U12367 ( .A1(n9926), .A2(n9925), .ZN(n9924) );
  NAND2_X1 U12368 ( .A1(n11072), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n9848) );
  AND2_X1 U12369 ( .A1(n9924), .A2(n9848), .ZN(n9853) );
  INV_X1 U12370 ( .A(n9853), .ZN(n9849) );
  NOR3_X1 U12371 ( .A1(n9849), .A2(P1_REG2_REG_11__SCAN_IN), .A3(n15266), .ZN(
        n9850) );
  NOR3_X1 U12372 ( .A1(n9851), .A2(n14340), .A3(n9850), .ZN(n9864) );
  INV_X1 U12373 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n9857) );
  INV_X1 U12374 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n9854) );
  MUX2_X1 U12375 ( .A(n9854), .B(P1_REG2_REG_11__SCAN_IN), .S(n11282), .Z(
        n9852) );
  OAI21_X1 U12376 ( .B1(n11282), .B2(n9854), .A(n9853), .ZN(n9855) );
  NAND3_X1 U12377 ( .A1(n10056), .A2(n14377), .A3(n9855), .ZN(n9856) );
  NAND2_X1 U12378 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n14178)
         );
  OAI211_X1 U12379 ( .C1(n9857), .C2(n15271), .A(n9856), .B(n14178), .ZN(n9858) );
  INV_X1 U12380 ( .A(n9858), .ZN(n9863) );
  NOR3_X1 U12381 ( .A1(n9860), .A2(n11282), .A3(P1_REG1_REG_11__SCAN_IN), .ZN(
        n9861) );
  MUX2_X1 U12382 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n15227), .S(n11282), .Z(
        n9859) );
  OAI21_X1 U12383 ( .B1(n9861), .B2(n10060), .A(n14378), .ZN(n9862) );
  OAI211_X1 U12384 ( .C1(n9864), .C2(n10061), .A(n9863), .B(n9862), .ZN(
        P1_U3254) );
  INV_X1 U12385 ( .A(n9865), .ZN(n9866) );
  NAND2_X1 U12386 ( .A1(n9878), .A2(n9866), .ZN(n9871) );
  AND3_X1 U12387 ( .A1(n9868), .A2(n9867), .A3(n10019), .ZN(n9870) );
  NAND2_X1 U12388 ( .A1(n9879), .A2(n9872), .ZN(n9869) );
  NAND3_X1 U12389 ( .A1(n9871), .A2(n9870), .A3(n9869), .ZN(n10472) );
  NOR2_X1 U12390 ( .A1(n10472), .A2(P3_U3151), .ZN(n10487) );
  INV_X1 U12391 ( .A(P3_REG3_REG_0__SCAN_IN), .ZN(n9887) );
  NAND2_X1 U12392 ( .A1(n9872), .A2(n15744), .ZN(n9873) );
  OAI22_X1 U12393 ( .A1(n9878), .A2(n9874), .B1(n9879), .B2(n9873), .ZN(n9875)
         );
  INV_X1 U12394 ( .A(n15704), .ZN(n12441) );
  NAND2_X1 U12395 ( .A1(n12638), .A2(n9876), .ZN(n12436) );
  NAND2_X1 U12396 ( .A1(n12441), .A2(n12436), .ZN(n12416) );
  NAND2_X1 U12397 ( .A1(n12610), .A2(n12611), .ZN(n9877) );
  NOR2_X1 U12398 ( .A1(n15009), .A2(n15017), .ZN(n12347) );
  INV_X1 U12399 ( .A(n12347), .ZN(n12313) );
  INV_X1 U12400 ( .A(n9879), .ZN(n9881) );
  AND2_X1 U12401 ( .A1(n12610), .A2(n15770), .ZN(n9880) );
  NAND2_X1 U12402 ( .A1(n9881), .A2(n9880), .ZN(n9884) );
  INV_X1 U12403 ( .A(n15712), .ZN(n9882) );
  NOR2_X1 U12404 ( .A1(n15744), .A2(n9882), .ZN(n9883) );
  OAI22_X1 U12405 ( .A1(n12313), .A2(n7130), .B1(n9876), .B2(n15581), .ZN(
        n9885) );
  AOI21_X1 U12406 ( .B1(n15021), .B2(n12416), .A(n9885), .ZN(n9886) );
  OAI21_X1 U12407 ( .B1(n10487), .B2(n9887), .A(n9886), .ZN(P3_U3172) );
  AOI211_X1 U12408 ( .C1(n9889), .C2(n9888), .A(n15264), .B(n14313), .ZN(n9896) );
  MUX2_X1 U12409 ( .A(n10446), .B(P1_REG2_REG_6__SCAN_IN), .S(n10436), .Z(
        n9890) );
  NAND3_X1 U12410 ( .A1(n14304), .A2(n9891), .A3(n9890), .ZN(n9892) );
  AND3_X1 U12411 ( .A1(n14377), .A2(n14320), .A3(n9892), .ZN(n9895) );
  NAND2_X1 U12412 ( .A1(n14340), .A2(n10436), .ZN(n9893) );
  NAND2_X1 U12413 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n10947) );
  OAI211_X1 U12414 ( .C1(n14891), .C2(n15271), .A(n9893), .B(n10947), .ZN(
        n9894) );
  OR3_X1 U12415 ( .A1(n9896), .A2(n9895), .A3(n9894), .ZN(P1_U3249) );
  NOR2_X1 U12416 ( .A1(n9898), .A2(n9897), .ZN(n9900) );
  NAND2_X1 U12417 ( .A1(n9902), .A2(n9901), .ZN(n9904) );
  XNOR2_X1 U12418 ( .A(n9956), .B(n9958), .ZN(n10563) );
  NAND2_X1 U12419 ( .A1(n9905), .A2(n10668), .ZN(n9906) );
  NAND2_X1 U12420 ( .A1(n9907), .A2(n9906), .ZN(n9908) );
  NAND2_X1 U12421 ( .A1(n9908), .A2(n9956), .ZN(n9963) );
  OAI21_X1 U12422 ( .B1(n9908), .B2(n9956), .A(n9963), .ZN(n10560) );
  OR2_X1 U12423 ( .A1(n9909), .A2(n10556), .ZN(n9910) );
  AND3_X1 U12424 ( .A1(n9965), .A2(n15144), .A3(n9910), .ZN(n10559) );
  NAND2_X1 U12425 ( .A1(n13576), .A2(n13701), .ZN(n9912) );
  NAND2_X1 U12426 ( .A1(n13574), .A2(n13555), .ZN(n9911) );
  AND2_X1 U12427 ( .A1(n9912), .A2(n9911), .ZN(n10555) );
  OAI21_X1 U12428 ( .B1(n10556), .B2(n15548), .A(n10555), .ZN(n9913) );
  AOI211_X1 U12429 ( .C1(n10560), .C2(n15527), .A(n10559), .B(n9913), .ZN(
        n9914) );
  OAI21_X1 U12430 ( .B1(n15522), .B2(n10563), .A(n9914), .ZN(n9917) );
  NAND2_X1 U12431 ( .A1(n9917), .A2(n15576), .ZN(n9915) );
  OAI21_X1 U12432 ( .B1(n15576), .B2(n9916), .A(n9915), .ZN(P2_U3502) );
  INV_X1 U12433 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n9919) );
  NAND2_X1 U12434 ( .A1(n9917), .A2(n15561), .ZN(n9918) );
  OAI21_X1 U12435 ( .B1(n15561), .B2(n9919), .A(n9918), .ZN(P2_U3439) );
  AOI211_X1 U12436 ( .C1(n9922), .C2(n9921), .A(n15264), .B(n9920), .ZN(n9923)
         );
  AOI21_X1 U12437 ( .B1(n14340), .B2(n11072), .A(n9923), .ZN(n9930) );
  AND2_X1 U12438 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n11552) );
  OAI211_X1 U12439 ( .C1(n9926), .C2(n9925), .A(n14377), .B(n9924), .ZN(n9927)
         );
  OAI21_X1 U12440 ( .B1(n14862), .B2(n15271), .A(n9927), .ZN(n9928) );
  NOR2_X1 U12441 ( .A1(n11552), .A2(n9928), .ZN(n9929) );
  NAND2_X1 U12442 ( .A1(n9930), .A2(n9929), .ZN(P1_U3253) );
  XNOR2_X1 U12443 ( .A(n13107), .B(n10704), .ZN(n10155) );
  AND2_X1 U12444 ( .A1(n13574), .A2(n11865), .ZN(n10156) );
  XNOR2_X1 U12445 ( .A(n10155), .B(n10156), .ZN(n9944) );
  INV_X1 U12446 ( .A(n9931), .ZN(n9933) );
  NAND2_X1 U12447 ( .A1(n9933), .A2(n9932), .ZN(n9934) );
  AND2_X1 U12448 ( .A1(n13575), .A2(n11865), .ZN(n9937) );
  XNOR2_X1 U12449 ( .A(n13107), .B(n13094), .ZN(n9936) );
  NAND2_X1 U12450 ( .A1(n9937), .A2(n9936), .ZN(n9941) );
  INV_X1 U12451 ( .A(n9936), .ZN(n9939) );
  INV_X1 U12452 ( .A(n9937), .ZN(n9938) );
  NAND2_X1 U12453 ( .A1(n9939), .A2(n9938), .ZN(n9940) );
  AND2_X1 U12454 ( .A1(n9941), .A2(n9940), .ZN(n13091) );
  NAND2_X1 U12455 ( .A1(n13090), .A2(n9941), .ZN(n9943) );
  INV_X1 U12456 ( .A(n10160), .ZN(n9942) );
  AOI21_X1 U12457 ( .B1(n9944), .B2(n9943), .A(n9942), .ZN(n9953) );
  NAND2_X1 U12458 ( .A1(n9946), .A2(n9945), .ZN(n9947) );
  NAND2_X1 U12459 ( .A1(n13575), .A2(n13701), .ZN(n9949) );
  NAND2_X1 U12460 ( .A1(n13573), .A2(n13555), .ZN(n9948) );
  AOI22_X1 U12461 ( .A1(n15125), .A2(n6813), .B1(P2_REG3_REG_4__SCAN_IN), .B2(
        P2_U3088), .ZN(n9950) );
  AOI21_X1 U12462 ( .B1(n10703), .B2(n13556), .A(n9951), .ZN(n9952) );
  OAI21_X1 U12463 ( .B1(n9953), .B2(n13561), .A(n9952), .ZN(P2_U3202) );
  INV_X1 U12464 ( .A(n15576), .ZN(n15573) );
  NAND2_X1 U12465 ( .A1(n9954), .A2(n15576), .ZN(n9955) );
  OAI21_X1 U12466 ( .B1(n15158), .B2(n9410), .A(n9955), .ZN(P2_U3501) );
  INV_X1 U12467 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n9970) );
  INV_X1 U12468 ( .A(n9956), .ZN(n9957) );
  NAND2_X1 U12469 ( .A1(n9958), .A2(n9957), .ZN(n9960) );
  NAND2_X1 U12470 ( .A1(n9961), .A2(n13094), .ZN(n9959) );
  NAND2_X1 U12471 ( .A1(n9960), .A2(n9959), .ZN(n10241) );
  XNOR2_X1 U12472 ( .A(n10241), .B(n10239), .ZN(n10711) );
  NAND2_X1 U12473 ( .A1(n9961), .A2(n10556), .ZN(n9962) );
  OAI21_X1 U12474 ( .B1(n9964), .B2(n10239), .A(n10238), .ZN(n10709) );
  AOI21_X1 U12475 ( .B1(n9965), .B2(n10704), .A(n11865), .ZN(n9966) );
  NAND2_X1 U12476 ( .A1(n9966), .A2(n10248), .ZN(n10706) );
  AOI21_X1 U12477 ( .B1(n10709), .B2(n15527), .A(n9967), .ZN(n9968) );
  OAI21_X1 U12478 ( .B1(n15522), .B2(n10711), .A(n9968), .ZN(n13999) );
  NAND2_X1 U12479 ( .A1(n13999), .A2(n15561), .ZN(n9969) );
  OAI21_X1 U12480 ( .B1(n15561), .B2(n9970), .A(n9969), .ZN(P2_U3442) );
  INV_X1 U12481 ( .A(n11613), .ZN(n10053) );
  OAI222_X1 U12482 ( .A1(n14031), .A2(n10053), .B1(n15478), .B2(P2_U3088), 
        .C1(n9971), .C2(n14038), .ZN(P2_U3312) );
  INV_X1 U12483 ( .A(n9974), .ZN(n9976) );
  XNOR2_X2 U12484 ( .A(n14229), .B(n15319), .ZN(n12150) );
  NAND2_X1 U12485 ( .A1(n14230), .A2(n10203), .ZN(n10198) );
  NAND2_X1 U12486 ( .A1(n12150), .A2(n10198), .ZN(n9979) );
  INV_X1 U12487 ( .A(n14229), .ZN(n10206) );
  NAND2_X1 U12488 ( .A1(n10206), .A2(n15319), .ZN(n9978) );
  NAND2_X1 U12489 ( .A1(n10128), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n9981) );
  NAND2_X1 U12490 ( .A1(n11657), .A2(n14258), .ZN(n9980) );
  XNOR2_X1 U12491 ( .A(n10126), .B(n10132), .ZN(n15327) );
  NAND2_X1 U12492 ( .A1(n14229), .A2(n15319), .ZN(n9983) );
  NAND2_X1 U12493 ( .A1(n11953), .A2(n9983), .ZN(n9985) );
  NAND2_X1 U12494 ( .A1(n10206), .A2(n11960), .ZN(n9984) );
  NAND2_X1 U12495 ( .A1(n9985), .A2(n9984), .ZN(n10133) );
  XNOR2_X1 U12496 ( .A(n10133), .B(n10132), .ZN(n9994) );
  NAND2_X1 U12497 ( .A1(n14229), .A2(n15378), .ZN(n9993) );
  NAND2_X1 U12498 ( .A1(n9986), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n9991) );
  INV_X1 U12499 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n9987) );
  NAND2_X1 U12500 ( .A1(n10117), .A2(n9987), .ZN(n9990) );
  NAND2_X1 U12501 ( .A1(n11088), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n9989) );
  NAND2_X1 U12502 ( .A1(n6658), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n9988) );
  NAND4_X1 U12503 ( .A1(n9991), .A2(n9990), .A3(n9989), .A4(n9988), .ZN(n14227) );
  NAND2_X1 U12504 ( .A1(n14227), .A2(n14966), .ZN(n9992) );
  NAND2_X1 U12505 ( .A1(n9993), .A2(n9992), .ZN(n10013) );
  AOI21_X1 U12506 ( .B1(n9994), .B2(n15375), .A(n10013), .ZN(n15329) );
  INV_X1 U12507 ( .A(n15329), .ZN(n10001) );
  NAND2_X1 U12508 ( .A1(n15319), .A2(n10225), .ZN(n10205) );
  AOI21_X1 U12509 ( .B1(n10205), .B2(n11957), .A(n15320), .ZN(n9995) );
  OR2_X1 U12510 ( .A1(n10205), .A2(n11957), .ZN(n10193) );
  NAND2_X1 U12511 ( .A1(n9995), .A2(n10193), .ZN(n15328) );
  NOR2_X1 U12512 ( .A1(n15328), .A2(n14550), .ZN(n10000) );
  NAND2_X1 U12513 ( .A1(n9996), .A2(n12140), .ZN(n9997) );
  INV_X1 U12514 ( .A(n11957), .ZN(n15330) );
  INV_X1 U12515 ( .A(n14986), .ZN(n15293) );
  AOI22_X1 U12516 ( .A1(n6665), .A2(P1_REG2_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(n15293), .ZN(n9998) );
  OAI21_X1 U12517 ( .B1(n15297), .B2(n15330), .A(n9998), .ZN(n9999) );
  AOI211_X1 U12518 ( .C1(n10001), .C2(n14969), .A(n10000), .B(n9999), .ZN(
        n10002) );
  OAI21_X1 U12519 ( .B1(n14982), .B2(n15327), .A(n10002), .ZN(P1_U3291) );
  NAND2_X1 U12520 ( .A1(n6659), .A2(n6664), .ZN(n10004) );
  NAND2_X1 U12521 ( .A1(n11957), .A2(n11832), .ZN(n10003) );
  NAND2_X1 U12522 ( .A1(n10004), .A2(n10003), .ZN(n10005) );
  XNOR2_X1 U12523 ( .A(n10005), .B(n11830), .ZN(n10674) );
  AND2_X1 U12524 ( .A1(n11957), .A2(n6664), .ZN(n10006) );
  AOI21_X1 U12525 ( .B1(n6659), .B2(n10688), .A(n10006), .ZN(n10675) );
  XNOR2_X1 U12526 ( .A(n10674), .B(n10675), .ZN(n10010) );
  OAI21_X1 U12527 ( .B1(n10010), .B2(n10009), .A(n10678), .ZN(n10011) );
  NAND2_X1 U12528 ( .A1(n10011), .A2(n14195), .ZN(n10015) );
  AOI22_X1 U12529 ( .A1(n10013), .A2(n14115), .B1(P1_REG3_REG_2__SCAN_IN), 
        .B2(n10012), .ZN(n10014) );
  OAI211_X1 U12530 ( .C1(n15330), .C2(n14191), .A(n10015), .B(n10014), .ZN(
        P1_U3237) );
  MUX2_X1 U12531 ( .A(P3_REG2_REG_2__SCAN_IN), .B(P3_REG1_REG_2__SCAN_IN), .S(
        n12694), .Z(n10105) );
  XNOR2_X1 U12532 ( .A(n10105), .B(n10107), .ZN(n10108) );
  MUX2_X1 U12533 ( .A(P3_REG2_REG_1__SCAN_IN), .B(P3_REG1_REG_1__SCAN_IN), .S(
        n12694), .Z(n10017) );
  XOR2_X1 U12534 ( .A(n10365), .B(n10017), .Z(n10361) );
  OAI21_X1 U12535 ( .B1(n10017), .B2(n10365), .A(n10360), .ZN(n10109) );
  XOR2_X1 U12536 ( .A(n10108), .B(n10109), .Z(n10045) );
  INV_X1 U12537 ( .A(n12610), .ZN(n10018) );
  OR2_X1 U12538 ( .A1(n10019), .A2(P3_U3151), .ZN(n12615) );
  NAND2_X1 U12539 ( .A1(n10018), .A2(n12615), .ZN(n10032) );
  NAND2_X1 U12540 ( .A1(n12593), .A2(n10019), .ZN(n10020) );
  AND2_X1 U12541 ( .A1(n10021), .A2(n10020), .ZN(n10031) );
  AND2_X1 U12542 ( .A1(n10032), .A2(n10031), .ZN(n10034) );
  MUX2_X1 U12543 ( .A(n10034), .B(n15577), .S(n10022), .Z(n15604) );
  INV_X1 U12544 ( .A(n10023), .ZN(n10024) );
  INV_X1 U12545 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n13254) );
  NOR3_X1 U12546 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), .A3(
        n13254), .ZN(n10027) );
  NOR2_X1 U12547 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(n13254), .ZN(n10524) );
  INV_X1 U12548 ( .A(n10027), .ZN(n10025) );
  INV_X1 U12549 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n15720) );
  NOR2_X1 U12550 ( .A1(n10355), .A2(n15720), .ZN(n10026) );
  OAI21_X1 U12551 ( .B1(P3_REG2_REG_2__SCAN_IN), .B2(n10092), .A(n10028), .ZN(
        n10029) );
  AOI21_X1 U12552 ( .B1(n10030), .B2(n10029), .A(n10093), .ZN(n10042) );
  INV_X1 U12553 ( .A(n10031), .ZN(n10033) );
  AND2_X1 U12554 ( .A1(n10033), .A2(n10032), .ZN(n15674) );
  AOI22_X1 U12555 ( .A1(n15674), .A2(P3_ADDR_REG_2__SCAN_IN), .B1(
        P3_REG3_REG_2__SCAN_IN), .B2(P3_U3151), .ZN(n10041) );
  NAND2_X1 U12556 ( .A1(n10034), .A2(n12694), .ZN(n12709) );
  INV_X1 U12557 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n15776) );
  AOI22_X1 U12558 ( .A1(n10107), .A2(n15776), .B1(P3_REG1_REG_2__SCAN_IN), 
        .B2(n10092), .ZN(n10038) );
  NAND2_X1 U12559 ( .A1(P3_REG1_REG_0__SCAN_IN), .A2(n10519), .ZN(n10522) );
  INV_X1 U12560 ( .A(n10365), .ZN(n10036) );
  NOR2_X1 U12561 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(n10522), .ZN(n10035) );
  AOI21_X1 U12562 ( .B1(n10036), .B2(n10522), .A(n10035), .ZN(n10353) );
  NAND2_X1 U12563 ( .A1(n10353), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n10352) );
  OAI21_X1 U12564 ( .B1(P3_IR_REG_1__SCAN_IN), .B2(n10522), .A(n10352), .ZN(
        n10037) );
  NAND2_X1 U12565 ( .A1(n10038), .A2(n10037), .ZN(n10084) );
  OAI21_X1 U12566 ( .B1(n10038), .B2(n10037), .A(n10084), .ZN(n10039) );
  NAND2_X1 U12567 ( .A1(n15679), .A2(n10039), .ZN(n10040) );
  OAI211_X1 U12568 ( .C1(n15687), .C2(n10042), .A(n10041), .B(n10040), .ZN(
        n10043) );
  AOI21_X1 U12569 ( .B1(n10107), .B2(n15604), .A(n10043), .ZN(n10044) );
  OAI21_X1 U12570 ( .B1(n10045), .B2(n15661), .A(n10044), .ZN(P3_U3184) );
  INV_X1 U12571 ( .A(P3_DATAO_REG_24__SCAN_IN), .ZN(n13470) );
  NAND2_X1 U12572 ( .A1(n6985), .A2(n15577), .ZN(n10046) );
  OAI21_X1 U12573 ( .B1(n15577), .B2(n13470), .A(n10046), .ZN(P3_U3515) );
  NAND3_X1 U12574 ( .A1(n10049), .A2(n10048), .A3(n10047), .ZN(n10050) );
  OAI21_X1 U12575 ( .B1(n10051), .B2(n10050), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n10052) );
  XNOR2_X1 U12576 ( .A(n10052), .B(P1_IR_REG_15__SCAN_IN), .ZN(n11614) );
  INV_X1 U12577 ( .A(n11614), .ZN(n10963) );
  OAI222_X1 U12578 ( .A1(n14817), .A2(n10054), .B1(n14815), .B2(n10053), .C1(
        n10963), .C2(P1_U3086), .ZN(P1_U3340) );
  INV_X1 U12579 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n10055) );
  AOI22_X1 U12580 ( .A1(P1_REG2_REG_12__SCAN_IN), .A2(n10065), .B1(n11288), 
        .B2(n10055), .ZN(n10059) );
  NAND2_X1 U12581 ( .A1(P1_REG2_REG_11__SCAN_IN), .A2(n11282), .ZN(n10057) );
  NAND2_X1 U12582 ( .A1(n10057), .A2(n10056), .ZN(n10058) );
  NOR2_X1 U12583 ( .A1(n10059), .A2(n10058), .ZN(n10488) );
  AOI21_X1 U12584 ( .B1(n10059), .B2(n10058), .A(n10488), .ZN(n10069) );
  INV_X1 U12585 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n14964) );
  AOI22_X1 U12586 ( .A1(P1_REG1_REG_12__SCAN_IN), .A2(n10065), .B1(n11288), 
        .B2(n14964), .ZN(n10062) );
  AOI21_X1 U12587 ( .B1(n10063), .B2(n10062), .A(n10495), .ZN(n10064) );
  OR2_X1 U12588 ( .A1(n10064), .A2(n15264), .ZN(n10068) );
  AND2_X1 U12589 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n14091) );
  NOR2_X1 U12590 ( .A1(n15267), .A2(n10065), .ZN(n10066) );
  AOI211_X1 U12591 ( .C1(n14360), .C2(P1_ADDR_REG_12__SCAN_IN), .A(n14091), 
        .B(n10066), .ZN(n10067) );
  OAI211_X1 U12592 ( .C1(n10069), .C2(n15266), .A(n10068), .B(n10067), .ZN(
        P1_U3255) );
  INV_X1 U12593 ( .A(n15490), .ZN(n10070) );
  NAND2_X1 U12594 ( .A1(n10071), .A2(n10070), .ZN(n10072) );
  INV_X4 U12595 ( .A(n13852), .ZN(n15151) );
  AOI21_X1 U12596 ( .B1(n9247), .B2(n13852), .A(n15147), .ZN(n10080) );
  NAND2_X1 U12597 ( .A1(n10295), .A2(n10073), .ZN(n15492) );
  AOI21_X1 U12598 ( .B1(n15522), .B2(n9794), .A(n15494), .ZN(n10075) );
  NOR2_X1 U12599 ( .A1(n10075), .A2(n10074), .ZN(n15493) );
  INV_X1 U12600 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n10076) );
  OAI22_X1 U12601 ( .A1(n15151), .A2(n15493), .B1(n10076), .B2(n13865), .ZN(
        n10078) );
  OR2_X1 U12602 ( .A1(n15151), .A2(n10235), .ZN(n10581) );
  NOR2_X1 U12603 ( .A1(n10581), .A2(n15494), .ZN(n10077) );
  AOI211_X1 U12604 ( .C1(n15151), .C2(P2_REG2_REG_0__SCAN_IN), .A(n10078), .B(
        n10077), .ZN(n10079) );
  OAI21_X1 U12605 ( .B1(n10080), .B2(n15492), .A(n10079), .ZN(P2_U3265) );
  INV_X1 U12606 ( .A(n10081), .ZN(n10083) );
  OAI222_X1 U12607 ( .A1(P3_U3151), .A2(n12666), .B1(n14938), .B2(n10083), 
        .C1(n10082), .C2(n14936), .ZN(P3_U3276) );
  NAND2_X1 U12608 ( .A1(P3_REG1_REG_2__SCAN_IN), .A2(n10092), .ZN(n10085) );
  NAND2_X1 U12609 ( .A1(n10085), .A2(n10084), .ZN(n10086) );
  XNOR2_X1 U12610 ( .A(n10086), .B(n10280), .ZN(n10285) );
  NAND2_X1 U12611 ( .A1(n10285), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n10088) );
  INV_X1 U12612 ( .A(n10280), .ZN(n10110) );
  NAND2_X1 U12613 ( .A1(n10086), .A2(n10110), .ZN(n10087) );
  NAND2_X1 U12614 ( .A1(n10088), .A2(n10087), .ZN(n10090) );
  AOI22_X1 U12615 ( .A1(P3_REG1_REG_4__SCAN_IN), .A2(n10264), .B1(n10258), 
        .B2(n8060), .ZN(n10089) );
  NAND2_X1 U12616 ( .A1(n10089), .A2(n10090), .ZN(n10265) );
  OAI21_X1 U12617 ( .B1(n10090), .B2(n10089), .A(n10265), .ZN(n10091) );
  INV_X1 U12618 ( .A(n10091), .ZN(n10104) );
  AND2_X1 U12619 ( .A1(P3_U3151), .A2(P3_REG3_REG_4__SCAN_IN), .ZN(n10780) );
  AOI21_X1 U12620 ( .B1(n15674), .B2(P3_ADDR_REG_4__SCAN_IN), .A(n10780), .ZN(
        n10103) );
  OAI21_X1 U12621 ( .B1(n10094), .B2(n10110), .A(n10095), .ZN(n10281) );
  NOR2_X1 U12622 ( .A1(n10281), .A2(n8047), .ZN(n10283) );
  INV_X1 U12623 ( .A(n10095), .ZN(n10096) );
  NOR2_X1 U12624 ( .A1(n10283), .A2(n10096), .ZN(n10099) );
  NAND2_X1 U12625 ( .A1(P3_REG2_REG_4__SCAN_IN), .A2(n10264), .ZN(n10097) );
  OAI21_X1 U12626 ( .B1(P3_REG2_REG_4__SCAN_IN), .B2(n10264), .A(n10097), .ZN(
        n10098) );
  AOI21_X1 U12627 ( .B1(n10099), .B2(n10098), .A(n10261), .ZN(n10100) );
  INV_X1 U12628 ( .A(n10100), .ZN(n10101) );
  NAND2_X1 U12629 ( .A1(n15082), .A2(n10101), .ZN(n10102) );
  OAI211_X1 U12630 ( .C1(n10104), .C2(n12709), .A(n10103), .B(n10102), .ZN(
        n10114) );
  MUX2_X1 U12631 ( .A(P3_REG2_REG_4__SCAN_IN), .B(P3_REG1_REG_4__SCAN_IN), .S(
        n12694), .Z(n10256) );
  XNOR2_X1 U12632 ( .A(n10256), .B(n10258), .ZN(n10259) );
  INV_X1 U12633 ( .A(n10105), .ZN(n10106) );
  AOI22_X1 U12634 ( .A1(n10109), .A2(n10108), .B1(n10107), .B2(n10106), .ZN(
        n10279) );
  MUX2_X1 U12635 ( .A(P3_REG2_REG_3__SCAN_IN), .B(P3_REG1_REG_3__SCAN_IN), .S(
        n12696), .Z(n10111) );
  XOR2_X1 U12636 ( .A(n10280), .B(n10111), .Z(n10278) );
  OAI22_X1 U12637 ( .A1(n10279), .A2(n10278), .B1(n10111), .B2(n10110), .ZN(
        n10260) );
  XOR2_X1 U12638 ( .A(n10259), .B(n10260), .Z(n10112) );
  NOR2_X1 U12639 ( .A1(n10112), .A2(n15661), .ZN(n10113) );
  AOI211_X1 U12640 ( .C1(n15604), .C2(n10258), .A(n10114), .B(n10113), .ZN(
        n10115) );
  INV_X1 U12641 ( .A(n10115), .ZN(P3_U3186) );
  NAND2_X1 U12642 ( .A1(n11837), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n10122) );
  INV_X1 U12643 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n10118) );
  XNOR2_X1 U12644 ( .A(n10118), .B(P1_REG3_REG_3__SCAN_IN), .ZN(n10148) );
  NAND2_X1 U12645 ( .A1(n11839), .A2(n10148), .ZN(n10121) );
  NAND2_X1 U12646 ( .A1(n11808), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n10120) );
  NAND2_X1 U12647 ( .A1(n11088), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n10119) );
  NAND4_X1 U12648 ( .A1(n10122), .A2(n10121), .A3(n10120), .A4(n10119), .ZN(
        n14226) );
  NAND2_X1 U12649 ( .A1(n12110), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n10124) );
  NAND2_X1 U12650 ( .A1(n11657), .A2(n14284), .ZN(n10123) );
  OAI211_X1 U12651 ( .C1(n12109), .C2(n10125), .A(n10124), .B(n10123), .ZN(
        n11982) );
  NOR2_X1 U12652 ( .A1(n14226), .A2(n11982), .ZN(n10422) );
  NOR2_X1 U12653 ( .A1(n10422), .A2(n6709), .ZN(n12149) );
  NAND2_X1 U12654 ( .A1(n10201), .A2(n15330), .ZN(n10127) );
  NAND2_X1 U12655 ( .A1(n10128), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n10129) );
  INV_X1 U12656 ( .A(n14064), .ZN(n10194) );
  INV_X1 U12657 ( .A(n14227), .ZN(n10136) );
  NAND2_X1 U12658 ( .A1(n10136), .A2(n10194), .ZN(n10131) );
  XOR2_X1 U12659 ( .A(n12149), .B(n10423), .Z(n10386) );
  NAND2_X1 U12660 ( .A1(n10133), .A2(n10132), .ZN(n10135) );
  NAND2_X1 U12661 ( .A1(n10201), .A2(n11957), .ZN(n10134) );
  NAND2_X1 U12662 ( .A1(n10135), .A2(n10134), .ZN(n10186) );
  NAND2_X1 U12663 ( .A1(n14227), .A2(n10194), .ZN(n11972) );
  NAND2_X1 U12664 ( .A1(n10186), .A2(n11972), .ZN(n10137) );
  NAND2_X1 U12665 ( .A1(n10136), .A2(n14064), .ZN(n11970) );
  XOR2_X1 U12666 ( .A(n10453), .B(n12149), .Z(n10138) );
  NAND2_X1 U12667 ( .A1(n10138), .A2(n15375), .ZN(n10384) );
  INV_X1 U12668 ( .A(n10384), .ZN(n10146) );
  NAND2_X1 U12669 ( .A1(n14227), .A2(n15378), .ZN(n10145) );
  NAND2_X1 U12670 ( .A1(n12112), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n10143) );
  AOI21_X1 U12671 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(P1_REG3_REG_5__SCAN_IN), .ZN(n10139) );
  AND3_X1 U12672 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n10429) );
  NOR2_X1 U12673 ( .A1(n10139), .A2(n10429), .ZN(n15294) );
  NAND2_X1 U12674 ( .A1(n10117), .A2(n15294), .ZN(n10142) );
  NAND2_X1 U12675 ( .A1(n11808), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n10141) );
  NAND2_X1 U12676 ( .A1(n11088), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n10140) );
  NAND4_X1 U12677 ( .A1(n10143), .A2(n10142), .A3(n10141), .A4(n10140), .ZN(
        n14225) );
  NAND2_X1 U12678 ( .A1(n14225), .A2(n14966), .ZN(n10144) );
  NAND2_X1 U12679 ( .A1(n10145), .A2(n10144), .ZN(n10696) );
  OAI21_X1 U12680 ( .B1(n10146), .B2(n10696), .A(n14969), .ZN(n10152) );
  INV_X1 U12681 ( .A(n11982), .ZN(n10451) );
  OR2_X1 U12682 ( .A1(n10192), .A2(n10451), .ZN(n10147) );
  AND3_X1 U12683 ( .A1(n10592), .A2(n15288), .A3(n10147), .ZN(n10383) );
  NOR2_X1 U12684 ( .A1(n15297), .A2(n10451), .ZN(n10150) );
  INV_X1 U12685 ( .A(n10148), .ZN(n10699) );
  OAI22_X1 U12686 ( .A1(n14969), .A2(n9734), .B1(n10699), .B2(n14986), .ZN(
        n10149) );
  AOI211_X1 U12687 ( .C1(n10383), .C2(n15299), .A(n10150), .B(n10149), .ZN(
        n10151) );
  OAI211_X1 U12688 ( .C1(n10386), .C2(n14982), .A(n10152), .B(n10151), .ZN(
        P1_U3289) );
  INV_X1 U12689 ( .A(n11620), .ZN(n10233) );
  INV_X1 U12690 ( .A(n10870), .ZN(n11106) );
  OAI222_X1 U12691 ( .A1(n14031), .A2(n10233), .B1(n11106), .B2(P2_U3088), 
        .C1(n10153), .C2(n14038), .ZN(P2_U3311) );
  INV_X1 U12692 ( .A(n10154), .ZN(n10251) );
  XNOR2_X1 U12693 ( .A(n10543), .B(n13107), .ZN(n10366) );
  NAND2_X1 U12694 ( .A1(n13573), .A2(n11865), .ZN(n10367) );
  XNOR2_X1 U12695 ( .A(n10366), .B(n10367), .ZN(n10162) );
  INV_X1 U12696 ( .A(n10155), .ZN(n10158) );
  INV_X1 U12697 ( .A(n10156), .ZN(n10157) );
  NAND2_X1 U12698 ( .A1(n10158), .A2(n10157), .ZN(n10159) );
  OAI21_X1 U12699 ( .B1(n10162), .B2(n10161), .A(n10376), .ZN(n10163) );
  NAND2_X1 U12700 ( .A1(n10163), .A2(n15123), .ZN(n10169) );
  NAND2_X1 U12701 ( .A1(n13574), .A2(n13701), .ZN(n10165) );
  NAND2_X1 U12702 ( .A1(n13572), .A2(n13555), .ZN(n10164) );
  AND2_X1 U12703 ( .A1(n10165), .A2(n10164), .ZN(n10245) );
  OAI21_X1 U12704 ( .B1(n13558), .B2(n10245), .A(n10166), .ZN(n10167) );
  AOI21_X1 U12705 ( .B1(n10543), .B2(n15128), .A(n10167), .ZN(n10168) );
  OAI211_X1 U12706 ( .C1(n15131), .C2(n10251), .A(n10169), .B(n10168), .ZN(
        P2_U3199) );
  NAND2_X1 U12707 ( .A1(n15454), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n10176) );
  AOI21_X1 U12708 ( .B1(n10172), .B2(n10171), .A(n10170), .ZN(n15457) );
  INV_X1 U12709 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n10175) );
  INV_X1 U12710 ( .A(n10176), .ZN(n10173) );
  AOI21_X1 U12711 ( .B1(n10175), .B2(n10174), .A(n10173), .ZN(n15456) );
  NAND2_X1 U12712 ( .A1(n15457), .A2(n15456), .ZN(n15455) );
  NAND2_X1 U12713 ( .A1(n10176), .A2(n15455), .ZN(n10864) );
  XNOR2_X1 U12714 ( .A(n10864), .B(n10865), .ZN(n10866) );
  XOR2_X1 U12715 ( .A(P2_REG2_REG_14__SCAN_IN), .B(n10866), .Z(n10183) );
  AOI22_X1 U12716 ( .A1(n15453), .A2(n10865), .B1(n15472), .B2(
        P2_ADDR_REG_14__SCAN_IN), .ZN(n10182) );
  NAND2_X1 U12717 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3088), .ZN(n15129)
         );
  XNOR2_X1 U12718 ( .A(n10865), .B(P2_REG1_REG_14__SCAN_IN), .ZN(n10877) );
  OAI21_X1 U12719 ( .B1(n10178), .B2(P2_REG1_REG_12__SCAN_IN), .A(n10177), 
        .ZN(n15460) );
  INV_X1 U12720 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n11435) );
  MUX2_X1 U12721 ( .A(n11435), .B(P2_REG1_REG_13__SCAN_IN), .S(n15454), .Z(
        n15461) );
  NOR2_X1 U12722 ( .A1(n15460), .A2(n15461), .ZN(n15458) );
  AOI21_X1 U12723 ( .B1(n15454), .B2(P2_REG1_REG_13__SCAN_IN), .A(n15458), 
        .ZN(n10878) );
  XOR2_X1 U12724 ( .A(n10877), .B(n10878), .Z(n10179) );
  NAND2_X1 U12725 ( .A1(n10179), .A2(n15467), .ZN(n10180) );
  AND2_X1 U12726 ( .A1(n15129), .A2(n10180), .ZN(n10181) );
  OAI211_X1 U12727 ( .C1(n10183), .C2(n15442), .A(n10182), .B(n10181), .ZN(
        P2_U3228) );
  XNOR2_X1 U12728 ( .A(n10184), .B(n11976), .ZN(n10190) );
  INV_X1 U12729 ( .A(n10190), .ZN(n10217) );
  NAND2_X1 U12730 ( .A1(n10185), .A2(n14612), .ZN(n12132) );
  OR2_X1 U12731 ( .A1(n6665), .A2(n12132), .ZN(n15284) );
  INV_X1 U12732 ( .A(n15318), .ZN(n15345) );
  XNOR2_X1 U12733 ( .A(n11976), .B(n10186), .ZN(n10188) );
  AOI22_X1 U12734 ( .A1(n15378), .A2(n6659), .B1(n14226), .B2(n14966), .ZN(
        n10187) );
  OAI21_X1 U12735 ( .B1(n10188), .B2(n15351), .A(n10187), .ZN(n10189) );
  AOI21_X1 U12736 ( .B1(n15345), .B2(n10190), .A(n10189), .ZN(n10216) );
  MUX2_X1 U12737 ( .A(n10191), .B(n10216), .S(n14969), .Z(n10197) );
  AOI21_X1 U12738 ( .B1(n14064), .B2(n10193), .A(n10192), .ZN(n10214) );
  NAND2_X1 U12739 ( .A1(n15299), .A2(n15288), .ZN(n14675) );
  INV_X1 U12740 ( .A(n14675), .ZN(n14628) );
  OAI22_X1 U12741 ( .A1(n15297), .A2(n10194), .B1(P1_REG3_REG_3__SCAN_IN), 
        .B2(n14986), .ZN(n10195) );
  AOI21_X1 U12742 ( .B1(n10214), .B2(n14628), .A(n10195), .ZN(n10196) );
  OAI211_X1 U12743 ( .C1(n10217), .C2(n15284), .A(n10197), .B(n10196), .ZN(
        P1_U3290) );
  INV_X1 U12744 ( .A(n10198), .ZN(n10199) );
  XNOR2_X1 U12745 ( .A(n12150), .B(n10199), .ZN(n15317) );
  INV_X1 U12746 ( .A(n14230), .ZN(n10202) );
  OAI21_X1 U12747 ( .B1(n12150), .B2(n10202), .A(n15375), .ZN(n10200) );
  AND2_X1 U12748 ( .A1(n10200), .A2(n15212), .ZN(n15316) );
  OAI22_X1 U12749 ( .A1(n15316), .A2(n10202), .B1(n10201), .B2(n14607), .ZN(
        n15324) );
  NAND2_X1 U12750 ( .A1(n15324), .A2(n14969), .ZN(n10213) );
  INV_X1 U12751 ( .A(n15316), .ZN(n10211) );
  NAND2_X1 U12752 ( .A1(n10203), .A2(n11960), .ZN(n10204) );
  NAND2_X1 U12753 ( .A1(n10205), .A2(n10204), .ZN(n15321) );
  XNOR2_X1 U12754 ( .A(n10206), .B(n15321), .ZN(n15315) );
  NOR2_X1 U12755 ( .A1(n15315), .A2(n14599), .ZN(n10210) );
  NAND2_X1 U12756 ( .A1(n15282), .A2(n11960), .ZN(n10208) );
  AOI22_X1 U12757 ( .A1(n6665), .A2(P1_REG2_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(n15293), .ZN(n10207) );
  OAI211_X1 U12758 ( .C1(n15321), .C2(n14675), .A(n10208), .B(n10207), .ZN(
        n10209) );
  AOI21_X1 U12759 ( .B1(n10211), .B2(n10210), .A(n10209), .ZN(n10212) );
  OAI211_X1 U12760 ( .C1(n14982), .C2(n15317), .A(n10213), .B(n10212), .ZN(
        P1_U3292) );
  INV_X1 U12761 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n10219) );
  AOI22_X1 U12762 ( .A1(n10214), .A2(n15288), .B1(n15379), .B2(n14064), .ZN(
        n10215) );
  OAI211_X1 U12763 ( .C1(n15341), .C2(n10217), .A(n10216), .B(n10215), .ZN(
        n10220) );
  NAND2_X1 U12764 ( .A1(n10220), .A2(n15389), .ZN(n10218) );
  OAI21_X1 U12765 ( .B1(n15389), .B2(n10219), .A(n10218), .ZN(P1_U3468) );
  NAND2_X1 U12766 ( .A1(n10220), .A2(n15403), .ZN(n10221) );
  OAI21_X1 U12767 ( .B1(n15403), .B2(n10222), .A(n10221), .ZN(P1_U3531) );
  OAI22_X1 U12768 ( .A1(n6665), .A2(n10224), .B1(n10223), .B2(n14986), .ZN(
        n10227) );
  AOI21_X1 U12769 ( .B1(n14675), .B2(n15297), .A(n10225), .ZN(n10226) );
  AOI211_X1 U12770 ( .C1(n6665), .C2(P1_REG2_REG_0__SCAN_IN), .A(n10227), .B(
        n10226), .ZN(n10229) );
  INV_X1 U12771 ( .A(n14599), .ZN(n14654) );
  OAI21_X1 U12772 ( .B1(n15191), .B2(n14654), .A(n12148), .ZN(n10228) );
  NAND2_X1 U12773 ( .A1(n10229), .A2(n10228), .ZN(P1_U3293) );
  NAND2_X1 U12774 ( .A1(n10231), .A2(n10230), .ZN(n10410) );
  NAND2_X1 U12775 ( .A1(n10410), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10232) );
  XNOR2_X1 U12776 ( .A(n10232), .B(P1_IR_REG_16__SCAN_IN), .ZN(n11621) );
  INV_X1 U12777 ( .A(n11621), .ZN(n14353) );
  OAI222_X1 U12778 ( .A1(n14817), .A2(n10234), .B1(n14815), .B2(n10233), .C1(
        n14353), .C2(P1_U3086), .ZN(P1_U3339) );
  AND2_X1 U12779 ( .A1(n9794), .A2(n10235), .ZN(n10236) );
  INV_X1 U12780 ( .A(n13574), .ZN(n10242) );
  XNOR2_X1 U12781 ( .A(n10545), .B(n10244), .ZN(n15505) );
  INV_X1 U12782 ( .A(n10239), .ZN(n10240) );
  NAND2_X1 U12783 ( .A1(n10242), .A2(n10704), .ZN(n10243) );
  XOR2_X1 U12784 ( .A(n10533), .B(n10244), .Z(n10246) );
  OAI21_X1 U12785 ( .B1(n10246), .B2(n15522), .A(n10245), .ZN(n15509) );
  INV_X1 U12786 ( .A(n15509), .ZN(n10247) );
  MUX2_X1 U12787 ( .A(n6846), .B(n10247), .S(n13852), .Z(n10255) );
  INV_X1 U12788 ( .A(n10248), .ZN(n10249) );
  INV_X1 U12789 ( .A(n10543), .ZN(n15507) );
  OAI211_X1 U12790 ( .C1(n10249), .C2(n15507), .A(n15144), .B(n10575), .ZN(
        n15506) );
  INV_X1 U12791 ( .A(n15506), .ZN(n10253) );
  OAI22_X1 U12792 ( .A1(n13890), .A2(n15507), .B1(n13865), .B2(n10251), .ZN(
        n10252) );
  AOI21_X1 U12793 ( .B1(n15147), .B2(n10253), .A(n10252), .ZN(n10254) );
  OAI211_X1 U12794 ( .C1(n13874), .C2(n15505), .A(n10255), .B(n10254), .ZN(
        P2_U3260) );
  INV_X1 U12795 ( .A(n10256), .ZN(n10257) );
  AOI22_X1 U12796 ( .A1(n10260), .A2(n10259), .B1(n10258), .B2(n10257), .ZN(
        n10331) );
  MUX2_X1 U12797 ( .A(P3_REG2_REG_5__SCAN_IN), .B(P3_REG1_REG_5__SCAN_IN), .S(
        n12696), .Z(n10329) );
  XNOR2_X1 U12798 ( .A(n10329), .B(n10337), .ZN(n10330) );
  XNOR2_X1 U12799 ( .A(n10331), .B(n10330), .ZN(n10276) );
  XNOR2_X1 U12800 ( .A(n10332), .B(n10333), .ZN(n10263) );
  INV_X1 U12801 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n10262) );
  AOI21_X1 U12802 ( .B1(n10263), .B2(n10262), .A(n10334), .ZN(n10274) );
  NAND2_X1 U12803 ( .A1(P3_REG1_REG_4__SCAN_IN), .A2(n10264), .ZN(n10266) );
  NAND2_X1 U12804 ( .A1(P3_REG1_REG_5__SCAN_IN), .A2(n10267), .ZN(n10338) );
  OAI21_X1 U12805 ( .B1(P3_REG1_REG_5__SCAN_IN), .B2(n10267), .A(n10338), .ZN(
        n10268) );
  INV_X1 U12806 ( .A(n10268), .ZN(n10270) );
  NAND2_X1 U12807 ( .A1(P3_U3151), .A2(P3_REG3_REG_5__SCAN_IN), .ZN(n10976) );
  NAND2_X1 U12808 ( .A1(n15674), .A2(P3_ADDR_REG_5__SCAN_IN), .ZN(n10269) );
  OAI211_X1 U12809 ( .C1(n12709), .C2(n10270), .A(n10976), .B(n10269), .ZN(
        n10271) );
  INV_X1 U12810 ( .A(n10271), .ZN(n10273) );
  NAND2_X1 U12811 ( .A1(n15604), .A2(n10333), .ZN(n10272) );
  OAI211_X1 U12812 ( .C1(n15687), .C2(n10274), .A(n10273), .B(n10272), .ZN(
        n10275) );
  AOI21_X1 U12813 ( .B1(n10276), .B2(n15681), .A(n10275), .ZN(n10277) );
  INV_X1 U12814 ( .A(n10277), .ZN(P3_U3187) );
  XNOR2_X1 U12815 ( .A(n10279), .B(n10278), .ZN(n10292) );
  NAND2_X1 U12816 ( .A1(n15604), .A2(n10280), .ZN(n10290) );
  AOI22_X1 U12817 ( .A1(n15674), .A2(P3_ADDR_REG_3__SCAN_IN), .B1(
        P3_REG3_REG_3__SCAN_IN), .B2(P3_U3151), .ZN(n10289) );
  AND2_X1 U12818 ( .A1(n10281), .A2(n8047), .ZN(n10282) );
  OAI21_X1 U12819 ( .B1(n10283), .B2(n10282), .A(n15082), .ZN(n10288) );
  INV_X1 U12820 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n10284) );
  XNOR2_X1 U12821 ( .A(n10285), .B(n10284), .ZN(n10286) );
  OR2_X1 U12822 ( .A1(n12709), .A2(n10286), .ZN(n10287) );
  NAND4_X1 U12823 ( .A1(n10290), .A2(n10289), .A3(n10288), .A4(n10287), .ZN(
        n10291) );
  AOI21_X1 U12824 ( .B1(n10292), .B2(n15681), .A(n10291), .ZN(n10293) );
  INV_X1 U12825 ( .A(n10293), .ZN(P3_U3185) );
  XNOR2_X1 U12826 ( .A(n10299), .B(n10294), .ZN(n15501) );
  AOI21_X1 U12827 ( .B1(n10295), .B2(n6672), .A(n11865), .ZN(n10297) );
  AND2_X1 U12828 ( .A1(n10297), .A2(n10296), .ZN(n15497) );
  OAI21_X1 U12829 ( .B1(n10300), .B2(n10299), .A(n10298), .ZN(n10302) );
  AOI21_X1 U12830 ( .B1(n10302), .B2(n15551), .A(n10301), .ZN(n15500) );
  NOR2_X1 U12831 ( .A1(n15151), .A2(n15500), .ZN(n10305) );
  INV_X1 U12832 ( .A(n13865), .ZN(n15137) );
  AOI22_X1 U12833 ( .A1(n15151), .A2(P2_REG2_REG_1__SCAN_IN), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(n15137), .ZN(n10303) );
  OAI21_X1 U12834 ( .B1(n13890), .B2(n7362), .A(n10303), .ZN(n10304) );
  AOI211_X1 U12835 ( .C1(n15497), .C2(n15147), .A(n10305), .B(n10304), .ZN(
        n10306) );
  OAI21_X1 U12836 ( .B1(n13874), .B2(n15501), .A(n10306), .ZN(P2_U3264) );
  NAND3_X1 U12837 ( .A1(n12416), .A2(n15744), .A3(n10307), .ZN(n10308) );
  OAI21_X1 U12838 ( .B1(n7130), .B2(n15017), .A(n10308), .ZN(n10715) );
  INV_X1 U12839 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n10309) );
  OAI22_X1 U12840 ( .A1(n13049), .A2(n9876), .B1(n15773), .B2(n10309), .ZN(
        n10310) );
  AOI21_X1 U12841 ( .B1(n10715), .B2(n15773), .A(n10310), .ZN(n10311) );
  INV_X1 U12842 ( .A(n10311), .ZN(P3_U3390) );
  INV_X1 U12843 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n15710) );
  INV_X1 U12844 ( .A(n10312), .ZN(n10315) );
  INV_X1 U12845 ( .A(n12442), .ZN(n10314) );
  NOR2_X1 U12846 ( .A1(n10316), .A2(n12270), .ZN(n10317) );
  AND2_X1 U12847 ( .A1(n10318), .A2(n10317), .ZN(n10319) );
  NAND2_X1 U12848 ( .A1(n15706), .A2(n12234), .ZN(n10320) );
  NAND2_X1 U12849 ( .A1(n10321), .A2(n10320), .ZN(n10322) );
  NAND2_X1 U12850 ( .A1(n10324), .A2(n10322), .ZN(n10467) );
  NAND3_X1 U12851 ( .A1(n15705), .A2(n12441), .A3(n12270), .ZN(n10323) );
  OAI211_X1 U12852 ( .C1(n10324), .C2(n15706), .A(n10467), .B(n10323), .ZN(
        n10325) );
  NAND2_X1 U12853 ( .A1(n10325), .A2(n15021), .ZN(n10328) );
  INV_X1 U12854 ( .A(n12638), .ZN(n10326) );
  INV_X1 U12855 ( .A(n12867), .ZN(n15019) );
  INV_X1 U12856 ( .A(n12637), .ZN(n10473) );
  OAI22_X1 U12857 ( .A1(n10326), .A2(n15019), .B1(n10473), .B2(n15017), .ZN(
        n15721) );
  INV_X1 U12858 ( .A(n15009), .ZN(n15591) );
  INV_X1 U12859 ( .A(n15581), .ZN(n15012) );
  AOI22_X1 U12860 ( .A1(n15721), .A2(n15591), .B1(n7129), .B2(n15012), .ZN(
        n10327) );
  OAI211_X1 U12861 ( .C1(n10487), .C2(n15710), .A(n10328), .B(n10327), .ZN(
        P3_U3162) );
  MUX2_X1 U12862 ( .A(P3_REG2_REG_6__SCAN_IN), .B(P3_REG1_REG_6__SCAN_IN), .S(
        n12694), .Z(n10391) );
  XNOR2_X1 U12863 ( .A(n10391), .B(n10393), .ZN(n10394) );
  OAI22_X1 U12864 ( .A1(n10331), .A2(n10330), .B1(n10329), .B2(n10337), .ZN(
        n10395) );
  XOR2_X1 U12865 ( .A(n10394), .B(n10395), .Z(n10351) );
  NAND2_X1 U12866 ( .A1(P3_REG2_REG_6__SCAN_IN), .A2(n10401), .ZN(n10335) );
  OAI21_X1 U12867 ( .B1(P3_REG2_REG_6__SCAN_IN), .B2(n10401), .A(n10335), .ZN(
        n10400) );
  XNOR2_X1 U12868 ( .A(n6818), .B(n10400), .ZN(n10349) );
  INV_X1 U12869 ( .A(P3_ADDR_REG_6__SCAN_IN), .ZN(n10346) );
  INV_X1 U12870 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n15782) );
  AOI22_X1 U12871 ( .A1(n10393), .A2(n15782), .B1(P3_REG1_REG_6__SCAN_IN), 
        .B2(n10401), .ZN(n10341) );
  NAND2_X1 U12872 ( .A1(n10337), .A2(n10336), .ZN(n10339) );
  NAND2_X1 U12873 ( .A1(n10339), .A2(n10338), .ZN(n10340) );
  NAND2_X1 U12874 ( .A1(n10341), .A2(n10340), .ZN(n10396) );
  OAI21_X1 U12875 ( .B1(n10341), .B2(n10340), .A(n10396), .ZN(n10342) );
  NAND2_X1 U12876 ( .A1(n15679), .A2(n10342), .ZN(n10345) );
  INV_X1 U12877 ( .A(P3_REG3_REG_6__SCAN_IN), .ZN(n10343) );
  NOR2_X1 U12878 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10343), .ZN(n11045) );
  INV_X1 U12879 ( .A(n11045), .ZN(n10344) );
  OAI211_X1 U12880 ( .C1(n15613), .C2(n10346), .A(n10345), .B(n10344), .ZN(
        n10348) );
  INV_X1 U12881 ( .A(n15604), .ZN(n15677) );
  NOR2_X1 U12882 ( .A1(n15677), .A2(n10401), .ZN(n10347) );
  AOI211_X1 U12883 ( .C1(n15082), .C2(n10349), .A(n10348), .B(n10347), .ZN(
        n10350) );
  OAI21_X1 U12884 ( .B1(n10351), .B2(n15661), .A(n10350), .ZN(P3_U3188) );
  OAI21_X1 U12885 ( .B1(P3_REG1_REG_1__SCAN_IN), .B2(n10353), .A(n10352), .ZN(
        n10359) );
  INV_X1 U12886 ( .A(P3_ADDR_REG_1__SCAN_IN), .ZN(n10354) );
  OAI22_X1 U12887 ( .A1(n15613), .A2(n10354), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n15710), .ZN(n10358) );
  XOR2_X1 U12888 ( .A(n15720), .B(n10355), .Z(n10356) );
  NOR2_X1 U12889 ( .A1(n15687), .A2(n10356), .ZN(n10357) );
  AOI211_X1 U12890 ( .C1(n15679), .C2(n10359), .A(n10358), .B(n10357), .ZN(
        n10364) );
  OAI21_X1 U12891 ( .B1(n10361), .B2(n10521), .A(n10360), .ZN(n10362) );
  NAND2_X1 U12892 ( .A1(n10362), .A2(n15681), .ZN(n10363) );
  OAI211_X1 U12893 ( .C1(n15677), .C2(n10365), .A(n10364), .B(n10363), .ZN(
        P3_U3183) );
  INV_X1 U12894 ( .A(n10366), .ZN(n10368) );
  NAND2_X1 U12895 ( .A1(n10368), .A2(n10367), .ZN(n10374) );
  AND2_X1 U12896 ( .A1(n10376), .A2(n10374), .ZN(n10378) );
  XNOR2_X1 U12897 ( .A(n15513), .B(n13107), .ZN(n10369) );
  AND2_X1 U12898 ( .A1(n13572), .A2(n11865), .ZN(n10370) );
  NAND2_X1 U12899 ( .A1(n10369), .A2(n10370), .ZN(n10415) );
  INV_X1 U12900 ( .A(n10369), .ZN(n10372) );
  INV_X1 U12901 ( .A(n10370), .ZN(n10371) );
  NAND2_X1 U12902 ( .A1(n10372), .A2(n10371), .ZN(n10373) );
  AND2_X1 U12903 ( .A1(n10415), .A2(n10373), .ZN(n10377) );
  AND2_X1 U12904 ( .A1(n10377), .A2(n10374), .ZN(n10375) );
  NAND2_X1 U12905 ( .A1(n10376), .A2(n10375), .ZN(n10416) );
  OAI211_X1 U12906 ( .C1(n10378), .C2(n10377), .A(n10416), .B(n15123), .ZN(
        n10382) );
  INV_X1 U12907 ( .A(n13573), .ZN(n10546) );
  OAI22_X1 U12908 ( .A1(n10793), .A2(n13630), .B1(n10546), .B2(n13496), .ZN(
        n10572) );
  INV_X1 U12909 ( .A(n10572), .ZN(n10379) );
  NAND2_X1 U12910 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3088), .ZN(n15437) );
  OAI21_X1 U12911 ( .B1(n13558), .B2(n10379), .A(n15437), .ZN(n10380) );
  AOI21_X1 U12912 ( .B1(n10576), .B2(n13556), .A(n10380), .ZN(n10381) );
  OAI211_X1 U12913 ( .C1(n7435), .C2(n13542), .A(n10382), .B(n10381), .ZN(
        P2_U3211) );
  AOI211_X1 U12914 ( .C1(n15379), .C2(n11982), .A(n10696), .B(n10383), .ZN(
        n10385) );
  OAI211_X1 U12915 ( .C1(n10386), .C2(n15219), .A(n10385), .B(n10384), .ZN(
        n10388) );
  NAND2_X1 U12916 ( .A1(n10388), .A2(n15403), .ZN(n10387) );
  OAI21_X1 U12917 ( .B1(n15403), .B2(n9711), .A(n10387), .ZN(P1_U3532) );
  INV_X1 U12918 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n10390) );
  NAND2_X1 U12919 ( .A1(n10388), .A2(n15389), .ZN(n10389) );
  OAI21_X1 U12920 ( .B1(n15389), .B2(n10390), .A(n10389), .ZN(P1_U3471) );
  INV_X1 U12921 ( .A(n11637), .ZN(n10413) );
  INV_X1 U12922 ( .A(n11111), .ZN(n11200) );
  OAI222_X1 U12923 ( .A1(n14031), .A2(n10413), .B1(n11200), .B2(P2_U3088), 
        .C1(n7532), .C2(n14038), .ZN(P2_U3310) );
  MUX2_X1 U12924 ( .A(P3_REG2_REG_7__SCAN_IN), .B(P3_REG1_REG_7__SCAN_IN), .S(
        n12694), .Z(n10605) );
  XNOR2_X1 U12925 ( .A(n10605), .B(n10613), .ZN(n10606) );
  INV_X1 U12926 ( .A(n10391), .ZN(n10392) );
  AOI22_X1 U12927 ( .A1(n10395), .A2(n10394), .B1(n10393), .B2(n10392), .ZN(
        n10607) );
  XOR2_X1 U12928 ( .A(n10606), .B(n10607), .Z(n10409) );
  NAND2_X1 U12929 ( .A1(P3_REG1_REG_6__SCAN_IN), .A2(n10401), .ZN(n10397) );
  NAND2_X1 U12930 ( .A1(P3_REG1_REG_7__SCAN_IN), .A2(n10398), .ZN(n10614) );
  OAI21_X1 U12931 ( .B1(P3_REG1_REG_7__SCAN_IN), .B2(n10398), .A(n10614), .ZN(
        n10407) );
  AND2_X1 U12932 ( .A1(P3_U3151), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n11162) );
  AOI21_X1 U12933 ( .B1(n15674), .B2(P3_ADDR_REG_7__SCAN_IN), .A(n11162), .ZN(
        n10399) );
  OAI21_X1 U12934 ( .B1(n15677), .B2(n10613), .A(n10399), .ZN(n10406) );
  INV_X1 U12935 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n10402) );
  AOI21_X1 U12936 ( .B1(n10403), .B2(n10402), .A(n10600), .ZN(n10404) );
  NOR2_X1 U12937 ( .A1(n10404), .A2(n15687), .ZN(n10405) );
  AOI211_X1 U12938 ( .C1(n15679), .C2(n10407), .A(n10406), .B(n10405), .ZN(
        n10408) );
  OAI21_X1 U12939 ( .B1(n10409), .B2(n15661), .A(n10408), .ZN(P3_U3189) );
  OAI21_X1 U12940 ( .B1(n10410), .B2(P1_IR_REG_16__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n10411) );
  MUX2_X1 U12941 ( .A(P1_IR_REG_31__SCAN_IN), .B(n10411), .S(
        P1_IR_REG_17__SCAN_IN), .Z(n10412) );
  AND2_X1 U12942 ( .A1(n10412), .A2(n10719), .ZN(n14347) );
  INV_X1 U12943 ( .A(n14347), .ZN(n14364) );
  OAI222_X1 U12944 ( .A1(n14817), .A2(n10414), .B1(n14815), .B2(n10413), .C1(
        n14364), .C2(P1_U3086), .ZN(P1_U3338) );
  INV_X1 U12945 ( .A(n10794), .ZN(n15521) );
  NAND2_X1 U12946 ( .A1(n10416), .A2(n10415), .ZN(n10418) );
  XNOR2_X1 U12947 ( .A(n10794), .B(n13107), .ZN(n10631) );
  NAND2_X1 U12948 ( .A1(n13571), .A2(n11865), .ZN(n10629) );
  XNOR2_X1 U12949 ( .A(n10631), .B(n10629), .ZN(n10417) );
  NAND2_X1 U12950 ( .A1(n10418), .A2(n10417), .ZN(n10633) );
  OAI211_X1 U12951 ( .C1(n10418), .C2(n10417), .A(n10633), .B(n15123), .ZN(
        n10421) );
  AOI22_X1 U12952 ( .A1(n13701), .A2(n13572), .B1(n13570), .B2(n13555), .ZN(
        n15519) );
  NAND2_X1 U12953 ( .A1(P2_U3088), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n13584) );
  OAI21_X1 U12954 ( .B1(n13558), .B2(n15519), .A(n13584), .ZN(n10419) );
  AOI21_X1 U12955 ( .B1(n10537), .B2(n13556), .A(n10419), .ZN(n10420) );
  OAI211_X1 U12956 ( .C1(n15521), .C2(n13542), .A(n10421), .B(n10420), .ZN(
        P2_U3185) );
  NAND2_X1 U12957 ( .A1(n11286), .A2(n10424), .ZN(n10426) );
  NAND2_X1 U12958 ( .A1(n11657), .A2(n14299), .ZN(n10425) );
  OAI211_X1 U12959 ( .C1(n10435), .C2(n10427), .A(n10426), .B(n10425), .ZN(
        n11988) );
  XNOR2_X1 U12960 ( .A(n14225), .B(n11988), .ZN(n12151) );
  INV_X1 U12961 ( .A(n11988), .ZN(n15296) );
  NAND2_X1 U12962 ( .A1(n10456), .A2(n15296), .ZN(n10428) );
  NAND2_X1 U12963 ( .A1(n11837), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n10434) );
  NAND2_X1 U12964 ( .A1(n10429), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n10747) );
  OAI21_X1 U12965 ( .B1(n10429), .B2(P1_REG3_REG_6__SCAN_IN), .A(n10747), .ZN(
        n10949) );
  INV_X1 U12966 ( .A(n10949), .ZN(n10430) );
  NAND2_X1 U12967 ( .A1(n11839), .A2(n10430), .ZN(n10433) );
  NAND2_X1 U12968 ( .A1(n11808), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n10432) );
  NAND2_X1 U12969 ( .A1(n11088), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n10431) );
  NAND4_X1 U12970 ( .A1(n10434), .A2(n10433), .A3(n10432), .A4(n10431), .ZN(
        n14224) );
  AOI22_X1 U12971 ( .A1(n12110), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n11657), 
        .B2(n10436), .ZN(n10439) );
  NAND2_X1 U12972 ( .A1(n10437), .A2(n11286), .ZN(n10438) );
  NAND2_X1 U12973 ( .A1(n10439), .A2(n10438), .ZN(n15337) );
  XNOR2_X1 U12974 ( .A(n14224), .B(n15337), .ZN(n12152) );
  XNOR2_X1 U12975 ( .A(n10760), .B(n12152), .ZN(n15342) );
  AOI211_X1 U12976 ( .C1(n15337), .C2(n10590), .A(n15320), .B(n10743), .ZN(
        n15335) );
  INV_X1 U12977 ( .A(n15337), .ZN(n10758) );
  NOR2_X1 U12978 ( .A1(n15297), .A2(n10758), .ZN(n10450) );
  NAND2_X1 U12979 ( .A1(n14225), .A2(n15378), .ZN(n10445) );
  NAND2_X1 U12980 ( .A1(n11837), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n10443) );
  XNOR2_X1 U12981 ( .A(n10747), .B(P1_REG3_REG_7__SCAN_IN), .ZN(n10742) );
  NAND2_X1 U12982 ( .A1(n11839), .A2(n10742), .ZN(n10442) );
  NAND2_X1 U12983 ( .A1(n11808), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n10441) );
  NAND2_X1 U12984 ( .A1(n11088), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n10440) );
  NAND4_X1 U12985 ( .A1(n10443), .A2(n10442), .A3(n10441), .A4(n10440), .ZN(
        n14223) );
  NAND2_X1 U12986 ( .A1(n14223), .A2(n14966), .ZN(n10444) );
  NAND2_X1 U12987 ( .A1(n10445), .A2(n10444), .ZN(n15336) );
  INV_X1 U12988 ( .A(n15336), .ZN(n10447) );
  MUX2_X1 U12989 ( .A(n10447), .B(n10446), .S(n6665), .Z(n10448) );
  OAI21_X1 U12990 ( .B1(n14986), .B2(n10949), .A(n10448), .ZN(n10449) );
  AOI211_X1 U12991 ( .C1(n15335), .C2(n15299), .A(n10450), .B(n10449), .ZN(
        n10460) );
  NAND2_X1 U12992 ( .A1(n14226), .A2(n10451), .ZN(n10452) );
  NAND2_X1 U12993 ( .A1(n10453), .A2(n10452), .ZN(n10455) );
  INV_X1 U12994 ( .A(n14226), .ZN(n14061) );
  NAND2_X1 U12995 ( .A1(n14061), .A2(n11982), .ZN(n10454) );
  NAND2_X1 U12996 ( .A1(n10455), .A2(n10454), .ZN(n10587) );
  NAND2_X1 U12997 ( .A1(n10587), .A2(n12151), .ZN(n10458) );
  NAND2_X1 U12998 ( .A1(n10456), .A2(n11988), .ZN(n10457) );
  XNOR2_X1 U12999 ( .A(n10740), .B(n12152), .ZN(n15338) );
  NAND2_X1 U13000 ( .A1(n15338), .A2(n14654), .ZN(n10459) );
  OAI211_X1 U13001 ( .C1(n15342), .C2(n14982), .A(n10460), .B(n10459), .ZN(
        P1_U3287) );
  INV_X1 U13002 ( .A(n10461), .ZN(n10464) );
  OAI222_X1 U13003 ( .A1(n14938), .A2(n10464), .B1(n14936), .B2(n10463), .C1(
        P3_U3151), .C2(n10462), .ZN(P3_U3275) );
  INV_X1 U13004 ( .A(n10465), .ZN(n10466) );
  XNOR2_X1 U13005 ( .A(n15690), .B(n12234), .ZN(n10468) );
  XNOR2_X1 U13006 ( .A(n10468), .B(n12637), .ZN(n10481) );
  NAND2_X1 U13007 ( .A1(n10480), .A2(n10481), .ZN(n10479) );
  INV_X1 U13008 ( .A(n10468), .ZN(n10469) );
  OR2_X1 U13009 ( .A1(n10469), .A2(n12637), .ZN(n10471) );
  NAND2_X1 U13010 ( .A1(n10773), .A2(n15021), .ZN(n10478) );
  INV_X1 U13011 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n10659) );
  OAI22_X1 U13012 ( .A1(n15581), .A2(n15732), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n10659), .ZN(n10475) );
  NOR2_X1 U13013 ( .A1(n15009), .A2(n15019), .ZN(n12311) );
  INV_X1 U13014 ( .A(n12311), .ZN(n12349) );
  OAI22_X1 U13015 ( .A1(n10473), .A2(n12349), .B1(n12313), .B2(n10775), .ZN(
        n10474) );
  AOI211_X1 U13016 ( .C1(n15002), .C2(n10659), .A(n10475), .B(n10474), .ZN(
        n10476) );
  OAI21_X1 U13017 ( .B1(n10478), .B2(n10477), .A(n10476), .ZN(P3_U3158) );
  INV_X1 U13018 ( .A(P3_REG3_REG_2__SCAN_IN), .ZN(n10486) );
  OAI21_X1 U13019 ( .B1(n10481), .B2(n10480), .A(n10479), .ZN(n10482) );
  NAND2_X1 U13020 ( .A1(n10482), .A2(n15021), .ZN(n10485) );
  OAI22_X1 U13021 ( .A1(n7130), .A2(n15019), .B1(n10851), .B2(n15017), .ZN(
        n15694) );
  AOI22_X1 U13022 ( .A1(n15694), .A2(n15591), .B1(n10483), .B2(n15012), .ZN(
        n10484) );
  OAI211_X1 U13023 ( .C1(n10487), .C2(n10486), .A(n10485), .B(n10484), .ZN(
        P3_U3177) );
  NOR2_X1 U13024 ( .A1(P1_REG2_REG_12__SCAN_IN), .A2(n11288), .ZN(n10489) );
  NOR2_X1 U13025 ( .A1(n10489), .A2(n10488), .ZN(n10493) );
  INV_X1 U13026 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n10490) );
  MUX2_X1 U13027 ( .A(n10490), .B(P1_REG2_REG_13__SCAN_IN), .S(n11446), .Z(
        n10491) );
  INV_X1 U13028 ( .A(n10491), .ZN(n10492) );
  NAND2_X1 U13029 ( .A1(n10492), .A2(n10493), .ZN(n10509) );
  OAI211_X1 U13030 ( .C1(n10493), .C2(n10492), .A(n14377), .B(n10509), .ZN(
        n10502) );
  NAND2_X1 U13031 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3086), .ZN(n14153)
         );
  NOR2_X1 U13032 ( .A1(n11288), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n10494) );
  INV_X1 U13033 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n10496) );
  MUX2_X1 U13034 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n10496), .S(n11446), .Z(
        n10497) );
  NAND2_X1 U13035 ( .A1(n10498), .A2(n10497), .ZN(n10503) );
  OAI211_X1 U13036 ( .C1(n10498), .C2(n10497), .A(n14378), .B(n10503), .ZN(
        n10499) );
  NAND2_X1 U13037 ( .A1(n14153), .A2(n10499), .ZN(n10500) );
  AOI21_X1 U13038 ( .B1(n14360), .B2(P1_ADDR_REG_13__SCAN_IN), .A(n10500), 
        .ZN(n10501) );
  OAI211_X1 U13039 ( .C1(n15267), .C2(n10504), .A(n10502), .B(n10501), .ZN(
        P1_U3256) );
  INV_X1 U13040 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n15210) );
  AOI22_X1 U13041 ( .A1(n11451), .A2(n15210), .B1(P1_REG1_REG_14__SCAN_IN), 
        .B2(n10954), .ZN(n10506) );
  OAI21_X1 U13042 ( .B1(n10504), .B2(n10496), .A(n10503), .ZN(n10505) );
  NOR2_X1 U13043 ( .A1(n10506), .A2(n10505), .ZN(n10953) );
  AOI21_X1 U13044 ( .B1(n10506), .B2(n10505), .A(n10953), .ZN(n10517) );
  INV_X1 U13045 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n10507) );
  NAND2_X1 U13046 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n15173)
         );
  OAI21_X1 U13047 ( .B1(n15271), .B2(n10507), .A(n15173), .ZN(n10508) );
  AOI21_X1 U13048 ( .B1(n11451), .B2(n14340), .A(n10508), .ZN(n10516) );
  NAND2_X1 U13049 ( .A1(P1_REG2_REG_13__SCAN_IN), .A2(n11446), .ZN(n10510) );
  NAND2_X1 U13050 ( .A1(n10510), .A2(n10509), .ZN(n10514) );
  INV_X1 U13051 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n10511) );
  MUX2_X1 U13052 ( .A(n10511), .B(P1_REG2_REG_14__SCAN_IN), .S(n11451), .Z(
        n10512) );
  INV_X1 U13053 ( .A(n10512), .ZN(n10513) );
  NAND2_X1 U13054 ( .A1(n10513), .A2(n10514), .ZN(n10956) );
  OAI211_X1 U13055 ( .C1(n10514), .C2(n10513), .A(n14377), .B(n10956), .ZN(
        n10515) );
  OAI211_X1 U13056 ( .C1(n10517), .C2(n15264), .A(n10516), .B(n10515), .ZN(
        P1_U3257) );
  NAND3_X1 U13057 ( .A1(n15681), .A2(n10519), .A3(n10518), .ZN(n10520) );
  OAI21_X1 U13058 ( .B1(P3_STATE_REG_SCAN_IN), .B2(n9887), .A(n10520), .ZN(
        n10530) );
  NOR3_X1 U13059 ( .A1(n15679), .A2(n15082), .A3(n15681), .ZN(n10528) );
  INV_X1 U13060 ( .A(n10521), .ZN(n10527) );
  INV_X1 U13061 ( .A(n10522), .ZN(n10523) );
  AOI22_X1 U13062 ( .A1(n15679), .A2(n10523), .B1(n15674), .B2(
        P3_ADDR_REG_0__SCAN_IN), .ZN(n10526) );
  NAND2_X1 U13063 ( .A1(n15082), .A2(n10524), .ZN(n10525) );
  OAI211_X1 U13064 ( .C1(n10528), .C2(n10527), .A(n10526), .B(n10525), .ZN(
        n10529) );
  AOI211_X1 U13065 ( .C1(n15604), .C2(P3_IR_REG_0__SCAN_IN), .A(n10530), .B(
        n10529), .ZN(n10531) );
  INV_X1 U13066 ( .A(n10531), .ZN(P3_U3182) );
  NOR2_X1 U13067 ( .A1(n15507), .A2(n13573), .ZN(n10532) );
  NAND2_X1 U13068 ( .A1(n15507), .A2(n13573), .ZN(n10534) );
  XOR2_X1 U13069 ( .A(n10552), .B(n10792), .Z(n15523) );
  INV_X1 U13070 ( .A(n10537), .ZN(n10540) );
  MUX2_X1 U13071 ( .A(n15519), .B(n10538), .S(n15151), .Z(n10539) );
  OAI21_X1 U13072 ( .B1(n13865), .B2(n10540), .A(n10539), .ZN(n10542) );
  OAI211_X1 U13073 ( .C1(n10574), .C2(n15521), .A(n15144), .B(n10893), .ZN(
        n15520) );
  NOR2_X1 U13074 ( .A1(n15520), .A2(n13870), .ZN(n10541) );
  AOI211_X1 U13075 ( .C1(n15139), .C2(n10794), .A(n10542), .B(n10541), .ZN(
        n10554) );
  NAND2_X1 U13076 ( .A1(n13573), .A2(n10543), .ZN(n10544) );
  NAND2_X1 U13077 ( .A1(n10546), .A2(n15507), .ZN(n10547) );
  NAND2_X1 U13078 ( .A1(n10548), .A2(n10547), .ZN(n10566) );
  NOR2_X1 U13079 ( .A1(n15513), .A2(n13572), .ZN(n10549) );
  OR2_X1 U13080 ( .A1(n10566), .A2(n10549), .ZN(n10551) );
  NAND2_X1 U13081 ( .A1(n15513), .A2(n13572), .ZN(n10550) );
  NAND2_X1 U13082 ( .A1(n10551), .A2(n10550), .ZN(n10786) );
  XNOR2_X1 U13083 ( .A(n10786), .B(n10552), .ZN(n15526) );
  NAND2_X1 U13084 ( .A1(n15526), .A2(n15148), .ZN(n10553) );
  OAI211_X1 U13085 ( .C1(n15523), .C2(n13859), .A(n10554), .B(n10553), .ZN(
        P2_U3258) );
  INV_X1 U13086 ( .A(n10555), .ZN(n13093) );
  MUX2_X1 U13087 ( .A(n13093), .B(P2_REG2_REG_3__SCAN_IN), .S(n15151), .Z(
        n10558) );
  OAI22_X1 U13088 ( .A1(n13890), .A2(n10556), .B1(P2_REG3_REG_3__SCAN_IN), 
        .B2(n13865), .ZN(n10557) );
  AOI211_X1 U13089 ( .C1(n10559), .C2(n15147), .A(n10558), .B(n10557), .ZN(
        n10562) );
  NAND2_X1 U13090 ( .A1(n10560), .A2(n15148), .ZN(n10561) );
  OAI211_X1 U13091 ( .C1(n10563), .C2(n13859), .A(n10562), .B(n10561), .ZN(
        P2_U3262) );
  OAI222_X1 U13092 ( .A1(n14938), .A2(n10565), .B1(n14936), .B2(n10564), .C1(
        P3_U3151), .C2(n12440), .ZN(P3_U3274) );
  XNOR2_X1 U13093 ( .A(n10566), .B(n10567), .ZN(n10573) );
  INV_X1 U13094 ( .A(n10573), .ZN(n15516) );
  INV_X1 U13095 ( .A(n9794), .ZN(n15558) );
  NAND2_X1 U13096 ( .A1(n10568), .A2(n10567), .ZN(n10569) );
  AOI21_X1 U13097 ( .B1(n10570), .B2(n10569), .A(n15522), .ZN(n10571) );
  AOI211_X1 U13098 ( .C1(n15558), .C2(n10573), .A(n10572), .B(n10571), .ZN(
        n15515) );
  MUX2_X1 U13099 ( .A(n9478), .B(n15515), .S(n13852), .Z(n10580) );
  AOI211_X1 U13100 ( .C1(n15513), .C2(n10575), .A(n11865), .B(n10574), .ZN(
        n15512) );
  INV_X1 U13101 ( .A(n10576), .ZN(n10577) );
  OAI22_X1 U13102 ( .A1(n13890), .A2(n7435), .B1(n10577), .B2(n13865), .ZN(
        n10578) );
  AOI21_X1 U13103 ( .B1(n15512), .B2(n15147), .A(n10578), .ZN(n10579) );
  OAI211_X1 U13104 ( .C1(n15516), .C2(n10581), .A(n10580), .B(n10579), .ZN(
        P2_U3259) );
  INV_X1 U13105 ( .A(P3_DATAO_REG_28__SCAN_IN), .ZN(n13258) );
  NAND2_X1 U13106 ( .A1(n12245), .A2(n15577), .ZN(n10582) );
  OAI21_X1 U13107 ( .B1(n15577), .B2(n13258), .A(n10582), .ZN(P3_U3519) );
  INV_X1 U13108 ( .A(P3_DATAO_REG_29__SCAN_IN), .ZN(n13319) );
  NAND2_X1 U13109 ( .A1(n12721), .A2(n15577), .ZN(n10583) );
  OAI21_X1 U13110 ( .B1(n15577), .B2(n13319), .A(n10583), .ZN(P3_U3520) );
  INV_X1 U13111 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n13483) );
  OAI21_X1 U13112 ( .B1(n10585), .B2(n10586), .A(n7139), .ZN(n15302) );
  INV_X1 U13113 ( .A(n15302), .ZN(n10594) );
  XNOR2_X1 U13114 ( .A(n10587), .B(n10586), .ZN(n10588) );
  AOI22_X1 U13115 ( .A1(n14966), .A2(n14224), .B1(n14226), .B2(n15378), .ZN(
        n10931) );
  OAI21_X1 U13116 ( .B1(n10588), .B2(n15351), .A(n10931), .ZN(n10589) );
  AOI21_X1 U13117 ( .B1(n15345), .B2(n15302), .A(n10589), .ZN(n15305) );
  INV_X1 U13118 ( .A(n10590), .ZN(n10591) );
  AOI211_X1 U13119 ( .C1(n11988), .C2(n10592), .A(n15320), .B(n10591), .ZN(
        n15300) );
  AOI21_X1 U13120 ( .B1(n15379), .B2(n11988), .A(n15300), .ZN(n10593) );
  OAI211_X1 U13121 ( .C1(n10594), .C2(n15341), .A(n15305), .B(n10593), .ZN(
        n10596) );
  NAND2_X1 U13122 ( .A1(n10596), .A2(n15389), .ZN(n10595) );
  OAI21_X1 U13123 ( .B1(n15389), .B2(n13483), .A(n10595), .ZN(P1_U3474) );
  NAND2_X1 U13124 ( .A1(n10596), .A2(n15403), .ZN(n10597) );
  OAI21_X1 U13125 ( .B1(n15403), .B2(n6957), .A(n10597), .ZN(P1_U3533) );
  NOR2_X1 U13126 ( .A1(n10599), .A2(n10598), .ZN(n10601) );
  NAND2_X1 U13127 ( .A1(P3_REG2_REG_8__SCAN_IN), .A2(n11024), .ZN(n10602) );
  OAI21_X1 U13128 ( .B1(P3_REG2_REG_8__SCAN_IN), .B2(n11024), .A(n10602), .ZN(
        n10603) );
  AOI21_X1 U13129 ( .B1(n10604), .B2(n10603), .A(n11013), .ZN(n10623) );
  OAI22_X1 U13130 ( .A1(n10607), .A2(n10606), .B1(n10605), .B2(n10613), .ZN(
        n10609) );
  MUX2_X1 U13131 ( .A(P3_REG2_REG_8__SCAN_IN), .B(P3_REG1_REG_8__SCAN_IN), .S(
        n12696), .Z(n11025) );
  XNOR2_X1 U13132 ( .A(n11025), .B(n10611), .ZN(n10608) );
  NAND2_X1 U13133 ( .A1(n10609), .A2(n10608), .ZN(n11026) );
  OAI21_X1 U13134 ( .B1(n10609), .B2(n10608), .A(n11026), .ZN(n10610) );
  NAND2_X1 U13135 ( .A1(n10610), .A2(n15681), .ZN(n10622) );
  AOI22_X1 U13136 ( .A1(P3_REG1_REG_8__SCAN_IN), .A2(n11024), .B1(n10611), 
        .B2(n8117), .ZN(n10617) );
  NAND2_X1 U13137 ( .A1(n10613), .A2(n10612), .ZN(n10615) );
  NAND2_X1 U13138 ( .A1(n10615), .A2(n10614), .ZN(n10616) );
  NAND2_X1 U13139 ( .A1(n10617), .A2(n10616), .ZN(n11018) );
  OAI21_X1 U13140 ( .B1(n10617), .B2(n10616), .A(n11018), .ZN(n10620) );
  NAND2_X1 U13141 ( .A1(P3_U3151), .A2(P3_REG3_REG_8__SCAN_IN), .ZN(n11252) );
  NAND2_X1 U13142 ( .A1(n15674), .A2(P3_ADDR_REG_8__SCAN_IN), .ZN(n10618) );
  OAI211_X1 U13143 ( .C1(n15677), .C2(n11024), .A(n11252), .B(n10618), .ZN(
        n10619) );
  AOI21_X1 U13144 ( .B1(n10620), .B2(n15679), .A(n10619), .ZN(n10621) );
  OAI211_X1 U13145 ( .C1(n10623), .C2(n15687), .A(n10622), .B(n10621), .ZN(
        P3_U3190) );
  XNOR2_X1 U13146 ( .A(n15530), .B(n13075), .ZN(n10625) );
  NAND2_X1 U13147 ( .A1(n13570), .A2(n11865), .ZN(n10626) );
  NAND2_X1 U13148 ( .A1(n10625), .A2(n10626), .ZN(n10812) );
  INV_X1 U13149 ( .A(n10625), .ZN(n10628) );
  INV_X1 U13150 ( .A(n10626), .ZN(n10627) );
  NAND2_X1 U13151 ( .A1(n10628), .A2(n10627), .ZN(n10814) );
  NAND2_X1 U13152 ( .A1(n10812), .A2(n10814), .ZN(n10634) );
  INV_X1 U13153 ( .A(n10629), .ZN(n10630) );
  NAND2_X1 U13154 ( .A1(n10631), .A2(n10630), .ZN(n10632) );
  NAND2_X1 U13155 ( .A1(n10633), .A2(n10632), .ZN(n10813) );
  XOR2_X1 U13156 ( .A(n10634), .B(n10813), .Z(n10641) );
  NAND2_X1 U13157 ( .A1(n13571), .A2(n13701), .ZN(n10636) );
  NAND2_X1 U13158 ( .A1(n13569), .A2(n13555), .ZN(n10635) );
  AND2_X1 U13159 ( .A1(n10636), .A2(n10635), .ZN(n10899) );
  NAND2_X1 U13160 ( .A1(n13556), .A2(n10894), .ZN(n10638) );
  OAI211_X1 U13161 ( .C1(n10899), .C2(n13558), .A(n10638), .B(n10637), .ZN(
        n10639) );
  AOI21_X1 U13162 ( .B1(n15530), .B2(n15128), .A(n10639), .ZN(n10640) );
  OAI21_X1 U13163 ( .B1(n10641), .B2(n13561), .A(n10640), .ZN(P2_U3193) );
  OAI21_X1 U13164 ( .B1(n10644), .B2(n10643), .A(n10642), .ZN(n15735) );
  INV_X1 U13165 ( .A(n15735), .ZN(n10649) );
  AOI22_X1 U13166 ( .A1(n12636), .A2(n12869), .B1(n12867), .B2(n12637), .ZN(
        n10648) );
  OAI211_X1 U13167 ( .C1(n10646), .C2(n12417), .A(n10645), .B(n15695), .ZN(
        n10647) );
  OAI211_X1 U13168 ( .C1(n10649), .C2(n15766), .A(n10648), .B(n10647), .ZN(
        n15733) );
  INV_X1 U13169 ( .A(n15733), .ZN(n10664) );
  NAND2_X1 U13170 ( .A1(n13050), .A2(n10650), .ZN(n10651) );
  OAI21_X1 U13171 ( .B1(n13050), .B2(n10652), .A(n10651), .ZN(n10653) );
  INV_X1 U13172 ( .A(n10653), .ZN(n10654) );
  NAND2_X1 U13173 ( .A1(n10655), .A2(n10654), .ZN(n10658) );
  NAND2_X1 U13174 ( .A1(n10656), .A2(n15712), .ZN(n10722) );
  INV_X1 U13175 ( .A(n10722), .ZN(n15700) );
  OR2_X1 U13176 ( .A1(n15712), .A2(n15744), .ZN(n10657) );
  NOR2_X2 U13177 ( .A1(n10658), .A2(n10657), .ZN(n15097) );
  AOI22_X1 U13178 ( .A1(n15097), .A2(n10660), .B1(n12911), .B2(n10659), .ZN(
        n10661) );
  OAI21_X1 U13179 ( .B1(n8047), .B2(n15719), .A(n10661), .ZN(n10662) );
  AOI21_X1 U13180 ( .B1(n15735), .B2(n15716), .A(n10662), .ZN(n10663) );
  OAI21_X1 U13181 ( .B1(n10664), .B2(n15703), .A(n10663), .ZN(P3_U3230) );
  NOR2_X1 U13182 ( .A1(n13870), .A2(n10665), .ZN(n10670) );
  AOI22_X1 U13183 ( .A1(n15151), .A2(P2_REG2_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(n15137), .ZN(n10667) );
  OAI21_X1 U13184 ( .B1(n13890), .B2(n10668), .A(n10667), .ZN(n10669) );
  AOI211_X1 U13185 ( .C1(n15148), .C2(n10671), .A(n10670), .B(n10669), .ZN(
        n10672) );
  OAI21_X1 U13186 ( .B1(n15151), .B2(n10673), .A(n10672), .ZN(P2_U3263) );
  INV_X1 U13187 ( .A(n10674), .ZN(n10676) );
  NAND2_X1 U13188 ( .A1(n10676), .A2(n10675), .ZN(n10677) );
  NAND2_X1 U13189 ( .A1(n14227), .A2(n6664), .ZN(n10680) );
  NAND2_X1 U13190 ( .A1(n14064), .A2(n11832), .ZN(n10679) );
  NAND2_X1 U13191 ( .A1(n10680), .A2(n10679), .ZN(n10681) );
  XNOR2_X1 U13192 ( .A(n10681), .B(n11778), .ZN(n10683) );
  AND2_X1 U13193 ( .A1(n14064), .A2(n6664), .ZN(n10682) );
  AOI21_X1 U13194 ( .B1(n14227), .B2(n10688), .A(n10682), .ZN(n10684) );
  XNOR2_X1 U13195 ( .A(n10683), .B(n10684), .ZN(n14057) );
  INV_X1 U13196 ( .A(n10683), .ZN(n10686) );
  INV_X1 U13197 ( .A(n10684), .ZN(n10685) );
  NAND2_X1 U13198 ( .A1(n10686), .A2(n10685), .ZN(n10687) );
  AND2_X1 U13199 ( .A1(n11982), .A2(n6664), .ZN(n10689) );
  AOI21_X1 U13200 ( .B1(n14226), .B2(n10688), .A(n10689), .ZN(n10922) );
  NAND2_X1 U13201 ( .A1(n14226), .A2(n6664), .ZN(n10691) );
  NAND2_X1 U13202 ( .A1(n11982), .A2(n11832), .ZN(n10690) );
  NAND2_X1 U13203 ( .A1(n10691), .A2(n10690), .ZN(n10692) );
  XNOR2_X1 U13204 ( .A(n10692), .B(n11830), .ZN(n10920) );
  XNOR2_X1 U13205 ( .A(n10921), .B(n10920), .ZN(n10702) );
  NAND2_X1 U13206 ( .A1(n10694), .A2(n10693), .ZN(n10695) );
  NAND2_X1 U13207 ( .A1(n10695), .A2(P1_STATE_REG_SCAN_IN), .ZN(n15176) );
  NAND2_X1 U13208 ( .A1(n10696), .A2(n14115), .ZN(n10698) );
  AND2_X1 U13209 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n14277) );
  INV_X1 U13210 ( .A(n14277), .ZN(n10697) );
  OAI211_X1 U13211 ( .C1(n15176), .C2(n10699), .A(n10698), .B(n10697), .ZN(
        n10700) );
  AOI21_X1 U13212 ( .B1(n15172), .B2(n11982), .A(n10700), .ZN(n10701) );
  OAI21_X1 U13213 ( .B1(n10702), .B2(n15167), .A(n10701), .ZN(P1_U3230) );
  MUX2_X1 U13214 ( .A(n6813), .B(P2_REG2_REG_4__SCAN_IN), .S(n15151), .Z(
        n10708) );
  AOI22_X1 U13215 ( .A1(n15139), .A2(n10704), .B1(n10703), .B2(n15137), .ZN(
        n10705) );
  OAI21_X1 U13216 ( .B1(n13870), .B2(n10706), .A(n10705), .ZN(n10707) );
  AOI211_X1 U13217 ( .C1(n15148), .C2(n10709), .A(n10708), .B(n10707), .ZN(
        n10710) );
  OAI21_X1 U13218 ( .B1(n10711), .B2(n13859), .A(n10710), .ZN(P2_U3261) );
  INV_X1 U13219 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n10712) );
  OAI22_X1 U13220 ( .A1(n12986), .A2(n9876), .B1(n15788), .B2(n10712), .ZN(
        n10713) );
  AOI21_X1 U13221 ( .B1(n10715), .B2(n15788), .A(n10713), .ZN(n10714) );
  INV_X1 U13222 ( .A(n10714), .ZN(P3_U3459) );
  AOI21_X1 U13223 ( .B1(P3_REG3_REG_0__SCAN_IN), .B2(n12911), .A(n10715), .ZN(
        n10718) );
  AOI22_X1 U13224 ( .A1(n15703), .A2(P3_REG2_REG_0__SCAN_IN), .B1(n15097), 
        .B2(n10716), .ZN(n10717) );
  OAI21_X1 U13225 ( .B1(n10718), .B2(n15703), .A(n10717), .ZN(P3_U3233) );
  INV_X1 U13226 ( .A(n11561), .ZN(n10733) );
  NAND2_X1 U13227 ( .A1(n10719), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10720) );
  XNOR2_X1 U13228 ( .A(n10720), .B(P1_IR_REG_18__SCAN_IN), .ZN(n14372) );
  OAI222_X1 U13229 ( .A1(n14817), .A2(n10721), .B1(n14815), .B2(n10733), .C1(
        n7164), .C2(P1_U3086), .ZN(P1_U3337) );
  NAND2_X1 U13230 ( .A1(n15766), .A2(n10722), .ZN(n10723) );
  XNOR2_X1 U13231 ( .A(n10724), .B(n12468), .ZN(n15741) );
  AND2_X1 U13232 ( .A1(n10853), .A2(n10725), .ZN(n10727) );
  OAI21_X1 U13233 ( .B1(n10727), .B2(n12468), .A(n10726), .ZN(n10729) );
  INV_X1 U13234 ( .A(n12634), .ZN(n10728) );
  OAI22_X1 U13235 ( .A1(n10728), .A2(n15017), .B1(n10775), .B2(n15019), .ZN(
        n10978) );
  AOI21_X1 U13236 ( .B1(n10729), .B2(n15695), .A(n10978), .ZN(n15742) );
  MUX2_X1 U13237 ( .A(n10262), .B(n15742), .S(n15719), .Z(n10732) );
  INV_X1 U13238 ( .A(n15743), .ZN(n10730) );
  AOI22_X1 U13239 ( .A1(n15097), .A2(n10730), .B1(n12911), .B2(n10970), .ZN(
        n10731) );
  OAI211_X1 U13240 ( .C1(n12827), .C2(n15741), .A(n10732), .B(n10731), .ZN(
        P3_U3228) );
  INV_X1 U13241 ( .A(n13618), .ZN(n10734) );
  OAI222_X1 U13242 ( .A1(n14038), .A2(n10735), .B1(n10734), .B2(P2_U3088), 
        .C1(n14031), .C2(n10733), .ZN(P2_U3309) );
  NAND2_X1 U13243 ( .A1(n10736), .A2(n11286), .ZN(n10738) );
  AOI22_X1 U13244 ( .A1(n12110), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n11657), 
        .B2(n14317), .ZN(n10737) );
  NAND2_X2 U13245 ( .A1(n10738), .A2(n10737), .ZN(n11995) );
  NOR2_X1 U13246 ( .A1(n14224), .A2(n10758), .ZN(n10739) );
  NAND2_X1 U13247 ( .A1(n14224), .A2(n10758), .ZN(n10741) );
  XOR2_X1 U13248 ( .A(n12157), .B(n10845), .Z(n15352) );
  INV_X1 U13249 ( .A(n10742), .ZN(n11262) );
  OAI22_X1 U13250 ( .A1(n14969), .A2(n9742), .B1(n11262), .B2(n14986), .ZN(
        n10757) );
  INV_X1 U13251 ( .A(n10743), .ZN(n10744) );
  INV_X1 U13252 ( .A(n11995), .ZN(n11260) );
  AND2_X2 U13253 ( .A1(n10743), .A2(n11260), .ZN(n10839) );
  AOI211_X1 U13254 ( .C1(n11995), .C2(n10744), .A(n15320), .B(n10839), .ZN(
        n15349) );
  NAND2_X1 U13255 ( .A1(n14224), .A2(n15378), .ZN(n10754) );
  NAND2_X1 U13256 ( .A1(n11837), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n10752) );
  INV_X1 U13257 ( .A(n10747), .ZN(n10745) );
  AOI21_X1 U13258 ( .B1(n10745), .B2(P1_REG3_REG_7__SCAN_IN), .A(
        P1_REG3_REG_8__SCAN_IN), .ZN(n10748) );
  NAND2_X1 U13259 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_REG3_REG_7__SCAN_IN), 
        .ZN(n10746) );
  NOR2_X1 U13260 ( .A1(n10747), .A2(n10746), .ZN(n10832) );
  NAND2_X1 U13261 ( .A1(n11839), .A2(n7912), .ZN(n10751) );
  NAND2_X1 U13262 ( .A1(n6658), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n10750) );
  NAND2_X1 U13263 ( .A1(n11088), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n10749) );
  NAND4_X1 U13264 ( .A1(n10752), .A2(n10751), .A3(n10750), .A4(n10749), .ZN(
        n14222) );
  NAND2_X1 U13265 ( .A1(n14222), .A2(n14966), .ZN(n10753) );
  NAND2_X1 U13266 ( .A1(n10754), .A2(n10753), .ZN(n15347) );
  AOI21_X1 U13267 ( .B1(n15349), .B2(n7108), .A(n15347), .ZN(n10755) );
  NOR2_X1 U13268 ( .A1(n10755), .A2(n6665), .ZN(n10756) );
  AOI211_X1 U13269 ( .C1(n15282), .C2(n11995), .A(n10757), .B(n10756), .ZN(
        n10762) );
  INV_X1 U13270 ( .A(n14224), .ZN(n10759) );
  XNOR2_X1 U13271 ( .A(n10825), .B(n12157), .ZN(n15354) );
  NAND2_X1 U13272 ( .A1(n15354), .A2(n15191), .ZN(n10761) );
  OAI211_X1 U13273 ( .C1(n15352), .C2(n14599), .A(n10762), .B(n10761), .ZN(
        P1_U3286) );
  INV_X1 U13274 ( .A(n11656), .ZN(n10769) );
  OAI222_X1 U13275 ( .A1(n14031), .A2(n10769), .B1(n10763), .B2(P2_U3088), 
        .C1(n13423), .C2(n14038), .ZN(P2_U3308) );
  NOR2_X1 U13276 ( .A1(n14936), .A2(SI_22_), .ZN(n10764) );
  AOI21_X1 U13277 ( .B1(n10765), .B2(P3_STATE_REG_SCAN_IN), .A(n10764), .ZN(
        n10766) );
  OAI21_X1 U13278 ( .B1(n10767), .B2(n14938), .A(n10766), .ZN(n10768) );
  INV_X1 U13279 ( .A(n10768), .ZN(P3_U3273) );
  OAI222_X1 U13280 ( .A1(n14817), .A2(n10770), .B1(n14815), .B2(n10769), .C1(
        n7108), .C2(P1_U3086), .ZN(P1_U3336) );
  NAND2_X1 U13281 ( .A1(n8394), .A2(n10771), .ZN(n10772) );
  XNOR2_X1 U13282 ( .A(n15736), .B(n12270), .ZN(n10774) );
  NAND2_X1 U13283 ( .A1(n10775), .A2(n10774), .ZN(n10971) );
  OAI21_X1 U13284 ( .B1(n10775), .B2(n10774), .A(n10971), .ZN(n10777) );
  INV_X1 U13285 ( .A(n10972), .ZN(n10776) );
  AOI21_X1 U13286 ( .B1(n10778), .B2(n10777), .A(n10776), .ZN(n10784) );
  OAI22_X1 U13287 ( .A1(n10851), .A2(n12349), .B1(n12313), .B2(n11050), .ZN(
        n10779) );
  AOI211_X1 U13288 ( .C1(n15736), .C2(n15012), .A(n10780), .B(n10779), .ZN(
        n10783) );
  INV_X1 U13289 ( .A(n10781), .ZN(n10860) );
  NAND2_X1 U13290 ( .A1(n15002), .A2(n10860), .ZN(n10782) );
  OAI211_X1 U13291 ( .C1(n10784), .C2(n15585), .A(n10783), .B(n10782), .ZN(
        P3_U3170) );
  AND2_X1 U13292 ( .A1(n10794), .A2(n13571), .ZN(n10785) );
  OR2_X1 U13293 ( .A1(n10794), .A2(n13571), .ZN(n10787) );
  OR2_X1 U13294 ( .A1(n10789), .A2(n10798), .ZN(n10790) );
  NAND2_X1 U13295 ( .A1(n10987), .A2(n10790), .ZN(n15541) );
  OR2_X1 U13296 ( .A1(n10794), .A2(n10793), .ZN(n10791) );
  NAND2_X1 U13297 ( .A1(n10794), .A2(n10793), .ZN(n10795) );
  AND2_X1 U13298 ( .A1(n15530), .A2(n10796), .ZN(n10797) );
  XNOR2_X1 U13299 ( .A(n10991), .B(n10798), .ZN(n10799) );
  NAND2_X1 U13300 ( .A1(n10799), .A2(n15551), .ZN(n10802) );
  NAND2_X1 U13301 ( .A1(n13570), .A2(n13701), .ZN(n10801) );
  NAND2_X1 U13302 ( .A1(n13568), .A2(n13555), .ZN(n10800) );
  AND2_X1 U13303 ( .A1(n10801), .A2(n10800), .ZN(n10821) );
  NAND2_X1 U13304 ( .A1(n10802), .A2(n10821), .ZN(n15543) );
  NAND2_X1 U13305 ( .A1(n15543), .A2(n13852), .ZN(n10806) );
  AOI211_X1 U13306 ( .C1(n15538), .C2(n10891), .A(n11865), .B(n10993), .ZN(
        n15537) );
  INV_X1 U13307 ( .A(n15538), .ZN(n10989) );
  AOI22_X1 U13308 ( .A1(n15151), .A2(P2_REG2_REG_9__SCAN_IN), .B1(n10819), 
        .B2(n15137), .ZN(n10803) );
  OAI21_X1 U13309 ( .B1(n13890), .B2(n10989), .A(n10803), .ZN(n10804) );
  AOI21_X1 U13310 ( .B1(n15537), .B2(n15147), .A(n10804), .ZN(n10805) );
  OAI211_X1 U13311 ( .C1(n13874), .C2(n15541), .A(n10806), .B(n10805), .ZN(
        P2_U3256) );
  XNOR2_X1 U13312 ( .A(n15538), .B(n13075), .ZN(n10807) );
  NAND2_X1 U13313 ( .A1(n13569), .A2(n11865), .ZN(n10808) );
  NAND2_X1 U13314 ( .A1(n10807), .A2(n10808), .ZN(n10904) );
  INV_X1 U13315 ( .A(n10807), .ZN(n10810) );
  INV_X1 U13316 ( .A(n10808), .ZN(n10809) );
  NAND2_X1 U13317 ( .A1(n10810), .A2(n10809), .ZN(n10811) );
  NAND2_X1 U13318 ( .A1(n10904), .A2(n10811), .ZN(n10818) );
  NAND2_X1 U13319 ( .A1(n10813), .A2(n10812), .ZN(n10815) );
  NAND2_X1 U13320 ( .A1(n10815), .A2(n10814), .ZN(n10817) );
  INV_X1 U13321 ( .A(n10905), .ZN(n10816) );
  AOI21_X1 U13322 ( .B1(n10818), .B2(n10817), .A(n10816), .ZN(n10824) );
  NAND2_X1 U13323 ( .A1(n13556), .A2(n10819), .ZN(n10820) );
  NAND2_X1 U13324 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3088), .ZN(n13611) );
  OAI211_X1 U13325 ( .C1(n10821), .C2(n13558), .A(n10820), .B(n13611), .ZN(
        n10822) );
  AOI21_X1 U13326 ( .B1(n15538), .B2(n15128), .A(n10822), .ZN(n10823) );
  OAI21_X1 U13327 ( .B1(n10824), .B2(n13561), .A(n10823), .ZN(P2_U3203) );
  NAND2_X1 U13328 ( .A1(n11260), .A2(n10842), .ZN(n10826) );
  NAND2_X1 U13329 ( .A1(n10827), .A2(n10826), .ZN(n11062) );
  NAND2_X1 U13330 ( .A1(n10828), .A2(n11286), .ZN(n10831) );
  AOI22_X1 U13331 ( .A1(n12110), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n11657), 
        .B2(n10829), .ZN(n10830) );
  INV_X1 U13332 ( .A(n14222), .ZN(n11096) );
  XNOR2_X1 U13333 ( .A(n11998), .B(n11096), .ZN(n12156) );
  XNOR2_X1 U13334 ( .A(n11062), .B(n12156), .ZN(n15363) );
  INV_X1 U13335 ( .A(n15363), .ZN(n10849) );
  NAND2_X1 U13336 ( .A1(n11837), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n10837) );
  NAND2_X1 U13337 ( .A1(n10832), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n11076) );
  OR2_X1 U13338 ( .A1(n10832), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n10833) );
  AND2_X1 U13339 ( .A1(n11076), .A2(n10833), .ZN(n15281) );
  NAND2_X1 U13340 ( .A1(n11839), .A2(n15281), .ZN(n10836) );
  NAND2_X1 U13341 ( .A1(n6658), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n10835) );
  NAND2_X1 U13342 ( .A1(n11088), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n10834) );
  NAND4_X1 U13343 ( .A1(n10837), .A2(n10836), .A3(n10835), .A4(n10834), .ZN(
        n15377) );
  AOI22_X1 U13344 ( .A1(n14966), .A2(n15377), .B1(n14223), .B2(n15378), .ZN(
        n15356) );
  AOI22_X1 U13345 ( .A1(n6665), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n7912), .B2(
        n15293), .ZN(n10838) );
  OAI21_X1 U13346 ( .B1(n15356), .B2(n6665), .A(n10838), .ZN(n10841) );
  INV_X1 U13347 ( .A(n11998), .ZN(n15358) );
  NAND2_X1 U13348 ( .A1(n10839), .A2(n15358), .ZN(n15285) );
  OAI211_X1 U13349 ( .C1(n10839), .C2(n15358), .A(n15288), .B(n15285), .ZN(
        n15357) );
  NOR2_X1 U13350 ( .A1(n15357), .A2(n14550), .ZN(n10840) );
  AOI211_X1 U13351 ( .C1(n15282), .C2(n11998), .A(n10841), .B(n10840), .ZN(
        n10848) );
  NOR2_X1 U13352 ( .A1(n10842), .A2(n11995), .ZN(n10844) );
  NAND2_X1 U13353 ( .A1(n10842), .A2(n11995), .ZN(n10843) );
  NAND2_X1 U13354 ( .A1(n10846), .A2(n12156), .ZN(n15359) );
  NAND3_X1 U13355 ( .A1(n15360), .A2(n15359), .A3(n14654), .ZN(n10847) );
  OAI211_X1 U13356 ( .C1(n10849), .C2(n14982), .A(n10848), .B(n10847), .ZN(
        P1_U3285) );
  XNOR2_X1 U13357 ( .A(n10850), .B(n10856), .ZN(n15737) );
  INV_X1 U13358 ( .A(n15737), .ZN(n10863) );
  INV_X1 U13359 ( .A(n15716), .ZN(n11060) );
  INV_X1 U13360 ( .A(n15766), .ZN(n15760) );
  OAI22_X1 U13361 ( .A1(n11050), .A2(n15017), .B1(n10851), .B2(n15019), .ZN(
        n10858) );
  INV_X1 U13362 ( .A(n10852), .ZN(n10855) );
  INV_X1 U13363 ( .A(n10853), .ZN(n10854) );
  AOI211_X1 U13364 ( .C1(n10856), .C2(n10855), .A(n15708), .B(n10854), .ZN(
        n10857) );
  AOI211_X1 U13365 ( .C1(n15737), .C2(n15760), .A(n10858), .B(n10857), .ZN(
        n15739) );
  MUX2_X1 U13366 ( .A(n10859), .B(n15739), .S(n15719), .Z(n10862) );
  AOI22_X1 U13367 ( .A1(n15097), .A2(n15736), .B1(n12911), .B2(n10860), .ZN(
        n10861) );
  OAI211_X1 U13368 ( .C1(n10863), .C2(n11060), .A(n10862), .B(n10861), .ZN(
        P3_U3229) );
  NAND2_X1 U13369 ( .A1(n10865), .A2(n10864), .ZN(n10867) );
  NAND2_X1 U13370 ( .A1(n10879), .A2(n10868), .ZN(n10869) );
  NAND2_X1 U13371 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n15475), .ZN(n15473) );
  NAND2_X1 U13372 ( .A1(n10869), .A2(n15473), .ZN(n10874) );
  INV_X1 U13373 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n10872) );
  NAND2_X1 U13374 ( .A1(n10870), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n11110) );
  INV_X1 U13375 ( .A(n11110), .ZN(n10871) );
  AOI21_X1 U13376 ( .B1(n10872), .B2(n11106), .A(n10871), .ZN(n10873) );
  NAND2_X1 U13377 ( .A1(n10873), .A2(n10874), .ZN(n11109) );
  OAI211_X1 U13378 ( .C1(n10874), .C2(n10873), .A(n15474), .B(n11109), .ZN(
        n10887) );
  NAND2_X1 U13379 ( .A1(P2_U3088), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n13512)
         );
  INV_X1 U13380 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n10876) );
  OAI22_X1 U13381 ( .A1(n10878), .A2(n10877), .B1(n10876), .B2(n10875), .ZN(
        n10880) );
  NAND2_X1 U13382 ( .A1(n10879), .A2(n10880), .ZN(n10881) );
  XNOR2_X1 U13383 ( .A(n10880), .B(n15478), .ZN(n15468) );
  NAND2_X1 U13384 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n15468), .ZN(n15466) );
  NAND2_X1 U13385 ( .A1(n10881), .A2(n15466), .ZN(n10883) );
  XNOR2_X1 U13386 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n11106), .ZN(n10882) );
  NAND2_X1 U13387 ( .A1(n10882), .A2(n10883), .ZN(n11104) );
  OAI211_X1 U13388 ( .C1(n10883), .C2(n10882), .A(n15467), .B(n11104), .ZN(
        n10884) );
  NAND2_X1 U13389 ( .A1(n13512), .A2(n10884), .ZN(n10885) );
  AOI21_X1 U13390 ( .B1(n15472), .B2(P2_ADDR_REG_16__SCAN_IN), .A(n10885), 
        .ZN(n10886) );
  OAI211_X1 U13391 ( .C1(n15479), .C2(n11106), .A(n10887), .B(n10886), .ZN(
        P2_U3230) );
  INV_X1 U13392 ( .A(n11674), .ZN(n11861) );
  OAI222_X1 U13393 ( .A1(n14817), .A2(n10888), .B1(n14815), .B2(n11861), .C1(
        n12130), .C2(P1_U3086), .ZN(P1_U3335) );
  AOI21_X1 U13394 ( .B1(n10890), .B2(n10889), .A(n6808), .ZN(n15535) );
  INV_X1 U13395 ( .A(n15535), .ZN(n15532) );
  INV_X1 U13396 ( .A(n10891), .ZN(n10892) );
  AOI211_X1 U13397 ( .C1(n15530), .C2(n10893), .A(n11865), .B(n10892), .ZN(
        n15529) );
  INV_X1 U13398 ( .A(n10894), .ZN(n10895) );
  OAI22_X1 U13399 ( .A1(n13890), .A2(n7447), .B1(n10895), .B2(n13865), .ZN(
        n10896) );
  AOI21_X1 U13400 ( .B1(n15529), .B2(n15147), .A(n10896), .ZN(n10903) );
  XNOR2_X1 U13401 ( .A(n10898), .B(n10897), .ZN(n10900) );
  OAI21_X1 U13402 ( .B1(n10900), .B2(n15522), .A(n10899), .ZN(n15534) );
  INV_X1 U13403 ( .A(n15534), .ZN(n10901) );
  MUX2_X1 U13404 ( .A(n9480), .B(n10901), .S(n13852), .Z(n10902) );
  OAI211_X1 U13405 ( .C1(n15532), .C2(n13874), .A(n10903), .B(n10902), .ZN(
        P2_U3257) );
  XNOR2_X1 U13406 ( .A(n11229), .B(n13075), .ZN(n11003) );
  NAND2_X1 U13407 ( .A1(n13568), .A2(n11865), .ZN(n11004) );
  XNOR2_X1 U13408 ( .A(n11003), .B(n11004), .ZN(n11001) );
  XNOR2_X1 U13409 ( .A(n11002), .B(n11001), .ZN(n10910) );
  AOI22_X1 U13410 ( .A1(n13555), .A2(n13567), .B1(n13569), .B2(n13701), .ZN(
        n15546) );
  NAND2_X1 U13411 ( .A1(n13556), .A2(n10994), .ZN(n10907) );
  OAI211_X1 U13412 ( .C1(n15546), .C2(n13558), .A(n10907), .B(n10906), .ZN(
        n10908) );
  AOI21_X1 U13413 ( .B1(n11229), .B2(n15128), .A(n10908), .ZN(n10909) );
  OAI21_X1 U13414 ( .B1(n10910), .B2(n13561), .A(n10909), .ZN(P2_U3189) );
  NAND2_X1 U13415 ( .A1(n14225), .A2(n6664), .ZN(n10912) );
  NAND2_X1 U13416 ( .A1(n11988), .A2(n11832), .ZN(n10911) );
  NAND2_X1 U13417 ( .A1(n10912), .A2(n10911), .ZN(n10913) );
  XNOR2_X1 U13418 ( .A(n10913), .B(n11778), .ZN(n10915) );
  AND2_X1 U13419 ( .A1(n11988), .A2(n6664), .ZN(n10914) );
  AOI21_X1 U13420 ( .B1(n14225), .B2(n10688), .A(n10914), .ZN(n10916) );
  NAND2_X1 U13421 ( .A1(n10915), .A2(n10916), .ZN(n10935) );
  INV_X1 U13422 ( .A(n10915), .ZN(n10918) );
  INV_X1 U13423 ( .A(n10916), .ZN(n10917) );
  NAND2_X1 U13424 ( .A1(n10918), .A2(n10917), .ZN(n10919) );
  NAND2_X1 U13425 ( .A1(n10935), .A2(n10919), .ZN(n10929) );
  INV_X1 U13426 ( .A(n10922), .ZN(n10923) );
  NAND2_X1 U13427 ( .A1(n10924), .A2(n10923), .ZN(n10925) );
  INV_X1 U13428 ( .A(n10936), .ZN(n10927) );
  AOI21_X1 U13429 ( .B1(n10929), .B2(n10928), .A(n10927), .ZN(n10934) );
  NAND2_X1 U13430 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n14293) );
  INV_X1 U13431 ( .A(n15176), .ZN(n14208) );
  NAND2_X1 U13432 ( .A1(n14208), .A2(n15294), .ZN(n10930) );
  OAI211_X1 U13433 ( .C1(n10931), .C2(n14200), .A(n14293), .B(n10930), .ZN(
        n10932) );
  AOI21_X1 U13434 ( .B1(n15172), .B2(n11988), .A(n10932), .ZN(n10933) );
  OAI21_X1 U13435 ( .B1(n10934), .B2(n15167), .A(n10933), .ZN(P1_U3227) );
  NAND2_X1 U13436 ( .A1(n14224), .A2(n6664), .ZN(n10938) );
  NAND2_X1 U13437 ( .A1(n15337), .A2(n11832), .ZN(n10937) );
  NAND2_X1 U13438 ( .A1(n10938), .A2(n10937), .ZN(n10939) );
  XNOR2_X1 U13439 ( .A(n10939), .B(n11830), .ZN(n10942) );
  NAND2_X1 U13440 ( .A1(n14224), .A2(n10688), .ZN(n10941) );
  NAND2_X1 U13441 ( .A1(n15337), .A2(n6664), .ZN(n10940) );
  NAND2_X1 U13442 ( .A1(n10941), .A2(n10940), .ZN(n10943) );
  NAND2_X1 U13443 ( .A1(n10942), .A2(n10943), .ZN(n11268) );
  INV_X1 U13444 ( .A(n10942), .ZN(n10945) );
  INV_X1 U13445 ( .A(n10943), .ZN(n10944) );
  NAND2_X1 U13446 ( .A1(n10945), .A2(n10944), .ZN(n11270) );
  NAND2_X1 U13447 ( .A1(n11268), .A2(n11270), .ZN(n10946) );
  XNOR2_X1 U13448 ( .A(n11269), .B(n10946), .ZN(n10952) );
  NAND2_X1 U13449 ( .A1(n15336), .A2(n14115), .ZN(n10948) );
  OAI211_X1 U13450 ( .C1(n15176), .C2(n10949), .A(n10948), .B(n10947), .ZN(
        n10950) );
  AOI21_X1 U13451 ( .B1(n15172), .B2(n15337), .A(n10950), .ZN(n10951) );
  OAI21_X1 U13452 ( .B1(n10952), .B2(n15167), .A(n10951), .ZN(P1_U3239) );
  XNOR2_X1 U13453 ( .A(n11614), .B(n11215), .ZN(n10955) );
  NOR2_X1 U13454 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(n10955), .ZN(n11216) );
  AOI21_X1 U13455 ( .B1(P1_REG1_REG_15__SCAN_IN), .B2(n10955), .A(n11216), 
        .ZN(n10966) );
  NAND2_X1 U13456 ( .A1(n11451), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n10957) );
  NAND2_X1 U13457 ( .A1(n10957), .A2(n10956), .ZN(n11208) );
  XNOR2_X1 U13458 ( .A(n11614), .B(n11208), .ZN(n10958) );
  NOR2_X1 U13459 ( .A1(P1_REG2_REG_15__SCAN_IN), .A2(n10958), .ZN(n11209) );
  AOI21_X1 U13460 ( .B1(P1_REG2_REG_15__SCAN_IN), .B2(n10958), .A(n11209), 
        .ZN(n10959) );
  OR2_X1 U13461 ( .A1(n10959), .A2(n15266), .ZN(n10962) );
  NOR2_X1 U13462 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n13404), .ZN(n10960) );
  AOI21_X1 U13463 ( .B1(n14360), .B2(P1_ADDR_REG_15__SCAN_IN), .A(n10960), 
        .ZN(n10961) );
  OAI211_X1 U13464 ( .C1(n15267), .C2(n10963), .A(n10962), .B(n10961), .ZN(
        n10964) );
  INV_X1 U13465 ( .A(n10964), .ZN(n10965) );
  OAI21_X1 U13466 ( .B1(n10966), .B2(n15264), .A(n10965), .ZN(P1_U3258) );
  NAND2_X1 U13467 ( .A1(n10967), .A2(n14945), .ZN(n10968) );
  OAI211_X1 U13468 ( .C1(n10969), .C2(n14936), .A(n10968), .B(n12615), .ZN(
        P3_U3272) );
  INV_X1 U13469 ( .A(n10970), .ZN(n10981) );
  XNOR2_X1 U13470 ( .A(n12234), .B(n15743), .ZN(n11039) );
  XNOR2_X1 U13471 ( .A(n11039), .B(n12635), .ZN(n10974) );
  OAI21_X1 U13472 ( .B1(n10974), .B2(n10973), .A(n11124), .ZN(n10975) );
  NAND2_X1 U13473 ( .A1(n10975), .A2(n15021), .ZN(n10980) );
  OAI21_X1 U13474 ( .B1(n15581), .B2(n15743), .A(n10976), .ZN(n10977) );
  AOI21_X1 U13475 ( .B1(n10978), .B2(n15591), .A(n10977), .ZN(n10979) );
  OAI211_X1 U13476 ( .C1(n10981), .C2(n15593), .A(n10980), .B(n10979), .ZN(
        P3_U3167) );
  INV_X1 U13477 ( .A(n11696), .ZN(n10984) );
  OAI222_X1 U13478 ( .A1(n14817), .A2(n10982), .B1(n14815), .B2(n10984), .C1(
        P1_U3086), .C2(n12141), .ZN(P1_U3334) );
  OAI222_X1 U13479 ( .A1(n14038), .A2(n10985), .B1(n14031), .B2(n10984), .C1(
        P2_U3088), .C2(n10983), .ZN(P2_U3306) );
  NAND2_X1 U13480 ( .A1(n15538), .A2(n13569), .ZN(n10986) );
  XOR2_X1 U13481 ( .A(n10992), .B(n11225), .Z(n15555) );
  NAND2_X1 U13482 ( .A1(n15538), .A2(n10988), .ZN(n10990) );
  AOI22_X1 U13483 ( .A1(n10991), .A2(n10990), .B1(n10989), .B2(n13569), .ZN(
        n11228) );
  XNOR2_X1 U13484 ( .A(n11228), .B(n10992), .ZN(n15552) );
  INV_X1 U13485 ( .A(n11235), .ZN(n11236) );
  OAI211_X1 U13486 ( .C1(n15549), .C2(n10993), .A(n11236), .B(n15144), .ZN(
        n15547) );
  INV_X1 U13487 ( .A(n10994), .ZN(n10995) );
  OAI22_X1 U13488 ( .A1(n15151), .A2(n15546), .B1(n10995), .B2(n13865), .ZN(
        n10997) );
  NOR2_X1 U13489 ( .A1(n15549), .A2(n13890), .ZN(n10996) );
  AOI211_X1 U13490 ( .C1(n15151), .C2(P2_REG2_REG_10__SCAN_IN), .A(n10997), 
        .B(n10996), .ZN(n10998) );
  OAI21_X1 U13491 ( .B1(n15547), .B2(n13870), .A(n10998), .ZN(n10999) );
  AOI21_X1 U13492 ( .B1(n15552), .B2(n13872), .A(n10999), .ZN(n11000) );
  OAI21_X1 U13493 ( .B1(n15555), .B2(n13874), .A(n11000), .ZN(P2_U3255) );
  INV_X1 U13494 ( .A(n11003), .ZN(n11006) );
  INV_X1 U13495 ( .A(n11004), .ZN(n11005) );
  XNOR2_X1 U13496 ( .A(n11323), .B(n13107), .ZN(n11177) );
  NAND2_X1 U13497 ( .A1(n13567), .A2(n11865), .ZN(n11175) );
  XNOR2_X1 U13498 ( .A(n11177), .B(n11175), .ZN(n11178) );
  XNOR2_X1 U13499 ( .A(n11179), .B(n11178), .ZN(n11012) );
  NAND2_X1 U13500 ( .A1(n13568), .A2(n13701), .ZN(n11008) );
  NAND2_X1 U13501 ( .A1(n13566), .A2(n13555), .ZN(n11007) );
  AND2_X1 U13502 ( .A1(n11008), .A2(n11007), .ZN(n11232) );
  OAI22_X1 U13503 ( .A1(n13558), .A2(n11232), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8783), .ZN(n11010) );
  INV_X1 U13504 ( .A(n11323), .ZN(n11395) );
  NOR2_X1 U13505 ( .A1(n11395), .A2(n13542), .ZN(n11009) );
  AOI211_X1 U13506 ( .C1(n13556), .C2(n11393), .A(n11010), .B(n11009), .ZN(
        n11011) );
  OAI21_X1 U13507 ( .B1(n11012), .B2(n13561), .A(n11011), .ZN(P2_U3208) );
  NOR2_X1 U13508 ( .A1(n15605), .A2(n11014), .ZN(n11015) );
  INV_X1 U13509 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n15600) );
  AOI22_X1 U13510 ( .A1(n12679), .A2(P3_REG2_REG_10__SCAN_IN), .B1(n11343), 
        .B2(n12655), .ZN(n11016) );
  OAI221_X1 U13511 ( .B1(n12654), .B2(n11017), .C1(n12654), .C2(n11016), .A(
        n15082), .ZN(n11038) );
  AOI22_X1 U13512 ( .A1(n12679), .A2(n8143), .B1(P3_REG1_REG_10__SCAN_IN), 
        .B2(n12655), .ZN(n11023) );
  NAND2_X1 U13513 ( .A1(P3_REG1_REG_8__SCAN_IN), .A2(n11024), .ZN(n11019) );
  NAND2_X1 U13514 ( .A1(n11019), .A2(n11018), .ZN(n11020) );
  NAND2_X1 U13515 ( .A1(n14928), .A2(n11020), .ZN(n11021) );
  XNOR2_X1 U13516 ( .A(n15605), .B(n11020), .ZN(n15603) );
  NAND2_X1 U13517 ( .A1(P3_REG1_REG_9__SCAN_IN), .A2(n15603), .ZN(n15602) );
  NAND2_X1 U13518 ( .A1(n11021), .A2(n15602), .ZN(n11022) );
  NAND2_X1 U13519 ( .A1(n11023), .A2(n11022), .ZN(n12642) );
  OAI21_X1 U13520 ( .B1(n11023), .B2(n11022), .A(n12642), .ZN(n11036) );
  OR2_X1 U13521 ( .A1(n11025), .A2(n11024), .ZN(n11027) );
  INV_X1 U13522 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n11370) );
  MUX2_X1 U13523 ( .A(n15600), .B(n11370), .S(n12694), .Z(n11028) );
  OR2_X1 U13524 ( .A1(n11028), .A2(n15605), .ZN(n15595) );
  NAND2_X1 U13525 ( .A1(n11028), .A2(n15605), .ZN(n15596) );
  INV_X1 U13526 ( .A(n15596), .ZN(n11029) );
  MUX2_X1 U13527 ( .A(P3_REG2_REG_10__SCAN_IN), .B(P3_REG1_REG_10__SCAN_IN), 
        .S(n12694), .Z(n12676) );
  XNOR2_X1 U13528 ( .A(n12676), .B(n12655), .ZN(n11030) );
  AOI21_X1 U13529 ( .B1(n11031), .B2(n11030), .A(n12677), .ZN(n11034) );
  INV_X1 U13530 ( .A(P3_ADDR_REG_10__SCAN_IN), .ZN(n14840) );
  NAND2_X1 U13531 ( .A1(P3_REG3_REG_10__SCAN_IN), .A2(P3_U3151), .ZN(n15579)
         );
  OAI21_X1 U13532 ( .B1(n15613), .B2(n14840), .A(n15579), .ZN(n11032) );
  AOI21_X1 U13533 ( .B1(n12679), .B2(n15604), .A(n11032), .ZN(n11033) );
  OAI21_X1 U13534 ( .B1(n11034), .B2(n15661), .A(n11033), .ZN(n11035) );
  AOI21_X1 U13535 ( .B1(n11036), .B2(n15679), .A(n11035), .ZN(n11037) );
  NAND2_X1 U13536 ( .A1(n11038), .A2(n11037), .ZN(P3_U3192) );
  INV_X1 U13537 ( .A(n11057), .ZN(n11048) );
  INV_X1 U13538 ( .A(n11039), .ZN(n11040) );
  OR2_X1 U13539 ( .A1(n11040), .A2(n12635), .ZN(n11121) );
  AND2_X1 U13540 ( .A1(n11124), .A2(n11121), .ZN(n11043) );
  XNOR2_X1 U13541 ( .A(n11041), .B(n12270), .ZN(n11125) );
  XOR2_X1 U13542 ( .A(n11125), .B(n12634), .Z(n11042) );
  NAND2_X1 U13543 ( .A1(n11043), .A2(n11042), .ZN(n11158) );
  OAI211_X1 U13544 ( .C1(n11043), .C2(n11042), .A(n11158), .B(n15021), .ZN(
        n11047) );
  OAI22_X1 U13545 ( .A1(n11050), .A2(n12349), .B1(n12313), .B2(n11144), .ZN(
        n11044) );
  AOI211_X1 U13546 ( .C1(n15749), .C2(n15012), .A(n11045), .B(n11044), .ZN(
        n11046) );
  OAI211_X1 U13547 ( .C1(n11048), .C2(n15593), .A(n11047), .B(n11046), .ZN(
        P3_U3179) );
  XNOR2_X1 U13548 ( .A(n11049), .B(n12412), .ZN(n15751) );
  INV_X1 U13549 ( .A(n15751), .ZN(n11061) );
  INV_X1 U13550 ( .A(P3_REG2_REG_6__SCAN_IN), .ZN(n11056) );
  OAI22_X1 U13551 ( .A1(n11050), .A2(n15019), .B1(n11144), .B2(n15017), .ZN(
        n11055) );
  INV_X1 U13552 ( .A(n11051), .ZN(n11052) );
  AOI211_X1 U13553 ( .C1(n12412), .C2(n11053), .A(n15708), .B(n11052), .ZN(
        n11054) );
  AOI211_X1 U13554 ( .C1(n15751), .C2(n15760), .A(n11055), .B(n11054), .ZN(
        n15753) );
  MUX2_X1 U13555 ( .A(n11056), .B(n15753), .S(n15719), .Z(n11059) );
  AOI22_X1 U13556 ( .A1(n15097), .A2(n15749), .B1(n12911), .B2(n11057), .ZN(
        n11058) );
  OAI211_X1 U13557 ( .C1(n11061), .C2(n11060), .A(n11059), .B(n11058), .ZN(
        P3_U3227) );
  NAND2_X1 U13558 ( .A1(n11062), .A2(n12156), .ZN(n11064) );
  OR2_X1 U13559 ( .A1(n11998), .A2(n14222), .ZN(n11063) );
  NAND2_X1 U13560 ( .A1(n11064), .A2(n11063), .ZN(n15277) );
  NAND2_X1 U13561 ( .A1(n11065), .A2(n11286), .ZN(n11067) );
  AOI22_X1 U13562 ( .A1(n12110), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n11657), 
        .B2(n14339), .ZN(n11066) );
  XNOR2_X1 U13563 ( .A(n15286), .B(n15377), .ZN(n15276) );
  INV_X1 U13564 ( .A(n15276), .ZN(n11068) );
  NAND2_X1 U13565 ( .A1(n15277), .A2(n11068), .ZN(n11070) );
  OR2_X1 U13566 ( .A1(n15286), .A2(n15377), .ZN(n11069) );
  NAND2_X1 U13567 ( .A1(n11070), .A2(n11069), .ZN(n11312) );
  NAND2_X1 U13568 ( .A1(n11071), .A2(n11286), .ZN(n11074) );
  AOI22_X1 U13569 ( .A1(n12110), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n11657), 
        .B2(n11072), .ZN(n11073) );
  NAND2_X1 U13570 ( .A1(n11837), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n11081) );
  INV_X1 U13571 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n11075) );
  NAND2_X1 U13572 ( .A1(n11076), .A2(n11075), .ZN(n11077) );
  AND2_X1 U13573 ( .A1(n11086), .A2(n11077), .ZN(n11553) );
  NAND2_X1 U13574 ( .A1(n11839), .A2(n11553), .ZN(n11080) );
  NAND2_X1 U13575 ( .A1(n11088), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n11079) );
  NAND2_X1 U13576 ( .A1(n11808), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n11078) );
  NAND4_X1 U13577 ( .A1(n11081), .A2(n11080), .A3(n11079), .A4(n11078), .ZN(
        n14221) );
  INV_X1 U13578 ( .A(n14221), .ZN(n11082) );
  OR2_X1 U13579 ( .A1(n15380), .A2(n11082), .ZN(n11280) );
  NAND2_X1 U13580 ( .A1(n15380), .A2(n11082), .ZN(n11083) );
  XNOR2_X1 U13581 ( .A(n11312), .B(n12158), .ZN(n15385) );
  INV_X1 U13582 ( .A(n15385), .ZN(n11103) );
  OR2_X1 U13583 ( .A1(n6665), .A2(n15212), .ZN(n14978) );
  INV_X1 U13584 ( .A(n15377), .ZN(n11556) );
  AOI22_X1 U13585 ( .A1(n6665), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n11553), 
        .B2(n15293), .ZN(n11084) );
  OAI21_X1 U13586 ( .B1(n14978), .B2(n11556), .A(n11084), .ZN(n11095) );
  XOR2_X1 U13587 ( .A(n15380), .B(n15287), .Z(n11093) );
  INV_X1 U13588 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n11085) );
  NAND2_X1 U13589 ( .A1(n11086), .A2(n11085), .ZN(n11087) );
  AND2_X1 U13590 ( .A1(n11292), .A2(n11087), .ZN(n15182) );
  NAND2_X1 U13591 ( .A1(n11839), .A2(n15182), .ZN(n11092) );
  NAND2_X1 U13592 ( .A1(n12112), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n11091) );
  NAND2_X1 U13593 ( .A1(n12113), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n11090) );
  NAND2_X1 U13594 ( .A1(n11808), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n11089) );
  NAND4_X1 U13595 ( .A1(n11092), .A2(n11091), .A3(n11090), .A4(n11089), .ZN(
        n14220) );
  AOI22_X1 U13596 ( .A1(n11093), .A2(n15288), .B1(n14966), .B2(n14220), .ZN(
        n15382) );
  NOR2_X1 U13597 ( .A1(n15382), .A2(n14550), .ZN(n11094) );
  AOI211_X1 U13598 ( .C1(n15282), .C2(n15380), .A(n11095), .B(n11094), .ZN(
        n11102) );
  OR2_X1 U13599 ( .A1(n11096), .A2(n11998), .ZN(n11097) );
  NAND2_X1 U13600 ( .A1(n15286), .A2(n11556), .ZN(n11098) );
  OR2_X1 U13601 ( .A1(n11100), .A2(n11099), .ZN(n15376) );
  NAND3_X1 U13602 ( .A1(n15376), .A2(n14654), .A3(n15374), .ZN(n11101) );
  OAI211_X1 U13603 ( .C1(n11103), .C2(n14982), .A(n11102), .B(n11101), .ZN(
        P1_U3283) );
  XNOR2_X1 U13604 ( .A(n11200), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n11108) );
  INV_X1 U13605 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n11105) );
  OAI21_X1 U13606 ( .B1(n11106), .B2(n11105), .A(n11104), .ZN(n11107) );
  NAND2_X1 U13607 ( .A1(n11108), .A2(n11107), .ZN(n11199) );
  OAI211_X1 U13608 ( .C1(n11108), .C2(n11107), .A(n15467), .B(n11199), .ZN(
        n11119) );
  NAND2_X1 U13609 ( .A1(P2_U3088), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n13520)
         );
  INV_X1 U13610 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n11113) );
  NAND2_X1 U13611 ( .A1(n11111), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n11196) );
  INV_X1 U13612 ( .A(n11196), .ZN(n11112) );
  AOI21_X1 U13613 ( .B1(n11113), .B2(n11200), .A(n11112), .ZN(n11114) );
  OAI211_X1 U13614 ( .C1(n11115), .C2(n11114), .A(n15474), .B(n11195), .ZN(
        n11116) );
  NAND2_X1 U13615 ( .A1(n13520), .A2(n11116), .ZN(n11117) );
  AOI21_X1 U13616 ( .B1(n15472), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n11117), 
        .ZN(n11118) );
  OAI211_X1 U13617 ( .C1(n15479), .C2(n11200), .A(n11119), .B(n11118), .ZN(
        P2_U3231) );
  XNOR2_X1 U13618 ( .A(n11120), .B(n12234), .ZN(n11374) );
  XNOR2_X1 U13619 ( .A(n11374), .B(n12631), .ZN(n11135) );
  XNOR2_X1 U13620 ( .A(n12234), .B(n15769), .ZN(n11128) );
  XNOR2_X1 U13621 ( .A(n11136), .B(n11128), .ZN(n11250) );
  OAI211_X1 U13622 ( .C1(n11125), .C2(n12634), .A(n11250), .B(n11121), .ZN(
        n11122) );
  NOR2_X1 U13623 ( .A1(n11248), .A2(n11122), .ZN(n11123) );
  NAND2_X1 U13624 ( .A1(n11124), .A2(n11123), .ZN(n11132) );
  INV_X1 U13625 ( .A(n11250), .ZN(n11127) );
  OAI21_X1 U13626 ( .B1(n11144), .B2(n11127), .A(n11248), .ZN(n11130) );
  NAND2_X1 U13627 ( .A1(n11125), .A2(n12634), .ZN(n11157) );
  INV_X1 U13628 ( .A(n11248), .ZN(n11126) );
  OAI21_X1 U13629 ( .B1(n11127), .B2(n11157), .A(n11126), .ZN(n11129) );
  AOI22_X1 U13630 ( .A1(n11130), .A2(n11129), .B1(n11128), .B2(n12632), .ZN(
        n11131) );
  INV_X1 U13631 ( .A(n15584), .ZN(n11133) );
  AOI21_X1 U13632 ( .B1(n11135), .B2(n11134), .A(n11133), .ZN(n11141) );
  OAI22_X1 U13633 ( .A1(n11136), .A2(n15019), .B1(n12498), .B2(n15017), .ZN(
        n11365) );
  OAI22_X1 U13634 ( .A1(n15581), .A2(n11403), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n13429), .ZN(n11139) );
  INV_X1 U13635 ( .A(n11137), .ZN(n11402) );
  NOR2_X1 U13636 ( .A1(n15593), .A2(n11402), .ZN(n11138) );
  AOI211_X1 U13637 ( .C1(n15591), .C2(n11365), .A(n11139), .B(n11138), .ZN(
        n11140) );
  OAI21_X1 U13638 ( .B1(n11141), .B2(n15585), .A(n11140), .ZN(P3_U3171) );
  XOR2_X1 U13639 ( .A(n11142), .B(n12483), .Z(n15764) );
  OAI21_X1 U13640 ( .B1(n6811), .B2(n7384), .A(n11143), .ZN(n11145) );
  INV_X1 U13641 ( .A(n12631), .ZN(n11376) );
  OAI22_X1 U13642 ( .A1(n11144), .A2(n15019), .B1(n11376), .B2(n15017), .ZN(
        n11257) );
  AOI21_X1 U13643 ( .B1(n11145), .B2(n15695), .A(n11257), .ZN(n15763) );
  MUX2_X1 U13644 ( .A(n11146), .B(n15763), .S(n15719), .Z(n11149) );
  INV_X1 U13645 ( .A(n11254), .ZN(n11147) );
  AOI22_X1 U13646 ( .A1(n15097), .A2(n15769), .B1(n11147), .B2(n12911), .ZN(
        n11148) );
  OAI211_X1 U13647 ( .C1(n12827), .C2(n15764), .A(n11149), .B(n11148), .ZN(
        P3_U3225) );
  INV_X1 U13648 ( .A(n15758), .ZN(n15761) );
  OAI22_X1 U13649 ( .A1(n12898), .A2(n12479), .B1(n11165), .B2(n15711), .ZN(
        n11155) );
  AOI22_X1 U13650 ( .A1(n12632), .A2(n12869), .B1(n12867), .B2(n12634), .ZN(
        n11160) );
  NAND2_X1 U13651 ( .A1(n11153), .A2(n11160), .ZN(n15755) );
  MUX2_X1 U13652 ( .A(P3_REG2_REG_7__SCAN_IN), .B(n15755), .S(n15719), .Z(
        n11154) );
  AOI211_X1 U13653 ( .C1(n15761), .C2(n15098), .A(n11155), .B(n11154), .ZN(
        n11156) );
  INV_X1 U13654 ( .A(n11156), .ZN(P3_U3226) );
  NAND2_X1 U13655 ( .A1(n11158), .A2(n11157), .ZN(n11249) );
  XNOR2_X1 U13656 ( .A(n11249), .B(n11248), .ZN(n11159) );
  NAND2_X1 U13657 ( .A1(n11159), .A2(n15021), .ZN(n11164) );
  NOR2_X1 U13658 ( .A1(n11160), .A2(n15009), .ZN(n11161) );
  AOI211_X1 U13659 ( .C1(n15756), .C2(n15012), .A(n11162), .B(n11161), .ZN(
        n11163) );
  OAI211_X1 U13660 ( .C1(n11165), .C2(n15593), .A(n11164), .B(n11163), .ZN(
        P3_U3153) );
  INV_X1 U13661 ( .A(n11166), .ZN(n11168) );
  OAI222_X1 U13662 ( .A1(n11169), .A2(P3_U3151), .B1(n14938), .B2(n11168), 
        .C1(n11167), .C2(n14936), .ZN(P3_U3271) );
  INV_X1 U13663 ( .A(n15140), .ZN(n15154) );
  XNOR2_X1 U13664 ( .A(n15140), .B(n13075), .ZN(n11170) );
  NAND2_X1 U13665 ( .A1(n13566), .A2(n11865), .ZN(n11171) );
  NAND2_X1 U13666 ( .A1(n11170), .A2(n11171), .ZN(n11189) );
  INV_X1 U13667 ( .A(n11170), .ZN(n11173) );
  INV_X1 U13668 ( .A(n11171), .ZN(n11172) );
  NAND2_X1 U13669 ( .A1(n11173), .A2(n11172), .ZN(n11174) );
  AND2_X1 U13670 ( .A1(n11189), .A2(n11174), .ZN(n11181) );
  INV_X1 U13671 ( .A(n11175), .ZN(n11176) );
  OAI21_X1 U13672 ( .B1(n11181), .B2(n11180), .A(n11190), .ZN(n11182) );
  NAND2_X1 U13673 ( .A1(n11182), .A2(n15123), .ZN(n11188) );
  NAND2_X1 U13674 ( .A1(n13567), .A2(n13701), .ZN(n11184) );
  NAND2_X1 U13675 ( .A1(n13565), .A2(n13555), .ZN(n11183) );
  AND2_X1 U13676 ( .A1(n11184), .A2(n11183), .ZN(n15134) );
  OAI21_X1 U13677 ( .B1(n13558), .B2(n15134), .A(n11185), .ZN(n11186) );
  AOI21_X1 U13678 ( .B1(n15138), .B2(n13556), .A(n11186), .ZN(n11187) );
  OAI211_X1 U13679 ( .C1(n15154), .C2(n13542), .A(n11188), .B(n11187), .ZN(
        P2_U3196) );
  XNOR2_X1 U13680 ( .A(n11491), .B(n13075), .ZN(n11868) );
  NAND2_X1 U13681 ( .A1(n13565), .A2(n11865), .ZN(n11869) );
  XNOR2_X1 U13682 ( .A(n11868), .B(n11869), .ZN(n11867) );
  XNOR2_X1 U13683 ( .A(n11866), .B(n11867), .ZN(n11194) );
  AOI22_X1 U13684 ( .A1(n13555), .A2(n13564), .B1(n13566), .B2(n13701), .ZN(
        n11428) );
  OAI22_X1 U13685 ( .A1(n13558), .A2(n11428), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n15451), .ZN(n11192) );
  INV_X1 U13686 ( .A(n11491), .ZN(n11490) );
  NOR2_X1 U13687 ( .A1(n11490), .A2(n13542), .ZN(n11191) );
  AOI211_X1 U13688 ( .C1(n13556), .C2(n11330), .A(n11192), .B(n11191), .ZN(
        n11193) );
  OAI21_X1 U13689 ( .B1(n11194), .B2(n13561), .A(n11193), .ZN(P2_U3206) );
  NOR2_X1 U13690 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n11197), .ZN(n13615) );
  AOI21_X1 U13691 ( .B1(P2_REG2_REG_18__SCAN_IN), .B2(n11197), .A(n13615), 
        .ZN(n11207) );
  INV_X1 U13692 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n11198) );
  NAND2_X1 U13693 ( .A1(P2_U3088), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n13547)
         );
  OAI21_X1 U13694 ( .B1(n15450), .B2(n11198), .A(n13547), .ZN(n11205) );
  INV_X1 U13695 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n11201) );
  OAI21_X1 U13696 ( .B1(n11201), .B2(n11200), .A(n11199), .ZN(n13617) );
  XOR2_X1 U13697 ( .A(n13618), .B(n13617), .Z(n11202) );
  NAND2_X1 U13698 ( .A1(P2_REG1_REG_18__SCAN_IN), .A2(n11202), .ZN(n13620) );
  OAI21_X1 U13699 ( .B1(P2_REG1_REG_18__SCAN_IN), .B2(n11202), .A(n13620), 
        .ZN(n11203) );
  NOR2_X1 U13700 ( .A1(n11203), .A2(n15459), .ZN(n11204) );
  AOI211_X1 U13701 ( .C1(n15453), .C2(n13618), .A(n11205), .B(n11204), .ZN(
        n11206) );
  OAI21_X1 U13702 ( .B1(n11207), .B2(n15442), .A(n11206), .ZN(P2_U3232) );
  NOR2_X1 U13703 ( .A1(n11614), .A2(n11208), .ZN(n11210) );
  NOR2_X1 U13704 ( .A1(n11210), .A2(n11209), .ZN(n11214) );
  INV_X1 U13705 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n11212) );
  NAND2_X1 U13706 ( .A1(n11621), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n14346) );
  INV_X1 U13707 ( .A(n14346), .ZN(n11211) );
  AOI21_X1 U13708 ( .B1(n11212), .B2(n14353), .A(n11211), .ZN(n11213) );
  NAND2_X1 U13709 ( .A1(n11213), .A2(n11214), .ZN(n14345) );
  OAI211_X1 U13710 ( .C1(n11214), .C2(n11213), .A(n14377), .B(n14345), .ZN(
        n11223) );
  NAND2_X1 U13711 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n14116)
         );
  NOR2_X1 U13712 ( .A1(n11614), .A2(n11215), .ZN(n11217) );
  XOR2_X1 U13713 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n11621), .Z(n11218) );
  OAI211_X1 U13714 ( .C1(n11219), .C2(n11218), .A(n14378), .B(n14352), .ZN(
        n11220) );
  NAND2_X1 U13715 ( .A1(n14116), .A2(n11220), .ZN(n11221) );
  AOI21_X1 U13716 ( .B1(n14360), .B2(P1_ADDR_REG_16__SCAN_IN), .A(n11221), 
        .ZN(n11222) );
  OAI211_X1 U13717 ( .C1(n15267), .C2(n14353), .A(n11223), .B(n11222), .ZN(
        P1_U3259) );
  OR2_X1 U13718 ( .A1(n11229), .A2(n13568), .ZN(n11224) );
  INV_X1 U13719 ( .A(n11320), .ZN(n11226) );
  AOI21_X1 U13720 ( .B1(n11325), .B2(n11227), .A(n11226), .ZN(n11396) );
  INV_X1 U13721 ( .A(n13568), .ZN(n11230) );
  OAI21_X1 U13722 ( .B1(n11230), .B2(n11229), .A(n11228), .ZN(n11231) );
  XNOR2_X1 U13723 ( .A(n11326), .B(n11325), .ZN(n11234) );
  INV_X1 U13724 ( .A(n11232), .ZN(n11233) );
  AOI21_X1 U13725 ( .B1(n11234), .B2(n15551), .A(n11233), .ZN(n11401) );
  NAND2_X1 U13726 ( .A1(n11235), .A2(n11395), .ZN(n11329) );
  INV_X1 U13727 ( .A(n11329), .ZN(n15145) );
  AOI211_X1 U13728 ( .C1(n11323), .C2(n11236), .A(n11865), .B(n15145), .ZN(
        n11399) );
  AOI21_X1 U13729 ( .B1(n15539), .B2(n11323), .A(n11399), .ZN(n11237) );
  OAI211_X1 U13730 ( .C1(n11396), .C2(n13998), .A(n11401), .B(n11237), .ZN(
        n11240) );
  NAND2_X1 U13731 ( .A1(n11240), .A2(n15576), .ZN(n11238) );
  OAI21_X1 U13732 ( .B1(n15158), .B2(n11239), .A(n11238), .ZN(P2_U3510) );
  INV_X1 U13733 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n11242) );
  NAND2_X1 U13734 ( .A1(n11240), .A2(n15561), .ZN(n11241) );
  OAI21_X1 U13735 ( .B1(n15561), .B2(n11242), .A(n11241), .ZN(P2_U3463) );
  INV_X1 U13736 ( .A(n11731), .ZN(n11247) );
  AOI21_X1 U13737 ( .B1(P2_DATAO_REG_23__SCAN_IN), .B2(n14797), .A(n11243), 
        .ZN(n11244) );
  OAI21_X1 U13738 ( .B1(n11247), .B2(n14815), .A(n11244), .ZN(P1_U3332) );
  AOI21_X1 U13739 ( .B1(P1_DATAO_REG_23__SCAN_IN), .B2(n14026), .A(n11245), 
        .ZN(n11246) );
  OAI21_X1 U13740 ( .B1(n11247), .B2(n14031), .A(n11246), .ZN(P2_U3304) );
  MUX2_X1 U13741 ( .A(n11249), .B(n12633), .S(n11248), .Z(n11251) );
  XNOR2_X1 U13742 ( .A(n11251), .B(n11250), .ZN(n11259) );
  OAI21_X1 U13743 ( .B1(n15581), .B2(n11253), .A(n11252), .ZN(n11256) );
  NOR2_X1 U13744 ( .A1(n15593), .A2(n11254), .ZN(n11255) );
  AOI211_X1 U13745 ( .C1(n15591), .C2(n11257), .A(n11256), .B(n11255), .ZN(
        n11258) );
  OAI21_X1 U13746 ( .B1(n11259), .B2(n15585), .A(n11258), .ZN(P3_U3161) );
  NOR2_X1 U13747 ( .A1(n11260), .A2(n15366), .ZN(n15348) );
  NAND2_X1 U13748 ( .A1(n15347), .A2(n14115), .ZN(n11261) );
  NAND2_X1 U13749 ( .A1(P1_U3086), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n14314) );
  OAI211_X1 U13750 ( .C1(n15176), .C2(n11262), .A(n11261), .B(n14314), .ZN(
        n11278) );
  NAND2_X1 U13751 ( .A1(n11995), .A2(n11832), .ZN(n11264) );
  NAND2_X1 U13752 ( .A1(n14223), .A2(n6664), .ZN(n11263) );
  NAND2_X1 U13753 ( .A1(n11264), .A2(n11263), .ZN(n11265) );
  XNOR2_X1 U13754 ( .A(n11265), .B(n11830), .ZN(n11353) );
  NAND2_X1 U13755 ( .A1(n11995), .A2(n6664), .ZN(n11267) );
  NAND2_X1 U13756 ( .A1(n14223), .A2(n10688), .ZN(n11266) );
  NAND2_X1 U13757 ( .A1(n11267), .A2(n11266), .ZN(n11352) );
  XNOR2_X1 U13758 ( .A(n11353), .B(n11352), .ZN(n11276) );
  NAND2_X1 U13759 ( .A1(n11271), .A2(n11270), .ZN(n11275) );
  INV_X1 U13760 ( .A(n11355), .ZN(n11274) );
  AOI211_X1 U13761 ( .C1(n11276), .C2(n11275), .A(n15167), .B(n11274), .ZN(
        n11277) );
  AOI211_X1 U13762 ( .C1(n14159), .C2(n15348), .A(n11278), .B(n11277), .ZN(
        n11279) );
  INV_X1 U13763 ( .A(n11279), .ZN(P1_U3213) );
  NAND2_X1 U13764 ( .A1(n15374), .A2(n11280), .ZN(n15179) );
  NAND2_X1 U13765 ( .A1(n11281), .A2(n11286), .ZN(n11284) );
  AOI22_X1 U13766 ( .A1(n12110), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n11657), 
        .B2(n11282), .ZN(n11283) );
  XNOR2_X1 U13767 ( .A(n15183), .B(n14220), .ZN(n15178) );
  NAND2_X1 U13768 ( .A1(n15179), .A2(n15178), .ZN(n15177) );
  INV_X1 U13769 ( .A(n14220), .ZN(n14093) );
  OR2_X1 U13770 ( .A1(n15183), .A2(n14093), .ZN(n11285) );
  NAND2_X1 U13771 ( .A1(n15177), .A2(n11285), .ZN(n11298) );
  NAND2_X1 U13772 ( .A1(n11287), .A2(n11286), .ZN(n11290) );
  AOI22_X1 U13773 ( .A1(n12110), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n11657), 
        .B2(n11288), .ZN(n11289) );
  NAND2_X1 U13774 ( .A1(n11837), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n11297) );
  AND2_X1 U13775 ( .A1(n11292), .A2(n11291), .ZN(n11293) );
  NOR2_X1 U13776 ( .A1(n11299), .A2(n11293), .ZN(n14095) );
  NAND2_X1 U13777 ( .A1(n11839), .A2(n14095), .ZN(n11296) );
  NAND2_X1 U13778 ( .A1(n11808), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n11295) );
  NAND2_X1 U13779 ( .A1(n12113), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n11294) );
  NAND4_X1 U13780 ( .A1(n11297), .A2(n11296), .A3(n11295), .A4(n11294), .ZN(
        n14219) );
  XNOR2_X1 U13781 ( .A(n14955), .B(n14219), .ZN(n12159) );
  NAND2_X1 U13782 ( .A1(n11298), .A2(n12159), .ZN(n11444) );
  OAI211_X1 U13783 ( .C1(n11298), .C2(n12159), .A(n11444), .B(n15375), .ZN(
        n11307) );
  NAND2_X1 U13784 ( .A1(n11299), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n11455) );
  OR2_X1 U13785 ( .A1(n11299), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n11300) );
  NAND2_X1 U13786 ( .A1(n11455), .A2(n11300), .ZN(n14987) );
  INV_X1 U13787 ( .A(n14987), .ZN(n11301) );
  NAND2_X1 U13788 ( .A1(n11839), .A2(n11301), .ZN(n11305) );
  NAND2_X1 U13789 ( .A1(n11837), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n11304) );
  NAND2_X1 U13790 ( .A1(n12113), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n11303) );
  NAND2_X1 U13791 ( .A1(n11808), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n11302) );
  NAND4_X1 U13792 ( .A1(n11305), .A2(n11304), .A3(n11303), .A4(n11302), .ZN(
        n14218) );
  AOI22_X1 U13793 ( .A1(n14966), .A2(n14218), .B1(n14220), .B2(n15378), .ZN(
        n11306) );
  AND2_X1 U13794 ( .A1(n11307), .A2(n11306), .ZN(n14962) );
  XNOR2_X1 U13795 ( .A(n15187), .B(n14955), .ZN(n11308) );
  NAND2_X1 U13796 ( .A1(n11308), .A2(n15288), .ZN(n14957) );
  INV_X1 U13797 ( .A(n14957), .ZN(n11311) );
  INV_X1 U13798 ( .A(n14955), .ZN(n14098) );
  AOI22_X1 U13799 ( .A1(n6665), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n14095), 
        .B2(n15293), .ZN(n11309) );
  OAI21_X1 U13800 ( .B1(n14098), .B2(n15297), .A(n11309), .ZN(n11310) );
  AOI21_X1 U13801 ( .B1(n11311), .B2(n15299), .A(n11310), .ZN(n11318) );
  NAND2_X1 U13802 ( .A1(n11312), .A2(n12158), .ZN(n11314) );
  OR2_X1 U13803 ( .A1(n15380), .A2(n14221), .ZN(n11313) );
  NAND2_X1 U13804 ( .A1(n11314), .A2(n11313), .ZN(n15185) );
  INV_X1 U13805 ( .A(n15178), .ZN(n15184) );
  NAND2_X1 U13806 ( .A1(n15185), .A2(n15184), .ZN(n11316) );
  OR2_X1 U13807 ( .A1(n15183), .A2(n14220), .ZN(n11315) );
  NAND2_X1 U13808 ( .A1(n11316), .A2(n11315), .ZN(n11476) );
  INV_X1 U13809 ( .A(n12159), .ZN(n11475) );
  XNOR2_X1 U13810 ( .A(n11476), .B(n11475), .ZN(n14958) );
  NAND2_X1 U13811 ( .A1(n14958), .A2(n15191), .ZN(n11317) );
  OAI211_X1 U13812 ( .C1(n14962), .C2(n6665), .A(n11318), .B(n11317), .ZN(
        P1_U3281) );
  OR2_X1 U13813 ( .A1(n11323), .A2(n13567), .ZN(n11319) );
  NAND2_X1 U13814 ( .A1(n11320), .A2(n11319), .ZN(n15142) );
  NAND2_X1 U13815 ( .A1(n15140), .A2(n13566), .ZN(n11321) );
  OR2_X1 U13816 ( .A1(n15140), .A2(n13566), .ZN(n11322) );
  XOR2_X1 U13817 ( .A(n11328), .B(n11487), .Z(n11433) );
  XNOR2_X1 U13818 ( .A(n11489), .B(n11328), .ZN(n11431) );
  OR2_X2 U13819 ( .A1(n11329), .A2(n15140), .ZN(n15143) );
  AOI211_X1 U13820 ( .C1(n11491), .C2(n15143), .A(n11865), .B(n11499), .ZN(
        n11430) );
  NAND2_X1 U13821 ( .A1(n11430), .A2(n15147), .ZN(n11334) );
  INV_X1 U13822 ( .A(n11330), .ZN(n11331) );
  OAI22_X1 U13823 ( .A1(n15151), .A2(n11428), .B1(n11331), .B2(n13865), .ZN(
        n11332) );
  AOI21_X1 U13824 ( .B1(P2_REG2_REG_13__SCAN_IN), .B2(n15151), .A(n11332), 
        .ZN(n11333) );
  OAI211_X1 U13825 ( .C1(n11490), .C2(n13890), .A(n11334), .B(n11333), .ZN(
        n11335) );
  AOI21_X1 U13826 ( .B1(n11431), .B2(n13872), .A(n11335), .ZN(n11336) );
  OAI21_X1 U13827 ( .B1(n13874), .B2(n11433), .A(n11336), .ZN(P2_U3252) );
  OAI211_X1 U13828 ( .C1(n11341), .C2(n11337), .A(n11411), .B(n15695), .ZN(
        n11340) );
  NAND2_X1 U13829 ( .A1(n12631), .A2(n12867), .ZN(n11339) );
  NAND2_X1 U13830 ( .A1(n12629), .A2(n12869), .ZN(n11338) );
  AND2_X1 U13831 ( .A1(n11339), .A2(n11338), .ZN(n15578) );
  NAND2_X1 U13832 ( .A1(n11340), .A2(n15578), .ZN(n11439) );
  INV_X1 U13833 ( .A(n11439), .ZN(n11347) );
  XNOR2_X1 U13834 ( .A(n11342), .B(n11341), .ZN(n11440) );
  NOR2_X1 U13835 ( .A1(n15719), .A2(n11343), .ZN(n11345) );
  OAI22_X1 U13836 ( .A1(n12898), .A2(n15580), .B1(n15594), .B2(n15711), .ZN(
        n11344) );
  AOI211_X1 U13837 ( .C1(n11440), .C2(n15098), .A(n11345), .B(n11344), .ZN(
        n11346) );
  OAI21_X1 U13838 ( .B1(n11347), .B2(n15703), .A(n11346), .ZN(P3_U3223) );
  NAND2_X1 U13839 ( .A1(n11998), .A2(n11832), .ZN(n11349) );
  NAND2_X1 U13840 ( .A1(n14222), .A2(n6664), .ZN(n11348) );
  NAND2_X1 U13841 ( .A1(n11349), .A2(n11348), .ZN(n11350) );
  XNOR2_X1 U13842 ( .A(n11350), .B(n11830), .ZN(n11516) );
  AND2_X1 U13843 ( .A1(n14222), .A2(n10688), .ZN(n11351) );
  AOI21_X1 U13844 ( .B1(n11998), .B2(n6664), .A(n11351), .ZN(n11517) );
  XNOR2_X1 U13845 ( .A(n11516), .B(n11517), .ZN(n11357) );
  NAND2_X1 U13846 ( .A1(n11353), .A2(n11352), .ZN(n11354) );
  OAI21_X1 U13847 ( .B1(n11357), .B2(n11356), .A(n11519), .ZN(n11358) );
  NAND2_X1 U13848 ( .A1(n11358), .A2(n14195), .ZN(n11362) );
  INV_X1 U13849 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n11359) );
  OAI22_X1 U13850 ( .A1(n15356), .A2(n14200), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n11359), .ZN(n11360) );
  AOI21_X1 U13851 ( .B1(n7912), .B2(n14208), .A(n11360), .ZN(n11361) );
  OAI211_X1 U13852 ( .C1(n15358), .C2(n14191), .A(n11362), .B(n11361), .ZN(
        P1_U3221) );
  XOR2_X1 U13853 ( .A(n11363), .B(n12489), .Z(n11404) );
  AOI21_X1 U13854 ( .B1(n11364), .B2(n12489), .A(n15708), .ZN(n11367) );
  AOI21_X1 U13855 ( .B1(n11367), .B2(n11366), .A(n11365), .ZN(n11408) );
  OAI21_X1 U13856 ( .B1(n11404), .B2(n15106), .A(n11408), .ZN(n11372) );
  INV_X1 U13857 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n13408) );
  OAI22_X1 U13858 ( .A1(n13049), .A2(n11403), .B1(n15773), .B2(n13408), .ZN(
        n11368) );
  AOI21_X1 U13859 ( .B1(n11372), .B2(n15773), .A(n11368), .ZN(n11369) );
  INV_X1 U13860 ( .A(n11369), .ZN(P3_U3417) );
  OAI22_X1 U13861 ( .A1(n12986), .A2(n11403), .B1(n15788), .B2(n11370), .ZN(
        n11371) );
  AOI21_X1 U13862 ( .B1(n11372), .B2(n15788), .A(n11371), .ZN(n11373) );
  INV_X1 U13863 ( .A(n11373), .ZN(P3_U3468) );
  XNOR2_X1 U13864 ( .A(n15580), .B(n12270), .ZN(n11378) );
  XNOR2_X1 U13865 ( .A(n12498), .B(n11378), .ZN(n15582) );
  INV_X1 U13866 ( .A(n11374), .ZN(n11375) );
  NAND2_X1 U13867 ( .A1(n11376), .A2(n11375), .ZN(n15583) );
  AND2_X1 U13868 ( .A1(n15582), .A2(n15583), .ZN(n11377) );
  NAND2_X1 U13869 ( .A1(n12630), .A2(n11378), .ZN(n11382) );
  XNOR2_X1 U13870 ( .A(n13048), .B(n12270), .ZN(n11380) );
  INV_X1 U13871 ( .A(n11380), .ZN(n11381) );
  AND2_X1 U13872 ( .A1(n11382), .A2(n11381), .ZN(n11383) );
  NAND2_X1 U13873 ( .A1(n11379), .A2(n11383), .ZN(n12288) );
  NAND2_X1 U13874 ( .A1(n12194), .A2(n12288), .ZN(n11384) );
  INV_X1 U13875 ( .A(n12629), .ZN(n12193) );
  XNOR2_X1 U13876 ( .A(n11384), .B(n12193), .ZN(n11388) );
  NOR2_X1 U13877 ( .A1(n15581), .A2(n13048), .ZN(n11386) );
  AOI22_X1 U13878 ( .A1(n12630), .A2(n12867), .B1(n12869), .B2(n12628), .ZN(
        n11413) );
  INV_X1 U13879 ( .A(P3_REG3_REG_11__SCAN_IN), .ZN(n15619) );
  OAI22_X1 U13880 ( .A1(n11413), .A2(n15009), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n15619), .ZN(n11385) );
  AOI211_X1 U13881 ( .C1(n15002), .C2(n11417), .A(n11386), .B(n11385), .ZN(
        n11387) );
  OAI21_X1 U13882 ( .B1(n11388), .B2(n15585), .A(n11387), .ZN(P3_U3176) );
  INV_X1 U13883 ( .A(n11389), .ZN(n11390) );
  OAI222_X1 U13884 ( .A1(P3_U3151), .A2(n11392), .B1(n14936), .B2(n11391), 
        .C1(n14938), .C2(n11390), .ZN(P3_U3270) );
  AOI22_X1 U13885 ( .A1(n15151), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n11393), 
        .B2(n15137), .ZN(n11394) );
  OAI21_X1 U13886 ( .B1(n11395), .B2(n13890), .A(n11394), .ZN(n11398) );
  NOR2_X1 U13887 ( .A1(n11396), .A2(n13874), .ZN(n11397) );
  AOI211_X1 U13888 ( .C1(n11399), .C2(n15147), .A(n11398), .B(n11397), .ZN(
        n11400) );
  OAI21_X1 U13889 ( .B1(n15151), .B2(n11401), .A(n11400), .ZN(P2_U3254) );
  OAI22_X1 U13890 ( .A1(n12898), .A2(n11403), .B1(n11402), .B2(n15711), .ZN(
        n11406) );
  NOR2_X1 U13891 ( .A1(n11404), .A2(n12827), .ZN(n11405) );
  AOI211_X1 U13892 ( .C1(n15703), .C2(P3_REG2_REG_9__SCAN_IN), .A(n11406), .B(
        n11405), .ZN(n11407) );
  OAI21_X1 U13893 ( .B1(n15703), .B2(n11408), .A(n11407), .ZN(P3_U3224) );
  NAND3_X1 U13894 ( .A1(n11411), .A2(n8172), .A3(n11410), .ZN(n11412) );
  NAND3_X1 U13895 ( .A1(n11409), .A2(n15695), .A3(n11412), .ZN(n11414) );
  NAND2_X1 U13896 ( .A1(n11414), .A2(n11413), .ZN(n12982) );
  INV_X1 U13897 ( .A(n12982), .ZN(n11423) );
  OAI21_X1 U13898 ( .B1(n11416), .B2(n8172), .A(n11415), .ZN(n12983) );
  INV_X1 U13899 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n11420) );
  AOI22_X1 U13900 ( .A1(n15097), .A2(n11418), .B1(n12911), .B2(n11417), .ZN(
        n11419) );
  OAI21_X1 U13901 ( .B1(n11420), .B2(n15719), .A(n11419), .ZN(n11421) );
  AOI21_X1 U13902 ( .B1(n12983), .B2(n15098), .A(n11421), .ZN(n11422) );
  OAI21_X1 U13903 ( .B1(n11423), .B2(n15703), .A(n11422), .ZN(P3_U3222) );
  INV_X1 U13904 ( .A(n11424), .ZN(n11426) );
  OAI222_X1 U13905 ( .A1(n11427), .A2(P3_U3151), .B1(n14938), .B2(n11426), 
        .C1(n11425), .C2(n14936), .ZN(P3_U3269) );
  OAI21_X1 U13906 ( .B1(n11490), .B2(n15548), .A(n11428), .ZN(n11429) );
  AOI211_X1 U13907 ( .C1(n11431), .C2(n15551), .A(n11430), .B(n11429), .ZN(
        n11432) );
  OAI21_X1 U13908 ( .B1(n13998), .B2(n11433), .A(n11432), .ZN(n11436) );
  NAND2_X1 U13909 ( .A1(n11436), .A2(n15576), .ZN(n11434) );
  OAI21_X1 U13910 ( .B1(n15576), .B2(n11435), .A(n11434), .ZN(P2_U3512) );
  INV_X1 U13911 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n11438) );
  NAND2_X1 U13912 ( .A1(n11436), .A2(n15561), .ZN(n11437) );
  OAI21_X1 U13913 ( .B1(n15561), .B2(n11438), .A(n11437), .ZN(P2_U3469) );
  INV_X1 U13914 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n11441) );
  AOI21_X1 U13915 ( .B1(n11440), .B2(n15746), .A(n11439), .ZN(n11484) );
  MUX2_X1 U13916 ( .A(n11441), .B(n11484), .S(n15773), .Z(n11442) );
  OAI21_X1 U13917 ( .B1(n13049), .B2(n15580), .A(n11442), .ZN(P3_U3420) );
  INV_X1 U13918 ( .A(n14219), .ZN(n15213) );
  OR2_X1 U13919 ( .A1(n14955), .A2(n15213), .ZN(n11443) );
  NAND2_X1 U13920 ( .A1(n11444), .A2(n11443), .ZN(n14973) );
  NAND2_X1 U13921 ( .A1(n11445), .A2(n11286), .ZN(n11448) );
  AOI22_X1 U13922 ( .A1(n12110), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n11446), 
        .B2(n11657), .ZN(n11447) );
  XNOR2_X1 U13923 ( .A(n15216), .B(n14218), .ZN(n14972) );
  NAND2_X1 U13924 ( .A1(n14973), .A2(n14972), .ZN(n14971) );
  INV_X1 U13925 ( .A(n14218), .ZN(n15162) );
  OR2_X1 U13926 ( .A1(n15216), .A2(n15162), .ZN(n11449) );
  NAND2_X1 U13927 ( .A1(n11450), .A2(n11286), .ZN(n11453) );
  AOI22_X1 U13928 ( .A1(n11451), .A2(n11657), .B1(n12110), .B2(
        P2_DATAO_REG_14__SCAN_IN), .ZN(n11452) );
  INV_X1 U13929 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n11454) );
  NAND2_X1 U13930 ( .A1(n11455), .A2(n11454), .ZN(n11456) );
  NAND2_X1 U13931 ( .A1(n11464), .A2(n11456), .ZN(n15175) );
  INV_X1 U13932 ( .A(n15175), .ZN(n11470) );
  NAND2_X1 U13933 ( .A1(n11839), .A2(n11470), .ZN(n11460) );
  NAND2_X1 U13934 ( .A1(n11837), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n11459) );
  NAND2_X1 U13935 ( .A1(n12113), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n11458) );
  NAND2_X1 U13936 ( .A1(n11808), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n11457) );
  NAND4_X1 U13937 ( .A1(n11460), .A2(n11459), .A3(n11458), .A4(n11457), .ZN(
        n14967) );
  INV_X1 U13938 ( .A(n14967), .ZN(n14211) );
  NAND2_X1 U13939 ( .A1(n15203), .A2(n14211), .ZN(n12025) );
  OAI21_X1 U13940 ( .B1(n11461), .B2(n12147), .A(n14661), .ZN(n15208) );
  NOR2_X1 U13942 ( .A1(n14975), .A2(n15203), .ZN(n14668) );
  NAND2_X1 U13943 ( .A1(n14975), .A2(n15203), .ZN(n11462) );
  NAND2_X1 U13944 ( .A1(n11462), .A2(n15288), .ZN(n11463) );
  NOR2_X1 U13945 ( .A1(n14668), .A2(n11463), .ZN(n15201) );
  NAND2_X1 U13946 ( .A1(n12112), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n11469) );
  AND2_X1 U13947 ( .A1(n11464), .A2(n13404), .ZN(n11465) );
  NOR2_X1 U13948 ( .A1(n11624), .A2(n11465), .ZN(n14671) );
  NAND2_X1 U13949 ( .A1(n11839), .A2(n14671), .ZN(n11468) );
  NAND2_X1 U13950 ( .A1(n11808), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n11467) );
  NAND2_X1 U13951 ( .A1(n12113), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n11466) );
  NAND4_X1 U13952 ( .A1(n11469), .A2(n11468), .A3(n11467), .A4(n11466), .ZN(
        n14421) );
  INV_X1 U13953 ( .A(n14421), .ZN(n15163) );
  OAI22_X1 U13954 ( .A1(n15163), .A2(n14607), .B1(n15162), .B2(n15212), .ZN(
        n15202) );
  AOI21_X1 U13955 ( .B1(n11470), .B2(n15293), .A(n15202), .ZN(n11473) );
  NAND2_X1 U13956 ( .A1(n15203), .A2(n15282), .ZN(n11472) );
  NAND2_X1 U13957 ( .A1(n6665), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n11471) );
  OAI211_X1 U13958 ( .C1(n6665), .C2(n11473), .A(n11472), .B(n11471), .ZN(
        n11474) );
  AOI21_X1 U13959 ( .B1(n15201), .B2(n15299), .A(n11474), .ZN(n11483) );
  NAND2_X1 U13960 ( .A1(n11476), .A2(n11475), .ZN(n11478) );
  OR2_X1 U13961 ( .A1(n14955), .A2(n14219), .ZN(n11477) );
  INV_X1 U13962 ( .A(n14972), .ZN(n12162) );
  OR2_X1 U13963 ( .A1(n15216), .A2(n14218), .ZN(n11479) );
  NAND2_X1 U13964 ( .A1(n11481), .A2(n12147), .ZN(n15204) );
  NAND3_X1 U13965 ( .A1(n15205), .A2(n15204), .A3(n15191), .ZN(n11482) );
  OAI211_X1 U13966 ( .C1(n15208), .C2(n14599), .A(n11483), .B(n11482), .ZN(
        P1_U3279) );
  MUX2_X1 U13967 ( .A(n8143), .B(n11484), .S(n15788), .Z(n11485) );
  OAI21_X1 U13968 ( .B1(n12986), .B2(n15580), .A(n11485), .ZN(P3_U3469) );
  NOR2_X1 U13969 ( .A1(n11491), .A2(n13565), .ZN(n11486) );
  NAND2_X1 U13970 ( .A1(n11491), .A2(n13565), .ZN(n11488) );
  XNOR2_X1 U13971 ( .A(n11527), .B(n11492), .ZN(n13997) );
  INV_X1 U13972 ( .A(n11492), .ZN(n11493) );
  OAI211_X1 U13973 ( .C1(n11494), .C2(n11493), .A(n11529), .B(n15551), .ZN(
        n11497) );
  OAI22_X1 U13974 ( .A1(n13667), .A2(n13630), .B1(n11495), .B2(n13496), .ZN(
        n15126) );
  INV_X1 U13975 ( .A(n15126), .ZN(n11496) );
  NAND2_X1 U13976 ( .A1(n11497), .A2(n11496), .ZN(n13994) );
  INV_X1 U13977 ( .A(n15127), .ZN(n11498) );
  OAI21_X1 U13978 ( .B1(n11499), .B2(n11498), .A(n15144), .ZN(n11500) );
  AND2_X2 U13979 ( .A1(n11499), .A2(n11498), .ZN(n11532) );
  NOR2_X1 U13980 ( .A1(n11500), .A2(n11532), .ZN(n13995) );
  NAND2_X1 U13981 ( .A1(n13995), .A2(n15147), .ZN(n11504) );
  NAND2_X1 U13982 ( .A1(n15151), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n11501) );
  OAI21_X1 U13983 ( .B1(n13865), .B2(n15132), .A(n11501), .ZN(n11502) );
  AOI21_X1 U13984 ( .B1(n15127), .B2(n15139), .A(n11502), .ZN(n11503) );
  NAND2_X1 U13985 ( .A1(n11504), .A2(n11503), .ZN(n11505) );
  AOI21_X1 U13986 ( .B1(n13994), .B2(n13852), .A(n11505), .ZN(n11506) );
  OAI21_X1 U13987 ( .B1(n13874), .B2(n13997), .A(n11506), .ZN(P2_U3251) );
  INV_X1 U13988 ( .A(n11507), .ZN(n11508) );
  OAI222_X1 U13989 ( .A1(n14938), .A2(n11508), .B1(n14936), .B2(n13471), .C1(
        P3_U3151), .C2(n12696), .ZN(P3_U3268) );
  INV_X1 U13990 ( .A(n11750), .ZN(n11512) );
  OAI222_X1 U13991 ( .A1(n14817), .A2(n11510), .B1(n14815), .B2(n11512), .C1(
        n11509), .C2(P1_U3086), .ZN(P1_U3331) );
  OAI222_X1 U13992 ( .A1(n14038), .A2(n6982), .B1(n14031), .B2(n11512), .C1(
        P2_U3088), .C2(n11511), .ZN(P2_U3303) );
  NAND2_X1 U13993 ( .A1(n15286), .A2(n11832), .ZN(n11514) );
  NAND2_X1 U13994 ( .A1(n15377), .A2(n6664), .ZN(n11513) );
  NAND2_X1 U13995 ( .A1(n11514), .A2(n11513), .ZN(n11515) );
  XNOR2_X1 U13996 ( .A(n11515), .B(n11778), .ZN(n11540) );
  INV_X1 U13997 ( .A(n11516), .ZN(n11518) );
  NAND2_X1 U13998 ( .A1(n15286), .A2(n6664), .ZN(n11521) );
  NAND2_X1 U13999 ( .A1(n15377), .A2(n10688), .ZN(n11520) );
  NAND2_X1 U14000 ( .A1(n11521), .A2(n11520), .ZN(n11542) );
  XOR2_X1 U14001 ( .A(n11540), .B(n11541), .Z(n11525) );
  AOI22_X1 U14002 ( .A1(n14966), .A2(n14221), .B1(n14222), .B2(n15378), .ZN(
        n15275) );
  INV_X1 U14003 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n14332) );
  OAI22_X1 U14004 ( .A1(n15275), .A2(n14200), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14332), .ZN(n11522) );
  AOI21_X1 U14005 ( .B1(n15281), .B2(n14208), .A(n11522), .ZN(n11524) );
  NAND2_X1 U14006 ( .A1(n15286), .A2(n15172), .ZN(n11523) );
  OAI211_X1 U14007 ( .C1(n11525), .C2(n15167), .A(n11524), .B(n11523), .ZN(
        P1_U3231) );
  AND2_X1 U14008 ( .A1(n15127), .A2(n13564), .ZN(n11526) );
  XNOR2_X1 U14009 ( .A(n13642), .B(n7216), .ZN(n13993) );
  OAI211_X1 U14010 ( .C1(n11530), .C2(n7216), .A(n13669), .B(n15551), .ZN(
        n11531) );
  AOI22_X1 U14011 ( .A1(n13555), .A2(n13670), .B1(n13564), .B2(n13701), .ZN(
        n11927) );
  NAND2_X1 U14012 ( .A1(n11531), .A2(n11927), .ZN(n13989) );
  INV_X1 U14013 ( .A(n13991), .ZN(n11537) );
  INV_X1 U14014 ( .A(n11532), .ZN(n11534) );
  NAND2_X1 U14015 ( .A1(n11532), .A2(n11537), .ZN(n13884) );
  INV_X1 U14016 ( .A(n13884), .ZN(n11533) );
  AOI211_X1 U14017 ( .C1(n13991), .C2(n11534), .A(n11865), .B(n11533), .ZN(
        n13990) );
  NAND2_X1 U14018 ( .A1(n13990), .A2(n15147), .ZN(n11536) );
  AOI22_X1 U14019 ( .A1(n15151), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n11925), 
        .B2(n15137), .ZN(n11535) );
  OAI211_X1 U14020 ( .C1(n11537), .C2(n13890), .A(n11536), .B(n11535), .ZN(
        n11538) );
  AOI21_X1 U14021 ( .B1(n13989), .B2(n13852), .A(n11538), .ZN(n11539) );
  OAI21_X1 U14022 ( .B1(n13874), .B2(n13993), .A(n11539), .ZN(P2_U3250) );
  INV_X1 U14023 ( .A(n11542), .ZN(n11543) );
  NAND2_X1 U14024 ( .A1(n11544), .A2(n11543), .ZN(n11545) );
  NAND2_X1 U14025 ( .A1(n15380), .A2(n11832), .ZN(n11548) );
  NAND2_X1 U14026 ( .A1(n14221), .A2(n6664), .ZN(n11547) );
  NAND2_X1 U14027 ( .A1(n11548), .A2(n11547), .ZN(n11549) );
  XNOR2_X1 U14028 ( .A(n11549), .B(n11778), .ZN(n11573) );
  AND2_X1 U14029 ( .A1(n14221), .A2(n10688), .ZN(n11550) );
  AOI21_X1 U14030 ( .B1(n15380), .B2(n6664), .A(n11550), .ZN(n11574) );
  XNOR2_X1 U14031 ( .A(n11573), .B(n11574), .ZN(n11551) );
  XNOR2_X1 U14032 ( .A(n11572), .B(n11551), .ZN(n11559) );
  AOI21_X1 U14033 ( .B1(n14207), .B2(n14220), .A(n11552), .ZN(n11555) );
  NAND2_X1 U14034 ( .A1(n14208), .A2(n11553), .ZN(n11554) );
  OAI211_X1 U14035 ( .C1(n11556), .C2(n15161), .A(n11555), .B(n11554), .ZN(
        n11557) );
  AOI21_X1 U14036 ( .B1(n15380), .B2(n15172), .A(n11557), .ZN(n11558) );
  OAI21_X1 U14037 ( .B1(n11559), .B2(n15167), .A(n11558), .ZN(P1_U3217) );
  INV_X1 U14038 ( .A(n11804), .ZN(n14030) );
  OAI222_X1 U14039 ( .A1(n14817), .A2(n11560), .B1(n14815), .B2(n14030), .C1(
        n6668), .C2(P1_U3086), .ZN(P1_U3328) );
  NAND2_X1 U14040 ( .A1(n11561), .A2(n11286), .ZN(n11563) );
  AOI22_X1 U14041 ( .A1(n12110), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n11657), 
        .B2(n14372), .ZN(n11562) );
  NAND2_X1 U14042 ( .A1(n12112), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n11567) );
  XNOR2_X1 U14043 ( .A(n11663), .B(P1_REG3_REG_18__SCAN_IN), .ZN(n14618) );
  NAND2_X1 U14044 ( .A1(n11839), .A2(n14618), .ZN(n11566) );
  NAND2_X1 U14045 ( .A1(n11808), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n11565) );
  NAND2_X1 U14046 ( .A1(n12113), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n11564) );
  NAND4_X1 U14047 ( .A1(n11567), .A2(n11566), .A3(n11565), .A4(n11564), .ZN(
        n14217) );
  AND2_X1 U14048 ( .A1(n14217), .A2(n10688), .ZN(n11568) );
  AOI21_X1 U14049 ( .B1(n14762), .B2(n6664), .A(n11568), .ZN(n11688) );
  NAND2_X1 U14050 ( .A1(n14762), .A2(n11832), .ZN(n11570) );
  NAND2_X1 U14051 ( .A1(n14217), .A2(n6664), .ZN(n11569) );
  NAND2_X1 U14052 ( .A1(n11570), .A2(n11569), .ZN(n11571) );
  XNOR2_X1 U14053 ( .A(n11571), .B(n11778), .ZN(n14069) );
  INV_X1 U14054 ( .A(n11573), .ZN(n11576) );
  INV_X1 U14055 ( .A(n11574), .ZN(n11575) );
  NAND2_X1 U14056 ( .A1(n11576), .A2(n11575), .ZN(n11577) );
  NAND2_X1 U14057 ( .A1(n15183), .A2(n11832), .ZN(n11579) );
  NAND2_X1 U14058 ( .A1(n14220), .A2(n6664), .ZN(n11578) );
  NAND2_X1 U14059 ( .A1(n11579), .A2(n11578), .ZN(n11580) );
  XNOR2_X1 U14060 ( .A(n11580), .B(n11830), .ZN(n11586) );
  AND2_X1 U14061 ( .A1(n14220), .A2(n10688), .ZN(n11581) );
  AOI21_X1 U14062 ( .B1(n15183), .B2(n6664), .A(n11581), .ZN(n11587) );
  XNOR2_X1 U14063 ( .A(n11586), .B(n11587), .ZN(n14174) );
  NAND2_X1 U14064 ( .A1(n14955), .A2(n11832), .ZN(n11583) );
  NAND2_X1 U14065 ( .A1(n14219), .A2(n6664), .ZN(n11582) );
  NAND2_X1 U14066 ( .A1(n11583), .A2(n11582), .ZN(n11584) );
  XNOR2_X1 U14067 ( .A(n11584), .B(n11830), .ZN(n11592) );
  AND2_X1 U14068 ( .A1(n14219), .A2(n10688), .ZN(n11585) );
  AOI21_X1 U14069 ( .B1(n14955), .B2(n6664), .A(n11585), .ZN(n11590) );
  XNOR2_X1 U14070 ( .A(n11592), .B(n11590), .ZN(n14089) );
  INV_X1 U14071 ( .A(n11586), .ZN(n11588) );
  NAND2_X1 U14072 ( .A1(n11588), .A2(n11587), .ZN(n14087) );
  AND2_X1 U14073 ( .A1(n14089), .A2(n14087), .ZN(n11589) );
  NAND2_X1 U14074 ( .A1(n14172), .A2(n11589), .ZN(n14088) );
  INV_X1 U14075 ( .A(n11590), .ZN(n11591) );
  NAND2_X1 U14076 ( .A1(n11592), .A2(n11591), .ZN(n11593) );
  NAND2_X1 U14077 ( .A1(n14088), .A2(n11593), .ZN(n14152) );
  NAND2_X1 U14078 ( .A1(n15216), .A2(n11832), .ZN(n11595) );
  NAND2_X1 U14079 ( .A1(n14218), .A2(n6664), .ZN(n11594) );
  NAND2_X1 U14080 ( .A1(n11595), .A2(n11594), .ZN(n11596) );
  XNOR2_X1 U14081 ( .A(n11596), .B(n11830), .ZN(n11600) );
  AND2_X1 U14082 ( .A1(n14218), .A2(n10688), .ZN(n11597) );
  AOI21_X1 U14083 ( .B1(n15216), .B2(n6664), .A(n11597), .ZN(n11598) );
  XNOR2_X1 U14084 ( .A(n11600), .B(n11598), .ZN(n14151) );
  INV_X1 U14085 ( .A(n11598), .ZN(n11599) );
  NAND2_X1 U14086 ( .A1(n11600), .A2(n11599), .ZN(n11601) );
  NAND2_X1 U14087 ( .A1(n15203), .A2(n11832), .ZN(n11603) );
  NAND2_X1 U14088 ( .A1(n14967), .A2(n6664), .ZN(n11602) );
  NAND2_X1 U14089 ( .A1(n11603), .A2(n11602), .ZN(n11604) );
  XNOR2_X1 U14090 ( .A(n11604), .B(n11778), .ZN(n11606) );
  AND2_X1 U14091 ( .A1(n14967), .A2(n10688), .ZN(n11605) );
  AOI21_X1 U14092 ( .B1(n15203), .B2(n6664), .A(n11605), .ZN(n11607) );
  NAND2_X1 U14093 ( .A1(n11606), .A2(n11607), .ZN(n11612) );
  INV_X1 U14094 ( .A(n11606), .ZN(n11609) );
  INV_X1 U14095 ( .A(n11607), .ZN(n11608) );
  NAND2_X1 U14096 ( .A1(n11609), .A2(n11608), .ZN(n11610) );
  NAND2_X1 U14097 ( .A1(n11612), .A2(n11610), .ZN(n15166) );
  INV_X1 U14098 ( .A(n15166), .ZN(n11611) );
  NAND2_X1 U14099 ( .A1(n11613), .A2(n11286), .ZN(n11616) );
  AOI22_X1 U14100 ( .A1(n12110), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n11657), 
        .B2(n11614), .ZN(n11615) );
  AOI22_X1 U14101 ( .A1(n14672), .A2(n11832), .B1(n6664), .B2(n14421), .ZN(
        n11617) );
  XNOR2_X1 U14102 ( .A(n11617), .B(n11830), .ZN(n11619) );
  AOI22_X1 U14103 ( .A1(n14672), .A2(n6664), .B1(n10688), .B2(n14421), .ZN(
        n14205) );
  NAND2_X1 U14104 ( .A1(n11620), .A2(n11286), .ZN(n11623) );
  AOI22_X1 U14105 ( .A1(n12110), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n11657), 
        .B2(n11621), .ZN(n11622) );
  NAND2_X1 U14106 ( .A1(n14773), .A2(n11832), .ZN(n11631) );
  NAND2_X1 U14107 ( .A1(n11837), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n11629) );
  NOR2_X1 U14108 ( .A1(n11624), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n11625) );
  OR2_X1 U14109 ( .A1(n11640), .A2(n11625), .ZN(n14118) );
  INV_X1 U14110 ( .A(n14118), .ZN(n14648) );
  NAND2_X1 U14111 ( .A1(n11839), .A2(n14648), .ZN(n11628) );
  NAND2_X1 U14112 ( .A1(n11808), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n11627) );
  NAND2_X1 U14113 ( .A1(n12113), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n11626) );
  NAND4_X1 U14114 ( .A1(n11629), .A2(n11628), .A3(n11627), .A4(n11626), .ZN(
        n14665) );
  NAND2_X1 U14115 ( .A1(n14665), .A2(n6664), .ZN(n11630) );
  NAND2_X1 U14116 ( .A1(n11631), .A2(n11630), .ZN(n11632) );
  XNOR2_X1 U14117 ( .A(n11632), .B(n11778), .ZN(n11635) );
  AND2_X1 U14118 ( .A1(n14665), .A2(n10688), .ZN(n11633) );
  AOI21_X1 U14119 ( .B1(n14773), .B2(n6664), .A(n11633), .ZN(n11634) );
  NAND2_X1 U14120 ( .A1(n11635), .A2(n11634), .ZN(n11636) );
  OAI21_X1 U14121 ( .B1(n11635), .B2(n11634), .A(n11636), .ZN(n14112) );
  INV_X1 U14122 ( .A(n11636), .ZN(n14124) );
  NAND2_X1 U14123 ( .A1(n11637), .A2(n11286), .ZN(n11639) );
  AOI22_X1 U14124 ( .A1(n12110), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n11657), 
        .B2(n14347), .ZN(n11638) );
  NAND2_X1 U14125 ( .A1(n14769), .A2(n11832), .ZN(n11647) );
  NAND2_X1 U14126 ( .A1(n12112), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n11645) );
  OR2_X1 U14127 ( .A1(n11640), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n11641) );
  AND2_X1 U14128 ( .A1(n11663), .A2(n11641), .ZN(n14638) );
  NAND2_X1 U14129 ( .A1(n11839), .A2(n14638), .ZN(n11644) );
  NAND2_X1 U14130 ( .A1(n11808), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n11643) );
  NAND2_X1 U14131 ( .A1(n12113), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n11642) );
  NAND4_X1 U14132 ( .A1(n11645), .A2(n11644), .A3(n11643), .A4(n11642), .ZN(
        n14427) );
  NAND2_X1 U14133 ( .A1(n14427), .A2(n6664), .ZN(n11646) );
  NAND2_X1 U14134 ( .A1(n11647), .A2(n11646), .ZN(n11648) );
  XNOR2_X1 U14135 ( .A(n11648), .B(n11778), .ZN(n11650) );
  AND2_X1 U14136 ( .A1(n14427), .A2(n10688), .ZN(n11649) );
  AOI21_X1 U14137 ( .B1(n14769), .B2(n6664), .A(n11649), .ZN(n11651) );
  NAND2_X1 U14138 ( .A1(n11650), .A2(n11651), .ZN(n11655) );
  INV_X1 U14139 ( .A(n11650), .ZN(n11653) );
  INV_X1 U14140 ( .A(n11651), .ZN(n11652) );
  NAND2_X1 U14141 ( .A1(n11653), .A2(n11652), .ZN(n11654) );
  AND2_X1 U14142 ( .A1(n11655), .A2(n11654), .ZN(n14123) );
  OAI21_X1 U14143 ( .B1(n14110), .B2(n14124), .A(n14123), .ZN(n14122) );
  NAND2_X1 U14144 ( .A1(n11656), .A2(n11286), .ZN(n11659) );
  AOI22_X1 U14145 ( .A1(n12110), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n14612), 
        .B2(n11657), .ZN(n11658) );
  NAND2_X1 U14146 ( .A1(n14759), .A2(n11832), .ZN(n11670) );
  NAND2_X1 U14147 ( .A1(n11837), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n11668) );
  INV_X1 U14148 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n11661) );
  INV_X1 U14149 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n11660) );
  OAI21_X1 U14150 ( .B1(n11663), .B2(n11661), .A(n11660), .ZN(n11664) );
  NAND2_X1 U14151 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(P1_REG3_REG_19__SCAN_IN), 
        .ZN(n11662) );
  AND2_X1 U14152 ( .A1(n11664), .A2(n11678), .ZN(n14610) );
  NAND2_X1 U14153 ( .A1(n11839), .A2(n14610), .ZN(n11667) );
  NAND2_X1 U14154 ( .A1(n6658), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n11666) );
  NAND2_X1 U14155 ( .A1(n12113), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n11665) );
  NAND4_X1 U14156 ( .A1(n11668), .A2(n11667), .A3(n11666), .A4(n11665), .ZN(
        n14587) );
  NAND2_X1 U14157 ( .A1(n14587), .A2(n6664), .ZN(n11669) );
  NAND2_X1 U14158 ( .A1(n11670), .A2(n11669), .ZN(n11671) );
  XNOR2_X1 U14159 ( .A(n11671), .B(n11830), .ZN(n14070) );
  NAND2_X1 U14160 ( .A1(n14759), .A2(n6664), .ZN(n11673) );
  NAND2_X1 U14161 ( .A1(n14587), .A2(n10688), .ZN(n11672) );
  NAND2_X1 U14162 ( .A1(n11673), .A2(n11672), .ZN(n14071) );
  NAND2_X1 U14163 ( .A1(n14070), .A2(n14071), .ZN(n14141) );
  NAND2_X1 U14164 ( .A1(n11674), .A2(n11286), .ZN(n11676) );
  NAND2_X1 U14165 ( .A1(n12110), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n11675) );
  INV_X1 U14166 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n11677) );
  AND2_X1 U14167 ( .A1(n11678), .A2(n11677), .ZN(n11679) );
  OR2_X1 U14168 ( .A1(n11679), .A2(n11699), .ZN(n14589) );
  INV_X1 U14169 ( .A(n11839), .ZN(n11705) );
  INV_X1 U14170 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n13198) );
  OAI22_X1 U14171 ( .A1(n14589), .A2(n11705), .B1(n11680), .B2(n13198), .ZN(
        n11684) );
  INV_X1 U14172 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n11682) );
  NAND2_X1 U14173 ( .A1(n11808), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n11681) );
  OAI21_X1 U14174 ( .B1(n11682), .B2(n10116), .A(n11681), .ZN(n11683) );
  INV_X1 U14175 ( .A(n14606), .ZN(n14570) );
  AND2_X1 U14176 ( .A1(n14570), .A2(n10688), .ZN(n11685) );
  AOI21_X1 U14177 ( .B1(n14400), .B2(n6664), .A(n11685), .ZN(n11691) );
  OAI22_X1 U14178 ( .A1(n14749), .A2(n11722), .B1(n14606), .B2(n7915), .ZN(
        n11686) );
  XNOR2_X1 U14179 ( .A(n11686), .B(n11830), .ZN(n11692) );
  XOR2_X1 U14180 ( .A(n11691), .B(n11692), .Z(n14144) );
  INV_X1 U14181 ( .A(n14069), .ZN(n11687) );
  INV_X1 U14182 ( .A(n11688), .ZN(n14068) );
  NOR3_X1 U14183 ( .A1(n11687), .A2(n14071), .A3(n14068), .ZN(n11690) );
  NAND2_X1 U14184 ( .A1(n14069), .A2(n11688), .ZN(n14072) );
  AOI21_X1 U14185 ( .B1(n14071), .B2(n14072), .A(n14070), .ZN(n11689) );
  NOR3_X1 U14186 ( .A1(n14144), .A2(n11690), .A3(n11689), .ZN(n11694) );
  INV_X1 U14187 ( .A(n11691), .ZN(n11693) );
  NAND2_X1 U14188 ( .A1(n11696), .A2(n11286), .ZN(n11698) );
  NAND2_X1 U14189 ( .A1(n12110), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n11697) );
  NAND2_X1 U14190 ( .A1(n14743), .A2(n11832), .ZN(n11707) );
  OR2_X1 U14191 ( .A1(n11699), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n11700) );
  NAND2_X1 U14192 ( .A1(n11699), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n11717) );
  NAND2_X1 U14193 ( .A1(n11700), .A2(n11717), .ZN(n14082) );
  NAND2_X1 U14194 ( .A1(n12112), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n11702) );
  NAND2_X1 U14195 ( .A1(n6658), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n11701) );
  AND2_X1 U14196 ( .A1(n11702), .A2(n11701), .ZN(n11704) );
  NAND2_X1 U14197 ( .A1(n12113), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n11703) );
  OAI211_X1 U14198 ( .C1(n14082), .C2(n11705), .A(n11704), .B(n11703), .ZN(
        n14588) );
  NAND2_X1 U14199 ( .A1(n14588), .A2(n6664), .ZN(n11706) );
  NAND2_X1 U14200 ( .A1(n11707), .A2(n11706), .ZN(n11708) );
  XNOR2_X1 U14201 ( .A(n11708), .B(n11830), .ZN(n11712) );
  NAND2_X1 U14202 ( .A1(n14743), .A2(n6664), .ZN(n11710) );
  NAND2_X1 U14203 ( .A1(n14588), .A2(n10688), .ZN(n11709) );
  NAND2_X1 U14204 ( .A1(n11710), .A2(n11709), .ZN(n11711) );
  NOR2_X1 U14205 ( .A1(n11712), .A2(n11711), .ZN(n11713) );
  AOI21_X1 U14206 ( .B1(n11712), .B2(n11711), .A(n11713), .ZN(n14079) );
  INV_X1 U14207 ( .A(n11713), .ZN(n14162) );
  NAND2_X1 U14208 ( .A1(n11837), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n11721) );
  INV_X1 U14209 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n14168) );
  INV_X1 U14210 ( .A(n11717), .ZN(n11716) );
  NAND2_X1 U14211 ( .A1(n11716), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n11735) );
  AOI21_X1 U14212 ( .B1(n14168), .B2(n11717), .A(n11734), .ZN(n14557) );
  NAND2_X1 U14213 ( .A1(n11839), .A2(n14557), .ZN(n11720) );
  NAND2_X1 U14214 ( .A1(n11808), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n11719) );
  NAND2_X1 U14215 ( .A1(n12113), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n11718) );
  OAI22_X1 U14216 ( .A1(n14559), .A2(n11722), .B1(n14543), .B2(n7915), .ZN(
        n11723) );
  XNOR2_X1 U14217 ( .A(n11723), .B(n11778), .ZN(n11725) );
  INV_X1 U14218 ( .A(n14559), .ZN(n14160) );
  AND2_X1 U14219 ( .A1(n14569), .A2(n10688), .ZN(n11724) );
  AOI21_X1 U14220 ( .B1(n14160), .B2(n6664), .A(n11724), .ZN(n11726) );
  NAND2_X1 U14221 ( .A1(n11725), .A2(n11726), .ZN(n11730) );
  INV_X1 U14222 ( .A(n11725), .ZN(n11728) );
  INV_X1 U14223 ( .A(n11726), .ZN(n11727) );
  NAND2_X1 U14224 ( .A1(n11728), .A2(n11727), .ZN(n11729) );
  NAND2_X1 U14225 ( .A1(n11730), .A2(n11729), .ZN(n14161) );
  INV_X1 U14226 ( .A(n11730), .ZN(n14050) );
  NAND2_X1 U14227 ( .A1(n12110), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n11732) );
  NAND2_X1 U14228 ( .A1(n14730), .A2(n11832), .ZN(n11742) );
  NAND2_X1 U14229 ( .A1(n12112), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n11740) );
  INV_X1 U14230 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n11736) );
  AOI21_X1 U14231 ( .B1(n11736), .B2(n11735), .A(n11753), .ZN(n14544) );
  NAND2_X1 U14232 ( .A1(n11839), .A2(n14544), .ZN(n11739) );
  NAND2_X1 U14233 ( .A1(n12113), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n11738) );
  NAND2_X1 U14234 ( .A1(n11808), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n11737) );
  NAND4_X1 U14235 ( .A1(n11740), .A2(n11739), .A3(n11738), .A4(n11737), .ZN(
        n14440) );
  NAND2_X1 U14236 ( .A1(n14440), .A2(n6664), .ZN(n11741) );
  NAND2_X1 U14237 ( .A1(n11742), .A2(n11741), .ZN(n11743) );
  XNOR2_X1 U14238 ( .A(n11743), .B(n11778), .ZN(n11745) );
  AND2_X1 U14239 ( .A1(n14440), .A2(n10688), .ZN(n11744) );
  AOI21_X1 U14240 ( .B1(n14730), .B2(n6664), .A(n11744), .ZN(n11746) );
  NAND2_X1 U14241 ( .A1(n11745), .A2(n11746), .ZN(n14133) );
  INV_X1 U14242 ( .A(n11745), .ZN(n11748) );
  INV_X1 U14243 ( .A(n11746), .ZN(n11747) );
  NAND2_X1 U14244 ( .A1(n11748), .A2(n11747), .ZN(n11749) );
  AND2_X1 U14245 ( .A1(n14133), .A2(n11749), .ZN(n14049) );
  NAND2_X1 U14246 ( .A1(n11750), .A2(n11286), .ZN(n11752) );
  NAND2_X1 U14247 ( .A1(n12110), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n11751) );
  NAND2_X1 U14248 ( .A1(n14724), .A2(n11832), .ZN(n11760) );
  NAND2_X1 U14249 ( .A1(n11837), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n11758) );
  NAND2_X1 U14250 ( .A1(P1_REG3_REG_24__SCAN_IN), .A2(n11753), .ZN(n11771) );
  OAI21_X1 U14251 ( .B1(P1_REG3_REG_24__SCAN_IN), .B2(n11753), .A(n11771), 
        .ZN(n11754) );
  INV_X1 U14252 ( .A(n11754), .ZN(n14529) );
  NAND2_X1 U14253 ( .A1(n11839), .A2(n14529), .ZN(n11757) );
  NAND2_X1 U14254 ( .A1(n11808), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n11756) );
  NAND2_X1 U14255 ( .A1(n12113), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n11755) );
  NAND4_X1 U14256 ( .A1(n11758), .A2(n11757), .A3(n11756), .A4(n11755), .ZN(
        n14541) );
  NAND2_X1 U14257 ( .A1(n14541), .A2(n6664), .ZN(n11759) );
  NAND2_X1 U14258 ( .A1(n11760), .A2(n11759), .ZN(n11761) );
  XNOR2_X1 U14259 ( .A(n11761), .B(n11778), .ZN(n11763) );
  AND2_X1 U14260 ( .A1(n14541), .A2(n10688), .ZN(n11762) );
  AOI21_X1 U14261 ( .B1(n14724), .B2(n6664), .A(n11762), .ZN(n11764) );
  NAND2_X1 U14262 ( .A1(n11763), .A2(n11764), .ZN(n11768) );
  INV_X1 U14263 ( .A(n11763), .ZN(n11766) );
  INV_X1 U14264 ( .A(n11764), .ZN(n11765) );
  NAND2_X1 U14265 ( .A1(n11766), .A2(n11765), .ZN(n11767) );
  NAND2_X1 U14266 ( .A1(n11768), .A2(n11767), .ZN(n14132) );
  INV_X1 U14267 ( .A(n11768), .ZN(n14101) );
  NAND2_X1 U14268 ( .A1(n14035), .A2(n11286), .ZN(n11770) );
  NAND2_X1 U14269 ( .A1(n12110), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n11769) );
  NAND2_X1 U14270 ( .A1(n14514), .A2(n11832), .ZN(n11777) );
  NAND2_X1 U14271 ( .A1(n12112), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n11775) );
  INV_X1 U14272 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n14106) );
  AOI21_X1 U14273 ( .B1(n14106), .B2(n11771), .A(n11789), .ZN(n14508) );
  NAND2_X1 U14274 ( .A1(n11839), .A2(n14508), .ZN(n11774) );
  NAND2_X1 U14275 ( .A1(n6658), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n11773) );
  NAND2_X1 U14276 ( .A1(n12113), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n11772) );
  NAND4_X1 U14277 ( .A1(n11775), .A2(n11774), .A3(n11773), .A4(n11772), .ZN(
        n14443) );
  NAND2_X1 U14278 ( .A1(n14443), .A2(n6664), .ZN(n11776) );
  NAND2_X1 U14279 ( .A1(n11777), .A2(n11776), .ZN(n11779) );
  XNOR2_X1 U14280 ( .A(n11779), .B(n11778), .ZN(n11781) );
  AND2_X1 U14281 ( .A1(n14443), .A2(n10688), .ZN(n11780) );
  AOI21_X1 U14282 ( .B1(n14514), .B2(n6664), .A(n11780), .ZN(n11782) );
  NAND2_X1 U14283 ( .A1(n11781), .A2(n11782), .ZN(n11786) );
  INV_X1 U14284 ( .A(n11781), .ZN(n11784) );
  INV_X1 U14285 ( .A(n11782), .ZN(n11783) );
  NAND2_X1 U14286 ( .A1(n11784), .A2(n11783), .ZN(n11785) );
  OAI21_X1 U14287 ( .B1(n14136), .B2(n14101), .A(n14100), .ZN(n14099) );
  NAND2_X1 U14288 ( .A1(n14099), .A2(n11786), .ZN(n14193) );
  NAND2_X1 U14289 ( .A1(n14032), .A2(n11286), .ZN(n11788) );
  NAND2_X1 U14290 ( .A1(n12110), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n11787) );
  NAND2_X1 U14291 ( .A1(n14499), .A2(n11832), .ZN(n11796) );
  NAND2_X1 U14292 ( .A1(n12112), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n11794) );
  INV_X1 U14293 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n14199) );
  INV_X1 U14294 ( .A(n11789), .ZN(n11790) );
  NAND2_X1 U14295 ( .A1(n11789), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n11807) );
  AOI21_X1 U14296 ( .B1(n14199), .B2(n11790), .A(n11824), .ZN(n14495) );
  NAND2_X1 U14297 ( .A1(n11839), .A2(n14495), .ZN(n11793) );
  NAND2_X1 U14298 ( .A1(n11808), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n11792) );
  NAND2_X1 U14299 ( .A1(n12113), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n11791) );
  NAND4_X1 U14300 ( .A1(n11794), .A2(n11793), .A3(n11792), .A4(n11791), .ZN(
        n14444) );
  NAND2_X1 U14301 ( .A1(n14444), .A2(n6664), .ZN(n11795) );
  NAND2_X1 U14302 ( .A1(n11796), .A2(n11795), .ZN(n11797) );
  XNOR2_X1 U14303 ( .A(n11797), .B(n11830), .ZN(n11801) );
  NAND2_X1 U14304 ( .A1(n14499), .A2(n6664), .ZN(n11799) );
  NAND2_X1 U14305 ( .A1(n14444), .A2(n10688), .ZN(n11798) );
  NAND2_X1 U14306 ( .A1(n11799), .A2(n11798), .ZN(n11800) );
  NOR2_X1 U14307 ( .A1(n11801), .A2(n11800), .ZN(n11802) );
  AOI21_X1 U14308 ( .B1(n11801), .B2(n11800), .A(n11802), .ZN(n14194) );
  INV_X1 U14309 ( .A(n11802), .ZN(n11803) );
  NAND2_X1 U14310 ( .A1(n11804), .A2(n11286), .ZN(n11806) );
  NAND2_X1 U14311 ( .A1(n12110), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n11805) );
  NAND2_X1 U14312 ( .A1(n14705), .A2(n11832), .ZN(n11814) );
  NAND2_X1 U14313 ( .A1(n12112), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n11812) );
  XNOR2_X1 U14314 ( .A(P1_REG3_REG_27__SCAN_IN), .B(n11807), .ZN(n14479) );
  NAND2_X1 U14315 ( .A1(n11839), .A2(n14479), .ZN(n11811) );
  NAND2_X1 U14316 ( .A1(n11808), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n11810) );
  NAND2_X1 U14317 ( .A1(n12113), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n11809) );
  NAND4_X1 U14318 ( .A1(n11812), .A2(n11811), .A3(n11810), .A4(n11809), .ZN(
        n14447) );
  NAND2_X1 U14319 ( .A1(n14447), .A2(n6664), .ZN(n11813) );
  NAND2_X1 U14320 ( .A1(n11814), .A2(n11813), .ZN(n11815) );
  XNOR2_X1 U14321 ( .A(n11815), .B(n11830), .ZN(n11819) );
  NAND2_X1 U14322 ( .A1(n14705), .A2(n6664), .ZN(n11817) );
  NAND2_X1 U14323 ( .A1(n14447), .A2(n10688), .ZN(n11816) );
  NAND2_X1 U14324 ( .A1(n11817), .A2(n11816), .ZN(n11818) );
  NOR2_X1 U14325 ( .A1(n11819), .A2(n11818), .ZN(n11820) );
  AOI21_X1 U14326 ( .B1(n11819), .B2(n11818), .A(n11820), .ZN(n14043) );
  NAND2_X1 U14327 ( .A1(n14024), .A2(n11286), .ZN(n11822) );
  NAND2_X1 U14328 ( .A1(n12110), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n11821) );
  NAND2_X1 U14329 ( .A1(n11837), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n11829) );
  INV_X1 U14330 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n13441) );
  NAND2_X1 U14331 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(n11824), .ZN(n11823) );
  NAND2_X1 U14332 ( .A1(n13441), .A2(n11823), .ZN(n11825) );
  NAND3_X1 U14333 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .A3(n11824), .ZN(n11838) );
  AND2_X1 U14334 ( .A1(n11825), .A2(n11838), .ZN(n11844) );
  NAND2_X1 U14335 ( .A1(n11839), .A2(n11844), .ZN(n11828) );
  NAND2_X1 U14336 ( .A1(n6658), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n11827) );
  NAND2_X1 U14337 ( .A1(n12113), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n11826) );
  NAND4_X1 U14338 ( .A1(n11829), .A2(n11828), .A3(n11827), .A4(n11826), .ZN(
        n14687) );
  AOI22_X1 U14339 ( .A1(n14468), .A2(n6664), .B1(n10688), .B2(n14687), .ZN(
        n11831) );
  XNOR2_X1 U14340 ( .A(n11831), .B(n11830), .ZN(n11834) );
  AOI22_X1 U14341 ( .A1(n14468), .A2(n11832), .B1(n6664), .B2(n14687), .ZN(
        n11833) );
  XNOR2_X1 U14342 ( .A(n11834), .B(n11833), .ZN(n11835) );
  XNOR2_X1 U14343 ( .A(n11836), .B(n11835), .ZN(n11849) );
  NAND2_X1 U14344 ( .A1(n11837), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n11843) );
  INV_X1 U14345 ( .A(n11838), .ZN(n14410) );
  NAND2_X1 U14346 ( .A1(n11839), .A2(n14410), .ZN(n11842) );
  NAND2_X1 U14347 ( .A1(n6658), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n11841) );
  NAND2_X1 U14348 ( .A1(n12113), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n11840) );
  NAND4_X1 U14349 ( .A1(n11843), .A2(n11842), .A3(n11841), .A4(n11840), .ZN(
        n14216) );
  INV_X1 U14350 ( .A(n11844), .ZN(n14466) );
  NOR2_X1 U14351 ( .A1(n15176), .A2(n14466), .ZN(n11846) );
  INV_X1 U14352 ( .A(n14447), .ZN(n14456) );
  OAI22_X1 U14353 ( .A1(n14456), .A2(n15161), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13441), .ZN(n11845) );
  AOI211_X1 U14354 ( .C1(n14207), .C2(n14216), .A(n11846), .B(n11845), .ZN(
        n11848) );
  NAND2_X1 U14355 ( .A1(n14468), .A2(n15172), .ZN(n11847) );
  OAI211_X1 U14356 ( .C1(n11849), .C2(n15167), .A(n11848), .B(n11847), .ZN(
        P1_U3220) );
  NAND2_X1 U14357 ( .A1(n11850), .A2(n12578), .ZN(n11851) );
  NAND2_X1 U14358 ( .A1(n11852), .A2(n11851), .ZN(n11856) );
  AOI22_X1 U14359 ( .A1(n12867), .A2(n12618), .B1(n12245), .B2(n12869), .ZN(
        n11855) );
  NOR2_X1 U14360 ( .A1(n12996), .A2(n12898), .ZN(n11858) );
  INV_X1 U14361 ( .A(P3_REG2_REG_27__SCAN_IN), .ZN(n13373) );
  OAI22_X1 U14362 ( .A1(n15719), .A2(n13373), .B1(n12242), .B2(n15711), .ZN(
        n11857) );
  AOI211_X1 U14363 ( .C1(n12925), .C2(n15716), .A(n11858), .B(n11857), .ZN(
        n11859) );
  OAI21_X1 U14364 ( .B1(n12927), .B2(n15703), .A(n11859), .ZN(P3_U3206) );
  OAI222_X1 U14365 ( .A1(n14031), .A2(n11861), .B1(n6670), .B2(P2_U3088), .C1(
        n11860), .C2(n14038), .ZN(P2_U3307) );
  INV_X1 U14366 ( .A(n11862), .ZN(n11863) );
  OAI222_X1 U14367 ( .A1(n14038), .A2(n11864), .B1(n14031), .B2(n11863), .C1(
        P2_U3088), .C2(n9173), .ZN(P2_U3305) );
  INV_X1 U14368 ( .A(n11868), .ZN(n11871) );
  INV_X1 U14369 ( .A(n11869), .ZN(n11870) );
  XNOR2_X1 U14370 ( .A(n15127), .B(n13075), .ZN(n11872) );
  NAND2_X1 U14371 ( .A1(n13564), .A2(n11865), .ZN(n11873) );
  NAND2_X1 U14372 ( .A1(n11872), .A2(n11873), .ZN(n11877) );
  INV_X1 U14373 ( .A(n11872), .ZN(n11875) );
  INV_X1 U14374 ( .A(n11873), .ZN(n11874) );
  NAND2_X1 U14375 ( .A1(n11875), .A2(n11874), .ZN(n11876) );
  AND2_X1 U14376 ( .A1(n11877), .A2(n11876), .ZN(n15122) );
  XNOR2_X1 U14377 ( .A(n13991), .B(n13075), .ZN(n11879) );
  NOR2_X2 U14378 ( .A1(n11880), .A2(n11879), .ZN(n11878) );
  INV_X1 U14379 ( .A(n11878), .ZN(n11881) );
  NAND2_X1 U14380 ( .A1(n13643), .A2(n11865), .ZN(n11882) );
  XNOR2_X1 U14381 ( .A(n13985), .B(n13107), .ZN(n11883) );
  NAND2_X1 U14382 ( .A1(n13670), .A2(n11865), .ZN(n11884) );
  XNOR2_X1 U14383 ( .A(n11883), .B(n11884), .ZN(n13504) );
  INV_X1 U14384 ( .A(n11883), .ZN(n11885) );
  NAND2_X1 U14385 ( .A1(n11885), .A2(n11884), .ZN(n11886) );
  NAND2_X1 U14386 ( .A1(n13507), .A2(n11886), .ZN(n13517) );
  XNOR2_X1 U14387 ( .A(n13673), .B(n13075), .ZN(n11887) );
  NAND2_X1 U14388 ( .A1(n13672), .A2(n11865), .ZN(n11888) );
  NAND2_X1 U14389 ( .A1(n11887), .A2(n11888), .ZN(n11892) );
  INV_X1 U14390 ( .A(n11887), .ZN(n11890) );
  INV_X1 U14391 ( .A(n11888), .ZN(n11889) );
  NAND2_X1 U14392 ( .A1(n11890), .A2(n11889), .ZN(n11891) );
  AND2_X1 U14393 ( .A1(n11892), .A2(n11891), .ZN(n13518) );
  XNOR2_X1 U14394 ( .A(n13845), .B(n13075), .ZN(n11894) );
  NAND2_X1 U14395 ( .A1(n13675), .A2(n11865), .ZN(n11895) );
  XNOR2_X1 U14396 ( .A(n11894), .B(n11895), .ZN(n13543) );
  INV_X1 U14397 ( .A(n13543), .ZN(n11893) );
  INV_X1 U14398 ( .A(n11894), .ZN(n11897) );
  INV_X1 U14399 ( .A(n11895), .ZN(n11896) );
  NAND2_X1 U14400 ( .A1(n11897), .A2(n11896), .ZN(n11898) );
  XNOR2_X1 U14401 ( .A(n13965), .B(n13107), .ZN(n11901) );
  INV_X1 U14402 ( .A(n11901), .ZN(n11899) );
  NAND2_X1 U14403 ( .A1(n11900), .A2(n11899), .ZN(n11904) );
  NAND2_X1 U14404 ( .A1(n11902), .A2(n11901), .ZN(n11903) );
  XNOR2_X1 U14405 ( .A(n13681), .B(n13075), .ZN(n11907) );
  NAND2_X1 U14406 ( .A1(n13680), .A2(n11865), .ZN(n11906) );
  XNOR2_X1 U14407 ( .A(n11907), .B(n11906), .ZN(n13532) );
  XNOR2_X1 U14408 ( .A(n13953), .B(n13107), .ZN(n11911) );
  NAND2_X1 U14409 ( .A1(n13684), .A2(n11865), .ZN(n11909) );
  XNOR2_X1 U14410 ( .A(n11911), .B(n11909), .ZN(n13117) );
  INV_X1 U14411 ( .A(n11909), .ZN(n11910) );
  XNOR2_X1 U14412 ( .A(n13947), .B(n13107), .ZN(n13064) );
  OAI22_X1 U14413 ( .A1(n11913), .A2(n13630), .B1(n11912), .B2(n13496), .ZN(
        n13794) );
  AOI22_X1 U14414 ( .A1(n13794), .A2(n15125), .B1(P2_REG3_REG_22__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11914) );
  OAI21_X1 U14415 ( .B1(n13797), .B2(n15131), .A(n11914), .ZN(n11917) );
  NAND2_X1 U14416 ( .A1(n15123), .A2(n11865), .ZN(n11934) );
  NOR3_X1 U14417 ( .A1(n11915), .A2(n13685), .A3(n11934), .ZN(n11916) );
  AOI211_X1 U14418 ( .C1(n13947), .C2(n15128), .A(n11917), .B(n11916), .ZN(
        n11918) );
  OAI21_X1 U14419 ( .B1(n13063), .B2(n13561), .A(n11918), .ZN(P2_U3207) );
  NAND2_X1 U14420 ( .A1(n14806), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n11919) );
  NAND2_X1 U14421 ( .A1(n11920), .A2(n11919), .ZN(n12388) );
  INV_X1 U14422 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n14803) );
  NAND2_X1 U14423 ( .A1(n14803), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n12389) );
  INV_X1 U14424 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n12190) );
  NAND2_X1 U14425 ( .A1(n12190), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n11921) );
  AND2_X1 U14426 ( .A1(n12389), .A2(n11921), .ZN(n12387) );
  INV_X1 U14427 ( .A(n12387), .ZN(n11922) );
  XNOR2_X1 U14428 ( .A(n12388), .B(n11922), .ZN(n12380) );
  INV_X1 U14429 ( .A(n12380), .ZN(n11923) );
  INV_X1 U14430 ( .A(SI_30_), .ZN(n12378) );
  OAI222_X1 U14431 ( .A1(P3_U3151), .A2(n8014), .B1(n14938), .B2(n11923), .C1(
        n12378), .C2(n14936), .ZN(P3_U3265) );
  NAND2_X1 U14432 ( .A1(n13556), .A2(n11925), .ZN(n11926) );
  NAND2_X1 U14433 ( .A1(P2_U3088), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n15470)
         );
  OAI211_X1 U14434 ( .C1(n11927), .C2(n13558), .A(n11926), .B(n15470), .ZN(
        n11929) );
  NOR3_X1 U14435 ( .A1(n6783), .A2(n13667), .A3(n11934), .ZN(n11928) );
  AOI211_X1 U14436 ( .C1(n13991), .C2(n15128), .A(n11929), .B(n11928), .ZN(
        n11930) );
  OAI21_X1 U14437 ( .B1(n11924), .B2(n13561), .A(n11930), .ZN(P2_U3213) );
  NAND2_X1 U14438 ( .A1(P2_U3088), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n13626)
         );
  NAND2_X1 U14439 ( .A1(n13680), .A2(n13555), .ZN(n11932) );
  NAND2_X1 U14440 ( .A1(n13675), .A2(n13701), .ZN(n11931) );
  NAND2_X1 U14441 ( .A1(n11932), .A2(n11931), .ZN(n13964) );
  NAND2_X1 U14442 ( .A1(n15125), .A2(n13964), .ZN(n11933) );
  OAI211_X1 U14443 ( .C1(n15131), .C2(n13831), .A(n13626), .B(n11933), .ZN(
        n11937) );
  NOR3_X1 U14444 ( .A1(n11935), .A2(n7745), .A3(n11934), .ZN(n11936) );
  AOI211_X1 U14445 ( .C1(n13965), .C2(n15128), .A(n11937), .B(n11936), .ZN(
        n11938) );
  OAI21_X1 U14446 ( .B1(n13533), .B2(n13561), .A(n11938), .ZN(P2_U3191) );
  INV_X1 U14447 ( .A(P3_REG2_REG_29__SCAN_IN), .ZN(n11941) );
  INV_X1 U14448 ( .A(n11939), .ZN(n11940) );
  NAND2_X1 U14449 ( .A1(n12911), .A2(n11940), .ZN(n12714) );
  OAI21_X1 U14450 ( .B1(n15719), .B2(n11941), .A(n12714), .ZN(n11944) );
  NOR2_X1 U14451 ( .A1(n11942), .A2(n12827), .ZN(n11943) );
  OAI21_X1 U14452 ( .B1(n11947), .B2(n15703), .A(n11946), .ZN(P3_U3204) );
  NAND2_X1 U14453 ( .A1(n14021), .A2(n11286), .ZN(n11949) );
  NAND2_X1 U14454 ( .A1(n12110), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n11948) );
  NAND2_X1 U14455 ( .A1(n12131), .A2(n14612), .ZN(n11950) );
  NAND2_X1 U14456 ( .A1(n11951), .A2(n11950), .ZN(n11952) );
  MUX2_X1 U14457 ( .A(n14419), .B(n14216), .S(n6663), .Z(n12104) );
  INV_X1 U14458 ( .A(n12104), .ZN(n12108) );
  MUX2_X1 U14459 ( .A(n14588), .B(n14743), .S(n12117), .Z(n12071) );
  XNOR2_X1 U14460 ( .A(n11953), .B(n12117), .ZN(n11955) );
  INV_X1 U14461 ( .A(n12150), .ZN(n11954) );
  OAI211_X1 U14462 ( .C1(n12148), .C2(n11956), .A(n11955), .B(n11954), .ZN(
        n11967) );
  MUX2_X1 U14463 ( .A(n6659), .B(n11957), .S(n11959), .Z(n11968) );
  INV_X1 U14464 ( .A(n11968), .ZN(n11965) );
  AND2_X1 U14465 ( .A1(n11957), .A2(n12117), .ZN(n11958) );
  AOI21_X1 U14466 ( .B1(n6659), .B2(n6663), .A(n11958), .ZN(n11969) );
  INV_X1 U14467 ( .A(n11969), .ZN(n11964) );
  AND2_X1 U14468 ( .A1(n14229), .A2(n11959), .ZN(n11962) );
  NOR2_X1 U14469 ( .A1(n14229), .A2(n11959), .ZN(n11961) );
  INV_X1 U14470 ( .A(n11976), .ZN(n12153) );
  NAND3_X1 U14471 ( .A1(n11967), .A2(n11966), .A3(n12153), .ZN(n11980) );
  NAND2_X1 U14472 ( .A1(n11969), .A2(n11968), .ZN(n11977) );
  INV_X1 U14473 ( .A(n11970), .ZN(n11971) );
  NAND2_X1 U14474 ( .A1(n11971), .A2(n6663), .ZN(n11975) );
  INV_X1 U14475 ( .A(n11972), .ZN(n11973) );
  NAND2_X1 U14476 ( .A1(n11973), .A2(n12117), .ZN(n11974) );
  OAI211_X1 U14477 ( .C1(n11977), .C2(n11976), .A(n11975), .B(n11974), .ZN(
        n11978) );
  INV_X1 U14478 ( .A(n11978), .ZN(n11979) );
  NAND2_X1 U14479 ( .A1(n11980), .A2(n11979), .ZN(n11985) );
  MUX2_X1 U14480 ( .A(n14226), .B(n11982), .S(n12117), .Z(n11981) );
  INV_X1 U14481 ( .A(n11981), .ZN(n11984) );
  MUX2_X1 U14482 ( .A(n14226), .B(n11982), .S(n6663), .Z(n11983) );
  OAI21_X1 U14483 ( .B1(n11985), .B2(n11984), .A(n11983), .ZN(n11987) );
  NAND2_X1 U14484 ( .A1(n11985), .A2(n11984), .ZN(n11986) );
  MUX2_X1 U14485 ( .A(n14225), .B(n11988), .S(n6663), .Z(n11990) );
  MUX2_X1 U14486 ( .A(n11988), .B(n14225), .S(n6663), .Z(n11989) );
  INV_X1 U14487 ( .A(n11990), .ZN(n11991) );
  MUX2_X1 U14488 ( .A(n14224), .B(n15337), .S(n12117), .Z(n11994) );
  MUX2_X1 U14489 ( .A(n14224), .B(n15337), .S(n6663), .Z(n11992) );
  MUX2_X1 U14490 ( .A(n14223), .B(n11995), .S(n6663), .Z(n11997) );
  MUX2_X1 U14491 ( .A(n11995), .B(n14223), .S(n6663), .Z(n11996) );
  MUX2_X1 U14492 ( .A(n14222), .B(n11998), .S(n12117), .Z(n12002) );
  NAND2_X1 U14493 ( .A1(n12001), .A2(n12002), .ZN(n12000) );
  MUX2_X1 U14494 ( .A(n14222), .B(n11998), .S(n6663), .Z(n11999) );
  NAND2_X1 U14495 ( .A1(n12000), .A2(n11999), .ZN(n12006) );
  INV_X1 U14496 ( .A(n12001), .ZN(n12004) );
  INV_X1 U14497 ( .A(n12002), .ZN(n12003) );
  NAND2_X1 U14498 ( .A1(n12004), .A2(n12003), .ZN(n12005) );
  MUX2_X1 U14499 ( .A(n15377), .B(n15286), .S(n6663), .Z(n12008) );
  MUX2_X1 U14500 ( .A(n15377), .B(n15286), .S(n12117), .Z(n12007) );
  MUX2_X1 U14501 ( .A(n14221), .B(n15380), .S(n12117), .Z(n12010) );
  MUX2_X1 U14502 ( .A(n14221), .B(n15380), .S(n6663), .Z(n12009) );
  MUX2_X1 U14503 ( .A(n14220), .B(n15183), .S(n6663), .Z(n12015) );
  MUX2_X1 U14504 ( .A(n14220), .B(n15183), .S(n12117), .Z(n12012) );
  INV_X1 U14505 ( .A(n12014), .ZN(n12017) );
  INV_X1 U14506 ( .A(n12015), .ZN(n12016) );
  NAND2_X1 U14507 ( .A1(n12017), .A2(n12016), .ZN(n12019) );
  MUX2_X1 U14508 ( .A(n14219), .B(n14955), .S(n12117), .Z(n12021) );
  MUX2_X1 U14509 ( .A(n14219), .B(n14955), .S(n6663), .Z(n12018) );
  MUX2_X1 U14510 ( .A(n14218), .B(n15216), .S(n6663), .Z(n12028) );
  NAND2_X1 U14511 ( .A1(n15216), .A2(n12117), .ZN(n12022) );
  OAI211_X1 U14512 ( .C1(n12117), .C2(n15162), .A(n12028), .B(n12022), .ZN(
        n12023) );
  NAND2_X1 U14513 ( .A1(n14672), .A2(n15163), .ZN(n12146) );
  NAND2_X1 U14514 ( .A1(n12146), .A2(n12025), .ZN(n12030) );
  NAND2_X1 U14515 ( .A1(n15162), .A2(n6663), .ZN(n12026) );
  OAI21_X1 U14516 ( .B1(n15216), .B2(n6663), .A(n12026), .ZN(n12027) );
  NOR2_X1 U14517 ( .A1(n12028), .A2(n12027), .ZN(n12029) );
  AOI22_X1 U14518 ( .A1(n12030), .A2(n12117), .B1(n12147), .B2(n12029), .ZN(
        n12033) );
  NAND2_X1 U14519 ( .A1(n14394), .A2(n14660), .ZN(n12031) );
  NAND2_X1 U14520 ( .A1(n12031), .A2(n6663), .ZN(n12032) );
  MUX2_X1 U14521 ( .A(n12146), .B(n14394), .S(n12117), .Z(n12035) );
  XNOR2_X1 U14522 ( .A(n14769), .B(n14427), .ZN(n14632) );
  MUX2_X1 U14523 ( .A(n14665), .B(n14773), .S(n6663), .Z(n12043) );
  NAND2_X1 U14524 ( .A1(n14632), .A2(n12043), .ZN(n12040) );
  INV_X1 U14525 ( .A(n14427), .ZN(n12037) );
  OR2_X1 U14526 ( .A1(n14769), .A2(n12037), .ZN(n14396) );
  AND2_X1 U14527 ( .A1(n14665), .A2(n6663), .ZN(n12036) );
  AOI21_X1 U14528 ( .B1(n14773), .B2(n12117), .A(n12036), .ZN(n12039) );
  NAND2_X1 U14529 ( .A1(n14769), .A2(n12037), .ZN(n12038) );
  NAND3_X1 U14530 ( .A1(n14396), .A2(n12039), .A3(n12038), .ZN(n12048) );
  NAND2_X1 U14531 ( .A1(n12040), .A2(n12048), .ZN(n12041) );
  NAND2_X1 U14532 ( .A1(n12042), .A2(n12041), .ZN(n12051) );
  INV_X1 U14533 ( .A(n12043), .ZN(n12047) );
  AND2_X1 U14534 ( .A1(n14427), .A2(n12117), .ZN(n12045) );
  OAI21_X1 U14535 ( .B1(n12117), .B2(n14427), .A(n14769), .ZN(n12044) );
  OAI21_X1 U14536 ( .B1(n12045), .B2(n14769), .A(n12044), .ZN(n12046) );
  OAI21_X1 U14537 ( .B1(n12048), .B2(n12047), .A(n12046), .ZN(n12049) );
  INV_X1 U14538 ( .A(n12049), .ZN(n12050) );
  NAND2_X1 U14539 ( .A1(n12051), .A2(n12050), .ZN(n12054) );
  INV_X1 U14540 ( .A(n14587), .ZN(n14146) );
  NAND2_X1 U14541 ( .A1(n14759), .A2(n14146), .ZN(n14398) );
  OR2_X1 U14542 ( .A1(n14759), .A2(n14146), .ZN(n12052) );
  NAND2_X1 U14543 ( .A1(n14398), .A2(n12052), .ZN(n14604) );
  INV_X1 U14544 ( .A(n14604), .ZN(n14600) );
  INV_X1 U14545 ( .A(n14217), .ZN(n14608) );
  OR2_X1 U14546 ( .A1(n14762), .A2(n14608), .ZN(n14397) );
  NAND2_X1 U14547 ( .A1(n14762), .A2(n14608), .ZN(n12053) );
  INV_X1 U14548 ( .A(n14759), .ZN(n14381) );
  NAND2_X1 U14549 ( .A1(n14587), .A2(n12117), .ZN(n12056) );
  OAI21_X1 U14550 ( .B1(n14397), .B2(n6663), .A(n12056), .ZN(n12058) );
  NAND2_X1 U14551 ( .A1(n14762), .A2(n14217), .ZN(n14430) );
  NOR2_X1 U14552 ( .A1(n14587), .A2(n12117), .ZN(n12059) );
  NAND3_X1 U14553 ( .A1(n14430), .A2(n12059), .A3(n14762), .ZN(n12055) );
  OAI21_X1 U14554 ( .B1(n14397), .B2(n12056), .A(n12055), .ZN(n12057) );
  AOI21_X1 U14555 ( .B1(n14381), .B2(n12058), .A(n12057), .ZN(n12064) );
  NAND3_X1 U14556 ( .A1(n14430), .A2(n6663), .A3(n14762), .ZN(n12061) );
  INV_X1 U14557 ( .A(n12059), .ZN(n12060) );
  NAND2_X1 U14558 ( .A1(n12061), .A2(n12060), .ZN(n12062) );
  NAND2_X1 U14559 ( .A1(n12062), .A2(n14759), .ZN(n12063) );
  MUX2_X1 U14560 ( .A(n14570), .B(n14400), .S(n6663), .Z(n12066) );
  MUX2_X1 U14561 ( .A(n14606), .B(n14749), .S(n12117), .Z(n12065) );
  NAND2_X1 U14562 ( .A1(n12070), .A2(n12071), .ZN(n12068) );
  MUX2_X1 U14563 ( .A(n14588), .B(n14743), .S(n6663), .Z(n12067) );
  NAND2_X1 U14564 ( .A1(n12068), .A2(n12067), .ZN(n12069) );
  OAI21_X1 U14565 ( .B1(n12071), .B2(n12070), .A(n12069), .ZN(n12074) );
  MUX2_X1 U14566 ( .A(n14541), .B(n14724), .S(n6663), .Z(n12080) );
  MUX2_X1 U14567 ( .A(n14541), .B(n14724), .S(n12117), .Z(n12077) );
  NAND2_X1 U14568 ( .A1(n12078), .A2(n12077), .ZN(n12084) );
  INV_X1 U14569 ( .A(n12079), .ZN(n12082) );
  INV_X1 U14570 ( .A(n12080), .ZN(n12081) );
  MUX2_X1 U14571 ( .A(n14443), .B(n14514), .S(n12117), .Z(n12087) );
  MUX2_X1 U14572 ( .A(n14443), .B(n14514), .S(n6663), .Z(n12085) );
  INV_X1 U14573 ( .A(n12087), .ZN(n12088) );
  MUX2_X1 U14574 ( .A(n14444), .B(n14499), .S(n6663), .Z(n12090) );
  MUX2_X1 U14575 ( .A(n14444), .B(n14499), .S(n12117), .Z(n12089) );
  INV_X1 U14576 ( .A(n12090), .ZN(n12091) );
  MUX2_X1 U14577 ( .A(n14447), .B(n14705), .S(n12117), .Z(n12095) );
  MUX2_X1 U14578 ( .A(n14447), .B(n14705), .S(n6663), .Z(n12092) );
  NAND2_X1 U14579 ( .A1(n12093), .A2(n12092), .ZN(n12099) );
  INV_X1 U14580 ( .A(n12094), .ZN(n12097) );
  INV_X1 U14581 ( .A(n12095), .ZN(n12096) );
  NAND2_X1 U14582 ( .A1(n12097), .A2(n12096), .ZN(n12098) );
  INV_X1 U14583 ( .A(n14687), .ZN(n14414) );
  INV_X1 U14584 ( .A(n14468), .ZN(n14700) );
  MUX2_X1 U14585 ( .A(n14414), .B(n14700), .S(n6663), .Z(n12101) );
  MUX2_X1 U14586 ( .A(n14468), .B(n14687), .S(n6663), .Z(n12100) );
  INV_X1 U14587 ( .A(n12101), .ZN(n12102) );
  INV_X1 U14588 ( .A(n12105), .ZN(n12107) );
  INV_X1 U14589 ( .A(n14216), .ZN(n14457) );
  INV_X1 U14590 ( .A(n14419), .ZN(n14690) );
  MUX2_X1 U14591 ( .A(n14457), .B(n14690), .S(n6663), .Z(n12103) );
  AOI21_X1 U14592 ( .B1(n12105), .B2(n12104), .A(n12103), .ZN(n12106) );
  INV_X1 U14593 ( .A(n12124), .ZN(n12127) );
  NAND2_X1 U14594 ( .A1(n12110), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n12111) );
  NAND2_X1 U14595 ( .A1(n12112), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n12116) );
  NAND2_X1 U14596 ( .A1(n12113), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n12115) );
  NAND2_X1 U14597 ( .A1(n6658), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n12114) );
  NAND3_X1 U14598 ( .A1(n12116), .A2(n12115), .A3(n12114), .ZN(n14386) );
  NAND2_X1 U14599 ( .A1(n14386), .A2(n12117), .ZN(n12137) );
  AOI21_X1 U14600 ( .B1(n12118), .B2(n12137), .A(n14408), .ZN(n12119) );
  AOI21_X1 U14601 ( .B1(n14682), .B2(n11959), .A(n12119), .ZN(n12123) );
  INV_X1 U14602 ( .A(n12123), .ZN(n12126) );
  INV_X1 U14603 ( .A(n14386), .ZN(n12136) );
  AOI21_X1 U14604 ( .B1(n12136), .B2(n12120), .A(n14408), .ZN(n12121) );
  MUX2_X1 U14605 ( .A(n14682), .B(n12121), .S(n6663), .Z(n12122) );
  NAND2_X1 U14606 ( .A1(n14017), .A2(n11286), .ZN(n12129) );
  NAND2_X1 U14607 ( .A1(n12110), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n12128) );
  XNOR2_X1 U14608 ( .A(n14679), .B(n12136), .ZN(n12175) );
  AND2_X1 U14609 ( .A1(n12131), .A2(n12130), .ZN(n12133) );
  OAI21_X1 U14610 ( .B1(n12134), .B2(n12133), .A(n12132), .ZN(n12174) );
  INV_X1 U14611 ( .A(n12137), .ZN(n12138) );
  NOR2_X1 U14612 ( .A1(n12139), .A2(n12138), .ZN(n12178) );
  NAND2_X1 U14613 ( .A1(n12141), .A2(n12140), .ZN(n12173) );
  NAND2_X1 U14614 ( .A1(n12174), .A2(n12173), .ZN(n12176) );
  XOR2_X1 U14615 ( .A(n14408), .B(n14682), .Z(n12170) );
  INV_X1 U14616 ( .A(n14444), .ZN(n12142) );
  INV_X1 U14617 ( .A(n14541), .ZN(n12143) );
  NAND2_X1 U14618 ( .A1(n14559), .A2(n14569), .ZN(n12144) );
  NAND2_X1 U14619 ( .A1(n14403), .A2(n12144), .ZN(n14561) );
  INV_X1 U14620 ( .A(n14561), .ZN(n14553) );
  INV_X1 U14621 ( .A(n14440), .ZN(n12145) );
  XNOR2_X1 U14622 ( .A(n14730), .B(n12145), .ZN(n14535) );
  INV_X1 U14623 ( .A(n14535), .ZN(n14539) );
  OR2_X1 U14624 ( .A1(n14762), .A2(n14217), .ZN(n14432) );
  NAND2_X1 U14625 ( .A1(n14432), .A2(n14430), .ZN(n14622) );
  NAND2_X1 U14626 ( .A1(n14394), .A2(n12146), .ZN(n14659) );
  NOR4_X1 U14627 ( .A1(n12150), .A2(n12149), .A3(n12148), .A4(n7141), .ZN(
        n12154) );
  NAND4_X1 U14628 ( .A1(n12154), .A2(n12153), .A3(n12152), .A4(n12151), .ZN(
        n12155) );
  NOR4_X1 U14629 ( .A1(n12158), .A2(n12157), .A3(n12156), .A4(n12155), .ZN(
        n12160) );
  NAND4_X1 U14630 ( .A1(n12160), .A2(n12159), .A3(n15178), .A4(n15276), .ZN(
        n12161) );
  NOR4_X1 U14631 ( .A1(n14659), .A2(n12162), .A3(n11480), .A4(n12161), .ZN(
        n12163) );
  XNOR2_X1 U14632 ( .A(n14773), .B(n14665), .ZN(n14645) );
  NAND4_X1 U14633 ( .A1(n14622), .A2(n12163), .A3(n14632), .A4(n14645), .ZN(
        n12165) );
  XNOR2_X1 U14634 ( .A(n14749), .B(n14606), .ZN(n14595) );
  INV_X1 U14635 ( .A(n14595), .ZN(n12164) );
  NOR3_X1 U14636 ( .A1(n12165), .A2(n12164), .A3(n14604), .ZN(n12166) );
  XNOR2_X1 U14637 ( .A(n14743), .B(n14588), .ZN(n14579) );
  NAND4_X1 U14638 ( .A1(n14553), .A2(n14539), .A3(n12166), .A4(n14579), .ZN(
        n12167) );
  NOR4_X1 U14639 ( .A1(n14491), .A2(n14503), .A3(n14525), .A4(n12167), .ZN(
        n12169) );
  NAND2_X1 U14640 ( .A1(n14468), .A2(n14687), .ZN(n14449) );
  OR2_X1 U14641 ( .A1(n14468), .A2(n14687), .ZN(n12168) );
  NAND4_X1 U14642 ( .A1(n12170), .A2(n12169), .A3(n14454), .A4(n14484), .ZN(
        n12171) );
  XNOR2_X1 U14643 ( .A(n14419), .B(n14457), .ZN(n14450) );
  NOR3_X1 U14644 ( .A1(n12175), .A2(n12171), .A3(n14450), .ZN(n12172) );
  INV_X1 U14645 ( .A(n12174), .ZN(n12181) );
  INV_X1 U14646 ( .A(n12175), .ZN(n12177) );
  NOR2_X1 U14647 ( .A1(n12177), .A2(n12176), .ZN(n12180) );
  INV_X1 U14648 ( .A(n12178), .ZN(n12179) );
  NAND3_X1 U14649 ( .A1(n12186), .A2(n6667), .A3(n15378), .ZN(n12187) );
  OAI211_X1 U14650 ( .C1(n9763), .C2(n12189), .A(n12187), .B(P1_B_REG_SCAN_IN), 
        .ZN(n12188) );
  OAI222_X1 U14651 ( .A1(n14031), .A2(n14802), .B1(n12191), .B2(P2_U3088), 
        .C1(n12190), .C2(n14038), .ZN(P2_U3297) );
  XNOR2_X1 U14652 ( .A(n12582), .B(n12234), .ZN(n12192) );
  NOR2_X1 U14653 ( .A1(n12192), .A2(n12722), .ZN(n12269) );
  AOI21_X1 U14654 ( .B1(n12192), .B2(n12722), .A(n12269), .ZN(n12238) );
  NAND2_X1 U14655 ( .A1(n12194), .A2(n12193), .ZN(n12290) );
  NAND2_X1 U14656 ( .A1(n12290), .A2(n12288), .ZN(n12195) );
  XNOR2_X1 U14657 ( .A(n13044), .B(n12234), .ZN(n12196) );
  XNOR2_X1 U14658 ( .A(n12196), .B(n12628), .ZN(n12287) );
  NAND2_X1 U14659 ( .A1(n12195), .A2(n12287), .ZN(n12292) );
  INV_X1 U14660 ( .A(n12628), .ZN(n15020) );
  NAND2_X1 U14661 ( .A1(n15020), .A2(n12196), .ZN(n12197) );
  XNOR2_X1 U14662 ( .A(n12198), .B(n12234), .ZN(n15014) );
  XNOR2_X1 U14663 ( .A(n15105), .B(n12234), .ZN(n12247) );
  AND2_X1 U14664 ( .A1(n12247), .A2(n15018), .ZN(n12200) );
  INV_X1 U14665 ( .A(n12247), .ZN(n12201) );
  XNOR2_X1 U14666 ( .A(n13040), .B(n12270), .ZN(n12363) );
  INV_X1 U14667 ( .A(n12363), .ZN(n12203) );
  NAND2_X1 U14668 ( .A1(n12203), .A2(n12362), .ZN(n12204) );
  XNOR2_X1 U14669 ( .A(n15005), .B(n12270), .ZN(n12205) );
  XNOR2_X1 U14670 ( .A(n12205), .B(n12856), .ZN(n15004) );
  INV_X1 U14671 ( .A(n12205), .ZN(n12206) );
  XNOR2_X1 U14672 ( .A(n13032), .B(n12270), .ZN(n12207) );
  XNOR2_X1 U14673 ( .A(n12207), .B(n12844), .ZN(n12309) );
  NAND2_X1 U14674 ( .A1(n12310), .A2(n12309), .ZN(n12308) );
  NAND2_X1 U14675 ( .A1(n12207), .A2(n12870), .ZN(n12208) );
  XNOR2_X1 U14676 ( .A(n12343), .B(n12270), .ZN(n12209) );
  XNOR2_X1 U14677 ( .A(n12209), .B(n12625), .ZN(n12345) );
  INV_X1 U14678 ( .A(n12209), .ZN(n12210) );
  NAND2_X1 U14679 ( .A1(n12210), .A2(n12625), .ZN(n12211) );
  XNOR2_X1 U14680 ( .A(n12411), .B(n12234), .ZN(n12212) );
  AND2_X1 U14681 ( .A1(n12212), .A2(n12624), .ZN(n12261) );
  INV_X1 U14682 ( .A(n12212), .ZN(n12213) );
  NAND2_X1 U14683 ( .A1(n12213), .A2(n12845), .ZN(n12260) );
  XNOR2_X1 U14684 ( .A(n12954), .B(n12270), .ZN(n12215) );
  XNOR2_X1 U14685 ( .A(n12215), .B(n12216), .ZN(n12326) );
  XNOR2_X1 U14686 ( .A(n13018), .B(n12234), .ZN(n12218) );
  NAND2_X1 U14687 ( .A1(n12218), .A2(n12217), .ZN(n12221) );
  INV_X1 U14688 ( .A(n12218), .ZN(n12219) );
  NAND2_X1 U14689 ( .A1(n12219), .A2(n12622), .ZN(n12220) );
  NAND2_X1 U14690 ( .A1(n12221), .A2(n12220), .ZN(n12279) );
  XNOR2_X1 U14691 ( .A(n12338), .B(n12270), .ZN(n12223) );
  XNOR2_X1 U14692 ( .A(n12318), .B(n12270), .ZN(n12225) );
  NAND2_X1 U14693 ( .A1(n12225), .A2(n12224), .ZN(n12228) );
  INV_X1 U14694 ( .A(n12225), .ZN(n12226) );
  NAND2_X1 U14695 ( .A1(n12226), .A2(n6985), .ZN(n12227) );
  NAND2_X1 U14696 ( .A1(n12228), .A2(n12227), .ZN(n12319) );
  INV_X1 U14697 ( .A(n12228), .ZN(n12300) );
  XNOR2_X1 U14698 ( .A(n12296), .B(n12270), .ZN(n12230) );
  NAND2_X1 U14699 ( .A1(n12230), .A2(n12229), .ZN(n12233) );
  INV_X1 U14700 ( .A(n12230), .ZN(n12231) );
  NAND2_X1 U14701 ( .A1(n12231), .A2(n12619), .ZN(n12232) );
  OAI21_X1 U14702 ( .B1(n12298), .B2(n12300), .A(n12299), .ZN(n12297) );
  XNOR2_X1 U14703 ( .A(n12747), .B(n12234), .ZN(n12235) );
  NOR2_X1 U14704 ( .A1(n12235), .A2(n12618), .ZN(n12236) );
  AOI21_X1 U14705 ( .B1(n12235), .B2(n12618), .A(n12236), .ZN(n12355) );
  INV_X1 U14706 ( .A(n12236), .ZN(n12237) );
  OAI22_X1 U14707 ( .A1(n12349), .A2(n12241), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12240), .ZN(n12244) );
  NOR2_X1 U14708 ( .A1(n15593), .A2(n12242), .ZN(n12243) );
  AOI211_X1 U14709 ( .C1(n12347), .C2(n12245), .A(n12244), .B(n12243), .ZN(
        n12246) );
  XNOR2_X1 U14710 ( .A(n12247), .B(n15018), .ZN(n12248) );
  XNOR2_X1 U14711 ( .A(n12249), .B(n12248), .ZN(n12253) );
  NOR2_X1 U14712 ( .A1(n15105), .A2(n15581), .ZN(n12251) );
  AOI22_X1 U14713 ( .A1(n12867), .A2(n15013), .B1(n12868), .B2(n12869), .ZN(
        n12892) );
  NAND2_X1 U14714 ( .A1(P3_REG3_REG_14__SCAN_IN), .A2(P3_U3151), .ZN(n15672)
         );
  OAI21_X1 U14715 ( .B1(n12892), .B2(n15009), .A(n15672), .ZN(n12250) );
  AOI211_X1 U14716 ( .C1(n15002), .C2(n12896), .A(n12251), .B(n12250), .ZN(
        n12252) );
  OAI21_X1 U14717 ( .B1(n12253), .B2(n15585), .A(n12252), .ZN(P3_U3155) );
  INV_X1 U14718 ( .A(n12563), .ZN(n13010) );
  OAI21_X1 U14719 ( .B1(n12562), .B2(n12254), .A(n12320), .ZN(n12255) );
  NAND2_X1 U14720 ( .A1(n12255), .A2(n15021), .ZN(n12259) );
  INV_X1 U14721 ( .A(n12256), .ZN(n12789) );
  AOI22_X1 U14722 ( .A1(n6985), .A2(n12869), .B1(n12867), .B2(n12621), .ZN(
        n12786) );
  OAI22_X1 U14723 ( .A1(n12786), .A2(n15009), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n13426), .ZN(n12257) );
  AOI21_X1 U14724 ( .B1(n12789), .B2(n15002), .A(n12257), .ZN(n12258) );
  OAI211_X1 U14725 ( .C1(n13010), .C2(n15581), .A(n12259), .B(n12258), .ZN(
        P3_U3156) );
  NOR2_X1 U14726 ( .A1(n7289), .A2(n12261), .ZN(n12262) );
  XNOR2_X1 U14727 ( .A(n12263), .B(n12262), .ZN(n12268) );
  AOI22_X1 U14728 ( .A1(n12867), .A2(n12625), .B1(n12623), .B2(n12869), .ZN(
        n12831) );
  OAI22_X1 U14729 ( .A1(n12831), .A2(n15009), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12264), .ZN(n12266) );
  INV_X1 U14730 ( .A(n12411), .ZN(n13025) );
  NOR2_X1 U14731 ( .A1(n13025), .A2(n15581), .ZN(n12265) );
  AOI211_X1 U14732 ( .C1(n15002), .C2(n12835), .A(n12266), .B(n12265), .ZN(
        n12267) );
  OAI21_X1 U14733 ( .B1(n12268), .B2(n15585), .A(n12267), .ZN(P3_U3159) );
  XOR2_X1 U14734 ( .A(n12270), .B(n12728), .Z(n12271) );
  OR2_X1 U14735 ( .A1(n12993), .A2(n15581), .ZN(n12275) );
  AOI22_X1 U14736 ( .A1(n12311), .A2(n12722), .B1(P3_REG3_REG_28__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12274) );
  NAND2_X1 U14737 ( .A1(n15002), .A2(n12730), .ZN(n12273) );
  NAND2_X1 U14738 ( .A1(n12347), .A2(n12721), .ZN(n12272) );
  OAI21_X1 U14739 ( .B1(n12277), .B2(n15585), .A(n12276), .ZN(P3_U3160) );
  AOI21_X1 U14740 ( .B1(n12279), .B2(n12278), .A(n6794), .ZN(n12285) );
  NOR2_X1 U14741 ( .A1(n15593), .A2(n12810), .ZN(n12282) );
  AOI22_X1 U14742 ( .A1(n12623), .A2(n12867), .B1(n12869), .B2(n12621), .ZN(
        n12806) );
  INV_X1 U14743 ( .A(P3_REG3_REG_21__SCAN_IN), .ZN(n12280) );
  OAI22_X1 U14744 ( .A1(n12806), .A2(n15009), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12280), .ZN(n12281) );
  AOI211_X1 U14745 ( .C1(n12283), .C2(n15012), .A(n12282), .B(n12281), .ZN(
        n12284) );
  OAI21_X1 U14746 ( .B1(n12285), .B2(n15585), .A(n12284), .ZN(P3_U3163) );
  AOI22_X1 U14747 ( .A1(n15013), .A2(n12869), .B1(n12867), .B2(n12629), .ZN(
        n12905) );
  NAND2_X1 U14748 ( .A1(P3_REG3_REG_12__SCAN_IN), .A2(P3_U3151), .ZN(n15637)
         );
  NAND2_X1 U14749 ( .A1(n15012), .A2(n12912), .ZN(n12286) );
  OAI211_X1 U14750 ( .C1(n12905), .C2(n15009), .A(n15637), .B(n12286), .ZN(
        n12294) );
  INV_X1 U14751 ( .A(n12287), .ZN(n12289) );
  NAND3_X1 U14752 ( .A1(n12290), .A2(n12289), .A3(n12288), .ZN(n12291) );
  AOI21_X1 U14753 ( .B1(n12292), .B2(n12291), .A(n15585), .ZN(n12293) );
  AOI211_X1 U14754 ( .C1(n15002), .C2(n12910), .A(n12294), .B(n12293), .ZN(
        n12295) );
  INV_X1 U14755 ( .A(n12295), .ZN(P3_U3164) );
  INV_X1 U14756 ( .A(n12297), .ZN(n12302) );
  NOR3_X1 U14757 ( .A1(n12298), .A2(n12300), .A3(n12299), .ZN(n12301) );
  OAI21_X1 U14758 ( .B1(n12302), .B2(n12301), .A(n15021), .ZN(n12307) );
  INV_X1 U14759 ( .A(n12303), .ZN(n12760) );
  AOI22_X1 U14760 ( .A1(n6985), .A2(n12867), .B1(n12869), .B2(n12618), .ZN(
        n12755) );
  INV_X1 U14761 ( .A(P3_REG3_REG_25__SCAN_IN), .ZN(n12304) );
  OAI22_X1 U14762 ( .A1(n12755), .A2(n15009), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12304), .ZN(n12305) );
  AOI21_X1 U14763 ( .B1(n15002), .B2(n12760), .A(n12305), .ZN(n12306) );
  OAI211_X1 U14764 ( .C1(n13003), .C2(n15581), .A(n12307), .B(n12306), .ZN(
        P3_U3165) );
  OAI211_X1 U14765 ( .C1(n12310), .C2(n12309), .A(n12308), .B(n15021), .ZN(
        n12317) );
  INV_X1 U14766 ( .A(n12861), .ZN(n12315) );
  AOI22_X1 U14767 ( .A1(n12311), .A2(n12626), .B1(P3_REG3_REG_17__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12312) );
  OAI21_X1 U14768 ( .B1(n12857), .B2(n12313), .A(n12312), .ZN(n12314) );
  AOI21_X1 U14769 ( .B1(n15002), .B2(n12315), .A(n12314), .ZN(n12316) );
  OAI211_X1 U14770 ( .C1(n15581), .C2(n13032), .A(n12317), .B(n12316), .ZN(
        P3_U3168) );
  AND3_X1 U14771 ( .A1(n12320), .A2(n6679), .A3(n12319), .ZN(n12321) );
  OAI21_X1 U14772 ( .B1(n12298), .B2(n12321), .A(n15021), .ZN(n12325) );
  INV_X1 U14773 ( .A(n12322), .ZN(n12774) );
  AOI22_X1 U14774 ( .A1(n12619), .A2(n12869), .B1(n12867), .B2(n12620), .ZN(
        n12767) );
  INV_X1 U14775 ( .A(P3_REG3_REG_24__SCAN_IN), .ZN(n13454) );
  OAI22_X1 U14776 ( .A1(n12767), .A2(n15009), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n13454), .ZN(n12323) );
  AOI21_X1 U14777 ( .B1(n15002), .B2(n12774), .A(n12323), .ZN(n12324) );
  OAI211_X1 U14778 ( .C1(n6986), .C2(n15581), .A(n12325), .B(n12324), .ZN(
        P3_U3169) );
  XNOR2_X1 U14779 ( .A(n12327), .B(n12326), .ZN(n12332) );
  NOR2_X1 U14780 ( .A1(n15593), .A2(n12821), .ZN(n12330) );
  AOI22_X1 U14781 ( .A1(n12622), .A2(n12869), .B1(n12867), .B2(n12624), .ZN(
        n12819) );
  OAI22_X1 U14782 ( .A1(n12819), .A2(n15009), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12328), .ZN(n12329) );
  AOI211_X1 U14783 ( .C1(n12954), .C2(n15012), .A(n12330), .B(n12329), .ZN(
        n12331) );
  OAI21_X1 U14784 ( .B1(n12332), .B2(n15585), .A(n12331), .ZN(P3_U3173) );
  INV_X1 U14785 ( .A(n12333), .ZN(n12334) );
  AOI21_X1 U14786 ( .B1(n12621), .B2(n12335), .A(n12334), .ZN(n12342) );
  INV_X1 U14787 ( .A(n12336), .ZN(n12800) );
  AOI22_X1 U14788 ( .A1(n12622), .A2(n12867), .B1(n12869), .B2(n12620), .ZN(
        n12796) );
  INV_X1 U14789 ( .A(P3_REG3_REG_22__SCAN_IN), .ZN(n12337) );
  OAI22_X1 U14790 ( .A1(n12796), .A2(n15009), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12337), .ZN(n12340) );
  INV_X1 U14791 ( .A(n12338), .ZN(n13014) );
  NOR2_X1 U14792 ( .A1(n13014), .A2(n15581), .ZN(n12339) );
  AOI211_X1 U14793 ( .C1(n15002), .C2(n12800), .A(n12340), .B(n12339), .ZN(
        n12341) );
  OAI21_X1 U14794 ( .B1(n12342), .B2(n15585), .A(n12341), .ZN(P3_U3175) );
  INV_X1 U14795 ( .A(n12343), .ZN(n13029) );
  OAI211_X1 U14796 ( .C1(n12346), .C2(n12345), .A(n12344), .B(n15021), .ZN(
        n12352) );
  NAND2_X1 U14797 ( .A1(P3_U3151), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n15086)
         );
  NAND2_X1 U14798 ( .A1(n12347), .A2(n12624), .ZN(n12348) );
  OAI211_X1 U14799 ( .C1(n12349), .C2(n12844), .A(n15086), .B(n12348), .ZN(
        n12350) );
  AOI21_X1 U14800 ( .B1(n15002), .B2(n12848), .A(n12350), .ZN(n12351) );
  OAI211_X1 U14801 ( .C1(n13029), .C2(n15581), .A(n12352), .B(n12351), .ZN(
        P3_U3178) );
  OAI21_X1 U14802 ( .B1(n12355), .B2(n12354), .A(n12353), .ZN(n12356) );
  NAND2_X1 U14803 ( .A1(n12356), .A2(n15021), .ZN(n12361) );
  INV_X1 U14804 ( .A(n12744), .ZN(n12359) );
  AOI22_X1 U14805 ( .A1(n12619), .A2(n12867), .B1(n12869), .B2(n12722), .ZN(
        n12742) );
  INV_X1 U14806 ( .A(P3_REG3_REG_26__SCAN_IN), .ZN(n12357) );
  OAI22_X1 U14807 ( .A1(n12742), .A2(n15009), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12357), .ZN(n12358) );
  AOI21_X1 U14808 ( .B1(n15002), .B2(n12359), .A(n12358), .ZN(n12360) );
  OAI211_X1 U14809 ( .C1(n12999), .C2(n15581), .A(n12361), .B(n12360), .ZN(
        P3_U3180) );
  XNOR2_X1 U14810 ( .A(n12363), .B(n12362), .ZN(n12364) );
  XNOR2_X1 U14811 ( .A(n12365), .B(n12364), .ZN(n12375) );
  NAND2_X1 U14812 ( .A1(n12626), .A2(n12869), .ZN(n12367) );
  NAND2_X1 U14813 ( .A1(n12627), .A2(n12867), .ZN(n12366) );
  AND2_X1 U14814 ( .A1(n12367), .A2(n12366), .ZN(n12882) );
  INV_X1 U14815 ( .A(n12368), .ZN(n12886) );
  NAND2_X1 U14816 ( .A1(n15002), .A2(n12886), .ZN(n12371) );
  INV_X1 U14817 ( .A(P3_REG3_REG_15__SCAN_IN), .ZN(n12369) );
  NOR2_X1 U14818 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n12369), .ZN(n15030) );
  INV_X1 U14819 ( .A(n15030), .ZN(n12370) );
  OAI211_X1 U14820 ( .C1(n12882), .C2(n15009), .A(n12371), .B(n12370), .ZN(
        n12372) );
  AOI21_X1 U14821 ( .B1(n12373), .B2(n15012), .A(n12372), .ZN(n12374) );
  OAI21_X1 U14822 ( .B1(n12375), .B2(n15585), .A(n12374), .ZN(P3_U3181) );
  INV_X1 U14823 ( .A(n12591), .ZN(n12376) );
  NOR2_X1 U14824 ( .A1(n12377), .A2(n12376), .ZN(n12400) );
  NOR2_X1 U14825 ( .A1(n8066), .A2(n12378), .ZN(n12379) );
  AOI21_X1 U14826 ( .B1(n12380), .B2(n12394), .A(n12379), .ZN(n12432) );
  NAND2_X1 U14827 ( .A1(n12381), .A2(P3_REG1_REG_31__SCAN_IN), .ZN(n12385) );
  NAND2_X1 U14828 ( .A1(n8059), .A2(P3_REG0_REG_31__SCAN_IN), .ZN(n12384) );
  NAND2_X1 U14829 ( .A1(n12382), .A2(P3_REG2_REG_31__SCAN_IN), .ZN(n12383) );
  INV_X1 U14830 ( .A(n12713), .ZN(n12616) );
  AND2_X1 U14831 ( .A1(n12617), .A2(n12616), .ZN(n12397) );
  NAND2_X1 U14832 ( .A1(n12388), .A2(n12387), .ZN(n12390) );
  NAND2_X1 U14833 ( .A1(n12390), .A2(n12389), .ZN(n12393) );
  INV_X1 U14834 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n12391) );
  XNOR2_X1 U14835 ( .A(n12391), .B(P2_DATAO_REG_31__SCAN_IN), .ZN(n12392) );
  XNOR2_X1 U14836 ( .A(n12393), .B(n12392), .ZN(n13053) );
  NAND2_X1 U14837 ( .A1(n13053), .A2(n12394), .ZN(n12396) );
  INV_X1 U14838 ( .A(SI_31_), .ZN(n13057) );
  OR2_X1 U14839 ( .A1(n8066), .A2(n13057), .ZN(n12395) );
  NAND2_X1 U14840 ( .A1(n12396), .A2(n12395), .ZN(n12404) );
  OR2_X1 U14841 ( .A1(n12404), .A2(n12713), .ZN(n12403) );
  OAI211_X1 U14842 ( .C1(n12432), .C2(n12397), .A(n12403), .B(n12590), .ZN(
        n12399) );
  AND2_X1 U14843 ( .A1(n12432), .A2(n12617), .ZN(n12405) );
  NOR2_X1 U14844 ( .A1(n12405), .A2(n12713), .ZN(n12398) );
  OAI22_X1 U14845 ( .A1(n12400), .A2(n12399), .B1(n12990), .B2(n12398), .ZN(
        n12401) );
  XNOR2_X1 U14846 ( .A(n12401), .B(n12706), .ZN(n12609) );
  INV_X1 U14847 ( .A(n12402), .ZN(n12608) );
  INV_X1 U14848 ( .A(n12403), .ZN(n12599) );
  NAND2_X1 U14849 ( .A1(n12404), .A2(n12713), .ZN(n12407) );
  INV_X1 U14850 ( .A(n12405), .ZN(n12406) );
  NAND2_X1 U14851 ( .A1(n12407), .A2(n12406), .ZN(n12598) );
  NAND2_X1 U14852 ( .A1(n12558), .A2(n12559), .ZN(n12798) );
  INV_X1 U14853 ( .A(n12408), .ZN(n12410) );
  NAND2_X1 U14854 ( .A1(n12410), .A2(n12409), .ZN(n12808) );
  XNOR2_X1 U14855 ( .A(n12411), .B(n12845), .ZN(n12833) );
  NOR2_X1 U14856 ( .A1(n12457), .A2(n15692), .ZN(n12413) );
  INV_X1 U14857 ( .A(n15705), .ZN(n15707) );
  NAND4_X1 U14858 ( .A1(n12413), .A2(n12503), .A3(n12412), .A4(n15707), .ZN(
        n12415) );
  NOR2_X1 U14859 ( .A1(n12415), .A2(n12414), .ZN(n12423) );
  NOR2_X1 U14860 ( .A1(n12417), .A2(n12416), .ZN(n12418) );
  NAND4_X1 U14861 ( .A1(n12418), .A2(n12477), .A3(n12462), .A4(n12483), .ZN(
        n12420) );
  NAND2_X1 U14862 ( .A1(n12908), .A2(n12489), .ZN(n12419) );
  NOR2_X1 U14863 ( .A1(n12420), .A2(n12419), .ZN(n12422) );
  INV_X1 U14864 ( .A(n12516), .ZN(n12421) );
  NAND4_X1 U14865 ( .A1(n12884), .A2(n12423), .A3(n12422), .A4(n6693), .ZN(
        n12424) );
  NOR2_X1 U14866 ( .A1(n12424), .A2(n12894), .ZN(n12425) );
  NAND4_X1 U14867 ( .A1(n12846), .A2(n12859), .A3(n12874), .A4(n12425), .ZN(
        n12426) );
  NOR2_X1 U14868 ( .A1(n12833), .A2(n12426), .ZN(n12427) );
  NAND3_X1 U14869 ( .A1(n12808), .A2(n12825), .A3(n12427), .ZN(n12428) );
  NOR2_X1 U14870 ( .A1(n12798), .A2(n12428), .ZN(n12429) );
  NAND4_X1 U14871 ( .A1(n12757), .A2(n7853), .A3(n12429), .A4(n12782), .ZN(
        n12430) );
  NOR2_X1 U14872 ( .A1(n12430), .A2(n12740), .ZN(n12431) );
  NAND4_X1 U14873 ( .A1(n6713), .A2(n12728), .A3(n12431), .A4(n12578), .ZN(
        n12434) );
  INV_X1 U14874 ( .A(n12432), .ZN(n15102) );
  INV_X1 U14875 ( .A(n12617), .ZN(n12433) );
  AND2_X1 U14876 ( .A1(n15102), .A2(n12433), .ZN(n12596) );
  XNOR2_X1 U14877 ( .A(n12435), .B(n12706), .ZN(n12603) );
  NAND2_X1 U14878 ( .A1(n12722), .A2(n12585), .ZN(n12581) );
  INV_X1 U14879 ( .A(n12436), .ZN(n12437) );
  NAND2_X1 U14880 ( .A1(n12437), .A2(n12442), .ZN(n12439) );
  AND2_X1 U14881 ( .A1(n12439), .A2(n12438), .ZN(n12446) );
  NAND3_X1 U14882 ( .A1(n12442), .A2(n12441), .A3(n12440), .ZN(n12443) );
  NAND3_X1 U14883 ( .A1(n12446), .A2(n12448), .A3(n12443), .ZN(n12445) );
  NAND3_X1 U14884 ( .A1(n12445), .A2(n12455), .A3(n12444), .ZN(n12450) );
  INV_X1 U14885 ( .A(n12446), .ZN(n12447) );
  AND2_X1 U14886 ( .A1(n12448), .A2(n12447), .ZN(n12449) );
  MUX2_X1 U14887 ( .A(n12450), .B(n12449), .S(n12593), .Z(n12451) );
  NAND2_X1 U14888 ( .A1(n12451), .A2(n12453), .ZN(n12460) );
  NAND2_X1 U14889 ( .A1(n12453), .A2(n12452), .ZN(n12454) );
  NAND2_X1 U14890 ( .A1(n12454), .A2(n12593), .ZN(n12459) );
  NOR2_X1 U14891 ( .A1(n12455), .A2(n12585), .ZN(n12456) );
  OR2_X1 U14892 ( .A1(n12457), .A2(n12456), .ZN(n12458) );
  AOI21_X1 U14893 ( .B1(n12460), .B2(n12459), .A(n12458), .ZN(n12466) );
  NAND2_X1 U14894 ( .A1(n12462), .A2(n12461), .ZN(n12464) );
  OAI211_X1 U14895 ( .C1(n12466), .C2(n12464), .A(n12478), .B(n12463), .ZN(
        n12465) );
  NAND2_X1 U14896 ( .A1(n12465), .A2(n12471), .ZN(n12476) );
  INV_X1 U14897 ( .A(n12466), .ZN(n12474) );
  INV_X1 U14898 ( .A(n12467), .ZN(n12469) );
  NOR2_X1 U14899 ( .A1(n12469), .A2(n12468), .ZN(n12473) );
  NAND2_X1 U14900 ( .A1(n12471), .A2(n12470), .ZN(n12472) );
  AOI21_X1 U14901 ( .B1(n12474), .B2(n12473), .A(n12472), .ZN(n12475) );
  MUX2_X1 U14902 ( .A(n12476), .B(n12475), .S(n12585), .Z(n12485) );
  OAI21_X1 U14903 ( .B1(n12593), .B2(n12478), .A(n12477), .ZN(n12484) );
  NAND2_X1 U14904 ( .A1(n15756), .A2(n12593), .ZN(n12481) );
  NAND2_X1 U14905 ( .A1(n12479), .A2(n12585), .ZN(n12480) );
  MUX2_X1 U14906 ( .A(n12481), .B(n12480), .S(n12633), .Z(n12482) );
  OAI211_X1 U14907 ( .C1(n12485), .C2(n12484), .A(n12483), .B(n12482), .ZN(
        n12490) );
  MUX2_X1 U14908 ( .A(n12487), .B(n12486), .S(n12593), .Z(n12488) );
  NAND3_X1 U14909 ( .A1(n12490), .A2(n12489), .A3(n12488), .ZN(n12496) );
  INV_X1 U14910 ( .A(n12491), .ZN(n12493) );
  MUX2_X1 U14911 ( .A(n12493), .B(n12492), .S(n12593), .Z(n12494) );
  INV_X1 U14912 ( .A(n12494), .ZN(n12495) );
  NAND2_X1 U14913 ( .A1(n12496), .A2(n12495), .ZN(n12504) );
  NAND2_X1 U14914 ( .A1(n15580), .A2(n12585), .ZN(n12500) );
  NAND2_X1 U14915 ( .A1(n12497), .A2(n12593), .ZN(n12499) );
  MUX2_X1 U14916 ( .A(n12500), .B(n12499), .S(n12498), .Z(n12501) );
  NAND2_X1 U14917 ( .A1(n12501), .A2(n8172), .ZN(n12502) );
  AOI21_X1 U14918 ( .B1(n12504), .B2(n12503), .A(n12502), .ZN(n12513) );
  NAND2_X1 U14919 ( .A1(n12510), .A2(n12505), .ZN(n12508) );
  NAND2_X1 U14920 ( .A1(n12509), .A2(n12506), .ZN(n12507) );
  MUX2_X1 U14921 ( .A(n12508), .B(n12507), .S(n12593), .Z(n12512) );
  MUX2_X1 U14922 ( .A(n12510), .B(n12509), .S(n12585), .Z(n12511) );
  OAI211_X1 U14923 ( .C1(n12513), .C2(n12512), .A(n6693), .B(n12511), .ZN(
        n12519) );
  INV_X1 U14924 ( .A(n12894), .ZN(n12518) );
  INV_X1 U14925 ( .A(n12514), .ZN(n12515) );
  MUX2_X1 U14926 ( .A(n12516), .B(n12515), .S(n12585), .Z(n12517) );
  NAND3_X1 U14927 ( .A1(n12519), .A2(n12518), .A3(n12517), .ZN(n12522) );
  NAND2_X1 U14928 ( .A1(n7408), .A2(n12593), .ZN(n12521) );
  INV_X1 U14929 ( .A(n12884), .ZN(n12880) );
  AOI21_X1 U14930 ( .B1(n12522), .B2(n12521), .A(n12880), .ZN(n12528) );
  INV_X1 U14931 ( .A(n12524), .ZN(n12525) );
  AOI21_X1 U14932 ( .B1(n12884), .B2(n8219), .A(n12525), .ZN(n12526) );
  AOI21_X1 U14933 ( .B1(n12526), .B2(n12532), .A(n12593), .ZN(n12527) );
  OAI21_X1 U14934 ( .B1(n12528), .B2(n12527), .A(n12530), .ZN(n12535) );
  NAND2_X1 U14935 ( .A1(n12530), .A2(n12529), .ZN(n12531) );
  NAND2_X1 U14936 ( .A1(n12531), .A2(n12593), .ZN(n12534) );
  NOR2_X1 U14937 ( .A1(n12532), .A2(n12585), .ZN(n12533) );
  AOI21_X1 U14938 ( .B1(n12535), .B2(n12534), .A(n12533), .ZN(n12540) );
  NAND3_X1 U14939 ( .A1(n12542), .A2(n12870), .A3(n13032), .ZN(n12537) );
  NAND3_X1 U14940 ( .A1(n12537), .A2(n12593), .A3(n12536), .ZN(n12538) );
  NOR2_X1 U14941 ( .A1(n12547), .A2(n12538), .ZN(n12541) );
  OAI22_X1 U14942 ( .A1(n12540), .A2(n12854), .B1(n12541), .B2(n12539), .ZN(
        n12545) );
  INV_X1 U14943 ( .A(n12541), .ZN(n12544) );
  NAND3_X1 U14944 ( .A1(n12546), .A2(n12542), .A3(n12585), .ZN(n12543) );
  AOI22_X1 U14945 ( .A1(n12545), .A2(n12846), .B1(n12544), .B2(n12543), .ZN(
        n12549) );
  MUX2_X1 U14946 ( .A(n12547), .B(n8291), .S(n12593), .Z(n12548) );
  OR3_X1 U14947 ( .A1(n12549), .A2(n12548), .A3(n7058), .ZN(n12553) );
  MUX2_X1 U14948 ( .A(n12551), .B(n12550), .S(n12593), .Z(n12552) );
  NAND3_X1 U14949 ( .A1(n12553), .A2(n12552), .A3(n12808), .ZN(n12557) );
  INV_X1 U14950 ( .A(n12798), .ZN(n12794) );
  MUX2_X1 U14951 ( .A(n12555), .B(n12554), .S(n12593), .Z(n12556) );
  NAND3_X1 U14952 ( .A1(n12557), .A2(n12794), .A3(n12556), .ZN(n12561) );
  MUX2_X1 U14953 ( .A(n12559), .B(n12558), .S(n12593), .Z(n12560) );
  NAND3_X1 U14954 ( .A1(n12561), .A2(n12782), .A3(n12560), .ZN(n12565) );
  NAND3_X1 U14955 ( .A1(n12563), .A2(n12562), .A3(n12593), .ZN(n12564) );
  AOI21_X1 U14956 ( .B1(n12565), .B2(n12564), .A(n12769), .ZN(n12570) );
  XNOR2_X1 U14957 ( .A(n12566), .B(n12593), .ZN(n12567) );
  NOR2_X1 U14958 ( .A1(n12568), .A2(n12567), .ZN(n12569) );
  OAI21_X1 U14959 ( .B1(n12570), .B2(n12569), .A(n12757), .ZN(n12574) );
  INV_X1 U14960 ( .A(n12740), .ZN(n12573) );
  MUX2_X1 U14961 ( .A(n12571), .B(n12736), .S(n12593), .Z(n12572) );
  NAND3_X1 U14962 ( .A1(n12574), .A2(n12573), .A3(n12572), .ZN(n12579) );
  MUX2_X1 U14963 ( .A(n12576), .B(n12575), .S(n12593), .Z(n12577) );
  NAND3_X1 U14964 ( .A1(n12579), .A2(n12578), .A3(n12577), .ZN(n12580) );
  OAI21_X1 U14965 ( .B1(n12582), .B2(n12581), .A(n12580), .ZN(n12583) );
  NAND2_X1 U14966 ( .A1(n12583), .A2(n12728), .ZN(n12589) );
  NAND2_X1 U14967 ( .A1(n12584), .A2(n12586), .ZN(n12587) );
  NAND3_X1 U14968 ( .A1(n12589), .A2(n6713), .A3(n12588), .ZN(n12592) );
  AND2_X1 U14969 ( .A1(n12592), .A2(n12590), .ZN(n12595) );
  NAND2_X1 U14970 ( .A1(n12592), .A2(n12591), .ZN(n12594) );
  INV_X1 U14971 ( .A(n12596), .ZN(n12597) );
  INV_X1 U14972 ( .A(n12598), .ZN(n12600) );
  AOI21_X1 U14973 ( .B1(n12601), .B2(n12600), .A(n12599), .ZN(n12606) );
  OAI22_X1 U14974 ( .A1(n12604), .A2(n12603), .B1(n12606), .B2(n12602), .ZN(
        n12605) );
  NAND4_X1 U14975 ( .A1(n12867), .A2(n12611), .A3(n12610), .A4(n12696), .ZN(
        n12612) );
  OAI211_X1 U14976 ( .C1(n12613), .C2(n12615), .A(n12612), .B(P3_B_REG_SCAN_IN), .ZN(n12614) );
  MUX2_X1 U14977 ( .A(P3_DATAO_REG_31__SCAN_IN), .B(n12616), .S(n15577), .Z(
        P3_U3522) );
  MUX2_X1 U14978 ( .A(P3_DATAO_REG_30__SCAN_IN), .B(n12617), .S(n15577), .Z(
        P3_U3521) );
  MUX2_X1 U14979 ( .A(P3_DATAO_REG_27__SCAN_IN), .B(n12722), .S(n15577), .Z(
        P3_U3518) );
  MUX2_X1 U14980 ( .A(P3_DATAO_REG_26__SCAN_IN), .B(n12618), .S(n15577), .Z(
        P3_U3517) );
  MUX2_X1 U14981 ( .A(P3_DATAO_REG_25__SCAN_IN), .B(n12619), .S(n15577), .Z(
        P3_U3516) );
  MUX2_X1 U14982 ( .A(P3_DATAO_REG_23__SCAN_IN), .B(n12620), .S(n15577), .Z(
        P3_U3514) );
  MUX2_X1 U14983 ( .A(P3_DATAO_REG_22__SCAN_IN), .B(n12621), .S(n15577), .Z(
        P3_U3513) );
  MUX2_X1 U14984 ( .A(P3_DATAO_REG_21__SCAN_IN), .B(n12622), .S(n15577), .Z(
        P3_U3512) );
  MUX2_X1 U14985 ( .A(P3_DATAO_REG_20__SCAN_IN), .B(n12623), .S(P3_U3897), .Z(
        P3_U3511) );
  MUX2_X1 U14986 ( .A(P3_DATAO_REG_19__SCAN_IN), .B(n12624), .S(n15577), .Z(
        P3_U3510) );
  MUX2_X1 U14987 ( .A(P3_DATAO_REG_18__SCAN_IN), .B(n12625), .S(P3_U3897), .Z(
        P3_U3509) );
  MUX2_X1 U14988 ( .A(P3_DATAO_REG_17__SCAN_IN), .B(n12870), .S(P3_U3897), .Z(
        P3_U3508) );
  MUX2_X1 U14989 ( .A(P3_DATAO_REG_16__SCAN_IN), .B(n12626), .S(P3_U3897), .Z(
        P3_U3507) );
  MUX2_X1 U14990 ( .A(P3_DATAO_REG_15__SCAN_IN), .B(n12868), .S(P3_U3897), .Z(
        P3_U3506) );
  MUX2_X1 U14991 ( .A(P3_DATAO_REG_14__SCAN_IN), .B(n12627), .S(P3_U3897), .Z(
        P3_U3505) );
  MUX2_X1 U14992 ( .A(P3_DATAO_REG_13__SCAN_IN), .B(n15013), .S(P3_U3897), .Z(
        P3_U3504) );
  MUX2_X1 U14993 ( .A(P3_DATAO_REG_12__SCAN_IN), .B(n12628), .S(P3_U3897), .Z(
        P3_U3503) );
  MUX2_X1 U14994 ( .A(P3_DATAO_REG_11__SCAN_IN), .B(n12629), .S(n15577), .Z(
        P3_U3502) );
  MUX2_X1 U14995 ( .A(P3_DATAO_REG_10__SCAN_IN), .B(n12630), .S(n15577), .Z(
        P3_U3501) );
  MUX2_X1 U14996 ( .A(P3_DATAO_REG_9__SCAN_IN), .B(n12631), .S(n15577), .Z(
        P3_U3500) );
  MUX2_X1 U14997 ( .A(P3_DATAO_REG_8__SCAN_IN), .B(n12632), .S(n15577), .Z(
        P3_U3499) );
  MUX2_X1 U14998 ( .A(P3_DATAO_REG_7__SCAN_IN), .B(n12633), .S(n15577), .Z(
        P3_U3498) );
  MUX2_X1 U14999 ( .A(P3_DATAO_REG_6__SCAN_IN), .B(n12634), .S(P3_U3897), .Z(
        P3_U3497) );
  MUX2_X1 U15000 ( .A(P3_DATAO_REG_5__SCAN_IN), .B(n12635), .S(n15577), .Z(
        P3_U3496) );
  MUX2_X1 U15001 ( .A(P3_DATAO_REG_4__SCAN_IN), .B(n12636), .S(n15577), .Z(
        P3_U3495) );
  MUX2_X1 U15002 ( .A(P3_DATAO_REG_2__SCAN_IN), .B(n12637), .S(n15577), .Z(
        P3_U3493) );
  MUX2_X1 U15003 ( .A(P3_DATAO_REG_0__SCAN_IN), .B(n12638), .S(n15577), .Z(
        P3_U3491) );
  XNOR2_X1 U15004 ( .A(n12706), .B(P3_REG1_REG_19__SCAN_IN), .ZN(n12672) );
  INV_X1 U15005 ( .A(n15073), .ZN(n14948) );
  AOI22_X1 U15006 ( .A1(P3_REG1_REG_18__SCAN_IN), .A2(n14948), .B1(n15073), 
        .B2(n13425), .ZN(n15076) );
  NAND2_X1 U15007 ( .A1(P3_REG1_REG_16__SCAN_IN), .A2(n12674), .ZN(n12651) );
  AOI22_X1 U15008 ( .A1(P3_REG1_REG_16__SCAN_IN), .A2(n12674), .B1(n15042), 
        .B2(n12972), .ZN(n15050) );
  NAND2_X1 U15009 ( .A1(n15676), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n12690) );
  INV_X1 U15010 ( .A(n15676), .ZN(n12641) );
  INV_X1 U15011 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n12640) );
  INV_X1 U15012 ( .A(n12690), .ZN(n12639) );
  AOI21_X1 U15013 ( .B1(n12641), .B2(n12640), .A(n12639), .ZN(n15671) );
  NAND2_X1 U15014 ( .A1(P3_REG1_REG_12__SCAN_IN), .A2(n15640), .ZN(n12646) );
  INV_X1 U15015 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n12980) );
  AOI22_X1 U15016 ( .A1(P3_REG1_REG_12__SCAN_IN), .A2(n15640), .B1(n12685), 
        .B2(n12980), .ZN(n15636) );
  NAND2_X1 U15017 ( .A1(P3_REG1_REG_10__SCAN_IN), .A2(n12655), .ZN(n12643) );
  NAND2_X1 U15018 ( .A1(n15622), .A2(n12644), .ZN(n12645) );
  NAND2_X1 U15019 ( .A1(P3_REG1_REG_11__SCAN_IN), .A2(n15618), .ZN(n15617) );
  NAND2_X1 U15020 ( .A1(n12645), .A2(n15617), .ZN(n15635) );
  NAND2_X1 U15021 ( .A1(n15636), .A2(n15635), .ZN(n15634) );
  NAND2_X1 U15022 ( .A1(n12646), .A2(n15634), .ZN(n12647) );
  NAND2_X1 U15023 ( .A1(n15655), .A2(n12647), .ZN(n12648) );
  INV_X1 U15024 ( .A(n15655), .ZN(n12688) );
  XNOR2_X1 U15025 ( .A(n12688), .B(n12647), .ZN(n15652) );
  NAND2_X1 U15026 ( .A1(P3_REG1_REG_13__SCAN_IN), .A2(n15652), .ZN(n15651) );
  NAND2_X1 U15027 ( .A1(n12648), .A2(n15651), .ZN(n15670) );
  NAND2_X1 U15028 ( .A1(n15671), .A2(n15670), .ZN(n15669) );
  NAND2_X1 U15029 ( .A1(n15032), .A2(n12649), .ZN(n12650) );
  NAND2_X1 U15030 ( .A1(P3_REG1_REG_15__SCAN_IN), .A2(n15029), .ZN(n15028) );
  NAND2_X1 U15031 ( .A1(n12650), .A2(n15028), .ZN(n15049) );
  NAND2_X1 U15032 ( .A1(n12699), .A2(n12652), .ZN(n12653) );
  XNOR2_X1 U15033 ( .A(n7689), .B(n12652), .ZN(n15060) );
  NAND2_X1 U15034 ( .A1(P3_REG1_REG_17__SCAN_IN), .A2(n15060), .ZN(n15059) );
  NAND2_X1 U15035 ( .A1(n15076), .A2(n15075), .ZN(n15074) );
  NAND2_X1 U15036 ( .A1(n15676), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n12691) );
  NOR2_X1 U15037 ( .A1(n12682), .A2(n12656), .ZN(n12657) );
  NAND2_X1 U15038 ( .A1(P3_REG2_REG_12__SCAN_IN), .A2(n15640), .ZN(n12658) );
  OAI21_X1 U15039 ( .B1(P3_REG2_REG_12__SCAN_IN), .B2(n15640), .A(n12658), 
        .ZN(n15633) );
  OR2_X1 U15040 ( .A1(n15676), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n12660) );
  NAND2_X1 U15041 ( .A1(n12691), .A2(n12660), .ZN(n15667) );
  AND2_X1 U15042 ( .A1(n15032), .A2(n12661), .ZN(n12662) );
  AOI22_X1 U15043 ( .A1(P3_REG2_REG_16__SCAN_IN), .A2(n15042), .B1(n12674), 
        .B2(n13407), .ZN(n15053) );
  NOR2_X1 U15044 ( .A1(n7689), .A2(n12663), .ZN(n12664) );
  INV_X1 U15045 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n15067) );
  INV_X1 U15046 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n12665) );
  AOI22_X1 U15047 ( .A1(P3_REG2_REG_18__SCAN_IN), .A2(n15073), .B1(n14948), 
        .B2(n12665), .ZN(n15083) );
  XNOR2_X1 U15048 ( .A(n12666), .B(P3_REG2_REG_19__SCAN_IN), .ZN(n12671) );
  XNOR2_X1 U15049 ( .A(n12667), .B(n12671), .ZN(n12668) );
  NAND2_X1 U15050 ( .A1(n12668), .A2(n15082), .ZN(n12708) );
  NAND2_X1 U15051 ( .A1(P3_REG3_REG_19__SCAN_IN), .A2(P3_U3151), .ZN(n12669)
         );
  OAI21_X1 U15052 ( .B1(n15613), .B2(n12670), .A(n12669), .ZN(n12705) );
  INV_X1 U15053 ( .A(n12671), .ZN(n12673) );
  MUX2_X1 U15054 ( .A(n12673), .B(n12672), .S(n12696), .Z(n12704) );
  MUX2_X1 U15055 ( .A(n12665), .B(n13425), .S(n12696), .Z(n15078) );
  MUX2_X1 U15056 ( .A(P3_REG2_REG_17__SCAN_IN), .B(P3_REG1_REG_17__SCAN_IN), 
        .S(n12694), .Z(n12700) );
  AND2_X1 U15057 ( .A1(n12700), .A2(n12699), .ZN(n12701) );
  MUX2_X1 U15058 ( .A(P3_REG2_REG_16__SCAN_IN), .B(P3_REG1_REG_16__SCAN_IN), 
        .S(n12694), .Z(n12675) );
  AND2_X1 U15059 ( .A1(n12675), .A2(n12674), .ZN(n15043) );
  MUX2_X1 U15060 ( .A(P3_REG2_REG_13__SCAN_IN), .B(P3_REG1_REG_13__SCAN_IN), 
        .S(n12696), .Z(n12686) );
  INV_X1 U15061 ( .A(n12686), .ZN(n12687) );
  MUX2_X1 U15062 ( .A(P3_REG2_REG_12__SCAN_IN), .B(P3_REG1_REG_12__SCAN_IN), 
        .S(n12696), .Z(n12683) );
  INV_X1 U15063 ( .A(n12683), .ZN(n12684) );
  MUX2_X1 U15064 ( .A(P3_REG2_REG_11__SCAN_IN), .B(P3_REG1_REG_11__SCAN_IN), 
        .S(n12696), .Z(n12680) );
  INV_X1 U15065 ( .A(n12680), .ZN(n12681) );
  INV_X1 U15066 ( .A(n12676), .ZN(n12678) );
  XNOR2_X1 U15067 ( .A(n12680), .B(n15622), .ZN(n15626) );
  NOR2_X1 U15068 ( .A1(n15627), .A2(n15626), .ZN(n15625) );
  AOI21_X1 U15069 ( .B1(n12682), .B2(n12681), .A(n15625), .ZN(n15645) );
  XNOR2_X1 U15070 ( .A(n12683), .B(n12685), .ZN(n15644) );
  NAND2_X1 U15071 ( .A1(n15645), .A2(n15644), .ZN(n15643) );
  OAI21_X1 U15072 ( .B1(n12685), .B2(n12684), .A(n15643), .ZN(n15659) );
  XNOR2_X1 U15073 ( .A(n12686), .B(n15655), .ZN(n15660) );
  NOR2_X1 U15074 ( .A1(n15659), .A2(n15660), .ZN(n15658) );
  AOI21_X1 U15075 ( .B1(n12688), .B2(n12687), .A(n15658), .ZN(n15684) );
  INV_X1 U15076 ( .A(n15667), .ZN(n12689) );
  MUX2_X1 U15077 ( .A(n12689), .B(n15671), .S(n12696), .Z(n15683) );
  NAND2_X1 U15078 ( .A1(n15684), .A2(n15683), .ZN(n15682) );
  MUX2_X1 U15079 ( .A(n12691), .B(n12690), .S(n12696), .Z(n12692) );
  NAND2_X1 U15080 ( .A1(n15682), .A2(n12692), .ZN(n12693) );
  MUX2_X1 U15081 ( .A(P3_REG2_REG_15__SCAN_IN), .B(P3_REG1_REG_15__SCAN_IN), 
        .S(n12694), .Z(n15037) );
  NOR2_X1 U15082 ( .A1(n12695), .A2(n15035), .ZN(n15047) );
  MUX2_X1 U15083 ( .A(n13407), .B(n12972), .S(n12696), .Z(n12697) );
  NAND2_X1 U15084 ( .A1(n12697), .A2(n15042), .ZN(n15045) );
  INV_X1 U15085 ( .A(n12701), .ZN(n12698) );
  OAI21_X1 U15086 ( .B1(n12700), .B2(n12699), .A(n12698), .ZN(n15062) );
  NAND2_X1 U15087 ( .A1(n15078), .A2(n15079), .ZN(n15077) );
  NAND2_X1 U15088 ( .A1(n15073), .A2(n12702), .ZN(n12703) );
  OAI211_X1 U15089 ( .C1(n12710), .C2(n12709), .A(n12708), .B(n12707), .ZN(
        P3_U3201) );
  INV_X1 U15090 ( .A(n12711), .ZN(n12712) );
  NOR2_X1 U15091 ( .A1(n12713), .A2(n12712), .ZN(n15101) );
  INV_X1 U15092 ( .A(n12714), .ZN(n12715) );
  AOI21_X1 U15093 ( .B1(n15101), .B2(n15719), .A(n12715), .ZN(n15090) );
  NAND2_X1 U15094 ( .A1(n15703), .A2(P3_REG2_REG_31__SCAN_IN), .ZN(n12716) );
  OAI211_X1 U15095 ( .C1(n12990), .C2(n12898), .A(n15090), .B(n12716), .ZN(
        P3_U3202) );
  NAND2_X1 U15096 ( .A1(n12717), .A2(n12728), .ZN(n12718) );
  NAND2_X1 U15097 ( .A1(n12718), .A2(n15695), .ZN(n12720) );
  OR2_X1 U15098 ( .A1(n12720), .A2(n12719), .ZN(n12724) );
  AOI22_X1 U15099 ( .A1(n12867), .A2(n12722), .B1(n12721), .B2(n12869), .ZN(
        n12723) );
  NAND2_X1 U15100 ( .A1(n12724), .A2(n12723), .ZN(n12923) );
  INV_X1 U15101 ( .A(n12923), .ZN(n12734) );
  INV_X1 U15102 ( .A(n12725), .ZN(n12726) );
  OR2_X1 U15103 ( .A1(n12727), .A2(n12726), .ZN(n12729) );
  XNOR2_X1 U15104 ( .A(n12729), .B(n12728), .ZN(n12921) );
  AOI22_X1 U15105 ( .A1(n15703), .A2(P3_REG2_REG_28__SCAN_IN), .B1(n12911), 
        .B2(n12730), .ZN(n12731) );
  OAI21_X1 U15106 ( .B1(n12993), .B2(n12898), .A(n12731), .ZN(n12732) );
  AOI21_X1 U15107 ( .B1(n12921), .B2(n15098), .A(n12732), .ZN(n12733) );
  OAI21_X1 U15108 ( .B1(n12734), .B2(n15703), .A(n12733), .ZN(P3_U3205) );
  NAND2_X1 U15109 ( .A1(n12735), .A2(n12736), .ZN(n12737) );
  NAND2_X1 U15110 ( .A1(n12737), .A2(n12740), .ZN(n12739) );
  INV_X1 U15111 ( .A(n12931), .ZN(n12750) );
  XNOR2_X1 U15112 ( .A(n12741), .B(n12740), .ZN(n12743) );
  OAI21_X1 U15113 ( .B1(n12743), .B2(n15708), .A(n12742), .ZN(n12930) );
  NAND2_X1 U15114 ( .A1(n12930), .A2(n15719), .ZN(n12749) );
  INV_X1 U15115 ( .A(P3_REG2_REG_26__SCAN_IN), .ZN(n12745) );
  OAI22_X1 U15116 ( .A1(n15719), .A2(n12745), .B1(n12744), .B2(n15711), .ZN(
        n12746) );
  AOI21_X1 U15117 ( .B1(n12747), .B2(n15097), .A(n12746), .ZN(n12748) );
  OAI211_X1 U15118 ( .C1(n12750), .C2(n12827), .A(n12749), .B(n12748), .ZN(
        P3_U3207) );
  AND2_X1 U15119 ( .A1(n12764), .A2(n12751), .ZN(n12754) );
  OAI211_X1 U15120 ( .C1(n12754), .C2(n12753), .A(n12752), .B(n15695), .ZN(
        n12756) );
  AND2_X1 U15121 ( .A1(n12756), .A2(n12755), .ZN(n12936) );
  OR2_X1 U15122 ( .A1(n12758), .A2(n12757), .ZN(n12759) );
  NAND2_X1 U15123 ( .A1(n12735), .A2(n12759), .ZN(n12934) );
  AOI22_X1 U15124 ( .A1(n15703), .A2(P3_REG2_REG_25__SCAN_IN), .B1(n12911), 
        .B2(n12760), .ZN(n12761) );
  OAI21_X1 U15125 ( .B1(n13003), .B2(n12898), .A(n12761), .ZN(n12762) );
  AOI21_X1 U15126 ( .B1(n12934), .B2(n15098), .A(n12762), .ZN(n12763) );
  OAI21_X1 U15127 ( .B1(n12936), .B2(n15703), .A(n12763), .ZN(P3_U3208) );
  INV_X1 U15128 ( .A(n12764), .ZN(n12765) );
  AOI21_X1 U15129 ( .B1(n7853), .B2(n12766), .A(n12765), .ZN(n12768) );
  OAI21_X1 U15130 ( .B1(n12768), .B2(n15708), .A(n12767), .ZN(n12938) );
  INV_X1 U15131 ( .A(n12938), .ZN(n12778) );
  INV_X1 U15132 ( .A(n12779), .ZN(n12771) );
  OAI21_X1 U15133 ( .B1(n12771), .B2(n12770), .A(n12769), .ZN(n12773) );
  NAND2_X1 U15134 ( .A1(n12773), .A2(n12772), .ZN(n12939) );
  AOI22_X1 U15135 ( .A1(n15703), .A2(P3_REG2_REG_24__SCAN_IN), .B1(n12911), 
        .B2(n12774), .ZN(n12775) );
  OAI21_X1 U15136 ( .B1(n6986), .B2(n12898), .A(n12775), .ZN(n12776) );
  AOI21_X1 U15137 ( .B1(n12939), .B2(n15098), .A(n12776), .ZN(n12777) );
  OAI21_X1 U15138 ( .B1(n12778), .B2(n15703), .A(n12777), .ZN(P3_U3209) );
  OAI21_X1 U15139 ( .B1(n12780), .B2(n12782), .A(n12779), .ZN(n12788) );
  INV_X1 U15140 ( .A(n12781), .ZN(n12785) );
  INV_X1 U15141 ( .A(n12782), .ZN(n12784) );
  OAI211_X1 U15142 ( .C1(n12785), .C2(n12784), .A(n12783), .B(n15695), .ZN(
        n12787) );
  OAI211_X1 U15143 ( .C1(n15766), .C2(n12788), .A(n12787), .B(n12786), .ZN(
        n12942) );
  INV_X1 U15144 ( .A(n12942), .ZN(n12793) );
  INV_X1 U15145 ( .A(n12788), .ZN(n12943) );
  AOI22_X1 U15146 ( .A1(n15703), .A2(P3_REG2_REG_23__SCAN_IN), .B1(n12789), 
        .B2(n12911), .ZN(n12790) );
  OAI21_X1 U15147 ( .B1(n13010), .B2(n12898), .A(n12790), .ZN(n12791) );
  AOI21_X1 U15148 ( .B1(n12943), .B2(n15716), .A(n12791), .ZN(n12792) );
  OAI21_X1 U15149 ( .B1(n12793), .B2(n15703), .A(n12792), .ZN(P3_U3210) );
  XNOR2_X1 U15150 ( .A(n12795), .B(n12794), .ZN(n12797) );
  OAI21_X1 U15151 ( .B1(n12797), .B2(n15708), .A(n12796), .ZN(n12946) );
  INV_X1 U15152 ( .A(n12946), .ZN(n12804) );
  XNOR2_X1 U15153 ( .A(n12799), .B(n12798), .ZN(n12947) );
  AOI22_X1 U15154 ( .A1(n15703), .A2(P3_REG2_REG_22__SCAN_IN), .B1(n12911), 
        .B2(n12800), .ZN(n12801) );
  OAI21_X1 U15155 ( .B1(n13014), .B2(n12898), .A(n12801), .ZN(n12802) );
  AOI21_X1 U15156 ( .B1(n12947), .B2(n15098), .A(n12802), .ZN(n12803) );
  OAI21_X1 U15157 ( .B1(n12804), .B2(n15703), .A(n12803), .ZN(P3_U3211) );
  XOR2_X1 U15158 ( .A(n12805), .B(n12808), .Z(n12807) );
  OAI21_X1 U15159 ( .B1(n12807), .B2(n15708), .A(n12806), .ZN(n12950) );
  INV_X1 U15160 ( .A(n12950), .ZN(n12815) );
  XOR2_X1 U15161 ( .A(n12809), .B(n12808), .Z(n12951) );
  NOR2_X1 U15162 ( .A1(n13018), .A2(n12898), .ZN(n12813) );
  OAI22_X1 U15163 ( .A1(n15719), .A2(n12811), .B1(n12810), .B2(n15711), .ZN(
        n12812) );
  AOI211_X1 U15164 ( .C1(n12951), .C2(n15098), .A(n12813), .B(n12812), .ZN(
        n12814) );
  OAI21_X1 U15165 ( .B1(n12815), .B2(n15703), .A(n12814), .ZN(P3_U3212) );
  NAND2_X1 U15166 ( .A1(n12816), .A2(n12825), .ZN(n12817) );
  NAND3_X1 U15167 ( .A1(n12818), .A2(n15695), .A3(n12817), .ZN(n12820) );
  INV_X1 U15168 ( .A(P3_REG2_REG_20__SCAN_IN), .ZN(n12822) );
  OAI22_X1 U15169 ( .A1(n15719), .A2(n12822), .B1(n12821), .B2(n15711), .ZN(
        n12823) );
  AOI21_X1 U15170 ( .B1(n12954), .B2(n15097), .A(n12823), .ZN(n12829) );
  OAI21_X1 U15171 ( .B1(n12826), .B2(n12825), .A(n12824), .ZN(n12955) );
  OR2_X1 U15172 ( .A1(n12955), .A2(n12827), .ZN(n12828) );
  OAI211_X1 U15173 ( .C1(n12957), .C2(n15703), .A(n12829), .B(n12828), .ZN(
        P3_U3213) );
  XOR2_X1 U15174 ( .A(n12833), .B(n12830), .Z(n12832) );
  OAI21_X1 U15175 ( .B1(n12832), .B2(n15708), .A(n12831), .ZN(n12959) );
  INV_X1 U15176 ( .A(n12959), .ZN(n12839) );
  XNOR2_X1 U15177 ( .A(n12834), .B(n12833), .ZN(n12960) );
  AOI22_X1 U15178 ( .A1(n15703), .A2(P3_REG2_REG_19__SCAN_IN), .B1(n12911), 
        .B2(n12835), .ZN(n12836) );
  OAI21_X1 U15179 ( .B1(n13025), .B2(n12898), .A(n12836), .ZN(n12837) );
  AOI21_X1 U15180 ( .B1(n12960), .B2(n15098), .A(n12837), .ZN(n12838) );
  OAI21_X1 U15181 ( .B1(n12839), .B2(n15703), .A(n12838), .ZN(P3_U3214) );
  INV_X1 U15182 ( .A(n12840), .ZN(n12841) );
  AOI21_X1 U15183 ( .B1(n12846), .B2(n12842), .A(n12841), .ZN(n12843) );
  OAI222_X1 U15184 ( .A1(n15017), .A2(n12845), .B1(n15019), .B2(n12844), .C1(
        n15708), .C2(n12843), .ZN(n12963) );
  INV_X1 U15185 ( .A(n12963), .ZN(n12852) );
  XNOR2_X1 U15186 ( .A(n12847), .B(n12846), .ZN(n12964) );
  AOI22_X1 U15187 ( .A1(n15703), .A2(P3_REG2_REG_18__SCAN_IN), .B1(n12911), 
        .B2(n12848), .ZN(n12849) );
  OAI21_X1 U15188 ( .B1(n13029), .B2(n12898), .A(n12849), .ZN(n12850) );
  AOI21_X1 U15189 ( .B1(n12964), .B2(n15098), .A(n12850), .ZN(n12851) );
  OAI21_X1 U15190 ( .B1(n12852), .B2(n15703), .A(n12851), .ZN(P3_U3215) );
  XNOR2_X1 U15191 ( .A(n12853), .B(n12854), .ZN(n12855) );
  OAI222_X1 U15192 ( .A1(n15017), .A2(n12857), .B1(n15019), .B2(n12856), .C1(
        n12855), .C2(n15708), .ZN(n12966) );
  INV_X1 U15193 ( .A(n12966), .ZN(n12865) );
  OAI21_X1 U15194 ( .B1(n12860), .B2(n12859), .A(n12858), .ZN(n12967) );
  NOR2_X1 U15195 ( .A1(n13032), .A2(n12898), .ZN(n12863) );
  OAI22_X1 U15196 ( .A1(n15719), .A2(n15067), .B1(n12861), .B2(n15711), .ZN(
        n12862) );
  AOI211_X1 U15197 ( .C1(n12967), .C2(n15098), .A(n12863), .B(n12862), .ZN(
        n12864) );
  OAI21_X1 U15198 ( .B1(n12865), .B2(n15703), .A(n12864), .ZN(P3_U3216) );
  XNOR2_X1 U15199 ( .A(n12866), .B(n12874), .ZN(n12873) );
  NAND2_X1 U15200 ( .A1(n12868), .A2(n12867), .ZN(n12872) );
  NAND2_X1 U15201 ( .A1(n12870), .A2(n12869), .ZN(n12871) );
  AND2_X1 U15202 ( .A1(n12872), .A2(n12871), .ZN(n15010) );
  OAI21_X1 U15203 ( .B1(n12873), .B2(n15708), .A(n15010), .ZN(n12970) );
  INV_X1 U15204 ( .A(n12970), .ZN(n12879) );
  XNOR2_X1 U15205 ( .A(n12875), .B(n12874), .ZN(n12971) );
  AOI22_X1 U15206 ( .A1(n15703), .A2(P3_REG2_REG_16__SCAN_IN), .B1(n12911), 
        .B2(n15001), .ZN(n12876) );
  OAI21_X1 U15207 ( .B1(n13036), .B2(n12898), .A(n12876), .ZN(n12877) );
  AOI21_X1 U15208 ( .B1(n12971), .B2(n15098), .A(n12877), .ZN(n12878) );
  OAI21_X1 U15209 ( .B1(n12879), .B2(n15703), .A(n12878), .ZN(P3_U3217) );
  XNOR2_X1 U15210 ( .A(n12881), .B(n12880), .ZN(n12883) );
  OAI21_X1 U15211 ( .B1(n12883), .B2(n15708), .A(n12882), .ZN(n12974) );
  INV_X1 U15212 ( .A(n12974), .ZN(n12890) );
  XNOR2_X1 U15213 ( .A(n12885), .B(n12884), .ZN(n12975) );
  AOI22_X1 U15214 ( .A1(n15703), .A2(P3_REG2_REG_15__SCAN_IN), .B1(n12911), 
        .B2(n12886), .ZN(n12887) );
  OAI21_X1 U15215 ( .B1(n13040), .B2(n12898), .A(n12887), .ZN(n12888) );
  AOI21_X1 U15216 ( .B1(n12975), .B2(n15098), .A(n12888), .ZN(n12889) );
  OAI21_X1 U15217 ( .B1(n12890), .B2(n15703), .A(n12889), .ZN(P3_U3218) );
  XNOR2_X1 U15218 ( .A(n12891), .B(n12894), .ZN(n12893) );
  OAI21_X1 U15219 ( .B1(n12893), .B2(n15708), .A(n12892), .ZN(n15109) );
  INV_X1 U15220 ( .A(n15109), .ZN(n12901) );
  XNOR2_X1 U15221 ( .A(n12895), .B(n12894), .ZN(n15104) );
  AOI22_X1 U15222 ( .A1(n15703), .A2(P3_REG2_REG_14__SCAN_IN), .B1(n12911), 
        .B2(n12896), .ZN(n12897) );
  OAI21_X1 U15223 ( .B1(n15105), .B2(n12898), .A(n12897), .ZN(n12899) );
  AOI21_X1 U15224 ( .B1(n15104), .B2(n15098), .A(n12899), .ZN(n12900) );
  OAI21_X1 U15225 ( .B1(n12901), .B2(n15703), .A(n12900), .ZN(P3_U3219) );
  NAND3_X1 U15226 ( .A1(n11409), .A2(n12908), .A3(n12902), .ZN(n12903) );
  NAND3_X1 U15227 ( .A1(n12904), .A2(n15695), .A3(n12903), .ZN(n12906) );
  NAND2_X1 U15228 ( .A1(n12906), .A2(n12905), .ZN(n12978) );
  INV_X1 U15229 ( .A(n12978), .ZN(n12917) );
  OAI21_X1 U15230 ( .B1(n12909), .B2(n12908), .A(n12907), .ZN(n12979) );
  INV_X1 U15231 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n12914) );
  AOI22_X1 U15232 ( .A1(n15097), .A2(n12912), .B1(n12911), .B2(n12910), .ZN(
        n12913) );
  OAI21_X1 U15233 ( .B1(n12914), .B2(n15719), .A(n12913), .ZN(n12915) );
  AOI21_X1 U15234 ( .B1(n12979), .B2(n15098), .A(n12915), .ZN(n12916) );
  OAI21_X1 U15235 ( .B1(n12917), .B2(n15703), .A(n12916), .ZN(P3_U3221) );
  INV_X1 U15236 ( .A(P3_REG1_REG_31__SCAN_IN), .ZN(n12918) );
  NOR2_X1 U15237 ( .A1(n15788), .A2(n12918), .ZN(n12919) );
  AOI21_X1 U15238 ( .B1(n15101), .B2(n15788), .A(n12919), .ZN(n12920) );
  OAI21_X1 U15239 ( .B1(n12990), .B2(n12986), .A(n12920), .ZN(P3_U3490) );
  INV_X1 U15240 ( .A(P3_REG1_REG_28__SCAN_IN), .ZN(n12924) );
  AND2_X1 U15241 ( .A1(n12921), .A2(n15746), .ZN(n12922) );
  NOR2_X1 U15242 ( .A1(n12923), .A2(n12922), .ZN(n12991) );
  INV_X1 U15243 ( .A(n15765), .ZN(n15750) );
  NAND2_X1 U15244 ( .A1(n12925), .A2(n15750), .ZN(n12926) );
  MUX2_X1 U15245 ( .A(P3_REG1_REG_27__SCAN_IN), .B(n12994), .S(n15788), .Z(
        n12928) );
  INV_X1 U15246 ( .A(n12928), .ZN(n12929) );
  OAI21_X1 U15247 ( .B1(n12996), .B2(n12986), .A(n12929), .ZN(P3_U3486) );
  INV_X1 U15248 ( .A(P3_REG1_REG_26__SCAN_IN), .ZN(n12932) );
  AOI21_X1 U15249 ( .B1(n12931), .B2(n15746), .A(n12930), .ZN(n12997) );
  MUX2_X1 U15250 ( .A(n12932), .B(n12997), .S(n15788), .Z(n12933) );
  OAI21_X1 U15251 ( .B1(n12999), .B2(n12986), .A(n12933), .ZN(P3_U3485) );
  NAND2_X1 U15252 ( .A1(n12934), .A2(n15746), .ZN(n12935) );
  AND2_X1 U15253 ( .A1(n12936), .A2(n12935), .ZN(n13001) );
  MUX2_X1 U15254 ( .A(n13001), .B(n13229), .S(n15786), .Z(n12937) );
  OAI21_X1 U15255 ( .B1(n13003), .B2(n12986), .A(n12937), .ZN(P3_U3484) );
  INV_X1 U15256 ( .A(P3_REG1_REG_24__SCAN_IN), .ZN(n12940) );
  AOI21_X1 U15257 ( .B1(n15746), .B2(n12939), .A(n12938), .ZN(n13004) );
  MUX2_X1 U15258 ( .A(n12940), .B(n13004), .S(n15788), .Z(n12941) );
  OAI21_X1 U15259 ( .B1(n6986), .B2(n12986), .A(n12941), .ZN(P3_U3483) );
  INV_X1 U15260 ( .A(P3_REG1_REG_23__SCAN_IN), .ZN(n12944) );
  AOI21_X1 U15261 ( .B1(n15750), .B2(n12943), .A(n12942), .ZN(n13007) );
  MUX2_X1 U15262 ( .A(n12944), .B(n13007), .S(n15788), .Z(n12945) );
  OAI21_X1 U15263 ( .B1(n13010), .B2(n12986), .A(n12945), .ZN(P3_U3482) );
  INV_X1 U15264 ( .A(P3_REG1_REG_22__SCAN_IN), .ZN(n12948) );
  AOI21_X1 U15265 ( .B1(n15746), .B2(n12947), .A(n12946), .ZN(n13011) );
  MUX2_X1 U15266 ( .A(n12948), .B(n13011), .S(n15788), .Z(n12949) );
  OAI21_X1 U15267 ( .B1(n13014), .B2(n12986), .A(n12949), .ZN(P3_U3481) );
  INV_X1 U15268 ( .A(P3_REG1_REG_21__SCAN_IN), .ZN(n12952) );
  AOI21_X1 U15269 ( .B1(n12951), .B2(n15746), .A(n12950), .ZN(n13015) );
  MUX2_X1 U15270 ( .A(n12952), .B(n13015), .S(n15788), .Z(n12953) );
  OAI21_X1 U15271 ( .B1(n13018), .B2(n12986), .A(n12953), .ZN(P3_U3480) );
  INV_X1 U15272 ( .A(n12954), .ZN(n13022) );
  OR2_X1 U15273 ( .A1(n12955), .A2(n15106), .ZN(n12956) );
  MUX2_X1 U15274 ( .A(n13020), .B(n13219), .S(n15786), .Z(n12958) );
  OAI21_X1 U15275 ( .B1(n13022), .B2(n12986), .A(n12958), .ZN(P3_U3479) );
  INV_X1 U15276 ( .A(P3_REG1_REG_19__SCAN_IN), .ZN(n12961) );
  AOI21_X1 U15277 ( .B1(n12960), .B2(n15746), .A(n12959), .ZN(n13023) );
  MUX2_X1 U15278 ( .A(n12961), .B(n13023), .S(n15788), .Z(n12962) );
  OAI21_X1 U15279 ( .B1(n13025), .B2(n12986), .A(n12962), .ZN(P3_U3478) );
  AOI21_X1 U15280 ( .B1(n12964), .B2(n15746), .A(n12963), .ZN(n13026) );
  MUX2_X1 U15281 ( .A(n13425), .B(n13026), .S(n15788), .Z(n12965) );
  OAI21_X1 U15282 ( .B1(n13029), .B2(n12986), .A(n12965), .ZN(P3_U3477) );
  INV_X1 U15283 ( .A(P3_REG1_REG_17__SCAN_IN), .ZN(n12968) );
  AOI21_X1 U15284 ( .B1(n15746), .B2(n12967), .A(n12966), .ZN(n13030) );
  MUX2_X1 U15285 ( .A(n12968), .B(n13030), .S(n15788), .Z(n12969) );
  OAI21_X1 U15286 ( .B1(n12986), .B2(n13032), .A(n12969), .ZN(P3_U3476) );
  AOI21_X1 U15287 ( .B1(n12971), .B2(n15746), .A(n12970), .ZN(n13033) );
  MUX2_X1 U15288 ( .A(n12972), .B(n13033), .S(n15788), .Z(n12973) );
  OAI21_X1 U15289 ( .B1(n13036), .B2(n12986), .A(n12973), .ZN(P3_U3475) );
  AOI21_X1 U15290 ( .B1(n12975), .B2(n15746), .A(n12974), .ZN(n13037) );
  MUX2_X1 U15291 ( .A(n12976), .B(n13037), .S(n15788), .Z(n12977) );
  OAI21_X1 U15292 ( .B1(n12986), .B2(n13040), .A(n12977), .ZN(P3_U3474) );
  AOI21_X1 U15293 ( .B1(n15746), .B2(n12979), .A(n12978), .ZN(n13041) );
  MUX2_X1 U15294 ( .A(n12980), .B(n13041), .S(n15788), .Z(n12981) );
  OAI21_X1 U15295 ( .B1(n13044), .B2(n12986), .A(n12981), .ZN(P3_U3471) );
  INV_X1 U15296 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n12984) );
  AOI21_X1 U15297 ( .B1(n15746), .B2(n12983), .A(n12982), .ZN(n13045) );
  MUX2_X1 U15298 ( .A(n12984), .B(n13045), .S(n15788), .Z(n12985) );
  OAI21_X1 U15299 ( .B1(n12986), .B2(n13048), .A(n12985), .ZN(P3_U3470) );
  INV_X1 U15300 ( .A(P3_REG0_REG_31__SCAN_IN), .ZN(n12987) );
  NOR2_X1 U15301 ( .A1(n15773), .A2(n12987), .ZN(n12988) );
  AOI21_X1 U15302 ( .B1(n15101), .B2(n15773), .A(n12988), .ZN(n12989) );
  OAI21_X1 U15303 ( .B1(n12990), .B2(n13049), .A(n12989), .ZN(P3_U3458) );
  INV_X1 U15304 ( .A(P3_REG0_REG_28__SCAN_IN), .ZN(n12992) );
  OAI21_X1 U15305 ( .B1(n12996), .B2(n13049), .A(n12995), .ZN(P3_U3454) );
  MUX2_X1 U15306 ( .A(n13428), .B(n12997), .S(n15773), .Z(n12998) );
  OAI21_X1 U15307 ( .B1(n12999), .B2(n13049), .A(n12998), .ZN(P3_U3453) );
  MUX2_X1 U15308 ( .A(n13001), .B(n13000), .S(n15771), .Z(n13002) );
  OAI21_X1 U15309 ( .B1(n13003), .B2(n13049), .A(n13002), .ZN(P3_U3452) );
  MUX2_X1 U15310 ( .A(n13005), .B(n13004), .S(n15773), .Z(n13006) );
  OAI21_X1 U15311 ( .B1(n6986), .B2(n13049), .A(n13006), .ZN(P3_U3451) );
  INV_X1 U15312 ( .A(P3_REG0_REG_23__SCAN_IN), .ZN(n13008) );
  MUX2_X1 U15313 ( .A(n13008), .B(n13007), .S(n15773), .Z(n13009) );
  OAI21_X1 U15314 ( .B1(n13010), .B2(n13049), .A(n13009), .ZN(P3_U3450) );
  INV_X1 U15315 ( .A(P3_REG0_REG_22__SCAN_IN), .ZN(n13012) );
  MUX2_X1 U15316 ( .A(n13012), .B(n13011), .S(n15773), .Z(n13013) );
  OAI21_X1 U15317 ( .B1(n13014), .B2(n13049), .A(n13013), .ZN(P3_U3449) );
  MUX2_X1 U15318 ( .A(n13016), .B(n13015), .S(n15773), .Z(n13017) );
  OAI21_X1 U15319 ( .B1(n13018), .B2(n13049), .A(n13017), .ZN(P3_U3448) );
  MUX2_X1 U15320 ( .A(n13020), .B(n13019), .S(n15771), .Z(n13021) );
  OAI21_X1 U15321 ( .B1(n13022), .B2(n13049), .A(n13021), .ZN(P3_U3447) );
  MUX2_X1 U15322 ( .A(n13243), .B(n13023), .S(n15773), .Z(n13024) );
  OAI21_X1 U15323 ( .B1(n13025), .B2(n13049), .A(n13024), .ZN(P3_U3446) );
  MUX2_X1 U15324 ( .A(n13027), .B(n13026), .S(n15773), .Z(n13028) );
  OAI21_X1 U15325 ( .B1(n13029), .B2(n13049), .A(n13028), .ZN(P3_U3444) );
  MUX2_X1 U15326 ( .A(n13421), .B(n13030), .S(n15773), .Z(n13031) );
  OAI21_X1 U15327 ( .B1(n13049), .B2(n13032), .A(n13031), .ZN(P3_U3441) );
  INV_X1 U15328 ( .A(P3_REG0_REG_16__SCAN_IN), .ZN(n13034) );
  MUX2_X1 U15329 ( .A(n13034), .B(n13033), .S(n15773), .Z(n13035) );
  OAI21_X1 U15330 ( .B1(n13036), .B2(n13049), .A(n13035), .ZN(P3_U3438) );
  INV_X1 U15331 ( .A(P3_REG0_REG_15__SCAN_IN), .ZN(n13038) );
  MUX2_X1 U15332 ( .A(n13038), .B(n13037), .S(n15773), .Z(n13039) );
  OAI21_X1 U15333 ( .B1(n13049), .B2(n13040), .A(n13039), .ZN(P3_U3435) );
  INV_X1 U15334 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n13042) );
  MUX2_X1 U15335 ( .A(n13042), .B(n13041), .S(n15773), .Z(n13043) );
  OAI21_X1 U15336 ( .B1(n13044), .B2(n13049), .A(n13043), .ZN(P3_U3426) );
  INV_X1 U15337 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n13046) );
  MUX2_X1 U15338 ( .A(n13046), .B(n13045), .S(n15773), .Z(n13047) );
  OAI21_X1 U15339 ( .B1(n13049), .B2(n13048), .A(n13047), .ZN(P3_U3423) );
  MUX2_X1 U15340 ( .A(n13050), .B(P3_D_REG_1__SCAN_IN), .S(n13051), .Z(
        P3_U3377) );
  MUX2_X1 U15341 ( .A(n13052), .B(P3_D_REG_0__SCAN_IN), .S(n13051), .Z(
        P3_U3376) );
  NAND2_X1 U15342 ( .A1(n13053), .A2(n14945), .ZN(n13056) );
  OR4_X1 U15343 ( .A1(n7078), .A2(P3_IR_REG_30__SCAN_IN), .A3(n13054), .A4(
        P3_U3151), .ZN(n13055) );
  OAI211_X1 U15344 ( .C1(n13057), .C2(n14936), .A(n13056), .B(n13055), .ZN(
        P3_U3264) );
  OAI222_X1 U15345 ( .A1(n14936), .A2(n13329), .B1(P3_U3151), .B2(n13058), 
        .C1(n14938), .C2(n6797), .ZN(P3_U3266) );
  INV_X1 U15346 ( .A(n13059), .ZN(n13060) );
  OAI222_X1 U15347 ( .A1(n14936), .A2(n13061), .B1(n14938), .B2(n13060), .C1(
        n8427), .C2(P3_U3151), .ZN(P3_U3267) );
  XNOR2_X1 U15348 ( .A(n13942), .B(n13075), .ZN(n13066) );
  NAND2_X1 U15349 ( .A1(n13686), .A2(n11865), .ZN(n13084) );
  XNOR2_X1 U15350 ( .A(n13935), .B(n13107), .ZN(n13067) );
  NAND2_X1 U15351 ( .A1(n13660), .A2(n11865), .ZN(n13068) );
  XNOR2_X1 U15352 ( .A(n13067), .B(n13068), .ZN(n13525) );
  INV_X1 U15353 ( .A(n13068), .ZN(n13069) );
  XNOR2_X1 U15354 ( .A(n13927), .B(n13107), .ZN(n13073) );
  NAND2_X1 U15355 ( .A1(n13688), .A2(n11865), .ZN(n13071) );
  XNOR2_X1 U15356 ( .A(n13073), .B(n13071), .ZN(n13494) );
  INV_X1 U15357 ( .A(n13071), .ZN(n13072) );
  NAND2_X1 U15358 ( .A1(n13073), .A2(n13072), .ZN(n13074) );
  XNOR2_X1 U15359 ( .A(n13918), .B(n13075), .ZN(n13077) );
  NAND2_X1 U15360 ( .A1(n13663), .A2(n11865), .ZN(n13076) );
  NAND2_X1 U15361 ( .A1(n13077), .A2(n13076), .ZN(n13078) );
  OAI21_X1 U15362 ( .B1(n13077), .B2(n13076), .A(n13078), .ZN(n13553) );
  NAND2_X1 U15363 ( .A1(n13694), .A2(n11865), .ZN(n13103) );
  XNOR2_X1 U15364 ( .A(n13912), .B(n13107), .ZN(n13105) );
  XOR2_X1 U15365 ( .A(n13103), .B(n13105), .Z(n13100) );
  XNOR2_X1 U15366 ( .A(n13099), .B(n13100), .ZN(n13083) );
  AOI22_X1 U15367 ( .A1(n13702), .A2(n13555), .B1(n13701), .B2(n13663), .ZN(
        n13909) );
  INV_X1 U15368 ( .A(n13079), .ZN(n13733) );
  AOI22_X1 U15369 ( .A1(n13733), .A2(n13556), .B1(P2_REG3_REG_27__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13080) );
  OAI21_X1 U15370 ( .B1(n13909), .B2(n13558), .A(n13080), .ZN(n13081) );
  AOI21_X1 U15371 ( .B1(n13912), .B2(n15128), .A(n13081), .ZN(n13082) );
  OAI21_X1 U15372 ( .B1(n13083), .B2(n13561), .A(n13082), .ZN(P2_U3186) );
  XNOR2_X1 U15373 ( .A(n13085), .B(n13084), .ZN(n13089) );
  OAI22_X1 U15374 ( .A1(n13497), .A2(n13630), .B1(n13685), .B2(n13496), .ZN(
        n13941) );
  AOI22_X1 U15375 ( .A1(n13941), .A2(n15125), .B1(P2_REG3_REG_23__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13086) );
  OAI21_X1 U15376 ( .B1(n13786), .B2(n15131), .A(n13086), .ZN(n13087) );
  AOI21_X1 U15377 ( .B1(n13942), .B2(n15128), .A(n13087), .ZN(n13088) );
  OAI21_X1 U15378 ( .B1(n13089), .B2(n13561), .A(n13088), .ZN(P2_U3188) );
  OAI211_X1 U15379 ( .C1(n13092), .C2(n13091), .A(n13090), .B(n15123), .ZN(
        n13098) );
  AOI22_X1 U15380 ( .A1(n15128), .A2(n13094), .B1(n15125), .B2(n13093), .ZN(
        n13097) );
  MUX2_X1 U15381 ( .A(P2_STATE_REG_SCAN_IN), .B(n15131), .S(n13095), .Z(n13096) );
  NAND3_X1 U15382 ( .A1(n13098), .A2(n13097), .A3(n13096), .ZN(P2_U3190) );
  INV_X1 U15383 ( .A(n13099), .ZN(n13102) );
  INV_X1 U15384 ( .A(n13100), .ZN(n13101) );
  INV_X1 U15385 ( .A(n13103), .ZN(n13104) );
  NAND2_X1 U15386 ( .A1(n13105), .A2(n13104), .ZN(n13106) );
  NAND2_X1 U15387 ( .A1(n13702), .A2(n11865), .ZN(n13108) );
  XNOR2_X1 U15388 ( .A(n13108), .B(n13107), .ZN(n13111) );
  NOR3_X1 U15389 ( .A1(n13725), .A2(n13111), .A3(n15128), .ZN(n13109) );
  AOI21_X1 U15390 ( .B1(n13725), .B2(n13111), .A(n13109), .ZN(n13114) );
  NAND3_X1 U15391 ( .A1(n13905), .A2(n13542), .A3(n13111), .ZN(n13110) );
  OAI21_X1 U15392 ( .B1(n13905), .B2(n13111), .A(n13110), .ZN(n13112) );
  OAI21_X1 U15393 ( .B1(n13725), .B2(n13542), .A(n13561), .ZN(n13113) );
  AOI22_X1 U15394 ( .A1(n13722), .A2(n13556), .B1(P2_REG3_REG_28__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13116) );
  OAI22_X1 U15395 ( .A1(n13115), .A2(n13630), .B1(n13665), .B2(n13496), .ZN(
        n13715) );
  XNOR2_X1 U15396 ( .A(n6768), .B(n13117), .ZN(n13123) );
  AND2_X1 U15397 ( .A1(n13680), .A2(n13701), .ZN(n13118) );
  AOI21_X1 U15398 ( .B1(n13656), .B2(n13555), .A(n13118), .ZN(n13808) );
  OAI22_X1 U15399 ( .A1(n13808), .A2(n13558), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13119), .ZN(n13121) );
  INV_X1 U15400 ( .A(n13953), .ZN(n13815) );
  NOR2_X1 U15401 ( .A1(n13815), .A2(n13542), .ZN(n13120) );
  AOI211_X1 U15402 ( .C1(n13556), .C2(n13812), .A(n13121), .B(n13120), .ZN(
        n13122) );
  OAI21_X1 U15403 ( .B1(n13123), .B2(n13561), .A(n13122), .ZN(n13493) );
  AOI22_X1 U15404 ( .A1(P3_ADDR_REG_13__SCAN_IN), .A2(keyinput235), .B1(
        P2_D_REG_25__SCAN_IN), .B2(keyinput173), .ZN(n13124) );
  OAI221_X1 U15405 ( .B1(P3_ADDR_REG_13__SCAN_IN), .B2(keyinput235), .C1(
        P2_D_REG_25__SCAN_IN), .C2(keyinput173), .A(n13124), .ZN(n13131) );
  AOI22_X1 U15406 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(keyinput160), .B1(SI_27_), 
        .B2(keyinput130), .ZN(n13125) );
  OAI221_X1 U15407 ( .B1(P1_IR_REG_31__SCAN_IN), .B2(keyinput160), .C1(SI_27_), 
        .C2(keyinput130), .A(n13125), .ZN(n13130) );
  AOI22_X1 U15408 ( .A1(P3_REG3_REG_27__SCAN_IN), .A2(keyinput178), .B1(
        P3_D_REG_30__SCAN_IN), .B2(keyinput180), .ZN(n13126) );
  OAI221_X1 U15409 ( .B1(P3_REG3_REG_27__SCAN_IN), .B2(keyinput178), .C1(
        P3_D_REG_30__SCAN_IN), .C2(keyinput180), .A(n13126), .ZN(n13129) );
  AOI22_X1 U15410 ( .A1(P3_DATAO_REG_29__SCAN_IN), .A2(keyinput150), .B1(
        P2_IR_REG_28__SCAN_IN), .B2(keyinput252), .ZN(n13127) );
  OAI221_X1 U15411 ( .B1(P3_DATAO_REG_29__SCAN_IN), .B2(keyinput150), .C1(
        P2_IR_REG_28__SCAN_IN), .C2(keyinput252), .A(n13127), .ZN(n13128) );
  NOR4_X1 U15412 ( .A1(n13131), .A2(n13130), .A3(n13129), .A4(n13128), .ZN(
        n13159) );
  AOI22_X1 U15413 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(keyinput212), .B1(
        P2_IR_REG_9__SCAN_IN), .B2(keyinput138), .ZN(n13132) );
  OAI221_X1 U15414 ( .B1(P2_IR_REG_7__SCAN_IN), .B2(keyinput212), .C1(
        P2_IR_REG_9__SCAN_IN), .C2(keyinput138), .A(n13132), .ZN(n13139) );
  AOI22_X1 U15415 ( .A1(P1_REG0_REG_13__SCAN_IN), .A2(keyinput147), .B1(
        P2_REG0_REG_15__SCAN_IN), .B2(keyinput187), .ZN(n13133) );
  OAI221_X1 U15416 ( .B1(P1_REG0_REG_13__SCAN_IN), .B2(keyinput147), .C1(
        P2_REG0_REG_15__SCAN_IN), .C2(keyinput187), .A(n13133), .ZN(n13138) );
  AOI22_X1 U15417 ( .A1(P3_DATAO_REG_30__SCAN_IN), .A2(keyinput142), .B1(
        P3_D_REG_14__SCAN_IN), .B2(keyinput211), .ZN(n13134) );
  OAI221_X1 U15418 ( .B1(P3_DATAO_REG_30__SCAN_IN), .B2(keyinput142), .C1(
        P3_D_REG_14__SCAN_IN), .C2(keyinput211), .A(n13134), .ZN(n13137) );
  AOI22_X1 U15419 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(keyinput249), .B1(
        P3_D_REG_2__SCAN_IN), .B2(keyinput215), .ZN(n13135) );
  OAI221_X1 U15420 ( .B1(P1_DATAO_REG_19__SCAN_IN), .B2(keyinput249), .C1(
        P3_D_REG_2__SCAN_IN), .C2(keyinput215), .A(n13135), .ZN(n13136) );
  NOR4_X1 U15421 ( .A1(n13139), .A2(n13138), .A3(n13137), .A4(n13136), .ZN(
        n13158) );
  AOI22_X1 U15422 ( .A1(P1_D_REG_29__SCAN_IN), .A2(keyinput163), .B1(SI_24_), 
        .B2(keyinput169), .ZN(n13140) );
  OAI221_X1 U15423 ( .B1(P1_D_REG_29__SCAN_IN), .B2(keyinput163), .C1(SI_24_), 
        .C2(keyinput169), .A(n13140), .ZN(n13147) );
  AOI22_X1 U15424 ( .A1(P1_REG1_REG_14__SCAN_IN), .A2(keyinput223), .B1(
        P2_D_REG_7__SCAN_IN), .B2(keyinput132), .ZN(n13141) );
  OAI221_X1 U15425 ( .B1(P1_REG1_REG_14__SCAN_IN), .B2(keyinput223), .C1(
        P2_D_REG_7__SCAN_IN), .C2(keyinput132), .A(n13141), .ZN(n13146) );
  AOI22_X1 U15426 ( .A1(P1_REG0_REG_5__SCAN_IN), .A2(keyinput200), .B1(
        P3_REG3_REG_7__SCAN_IN), .B2(keyinput238), .ZN(n13142) );
  OAI221_X1 U15427 ( .B1(P1_REG0_REG_5__SCAN_IN), .B2(keyinput200), .C1(
        P3_REG3_REG_7__SCAN_IN), .C2(keyinput238), .A(n13142), .ZN(n13145) );
  AOI22_X1 U15428 ( .A1(P3_REG3_REG_0__SCAN_IN), .A2(keyinput198), .B1(
        P3_REG2_REG_10__SCAN_IN), .B2(keyinput131), .ZN(n13143) );
  OAI221_X1 U15429 ( .B1(P3_REG3_REG_0__SCAN_IN), .B2(keyinput198), .C1(
        P3_REG2_REG_10__SCAN_IN), .C2(keyinput131), .A(n13143), .ZN(n13144) );
  NOR4_X1 U15430 ( .A1(n13147), .A2(n13146), .A3(n13145), .A4(n13144), .ZN(
        n13157) );
  AOI22_X1 U15431 ( .A1(P2_REG0_REG_3__SCAN_IN), .A2(keyinput128), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(keyinput177), .ZN(n13148) );
  OAI221_X1 U15432 ( .B1(P2_REG0_REG_3__SCAN_IN), .B2(keyinput128), .C1(
        P2_DATAO_REG_12__SCAN_IN), .C2(keyinput177), .A(n13148), .ZN(n13155)
         );
  AOI22_X1 U15433 ( .A1(P2_REG3_REG_20__SCAN_IN), .A2(keyinput241), .B1(
        P3_REG0_REG_30__SCAN_IN), .B2(keyinput129), .ZN(n13149) );
  OAI221_X1 U15434 ( .B1(P2_REG3_REG_20__SCAN_IN), .B2(keyinput241), .C1(
        P3_REG0_REG_30__SCAN_IN), .C2(keyinput129), .A(n13149), .ZN(n13154) );
  AOI22_X1 U15435 ( .A1(P3_REG2_REG_27__SCAN_IN), .A2(keyinput179), .B1(
        P1_DATAO_REG_5__SCAN_IN), .B2(keyinput151), .ZN(n13150) );
  OAI221_X1 U15436 ( .B1(P3_REG2_REG_27__SCAN_IN), .B2(keyinput179), .C1(
        P1_DATAO_REG_5__SCAN_IN), .C2(keyinput151), .A(n13150), .ZN(n13153) );
  AOI22_X1 U15437 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(keyinput245), .B1(
        P1_D_REG_11__SCAN_IN), .B2(keyinput204), .ZN(n13151) );
  OAI221_X1 U15438 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(keyinput245), .C1(
        P1_D_REG_11__SCAN_IN), .C2(keyinput204), .A(n13151), .ZN(n13152) );
  NOR4_X1 U15439 ( .A1(n13155), .A2(n13154), .A3(n13153), .A4(n13152), .ZN(
        n13156) );
  NAND4_X1 U15440 ( .A1(n13159), .A2(n13158), .A3(n13157), .A4(n13156), .ZN(
        n13289) );
  AOI22_X1 U15441 ( .A1(P3_ADDR_REG_8__SCAN_IN), .A2(keyinput201), .B1(
        P2_REG1_REG_7__SCAN_IN), .B2(keyinput152), .ZN(n13160) );
  OAI221_X1 U15442 ( .B1(P3_ADDR_REG_8__SCAN_IN), .B2(keyinput201), .C1(
        P2_REG1_REG_7__SCAN_IN), .C2(keyinput152), .A(n13160), .ZN(n13167) );
  AOI22_X1 U15443 ( .A1(P3_DATAO_REG_24__SCAN_IN), .A2(keyinput136), .B1(
        P1_REG1_REG_6__SCAN_IN), .B2(keyinput139), .ZN(n13161) );
  OAI221_X1 U15444 ( .B1(P3_DATAO_REG_24__SCAN_IN), .B2(keyinput136), .C1(
        P1_REG1_REG_6__SCAN_IN), .C2(keyinput139), .A(n13161), .ZN(n13166) );
  AOI22_X1 U15445 ( .A1(P1_REG2_REG_27__SCAN_IN), .A2(keyinput190), .B1(
        P2_D_REG_24__SCAN_IN), .B2(keyinput202), .ZN(n13162) );
  OAI221_X1 U15446 ( .B1(P1_REG2_REG_27__SCAN_IN), .B2(keyinput190), .C1(
        P2_D_REG_24__SCAN_IN), .C2(keyinput202), .A(n13162), .ZN(n13165) );
  AOI22_X1 U15447 ( .A1(P2_D_REG_29__SCAN_IN), .A2(keyinput222), .B1(
        P1_DATAO_REG_11__SCAN_IN), .B2(keyinput233), .ZN(n13163) );
  OAI221_X1 U15448 ( .B1(P2_D_REG_29__SCAN_IN), .B2(keyinput222), .C1(
        P1_DATAO_REG_11__SCAN_IN), .C2(keyinput233), .A(n13163), .ZN(n13164)
         );
  NOR4_X1 U15449 ( .A1(n13167), .A2(n13166), .A3(n13165), .A4(n13164), .ZN(
        n13195) );
  AOI22_X1 U15450 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(keyinput194), .B1(
        P2_IR_REG_29__SCAN_IN), .B2(keyinput228), .ZN(n13168) );
  OAI221_X1 U15451 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(keyinput194), .C1(
        P2_IR_REG_29__SCAN_IN), .C2(keyinput228), .A(n13168), .ZN(n13175) );
  AOI22_X1 U15452 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(keyinput251), .B1(
        P1_D_REG_30__SCAN_IN), .B2(keyinput153), .ZN(n13169) );
  OAI221_X1 U15453 ( .B1(P1_ADDR_REG_2__SCAN_IN), .B2(keyinput251), .C1(
        P1_D_REG_30__SCAN_IN), .C2(keyinput153), .A(n13169), .ZN(n13174) );
  AOI22_X1 U15454 ( .A1(P1_REG0_REG_15__SCAN_IN), .A2(keyinput189), .B1(
        P2_REG2_REG_3__SCAN_IN), .B2(keyinput133), .ZN(n13170) );
  OAI221_X1 U15455 ( .B1(P1_REG0_REG_15__SCAN_IN), .B2(keyinput189), .C1(
        P2_REG2_REG_3__SCAN_IN), .C2(keyinput133), .A(n13170), .ZN(n13173) );
  AOI22_X1 U15456 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(keyinput149), .B1(
        P2_REG1_REG_27__SCAN_IN), .B2(keyinput242), .ZN(n13171) );
  OAI221_X1 U15457 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(keyinput149), .C1(
        P2_REG1_REG_27__SCAN_IN), .C2(keyinput242), .A(n13171), .ZN(n13172) );
  NOR4_X1 U15458 ( .A1(n13175), .A2(n13174), .A3(n13173), .A4(n13172), .ZN(
        n13194) );
  AOI22_X1 U15459 ( .A1(P3_REG2_REG_24__SCAN_IN), .A2(keyinput206), .B1(SI_17_), .B2(keyinput248), .ZN(n13176) );
  OAI221_X1 U15460 ( .B1(P3_REG2_REG_24__SCAN_IN), .B2(keyinput206), .C1(
        SI_17_), .C2(keyinput248), .A(n13176), .ZN(n13183) );
  AOI22_X1 U15461 ( .A1(P1_REG2_REG_2__SCAN_IN), .A2(keyinput159), .B1(
        P3_REG2_REG_16__SCAN_IN), .B2(keyinput134), .ZN(n13177) );
  OAI221_X1 U15462 ( .B1(P1_REG2_REG_2__SCAN_IN), .B2(keyinput159), .C1(
        P3_REG2_REG_16__SCAN_IN), .C2(keyinput134), .A(n13177), .ZN(n13182) );
  AOI22_X1 U15463 ( .A1(P1_REG3_REG_25__SCAN_IN), .A2(keyinput217), .B1(
        P1_REG3_REG_28__SCAN_IN), .B2(keyinput154), .ZN(n13178) );
  OAI221_X1 U15464 ( .B1(P1_REG3_REG_25__SCAN_IN), .B2(keyinput217), .C1(
        P1_REG3_REG_28__SCAN_IN), .C2(keyinput154), .A(n13178), .ZN(n13181) );
  AOI22_X1 U15465 ( .A1(P1_DATAO_REG_0__SCAN_IN), .A2(keyinput145), .B1(
        P3_IR_REG_19__SCAN_IN), .B2(keyinput135), .ZN(n13179) );
  OAI221_X1 U15466 ( .B1(P1_DATAO_REG_0__SCAN_IN), .B2(keyinput145), .C1(
        P3_IR_REG_19__SCAN_IN), .C2(keyinput135), .A(n13179), .ZN(n13180) );
  NOR4_X1 U15467 ( .A1(n13183), .A2(n13182), .A3(n13181), .A4(n13180), .ZN(
        n13193) );
  AOI22_X1 U15468 ( .A1(P2_REG3_REG_28__SCAN_IN), .A2(keyinput197), .B1(
        P3_REG2_REG_21__SCAN_IN), .B2(keyinput205), .ZN(n13184) );
  OAI221_X1 U15469 ( .B1(P2_REG3_REG_28__SCAN_IN), .B2(keyinput197), .C1(
        P3_REG2_REG_21__SCAN_IN), .C2(keyinput205), .A(n13184), .ZN(n13191) );
  AOI22_X1 U15470 ( .A1(P2_REG0_REG_25__SCAN_IN), .A2(keyinput158), .B1(
        P3_REG3_REG_8__SCAN_IN), .B2(keyinput157), .ZN(n13185) );
  OAI221_X1 U15471 ( .B1(P2_REG0_REG_25__SCAN_IN), .B2(keyinput158), .C1(
        P3_REG3_REG_8__SCAN_IN), .C2(keyinput157), .A(n13185), .ZN(n13190) );
  AOI22_X1 U15472 ( .A1(P1_REG3_REG_15__SCAN_IN), .A2(keyinput216), .B1(
        P3_REG1_REG_7__SCAN_IN), .B2(keyinput162), .ZN(n13186) );
  OAI221_X1 U15473 ( .B1(P1_REG3_REG_15__SCAN_IN), .B2(keyinput216), .C1(
        P3_REG1_REG_7__SCAN_IN), .C2(keyinput162), .A(n13186), .ZN(n13189) );
  INV_X1 U15474 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n13481) );
  AOI22_X1 U15475 ( .A1(n13426), .A2(keyinput246), .B1(keyinput181), .B2(
        n13481), .ZN(n13187) );
  OAI221_X1 U15476 ( .B1(n13426), .B2(keyinput246), .C1(n13481), .C2(
        keyinput181), .A(n13187), .ZN(n13188) );
  NOR4_X1 U15477 ( .A1(n13191), .A2(n13190), .A3(n13189), .A4(n13188), .ZN(
        n13192) );
  NAND4_X1 U15478 ( .A1(n13195), .A2(n13194), .A3(n13193), .A4(n13192), .ZN(
        n13288) );
  INV_X1 U15479 ( .A(P3_ADDR_REG_18__SCAN_IN), .ZN(n14995) );
  AOI22_X1 U15480 ( .A1(n14995), .A2(keyinput196), .B1(keyinput174), .B2(
        n13405), .ZN(n13196) );
  OAI221_X1 U15481 ( .B1(n14995), .B2(keyinput196), .C1(n13405), .C2(
        keyinput174), .A(n13196), .ZN(n13205) );
  AOI22_X1 U15482 ( .A1(n8707), .A2(keyinput219), .B1(keyinput227), .B2(n13198), .ZN(n13197) );
  OAI221_X1 U15483 ( .B1(n8707), .B2(keyinput219), .C1(n13198), .C2(
        keyinput227), .A(n13197), .ZN(n13204) );
  XOR2_X1 U15484 ( .A(n11941), .B(keyinput240), .Z(n13202) );
  XOR2_X1 U15485 ( .A(n13408), .B(keyinput193), .Z(n13201) );
  XNOR2_X1 U15486 ( .A(P1_IR_REG_1__SCAN_IN), .B(keyinput164), .ZN(n13200) );
  XNOR2_X1 U15487 ( .A(P2_REG3_REG_5__SCAN_IN), .B(keyinput255), .ZN(n13199)
         );
  NAND4_X1 U15488 ( .A1(n13202), .A2(n13201), .A3(n13200), .A4(n13199), .ZN(
        n13203) );
  NOR3_X1 U15489 ( .A1(n13205), .A2(n13204), .A3(n13203), .ZN(n13241) );
  INV_X1 U15490 ( .A(P3_WR_REG_SCAN_IN), .ZN(n13409) );
  AOI22_X1 U15491 ( .A1(n13409), .A2(keyinput230), .B1(n14137), .B2(
        keyinput250), .ZN(n13206) );
  OAI221_X1 U15492 ( .B1(n13409), .B2(keyinput230), .C1(n14137), .C2(
        keyinput250), .A(n13206), .ZN(n13215) );
  INV_X1 U15493 ( .A(P1_D_REG_8__SCAN_IN), .ZN(n15312) );
  AOI22_X1 U15494 ( .A1(n15312), .A2(keyinput140), .B1(n6979), .B2(keyinput207), .ZN(n13207) );
  OAI221_X1 U15495 ( .B1(n15312), .B2(keyinput140), .C1(n6979), .C2(
        keyinput207), .A(n13207), .ZN(n13214) );
  AOI22_X1 U15496 ( .A1(n13209), .A2(keyinput253), .B1(keyinput168), .B2(
        n13421), .ZN(n13208) );
  OAI221_X1 U15497 ( .B1(n13209), .B2(keyinput253), .C1(n13421), .C2(
        keyinput168), .A(n13208), .ZN(n13213) );
  XNOR2_X1 U15498 ( .A(P2_IR_REG_27__SCAN_IN), .B(keyinput243), .ZN(n13211) );
  XNOR2_X1 U15499 ( .A(P2_IR_REG_3__SCAN_IN), .B(keyinput229), .ZN(n13210) );
  NAND2_X1 U15500 ( .A1(n13211), .A2(n13210), .ZN(n13212) );
  NOR4_X1 U15501 ( .A1(n13215), .A2(n13214), .A3(n13213), .A4(n13212), .ZN(
        n13240) );
  INV_X1 U15502 ( .A(P2_D_REG_8__SCAN_IN), .ZN(n15482) );
  INV_X1 U15503 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n13217) );
  AOI22_X1 U15504 ( .A1(n15482), .A2(keyinput176), .B1(keyinput185), .B2(
        n13217), .ZN(n13216) );
  OAI221_X1 U15505 ( .B1(n15482), .B2(keyinput176), .C1(n13217), .C2(
        keyinput185), .A(n13216), .ZN(n13227) );
  AOI22_X1 U15506 ( .A1(n13329), .A2(keyinput191), .B1(keyinput239), .B2(
        n13219), .ZN(n13218) );
  OAI221_X1 U15507 ( .B1(n13329), .B2(keyinput191), .C1(n13219), .C2(
        keyinput239), .A(n13218), .ZN(n13226) );
  INV_X1 U15508 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n13221) );
  INV_X1 U15509 ( .A(P3_REG2_REG_28__SCAN_IN), .ZN(n13376) );
  AOI22_X1 U15510 ( .A1(n13221), .A2(keyinput224), .B1(n13376), .B2(
        keyinput141), .ZN(n13220) );
  OAI221_X1 U15511 ( .B1(n13221), .B2(keyinput224), .C1(n13376), .C2(
        keyinput141), .A(n13220), .ZN(n13225) );
  INV_X1 U15512 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n13223) );
  AOI22_X1 U15513 ( .A1(n13223), .A2(keyinput234), .B1(n13429), .B2(
        keyinput209), .ZN(n13222) );
  OAI221_X1 U15514 ( .B1(n13223), .B2(keyinput234), .C1(n13429), .C2(
        keyinput209), .A(n13222), .ZN(n13224) );
  NOR4_X1 U15515 ( .A1(n13227), .A2(n13226), .A3(n13225), .A4(n13224), .ZN(
        n13239) );
  AOI22_X1 U15516 ( .A1(n8191), .A2(keyinput166), .B1(n13229), .B2(keyinput188), .ZN(n13228) );
  OAI221_X1 U15517 ( .B1(n8191), .B2(keyinput166), .C1(n13229), .C2(
        keyinput188), .A(n13228), .ZN(n13237) );
  INV_X1 U15518 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n13453) );
  XNOR2_X1 U15519 ( .A(keyinput210), .B(n13453), .ZN(n13236) );
  INV_X1 U15520 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n14963) );
  XNOR2_X1 U15521 ( .A(keyinput184), .B(n14963), .ZN(n13235) );
  XNOR2_X1 U15522 ( .A(P3_REG2_REG_19__SCAN_IN), .B(keyinput144), .ZN(n13233)
         );
  XNOR2_X1 U15523 ( .A(P3_IR_REG_26__SCAN_IN), .B(keyinput232), .ZN(n13232) );
  XNOR2_X1 U15524 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(keyinput221), .ZN(n13231)
         );
  XNOR2_X1 U15525 ( .A(P3_IR_REG_25__SCAN_IN), .B(keyinput156), .ZN(n13230) );
  NAND4_X1 U15526 ( .A1(n13233), .A2(n13232), .A3(n13231), .A4(n13230), .ZN(
        n13234) );
  NOR4_X1 U15527 ( .A1(n13237), .A2(n13236), .A3(n13235), .A4(n13234), .ZN(
        n13238) );
  NAND4_X1 U15528 ( .A1(n13241), .A2(n13240), .A3(n13239), .A4(n13238), .ZN(
        n13287) );
  INV_X1 U15529 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n13467) );
  AOI22_X1 U15530 ( .A1(n13467), .A2(keyinput213), .B1(n13243), .B2(
        keyinput171), .ZN(n13242) );
  OAI221_X1 U15531 ( .B1(n13467), .B2(keyinput213), .C1(n13243), .C2(
        keyinput171), .A(n13242), .ZN(n13251) );
  INV_X1 U15532 ( .A(P1_D_REG_20__SCAN_IN), .ZN(n15308) );
  INV_X1 U15533 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n13446) );
  AOI22_X1 U15534 ( .A1(n15308), .A2(keyinput172), .B1(keyinput192), .B2(
        n13446), .ZN(n13244) );
  OAI221_X1 U15535 ( .B1(n15308), .B2(keyinput172), .C1(n13446), .C2(
        keyinput192), .A(n13244), .ZN(n13250) );
  INV_X1 U15536 ( .A(P2_D_REG_17__SCAN_IN), .ZN(n15481) );
  AOI22_X1 U15537 ( .A1(n15481), .A2(keyinput175), .B1(n13246), .B2(
        keyinput254), .ZN(n13245) );
  OAI221_X1 U15538 ( .B1(n15481), .B2(keyinput175), .C1(n13246), .C2(
        keyinput254), .A(n13245), .ZN(n13249) );
  INV_X1 U15539 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n15748) );
  AOI22_X1 U15540 ( .A1(n15748), .A2(keyinput208), .B1(n13428), .B2(
        keyinput195), .ZN(n13247) );
  OAI221_X1 U15541 ( .B1(n15748), .B2(keyinput208), .C1(n13428), .C2(
        keyinput195), .A(n13247), .ZN(n13248) );
  NOR4_X1 U15542 ( .A1(n13251), .A2(n13250), .A3(n13249), .A4(n13248), .ZN(
        n13285) );
  AOI22_X1 U15543 ( .A1(n14803), .A2(keyinput167), .B1(keyinput143), .B2(
        n13310), .ZN(n13252) );
  OAI221_X1 U15544 ( .B1(n14803), .B2(keyinput167), .C1(n13310), .C2(
        keyinput143), .A(n13252), .ZN(n13262) );
  AOI22_X1 U15545 ( .A1(n13254), .A2(keyinput161), .B1(n14809), .B2(
        keyinput237), .ZN(n13253) );
  OAI221_X1 U15546 ( .B1(n13254), .B2(keyinput161), .C1(n14809), .C2(
        keyinput237), .A(n13253), .ZN(n13261) );
  XNOR2_X1 U15547 ( .A(P3_REG1_REG_29__SCAN_IN), .B(keyinput247), .ZN(n13257)
         );
  XNOR2_X1 U15548 ( .A(P2_IR_REG_14__SCAN_IN), .B(keyinput137), .ZN(n13256) );
  XNOR2_X1 U15549 ( .A(P2_IR_REG_25__SCAN_IN), .B(keyinput155), .ZN(n13255) );
  NAND3_X1 U15550 ( .A1(n13257), .A2(n13256), .A3(n13255), .ZN(n13260) );
  XNOR2_X1 U15551 ( .A(n13258), .B(keyinput218), .ZN(n13259) );
  NOR4_X1 U15552 ( .A1(n13262), .A2(n13261), .A3(n13260), .A4(n13259), .ZN(
        n13284) );
  INV_X1 U15553 ( .A(P1_D_REG_17__SCAN_IN), .ZN(n15309) );
  AOI22_X1 U15554 ( .A1(n13317), .A2(keyinput182), .B1(keyinput199), .B2(
        n15309), .ZN(n13263) );
  OAI221_X1 U15555 ( .B1(n13317), .B2(keyinput182), .C1(n15309), .C2(
        keyinput199), .A(n13263), .ZN(n13271) );
  AOI22_X1 U15556 ( .A1(n8046), .A2(keyinput244), .B1(n13311), .B2(keyinput231), .ZN(n13264) );
  OAI221_X1 U15557 ( .B1(n8046), .B2(keyinput244), .C1(n13311), .C2(
        keyinput231), .A(n13264), .ZN(n13270) );
  AOI22_X1 U15558 ( .A1(n13454), .A2(keyinput225), .B1(keyinput183), .B2(
        n13266), .ZN(n13265) );
  OAI221_X1 U15559 ( .B1(n13454), .B2(keyinput225), .C1(n13266), .C2(
        keyinput183), .A(n13265), .ZN(n13269) );
  INV_X1 U15560 ( .A(P1_D_REG_10__SCAN_IN), .ZN(n15311) );
  AOI22_X1 U15561 ( .A1(n13425), .A2(keyinput146), .B1(keyinput214), .B2(
        n15311), .ZN(n13267) );
  OAI221_X1 U15562 ( .B1(n13425), .B2(keyinput146), .C1(n15311), .C2(
        keyinput214), .A(n13267), .ZN(n13268) );
  NOR4_X1 U15563 ( .A1(n13271), .A2(n13270), .A3(n13269), .A4(n13268), .ZN(
        n13283) );
  INV_X1 U15564 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n15355) );
  AOI22_X1 U15565 ( .A1(n12670), .A2(keyinput165), .B1(keyinput226), .B2(
        n15355), .ZN(n13272) );
  OAI221_X1 U15566 ( .B1(n12670), .B2(keyinput165), .C1(n15355), .C2(
        keyinput226), .A(n13272), .ZN(n13281) );
  AOI22_X1 U15567 ( .A1(n13274), .A2(keyinput148), .B1(keyinput203), .B2(
        n15396), .ZN(n13273) );
  OAI221_X1 U15568 ( .B1(n13274), .B2(keyinput148), .C1(n15396), .C2(
        keyinput203), .A(n13273), .ZN(n13280) );
  AOI22_X1 U15569 ( .A1(n15027), .A2(keyinput220), .B1(n13466), .B2(
        keyinput186), .ZN(n13275) );
  OAI221_X1 U15570 ( .B1(n15027), .B2(keyinput220), .C1(n13466), .C2(
        keyinput186), .A(n13275), .ZN(n13279) );
  AOI22_X1 U15571 ( .A1(n13277), .A2(keyinput170), .B1(keyinput236), .B2(n9708), .ZN(n13276) );
  OAI221_X1 U15572 ( .B1(n13277), .B2(keyinput170), .C1(n9708), .C2(
        keyinput236), .A(n13276), .ZN(n13278) );
  NOR4_X1 U15573 ( .A1(n13281), .A2(n13280), .A3(n13279), .A4(n13278), .ZN(
        n13282) );
  NAND4_X1 U15574 ( .A1(n13285), .A2(n13284), .A3(n13283), .A4(n13282), .ZN(
        n13286) );
  OR4_X1 U15575 ( .A1(n13289), .A2(n13288), .A3(n13287), .A4(n13286), .ZN(
        n13491) );
  OAI22_X1 U15576 ( .A1(P2_DATAO_REG_30__SCAN_IN), .A2(keyinput39), .B1(
        keyinput95), .B2(P1_REG1_REG_14__SCAN_IN), .ZN(n13290) );
  AOI221_X1 U15577 ( .B1(P2_DATAO_REG_30__SCAN_IN), .B2(keyinput39), .C1(
        P1_REG1_REG_14__SCAN_IN), .C2(keyinput95), .A(n13290), .ZN(n13297) );
  OAI22_X1 U15578 ( .A1(P2_DATAO_REG_12__SCAN_IN), .A2(keyinput49), .B1(
        P1_D_REG_10__SCAN_IN), .B2(keyinput86), .ZN(n13291) );
  AOI221_X1 U15579 ( .B1(P2_DATAO_REG_12__SCAN_IN), .B2(keyinput49), .C1(
        keyinput86), .C2(P1_D_REG_10__SCAN_IN), .A(n13291), .ZN(n13296) );
  OAI22_X1 U15580 ( .A1(P3_D_REG_6__SCAN_IN), .A2(keyinput42), .B1(
        P3_REG1_REG_25__SCAN_IN), .B2(keyinput60), .ZN(n13292) );
  AOI221_X1 U15581 ( .B1(P3_D_REG_6__SCAN_IN), .B2(keyinput42), .C1(keyinput60), .C2(P3_REG1_REG_25__SCAN_IN), .A(n13292), .ZN(n13295) );
  OAI22_X1 U15582 ( .A1(P1_REG1_REG_27__SCAN_IN), .A2(keyinput106), .B1(
        P1_ADDR_REG_11__SCAN_IN), .B2(keyinput66), .ZN(n13293) );
  AOI221_X1 U15583 ( .B1(P1_REG1_REG_27__SCAN_IN), .B2(keyinput106), .C1(
        keyinput66), .C2(P1_ADDR_REG_11__SCAN_IN), .A(n13293), .ZN(n13294) );
  NAND4_X1 U15584 ( .A1(n13297), .A2(n13296), .A3(n13295), .A4(n13294), .ZN(
        n13307) );
  OAI22_X1 U15585 ( .A1(P1_DATAO_REG_5__SCAN_IN), .A2(keyinput23), .B1(
        P3_REG2_REG_0__SCAN_IN), .B2(keyinput33), .ZN(n13298) );
  AOI221_X1 U15586 ( .B1(P1_DATAO_REG_5__SCAN_IN), .B2(keyinput23), .C1(
        keyinput33), .C2(P3_REG2_REG_0__SCAN_IN), .A(n13298), .ZN(n13305) );
  OAI22_X1 U15587 ( .A1(P2_REG1_REG_27__SCAN_IN), .A2(keyinput114), .B1(
        keyinput36), .B2(P1_IR_REG_1__SCAN_IN), .ZN(n13299) );
  AOI221_X1 U15588 ( .B1(P2_REG1_REG_27__SCAN_IN), .B2(keyinput114), .C1(
        P1_IR_REG_1__SCAN_IN), .C2(keyinput36), .A(n13299), .ZN(n13304) );
  OAI22_X1 U15589 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(keyinput126), .B1(
        P1_REG1_REG_28__SCAN_IN), .B2(keyinput57), .ZN(n13300) );
  AOI221_X1 U15590 ( .B1(P1_DATAO_REG_28__SCAN_IN), .B2(keyinput126), .C1(
        keyinput57), .C2(P1_REG1_REG_28__SCAN_IN), .A(n13300), .ZN(n13303) );
  OAI22_X1 U15591 ( .A1(P3_REG2_REG_29__SCAN_IN), .A2(keyinput112), .B1(
        P3_REG2_REG_24__SCAN_IN), .B2(keyinput78), .ZN(n13301) );
  AOI221_X1 U15592 ( .B1(P3_REG2_REG_29__SCAN_IN), .B2(keyinput112), .C1(
        keyinput78), .C2(P3_REG2_REG_24__SCAN_IN), .A(n13301), .ZN(n13302) );
  NAND4_X1 U15593 ( .A1(n13305), .A2(n13304), .A3(n13303), .A4(n13302), .ZN(
        n13306) );
  NOR2_X1 U15594 ( .A1(n13307), .A2(n13306), .ZN(n13325) );
  INV_X1 U15595 ( .A(P1_D_REG_29__SCAN_IN), .ZN(n15307) );
  AOI22_X1 U15596 ( .A1(n15307), .A2(keyinput35), .B1(keyinput44), .B2(n15308), 
        .ZN(n13308) );
  OAI221_X1 U15597 ( .B1(n15307), .B2(keyinput35), .C1(n15308), .C2(keyinput44), .A(n13308), .ZN(n13313) );
  AOI22_X1 U15598 ( .A1(n13311), .A2(keyinput103), .B1(keyinput15), .B2(n13310), .ZN(n13309) );
  OAI221_X1 U15599 ( .B1(n13311), .B2(keyinput103), .C1(n13310), .C2(
        keyinput15), .A(n13309), .ZN(n13312) );
  NOR2_X1 U15600 ( .A1(n13313), .A2(n13312), .ZN(n13324) );
  INV_X1 U15601 ( .A(P2_D_REG_7__SCAN_IN), .ZN(n15483) );
  AOI22_X1 U15602 ( .A1(n15483), .A2(keyinput4), .B1(keyinput30), .B2(n13315), 
        .ZN(n13314) );
  OAI221_X1 U15603 ( .B1(n15483), .B2(keyinput4), .C1(n13315), .C2(keyinput30), 
        .A(n13314), .ZN(n13322) );
  AOI22_X1 U15604 ( .A1(n13318), .A2(keyinput52), .B1(keyinput54), .B2(n13317), 
        .ZN(n13316) );
  OAI221_X1 U15605 ( .B1(n13318), .B2(keyinput52), .C1(n13317), .C2(keyinput54), .A(n13316), .ZN(n13321) );
  XNOR2_X1 U15606 ( .A(n13319), .B(keyinput22), .ZN(n13320) );
  NOR3_X1 U15607 ( .A1(n13322), .A2(n13321), .A3(n13320), .ZN(n13323) );
  NAND3_X1 U15608 ( .A1(n13325), .A2(n13324), .A3(n13323), .ZN(n13354) );
  OAI22_X1 U15609 ( .A1(P1_D_REG_17__SCAN_IN), .A2(keyinput71), .B1(
        P1_REG2_REG_20__SCAN_IN), .B2(keyinput99), .ZN(n13326) );
  AOI221_X1 U15610 ( .B1(P1_D_REG_17__SCAN_IN), .B2(keyinput71), .C1(
        keyinput99), .C2(P1_REG2_REG_20__SCAN_IN), .A(n13326), .ZN(n13334) );
  OAI22_X1 U15611 ( .A1(P3_REG2_REG_19__SCAN_IN), .A2(keyinput16), .B1(
        P1_REG0_REG_7__SCAN_IN), .B2(keyinput98), .ZN(n13327) );
  AOI221_X1 U15612 ( .B1(P3_REG2_REG_19__SCAN_IN), .B2(keyinput16), .C1(
        keyinput98), .C2(P1_REG0_REG_7__SCAN_IN), .A(n13327), .ZN(n13333) );
  OAI22_X1 U15613 ( .A1(n13329), .A2(keyinput63), .B1(n15312), .B2(keyinput12), 
        .ZN(n13328) );
  AOI221_X1 U15614 ( .B1(n13329), .B2(keyinput63), .C1(keyinput12), .C2(n15312), .A(n13328), .ZN(n13332) );
  OAI22_X1 U15615 ( .A1(P1_DATAO_REG_2__SCAN_IN), .A2(keyinput93), .B1(
        P2_REG0_REG_3__SCAN_IN), .B2(keyinput0), .ZN(n13330) );
  AOI221_X1 U15616 ( .B1(P1_DATAO_REG_2__SCAN_IN), .B2(keyinput93), .C1(
        keyinput0), .C2(P2_REG0_REG_3__SCAN_IN), .A(n13330), .ZN(n13331) );
  NAND4_X1 U15617 ( .A1(n13334), .A2(n13333), .A3(n13332), .A4(n13331), .ZN(
        n13353) );
  OAI22_X1 U15618 ( .A1(P1_DATAO_REG_11__SCAN_IN), .A2(keyinput105), .B1(
        keyinput5), .B2(P2_REG2_REG_3__SCAN_IN), .ZN(n13335) );
  AOI221_X1 U15619 ( .B1(P1_DATAO_REG_11__SCAN_IN), .B2(keyinput105), .C1(
        P2_REG2_REG_3__SCAN_IN), .C2(keyinput5), .A(n13335), .ZN(n13342) );
  OAI22_X1 U15620 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(keyinput91), .B1(
        P3_ADDR_REG_18__SCAN_IN), .B2(keyinput68), .ZN(n13336) );
  AOI221_X1 U15621 ( .B1(P2_REG3_REG_9__SCAN_IN), .B2(keyinput91), .C1(
        keyinput68), .C2(P3_ADDR_REG_18__SCAN_IN), .A(n13336), .ZN(n13341) );
  OAI22_X1 U15622 ( .A1(P2_D_REG_25__SCAN_IN), .A2(keyinput45), .B1(
        P1_REG0_REG_15__SCAN_IN), .B2(keyinput61), .ZN(n13337) );
  AOI221_X1 U15623 ( .B1(P2_D_REG_25__SCAN_IN), .B2(keyinput45), .C1(
        keyinput61), .C2(P1_REG0_REG_15__SCAN_IN), .A(n13337), .ZN(n13340) );
  OAI22_X1 U15624 ( .A1(P3_REG1_REG_20__SCAN_IN), .A2(keyinput111), .B1(
        P2_IR_REG_29__SCAN_IN), .B2(keyinput100), .ZN(n13338) );
  AOI221_X1 U15625 ( .B1(P3_REG1_REG_20__SCAN_IN), .B2(keyinput111), .C1(
        keyinput100), .C2(P2_IR_REG_29__SCAN_IN), .A(n13338), .ZN(n13339) );
  NAND4_X1 U15626 ( .A1(n13342), .A2(n13341), .A3(n13340), .A4(n13339), .ZN(
        n13352) );
  OAI22_X1 U15627 ( .A1(P2_D_REG_17__SCAN_IN), .A2(keyinput47), .B1(keyinput94), .B2(P2_D_REG_29__SCAN_IN), .ZN(n13343) );
  AOI221_X1 U15628 ( .B1(P2_D_REG_17__SCAN_IN), .B2(keyinput47), .C1(
        P2_D_REG_29__SCAN_IN), .C2(keyinput94), .A(n13343), .ZN(n13350) );
  OAI22_X1 U15629 ( .A1(P3_D_REG_14__SCAN_IN), .A2(keyinput83), .B1(
        P1_REG2_REG_27__SCAN_IN), .B2(keyinput62), .ZN(n13344) );
  AOI221_X1 U15630 ( .B1(P3_D_REG_14__SCAN_IN), .B2(keyinput83), .C1(
        keyinput62), .C2(P1_REG2_REG_27__SCAN_IN), .A(n13344), .ZN(n13349) );
  OAI22_X1 U15631 ( .A1(P1_REG0_REG_18__SCAN_IN), .A2(keyinput96), .B1(
        keyinput56), .B2(P1_REG0_REG_12__SCAN_IN), .ZN(n13345) );
  AOI221_X1 U15632 ( .B1(P1_REG0_REG_18__SCAN_IN), .B2(keyinput96), .C1(
        P1_REG0_REG_12__SCAN_IN), .C2(keyinput56), .A(n13345), .ZN(n13348) );
  OAI22_X1 U15633 ( .A1(P1_DATAO_REG_4__SCAN_IN), .A2(keyinput20), .B1(
        P2_IR_REG_14__SCAN_IN), .B2(keyinput9), .ZN(n13346) );
  AOI221_X1 U15634 ( .B1(P1_DATAO_REG_4__SCAN_IN), .B2(keyinput20), .C1(
        keyinput9), .C2(P2_IR_REG_14__SCAN_IN), .A(n13346), .ZN(n13347) );
  NAND4_X1 U15635 ( .A1(n13350), .A2(n13349), .A3(n13348), .A4(n13347), .ZN(
        n13351) );
  NOR4_X1 U15636 ( .A1(n13354), .A2(n13353), .A3(n13352), .A4(n13351), .ZN(
        n13417) );
  INV_X1 U15637 ( .A(P1_D_REG_11__SCAN_IN), .ZN(n15310) );
  OAI22_X1 U15638 ( .A1(n9211), .A2(keyinput69), .B1(n15310), .B2(keyinput76), 
        .ZN(n13355) );
  AOI221_X1 U15639 ( .B1(n9211), .B2(keyinput69), .C1(keyinput76), .C2(n15310), 
        .A(n13355), .ZN(n13416) );
  XOR2_X1 U15640 ( .A(P3_REG3_REG_27__SCAN_IN), .B(keyinput50), .Z(n13359) );
  XOR2_X1 U15641 ( .A(P1_IR_REG_31__SCAN_IN), .B(keyinput32), .Z(n13358) );
  XOR2_X1 U15642 ( .A(P1_REG2_REG_2__SCAN_IN), .B(keyinput31), .Z(n13357) );
  XNOR2_X1 U15643 ( .A(n6979), .B(keyinput79), .ZN(n13356) );
  NOR4_X1 U15644 ( .A1(n13359), .A2(n13358), .A3(n13357), .A4(n13356), .ZN(
        n13384) );
  XOR2_X1 U15645 ( .A(P2_IR_REG_7__SCAN_IN), .B(keyinput84), .Z(n13364) );
  XOR2_X1 U15646 ( .A(P2_IR_REG_25__SCAN_IN), .B(keyinput27), .Z(n13363) );
  XNOR2_X1 U15647 ( .A(n8699), .B(keyinput10), .ZN(n13362) );
  XNOR2_X1 U15648 ( .A(n13360), .B(keyinput101), .ZN(n13361) );
  NOR4_X1 U15649 ( .A1(n13364), .A2(n13363), .A3(n13362), .A4(n13361), .ZN(
        n13383) );
  XNOR2_X1 U15650 ( .A(n13365), .B(keyinput124), .ZN(n13372) );
  XNOR2_X1 U15651 ( .A(n13366), .B(keyinput115), .ZN(n13371) );
  XNOR2_X1 U15652 ( .A(n13367), .B(keyinput7), .ZN(n13370) );
  XNOR2_X1 U15653 ( .A(n13368), .B(keyinput104), .ZN(n13369) );
  NOR4_X1 U15654 ( .A1(n13372), .A2(n13371), .A3(n13370), .A4(n13369), .ZN(
        n13382) );
  XNOR2_X1 U15655 ( .A(n13373), .B(keyinput51), .ZN(n13380) );
  XNOR2_X1 U15656 ( .A(n13374), .B(keyinput28), .ZN(n13379) );
  INV_X1 U15657 ( .A(P3_REG3_REG_7__SCAN_IN), .ZN(n13375) );
  XNOR2_X1 U15658 ( .A(keyinput110), .B(n13375), .ZN(n13378) );
  XNOR2_X1 U15659 ( .A(keyinput13), .B(n13376), .ZN(n13377) );
  NOR4_X1 U15660 ( .A1(n13380), .A2(n13379), .A3(n13378), .A4(n13377), .ZN(
        n13381) );
  NAND4_X1 U15661 ( .A1(n13384), .A2(n13383), .A3(n13382), .A4(n13381), .ZN(
        n13394) );
  OAI22_X1 U15662 ( .A1(P1_DATAO_REG_8__SCAN_IN), .A2(keyinput125), .B1(
        P2_REG3_REG_5__SCAN_IN), .B2(keyinput127), .ZN(n13385) );
  AOI221_X1 U15663 ( .B1(P1_DATAO_REG_8__SCAN_IN), .B2(keyinput125), .C1(
        keyinput127), .C2(P2_REG3_REG_5__SCAN_IN), .A(n13385), .ZN(n13392) );
  OAI22_X1 U15664 ( .A1(P3_ADDR_REG_19__SCAN_IN), .A2(keyinput37), .B1(
        P3_DATAO_REG_28__SCAN_IN), .B2(keyinput90), .ZN(n13386) );
  AOI221_X1 U15665 ( .B1(P3_ADDR_REG_19__SCAN_IN), .B2(keyinput37), .C1(
        keyinput90), .C2(P3_DATAO_REG_28__SCAN_IN), .A(n13386), .ZN(n13391) );
  OAI22_X1 U15666 ( .A1(P3_REG0_REG_19__SCAN_IN), .A2(keyinput43), .B1(
        keyinput117), .B2(P2_ADDR_REG_11__SCAN_IN), .ZN(n13387) );
  AOI221_X1 U15667 ( .B1(P3_REG0_REG_19__SCAN_IN), .B2(keyinput43), .C1(
        P2_ADDR_REG_11__SCAN_IN), .C2(keyinput117), .A(n13387), .ZN(n13390) );
  OAI22_X1 U15668 ( .A1(P3_REG0_REG_5__SCAN_IN), .A2(keyinput80), .B1(
        keyinput14), .B2(P3_DATAO_REG_30__SCAN_IN), .ZN(n13388) );
  AOI221_X1 U15669 ( .B1(P3_REG0_REG_5__SCAN_IN), .B2(keyinput80), .C1(
        P3_DATAO_REG_30__SCAN_IN), .C2(keyinput14), .A(n13388), .ZN(n13389) );
  NAND4_X1 U15670 ( .A1(n13392), .A2(n13391), .A3(n13390), .A4(n13389), .ZN(
        n13393) );
  NOR2_X1 U15671 ( .A1(n13394), .A2(n13393), .ZN(n13415) );
  OAI22_X1 U15672 ( .A1(SI_24_), .A2(keyinput41), .B1(keyinput74), .B2(
        P2_D_REG_24__SCAN_IN), .ZN(n13395) );
  AOI221_X1 U15673 ( .B1(SI_24_), .B2(keyinput41), .C1(P2_D_REG_24__SCAN_IN), 
        .C2(keyinput74), .A(n13395), .ZN(n13402) );
  OAI22_X1 U15674 ( .A1(P3_D_REG_2__SCAN_IN), .A2(keyinput87), .B1(
        P2_REG3_REG_10__SCAN_IN), .B2(keyinput55), .ZN(n13396) );
  AOI221_X1 U15675 ( .B1(P3_D_REG_2__SCAN_IN), .B2(keyinput87), .C1(keyinput55), .C2(P2_REG3_REG_10__SCAN_IN), .A(n13396), .ZN(n13401) );
  OAI22_X1 U15676 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(keyinput109), .B1(
        keyinput123), .B2(P1_ADDR_REG_2__SCAN_IN), .ZN(n13397) );
  AOI221_X1 U15677 ( .B1(P2_DATAO_REG_28__SCAN_IN), .B2(keyinput109), .C1(
        P1_ADDR_REG_2__SCAN_IN), .C2(keyinput123), .A(n13397), .ZN(n13400) );
  OAI22_X1 U15678 ( .A1(P2_D_REG_8__SCAN_IN), .A2(keyinput48), .B1(keyinput113), .B2(P2_REG3_REG_20__SCAN_IN), .ZN(n13398) );
  AOI221_X1 U15679 ( .B1(P2_D_REG_8__SCAN_IN), .B2(keyinput48), .C1(
        P2_REG3_REG_20__SCAN_IN), .C2(keyinput113), .A(n13398), .ZN(n13399) );
  NAND4_X1 U15680 ( .A1(n13402), .A2(n13401), .A3(n13400), .A4(n13399), .ZN(
        n13413) );
  AOI22_X1 U15681 ( .A1(n13405), .A2(keyinput46), .B1(n13404), .B2(keyinput88), 
        .ZN(n13403) );
  OAI221_X1 U15682 ( .B1(n13405), .B2(keyinput46), .C1(n13404), .C2(keyinput88), .A(n13403), .ZN(n13412) );
  AOI22_X1 U15683 ( .A1(n13408), .A2(keyinput65), .B1(n13407), .B2(keyinput6), 
        .ZN(n13406) );
  OAI221_X1 U15684 ( .B1(n13408), .B2(keyinput65), .C1(n13407), .C2(keyinput6), 
        .A(n13406), .ZN(n13411) );
  XNOR2_X1 U15685 ( .A(n13409), .B(keyinput102), .ZN(n13410) );
  NOR4_X1 U15686 ( .A1(n13413), .A2(n13412), .A3(n13411), .A4(n13410), .ZN(
        n13414) );
  AND4_X1 U15687 ( .A1(n13417), .A2(n13416), .A3(n13415), .A4(n13414), .ZN(
        n13464) );
  INV_X1 U15688 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n15784) );
  INV_X1 U15689 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n14846) );
  OAI22_X1 U15690 ( .A1(n15784), .A2(keyinput34), .B1(n14846), .B2(keyinput107), .ZN(n13418) );
  AOI221_X1 U15691 ( .B1(n15784), .B2(keyinput34), .C1(keyinput107), .C2(
        n14846), .A(n13418), .ZN(n13463) );
  INV_X1 U15692 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n13420) );
  OAI22_X1 U15693 ( .A1(n13421), .A2(keyinput40), .B1(n13420), .B2(keyinput59), 
        .ZN(n13419) );
  AOI221_X1 U15694 ( .B1(n13421), .B2(keyinput40), .C1(keyinput59), .C2(n13420), .A(n13419), .ZN(n13462) );
  AOI22_X1 U15695 ( .A1(n13423), .A2(keyinput121), .B1(keyinput70), .B2(n9887), 
        .ZN(n13422) );
  OAI221_X1 U15696 ( .B1(n13423), .B2(keyinput121), .C1(n9887), .C2(keyinput70), .A(n13422), .ZN(n13432) );
  AOI22_X1 U15697 ( .A1(n13426), .A2(keyinput118), .B1(keyinput18), .B2(n13425), .ZN(n13424) );
  OAI221_X1 U15698 ( .B1(n13426), .B2(keyinput118), .C1(n13425), .C2(
        keyinput18), .A(n13424), .ZN(n13431) );
  AOI22_X1 U15699 ( .A1(n13429), .A2(keyinput81), .B1(keyinput67), .B2(n13428), 
        .ZN(n13427) );
  OAI221_X1 U15700 ( .B1(n13429), .B2(keyinput81), .C1(n13428), .C2(keyinput67), .A(n13427), .ZN(n13430) );
  NOR3_X1 U15701 ( .A1(n13432), .A2(n13431), .A3(n13430), .ZN(n13460) );
  AOI22_X1 U15702 ( .A1(n14836), .A2(keyinput73), .B1(n13434), .B2(keyinput17), 
        .ZN(n13433) );
  OAI221_X1 U15703 ( .B1(n14836), .B2(keyinput73), .C1(n13434), .C2(keyinput17), .A(n13433), .ZN(n13437) );
  AOI22_X1 U15704 ( .A1(n8046), .A2(keyinput116), .B1(n15027), .B2(keyinput92), 
        .ZN(n13435) );
  OAI221_X1 U15705 ( .B1(n8046), .B2(keyinput116), .C1(n15027), .C2(keyinput92), .A(n13435), .ZN(n13436) );
  NOR2_X1 U15706 ( .A1(n13437), .A2(n13436), .ZN(n13459) );
  AOI22_X1 U15707 ( .A1(n15394), .A2(keyinput11), .B1(n13439), .B2(keyinput120), .ZN(n13438) );
  OAI221_X1 U15708 ( .B1(n15394), .B2(keyinput11), .C1(n13439), .C2(
        keyinput120), .A(n13438), .ZN(n13443) );
  AOI22_X1 U15709 ( .A1(n8191), .A2(keyinput38), .B1(keyinput26), .B2(n13441), 
        .ZN(n13440) );
  OAI221_X1 U15710 ( .B1(n8191), .B2(keyinput38), .C1(n13441), .C2(keyinput26), 
        .A(n13440), .ZN(n13442) );
  NOR2_X1 U15711 ( .A1(n13443), .A2(n13442), .ZN(n13458) );
  AOI22_X1 U15712 ( .A1(n13446), .A2(keyinput64), .B1(n13445), .B2(keyinput29), 
        .ZN(n13444) );
  OAI221_X1 U15713 ( .B1(n13446), .B2(keyinput64), .C1(n13445), .C2(keyinput29), .A(n13444), .ZN(n13447) );
  INV_X1 U15714 ( .A(n13447), .ZN(n13451) );
  INV_X1 U15715 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n15244) );
  XNOR2_X1 U15716 ( .A(keyinput21), .B(n15244), .ZN(n13449) );
  XNOR2_X1 U15717 ( .A(keyinput3), .B(n11343), .ZN(n13448) );
  NOR2_X1 U15718 ( .A1(n13449), .A2(n13448), .ZN(n13450) );
  NAND2_X1 U15719 ( .A1(n13451), .A2(n13450), .ZN(n13456) );
  AOI22_X1 U15720 ( .A1(n13454), .A2(keyinput97), .B1(keyinput82), .B2(n13453), 
        .ZN(n13452) );
  OAI221_X1 U15721 ( .B1(n13454), .B2(keyinput97), .C1(n13453), .C2(keyinput82), .A(n13452), .ZN(n13455) );
  NOR2_X1 U15722 ( .A1(n13456), .A2(n13455), .ZN(n13457) );
  AND4_X1 U15723 ( .A1(n13460), .A2(n13459), .A3(n13458), .A4(n13457), .ZN(
        n13461) );
  AND4_X1 U15724 ( .A1(n13464), .A2(n13463), .A3(n13462), .A4(n13461), .ZN(
        n13490) );
  AOI22_X1 U15725 ( .A1(n13467), .A2(keyinput85), .B1(n13466), .B2(keyinput58), 
        .ZN(n13465) );
  OAI221_X1 U15726 ( .B1(n13467), .B2(keyinput85), .C1(n13466), .C2(keyinput58), .A(n13465), .ZN(n13476) );
  INV_X1 U15727 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n15232) );
  AOI22_X1 U15728 ( .A1(n15232), .A2(keyinput19), .B1(n15114), .B2(keyinput1), 
        .ZN(n13468) );
  OAI221_X1 U15729 ( .B1(n15232), .B2(keyinput19), .C1(n15114), .C2(keyinput1), 
        .A(n13468), .ZN(n13475) );
  AOI22_X1 U15730 ( .A1(n13471), .A2(keyinput2), .B1(keyinput8), .B2(n13470), 
        .ZN(n13469) );
  OAI221_X1 U15731 ( .B1(n13471), .B2(keyinput2), .C1(n13470), .C2(keyinput8), 
        .A(n13469), .ZN(n13474) );
  AOI22_X1 U15732 ( .A1(n15396), .A2(keyinput75), .B1(n9708), .B2(keyinput108), 
        .ZN(n13472) );
  OAI221_X1 U15733 ( .B1(n15396), .B2(keyinput75), .C1(n9708), .C2(keyinput108), .A(n13472), .ZN(n13473) );
  NOR4_X1 U15734 ( .A1(n13476), .A2(n13475), .A3(n13474), .A4(n13473), .ZN(
        n13489) );
  INV_X1 U15735 ( .A(P1_D_REG_30__SCAN_IN), .ZN(n15306) );
  AOI22_X1 U15736 ( .A1(n15306), .A2(keyinput25), .B1(n9487), .B2(keyinput24), 
        .ZN(n13477) );
  OAI221_X1 U15737 ( .B1(n15306), .B2(keyinput25), .C1(n9487), .C2(keyinput24), 
        .A(n13477), .ZN(n13487) );
  AOI22_X1 U15738 ( .A1(n12811), .A2(keyinput77), .B1(n13479), .B2(keyinput119), .ZN(n13478) );
  OAI221_X1 U15739 ( .B1(n12811), .B2(keyinput77), .C1(n13479), .C2(
        keyinput119), .A(n13478), .ZN(n13486) );
  AOI22_X1 U15740 ( .A1(n14137), .A2(keyinput122), .B1(keyinput53), .B2(n13481), .ZN(n13480) );
  OAI221_X1 U15741 ( .B1(n14137), .B2(keyinput122), .C1(n13481), .C2(
        keyinput53), .A(n13480), .ZN(n13485) );
  AOI22_X1 U15742 ( .A1(n13483), .A2(keyinput72), .B1(n14106), .B2(keyinput89), 
        .ZN(n13482) );
  OAI221_X1 U15743 ( .B1(n13483), .B2(keyinput72), .C1(n14106), .C2(keyinput89), .A(n13482), .ZN(n13484) );
  NOR4_X1 U15744 ( .A1(n13487), .A2(n13486), .A3(n13485), .A4(n13484), .ZN(
        n13488) );
  NAND4_X1 U15745 ( .A1(n13491), .A2(n13490), .A3(n13489), .A4(n13488), .ZN(
        n13492) );
  XNOR2_X1 U15746 ( .A(n13493), .B(n13492), .ZN(P2_U3195) );
  XNOR2_X1 U15747 ( .A(n13495), .B(n13494), .ZN(n13502) );
  OAI22_X1 U15748 ( .A1(n13498), .A2(n13630), .B1(n13497), .B2(n13496), .ZN(
        n13758) );
  AOI22_X1 U15749 ( .A1(n13758), .A2(n15125), .B1(P2_REG3_REG_25__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13499) );
  OAI21_X1 U15750 ( .B1(n13762), .B2(n15131), .A(n13499), .ZN(n13500) );
  AOI21_X1 U15751 ( .B1(n13927), .B2(n15128), .A(n13500), .ZN(n13501) );
  OAI21_X1 U15752 ( .B1(n13502), .B2(n13561), .A(n13501), .ZN(P2_U3197) );
  INV_X1 U15753 ( .A(n13985), .ZN(n13891) );
  INV_X1 U15754 ( .A(n11924), .ZN(n13506) );
  INV_X1 U15755 ( .A(n13503), .ZN(n13505) );
  NOR3_X1 U15756 ( .A1(n13506), .A2(n13505), .A3(n13504), .ZN(n13509) );
  INV_X1 U15757 ( .A(n13507), .ZN(n13508) );
  OAI21_X1 U15758 ( .B1(n13509), .B2(n13508), .A(n15123), .ZN(n13515) );
  NAND2_X1 U15759 ( .A1(n13672), .A2(n13555), .ZN(n13511) );
  NAND2_X1 U15760 ( .A1(n13643), .A2(n13701), .ZN(n13510) );
  AND2_X1 U15761 ( .A1(n13511), .A2(n13510), .ZN(n13876) );
  OAI21_X1 U15762 ( .B1(n13558), .B2(n13876), .A(n13512), .ZN(n13513) );
  AOI21_X1 U15763 ( .B1(n13887), .B2(n13556), .A(n13513), .ZN(n13514) );
  OAI211_X1 U15764 ( .C1(n13891), .C2(n13542), .A(n13515), .B(n13514), .ZN(
        P2_U3198) );
  OAI21_X1 U15765 ( .B1(n13518), .B2(n13517), .A(n13516), .ZN(n13519) );
  NAND2_X1 U15766 ( .A1(n13519), .A2(n15123), .ZN(n13523) );
  AOI22_X1 U15767 ( .A1(n13555), .A2(n13675), .B1(n13670), .B2(n13701), .ZN(
        n13977) );
  OAI21_X1 U15768 ( .B1(n13558), .B2(n13977), .A(n13520), .ZN(n13521) );
  AOI21_X1 U15769 ( .B1(n13864), .B2(n13556), .A(n13521), .ZN(n13522) );
  OAI211_X1 U15770 ( .C1(n13979), .C2(n13542), .A(n13523), .B(n13522), .ZN(
        P2_U3200) );
  XNOR2_X1 U15771 ( .A(n13524), .B(n13525), .ZN(n13531) );
  AND2_X1 U15772 ( .A1(n13686), .A2(n13701), .ZN(n13526) );
  AOI21_X1 U15773 ( .B1(n13688), .B2(n13555), .A(n13526), .ZN(n13932) );
  OAI22_X1 U15774 ( .A1(n13932), .A2(n13558), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13527), .ZN(n13528) );
  AOI21_X1 U15775 ( .B1(n13776), .B2(n13556), .A(n13528), .ZN(n13530) );
  NAND2_X1 U15776 ( .A1(n13935), .A2(n15128), .ZN(n13529) );
  OAI211_X1 U15777 ( .C1(n13531), .C2(n13561), .A(n13530), .B(n13529), .ZN(
        P2_U3201) );
  AND3_X1 U15778 ( .A1(n13533), .A2(n13532), .A3(n11905), .ZN(n13534) );
  OAI21_X1 U15779 ( .B1(n13535), .B2(n13534), .A(n15123), .ZN(n13541) );
  INV_X1 U15780 ( .A(n13823), .ZN(n13539) );
  AND2_X1 U15781 ( .A1(n13679), .A2(n13701), .ZN(n13536) );
  AOI21_X1 U15782 ( .B1(n13684), .B2(n13555), .A(n13536), .ZN(n13956) );
  OAI22_X1 U15783 ( .A1(n13558), .A2(n13956), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13537), .ZN(n13538) );
  AOI21_X1 U15784 ( .B1(n13539), .B2(n13556), .A(n13538), .ZN(n13540) );
  OAI211_X1 U15785 ( .C1(n13958), .C2(n13542), .A(n13541), .B(n13540), .ZN(
        P2_U3205) );
  XNOR2_X1 U15786 ( .A(n13544), .B(n13543), .ZN(n13551) );
  NAND2_X1 U15787 ( .A1(n13679), .A2(n13555), .ZN(n13546) );
  NAND2_X1 U15788 ( .A1(n13672), .A2(n13701), .ZN(n13545) );
  AND2_X1 U15789 ( .A1(n13546), .A2(n13545), .ZN(n13970) );
  NAND2_X1 U15790 ( .A1(n13556), .A2(n13846), .ZN(n13548) );
  OAI211_X1 U15791 ( .C1(n13970), .C2(n13558), .A(n13548), .B(n13547), .ZN(
        n13549) );
  AOI21_X1 U15792 ( .B1(n13845), .B2(n15128), .A(n13549), .ZN(n13550) );
  OAI21_X1 U15793 ( .B1(n13551), .B2(n13561), .A(n13550), .ZN(P2_U3210) );
  AOI21_X1 U15794 ( .B1(n13553), .B2(n13552), .A(n6721), .ZN(n13562) );
  AND2_X1 U15795 ( .A1(n13688), .A2(n13701), .ZN(n13554) );
  AOI21_X1 U15796 ( .B1(n13694), .B2(n13555), .A(n13554), .ZN(n13919) );
  AOI22_X1 U15797 ( .A1(n13745), .A2(n13556), .B1(P2_REG3_REG_26__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13557) );
  OAI21_X1 U15798 ( .B1(n13919), .B2(n13558), .A(n13557), .ZN(n13559) );
  AOI21_X1 U15799 ( .B1(n13918), .B2(n15128), .A(n13559), .ZN(n13560) );
  OAI21_X1 U15800 ( .B1(n13562), .B2(n13561), .A(n13560), .ZN(P2_U3212) );
  MUX2_X1 U15801 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n13631), .S(n6666), .Z(
        P2_U3562) );
  MUX2_X1 U15802 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n13699), .S(n6666), .Z(
        P2_U3561) );
  MUX2_X1 U15803 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n13563), .S(n6666), .Z(
        P2_U3560) );
  MUX2_X1 U15804 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n13702), .S(P2_U3947), .Z(
        P2_U3559) );
  MUX2_X1 U15805 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n13694), .S(P2_U3947), .Z(
        P2_U3558) );
  MUX2_X1 U15806 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n13663), .S(P2_U3947), .Z(
        P2_U3557) );
  MUX2_X1 U15807 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n13688), .S(P2_U3947), .Z(
        P2_U3556) );
  MUX2_X1 U15808 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n13660), .S(P2_U3947), .Z(
        P2_U3555) );
  MUX2_X1 U15809 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(n13686), .S(P2_U3947), .Z(
        P2_U3554) );
  MUX2_X1 U15810 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n13656), .S(n6666), .Z(
        P2_U3553) );
  MUX2_X1 U15811 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n13684), .S(n6666), .Z(
        P2_U3552) );
  MUX2_X1 U15812 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n13680), .S(n6666), .Z(
        P2_U3551) );
  MUX2_X1 U15813 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n13679), .S(n6666), .Z(
        P2_U3550) );
  MUX2_X1 U15814 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n13675), .S(n6666), .Z(
        P2_U3549) );
  MUX2_X1 U15815 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n13672), .S(n6666), .Z(
        P2_U3548) );
  MUX2_X1 U15816 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n13670), .S(n6666), .Z(
        P2_U3547) );
  MUX2_X1 U15817 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n13643), .S(n6666), .Z(
        P2_U3546) );
  MUX2_X1 U15818 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n13564), .S(n6666), .Z(
        P2_U3545) );
  MUX2_X1 U15819 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n13565), .S(n6666), .Z(
        P2_U3544) );
  MUX2_X1 U15820 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n13566), .S(n6666), .Z(
        P2_U3543) );
  MUX2_X1 U15821 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n13567), .S(n6666), .Z(
        P2_U3542) );
  MUX2_X1 U15822 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n13568), .S(n6666), .Z(
        P2_U3541) );
  MUX2_X1 U15823 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n13569), .S(n6666), .Z(
        P2_U3540) );
  MUX2_X1 U15824 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n13570), .S(n6666), .Z(
        P2_U3539) );
  MUX2_X1 U15825 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n13571), .S(n6666), .Z(
        P2_U3538) );
  MUX2_X1 U15826 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n13572), .S(n6666), .Z(
        P2_U3537) );
  MUX2_X1 U15827 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(n13573), .S(n6666), .Z(
        P2_U3536) );
  MUX2_X1 U15828 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n13574), .S(n6666), .Z(
        P2_U3535) );
  MUX2_X1 U15829 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(n13575), .S(n6666), .Z(
        P2_U3534) );
  MUX2_X1 U15830 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(n13576), .S(n6666), .Z(
        P2_U3533) );
  MUX2_X1 U15831 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n13577), .S(n6666), .Z(
        P2_U3532) );
  MUX2_X1 U15832 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n13578), .S(n6666), .Z(
        P2_U3531) );
  MUX2_X1 U15833 ( .A(n10538), .B(P2_REG2_REG_7__SCAN_IN), .S(n13589), .Z(
        n13581) );
  INV_X1 U15834 ( .A(n13579), .ZN(n13580) );
  NAND2_X1 U15835 ( .A1(n13581), .A2(n13580), .ZN(n13583) );
  OAI211_X1 U15836 ( .C1(n15441), .C2(n13583), .A(n13582), .B(n15474), .ZN(
        n13596) );
  INV_X1 U15837 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n13585) );
  OAI21_X1 U15838 ( .B1(n15450), .B2(n13585), .A(n13584), .ZN(n13586) );
  AOI21_X1 U15839 ( .B1(n15453), .B2(n13589), .A(n13586), .ZN(n13595) );
  INV_X1 U15840 ( .A(n13587), .ZN(n15436) );
  INV_X1 U15841 ( .A(n13588), .ZN(n13591) );
  MUX2_X1 U15842 ( .A(n9487), .B(P2_REG1_REG_7__SCAN_IN), .S(n13589), .Z(
        n13590) );
  NAND3_X1 U15843 ( .A1(n15436), .A2(n13591), .A3(n13590), .ZN(n13592) );
  NAND3_X1 U15844 ( .A1(n15467), .A2(n13593), .A3(n13592), .ZN(n13594) );
  NAND3_X1 U15845 ( .A1(n13596), .A2(n13595), .A3(n13594), .ZN(P2_U3221) );
  NOR3_X1 U15846 ( .A1(n13602), .A2(n13597), .A3(n15442), .ZN(n13599) );
  NOR3_X1 U15847 ( .A1(n13606), .A2(n15571), .A3(n15459), .ZN(n13598) );
  OR3_X1 U15848 ( .A1(n13599), .A2(n15453), .A3(n13598), .ZN(n13604) );
  OAI21_X1 U15849 ( .B1(n13602), .B2(n13601), .A(n13600), .ZN(n13603) );
  AOI22_X1 U15850 ( .A1(n13604), .A2(n13605), .B1(n15474), .B2(n13603), .ZN(
        n13612) );
  NAND2_X1 U15851 ( .A1(n15472), .A2(P2_ADDR_REG_9__SCAN_IN), .ZN(n13610) );
  NOR3_X1 U15852 ( .A1(n13606), .A2(n13605), .A3(P2_REG1_REG_9__SCAN_IN), .ZN(
        n13608) );
  OAI21_X1 U15853 ( .B1(n13608), .B2(n13607), .A(n15467), .ZN(n13609) );
  NAND4_X1 U15854 ( .A1(n13612), .A2(n13611), .A3(n13610), .A4(n13609), .ZN(
        P2_U3223) );
  NOR2_X1 U15855 ( .A1(n13618), .A2(n13613), .ZN(n13614) );
  NOR2_X1 U15856 ( .A1(n13615), .A2(n13614), .ZN(n13616) );
  XOR2_X1 U15857 ( .A(n13616), .B(P2_REG2_REG_19__SCAN_IN), .Z(n13623) );
  NAND2_X1 U15858 ( .A1(n13618), .A2(n13617), .ZN(n13619) );
  NAND2_X1 U15859 ( .A1(n13620), .A2(n13619), .ZN(n13621) );
  XOR2_X1 U15860 ( .A(n13621), .B(P2_REG1_REG_19__SCAN_IN), .Z(n13622) );
  AOI22_X1 U15861 ( .A1(n13623), .A2(n15474), .B1(n15467), .B2(n13622), .ZN(
        n13625) );
  INV_X1 U15862 ( .A(n13622), .ZN(n13624) );
  INV_X1 U15863 ( .A(n13965), .ZN(n13835) );
  NAND2_X1 U15864 ( .A1(n13695), .A2(n13744), .ZN(n13730) );
  XNOR2_X1 U15865 ( .A(n13636), .B(n13632), .ZN(n13627) );
  NAND2_X1 U15866 ( .A1(n13627), .A2(n15144), .ZN(n13895) );
  NOR2_X1 U15867 ( .A1(n14029), .A2(n13628), .ZN(n13629) );
  NOR2_X1 U15868 ( .A1(n13630), .A2(n13629), .ZN(n13700) );
  NAND2_X1 U15869 ( .A1(n13631), .A2(n13700), .ZN(n13897) );
  NOR2_X1 U15870 ( .A1(n15151), .A2(n13897), .ZN(n13639) );
  INV_X1 U15871 ( .A(n13632), .ZN(n13896) );
  NOR2_X1 U15872 ( .A1(n13896), .A2(n13890), .ZN(n13633) );
  AOI211_X1 U15873 ( .C1(n15151), .C2(P2_REG2_REG_31__SCAN_IN), .A(n13639), 
        .B(n13633), .ZN(n13634) );
  OAI21_X1 U15874 ( .B1(n13895), .B2(n13870), .A(n13634), .ZN(P2_U3234) );
  INV_X1 U15875 ( .A(n13705), .ZN(n13637) );
  NOR2_X1 U15876 ( .A1(n13899), .A2(n13890), .ZN(n13638) );
  AOI211_X1 U15877 ( .C1(n15151), .C2(P2_REG2_REG_30__SCAN_IN), .A(n13639), 
        .B(n13638), .ZN(n13640) );
  OAI21_X1 U15878 ( .B1(n13870), .B2(n13898), .A(n13640), .ZN(P2_U3235) );
  OR2_X1 U15879 ( .A1(n13991), .A2(n13643), .ZN(n13644) );
  NAND2_X1 U15880 ( .A1(n13645), .A2(n13644), .ZN(n13879) );
  NAND2_X1 U15881 ( .A1(n13985), .A2(n13670), .ZN(n13646) );
  NAND2_X1 U15882 ( .A1(n13651), .A2(n13650), .ZN(n13818) );
  NAND2_X1 U15883 ( .A1(n13818), .A2(n13819), .ZN(n13653) );
  OR2_X1 U15884 ( .A1(n13681), .A2(n13680), .ZN(n13652) );
  NAND2_X1 U15885 ( .A1(n13653), .A2(n13652), .ZN(n13805) );
  NOR2_X1 U15886 ( .A1(n13953), .A2(n13684), .ZN(n13654) );
  NAND2_X1 U15887 ( .A1(n13953), .A2(n13684), .ZN(n13655) );
  AND2_X1 U15888 ( .A1(n13942), .A2(n13686), .ZN(n13657) );
  OR2_X1 U15889 ( .A1(n13782), .A2(n13657), .ZN(n13659) );
  OR2_X1 U15890 ( .A1(n13942), .A2(n13686), .ZN(n13658) );
  NAND2_X1 U15891 ( .A1(n13935), .A2(n13660), .ZN(n13661) );
  OR2_X1 U15892 ( .A1(n13927), .A2(n13688), .ZN(n13662) );
  NAND2_X1 U15893 ( .A1(n13918), .A2(n13663), .ZN(n13664) );
  OAI21_X1 U15894 ( .B1(n13695), .B2(n13665), .A(n13913), .ZN(n13719) );
  NAND2_X1 U15895 ( .A1(n13719), .A2(n13718), .ZN(n13717) );
  INV_X1 U15896 ( .A(n13672), .ZN(n13674) );
  INV_X1 U15897 ( .A(n13670), .ZN(n13671) );
  INV_X1 U15898 ( .A(n13845), .ZN(n13971) );
  INV_X1 U15899 ( .A(n13770), .ZN(n13772) );
  NAND2_X1 U15900 ( .A1(n13771), .A2(n13687), .ZN(n13757) );
  INV_X1 U15901 ( .A(n13753), .ZN(n13756) );
  NAND2_X1 U15902 ( .A1(n13757), .A2(n13756), .ZN(n13755) );
  INV_X1 U15903 ( .A(n13737), .ZN(n13692) );
  NAND2_X1 U15904 ( .A1(n13698), .A2(n15551), .ZN(n13704) );
  AOI22_X1 U15905 ( .A1(n13702), .A2(n13701), .B1(n13700), .B2(n13699), .ZN(
        n13703) );
  NAND2_X1 U15906 ( .A1(n13900), .A2(n13852), .ZN(n13713) );
  AOI21_X1 U15907 ( .B1(n13901), .B2(n13720), .A(n11865), .ZN(n13706) );
  NAND2_X1 U15908 ( .A1(n13706), .A2(n13705), .ZN(n13902) );
  INV_X1 U15909 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n13707) );
  OAI22_X1 U15910 ( .A1(n13708), .A2(n13865), .B1(n13707), .B2(n13852), .ZN(
        n13709) );
  AOI21_X1 U15911 ( .B1(n13901), .B2(n15139), .A(n13709), .ZN(n13710) );
  OAI21_X1 U15912 ( .B1(n13902), .B2(n13870), .A(n13710), .ZN(n13711) );
  INV_X1 U15913 ( .A(n13711), .ZN(n13712) );
  OAI211_X1 U15914 ( .C1(n13903), .C2(n13874), .A(n13713), .B(n13712), .ZN(
        P2_U3236) );
  AOI21_X1 U15915 ( .B1(n13714), .B2(n13718), .A(n15522), .ZN(n13716) );
  OAI21_X1 U15916 ( .B1(n13719), .B2(n13718), .A(n13717), .ZN(n13908) );
  INV_X1 U15917 ( .A(n13908), .ZN(n13727) );
  AOI21_X1 U15918 ( .B1(n13905), .B2(n13730), .A(n11865), .ZN(n13721) );
  NAND2_X1 U15919 ( .A1(n13904), .A2(n15147), .ZN(n13724) );
  AOI22_X1 U15920 ( .A1(n13722), .A2(n15137), .B1(P2_REG2_REG_28__SCAN_IN), 
        .B2(n15151), .ZN(n13723) );
  OAI211_X1 U15921 ( .C1(n13725), .C2(n13890), .A(n13724), .B(n13723), .ZN(
        n13726) );
  AOI21_X1 U15922 ( .B1(n13727), .B2(n15148), .A(n13726), .ZN(n13728) );
  OAI21_X1 U15923 ( .B1(n13907), .B2(n15151), .A(n13728), .ZN(P2_U3237) );
  XNOR2_X1 U15924 ( .A(n13729), .B(n13737), .ZN(n13917) );
  INV_X1 U15925 ( .A(n13744), .ZN(n13732) );
  INV_X1 U15926 ( .A(n13730), .ZN(n13731) );
  AOI211_X1 U15927 ( .C1(n13912), .C2(n13732), .A(n11865), .B(n13731), .ZN(
        n13910) );
  NAND2_X1 U15928 ( .A1(n13912), .A2(n15139), .ZN(n13735) );
  AOI22_X1 U15929 ( .A1(n13733), .A2(n15137), .B1(P2_REG2_REG_27__SCAN_IN), 
        .B2(n15151), .ZN(n13734) );
  OAI211_X1 U15930 ( .C1(n13909), .C2(n15151), .A(n13735), .B(n13734), .ZN(
        n13736) );
  AOI21_X1 U15931 ( .B1(n13910), .B2(n15147), .A(n13736), .ZN(n13740) );
  OR2_X1 U15932 ( .A1(n13738), .A2(n13737), .ZN(n13914) );
  NAND3_X1 U15933 ( .A1(n13914), .A2(n13913), .A3(n15148), .ZN(n13739) );
  OAI211_X1 U15934 ( .C1(n13917), .C2(n13859), .A(n13740), .B(n13739), .ZN(
        P2_U3238) );
  XNOR2_X1 U15935 ( .A(n13741), .B(n13749), .ZN(n13925) );
  NAND2_X1 U15936 ( .A1(n13918), .A2(n13760), .ZN(n13742) );
  NAND2_X1 U15937 ( .A1(n13742), .A2(n15144), .ZN(n13743) );
  NOR2_X1 U15938 ( .A1(n13744), .A2(n13743), .ZN(n13922) );
  NAND2_X1 U15939 ( .A1(n13918), .A2(n15139), .ZN(n13747) );
  AOI22_X1 U15940 ( .A1(n13745), .A2(n15137), .B1(P2_REG2_REG_26__SCAN_IN), 
        .B2(n15151), .ZN(n13746) );
  OAI211_X1 U15941 ( .C1(n15151), .C2(n13919), .A(n13747), .B(n13746), .ZN(
        n13748) );
  AOI21_X1 U15942 ( .B1(n13922), .B2(n15147), .A(n13748), .ZN(n13752) );
  XNOR2_X1 U15943 ( .A(n13750), .B(n13749), .ZN(n13923) );
  NAND2_X1 U15944 ( .A1(n13923), .A2(n15148), .ZN(n13751) );
  OAI211_X1 U15945 ( .C1(n13925), .C2(n13859), .A(n13752), .B(n13751), .ZN(
        P2_U3239) );
  XNOR2_X1 U15946 ( .A(n13754), .B(n13753), .ZN(n13930) );
  OAI21_X1 U15947 ( .B1(n13757), .B2(n13756), .A(n13755), .ZN(n13759) );
  AOI21_X1 U15948 ( .B1(n13759), .B2(n15551), .A(n13758), .ZN(n13929) );
  INV_X1 U15949 ( .A(n13929), .ZN(n13767) );
  AOI21_X1 U15950 ( .B1(n13927), .B2(n13774), .A(n11865), .ZN(n13761) );
  AND2_X1 U15951 ( .A1(n13761), .A2(n13760), .ZN(n13926) );
  NAND2_X1 U15952 ( .A1(n13926), .A2(n15147), .ZN(n13765) );
  INV_X1 U15953 ( .A(n13762), .ZN(n13763) );
  AOI22_X1 U15954 ( .A1(n13763), .A2(n15137), .B1(P2_REG2_REG_25__SCAN_IN), 
        .B2(n15151), .ZN(n13764) );
  OAI211_X1 U15955 ( .C1(n7449), .C2(n13890), .A(n13765), .B(n13764), .ZN(
        n13766) );
  AOI21_X1 U15956 ( .B1(n13767), .B2(n13852), .A(n13766), .ZN(n13768) );
  OAI21_X1 U15957 ( .B1(n13930), .B2(n13874), .A(n13768), .ZN(P2_U3240) );
  OAI21_X1 U15958 ( .B1(n6699), .B2(n13770), .A(n13769), .ZN(n13938) );
  OAI21_X1 U15959 ( .B1(n13773), .B2(n13772), .A(n13771), .ZN(n13931) );
  NAND2_X1 U15960 ( .A1(n13931), .A2(n13872), .ZN(n13781) );
  AOI21_X1 U15961 ( .B1(n13935), .B2(n6760), .A(n11865), .ZN(n13775) );
  AND2_X1 U15962 ( .A1(n13775), .A2(n13774), .ZN(n13933) );
  NAND2_X1 U15963 ( .A1(n13935), .A2(n15139), .ZN(n13778) );
  AOI22_X1 U15964 ( .A1(n15151), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n13776), 
        .B2(n15137), .ZN(n13777) );
  OAI211_X1 U15965 ( .C1(n15151), .C2(n13932), .A(n13778), .B(n13777), .ZN(
        n13779) );
  AOI21_X1 U15966 ( .B1(n13933), .B2(n15147), .A(n13779), .ZN(n13780) );
  OAI211_X1 U15967 ( .C1(n13938), .C2(n13874), .A(n13781), .B(n13780), .ZN(
        P2_U3241) );
  XNOR2_X1 U15968 ( .A(n13782), .B(n13783), .ZN(n13945) );
  XNOR2_X1 U15969 ( .A(n13784), .B(n13783), .ZN(n13939) );
  NAND2_X1 U15970 ( .A1(n13939), .A2(n13872), .ZN(n13792) );
  AOI21_X1 U15971 ( .B1(n13942), .B2(n13796), .A(n11865), .ZN(n13785) );
  AND2_X1 U15972 ( .A1(n13785), .A2(n6760), .ZN(n13940) );
  INV_X1 U15973 ( .A(n13941), .ZN(n13787) );
  OAI22_X1 U15974 ( .A1(n13787), .A2(n15151), .B1(n13786), .B2(n13865), .ZN(
        n13788) );
  AOI21_X1 U15975 ( .B1(P2_REG2_REG_23__SCAN_IN), .B2(n15151), .A(n13788), 
        .ZN(n13789) );
  OAI21_X1 U15976 ( .B1(n7451), .B2(n13890), .A(n13789), .ZN(n13790) );
  AOI21_X1 U15977 ( .B1(n15147), .B2(n13940), .A(n13790), .ZN(n13791) );
  OAI211_X1 U15978 ( .C1(n13945), .C2(n13874), .A(n13792), .B(n13791), .ZN(
        P2_U3242) );
  XOR2_X1 U15979 ( .A(n13800), .B(n13793), .Z(n13795) );
  AOI21_X1 U15980 ( .B1(n13795), .B2(n15551), .A(n13794), .ZN(n13949) );
  AOI211_X1 U15981 ( .C1(n13947), .C2(n13810), .A(n11865), .B(n7452), .ZN(
        n13946) );
  INV_X1 U15982 ( .A(n13797), .ZN(n13798) );
  AOI22_X1 U15983 ( .A1(n15151), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n13798), 
        .B2(n15137), .ZN(n13799) );
  OAI21_X1 U15984 ( .B1(n7233), .B2(n13890), .A(n13799), .ZN(n13803) );
  XNOR2_X1 U15985 ( .A(n13801), .B(n13800), .ZN(n13950) );
  NOR2_X1 U15986 ( .A1(n13950), .A2(n13874), .ZN(n13802) );
  AOI211_X1 U15987 ( .C1(n13946), .C2(n15147), .A(n13803), .B(n13802), .ZN(
        n13804) );
  OAI21_X1 U15988 ( .B1(n13949), .B2(n15151), .A(n13804), .ZN(P2_U3243) );
  XNOR2_X1 U15989 ( .A(n13805), .B(n13806), .ZN(n13955) );
  XNOR2_X1 U15990 ( .A(n13807), .B(n13806), .ZN(n13809) );
  OAI21_X1 U15991 ( .B1(n13809), .B2(n15522), .A(n13808), .ZN(n13951) );
  AOI21_X1 U15992 ( .B1(n13822), .B2(n13953), .A(n11865), .ZN(n13811) );
  AND2_X1 U15993 ( .A1(n13811), .A2(n13810), .ZN(n13952) );
  NAND2_X1 U15994 ( .A1(n13952), .A2(n15147), .ZN(n13814) );
  AOI22_X1 U15995 ( .A1(n15151), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n13812), 
        .B2(n15137), .ZN(n13813) );
  OAI211_X1 U15996 ( .C1(n13815), .C2(n13890), .A(n13814), .B(n13813), .ZN(
        n13816) );
  AOI21_X1 U15997 ( .B1(n13951), .B2(n13852), .A(n13816), .ZN(n13817) );
  OAI21_X1 U15998 ( .B1(n13874), .B2(n13955), .A(n13817), .ZN(P2_U3244) );
  XOR2_X1 U15999 ( .A(n13819), .B(n13818), .Z(n13962) );
  XNOR2_X1 U16000 ( .A(n13820), .B(n13819), .ZN(n13960) );
  INV_X1 U16001 ( .A(n13821), .ZN(n13830) );
  OAI211_X1 U16002 ( .C1(n13830), .C2(n13958), .A(n15144), .B(n13822), .ZN(
        n13957) );
  OAI22_X1 U16003 ( .A1(n15151), .A2(n13956), .B1(n13823), .B2(n13865), .ZN(
        n13825) );
  NOR2_X1 U16004 ( .A1(n13958), .A2(n13890), .ZN(n13824) );
  AOI211_X1 U16005 ( .C1(n15151), .C2(P2_REG2_REG_20__SCAN_IN), .A(n13825), 
        .B(n13824), .ZN(n13826) );
  OAI21_X1 U16006 ( .B1(n13870), .B2(n13957), .A(n13826), .ZN(n13827) );
  AOI21_X1 U16007 ( .B1(n13960), .B2(n13872), .A(n13827), .ZN(n13828) );
  OAI21_X1 U16008 ( .B1(n13874), .B2(n13962), .A(n13828), .ZN(P2_U3245) );
  XNOR2_X1 U16009 ( .A(n13829), .B(n13838), .ZN(n13969) );
  AOI211_X1 U16010 ( .C1(n13965), .C2(n6919), .A(n11865), .B(n13830), .ZN(
        n13963) );
  INV_X1 U16011 ( .A(n13964), .ZN(n13832) );
  OAI22_X1 U16012 ( .A1(n15151), .A2(n13832), .B1(n13831), .B2(n13865), .ZN(
        n13833) );
  AOI21_X1 U16013 ( .B1(P2_REG2_REG_19__SCAN_IN), .B2(n15151), .A(n13833), 
        .ZN(n13834) );
  OAI21_X1 U16014 ( .B1(n13835), .B2(n13890), .A(n13834), .ZN(n13836) );
  AOI21_X1 U16015 ( .B1(n13963), .B2(n15147), .A(n13836), .ZN(n13840) );
  XOR2_X1 U16016 ( .A(n13838), .B(n13837), .Z(n13966) );
  NAND2_X1 U16017 ( .A1(n13966), .A2(n15148), .ZN(n13839) );
  OAI211_X1 U16018 ( .C1(n13969), .C2(n13859), .A(n13840), .B(n13839), .ZN(
        P2_U3246) );
  XOR2_X1 U16019 ( .A(n13855), .B(n13841), .Z(n13976) );
  NAND2_X1 U16020 ( .A1(n13845), .A2(n13863), .ZN(n13842) );
  NAND2_X1 U16021 ( .A1(n13842), .A2(n15144), .ZN(n13843) );
  NOR2_X1 U16022 ( .A1(n13844), .A2(n13843), .ZN(n13973) );
  INV_X1 U16023 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n13851) );
  NAND2_X1 U16024 ( .A1(n13845), .A2(n15139), .ZN(n13850) );
  INV_X1 U16025 ( .A(n13846), .ZN(n13847) );
  OAI22_X1 U16026 ( .A1(n15151), .A2(n13970), .B1(n13847), .B2(n13865), .ZN(
        n13848) );
  INV_X1 U16027 ( .A(n13848), .ZN(n13849) );
  OAI211_X1 U16028 ( .C1(n13852), .C2(n13851), .A(n13850), .B(n13849), .ZN(
        n13853) );
  AOI21_X1 U16029 ( .B1(n13973), .B2(n15147), .A(n13853), .ZN(n13858) );
  OAI21_X1 U16030 ( .B1(n13856), .B2(n13855), .A(n13854), .ZN(n13974) );
  NAND2_X1 U16031 ( .A1(n13974), .A2(n15148), .ZN(n13857) );
  OAI211_X1 U16032 ( .C1(n13976), .C2(n13859), .A(n13858), .B(n13857), .ZN(
        P2_U3247) );
  XOR2_X1 U16033 ( .A(n13862), .B(n13860), .Z(n13983) );
  XOR2_X1 U16034 ( .A(n13862), .B(n13861), .Z(n13981) );
  OAI211_X1 U16035 ( .C1(n7448), .C2(n13979), .A(n15144), .B(n13863), .ZN(
        n13978) );
  INV_X1 U16036 ( .A(n13864), .ZN(n13866) );
  OAI22_X1 U16037 ( .A1(n15151), .A2(n13977), .B1(n13866), .B2(n13865), .ZN(
        n13868) );
  NOR2_X1 U16038 ( .A1(n13979), .A2(n13890), .ZN(n13867) );
  AOI211_X1 U16039 ( .C1(n15151), .C2(P2_REG2_REG_17__SCAN_IN), .A(n13868), 
        .B(n13867), .ZN(n13869) );
  OAI21_X1 U16040 ( .B1(n13870), .B2(n13978), .A(n13869), .ZN(n13871) );
  AOI21_X1 U16041 ( .B1(n13981), .B2(n13872), .A(n13871), .ZN(n13873) );
  OAI21_X1 U16042 ( .B1(n13983), .B2(n13874), .A(n13873), .ZN(P2_U3248) );
  XOR2_X1 U16043 ( .A(n13880), .B(n13875), .Z(n13878) );
  INV_X1 U16044 ( .A(n13876), .ZN(n13877) );
  AOI21_X1 U16045 ( .B1(n13878), .B2(n15551), .A(n13877), .ZN(n13987) );
  INV_X1 U16046 ( .A(n13879), .ZN(n13883) );
  INV_X1 U16047 ( .A(n13880), .ZN(n13882) );
  OAI21_X1 U16048 ( .B1(n13883), .B2(n13882), .A(n13881), .ZN(n13988) );
  INV_X1 U16049 ( .A(n13988), .ZN(n13893) );
  AOI21_X1 U16050 ( .B1(n13884), .B2(n13985), .A(n11865), .ZN(n13886) );
  AND2_X1 U16051 ( .A1(n13886), .A2(n13885), .ZN(n13984) );
  NAND2_X1 U16052 ( .A1(n13984), .A2(n15147), .ZN(n13889) );
  AOI22_X1 U16053 ( .A1(n15151), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n13887), 
        .B2(n15137), .ZN(n13888) );
  OAI211_X1 U16054 ( .C1(n13891), .C2(n13890), .A(n13889), .B(n13888), .ZN(
        n13892) );
  AOI21_X1 U16055 ( .B1(n13893), .B2(n15148), .A(n13892), .ZN(n13894) );
  OAI21_X1 U16056 ( .B1(n13987), .B2(n15151), .A(n13894), .ZN(P2_U3249) );
  OAI211_X1 U16057 ( .C1(n13896), .C2(n15548), .A(n13895), .B(n13897), .ZN(
        n14000) );
  MUX2_X1 U16058 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n14000), .S(n15158), .Z(
        P2_U3530) );
  MUX2_X1 U16059 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n14001), .S(n15576), .Z(
        P2_U3529) );
  AOI21_X1 U16060 ( .B1(n15539), .B2(n13905), .A(n13904), .ZN(n13906) );
  OAI211_X1 U16061 ( .C1(n13998), .C2(n13908), .A(n13907), .B(n13906), .ZN(
        n14002) );
  MUX2_X1 U16062 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n14002), .S(n15158), .Z(
        P2_U3527) );
  INV_X1 U16063 ( .A(n13909), .ZN(n13911) );
  AOI211_X1 U16064 ( .C1(n15539), .C2(n13912), .A(n13911), .B(n13910), .ZN(
        n13916) );
  NAND3_X1 U16065 ( .A1(n13914), .A2(n13913), .A3(n15527), .ZN(n13915) );
  OAI211_X1 U16066 ( .C1(n13917), .C2(n15522), .A(n13916), .B(n13915), .ZN(
        n14003) );
  MUX2_X1 U16067 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n14003), .S(n15158), .Z(
        P2_U3526) );
  INV_X1 U16068 ( .A(n13918), .ZN(n13920) );
  OAI21_X1 U16069 ( .B1(n13920), .B2(n15548), .A(n13919), .ZN(n13921) );
  AOI211_X1 U16070 ( .C1(n13923), .C2(n15527), .A(n13922), .B(n13921), .ZN(
        n13924) );
  OAI21_X1 U16071 ( .B1(n13925), .B2(n15522), .A(n13924), .ZN(n14004) );
  MUX2_X1 U16072 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n14004), .S(n15158), .Z(
        P2_U3525) );
  AOI21_X1 U16073 ( .B1(n15539), .B2(n13927), .A(n13926), .ZN(n13928) );
  OAI211_X1 U16074 ( .C1(n13998), .C2(n13930), .A(n13929), .B(n13928), .ZN(
        n14005) );
  MUX2_X1 U16075 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n14005), .S(n15158), .Z(
        P2_U3524) );
  NAND2_X1 U16076 ( .A1(n13931), .A2(n15551), .ZN(n13937) );
  INV_X1 U16077 ( .A(n13932), .ZN(n13934) );
  AOI211_X1 U16078 ( .C1(n15539), .C2(n13935), .A(n13934), .B(n13933), .ZN(
        n13936) );
  OAI211_X1 U16079 ( .C1(n13998), .C2(n13938), .A(n13937), .B(n13936), .ZN(
        n14006) );
  MUX2_X1 U16080 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n14006), .S(n15158), .Z(
        P2_U3523) );
  NAND2_X1 U16081 ( .A1(n13939), .A2(n15551), .ZN(n13944) );
  AOI211_X1 U16082 ( .C1(n15539), .C2(n13942), .A(n13941), .B(n13940), .ZN(
        n13943) );
  OAI211_X1 U16083 ( .C1(n13998), .C2(n13945), .A(n13944), .B(n13943), .ZN(
        n14007) );
  MUX2_X1 U16084 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n14007), .S(n15158), .Z(
        P2_U3522) );
  AOI21_X1 U16085 ( .B1(n15539), .B2(n13947), .A(n13946), .ZN(n13948) );
  OAI211_X1 U16086 ( .C1(n13998), .C2(n13950), .A(n13949), .B(n13948), .ZN(
        n14008) );
  MUX2_X1 U16087 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n14008), .S(n15158), .Z(
        P2_U3521) );
  AOI211_X1 U16088 ( .C1(n15539), .C2(n13953), .A(n13952), .B(n13951), .ZN(
        n13954) );
  OAI21_X1 U16089 ( .B1(n13998), .B2(n13955), .A(n13954), .ZN(n14009) );
  MUX2_X1 U16090 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n14009), .S(n15158), .Z(
        P2_U3520) );
  OAI211_X1 U16091 ( .C1(n13958), .C2(n15548), .A(n13957), .B(n13956), .ZN(
        n13959) );
  AOI21_X1 U16092 ( .B1(n13960), .B2(n15551), .A(n13959), .ZN(n13961) );
  OAI21_X1 U16093 ( .B1(n13998), .B2(n13962), .A(n13961), .ZN(n14010) );
  MUX2_X1 U16094 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n14010), .S(n15158), .Z(
        P2_U3519) );
  AOI211_X1 U16095 ( .C1(n15539), .C2(n13965), .A(n13964), .B(n13963), .ZN(
        n13968) );
  NAND2_X1 U16096 ( .A1(n13966), .A2(n15527), .ZN(n13967) );
  OAI211_X1 U16097 ( .C1(n13969), .C2(n15522), .A(n13968), .B(n13967), .ZN(
        n14011) );
  MUX2_X1 U16098 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n14011), .S(n15158), .Z(
        P2_U3518) );
  OAI21_X1 U16099 ( .B1(n13971), .B2(n15548), .A(n13970), .ZN(n13972) );
  AOI211_X1 U16100 ( .C1(n13974), .C2(n15527), .A(n13973), .B(n13972), .ZN(
        n13975) );
  OAI21_X1 U16101 ( .B1(n13976), .B2(n15522), .A(n13975), .ZN(n14012) );
  MUX2_X1 U16102 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n14012), .S(n15158), .Z(
        P2_U3517) );
  OAI211_X1 U16103 ( .C1(n13979), .C2(n15548), .A(n13978), .B(n13977), .ZN(
        n13980) );
  AOI21_X1 U16104 ( .B1(n13981), .B2(n15551), .A(n13980), .ZN(n13982) );
  OAI21_X1 U16105 ( .B1(n13998), .B2(n13983), .A(n13982), .ZN(n14013) );
  MUX2_X1 U16106 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n14013), .S(n15158), .Z(
        P2_U3516) );
  AOI21_X1 U16107 ( .B1(n15539), .B2(n13985), .A(n13984), .ZN(n13986) );
  OAI211_X1 U16108 ( .C1(n13998), .C2(n13988), .A(n13987), .B(n13986), .ZN(
        n14014) );
  MUX2_X1 U16109 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n14014), .S(n15158), .Z(
        P2_U3515) );
  AOI211_X1 U16110 ( .C1(n15539), .C2(n13991), .A(n13990), .B(n13989), .ZN(
        n13992) );
  OAI21_X1 U16111 ( .B1(n13998), .B2(n13993), .A(n13992), .ZN(n14015) );
  MUX2_X1 U16112 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n14015), .S(n15158), .Z(
        P2_U3514) );
  AOI211_X1 U16113 ( .C1(n15539), .C2(n15127), .A(n13995), .B(n13994), .ZN(
        n13996) );
  OAI21_X1 U16114 ( .B1(n13998), .B2(n13997), .A(n13996), .ZN(n14016) );
  MUX2_X1 U16115 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n14016), .S(n15576), .Z(
        P2_U3513) );
  MUX2_X1 U16116 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n13999), .S(n15576), .Z(
        P2_U3503) );
  MUX2_X1 U16117 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n14000), .S(n15561), .Z(
        P2_U3498) );
  MUX2_X1 U16118 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n14002), .S(n15561), .Z(
        P2_U3495) );
  MUX2_X1 U16119 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n14003), .S(n15561), .Z(
        P2_U3494) );
  MUX2_X1 U16120 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n14004), .S(n15561), .Z(
        P2_U3493) );
  MUX2_X1 U16121 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n14005), .S(n15561), .Z(
        P2_U3492) );
  MUX2_X1 U16122 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n14006), .S(n15561), .Z(
        P2_U3491) );
  MUX2_X1 U16123 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n14007), .S(n15561), .Z(
        P2_U3490) );
  MUX2_X1 U16124 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n14008), .S(n15561), .Z(
        P2_U3489) );
  MUX2_X1 U16125 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n14009), .S(n15561), .Z(
        P2_U3488) );
  MUX2_X1 U16126 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n14010), .S(n15561), .Z(
        P2_U3487) );
  MUX2_X1 U16127 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n14011), .S(n15561), .Z(
        P2_U3486) );
  MUX2_X1 U16128 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n14012), .S(n15561), .Z(
        P2_U3484) );
  MUX2_X1 U16129 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n14013), .S(n15561), .Z(
        P2_U3481) );
  MUX2_X1 U16130 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n14014), .S(n15561), .Z(
        P2_U3478) );
  MUX2_X1 U16131 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n14015), .S(n15561), .Z(
        P2_U3475) );
  MUX2_X1 U16132 ( .A(P2_REG0_REG_14__SCAN_IN), .B(n14016), .S(n15561), .Z(
        P2_U3472) );
  INV_X1 U16133 ( .A(n14017), .ZN(n14799) );
  NOR4_X1 U16134 ( .A1(n8505), .A2(P2_IR_REG_30__SCAN_IN), .A3(n14018), .A4(
        P2_U3088), .ZN(n14019) );
  AOI21_X1 U16135 ( .B1(P1_DATAO_REG_31__SCAN_IN), .B2(n14026), .A(n14019), 
        .ZN(n14020) );
  OAI21_X1 U16136 ( .B1(n14799), .B2(n14031), .A(n14020), .ZN(P2_U3296) );
  INV_X1 U16137 ( .A(n14021), .ZN(n14805) );
  OAI222_X1 U16138 ( .A1(n14031), .A2(n14805), .B1(n14023), .B2(P2_U3088), 
        .C1(n14022), .C2(n14038), .ZN(P2_U3298) );
  INV_X1 U16139 ( .A(n14024), .ZN(n14808) );
  AOI21_X1 U16140 ( .B1(n14026), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n14025), 
        .ZN(n14027) );
  OAI21_X1 U16141 ( .B1(n14808), .B2(n14031), .A(n14027), .ZN(P2_U3299) );
  OAI222_X1 U16142 ( .A1(n14031), .A2(n14030), .B1(n14029), .B2(P2_U3088), 
        .C1(n14028), .C2(n14038), .ZN(P2_U3300) );
  INV_X1 U16143 ( .A(n14032), .ZN(n14811) );
  OAI222_X1 U16144 ( .A1(n14038), .A2(n14034), .B1(n14033), .B2(P2_U3088), 
        .C1(n14031), .C2(n14811), .ZN(P2_U3301) );
  INV_X1 U16145 ( .A(n14035), .ZN(n14814) );
  OAI222_X1 U16146 ( .A1(n14038), .A2(n14037), .B1(n14031), .B2(n14814), .C1(
        P2_U3088), .C2(n14036), .ZN(P2_U3302) );
  INV_X1 U16147 ( .A(n14039), .ZN(n14040) );
  MUX2_X1 U16148 ( .A(n14040), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3327) );
  OAI21_X1 U16149 ( .B1(n14043), .B2(n14042), .A(n14041), .ZN(n14044) );
  NAND2_X1 U16150 ( .A1(n14044), .A2(n14195), .ZN(n14048) );
  AOI22_X1 U16151 ( .A1(n14966), .A2(n14687), .B1(n14444), .B2(n15378), .ZN(
        n14474) );
  INV_X1 U16152 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n14045) );
  OAI22_X1 U16153 ( .A1(n14474), .A2(n14200), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14045), .ZN(n14046) );
  AOI21_X1 U16154 ( .B1(n14208), .B2(n14479), .A(n14046), .ZN(n14047) );
  OAI211_X1 U16155 ( .C1(n7519), .C2(n14191), .A(n14048), .B(n14047), .ZN(
        P1_U3214) );
  INV_X1 U16156 ( .A(n14730), .ZN(n14404) );
  INV_X1 U16157 ( .A(n14134), .ZN(n14052) );
  NOR3_X1 U16158 ( .A1(n14165), .A2(n14050), .A3(n14049), .ZN(n14051) );
  OAI21_X1 U16159 ( .B1(n14052), .B2(n14051), .A(n14195), .ZN(n14056) );
  AOI22_X1 U16160 ( .A1(n14207), .A2(n14541), .B1(P1_REG3_REG_23__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14053) );
  OAI21_X1 U16161 ( .B1(n14543), .B2(n15161), .A(n14053), .ZN(n14054) );
  AOI21_X1 U16162 ( .B1(n14544), .B2(n14208), .A(n14054), .ZN(n14055) );
  OAI211_X1 U16163 ( .C1(n14404), .C2(n14191), .A(n14056), .B(n14055), .ZN(
        P1_U3216) );
  AOI21_X1 U16164 ( .B1(n14058), .B2(n14057), .A(n15167), .ZN(n14060) );
  NAND2_X1 U16165 ( .A1(n14060), .A2(n14059), .ZN(n14067) );
  NAND2_X1 U16166 ( .A1(P1_U3086), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n14262) );
  OAI21_X1 U16167 ( .B1(n15164), .B2(n14061), .A(n14262), .ZN(n14062) );
  AOI21_X1 U16168 ( .B1(n14063), .B2(n6659), .A(n14062), .ZN(n14066) );
  AOI22_X1 U16169 ( .A1(n15172), .A2(n14064), .B1(n14208), .B2(n9987), .ZN(
        n14065) );
  NAND3_X1 U16170 ( .A1(n14067), .A2(n14066), .A3(n14065), .ZN(P1_U3218) );
  XNOR2_X1 U16171 ( .A(n14069), .B(n14068), .ZN(n14184) );
  NAND2_X1 U16172 ( .A1(n14183), .A2(n14184), .ZN(n14182) );
  AND2_X1 U16173 ( .A1(n14182), .A2(n14072), .ZN(n14074) );
  XOR2_X1 U16174 ( .A(n14071), .B(n14070), .Z(n14073) );
  NAND3_X1 U16175 ( .A1(n14182), .A2(n14073), .A3(n14072), .ZN(n14142) );
  OAI211_X1 U16176 ( .C1(n14074), .C2(n14073), .A(n14195), .B(n14142), .ZN(
        n14078) );
  NAND2_X1 U16177 ( .A1(n14570), .A2(n14207), .ZN(n14075) );
  NAND2_X1 U16178 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n14379)
         );
  OAI211_X1 U16179 ( .C1(n14608), .C2(n15161), .A(n14075), .B(n14379), .ZN(
        n14076) );
  AOI21_X1 U16180 ( .B1(n14610), .B2(n14208), .A(n14076), .ZN(n14077) );
  OAI211_X1 U16181 ( .C1(n14381), .C2(n14191), .A(n14078), .B(n14077), .ZN(
        P1_U3219) );
  INV_X1 U16182 ( .A(n14743), .ZN(n14575) );
  OAI21_X1 U16183 ( .B1(n14080), .B2(n14079), .A(n14163), .ZN(n14081) );
  NAND2_X1 U16184 ( .A1(n14081), .A2(n14195), .ZN(n14086) );
  INV_X1 U16185 ( .A(n14082), .ZN(n14573) );
  AOI22_X1 U16186 ( .A1(n14569), .A2(n14207), .B1(P1_REG3_REG_21__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14083) );
  OAI21_X1 U16187 ( .B1(n14606), .B2(n15161), .A(n14083), .ZN(n14084) );
  AOI21_X1 U16188 ( .B1(n14573), .B2(n14208), .A(n14084), .ZN(n14085) );
  OAI211_X1 U16189 ( .C1(n14575), .C2(n14191), .A(n14086), .B(n14085), .ZN(
        P1_U3223) );
  AND2_X1 U16190 ( .A1(n14172), .A2(n14087), .ZN(n14090) );
  OAI211_X1 U16191 ( .C1(n14090), .C2(n14089), .A(n14195), .B(n14088), .ZN(
        n14097) );
  AOI21_X1 U16192 ( .B1(n14207), .B2(n14218), .A(n14091), .ZN(n14092) );
  OAI21_X1 U16193 ( .B1(n14093), .B2(n15161), .A(n14092), .ZN(n14094) );
  AOI21_X1 U16194 ( .B1(n14095), .B2(n14208), .A(n14094), .ZN(n14096) );
  OAI211_X1 U16195 ( .C1(n14098), .C2(n14191), .A(n14097), .B(n14096), .ZN(
        P1_U3224) );
  INV_X1 U16196 ( .A(n14514), .ZN(n14717) );
  INV_X1 U16197 ( .A(n14099), .ZN(n14103) );
  NOR3_X1 U16198 ( .A1(n14136), .A2(n14101), .A3(n14100), .ZN(n14102) );
  OAI21_X1 U16199 ( .B1(n14103), .B2(n14102), .A(n14195), .ZN(n14109) );
  NAND2_X1 U16200 ( .A1(n14541), .A2(n15378), .ZN(n14105) );
  NAND2_X1 U16201 ( .A1(n14444), .A2(n14966), .ZN(n14104) );
  AND2_X1 U16202 ( .A1(n14105), .A2(n14104), .ZN(n14715) );
  OAI22_X1 U16203 ( .A1(n14715), .A2(n14200), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14106), .ZN(n14107) );
  AOI21_X1 U16204 ( .B1(n14508), .B2(n14208), .A(n14107), .ZN(n14108) );
  OAI211_X1 U16205 ( .C1(n14717), .C2(n14191), .A(n14109), .B(n14108), .ZN(
        P1_U3225) );
  AOI21_X1 U16206 ( .B1(n14112), .B2(n14111), .A(n14110), .ZN(n14121) );
  NAND2_X1 U16207 ( .A1(n14427), .A2(n14966), .ZN(n14114) );
  NAND2_X1 U16208 ( .A1(n14421), .A2(n15378), .ZN(n14113) );
  NAND2_X1 U16209 ( .A1(n14114), .A2(n14113), .ZN(n14772) );
  NAND2_X1 U16210 ( .A1(n14772), .A2(n14115), .ZN(n14117) );
  OAI211_X1 U16211 ( .C1(n15176), .C2(n14118), .A(n14117), .B(n14116), .ZN(
        n14119) );
  AOI21_X1 U16212 ( .B1(n14773), .B2(n15172), .A(n14119), .ZN(n14120) );
  OAI21_X1 U16213 ( .B1(n14121), .B2(n15167), .A(n14120), .ZN(P1_U3226) );
  INV_X1 U16214 ( .A(n14769), .ZN(n14641) );
  INV_X1 U16215 ( .A(n14122), .ZN(n14126) );
  NOR3_X1 U16216 ( .A1(n14110), .A2(n14124), .A3(n14123), .ZN(n14125) );
  OAI21_X1 U16217 ( .B1(n14126), .B2(n14125), .A(n14195), .ZN(n14131) );
  NAND2_X1 U16218 ( .A1(n14217), .A2(n14966), .ZN(n14128) );
  NAND2_X1 U16219 ( .A1(n14665), .A2(n15378), .ZN(n14127) );
  AND2_X1 U16220 ( .A1(n14128), .A2(n14127), .ZN(n14634) );
  NAND2_X1 U16221 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n14358)
         );
  OAI21_X1 U16222 ( .B1(n14634), .B2(n14200), .A(n14358), .ZN(n14129) );
  AOI21_X1 U16223 ( .B1(n14638), .B2(n14208), .A(n14129), .ZN(n14130) );
  OAI211_X1 U16224 ( .C1(n14641), .C2(n14191), .A(n14131), .B(n14130), .ZN(
        P1_U3228) );
  INV_X1 U16225 ( .A(n14724), .ZN(n14532) );
  AND3_X1 U16226 ( .A1(n14134), .A2(n14133), .A3(n14132), .ZN(n14135) );
  OAI21_X1 U16227 ( .B1(n14136), .B2(n14135), .A(n14195), .ZN(n14140) );
  AOI22_X1 U16228 ( .A1(n14966), .A2(n14443), .B1(n14440), .B2(n15378), .ZN(
        n14520) );
  INV_X1 U16229 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n14137) );
  OAI22_X1 U16230 ( .A1(n14520), .A2(n14200), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14137), .ZN(n14138) );
  AOI21_X1 U16231 ( .B1(n14529), .B2(n14208), .A(n14138), .ZN(n14139) );
  OAI211_X1 U16232 ( .C1(n14532), .C2(n14191), .A(n14140), .B(n14139), .ZN(
        P1_U3229) );
  NAND2_X1 U16233 ( .A1(n14142), .A2(n14141), .ZN(n14143) );
  XOR2_X1 U16234 ( .A(n14144), .B(n14143), .Z(n14150) );
  NOR2_X1 U16235 ( .A1(n15176), .A2(n14589), .ZN(n14148) );
  AOI22_X1 U16236 ( .A1(n14588), .A2(n14207), .B1(P1_REG3_REG_20__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14145) );
  OAI21_X1 U16237 ( .B1(n14146), .B2(n15161), .A(n14145), .ZN(n14147) );
  AOI211_X1 U16238 ( .C1(n14400), .C2(n15172), .A(n14148), .B(n14147), .ZN(
        n14149) );
  OAI21_X1 U16239 ( .B1(n14150), .B2(n15167), .A(n14149), .ZN(P1_U3233) );
  XNOR2_X1 U16240 ( .A(n14152), .B(n14151), .ZN(n14158) );
  NOR2_X1 U16241 ( .A1(n15176), .A2(n14987), .ZN(n14156) );
  NAND2_X1 U16242 ( .A1(n14207), .A2(n14967), .ZN(n14154) );
  OAI211_X1 U16243 ( .C1(n15213), .C2(n15161), .A(n14154), .B(n14153), .ZN(
        n14155) );
  AOI211_X1 U16244 ( .C1(n15216), .C2(n15172), .A(n14156), .B(n14155), .ZN(
        n14157) );
  OAI21_X1 U16245 ( .B1(n14158), .B2(n15167), .A(n14157), .ZN(P1_U3234) );
  INV_X1 U16246 ( .A(n14159), .ZN(n14204) );
  NAND2_X1 U16247 ( .A1(n14160), .A2(n15379), .ZN(n14738) );
  AND3_X1 U16248 ( .A1(n14163), .A2(n14162), .A3(n14161), .ZN(n14164) );
  OAI21_X1 U16249 ( .B1(n14165), .B2(n14164), .A(n14195), .ZN(n14171) );
  NAND2_X1 U16250 ( .A1(n14588), .A2(n15378), .ZN(n14167) );
  NAND2_X1 U16251 ( .A1(n14440), .A2(n14966), .ZN(n14166) );
  AND2_X1 U16252 ( .A1(n14167), .A2(n14166), .ZN(n14739) );
  OAI22_X1 U16253 ( .A1(n14739), .A2(n14200), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14168), .ZN(n14169) );
  AOI21_X1 U16254 ( .B1(n14557), .B2(n14208), .A(n14169), .ZN(n14170) );
  OAI211_X1 U16255 ( .C1(n14204), .C2(n14738), .A(n14171), .B(n14170), .ZN(
        P1_U3235) );
  INV_X1 U16256 ( .A(n15183), .ZN(n15224) );
  OAI21_X1 U16257 ( .B1(n14174), .B2(n14173), .A(n14172), .ZN(n14175) );
  NAND2_X1 U16258 ( .A1(n14175), .A2(n14195), .ZN(n14181) );
  NAND2_X1 U16259 ( .A1(n14221), .A2(n15378), .ZN(n14177) );
  NAND2_X1 U16260 ( .A1(n14219), .A2(n14966), .ZN(n14176) );
  AND2_X1 U16261 ( .A1(n14177), .A2(n14176), .ZN(n15180) );
  OAI21_X1 U16262 ( .B1(n15180), .B2(n14200), .A(n14178), .ZN(n14179) );
  AOI21_X1 U16263 ( .B1(n15182), .B2(n14208), .A(n14179), .ZN(n14180) );
  OAI211_X1 U16264 ( .C1(n15224), .C2(n14191), .A(n14181), .B(n14180), .ZN(
        P1_U3236) );
  INV_X1 U16265 ( .A(n14762), .ZN(n14620) );
  OAI21_X1 U16266 ( .B1(n14184), .B2(n14183), .A(n14182), .ZN(n14185) );
  NAND2_X1 U16267 ( .A1(n14185), .A2(n14195), .ZN(n14190) );
  NAND2_X1 U16268 ( .A1(n14427), .A2(n15378), .ZN(n14187) );
  NAND2_X1 U16269 ( .A1(n14587), .A2(n14966), .ZN(n14186) );
  AND2_X1 U16270 ( .A1(n14187), .A2(n14186), .ZN(n14624) );
  NAND2_X1 U16271 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n15269)
         );
  OAI21_X1 U16272 ( .B1(n14624), .B2(n14200), .A(n15269), .ZN(n14188) );
  AOI21_X1 U16273 ( .B1(n14618), .B2(n14208), .A(n14188), .ZN(n14189) );
  OAI211_X1 U16274 ( .C1(n14620), .C2(n14191), .A(n14190), .B(n14189), .ZN(
        P1_U3238) );
  NAND2_X1 U16275 ( .A1(n14499), .A2(n15379), .ZN(n14709) );
  OAI21_X1 U16276 ( .B1(n14194), .B2(n14193), .A(n14192), .ZN(n14196) );
  NAND2_X1 U16277 ( .A1(n14196), .A2(n14195), .ZN(n14203) );
  NAND2_X1 U16278 ( .A1(n14447), .A2(n14966), .ZN(n14198) );
  NAND2_X1 U16279 ( .A1(n14443), .A2(n15378), .ZN(n14197) );
  AND2_X1 U16280 ( .A1(n14198), .A2(n14197), .ZN(n14711) );
  OAI22_X1 U16281 ( .A1(n14711), .A2(n14200), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14199), .ZN(n14201) );
  AOI21_X1 U16282 ( .B1(n14495), .B2(n14208), .A(n14201), .ZN(n14202) );
  OAI211_X1 U16283 ( .C1(n14709), .C2(n14204), .A(n14203), .B(n14202), .ZN(
        P1_U3240) );
  XNOR2_X1 U16284 ( .A(n14206), .B(n14205), .ZN(n14214) );
  AOI22_X1 U16285 ( .A1(n14207), .A2(n14665), .B1(P1_REG3_REG_15__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14210) );
  NAND2_X1 U16286 ( .A1(n14208), .A2(n14671), .ZN(n14209) );
  OAI211_X1 U16287 ( .C1(n14211), .C2(n15161), .A(n14210), .B(n14209), .ZN(
        n14212) );
  AOI21_X1 U16288 ( .B1(n14672), .B2(n15172), .A(n14212), .ZN(n14213) );
  OAI21_X1 U16289 ( .B1(n14214), .B2(n15167), .A(n14213), .ZN(P1_U3241) );
  MUX2_X1 U16290 ( .A(n14386), .B(P1_DATAO_REG_31__SCAN_IN), .S(n14215), .Z(
        P1_U3591) );
  MUX2_X1 U16291 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n14216), .S(P1_U4016), .Z(
        P1_U3589) );
  MUX2_X1 U16292 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n14687), .S(P1_U4016), .Z(
        P1_U3588) );
  MUX2_X1 U16293 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n14447), .S(P1_U4016), .Z(
        P1_U3587) );
  MUX2_X1 U16294 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n14444), .S(P1_U4016), .Z(
        P1_U3586) );
  MUX2_X1 U16295 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n14443), .S(P1_U4016), .Z(
        P1_U3585) );
  MUX2_X1 U16296 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n14541), .S(P1_U4016), .Z(
        P1_U3584) );
  MUX2_X1 U16297 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n14440), .S(P1_U4016), .Z(
        P1_U3583) );
  MUX2_X1 U16298 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n14569), .S(P1_U4016), .Z(
        P1_U3582) );
  MUX2_X1 U16299 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n14588), .S(P1_U4016), .Z(
        P1_U3581) );
  MUX2_X1 U16300 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n14570), .S(P1_U4016), .Z(
        P1_U3580) );
  MUX2_X1 U16301 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n14587), .S(P1_U4016), .Z(
        P1_U3579) );
  MUX2_X1 U16302 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n14217), .S(P1_U4016), .Z(
        P1_U3578) );
  MUX2_X1 U16303 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n14427), .S(P1_U4016), .Z(
        P1_U3577) );
  MUX2_X1 U16304 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n14665), .S(P1_U4016), .Z(
        P1_U3576) );
  MUX2_X1 U16305 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n14421), .S(P1_U4016), .Z(
        P1_U3575) );
  MUX2_X1 U16306 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n14967), .S(P1_U4016), .Z(
        P1_U3574) );
  MUX2_X1 U16307 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n14218), .S(P1_U4016), .Z(
        P1_U3573) );
  MUX2_X1 U16308 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n14219), .S(P1_U4016), .Z(
        P1_U3572) );
  MUX2_X1 U16309 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n14220), .S(P1_U4016), .Z(
        P1_U3571) );
  MUX2_X1 U16310 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n14221), .S(P1_U4016), .Z(
        P1_U3570) );
  MUX2_X1 U16311 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n15377), .S(P1_U4016), .Z(
        P1_U3569) );
  MUX2_X1 U16312 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n14222), .S(P1_U4016), .Z(
        P1_U3568) );
  MUX2_X1 U16313 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n14223), .S(P1_U4016), .Z(
        P1_U3567) );
  MUX2_X1 U16314 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n14224), .S(P1_U4016), .Z(
        P1_U3566) );
  MUX2_X1 U16315 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n14225), .S(P1_U4016), .Z(
        P1_U3565) );
  MUX2_X1 U16316 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n14226), .S(P1_U4016), .Z(
        P1_U3564) );
  MUX2_X1 U16317 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n14227), .S(P1_U4016), .Z(
        P1_U3563) );
  MUX2_X1 U16318 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n6659), .S(P1_U4016), .Z(
        P1_U3562) );
  MUX2_X1 U16319 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n14229), .S(P1_U4016), .Z(
        P1_U3561) );
  MUX2_X1 U16320 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n14230), .S(P1_U4016), .Z(
        P1_U3560) );
  OAI22_X1 U16321 ( .A1(n15271), .A2(n14232), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14231), .ZN(n14233) );
  AOI21_X1 U16322 ( .B1(n14234), .B2(n14340), .A(n14233), .ZN(n14243) );
  INV_X1 U16323 ( .A(n14235), .ZN(n14238) );
  OAI21_X1 U16324 ( .B1(n9709), .B2(n14247), .A(n14236), .ZN(n14237) );
  NAND3_X1 U16325 ( .A1(n14378), .A2(n14238), .A3(n14237), .ZN(n14242) );
  NAND2_X1 U16326 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n14245) );
  OAI211_X1 U16327 ( .C1(n9729), .C2(n14240), .A(n14377), .B(n14239), .ZN(
        n14241) );
  NAND3_X1 U16328 ( .A1(n14243), .A2(n14242), .A3(n14241), .ZN(P1_U3244) );
  MUX2_X1 U16329 ( .A(n14246), .B(n14245), .S(n6667), .Z(n14250) );
  NAND2_X1 U16330 ( .A1(n14248), .A2(n14247), .ZN(n14249) );
  OAI211_X1 U16331 ( .C1(n14250), .C2(n14807), .A(P1_U4016), .B(n14249), .ZN(
        n14292) );
  AOI22_X1 U16332 ( .A1(n14360), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n14261) );
  XNOR2_X1 U16333 ( .A(n14252), .B(n14251), .ZN(n14257) );
  AOI211_X1 U16334 ( .C1(n14255), .C2(n14254), .A(n14253), .B(n15264), .ZN(
        n14256) );
  AOI21_X1 U16335 ( .B1(n14377), .B2(n14257), .A(n14256), .ZN(n14260) );
  NAND2_X1 U16336 ( .A1(n14340), .A2(n14258), .ZN(n14259) );
  NAND4_X1 U16337 ( .A1(n14292), .A2(n14261), .A3(n14260), .A4(n14259), .ZN(
        P1_U3245) );
  INV_X1 U16338 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n14263) );
  OAI21_X1 U16339 ( .B1(n15271), .B2(n14263), .A(n14262), .ZN(n14264) );
  AOI21_X1 U16340 ( .B1(n14265), .B2(n14340), .A(n14264), .ZN(n14274) );
  OAI211_X1 U16341 ( .C1(n14267), .C2(n14266), .A(n14377), .B(n14287), .ZN(
        n14273) );
  NAND3_X1 U16342 ( .A1(n14270), .A2(n14269), .A3(n14268), .ZN(n14271) );
  NAND3_X1 U16343 ( .A1(n14378), .A2(n6947), .A3(n14271), .ZN(n14272) );
  NAND3_X1 U16344 ( .A1(n14274), .A2(n14273), .A3(n14272), .ZN(P1_U3246) );
  NOR2_X1 U16345 ( .A1(n15267), .A2(n14275), .ZN(n14276) );
  AOI211_X1 U16346 ( .C1(n14360), .C2(P1_ADDR_REG_4__SCAN_IN), .A(n14277), .B(
        n14276), .ZN(n14291) );
  MUX2_X1 U16347 ( .A(n9711), .B(P1_REG1_REG_4__SCAN_IN), .S(n14284), .Z(
        n14280) );
  INV_X1 U16348 ( .A(n14278), .ZN(n14279) );
  NAND2_X1 U16349 ( .A1(n14280), .A2(n14279), .ZN(n14282) );
  OAI211_X1 U16350 ( .C1(n14283), .C2(n14282), .A(n14378), .B(n14281), .ZN(
        n14290) );
  MUX2_X1 U16351 ( .A(n9734), .B(P1_REG2_REG_4__SCAN_IN), .S(n14284), .Z(
        n14285) );
  NAND3_X1 U16352 ( .A1(n14287), .A2(n14286), .A3(n14285), .ZN(n14288) );
  NAND3_X1 U16353 ( .A1(n14377), .A2(n14302), .A3(n14288), .ZN(n14289) );
  NAND4_X1 U16354 ( .A1(n14292), .A2(n14291), .A3(n14290), .A4(n14289), .ZN(
        P1_U3247) );
  OAI21_X1 U16355 ( .B1(n15271), .B2(n14867), .A(n14293), .ZN(n14294) );
  AOI21_X1 U16356 ( .B1(n14299), .B2(n14340), .A(n14294), .ZN(n14307) );
  OAI21_X1 U16357 ( .B1(n14297), .B2(n14296), .A(n14295), .ZN(n14298) );
  NAND2_X1 U16358 ( .A1(n14298), .A2(n14378), .ZN(n14306) );
  MUX2_X1 U16359 ( .A(n9737), .B(P1_REG2_REG_5__SCAN_IN), .S(n14299), .Z(
        n14300) );
  NAND3_X1 U16360 ( .A1(n14302), .A2(n14301), .A3(n14300), .ZN(n14303) );
  NAND3_X1 U16361 ( .A1(n14377), .A2(n14304), .A3(n14303), .ZN(n14305) );
  NAND3_X1 U16362 ( .A1(n14307), .A2(n14306), .A3(n14305), .ZN(P1_U3248) );
  INV_X1 U16363 ( .A(n14308), .ZN(n14310) );
  MUX2_X1 U16364 ( .A(n15396), .B(P1_REG1_REG_7__SCAN_IN), .S(n14317), .Z(
        n14309) );
  NAND2_X1 U16365 ( .A1(n14310), .A2(n14309), .ZN(n14312) );
  OAI211_X1 U16366 ( .C1(n14313), .C2(n14312), .A(n14311), .B(n14378), .ZN(
        n14325) );
  INV_X1 U16367 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n14315) );
  OAI21_X1 U16368 ( .B1(n15271), .B2(n14315), .A(n14314), .ZN(n14316) );
  AOI21_X1 U16369 ( .B1(n14317), .B2(n14340), .A(n14316), .ZN(n14324) );
  MUX2_X1 U16370 ( .A(n9742), .B(P1_REG2_REG_7__SCAN_IN), .S(n14317), .Z(
        n14318) );
  NAND3_X1 U16371 ( .A1(n14320), .A2(n14319), .A3(n14318), .ZN(n14321) );
  NAND3_X1 U16372 ( .A1(n14377), .A2(n14322), .A3(n14321), .ZN(n14323) );
  NAND3_X1 U16373 ( .A1(n14325), .A2(n14324), .A3(n14323), .ZN(P1_U3250) );
  INV_X1 U16374 ( .A(n14326), .ZN(n14331) );
  NOR3_X1 U16375 ( .A1(n14329), .A2(n14328), .A3(n14327), .ZN(n14330) );
  OAI21_X1 U16376 ( .B1(n14331), .B2(n14330), .A(n14378), .ZN(n14344) );
  NOR2_X1 U16377 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n14332), .ZN(n14333) );
  AOI21_X1 U16378 ( .B1(n14360), .B2(P1_ADDR_REG_9__SCAN_IN), .A(n14333), .ZN(
        n14343) );
  MUX2_X1 U16379 ( .A(n9843), .B(P1_REG2_REG_9__SCAN_IN), .S(n14339), .Z(
        n14334) );
  NAND3_X1 U16380 ( .A1(n14336), .A2(n14335), .A3(n14334), .ZN(n14337) );
  NAND3_X1 U16381 ( .A1(n14377), .A2(n14338), .A3(n14337), .ZN(n14342) );
  NAND2_X1 U16382 ( .A1(n14340), .A2(n14339), .ZN(n14341) );
  NAND4_X1 U16383 ( .A1(n14344), .A2(n14343), .A3(n14342), .A4(n14341), .ZN(
        P1_U3252) );
  NAND2_X1 U16384 ( .A1(n14346), .A2(n14345), .ZN(n14351) );
  INV_X1 U16385 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n14349) );
  NAND2_X1 U16386 ( .A1(n14347), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n14370) );
  INV_X1 U16387 ( .A(n14370), .ZN(n14348) );
  AOI21_X1 U16388 ( .B1(n14349), .B2(n14364), .A(n14348), .ZN(n14350) );
  NAND2_X1 U16389 ( .A1(n14350), .A2(n14351), .ZN(n14369) );
  OAI211_X1 U16390 ( .C1(n14351), .C2(n14350), .A(n14377), .B(n14369), .ZN(
        n14362) );
  XNOR2_X1 U16391 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n14364), .ZN(n14356) );
  INV_X1 U16392 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n14354) );
  OAI211_X1 U16393 ( .C1(n14356), .C2(n14355), .A(n14363), .B(n14378), .ZN(
        n14357) );
  NAND2_X1 U16394 ( .A1(n14358), .A2(n14357), .ZN(n14359) );
  AOI21_X1 U16395 ( .B1(n14360), .B2(P1_ADDR_REG_17__SCAN_IN), .A(n14359), 
        .ZN(n14361) );
  OAI211_X1 U16396 ( .C1(n15267), .C2(n14364), .A(n14362), .B(n14361), .ZN(
        P1_U3260) );
  INV_X1 U16397 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n14365) );
  NAND2_X1 U16398 ( .A1(n14372), .A2(n14366), .ZN(n14367) );
  NAND2_X1 U16399 ( .A1(n15261), .A2(n14367), .ZN(n14368) );
  NAND2_X1 U16400 ( .A1(n14370), .A2(n14369), .ZN(n14371) );
  NAND2_X1 U16401 ( .A1(n14372), .A2(n14371), .ZN(n14373) );
  XOR2_X1 U16402 ( .A(n14372), .B(n14371), .Z(n15260) );
  NAND2_X1 U16403 ( .A1(P1_REG2_REG_18__SCAN_IN), .A2(n15260), .ZN(n15259) );
  NAND2_X1 U16404 ( .A1(n14373), .A2(n15259), .ZN(n14374) );
  XOR2_X1 U16405 ( .A(P1_REG2_REG_19__SCAN_IN), .B(n14374), .Z(n14376) );
  OAI21_X1 U16406 ( .B1(n14376), .B2(n15266), .A(n15267), .ZN(n14375) );
  OAI211_X1 U16407 ( .C1(n8002), .C2(n15271), .A(n14380), .B(n14379), .ZN(
        P1_U3262) );
  INV_X1 U16408 ( .A(n14672), .ZN(n15195) );
  AND2_X2 U16409 ( .A1(n14668), .A2(n15195), .ZN(n14670) );
  INV_X1 U16410 ( .A(n14773), .ZN(n14651) );
  NAND2_X1 U16411 ( .A1(n14609), .A2(n14749), .ZN(n14586) );
  OR2_X2 U16412 ( .A1(n14514), .A2(n14527), .ZN(n14506) );
  NOR2_X1 U16413 ( .A1(n14415), .A2(n14682), .ZN(n14382) );
  XOR2_X1 U16414 ( .A(n14382), .B(n14679), .Z(n14681) );
  INV_X1 U16415 ( .A(P1_B_REG_SCAN_IN), .ZN(n14383) );
  OR2_X1 U16416 ( .A1(n6668), .A2(n14383), .ZN(n14384) );
  NAND2_X1 U16417 ( .A1(n14966), .A2(n14384), .ZN(n14407) );
  INV_X1 U16418 ( .A(n14407), .ZN(n14385) );
  NAND2_X1 U16419 ( .A1(n14386), .A2(n14385), .ZN(n14683) );
  NOR2_X1 U16420 ( .A1(n6665), .A2(n14683), .ZN(n14391) );
  AOI21_X1 U16421 ( .B1(n6665), .B2(P1_REG2_REG_31__SCAN_IN), .A(n14391), .ZN(
        n14388) );
  NAND2_X1 U16422 ( .A1(n14679), .A2(n15282), .ZN(n14387) );
  OAI211_X1 U16423 ( .C1(n14681), .C2(n14675), .A(n14388), .B(n14387), .ZN(
        P1_U3263) );
  XOR2_X1 U16424 ( .A(n14415), .B(n14682), .Z(n14389) );
  NAND2_X1 U16425 ( .A1(n14389), .A2(n15288), .ZN(n14684) );
  AND2_X1 U16426 ( .A1(n6665), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n14390) );
  NOR2_X1 U16427 ( .A1(n14391), .A2(n14390), .ZN(n14393) );
  NAND2_X1 U16428 ( .A1(n14682), .A2(n15282), .ZN(n14392) );
  OAI211_X1 U16429 ( .C1(n14684), .C2(n14550), .A(n14393), .B(n14392), .ZN(
        P1_U3264) );
  INV_X1 U16430 ( .A(n14665), .ZN(n14395) );
  NAND2_X1 U16431 ( .A1(n14633), .A2(n14632), .ZN(n14631) );
  NAND2_X1 U16432 ( .A1(n14631), .A2(n14396), .ZN(n14623) );
  INV_X1 U16433 ( .A(n14398), .ZN(n14399) );
  INV_X1 U16434 ( .A(n14588), .ZN(n14401) );
  INV_X1 U16435 ( .A(n14499), .ZN(n14406) );
  AOI22_X2 U16436 ( .A1(n14473), .A2(n14484), .B1(n14456), .B2(n14705), .ZN(
        n14455) );
  NOR2_X1 U16437 ( .A1(n14408), .A2(n14407), .ZN(n14686) );
  INV_X1 U16438 ( .A(n14409), .ZN(n14411) );
  AOI22_X1 U16439 ( .A1(n14686), .A2(n14411), .B1(n14410), .B2(n15293), .ZN(
        n14413) );
  NAND2_X1 U16440 ( .A1(n6665), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n14412) );
  OAI211_X1 U16441 ( .C1(n14414), .C2(n14978), .A(n14413), .B(n14412), .ZN(
        n14418) );
  AOI21_X1 U16442 ( .B1(n14419), .B2(n14461), .A(n15320), .ZN(n14416) );
  NAND2_X1 U16443 ( .A1(n14416), .A2(n14415), .ZN(n14689) );
  NOR2_X1 U16444 ( .A1(n14689), .A2(n14550), .ZN(n14417) );
  AOI211_X1 U16445 ( .C1(n15282), .C2(n14419), .A(n14418), .B(n14417), .ZN(
        n14453) );
  NAND2_X1 U16446 ( .A1(n15203), .A2(n14967), .ZN(n14420) );
  OR2_X1 U16447 ( .A1(n14672), .A2(n14421), .ZN(n14422) );
  INV_X1 U16448 ( .A(n14645), .ZN(n14423) );
  OR2_X1 U16449 ( .A1(n14773), .A2(n14665), .ZN(n14424) );
  NOR2_X1 U16450 ( .A1(n14769), .A2(n14427), .ZN(n14426) );
  NAND2_X1 U16451 ( .A1(n14769), .A2(n14427), .ZN(n14428) );
  INV_X1 U16452 ( .A(n14430), .ZN(n14431) );
  OR2_X1 U16453 ( .A1(n14759), .A2(n14587), .ZN(n14433) );
  NAND2_X1 U16454 ( .A1(n14434), .A2(n14433), .ZN(n14596) );
  OR2_X1 U16455 ( .A1(n14749), .A2(n14606), .ZN(n14436) );
  OR2_X1 U16456 ( .A1(n14743), .A2(n14588), .ZN(n14437) );
  NAND2_X1 U16457 ( .A1(n14559), .A2(n14543), .ZN(n14438) );
  NAND2_X1 U16458 ( .A1(n14439), .A2(n14438), .ZN(n14540) );
  NAND2_X1 U16459 ( .A1(n14730), .A2(n14440), .ZN(n14523) );
  OR2_X1 U16460 ( .A1(n14724), .A2(n14541), .ZN(n14442) );
  NAND2_X1 U16461 ( .A1(n14499), .A2(n14444), .ZN(n14445) );
  INV_X1 U16462 ( .A(n14484), .ZN(n14446) );
  OR2_X1 U16463 ( .A1(n14705), .A2(n14447), .ZN(n14448) );
  AND2_X2 U16464 ( .A1(n14481), .A2(n14448), .ZN(n14464) );
  NAND2_X1 U16465 ( .A1(n14692), .A2(n15191), .ZN(n14452) );
  OAI211_X1 U16466 ( .C1(n14694), .C2(n14599), .A(n14453), .B(n14452), .ZN(
        P1_U3356) );
  NOR2_X1 U16467 ( .A1(n14457), .A2(n14607), .ZN(n14458) );
  AOI21_X1 U16468 ( .B1(n14468), .B2(n14477), .A(n15320), .ZN(n14462) );
  NAND2_X1 U16469 ( .A1(n14462), .A2(n14461), .ZN(n14698) );
  NAND3_X1 U16470 ( .A1(n14697), .A2(n15191), .A3(n14696), .ZN(n14470) );
  NAND2_X1 U16471 ( .A1(n6665), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n14465) );
  OAI21_X1 U16472 ( .B1(n14986), .B2(n14466), .A(n14465), .ZN(n14467) );
  AOI21_X1 U16473 ( .B1(n14468), .B2(n15282), .A(n14467), .ZN(n14469) );
  OAI211_X1 U16474 ( .C1(n14550), .C2(n14698), .A(n14470), .B(n14469), .ZN(
        n14471) );
  AOI21_X1 U16475 ( .B1(n14695), .B2(n14969), .A(n14471), .ZN(n14472) );
  INV_X1 U16476 ( .A(n14472), .ZN(P1_U3265) );
  XNOR2_X1 U16477 ( .A(n14473), .B(n14484), .ZN(n14476) );
  INV_X1 U16478 ( .A(n14474), .ZN(n14475) );
  AOI21_X1 U16479 ( .B1(n14476), .B2(n15375), .A(n14475), .ZN(n14707) );
  INV_X1 U16480 ( .A(n14477), .ZN(n14478) );
  AOI211_X1 U16481 ( .C1(n14705), .C2(n14489), .A(n15320), .B(n14478), .ZN(
        n14704) );
  AOI22_X1 U16482 ( .A1(n6665), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n15293), 
        .B2(n14479), .ZN(n14480) );
  OAI21_X1 U16483 ( .B1(n7519), .B2(n15297), .A(n14480), .ZN(n14486) );
  INV_X1 U16484 ( .A(n14481), .ZN(n14482) );
  AOI21_X1 U16485 ( .B1(n14484), .B2(n14483), .A(n14482), .ZN(n14708) );
  NOR2_X1 U16486 ( .A1(n14708), .A2(n14982), .ZN(n14485) );
  AOI211_X1 U16487 ( .C1(n14704), .C2(n15299), .A(n14486), .B(n14485), .ZN(
        n14487) );
  OAI21_X1 U16488 ( .B1(n14707), .B2(n6665), .A(n14487), .ZN(P1_U3266) );
  XNOR2_X1 U16489 ( .A(n14488), .B(n14491), .ZN(n14714) );
  AOI21_X1 U16490 ( .B1(n14499), .B2(n14506), .A(n15320), .ZN(n14490) );
  NAND2_X1 U16491 ( .A1(n14490), .A2(n14489), .ZN(n14710) );
  XNOR2_X1 U16492 ( .A(n14492), .B(n14491), .ZN(n14493) );
  NAND2_X1 U16493 ( .A1(n14493), .A2(n15375), .ZN(n14712) );
  OAI211_X1 U16494 ( .C1(n14612), .C2(n14710), .A(n14712), .B(n14711), .ZN(
        n14494) );
  NAND2_X1 U16495 ( .A1(n14494), .A2(n14969), .ZN(n14501) );
  INV_X1 U16496 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n14497) );
  INV_X1 U16497 ( .A(n14495), .ZN(n14496) );
  OAI22_X1 U16498 ( .A1(n14969), .A2(n14497), .B1(n14496), .B2(n14986), .ZN(
        n14498) );
  AOI21_X1 U16499 ( .B1(n14499), .B2(n15282), .A(n14498), .ZN(n14500) );
  OAI211_X1 U16500 ( .C1(n14714), .C2(n14982), .A(n14501), .B(n14500), .ZN(
        P1_U3267) );
  XNOR2_X1 U16501 ( .A(n6765), .B(n14503), .ZN(n14721) );
  OAI21_X1 U16502 ( .B1(n14504), .B2(n14503), .A(n14502), .ZN(n14505) );
  INV_X1 U16503 ( .A(n14505), .ZN(n14719) );
  AOI21_X1 U16504 ( .B1(n14514), .B2(n14527), .A(n15320), .ZN(n14507) );
  NAND2_X1 U16505 ( .A1(n14507), .A2(n14506), .ZN(n14716) );
  INV_X1 U16506 ( .A(n14508), .ZN(n14509) );
  OAI21_X1 U16507 ( .B1(n14509), .B2(n14986), .A(n14715), .ZN(n14510) );
  NAND2_X1 U16508 ( .A1(n14510), .A2(n14969), .ZN(n14512) );
  NAND2_X1 U16509 ( .A1(n6665), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n14511) );
  NAND2_X1 U16510 ( .A1(n14512), .A2(n14511), .ZN(n14513) );
  AOI21_X1 U16511 ( .B1(n14514), .B2(n15282), .A(n14513), .ZN(n14515) );
  OAI21_X1 U16512 ( .B1(n14716), .B2(n14550), .A(n14515), .ZN(n14516) );
  AOI21_X1 U16513 ( .B1(n14719), .B2(n15191), .A(n14516), .ZN(n14517) );
  OAI21_X1 U16514 ( .B1(n14721), .B2(n14599), .A(n14517), .ZN(P1_U3268) );
  AOI211_X1 U16515 ( .C1(n14525), .C2(n14519), .A(n15351), .B(n14518), .ZN(
        n14522) );
  INV_X1 U16516 ( .A(n14520), .ZN(n14521) );
  NOR2_X1 U16517 ( .A1(n14522), .A2(n14521), .ZN(n14726) );
  AND2_X1 U16518 ( .A1(n14732), .A2(n14523), .ZN(n14526) );
  OAI21_X1 U16519 ( .B1(n14526), .B2(n14525), .A(n14524), .ZN(n14722) );
  INV_X1 U16520 ( .A(n14527), .ZN(n14528) );
  AOI211_X1 U16521 ( .C1(n14724), .C2(n14537), .A(n15320), .B(n14528), .ZN(
        n14723) );
  NAND2_X1 U16522 ( .A1(n14723), .A2(n15299), .ZN(n14531) );
  AOI22_X1 U16523 ( .A1(n6665), .A2(P1_REG2_REG_24__SCAN_IN), .B1(n14529), 
        .B2(n15293), .ZN(n14530) );
  OAI211_X1 U16524 ( .C1(n14532), .C2(n15297), .A(n14531), .B(n14530), .ZN(
        n14533) );
  AOI21_X1 U16525 ( .B1(n14722), .B2(n15191), .A(n14533), .ZN(n14534) );
  OAI21_X1 U16526 ( .B1(n14726), .B2(n6665), .A(n14534), .ZN(P1_U3269) );
  XNOR2_X1 U16527 ( .A(n14536), .B(n14535), .ZN(n14728) );
  AOI21_X1 U16528 ( .B1(n14730), .B2(n14555), .A(n15320), .ZN(n14538) );
  NAND2_X1 U16529 ( .A1(n14538), .A2(n14537), .ZN(n14733) );
  NAND2_X1 U16530 ( .A1(n14540), .A2(n14539), .ZN(n14731) );
  NAND3_X1 U16531 ( .A1(n14732), .A2(n14731), .A3(n15191), .ZN(n14549) );
  NAND2_X1 U16532 ( .A1(n14541), .A2(n14966), .ZN(n14542) );
  OAI21_X1 U16533 ( .B1(n14543), .B2(n15212), .A(n14542), .ZN(n14729) );
  NAND2_X1 U16534 ( .A1(n14729), .A2(n14969), .ZN(n14546) );
  AOI22_X1 U16535 ( .A1(n6665), .A2(P1_REG2_REG_23__SCAN_IN), .B1(n14544), 
        .B2(n15293), .ZN(n14545) );
  NAND2_X1 U16536 ( .A1(n14546), .A2(n14545), .ZN(n14547) );
  AOI21_X1 U16537 ( .B1(n14730), .B2(n15282), .A(n14547), .ZN(n14548) );
  OAI211_X1 U16538 ( .C1(n14733), .C2(n14550), .A(n14549), .B(n14548), .ZN(
        n14551) );
  AOI21_X1 U16539 ( .B1(n14728), .B2(n14654), .A(n14551), .ZN(n14552) );
  INV_X1 U16540 ( .A(n14552), .ZN(P1_U3270) );
  XNOR2_X1 U16541 ( .A(n14554), .B(n14553), .ZN(n14742) );
  OAI211_X1 U16542 ( .C1(n14559), .C2(n14556), .A(n15288), .B(n14555), .ZN(
        n14737) );
  INV_X1 U16543 ( .A(n14737), .ZN(n14565) );
  AOI22_X1 U16544 ( .A1(n6665), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n14557), 
        .B2(n15293), .ZN(n14558) );
  OAI21_X1 U16545 ( .B1(n14559), .B2(n15297), .A(n14558), .ZN(n14564) );
  AOI21_X1 U16546 ( .B1(n14561), .B2(n14560), .A(n6736), .ZN(n14562) );
  OR2_X1 U16547 ( .A1(n14562), .A2(n15351), .ZN(n14740) );
  AOI21_X1 U16548 ( .B1(n14740), .B2(n14739), .A(n6665), .ZN(n14563) );
  AOI211_X1 U16549 ( .C1(n14565), .C2(n15299), .A(n14564), .B(n14563), .ZN(
        n14566) );
  OAI21_X1 U16550 ( .B1(n14742), .B2(n14982), .A(n14566), .ZN(P1_U3271) );
  OAI211_X1 U16551 ( .C1(n14568), .C2(n14579), .A(n14567), .B(n15375), .ZN(
        n14572) );
  AOI22_X1 U16552 ( .A1(n14570), .A2(n15378), .B1(n14569), .B2(n14966), .ZN(
        n14571) );
  AND2_X1 U16553 ( .A1(n14572), .A2(n14571), .ZN(n14746) );
  XNOR2_X1 U16554 ( .A(n14575), .B(n14586), .ZN(n14744) );
  AOI22_X1 U16555 ( .A1(n6665), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n14573), 
        .B2(n15293), .ZN(n14574) );
  OAI21_X1 U16556 ( .B1(n14575), .B2(n15297), .A(n14574), .ZN(n14581) );
  INV_X1 U16557 ( .A(n14576), .ZN(n14577) );
  AOI21_X1 U16558 ( .B1(n14579), .B2(n14578), .A(n14577), .ZN(n14747) );
  NOR2_X1 U16559 ( .A1(n14747), .A2(n14982), .ZN(n14580) );
  AOI211_X1 U16560 ( .C1(n14744), .C2(n14628), .A(n14581), .B(n14580), .ZN(
        n14582) );
  OAI21_X1 U16561 ( .B1(n6665), .B2(n14746), .A(n14582), .ZN(P1_U3272) );
  OAI21_X1 U16562 ( .B1(n14584), .B2(n14595), .A(n14583), .ZN(n14756) );
  OR2_X1 U16563 ( .A1(n14609), .A2(n14749), .ZN(n14585) );
  AND2_X1 U16564 ( .A1(n14586), .A2(n14585), .ZN(n14751) );
  AOI22_X1 U16565 ( .A1(n14588), .A2(n14966), .B1(n14587), .B2(n15378), .ZN(
        n14748) );
  NOR2_X1 U16566 ( .A1(n14986), .A2(n14589), .ZN(n14590) );
  AOI21_X1 U16567 ( .B1(n6665), .B2(P1_REG2_REG_20__SCAN_IN), .A(n14590), .ZN(
        n14591) );
  OAI21_X1 U16568 ( .B1(n14748), .B2(n6665), .A(n14591), .ZN(n14592) );
  INV_X1 U16569 ( .A(n14592), .ZN(n14593) );
  OAI21_X1 U16570 ( .B1(n14749), .B2(n15297), .A(n14593), .ZN(n14594) );
  AOI21_X1 U16571 ( .B1(n14751), .B2(n14628), .A(n14594), .ZN(n14598) );
  NAND2_X1 U16572 ( .A1(n14596), .A2(n14595), .ZN(n14752) );
  NAND3_X1 U16573 ( .A1(n14753), .A2(n14752), .A3(n15191), .ZN(n14597) );
  OAI211_X1 U16574 ( .C1(n14756), .C2(n14599), .A(n14598), .B(n14597), .ZN(
        P1_U3273) );
  XNOR2_X1 U16575 ( .A(n14601), .B(n14600), .ZN(n14761) );
  AOI21_X1 U16576 ( .B1(n14604), .B2(n14603), .A(n14602), .ZN(n14605) );
  OAI222_X1 U16577 ( .A1(n15212), .A2(n14608), .B1(n14607), .B2(n14606), .C1(
        n15351), .C2(n14605), .ZN(n14757) );
  AOI211_X1 U16578 ( .C1(n14759), .C2(n6790), .A(n15320), .B(n14609), .ZN(
        n14758) );
  INV_X1 U16579 ( .A(n14758), .ZN(n14613) );
  INV_X1 U16580 ( .A(n14610), .ZN(n14611) );
  OAI22_X1 U16581 ( .A1(n14613), .A2(n14612), .B1(n14986), .B2(n14611), .ZN(
        n14614) );
  OAI21_X1 U16582 ( .B1(n14757), .B2(n14614), .A(n14969), .ZN(n14616) );
  AOI22_X1 U16583 ( .A1(n14759), .A2(n15282), .B1(n6665), .B2(
        P1_REG2_REG_19__SCAN_IN), .ZN(n14615) );
  OAI211_X1 U16584 ( .C1(n14761), .C2(n14982), .A(n14616), .B(n14615), .ZN(
        P1_U3274) );
  XOR2_X1 U16585 ( .A(n14617), .B(n14622), .Z(n14766) );
  XNOR2_X1 U16586 ( .A(n14636), .B(n14620), .ZN(n14763) );
  AOI22_X1 U16587 ( .A1(n6665), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n14618), 
        .B2(n15293), .ZN(n14619) );
  OAI21_X1 U16588 ( .B1(n14620), .B2(n15297), .A(n14619), .ZN(n14627) );
  OAI211_X1 U16589 ( .C1(n14623), .C2(n14622), .A(n14621), .B(n15375), .ZN(
        n14625) );
  NOR2_X1 U16590 ( .A1(n14765), .A2(n6665), .ZN(n14626) );
  AOI211_X1 U16591 ( .C1(n14763), .C2(n14628), .A(n14627), .B(n14626), .ZN(
        n14629) );
  OAI21_X1 U16592 ( .B1(n14982), .B2(n14766), .A(n14629), .ZN(P1_U3275) );
  XNOR2_X1 U16593 ( .A(n14630), .B(n14632), .ZN(n14771) );
  OAI211_X1 U16594 ( .C1(n14633), .C2(n14632), .A(n14631), .B(n15375), .ZN(
        n14635) );
  NAND2_X1 U16595 ( .A1(n14635), .A2(n14634), .ZN(n14767) );
  INV_X1 U16596 ( .A(n14636), .ZN(n14637) );
  AOI211_X1 U16597 ( .C1(n14769), .C2(n14647), .A(n15320), .B(n14637), .ZN(
        n14768) );
  NAND2_X1 U16598 ( .A1(n14768), .A2(n15299), .ZN(n14640) );
  AOI22_X1 U16599 ( .A1(n6665), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n14638), 
        .B2(n15293), .ZN(n14639) );
  OAI211_X1 U16600 ( .C1(n14641), .C2(n15297), .A(n14640), .B(n14639), .ZN(
        n14642) );
  AOI21_X1 U16601 ( .B1(n14767), .B2(n14969), .A(n14642), .ZN(n14643) );
  OAI21_X1 U16602 ( .B1(n14982), .B2(n14771), .A(n14643), .ZN(P1_U3276) );
  XNOR2_X1 U16603 ( .A(n14644), .B(n14645), .ZN(n14779) );
  XNOR2_X1 U16604 ( .A(n14646), .B(n14645), .ZN(n14777) );
  OAI21_X1 U16605 ( .B1(n14670), .B2(n14651), .A(n14647), .ZN(n14775) );
  NOR2_X1 U16606 ( .A1(n14775), .A2(n14675), .ZN(n14653) );
  AOI22_X1 U16607 ( .A1(n6665), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n14648), 
        .B2(n15293), .ZN(n14650) );
  NAND2_X1 U16608 ( .A1(n14969), .A2(n14772), .ZN(n14649) );
  OAI211_X1 U16609 ( .C1(n14651), .C2(n15297), .A(n14650), .B(n14649), .ZN(
        n14652) );
  AOI211_X1 U16610 ( .C1(n14777), .C2(n14654), .A(n14653), .B(n14652), .ZN(
        n14655) );
  OAI21_X1 U16611 ( .B1(n14982), .B2(n14779), .A(n14655), .ZN(P1_U3277) );
  NAND2_X1 U16612 ( .A1(n14656), .A2(n7476), .ZN(n14657) );
  NAND2_X1 U16613 ( .A1(n14658), .A2(n14657), .ZN(n15194) );
  INV_X1 U16614 ( .A(n15194), .ZN(n14678) );
  NAND3_X1 U16615 ( .A1(n14661), .A2(n14660), .A3(n14659), .ZN(n14662) );
  NAND2_X1 U16616 ( .A1(n14662), .A2(n15375), .ZN(n14663) );
  OR2_X1 U16617 ( .A1(n14664), .A2(n14663), .ZN(n14667) );
  AOI22_X1 U16618 ( .A1(n14966), .A2(n14665), .B1(n14967), .B2(n15378), .ZN(
        n14666) );
  NAND2_X1 U16619 ( .A1(n14667), .A2(n14666), .ZN(n15199) );
  NOR2_X1 U16620 ( .A1(n14668), .A2(n15195), .ZN(n14669) );
  OR2_X1 U16621 ( .A1(n14670), .A2(n14669), .ZN(n15196) );
  AOI22_X1 U16622 ( .A1(n6665), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n14671), 
        .B2(n15293), .ZN(n14674) );
  NAND2_X1 U16623 ( .A1(n14672), .A2(n15282), .ZN(n14673) );
  OAI211_X1 U16624 ( .C1(n15196), .C2(n14675), .A(n14674), .B(n14673), .ZN(
        n14676) );
  AOI21_X1 U16625 ( .B1(n15199), .B2(n14969), .A(n14676), .ZN(n14677) );
  OAI21_X1 U16626 ( .B1(n14678), .B2(n14982), .A(n14677), .ZN(P1_U3278) );
  NAND2_X1 U16627 ( .A1(n14679), .A2(n15379), .ZN(n14680) );
  OAI211_X1 U16628 ( .C1(n14681), .C2(n15320), .A(n14680), .B(n14683), .ZN(
        n14780) );
  MUX2_X1 U16629 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n14780), .S(n15403), .Z(
        P1_U3559) );
  INV_X1 U16630 ( .A(n14682), .ZN(n14685) );
  OAI211_X1 U16631 ( .C1(n14685), .C2(n15366), .A(n14684), .B(n14683), .ZN(
        n14781) );
  MUX2_X1 U16632 ( .A(n14781), .B(P1_REG1_REG_30__SCAN_IN), .S(n7026), .Z(
        P1_U3558) );
  AOI21_X1 U16633 ( .B1(n15378), .B2(n14687), .A(n14686), .ZN(n14688) );
  OAI211_X1 U16634 ( .C1(n14690), .C2(n15366), .A(n14689), .B(n14688), .ZN(
        n14691) );
  INV_X1 U16635 ( .A(n14695), .ZN(n14703) );
  NAND3_X1 U16636 ( .A1(n14697), .A2(n15386), .A3(n14696), .ZN(n14699) );
  OAI211_X1 U16637 ( .C1(n14700), .C2(n15366), .A(n14699), .B(n14698), .ZN(
        n14701) );
  INV_X1 U16638 ( .A(n14701), .ZN(n14702) );
  NAND2_X1 U16639 ( .A1(n14703), .A2(n14702), .ZN(n14782) );
  MUX2_X1 U16640 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n14782), .S(n15403), .Z(
        P1_U3556) );
  AOI21_X1 U16641 ( .B1(n15379), .B2(n14705), .A(n14704), .ZN(n14706) );
  OAI211_X1 U16642 ( .C1(n15219), .C2(n14708), .A(n14707), .B(n14706), .ZN(
        n14783) );
  MUX2_X1 U16643 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n14783), .S(n15403), .Z(
        P1_U3555) );
  OAI21_X1 U16644 ( .B1(n15219), .B2(n14714), .A(n14713), .ZN(n14784) );
  MUX2_X1 U16645 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n14784), .S(n15403), .Z(
        P1_U3554) );
  OAI211_X1 U16646 ( .C1(n14717), .C2(n15366), .A(n14716), .B(n14715), .ZN(
        n14718) );
  AOI21_X1 U16647 ( .B1(n14719), .B2(n15386), .A(n14718), .ZN(n14720) );
  OAI21_X1 U16648 ( .B1(n14721), .B2(n15351), .A(n14720), .ZN(n14785) );
  MUX2_X1 U16649 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n14785), .S(n15403), .Z(
        P1_U3553) );
  INV_X1 U16650 ( .A(n14722), .ZN(n14727) );
  AOI21_X1 U16651 ( .B1(n15379), .B2(n14724), .A(n14723), .ZN(n14725) );
  OAI211_X1 U16652 ( .C1(n15219), .C2(n14727), .A(n14726), .B(n14725), .ZN(
        n14786) );
  MUX2_X1 U16653 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n14786), .S(n15403), .Z(
        P1_U3552) );
  NAND2_X1 U16654 ( .A1(n14728), .A2(n15375), .ZN(n14736) );
  AOI21_X1 U16655 ( .B1(n14730), .B2(n15379), .A(n14729), .ZN(n14735) );
  NAND3_X1 U16656 ( .A1(n14732), .A2(n14731), .A3(n15386), .ZN(n14734) );
  NAND4_X1 U16657 ( .A1(n14736), .A2(n14735), .A3(n14734), .A4(n14733), .ZN(
        n14787) );
  MUX2_X1 U16658 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n14787), .S(n15403), .Z(
        P1_U3551) );
  OAI21_X1 U16659 ( .B1(n15219), .B2(n14742), .A(n14741), .ZN(n14788) );
  MUX2_X1 U16660 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n14788), .S(n15403), .Z(
        P1_U3550) );
  AOI22_X1 U16661 ( .A1(n14744), .A2(n15288), .B1(n15379), .B2(n14743), .ZN(
        n14745) );
  OAI211_X1 U16662 ( .C1(n15219), .C2(n14747), .A(n14746), .B(n14745), .ZN(
        n14789) );
  MUX2_X1 U16663 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n14789), .S(n15403), .Z(
        P1_U3549) );
  OAI21_X1 U16664 ( .B1(n14749), .B2(n15366), .A(n14748), .ZN(n14750) );
  AOI21_X1 U16665 ( .B1(n14751), .B2(n15288), .A(n14750), .ZN(n14755) );
  NAND3_X1 U16666 ( .A1(n14753), .A2(n14752), .A3(n15386), .ZN(n14754) );
  OAI211_X1 U16667 ( .C1(n14756), .C2(n15351), .A(n14755), .B(n14754), .ZN(
        n14790) );
  MUX2_X1 U16668 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n14790), .S(n15403), .Z(
        P1_U3548) );
  AOI211_X1 U16669 ( .C1(n15379), .C2(n14759), .A(n14758), .B(n14757), .ZN(
        n14760) );
  OAI21_X1 U16670 ( .B1(n15219), .B2(n14761), .A(n14760), .ZN(n14791) );
  MUX2_X1 U16671 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n14791), .S(n15403), .Z(
        P1_U3547) );
  AOI22_X1 U16672 ( .A1(n14763), .A2(n15288), .B1(n15379), .B2(n14762), .ZN(
        n14764) );
  OAI211_X1 U16673 ( .C1(n15219), .C2(n14766), .A(n14765), .B(n14764), .ZN(
        n14792) );
  MUX2_X1 U16674 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n14792), .S(n15403), .Z(
        P1_U3546) );
  AOI211_X1 U16675 ( .C1(n15379), .C2(n14769), .A(n14768), .B(n14767), .ZN(
        n14770) );
  OAI21_X1 U16676 ( .B1(n15219), .B2(n14771), .A(n14770), .ZN(n14793) );
  MUX2_X1 U16677 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n14793), .S(n15403), .Z(
        P1_U3545) );
  AOI21_X1 U16678 ( .B1(n14773), .B2(n15379), .A(n14772), .ZN(n14774) );
  OAI21_X1 U16679 ( .B1(n14775), .B2(n15320), .A(n14774), .ZN(n14776) );
  AOI21_X1 U16680 ( .B1(n14777), .B2(n15375), .A(n14776), .ZN(n14778) );
  OAI21_X1 U16681 ( .B1(n15219), .B2(n14779), .A(n14778), .ZN(n14794) );
  MUX2_X1 U16682 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n14794), .S(n15403), .Z(
        P1_U3544) );
  MUX2_X1 U16683 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n14780), .S(n15389), .Z(
        P1_U3527) );
  MUX2_X1 U16684 ( .A(n14781), .B(P1_REG0_REG_30__SCAN_IN), .S(n15387), .Z(
        P1_U3526) );
  MUX2_X1 U16685 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n14782), .S(n15389), .Z(
        P1_U3524) );
  MUX2_X1 U16686 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n14783), .S(n15389), .Z(
        P1_U3523) );
  MUX2_X1 U16687 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n14784), .S(n15389), .Z(
        P1_U3522) );
  MUX2_X1 U16688 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n14785), .S(n15389), .Z(
        P1_U3521) );
  MUX2_X1 U16689 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n14786), .S(n15389), .Z(
        P1_U3520) );
  MUX2_X1 U16690 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n14787), .S(n15389), .Z(
        P1_U3519) );
  MUX2_X1 U16691 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n14788), .S(n15389), .Z(
        P1_U3518) );
  MUX2_X1 U16692 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n14789), .S(n15389), .Z(
        P1_U3517) );
  MUX2_X1 U16693 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n14790), .S(n15389), .Z(
        P1_U3516) );
  MUX2_X1 U16694 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n14791), .S(n15389), .Z(
        P1_U3515) );
  MUX2_X1 U16695 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n14792), .S(n15389), .Z(
        P1_U3513) );
  MUX2_X1 U16696 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n14793), .S(n15389), .Z(
        P1_U3510) );
  MUX2_X1 U16697 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n14794), .S(n15389), .Z(
        P1_U3507) );
  NOR4_X1 U16698 ( .A1(n14795), .A2(P1_IR_REG_30__SCAN_IN), .A3(n9336), .A4(
        P1_U3086), .ZN(n14796) );
  AOI21_X1 U16699 ( .B1(P2_DATAO_REG_31__SCAN_IN), .B2(n14797), .A(n14796), 
        .ZN(n14798) );
  OAI21_X1 U16700 ( .B1(n14799), .B2(n14815), .A(n14798), .ZN(P1_U3324) );
  OAI222_X1 U16701 ( .A1(n14817), .A2(n14803), .B1(n14815), .B2(n14802), .C1(
        n14801), .C2(P1_U3086), .ZN(P1_U3325) );
  OAI222_X1 U16702 ( .A1(n14817), .A2(n14806), .B1(n14815), .B2(n14805), .C1(
        n14804), .C2(P1_U3086), .ZN(P1_U3326) );
  OAI222_X1 U16703 ( .A1(n14817), .A2(n14809), .B1(n14815), .B2(n14808), .C1(
        n14807), .C2(P1_U3086), .ZN(P1_U3327) );
  OAI222_X1 U16704 ( .A1(n14812), .A2(P1_U3086), .B1(n14815), .B2(n14811), 
        .C1(n14810), .C2(n14817), .ZN(P1_U3329) );
  OAI222_X1 U16705 ( .A1(n14817), .A2(n14816), .B1(n14815), .B2(n14814), .C1(
        n14813), .C2(P1_U3086), .ZN(P1_U3330) );
  MUX2_X1 U16706 ( .A(n9763), .B(n14818), .S(P1_U3086), .Z(P1_U3333) );
  INV_X1 U16707 ( .A(n14819), .ZN(n14820) );
  MUX2_X1 U16708 ( .A(n14820), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  INV_X1 U16709 ( .A(P3_ADDR_REG_17__SCAN_IN), .ZN(n14854) );
  INV_X1 U16710 ( .A(P3_ADDR_REG_16__SCAN_IN), .ZN(n14852) );
  XNOR2_X1 U16711 ( .A(P1_ADDR_REG_16__SCAN_IN), .B(n14852), .ZN(n14918) );
  INV_X1 U16712 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n14850) );
  XOR2_X1 U16713 ( .A(P1_ADDR_REG_15__SCAN_IN), .B(n14850), .Z(n14856) );
  INV_X1 U16714 ( .A(P3_ADDR_REG_14__SCAN_IN), .ZN(n14848) );
  NOR2_X1 U16715 ( .A1(P1_ADDR_REG_13__SCAN_IN), .A2(n14846), .ZN(n14821) );
  AOI21_X1 U16716 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(n14846), .A(n14821), 
        .ZN(n14912) );
  INV_X1 U16717 ( .A(P3_ADDR_REG_11__SCAN_IN), .ZN(n14842) );
  NOR2_X1 U16718 ( .A1(n14822), .A2(n7269), .ZN(n14824) );
  NOR2_X1 U16719 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(n14883), .ZN(n14823) );
  NOR2_X1 U16720 ( .A1(n14827), .A2(n14826), .ZN(n14829) );
  NOR2_X1 U16721 ( .A1(P3_ADDR_REG_6__SCAN_IN), .A2(n14891), .ZN(n14830) );
  NOR2_X1 U16722 ( .A1(P3_ADDR_REG_7__SCAN_IN), .A2(n14831), .ZN(n14833) );
  XOR2_X1 U16723 ( .A(P3_ADDR_REG_7__SCAN_IN), .B(n14831), .Z(n14895) );
  NAND2_X1 U16724 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n14836), .ZN(n14834) );
  OAI21_X1 U16725 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(n14836), .A(n14834), .ZN(
        n14897) );
  XOR2_X1 U16726 ( .A(n15614), .B(P1_ADDR_REG_9__SCAN_IN), .Z(n14865) );
  NAND2_X1 U16727 ( .A1(n14866), .A2(n14865), .ZN(n14837) );
  NAND2_X1 U16728 ( .A1(n14862), .A2(n14864), .ZN(n14839) );
  NOR2_X1 U16729 ( .A1(n14862), .A2(n14864), .ZN(n14838) );
  XNOR2_X1 U16730 ( .A(P1_ADDR_REG_11__SCAN_IN), .B(n14842), .ZN(n14909) );
  XOR2_X1 U16731 ( .A(n14844), .B(P1_ADDR_REG_12__SCAN_IN), .Z(n14861) );
  NAND2_X1 U16732 ( .A1(n14860), .A2(n14861), .ZN(n14843) );
  NAND2_X1 U16733 ( .A1(n14912), .A2(n14913), .ZN(n14845) );
  XNOR2_X1 U16734 ( .A(n14848), .B(P1_ADDR_REG_14__SCAN_IN), .ZN(n14858) );
  NAND2_X1 U16735 ( .A1(n14856), .A2(n14857), .ZN(n14849) );
  NOR2_X1 U16736 ( .A1(n14918), .A2(n14917), .ZN(n14851) );
  AOI21_X1 U16737 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(n14852), .A(n14851), 
        .ZN(n14920) );
  XNOR2_X1 U16738 ( .A(n14854), .B(P1_ADDR_REG_17__SCAN_IN), .ZN(n14919) );
  NOR2_X1 U16739 ( .A1(n14920), .A2(n14919), .ZN(n14853) );
  AOI21_X1 U16740 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(n14854), .A(n14853), 
        .ZN(n14993) );
  NAND2_X1 U16741 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n14995), .ZN(n14855) );
  OAI21_X1 U16742 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n14995), .A(n14855), 
        .ZN(n14992) );
  XNOR2_X1 U16743 ( .A(n14993), .B(n14992), .ZN(n14997) );
  XOR2_X1 U16744 ( .A(n14857), .B(n14856), .Z(n15253) );
  XNOR2_X1 U16745 ( .A(n14859), .B(n14858), .ZN(n15249) );
  XNOR2_X1 U16746 ( .A(n14861), .B(n14860), .ZN(n14910) );
  XNOR2_X1 U16747 ( .A(n14862), .B(P3_ADDR_REG_10__SCAN_IN), .ZN(n14863) );
  XNOR2_X1 U16748 ( .A(n14864), .B(n14863), .ZN(n14906) );
  XOR2_X1 U16749 ( .A(n14866), .B(n14865), .Z(n14902) );
  INV_X1 U16750 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n14871) );
  NAND2_X1 U16751 ( .A1(n14870), .A2(n14871), .ZN(n14885) );
  XNOR2_X1 U16752 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(n14872), .ZN(n14873) );
  XNOR2_X1 U16753 ( .A(n14873), .B(P3_ADDR_REG_2__SCAN_IN), .ZN(n14881) );
  INV_X1 U16754 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n14875) );
  NOR2_X1 U16755 ( .A1(n14878), .A2(n14875), .ZN(n14879) );
  OAI21_X1 U16756 ( .B1(P3_ADDR_REG_0__SCAN_IN), .B2(n14877), .A(n14876), .ZN(
        n15795) );
  NAND2_X1 U16757 ( .A1(P2_ADDR_REG_0__SCAN_IN), .A2(n15795), .ZN(n15805) );
  XOR2_X1 U16758 ( .A(P2_ADDR_REG_1__SCAN_IN), .B(n14878), .Z(n15804) );
  NOR2_X1 U16759 ( .A1(n14881), .A2(n14880), .ZN(n14882) );
  INV_X1 U16760 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n14924) );
  XOR2_X1 U16761 ( .A(n14883), .B(P1_ADDR_REG_3__SCAN_IN), .Z(n15800) );
  NOR2_X1 U16762 ( .A1(n15801), .A2(n15800), .ZN(n14884) );
  NAND2_X1 U16763 ( .A1(n15801), .A2(n15800), .ZN(n15799) );
  OAI21_X1 U16764 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(n14884), .A(n15799), .ZN(
        n15790) );
  NAND2_X1 U16765 ( .A1(n15791), .A2(n15790), .ZN(n15789) );
  NAND2_X1 U16766 ( .A1(n14886), .A2(n14888), .ZN(n14889) );
  INV_X1 U16767 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n15793) );
  INV_X1 U16768 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n15448) );
  NOR2_X1 U16769 ( .A1(n14890), .A2(n15448), .ZN(n14894) );
  XOR2_X1 U16770 ( .A(n14891), .B(P3_ADDR_REG_6__SCAN_IN), .Z(n14893) );
  XNOR2_X1 U16771 ( .A(n14893), .B(n14892), .ZN(n14934) );
  XNOR2_X1 U16772 ( .A(n14895), .B(P1_ADDR_REG_7__SCAN_IN), .ZN(n15798) );
  XNOR2_X1 U16773 ( .A(n14898), .B(n14897), .ZN(n14900) );
  NAND2_X1 U16774 ( .A1(n14899), .A2(n14900), .ZN(n14901) );
  NOR2_X1 U16775 ( .A1(n14902), .A2(n14903), .ZN(n14904) );
  INV_X1 U16776 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n14951) );
  NAND2_X1 U16777 ( .A1(n14906), .A2(n14905), .ZN(n14907) );
  INV_X1 U16778 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n14953) );
  XNOR2_X1 U16779 ( .A(n14909), .B(n14908), .ZN(n15238) );
  INV_X1 U16780 ( .A(n15241), .ZN(n15242) );
  NAND2_X1 U16781 ( .A1(n15244), .A2(n15243), .ZN(n15240) );
  XOR2_X1 U16782 ( .A(n14913), .B(n14912), .Z(n14915) );
  INV_X1 U16783 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n15449) );
  NAND2_X1 U16784 ( .A1(n14915), .A2(n14914), .ZN(n14916) );
  NAND2_X1 U16785 ( .A1(n15249), .A2(n15248), .ZN(n15247) );
  XNOR2_X1 U16786 ( .A(n14918), .B(n14917), .ZN(n15256) );
  XNOR2_X1 U16787 ( .A(n14920), .B(n14919), .ZN(n14990) );
  NAND2_X1 U16788 ( .A1(n14989), .A2(n14990), .ZN(n14988) );
  AOI21_X1 U16789 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n14921) );
  OAI21_X1 U16790 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(n14921), 
        .ZN(U28) );
  AOI21_X1 U16791 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(
        P3_RD_REG_SCAN_IN), .ZN(n14922) );
  OAI21_X1 U16792 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(n14922), 
        .ZN(U29) );
  AOI21_X1 U16793 ( .B1(n14925), .B2(n14924), .A(n14923), .ZN(SUB_1596_U61) );
  AOI22_X1 U16794 ( .A1(n14926), .A2(n14945), .B1(SI_9_), .B2(n14944), .ZN(
        n14927) );
  OAI21_X1 U16795 ( .B1(P3_U3151), .B2(n14928), .A(n14927), .ZN(P3_U3286) );
  OAI22_X1 U16796 ( .A1(n14930), .A2(n14938), .B1(n14929), .B2(n14936), .ZN(
        n14931) );
  INV_X1 U16797 ( .A(n14931), .ZN(n14932) );
  OAI21_X1 U16798 ( .B1(P3_U3151), .B2(n15655), .A(n14932), .ZN(P3_U3282) );
  AOI21_X1 U16799 ( .B1(n14935), .B2(n14934), .A(n14933), .ZN(SUB_1596_U57) );
  OAI22_X1 U16800 ( .A1(n14939), .A2(n14938), .B1(n14937), .B2(n14936), .ZN(
        n14940) );
  INV_X1 U16801 ( .A(n14940), .ZN(n14941) );
  OAI21_X1 U16802 ( .B1(P3_U3151), .B2(n15676), .A(n14941), .ZN(P3_U3281) );
  OAI21_X1 U16803 ( .B1(n14943), .B2(n9484), .A(n14942), .ZN(SUB_1596_U55) );
  AOI22_X1 U16804 ( .A1(n14946), .A2(n14945), .B1(SI_18_), .B2(n14944), .ZN(
        n14947) );
  OAI21_X1 U16805 ( .B1(P3_U3151), .B2(n14948), .A(n14947), .ZN(P3_U3277) );
  AOI21_X1 U16806 ( .B1(n14951), .B2(n14950), .A(n14949), .ZN(SUB_1596_U54) );
  OAI21_X1 U16807 ( .B1(n14954), .B2(n14953), .A(n14952), .ZN(SUB_1596_U70) );
  NAND2_X1 U16808 ( .A1(n14955), .A2(n15379), .ZN(n14956) );
  AND2_X1 U16809 ( .A1(n14957), .A2(n14956), .ZN(n14961) );
  NAND2_X1 U16810 ( .A1(n14958), .A2(n15345), .ZN(n14960) );
  INV_X1 U16811 ( .A(n15341), .ZN(n15372) );
  NAND2_X1 U16812 ( .A1(n14958), .A2(n15372), .ZN(n14959) );
  AOI22_X1 U16813 ( .A1(n15389), .A2(n14965), .B1(n14963), .B2(n15387), .ZN(
        P1_U3495) );
  AOI22_X1 U16814 ( .A1(n15403), .A2(n14965), .B1(n14964), .B2(n7026), .ZN(
        P1_U3540) );
  NAND2_X1 U16815 ( .A1(n14967), .A2(n14966), .ZN(n15211) );
  NAND2_X1 U16816 ( .A1(n14969), .A2(n15211), .ZN(n14968) );
  OAI21_X1 U16817 ( .B1(n14969), .B2(P1_REG2_REG_13__SCAN_IN), .A(n14968), 
        .ZN(n14985) );
  XNOR2_X1 U16818 ( .A(n14970), .B(n14972), .ZN(n15220) );
  OAI211_X1 U16819 ( .C1(n14973), .C2(n14972), .A(n15375), .B(n14971), .ZN(
        n15217) );
  OR2_X1 U16820 ( .A1(n15217), .A2(n6665), .ZN(n14981) );
  AOI21_X1 U16821 ( .B1(n14974), .B2(n15216), .A(n15320), .ZN(n14976) );
  AND2_X1 U16822 ( .A1(n14976), .A2(n14975), .ZN(n15214) );
  NAND2_X1 U16823 ( .A1(n15216), .A2(n15282), .ZN(n14977) );
  OAI21_X1 U16824 ( .B1(n15213), .B2(n14978), .A(n14977), .ZN(n14979) );
  AOI21_X1 U16825 ( .B1(n15214), .B2(n15299), .A(n14979), .ZN(n14980) );
  OAI211_X1 U16826 ( .C1(n15220), .C2(n14982), .A(n14981), .B(n14980), .ZN(
        n14983) );
  INV_X1 U16827 ( .A(n14983), .ZN(n14984) );
  OAI211_X1 U16828 ( .C1(n14987), .C2(n14986), .A(n14985), .B(n14984), .ZN(
        P1_U3280) );
  OAI21_X1 U16829 ( .B1(n14990), .B2(n14989), .A(n14988), .ZN(n14991) );
  XNOR2_X1 U16830 ( .A(n14991), .B(P2_ADDR_REG_17__SCAN_IN), .ZN(SUB_1596_U63)
         );
  NOR2_X1 U16831 ( .A1(n14993), .A2(n14992), .ZN(n14994) );
  AOI21_X1 U16832 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n14995), .A(n14994), 
        .ZN(n15000) );
  AOI22_X1 U16833 ( .A1(n15002), .A2(n15001), .B1(P3_REG3_REG_16__SCAN_IN), 
        .B2(P3_U3151), .ZN(n15008) );
  XOR2_X1 U16834 ( .A(n15004), .B(n15003), .Z(n15006) );
  AOI22_X1 U16835 ( .A1(n15006), .A2(n15021), .B1(n15005), .B2(n15012), .ZN(
        n15007) );
  OAI211_X1 U16836 ( .C1(n15010), .C2(n15009), .A(n15008), .B(n15007), .ZN(
        P3_U3166) );
  AOI22_X1 U16837 ( .A1(n15012), .A2(n15110), .B1(P3_REG3_REG_13__SCAN_IN), 
        .B2(P3_U3151), .ZN(n15024) );
  XNOR2_X1 U16838 ( .A(n15014), .B(n15013), .ZN(n15015) );
  XNOR2_X1 U16839 ( .A(n15016), .B(n15015), .ZN(n15022) );
  OAI22_X1 U16840 ( .A1(n15020), .A2(n15019), .B1(n15018), .B2(n15017), .ZN(
        n15092) );
  AOI22_X1 U16841 ( .A1(n15022), .A2(n15021), .B1(n15591), .B2(n15092), .ZN(
        n15023) );
  OAI211_X1 U16842 ( .C1(n15094), .C2(n15593), .A(n15024), .B(n15023), .ZN(
        P3_U3174) );
  AOI21_X1 U16843 ( .B1(n15027), .B2(n15026), .A(n15025), .ZN(n15041) );
  OAI21_X1 U16844 ( .B1(P3_REG1_REG_15__SCAN_IN), .B2(n15029), .A(n15028), 
        .ZN(n15034) );
  AOI21_X1 U16845 ( .B1(n15674), .B2(P3_ADDR_REG_15__SCAN_IN), .A(n15030), 
        .ZN(n15031) );
  OAI21_X1 U16846 ( .B1(n15677), .B2(n15032), .A(n15031), .ZN(n15033) );
  AOI21_X1 U16847 ( .B1(n15034), .B2(n15679), .A(n15033), .ZN(n15040) );
  AOI21_X1 U16848 ( .B1(n15037), .B2(n15036), .A(n15035), .ZN(n15038) );
  OR2_X1 U16849 ( .A1(n15038), .A2(n15661), .ZN(n15039) );
  OAI211_X1 U16850 ( .C1(n15041), .C2(n15687), .A(n15040), .B(n15039), .ZN(
        P3_U3197) );
  AOI22_X1 U16851 ( .A1(n15604), .A2(n15042), .B1(n15674), .B2(
        P3_ADDR_REG_16__SCAN_IN), .ZN(n15058) );
  INV_X1 U16852 ( .A(n15043), .ZN(n15044) );
  NAND2_X1 U16853 ( .A1(n15045), .A2(n15044), .ZN(n15046) );
  XNOR2_X1 U16854 ( .A(n15047), .B(n15046), .ZN(n15052) );
  OAI21_X1 U16855 ( .B1(n15050), .B2(n15049), .A(n15048), .ZN(n15051) );
  AOI22_X1 U16856 ( .A1(n15052), .A2(n15681), .B1(n15679), .B2(n15051), .ZN(
        n15057) );
  NAND2_X1 U16857 ( .A1(P3_REG3_REG_16__SCAN_IN), .A2(P3_U3151), .ZN(n15056)
         );
  OAI221_X1 U16858 ( .B1(n15054), .B2(n6770), .C1(n15054), .C2(n15053), .A(
        n15082), .ZN(n15055) );
  NAND4_X1 U16859 ( .A1(n15058), .A2(n15057), .A3(n15056), .A4(n15055), .ZN(
        P3_U3198) );
  AOI22_X1 U16860 ( .A1(n15604), .A2(n7689), .B1(n15674), .B2(
        P3_ADDR_REG_17__SCAN_IN), .ZN(n15072) );
  OAI21_X1 U16861 ( .B1(P3_REG1_REG_17__SCAN_IN), .B2(n15060), .A(n15059), 
        .ZN(n15065) );
  AOI211_X1 U16862 ( .C1(n15063), .C2(n15062), .A(n15061), .B(n15661), .ZN(
        n15064) );
  AOI21_X1 U16863 ( .B1(n15679), .B2(n15065), .A(n15064), .ZN(n15071) );
  NAND2_X1 U16864 ( .A1(P3_REG3_REG_17__SCAN_IN), .A2(P3_U3151), .ZN(n15070)
         );
  OAI221_X1 U16865 ( .B1(n15068), .B2(n15067), .C1(n15068), .C2(n15066), .A(
        n15082), .ZN(n15069) );
  NAND4_X1 U16866 ( .A1(n15072), .A2(n15071), .A3(n15070), .A4(n15069), .ZN(
        P3_U3199) );
  AOI22_X1 U16867 ( .A1(n15604), .A2(n15073), .B1(n15674), .B2(
        P3_ADDR_REG_18__SCAN_IN), .ZN(n15088) );
  OAI21_X1 U16868 ( .B1(n15076), .B2(n15075), .A(n15074), .ZN(n15081) );
  OAI21_X1 U16869 ( .B1(n15079), .B2(n15078), .A(n15077), .ZN(n15080) );
  AOI22_X1 U16870 ( .A1(n15081), .A2(n15679), .B1(n15681), .B2(n15080), .ZN(
        n15087) );
  OAI221_X1 U16871 ( .B1(n15084), .B2(n6741), .C1(n15084), .C2(n15083), .A(
        n15082), .ZN(n15085) );
  NAND4_X1 U16872 ( .A1(n15088), .A2(n15087), .A3(n15086), .A4(n15085), .ZN(
        P3_U3200) );
  AOI22_X1 U16873 ( .A1(n15102), .A2(n15097), .B1(P3_REG2_REG_30__SCAN_IN), 
        .B2(n15703), .ZN(n15089) );
  NAND2_X1 U16874 ( .A1(n15090), .A2(n15089), .ZN(P3_U3203) );
  XNOR2_X1 U16875 ( .A(n15091), .B(n6693), .ZN(n15093) );
  AOI21_X1 U16876 ( .B1(n15093), .B2(n15695), .A(n15092), .ZN(n15113) );
  OAI22_X1 U16877 ( .A1(n15719), .A2(n8190), .B1(n15711), .B2(n15094), .ZN(
        n15095) );
  INV_X1 U16878 ( .A(n15095), .ZN(n15100) );
  XNOR2_X1 U16879 ( .A(n15096), .B(n6693), .ZN(n15111) );
  AOI22_X1 U16880 ( .A1(n15111), .A2(n15098), .B1(n15110), .B2(n15097), .ZN(
        n15099) );
  OAI211_X1 U16881 ( .C1(n15703), .C2(n15113), .A(n15100), .B(n15099), .ZN(
        P3_U3220) );
  AOI21_X1 U16882 ( .B1(n15102), .B2(n15770), .A(n15101), .ZN(n15115) );
  INV_X1 U16883 ( .A(P3_REG1_REG_30__SCAN_IN), .ZN(n15103) );
  AOI22_X1 U16884 ( .A1(n15788), .A2(n15115), .B1(n15103), .B2(n15786), .ZN(
        P3_U3489) );
  INV_X1 U16885 ( .A(n15104), .ZN(n15107) );
  OAI22_X1 U16886 ( .A1(n15107), .A2(n15106), .B1(n15744), .B2(n15105), .ZN(
        n15108) );
  NOR2_X1 U16887 ( .A1(n15109), .A2(n15108), .ZN(n15117) );
  AOI22_X1 U16888 ( .A1(n15788), .A2(n15117), .B1(n12640), .B2(n15786), .ZN(
        P3_U3473) );
  AOI22_X1 U16889 ( .A1(n15111), .A2(n15746), .B1(n15770), .B2(n15110), .ZN(
        n15112) );
  AND2_X1 U16890 ( .A1(n15113), .A2(n15112), .ZN(n15119) );
  AOI22_X1 U16891 ( .A1(n15788), .A2(n15119), .B1(n8191), .B2(n15786), .ZN(
        P3_U3472) );
  AOI22_X1 U16892 ( .A1(n15773), .A2(n15115), .B1(n15114), .B2(n15771), .ZN(
        P3_U3457) );
  INV_X1 U16893 ( .A(P3_REG0_REG_14__SCAN_IN), .ZN(n15116) );
  AOI22_X1 U16894 ( .A1(n15773), .A2(n15117), .B1(n15116), .B2(n15771), .ZN(
        P3_U3432) );
  INV_X1 U16895 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n15118) );
  AOI22_X1 U16896 ( .A1(n15773), .A2(n15119), .B1(n15118), .B2(n15771), .ZN(
        P3_U3429) );
  OAI21_X1 U16897 ( .B1(n15122), .B2(n15121), .A(n15120), .ZN(n15124) );
  AOI222_X1 U16898 ( .A1(n15128), .A2(n15127), .B1(n15126), .B2(n15125), .C1(
        n15124), .C2(n15123), .ZN(n15130) );
  OAI211_X1 U16899 ( .C1(n15132), .C2(n15131), .A(n15130), .B(n15129), .ZN(
        P2_U3187) );
  XNOR2_X1 U16900 ( .A(n15133), .B(n15141), .ZN(n15136) );
  INV_X1 U16901 ( .A(n15134), .ZN(n15135) );
  AOI21_X1 U16902 ( .B1(n15136), .B2(n15551), .A(n15135), .ZN(n15153) );
  AOI222_X1 U16903 ( .A1(n15140), .A2(n15139), .B1(n15138), .B2(n15137), .C1(
        P2_REG2_REG_12__SCAN_IN), .C2(n15151), .ZN(n15150) );
  XNOR2_X1 U16904 ( .A(n15142), .B(n15141), .ZN(n15156) );
  OAI211_X1 U16905 ( .C1(n15145), .C2(n15154), .A(n15144), .B(n15143), .ZN(
        n15152) );
  INV_X1 U16906 ( .A(n15152), .ZN(n15146) );
  AOI22_X1 U16907 ( .A1(n15156), .A2(n15148), .B1(n15147), .B2(n15146), .ZN(
        n15149) );
  OAI211_X1 U16908 ( .C1(n15151), .C2(n15153), .A(n15150), .B(n15149), .ZN(
        P2_U3253) );
  OAI211_X1 U16909 ( .C1(n15154), .C2(n15548), .A(n15153), .B(n15152), .ZN(
        n15155) );
  AOI21_X1 U16910 ( .B1(n15156), .B2(n15527), .A(n15155), .ZN(n15160) );
  AOI22_X1 U16911 ( .A1(n15158), .A2(n15160), .B1(n15157), .B2(n15573), .ZN(
        P2_U3511) );
  INV_X1 U16912 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n15159) );
  AOI22_X1 U16913 ( .A1(n15561), .A2(n15160), .B1(n15159), .B2(n15559), .ZN(
        P2_U3466) );
  OAI22_X1 U16914 ( .A1(n15164), .A2(n15163), .B1(n15162), .B2(n15161), .ZN(
        n15171) );
  NAND2_X1 U16915 ( .A1(n15165), .A2(n15166), .ZN(n15168) );
  AOI21_X1 U16916 ( .B1(n15169), .B2(n15168), .A(n15167), .ZN(n15170) );
  AOI211_X1 U16917 ( .C1(n15172), .C2(n15203), .A(n15171), .B(n15170), .ZN(
        n15174) );
  OAI211_X1 U16918 ( .C1(n15176), .C2(n15175), .A(n15174), .B(n15173), .ZN(
        P1_U3215) );
  OAI211_X1 U16919 ( .C1(n15179), .C2(n15178), .A(n15177), .B(n15375), .ZN(
        n15181) );
  AND2_X1 U16920 ( .A1(n15181), .A2(n15180), .ZN(n15223) );
  AOI222_X1 U16921 ( .A1(n15183), .A2(n15282), .B1(P1_REG2_REG_11__SCAN_IN), 
        .B2(n6665), .C1(n15293), .C2(n15182), .ZN(n15193) );
  XNOR2_X1 U16922 ( .A(n15185), .B(n15184), .ZN(n15226) );
  INV_X1 U16923 ( .A(n15186), .ZN(n15189) );
  INV_X1 U16924 ( .A(n15187), .ZN(n15188) );
  OAI211_X1 U16925 ( .C1(n15224), .C2(n15189), .A(n15188), .B(n15288), .ZN(
        n15222) );
  INV_X1 U16926 ( .A(n15222), .ZN(n15190) );
  AOI22_X1 U16927 ( .A1(n15226), .A2(n15191), .B1(n15299), .B2(n15190), .ZN(
        n15192) );
  OAI211_X1 U16928 ( .C1(n6665), .C2(n15223), .A(n15193), .B(n15192), .ZN(
        P1_U3282) );
  AND2_X1 U16929 ( .A1(n15386), .A2(n15194), .ZN(n15198) );
  OAI22_X1 U16930 ( .A1(n15196), .A2(n15320), .B1(n15195), .B2(n15366), .ZN(
        n15197) );
  NOR3_X1 U16931 ( .A1(n15199), .A2(n15198), .A3(n15197), .ZN(n15229) );
  INV_X1 U16932 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n15200) );
  AOI22_X1 U16933 ( .A1(n15403), .A2(n15229), .B1(n15200), .B2(n7026), .ZN(
        P1_U3543) );
  AOI211_X1 U16934 ( .C1(n15379), .C2(n15203), .A(n15202), .B(n15201), .ZN(
        n15207) );
  NAND3_X1 U16935 ( .A1(n15205), .A2(n15204), .A3(n15386), .ZN(n15206) );
  OAI211_X1 U16936 ( .C1(n15208), .C2(n15351), .A(n15207), .B(n15206), .ZN(
        n15209) );
  INV_X1 U16937 ( .A(n15209), .ZN(n15231) );
  AOI22_X1 U16938 ( .A1(n15403), .A2(n15231), .B1(n15210), .B2(n7026), .ZN(
        P1_U3542) );
  OAI21_X1 U16939 ( .B1(n15213), .B2(n15212), .A(n15211), .ZN(n15215) );
  AOI211_X1 U16940 ( .C1(n15379), .C2(n15216), .A(n15215), .B(n15214), .ZN(
        n15218) );
  OAI211_X1 U16941 ( .C1(n15220), .C2(n15219), .A(n15218), .B(n15217), .ZN(
        n15221) );
  INV_X1 U16942 ( .A(n15221), .ZN(n15233) );
  AOI22_X1 U16943 ( .A1(n15403), .A2(n15233), .B1(n10496), .B2(n7026), .ZN(
        P1_U3541) );
  OAI211_X1 U16944 ( .C1(n15224), .C2(n15366), .A(n15223), .B(n15222), .ZN(
        n15225) );
  AOI21_X1 U16945 ( .B1(n15226), .B2(n15386), .A(n15225), .ZN(n15235) );
  AOI22_X1 U16946 ( .A1(n15403), .A2(n15235), .B1(n15227), .B2(n7026), .ZN(
        P1_U3539) );
  INV_X1 U16947 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n15228) );
  AOI22_X1 U16948 ( .A1(n15389), .A2(n15229), .B1(n15228), .B2(n15387), .ZN(
        P1_U3504) );
  INV_X1 U16949 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n15230) );
  AOI22_X1 U16950 ( .A1(n15389), .A2(n15231), .B1(n15230), .B2(n15387), .ZN(
        P1_U3501) );
  AOI22_X1 U16951 ( .A1(n15389), .A2(n15233), .B1(n15232), .B2(n15387), .ZN(
        P1_U3498) );
  INV_X1 U16952 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n15234) );
  AOI22_X1 U16953 ( .A1(n15389), .A2(n15235), .B1(n15234), .B2(n15387), .ZN(
        P1_U3492) );
  OAI21_X1 U16954 ( .B1(n15238), .B2(n15237), .A(n15236), .ZN(n15239) );
  XNOR2_X1 U16955 ( .A(n15239), .B(P2_ADDR_REG_11__SCAN_IN), .ZN(SUB_1596_U69)
         );
  OAI222_X1 U16956 ( .A1(n15244), .A2(n15243), .B1(n15244), .B2(n15242), .C1(
        n15241), .C2(n15240), .ZN(SUB_1596_U68) );
  OAI21_X1 U16957 ( .B1(n15246), .B2(n15449), .A(n15245), .ZN(SUB_1596_U67) );
  OAI21_X1 U16958 ( .B1(n15249), .B2(n15248), .A(n15247), .ZN(n15250) );
  XNOR2_X1 U16959 ( .A(n15250), .B(P2_ADDR_REG_14__SCAN_IN), .ZN(SUB_1596_U66)
         );
  AOI21_X1 U16960 ( .B1(n15253), .B2(n15252), .A(n15251), .ZN(n15254) );
  XOR2_X1 U16961 ( .A(P2_ADDR_REG_15__SCAN_IN), .B(n15254), .Z(SUB_1596_U65)
         );
  AOI21_X1 U16962 ( .B1(n15257), .B2(n15256), .A(n15255), .ZN(n15258) );
  XOR2_X1 U16963 ( .A(P2_ADDR_REG_16__SCAN_IN), .B(n15258), .Z(SUB_1596_U64)
         );
  INV_X1 U16964 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n15272) );
  OAI21_X1 U16965 ( .B1(P1_REG2_REG_18__SCAN_IN), .B2(n15260), .A(n15259), 
        .ZN(n15265) );
  OAI21_X1 U16966 ( .B1(P1_REG1_REG_18__SCAN_IN), .B2(n15262), .A(n15261), 
        .ZN(n15263) );
  OAI222_X1 U16967 ( .A1(n15267), .A2(n7164), .B1(n15266), .B2(n15265), .C1(
        n15264), .C2(n15263), .ZN(n15268) );
  INV_X1 U16968 ( .A(n15268), .ZN(n15270) );
  OAI211_X1 U16969 ( .C1(n15272), .C2(n15271), .A(n15270), .B(n15269), .ZN(
        P1_U3261) );
  OAI21_X1 U16970 ( .B1(n15274), .B2(n15276), .A(n15273), .ZN(n15280) );
  INV_X1 U16971 ( .A(n15275), .ZN(n15279) );
  XNOR2_X1 U16972 ( .A(n15277), .B(n15276), .ZN(n15283) );
  NOR2_X1 U16973 ( .A1(n15283), .A2(n15318), .ZN(n15278) );
  AOI211_X1 U16974 ( .C1(n15375), .C2(n15280), .A(n15279), .B(n15278), .ZN(
        n15368) );
  AOI222_X1 U16975 ( .A1(n15286), .A2(n15282), .B1(P1_REG2_REG_9__SCAN_IN), 
        .B2(n6665), .C1(n15293), .C2(n15281), .ZN(n15292) );
  INV_X1 U16976 ( .A(n15283), .ZN(n15371) );
  INV_X1 U16977 ( .A(n15284), .ZN(n15301) );
  INV_X1 U16978 ( .A(n15285), .ZN(n15289) );
  INV_X1 U16979 ( .A(n15286), .ZN(n15367) );
  OAI211_X1 U16980 ( .C1(n15289), .C2(n15367), .A(n15288), .B(n15287), .ZN(
        n15365) );
  INV_X1 U16981 ( .A(n15365), .ZN(n15290) );
  AOI22_X1 U16982 ( .A1(n15371), .A2(n15301), .B1(n15299), .B2(n15290), .ZN(
        n15291) );
  OAI211_X1 U16983 ( .C1(n6665), .C2(n15368), .A(n15292), .B(n15291), .ZN(
        P1_U3284) );
  AOI22_X1 U16984 ( .A1(n6665), .A2(P1_REG2_REG_5__SCAN_IN), .B1(n15294), .B2(
        n15293), .ZN(n15295) );
  OAI21_X1 U16985 ( .B1(n15297), .B2(n15296), .A(n15295), .ZN(n15298) );
  INV_X1 U16986 ( .A(n15298), .ZN(n15304) );
  AOI22_X1 U16987 ( .A1(n15302), .A2(n15301), .B1(n15300), .B2(n15299), .ZN(
        n15303) );
  OAI211_X1 U16988 ( .C1(n6665), .C2(n15305), .A(n15304), .B(n15303), .ZN(
        P1_U3288) );
  AND2_X1 U16989 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n15314), .ZN(P1_U3294) );
  NOR2_X1 U16990 ( .A1(n15313), .A2(n15306), .ZN(P1_U3295) );
  NOR2_X1 U16991 ( .A1(n15313), .A2(n15307), .ZN(P1_U3296) );
  AND2_X1 U16992 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n15314), .ZN(P1_U3297) );
  AND2_X1 U16993 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n15314), .ZN(P1_U3298) );
  AND2_X1 U16994 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n15314), .ZN(P1_U3299) );
  AND2_X1 U16995 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n15314), .ZN(P1_U3300) );
  AND2_X1 U16996 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n15314), .ZN(P1_U3301) );
  AND2_X1 U16997 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n15314), .ZN(P1_U3302) );
  AND2_X1 U16998 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n15314), .ZN(P1_U3303) );
  AND2_X1 U16999 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n15314), .ZN(P1_U3304) );
  NOR2_X1 U17000 ( .A1(n15313), .A2(n15308), .ZN(P1_U3305) );
  AND2_X1 U17001 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n15314), .ZN(P1_U3306) );
  AND2_X1 U17002 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n15314), .ZN(P1_U3307) );
  NOR2_X1 U17003 ( .A1(n15313), .A2(n15309), .ZN(P1_U3308) );
  AND2_X1 U17004 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n15314), .ZN(P1_U3309) );
  AND2_X1 U17005 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n15314), .ZN(P1_U3310) );
  AND2_X1 U17006 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n15314), .ZN(P1_U3311) );
  AND2_X1 U17007 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n15314), .ZN(P1_U3312) );
  AND2_X1 U17008 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n15314), .ZN(P1_U3313) );
  NOR2_X1 U17009 ( .A1(n15313), .A2(n15310), .ZN(P1_U3314) );
  NOR2_X1 U17010 ( .A1(n15313), .A2(n15311), .ZN(P1_U3315) );
  AND2_X1 U17011 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n15314), .ZN(P1_U3316) );
  NOR2_X1 U17012 ( .A1(n15313), .A2(n15312), .ZN(P1_U3317) );
  AND2_X1 U17013 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n15314), .ZN(P1_U3318) );
  AND2_X1 U17014 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n15314), .ZN(P1_U3319) );
  AND2_X1 U17015 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n15314), .ZN(P1_U3320) );
  AND2_X1 U17016 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n15314), .ZN(P1_U3321) );
  AND2_X1 U17017 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n15314), .ZN(P1_U3322) );
  AND2_X1 U17018 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n15314), .ZN(P1_U3323) );
  NOR3_X1 U17019 ( .A1(n15316), .A2(n15351), .A3(n15315), .ZN(n15325) );
  AOI21_X1 U17020 ( .B1(n15318), .B2(n15341), .A(n15317), .ZN(n15323) );
  OAI22_X1 U17021 ( .A1(n15321), .A2(n15320), .B1(n15319), .B2(n15366), .ZN(
        n15322) );
  NOR4_X1 U17022 ( .A1(n15325), .A2(n15324), .A3(n15323), .A4(n15322), .ZN(
        n15391) );
  INV_X1 U17023 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n15326) );
  AOI22_X1 U17024 ( .A1(n15389), .A2(n15391), .B1(n15326), .B2(n15387), .ZN(
        P1_U3462) );
  INV_X1 U17025 ( .A(n15327), .ZN(n15333) );
  NOR2_X1 U17026 ( .A1(n15327), .A2(n15341), .ZN(n15332) );
  OAI211_X1 U17027 ( .C1(n15330), .C2(n15366), .A(n15329), .B(n15328), .ZN(
        n15331) );
  AOI211_X1 U17028 ( .C1(n15333), .C2(n15345), .A(n15332), .B(n15331), .ZN(
        n15393) );
  INV_X1 U17029 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n15334) );
  AOI22_X1 U17030 ( .A1(n15389), .A2(n15393), .B1(n15334), .B2(n15387), .ZN(
        P1_U3465) );
  INV_X1 U17031 ( .A(n15342), .ZN(n15344) );
  AOI211_X1 U17032 ( .C1(n15379), .C2(n15337), .A(n15336), .B(n15335), .ZN(
        n15340) );
  NAND2_X1 U17033 ( .A1(n15338), .A2(n15375), .ZN(n15339) );
  OAI211_X1 U17034 ( .C1(n15342), .C2(n15341), .A(n15340), .B(n15339), .ZN(
        n15343) );
  AOI21_X1 U17035 ( .B1(n15345), .B2(n15344), .A(n15343), .ZN(n15395) );
  INV_X1 U17036 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n15346) );
  AOI22_X1 U17037 ( .A1(n15389), .A2(n15395), .B1(n15346), .B2(n15387), .ZN(
        P1_U3477) );
  NOR3_X1 U17038 ( .A1(n15349), .A2(n15348), .A3(n15347), .ZN(n15350) );
  OAI21_X1 U17039 ( .B1(n15352), .B2(n15351), .A(n15350), .ZN(n15353) );
  AOI21_X1 U17040 ( .B1(n15354), .B2(n15386), .A(n15353), .ZN(n15397) );
  AOI22_X1 U17041 ( .A1(n15389), .A2(n15397), .B1(n15355), .B2(n15387), .ZN(
        P1_U3480) );
  OAI211_X1 U17042 ( .C1(n15358), .C2(n15366), .A(n15357), .B(n15356), .ZN(
        n15362) );
  AND3_X1 U17043 ( .A1(n15360), .A2(n15375), .A3(n15359), .ZN(n15361) );
  AOI211_X1 U17044 ( .C1(n15363), .C2(n15386), .A(n15362), .B(n15361), .ZN(
        n15398) );
  INV_X1 U17045 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n15364) );
  AOI22_X1 U17046 ( .A1(n15389), .A2(n15398), .B1(n15364), .B2(n15387), .ZN(
        P1_U3483) );
  OAI21_X1 U17047 ( .B1(n15367), .B2(n15366), .A(n15365), .ZN(n15370) );
  INV_X1 U17048 ( .A(n15368), .ZN(n15369) );
  AOI211_X1 U17049 ( .C1(n15372), .C2(n15371), .A(n15370), .B(n15369), .ZN(
        n15400) );
  INV_X1 U17050 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n15373) );
  AOI22_X1 U17051 ( .A1(n15389), .A2(n15400), .B1(n15373), .B2(n15387), .ZN(
        P1_U3486) );
  NAND3_X1 U17052 ( .A1(n15376), .A2(n15375), .A3(n15374), .ZN(n15383) );
  AOI22_X1 U17053 ( .A1(n15380), .A2(n15379), .B1(n15378), .B2(n15377), .ZN(
        n15381) );
  NAND3_X1 U17054 ( .A1(n15383), .A2(n15382), .A3(n15381), .ZN(n15384) );
  AOI21_X1 U17055 ( .B1(n15386), .B2(n15385), .A(n15384), .ZN(n15402) );
  INV_X1 U17056 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n15388) );
  AOI22_X1 U17057 ( .A1(n15389), .A2(n15402), .B1(n15388), .B2(n15387), .ZN(
        P1_U3489) );
  AOI22_X1 U17058 ( .A1(n15403), .A2(n15391), .B1(n15390), .B2(n7026), .ZN(
        P1_U3529) );
  AOI22_X1 U17059 ( .A1(n15403), .A2(n15393), .B1(n15392), .B2(n7026), .ZN(
        P1_U3530) );
  AOI22_X1 U17060 ( .A1(n15403), .A2(n15395), .B1(n15394), .B2(n7026), .ZN(
        P1_U3534) );
  AOI22_X1 U17061 ( .A1(n15403), .A2(n15397), .B1(n15396), .B2(n7026), .ZN(
        P1_U3535) );
  AOI22_X1 U17062 ( .A1(n15403), .A2(n15398), .B1(n9708), .B2(n7026), .ZN(
        P1_U3536) );
  AOI22_X1 U17063 ( .A1(n15403), .A2(n15400), .B1(n15399), .B2(n7026), .ZN(
        P1_U3537) );
  AOI22_X1 U17064 ( .A1(n15403), .A2(n15402), .B1(n15401), .B2(n7026), .ZN(
        P1_U3538) );
  NOR2_X1 U17065 ( .A1(n15472), .A2(P2_U3947), .ZN(P2_U3087) );
  AOI22_X1 U17066 ( .A1(P2_REG2_REG_0__SCAN_IN), .A2(n15474), .B1(n15467), 
        .B2(P2_REG1_REG_0__SCAN_IN), .ZN(n15407) );
  AOI22_X1 U17067 ( .A1(n15472), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3088), .ZN(n15406) );
  OAI22_X1 U17068 ( .A1(n15459), .A2(P2_REG1_REG_0__SCAN_IN), .B1(
        P2_REG2_REG_0__SCAN_IN), .B2(n15442), .ZN(n15404) );
  OAI21_X1 U17069 ( .B1(n15453), .B2(n15404), .A(P2_IR_REG_0__SCAN_IN), .ZN(
        n15405) );
  OAI211_X1 U17070 ( .C1(P2_IR_REG_0__SCAN_IN), .C2(n15407), .A(n15406), .B(
        n15405), .ZN(P2_U3214) );
  OAI21_X1 U17071 ( .B1(n15420), .B2(n8537), .A(P2_STATE_REG_SCAN_IN), .ZN(
        n15408) );
  OAI21_X1 U17072 ( .B1(P2_STATE_REG_SCAN_IN), .B2(P2_REG3_REG_1__SCAN_IN), 
        .A(n15408), .ZN(n15418) );
  AND2_X1 U17073 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n15411) );
  OAI211_X1 U17074 ( .C1(n15411), .C2(n15410), .A(n15474), .B(n15409), .ZN(
        n15417) );
  NAND2_X1 U17075 ( .A1(P2_ADDR_REG_1__SCAN_IN), .A2(n15472), .ZN(n15416) );
  OAI211_X1 U17076 ( .C1(n15414), .C2(n15413), .A(n15467), .B(n15412), .ZN(
        n15415) );
  NAND4_X1 U17077 ( .A1(n15418), .A2(n15417), .A3(n15416), .A4(n15415), .ZN(
        P2_U3215) );
  OAI21_X1 U17078 ( .B1(n15420), .B2(n15419), .A(P2_STATE_REG_SCAN_IN), .ZN(
        n15421) );
  OAI21_X1 U17079 ( .B1(P2_STATE_REG_SCAN_IN), .B2(P2_REG3_REG_4__SCAN_IN), 
        .A(n15421), .ZN(n15431) );
  OAI211_X1 U17080 ( .C1(n15424), .C2(n15423), .A(n15474), .B(n15422), .ZN(
        n15430) );
  OAI211_X1 U17081 ( .C1(n15427), .C2(n15426), .A(n15467), .B(n15425), .ZN(
        n15429) );
  NAND2_X1 U17082 ( .A1(P2_ADDR_REG_4__SCAN_IN), .A2(n15472), .ZN(n15428) );
  NAND4_X1 U17083 ( .A1(n15431), .A2(n15430), .A3(n15429), .A4(n15428), .ZN(
        P2_U3218) );
  NAND3_X1 U17084 ( .A1(n15434), .A2(n15433), .A3(n15432), .ZN(n15435) );
  NAND3_X1 U17085 ( .A1(n15467), .A2(n15436), .A3(n15435), .ZN(n15438) );
  OAI211_X1 U17086 ( .C1(n15479), .C2(n15439), .A(n15438), .B(n15437), .ZN(
        n15440) );
  INV_X1 U17087 ( .A(n15440), .ZN(n15447) );
  AOI211_X1 U17088 ( .C1(n15444), .C2(n15443), .A(n15442), .B(n15441), .ZN(
        n15445) );
  INV_X1 U17089 ( .A(n15445), .ZN(n15446) );
  OAI211_X1 U17090 ( .C1(n15450), .C2(n15448), .A(n15447), .B(n15446), .ZN(
        P2_U3220) );
  OAI22_X1 U17091 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n15451), .B1(n15450), .B2(
        n15449), .ZN(n15452) );
  AOI21_X1 U17092 ( .B1(n15454), .B2(n15453), .A(n15452), .ZN(n15465) );
  OAI211_X1 U17093 ( .C1(n15457), .C2(n15456), .A(n15455), .B(n15474), .ZN(
        n15464) );
  AOI211_X1 U17094 ( .C1(n15461), .C2(n15460), .A(n15459), .B(n15458), .ZN(
        n15462) );
  INV_X1 U17095 ( .A(n15462), .ZN(n15463) );
  NAND3_X1 U17096 ( .A1(n15465), .A2(n15464), .A3(n15463), .ZN(P2_U3227) );
  OAI211_X1 U17097 ( .C1(n15468), .C2(P2_REG1_REG_15__SCAN_IN), .A(n15467), 
        .B(n15466), .ZN(n15469) );
  NAND2_X1 U17098 ( .A1(n15470), .A2(n15469), .ZN(n15471) );
  AOI21_X1 U17099 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(n15472), .A(n15471), 
        .ZN(n15477) );
  OAI211_X1 U17100 ( .C1(P2_REG2_REG_15__SCAN_IN), .C2(n15475), .A(n15474), 
        .B(n15473), .ZN(n15476) );
  OAI211_X1 U17101 ( .C1(n15479), .C2(n15478), .A(n15477), .B(n15476), .ZN(
        P2_U3229) );
  AND2_X1 U17102 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n15485), .ZN(P2_U3266) );
  AND2_X1 U17103 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n15485), .ZN(P2_U3267) );
  AND2_X1 U17104 ( .A1(n15485), .A2(P2_D_REG_29__SCAN_IN), .ZN(P2_U3268) );
  AND2_X1 U17105 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n15485), .ZN(P2_U3269) );
  AND2_X1 U17106 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n15485), .ZN(P2_U3270) );
  AND2_X1 U17107 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n15485), .ZN(P2_U3271) );
  AND2_X1 U17108 ( .A1(n15485), .A2(P2_D_REG_25__SCAN_IN), .ZN(P2_U3272) );
  AND2_X1 U17109 ( .A1(n15485), .A2(P2_D_REG_24__SCAN_IN), .ZN(P2_U3273) );
  AND2_X1 U17110 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n15485), .ZN(P2_U3274) );
  AND2_X1 U17111 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n15485), .ZN(P2_U3275) );
  AND2_X1 U17112 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n15485), .ZN(P2_U3276) );
  AND2_X1 U17113 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n15485), .ZN(P2_U3277) );
  AND2_X1 U17114 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n15485), .ZN(P2_U3278) );
  AND2_X1 U17115 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n15485), .ZN(P2_U3279) );
  NOR2_X1 U17116 ( .A1(n15484), .A2(n15481), .ZN(P2_U3280) );
  AND2_X1 U17117 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n15485), .ZN(P2_U3281) );
  AND2_X1 U17118 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n15485), .ZN(P2_U3282) );
  AND2_X1 U17119 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n15485), .ZN(P2_U3283) );
  AND2_X1 U17120 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n15485), .ZN(P2_U3284) );
  AND2_X1 U17121 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n15485), .ZN(P2_U3285) );
  AND2_X1 U17122 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n15485), .ZN(P2_U3286) );
  AND2_X1 U17123 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n15485), .ZN(P2_U3287) );
  AND2_X1 U17124 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n15485), .ZN(P2_U3288) );
  NOR2_X1 U17125 ( .A1(n15484), .A2(n15482), .ZN(P2_U3289) );
  NOR2_X1 U17126 ( .A1(n15484), .A2(n15483), .ZN(P2_U3290) );
  AND2_X1 U17127 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n15485), .ZN(P2_U3291) );
  AND2_X1 U17128 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n15485), .ZN(P2_U3292) );
  AND2_X1 U17129 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n15485), .ZN(P2_U3293) );
  AND2_X1 U17130 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n15485), .ZN(P2_U3294) );
  AND2_X1 U17131 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n15485), .ZN(P2_U3295) );
  AOI21_X1 U17132 ( .B1(n15488), .B2(n15487), .A(n15486), .ZN(P2_U3416) );
  AOI22_X1 U17133 ( .A1(n15491), .A2(n15490), .B1(n15489), .B2(n15488), .ZN(
        P2_U3417) );
  OAI211_X1 U17134 ( .C1(n15554), .C2(n15494), .A(n15493), .B(n15492), .ZN(
        n15495) );
  INV_X1 U17135 ( .A(n15495), .ZN(n15563) );
  INV_X1 U17136 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n15496) );
  AOI22_X1 U17137 ( .A1(n15561), .A2(n15563), .B1(n15496), .B2(n15559), .ZN(
        P2_U3430) );
  INV_X1 U17138 ( .A(n15501), .ZN(n15503) );
  AOI21_X1 U17139 ( .B1(n15539), .B2(n6672), .A(n15497), .ZN(n15499) );
  OAI211_X1 U17140 ( .C1(n15554), .C2(n15501), .A(n15500), .B(n15499), .ZN(
        n15502) );
  AOI21_X1 U17141 ( .B1(n15558), .B2(n15503), .A(n15502), .ZN(n15564) );
  INV_X1 U17142 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n15504) );
  AOI22_X1 U17143 ( .A1(n15561), .A2(n15564), .B1(n15504), .B2(n15559), .ZN(
        P2_U3433) );
  AOI21_X1 U17144 ( .B1(n9794), .B2(n15554), .A(n15505), .ZN(n15510) );
  OAI21_X1 U17145 ( .B1(n15507), .B2(n15548), .A(n15506), .ZN(n15508) );
  NOR3_X1 U17146 ( .A1(n15510), .A2(n15509), .A3(n15508), .ZN(n15565) );
  INV_X1 U17147 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n15511) );
  AOI22_X1 U17148 ( .A1(n15561), .A2(n15565), .B1(n15511), .B2(n15559), .ZN(
        P2_U3445) );
  AOI21_X1 U17149 ( .B1(n15539), .B2(n15513), .A(n15512), .ZN(n15514) );
  OAI211_X1 U17150 ( .C1(n15516), .C2(n15554), .A(n15515), .B(n15514), .ZN(
        n15517) );
  INV_X1 U17151 ( .A(n15517), .ZN(n15567) );
  INV_X1 U17152 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n15518) );
  AOI22_X1 U17153 ( .A1(n15561), .A2(n15567), .B1(n15518), .B2(n15559), .ZN(
        P2_U3448) );
  OAI211_X1 U17154 ( .C1(n15521), .C2(n15548), .A(n15520), .B(n15519), .ZN(
        n15525) );
  NOR2_X1 U17155 ( .A1(n15523), .A2(n15522), .ZN(n15524) );
  AOI211_X1 U17156 ( .C1(n15527), .C2(n15526), .A(n15525), .B(n15524), .ZN(
        n15568) );
  INV_X1 U17157 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n15528) );
  AOI22_X1 U17158 ( .A1(n15561), .A2(n15568), .B1(n15528), .B2(n15559), .ZN(
        P2_U3451) );
  AOI21_X1 U17159 ( .B1(n15539), .B2(n15530), .A(n15529), .ZN(n15531) );
  OAI21_X1 U17160 ( .B1(n15532), .B2(n15554), .A(n15531), .ZN(n15533) );
  AOI211_X1 U17161 ( .C1(n15558), .C2(n15535), .A(n15534), .B(n15533), .ZN(
        n15570) );
  INV_X1 U17162 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n15536) );
  AOI22_X1 U17163 ( .A1(n15561), .A2(n15570), .B1(n15536), .B2(n15559), .ZN(
        P2_U3454) );
  INV_X1 U17164 ( .A(n15541), .ZN(n15544) );
  AOI21_X1 U17165 ( .B1(n15539), .B2(n15538), .A(n15537), .ZN(n15540) );
  OAI21_X1 U17166 ( .B1(n15541), .B2(n15554), .A(n15540), .ZN(n15542) );
  AOI211_X1 U17167 ( .C1(n15558), .C2(n15544), .A(n15543), .B(n15542), .ZN(
        n15572) );
  INV_X1 U17168 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n15545) );
  AOI22_X1 U17169 ( .A1(n15561), .A2(n15572), .B1(n15545), .B2(n15559), .ZN(
        P2_U3457) );
  INV_X1 U17170 ( .A(n15555), .ZN(n15557) );
  OAI211_X1 U17171 ( .C1(n15549), .C2(n15548), .A(n15547), .B(n15546), .ZN(
        n15550) );
  AOI21_X1 U17172 ( .B1(n15552), .B2(n15551), .A(n15550), .ZN(n15553) );
  OAI21_X1 U17173 ( .B1(n15555), .B2(n15554), .A(n15553), .ZN(n15556) );
  AOI21_X1 U17174 ( .B1(n15558), .B2(n15557), .A(n15556), .ZN(n15575) );
  INV_X1 U17175 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n15560) );
  AOI22_X1 U17176 ( .A1(n15561), .A2(n15575), .B1(n15560), .B2(n15559), .ZN(
        P2_U3460) );
  INV_X1 U17177 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n15562) );
  AOI22_X1 U17178 ( .A1(n15576), .A2(n15563), .B1(n15562), .B2(n15573), .ZN(
        P2_U3499) );
  AOI22_X1 U17179 ( .A1(n15576), .A2(n15564), .B1(n9411), .B2(n15573), .ZN(
        P2_U3500) );
  AOI22_X1 U17180 ( .A1(n15576), .A2(n15565), .B1(n9419), .B2(n15573), .ZN(
        P2_U3504) );
  AOI22_X1 U17181 ( .A1(n15576), .A2(n15567), .B1(n15566), .B2(n15573), .ZN(
        P2_U3505) );
  AOI22_X1 U17182 ( .A1(n15576), .A2(n15568), .B1(n9487), .B2(n15573), .ZN(
        P2_U3506) );
  AOI22_X1 U17183 ( .A1(n15576), .A2(n15570), .B1(n15569), .B2(n15573), .ZN(
        P2_U3507) );
  AOI22_X1 U17184 ( .A1(n15576), .A2(n15572), .B1(n15571), .B2(n15573), .ZN(
        P2_U3508) );
  AOI22_X1 U17185 ( .A1(n15576), .A2(n15575), .B1(n15574), .B2(n15573), .ZN(
        P2_U3509) );
  NOR2_X1 U17186 ( .A1(n15577), .A2(n15674), .ZN(P3_U3150) );
  INV_X1 U17187 ( .A(n15578), .ZN(n15590) );
  OAI21_X1 U17188 ( .B1(n15581), .B2(n15580), .A(n15579), .ZN(n15589) );
  INV_X1 U17189 ( .A(n11379), .ZN(n15587) );
  AOI21_X1 U17190 ( .B1(n15584), .B2(n15583), .A(n15582), .ZN(n15586) );
  NOR3_X1 U17191 ( .A1(n15587), .A2(n15586), .A3(n15585), .ZN(n15588) );
  AOI211_X1 U17192 ( .C1(n15591), .C2(n15590), .A(n15589), .B(n15588), .ZN(
        n15592) );
  OAI21_X1 U17193 ( .B1(n15594), .B2(n15593), .A(n15592), .ZN(P3_U3157) );
  NAND2_X1 U17194 ( .A1(n15596), .A2(n15595), .ZN(n15597) );
  XNOR2_X1 U17195 ( .A(n15598), .B(n15597), .ZN(n15599) );
  NOR2_X1 U17196 ( .A1(n15599), .A2(n15661), .ZN(n15610) );
  AOI21_X1 U17197 ( .B1(n15601), .B2(n15600), .A(n6806), .ZN(n15608) );
  OAI21_X1 U17198 ( .B1(P3_REG1_REG_9__SCAN_IN), .B2(n15603), .A(n15602), .ZN(
        n15606) );
  AOI22_X1 U17199 ( .A1(n15606), .A2(n15679), .B1(n15605), .B2(n15604), .ZN(
        n15607) );
  OAI21_X1 U17200 ( .B1(n15608), .B2(n15687), .A(n15607), .ZN(n15609) );
  NOR2_X1 U17201 ( .A1(n15610), .A2(n15609), .ZN(n15612) );
  NAND2_X1 U17202 ( .A1(P3_REG3_REG_9__SCAN_IN), .A2(P3_U3151), .ZN(n15611) );
  OAI211_X1 U17203 ( .C1(n15614), .C2(n15613), .A(n15612), .B(n15611), .ZN(
        P3_U3191) );
  AOI21_X1 U17204 ( .B1(n11420), .B2(n15616), .A(n15615), .ZN(n15631) );
  OAI21_X1 U17205 ( .B1(P3_REG1_REG_11__SCAN_IN), .B2(n15618), .A(n15617), 
        .ZN(n15624) );
  NOR2_X1 U17206 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15619), .ZN(n15620) );
  AOI21_X1 U17207 ( .B1(n15674), .B2(P3_ADDR_REG_11__SCAN_IN), .A(n15620), 
        .ZN(n15621) );
  OAI21_X1 U17208 ( .B1(n15677), .B2(n15622), .A(n15621), .ZN(n15623) );
  AOI21_X1 U17209 ( .B1(n15624), .B2(n15679), .A(n15623), .ZN(n15630) );
  AOI21_X1 U17210 ( .B1(n15627), .B2(n15626), .A(n15625), .ZN(n15628) );
  OR2_X1 U17211 ( .A1(n15628), .A2(n15661), .ZN(n15629) );
  OAI211_X1 U17212 ( .C1(n15631), .C2(n15687), .A(n15630), .B(n15629), .ZN(
        P3_U3193) );
  AOI21_X1 U17213 ( .B1(n6805), .B2(n15633), .A(n15632), .ZN(n15648) );
  OAI21_X1 U17214 ( .B1(n15636), .B2(n15635), .A(n15634), .ZN(n15642) );
  INV_X1 U17215 ( .A(n15637), .ZN(n15638) );
  AOI21_X1 U17216 ( .B1(n15674), .B2(P3_ADDR_REG_12__SCAN_IN), .A(n15638), 
        .ZN(n15639) );
  OAI21_X1 U17217 ( .B1(n15677), .B2(n15640), .A(n15639), .ZN(n15641) );
  AOI21_X1 U17218 ( .B1(n15642), .B2(n15679), .A(n15641), .ZN(n15647) );
  OAI211_X1 U17219 ( .C1(n15645), .C2(n15644), .A(n15643), .B(n15681), .ZN(
        n15646) );
  OAI211_X1 U17220 ( .C1(n15648), .C2(n15687), .A(n15647), .B(n15646), .ZN(
        P3_U3194) );
  AOI21_X1 U17221 ( .B1(n8190), .B2(n15650), .A(n15649), .ZN(n15665) );
  OAI21_X1 U17222 ( .B1(P3_REG1_REG_13__SCAN_IN), .B2(n15652), .A(n15651), 
        .ZN(n15657) );
  AND2_X1 U17223 ( .A1(P3_U3151), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n15653) );
  AOI21_X1 U17224 ( .B1(n15674), .B2(P3_ADDR_REG_13__SCAN_IN), .A(n15653), 
        .ZN(n15654) );
  OAI21_X1 U17225 ( .B1(n15677), .B2(n15655), .A(n15654), .ZN(n15656) );
  AOI21_X1 U17226 ( .B1(n15657), .B2(n15679), .A(n15656), .ZN(n15664) );
  AOI21_X1 U17227 ( .B1(n15660), .B2(n15659), .A(n15658), .ZN(n15662) );
  OR2_X1 U17228 ( .A1(n15662), .A2(n15661), .ZN(n15663) );
  OAI211_X1 U17229 ( .C1(n15665), .C2(n15687), .A(n15664), .B(n15663), .ZN(
        P3_U3195) );
  AOI21_X1 U17230 ( .B1(n15668), .B2(n15667), .A(n15666), .ZN(n15688) );
  OAI21_X1 U17231 ( .B1(n15671), .B2(n15670), .A(n15669), .ZN(n15680) );
  INV_X1 U17232 ( .A(n15672), .ZN(n15673) );
  AOI21_X1 U17233 ( .B1(n15674), .B2(P3_ADDR_REG_14__SCAN_IN), .A(n15673), 
        .ZN(n15675) );
  OAI21_X1 U17234 ( .B1(n15677), .B2(n15676), .A(n15675), .ZN(n15678) );
  AOI21_X1 U17235 ( .B1(n15680), .B2(n15679), .A(n15678), .ZN(n15686) );
  OAI211_X1 U17236 ( .C1(n15684), .C2(n15683), .A(n15682), .B(n15681), .ZN(
        n15685) );
  OAI211_X1 U17237 ( .C1(n15688), .C2(n15687), .A(n15686), .B(n15685), .ZN(
        P3_U3196) );
  INV_X1 U17238 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n15702) );
  XNOR2_X1 U17239 ( .A(n15689), .B(n15692), .ZN(n15698) );
  INV_X1 U17240 ( .A(n15698), .ZN(n15730) );
  NOR2_X1 U17241 ( .A1(n15690), .A2(n15744), .ZN(n15729) );
  INV_X1 U17242 ( .A(n15729), .ZN(n15691) );
  OAI22_X1 U17243 ( .A1(n15691), .A2(n15712), .B1(n10486), .B2(n15711), .ZN(
        n15699) );
  XNOR2_X1 U17244 ( .A(n15693), .B(n15692), .ZN(n15696) );
  AOI21_X1 U17245 ( .B1(n15696), .B2(n15695), .A(n15694), .ZN(n15697) );
  OAI21_X1 U17246 ( .B1(n15698), .B2(n15766), .A(n15697), .ZN(n15728) );
  AOI211_X1 U17247 ( .C1(n15700), .C2(n15730), .A(n15699), .B(n15728), .ZN(
        n15701) );
  AOI22_X1 U17248 ( .A1(n15703), .A2(n15702), .B1(n15701), .B2(n15719), .ZN(
        P3_U3231) );
  XNOR2_X1 U17249 ( .A(n15705), .B(n15704), .ZN(n15715) );
  XNOR2_X1 U17250 ( .A(n15707), .B(n15706), .ZN(n15709) );
  NOR2_X1 U17251 ( .A1(n15709), .A2(n15708), .ZN(n15724) );
  NAND2_X1 U17252 ( .A1(n7129), .A2(n15770), .ZN(n15722) );
  OAI22_X1 U17253 ( .A1(n15722), .A2(n15712), .B1(n15711), .B2(n15710), .ZN(
        n15713) );
  NOR3_X1 U17254 ( .A1(n15724), .A2(n15721), .A3(n15713), .ZN(n15714) );
  OAI21_X1 U17255 ( .B1(n15766), .B2(n15715), .A(n15714), .ZN(n15717) );
  INV_X1 U17256 ( .A(n15715), .ZN(n15726) );
  AOI22_X1 U17257 ( .A1(n15717), .A2(n15719), .B1(n15716), .B2(n15726), .ZN(
        n15718) );
  OAI21_X1 U17258 ( .B1(n15720), .B2(n15719), .A(n15718), .ZN(P3_U3232) );
  INV_X1 U17259 ( .A(n15721), .ZN(n15723) );
  NAND2_X1 U17260 ( .A1(n15723), .A2(n15722), .ZN(n15725) );
  AOI211_X1 U17261 ( .C1(n15746), .C2(n15726), .A(n15725), .B(n15724), .ZN(
        n15775) );
  INV_X1 U17262 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n15727) );
  AOI22_X1 U17263 ( .A1(n15773), .A2(n15775), .B1(n15727), .B2(n15771), .ZN(
        P3_U3393) );
  AOI211_X1 U17264 ( .C1(n15730), .C2(n15750), .A(n15729), .B(n15728), .ZN(
        n15777) );
  INV_X1 U17265 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n15731) );
  AOI22_X1 U17266 ( .A1(n15773), .A2(n15777), .B1(n15731), .B2(n15771), .ZN(
        P3_U3396) );
  NOR2_X1 U17267 ( .A1(n15732), .A2(n15744), .ZN(n15734) );
  AOI211_X1 U17268 ( .C1(n15750), .C2(n15735), .A(n15734), .B(n15733), .ZN(
        n15778) );
  AOI22_X1 U17269 ( .A1(n15773), .A2(n15778), .B1(n8046), .B2(n15771), .ZN(
        P3_U3399) );
  AOI22_X1 U17270 ( .A1(n15737), .A2(n15750), .B1(n15770), .B2(n15736), .ZN(
        n15738) );
  AND2_X1 U17271 ( .A1(n15739), .A2(n15738), .ZN(n15779) );
  INV_X1 U17272 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n15740) );
  AOI22_X1 U17273 ( .A1(n15773), .A2(n15779), .B1(n15740), .B2(n15771), .ZN(
        P3_U3402) );
  INV_X1 U17274 ( .A(n15741), .ZN(n15747) );
  OAI21_X1 U17275 ( .B1(n15744), .B2(n15743), .A(n15742), .ZN(n15745) );
  AOI21_X1 U17276 ( .B1(n15747), .B2(n15746), .A(n15745), .ZN(n15781) );
  AOI22_X1 U17277 ( .A1(n15773), .A2(n15781), .B1(n15748), .B2(n15771), .ZN(
        P3_U3405) );
  AOI22_X1 U17278 ( .A1(n15751), .A2(n15750), .B1(n15770), .B2(n15749), .ZN(
        n15752) );
  AND2_X1 U17279 ( .A1(n15753), .A2(n15752), .ZN(n15783) );
  INV_X1 U17280 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n15754) );
  AOI22_X1 U17281 ( .A1(n15773), .A2(n15783), .B1(n15754), .B2(n15771), .ZN(
        P3_U3408) );
  AOI21_X1 U17282 ( .B1(n15770), .B2(n15756), .A(n15755), .ZN(n15757) );
  OAI21_X1 U17283 ( .B1(n15765), .B2(n15758), .A(n15757), .ZN(n15759) );
  AOI21_X1 U17284 ( .B1(n15761), .B2(n15760), .A(n15759), .ZN(n15785) );
  INV_X1 U17285 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n15762) );
  AOI22_X1 U17286 ( .A1(n15773), .A2(n15785), .B1(n15762), .B2(n15771), .ZN(
        P3_U3411) );
  INV_X1 U17287 ( .A(n15763), .ZN(n15768) );
  AOI21_X1 U17288 ( .B1(n15766), .B2(n15765), .A(n15764), .ZN(n15767) );
  AOI211_X1 U17289 ( .C1(n15770), .C2(n15769), .A(n15768), .B(n15767), .ZN(
        n15787) );
  INV_X1 U17290 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n15772) );
  AOI22_X1 U17291 ( .A1(n15773), .A2(n15787), .B1(n15772), .B2(n15771), .ZN(
        P3_U3414) );
  INV_X1 U17292 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n15774) );
  AOI22_X1 U17293 ( .A1(n15788), .A2(n15775), .B1(n15774), .B2(n15786), .ZN(
        P3_U3460) );
  AOI22_X1 U17294 ( .A1(n15788), .A2(n15777), .B1(n15776), .B2(n15786), .ZN(
        P3_U3461) );
  AOI22_X1 U17295 ( .A1(n15788), .A2(n15778), .B1(n10284), .B2(n15786), .ZN(
        P3_U3462) );
  AOI22_X1 U17296 ( .A1(n15788), .A2(n15779), .B1(n8060), .B2(n15786), .ZN(
        P3_U3463) );
  INV_X1 U17297 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n15780) );
  AOI22_X1 U17298 ( .A1(n15788), .A2(n15781), .B1(n15780), .B2(n15786), .ZN(
        P3_U3464) );
  AOI22_X1 U17299 ( .A1(n15788), .A2(n15783), .B1(n15782), .B2(n15786), .ZN(
        P3_U3465) );
  AOI22_X1 U17300 ( .A1(n15788), .A2(n15785), .B1(n15784), .B2(n15786), .ZN(
        P3_U3466) );
  AOI22_X1 U17301 ( .A1(n15788), .A2(n15787), .B1(n8117), .B2(n15786), .ZN(
        P3_U3467) );
  OAI21_X1 U17302 ( .B1(n15791), .B2(n15790), .A(n15789), .ZN(SUB_1596_U59) );
  OAI21_X1 U17303 ( .B1(n15794), .B2(n15793), .A(n15792), .ZN(SUB_1596_U58) );
  XOR2_X1 U17304 ( .A(P2_ADDR_REG_0__SCAN_IN), .B(n15795), .Z(SUB_1596_U53) );
  AOI21_X1 U17305 ( .B1(n15798), .B2(n15797), .A(n15796), .ZN(SUB_1596_U56) );
  OAI21_X1 U17306 ( .B1(n15801), .B2(n15800), .A(n15799), .ZN(n15802) );
  XNOR2_X1 U17307 ( .A(n15802), .B(P2_ADDR_REG_3__SCAN_IN), .ZN(SUB_1596_U60)
         );
  AOI21_X1 U17308 ( .B1(n15805), .B2(n15804), .A(n15803), .ZN(SUB_1596_U5) );
  CLKBUF_X1 U7419 ( .A(n10624), .Z(n13075) );
  CLKBUF_X1 U7444 ( .A(n8751), .Z(n6660) );
  OR2_X1 U7478 ( .A1(n14974), .A2(n15216), .ZN(n14975) );
  CLKBUF_X1 U8465 ( .A(n8386), .Z(n7128) );
  AND2_X2 U12202 ( .A1(n9620), .A2(n9619), .ZN(n10117) );
endmodule

