

module b14_C_SARLock_k_128_5 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, U3352, 
        U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343, U3342, 
        U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333, U3332, 
        U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323, U3322, 
        U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315, U3314, 
        U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305, U3304, 
        U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295, U3294, 
        U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477, U3479, 
        U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497, U3499, 
        U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511, U3512, 
        U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521, U3522, 
        U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531, U3532, 
        U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541, U3542, 
        U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289, U3288, 
        U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279, U3278, 
        U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269, U3268, 
        U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260, U3259, 
        U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250, U3249, 
        U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240, U3550, 
        U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559, U3560, 
        U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569, U3570, 
        U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579, U3580, 
        U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232, U3231, 
        U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222, U3221, 
        U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212, U3211, 
        U3210, U3149, U3148, U4043 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190,
         n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200,
         n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210,
         n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220,
         n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230,
         n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240,
         n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250,
         n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260,
         n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270,
         n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280,
         n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290,
         n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300,
         n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310,
         n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320,
         n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330,
         n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340,
         n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350,
         n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360,
         n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370,
         n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380,
         n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390,
         n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400,
         n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410,
         n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420,
         n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430,
         n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440,
         n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450,
         n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460,
         n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470,
         n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480,
         n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490,
         n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500,
         n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510,
         n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520,
         n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530,
         n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540,
         n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550,
         n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560,
         n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570,
         n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580,
         n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590,
         n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600,
         n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610,
         n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620,
         n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630,
         n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640,
         n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650,
         n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660,
         n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670,
         n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680,
         n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690,
         n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700,
         n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710,
         n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720,
         n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730,
         n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740,
         n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750,
         n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760,
         n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770,
         n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780,
         n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790,
         n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800,
         n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810,
         n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820,
         n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830,
         n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840,
         n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850,
         n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860,
         n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870,
         n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880,
         n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890,
         n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900,
         n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910,
         n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920,
         n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930,
         n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940,
         n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950,
         n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960,
         n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970,
         n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980,
         n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990,
         n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000,
         n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010,
         n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020,
         n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030,
         n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040,
         n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050,
         n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060,
         n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070,
         n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080,
         n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090,
         n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100,
         n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110,
         n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120,
         n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130,
         n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140,
         n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150,
         n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160,
         n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170,
         n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180,
         n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190,
         n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200,
         n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210,
         n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220,
         n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230,
         n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240,
         n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250,
         n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260,
         n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270,
         n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280,
         n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290,
         n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300,
         n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310,
         n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320,
         n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330,
         n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340,
         n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350,
         n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360,
         n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370,
         n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380,
         n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390,
         n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400,
         n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410,
         n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420,
         n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430,
         n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440,
         n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450,
         n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460,
         n3461, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471,
         n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481,
         n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491,
         n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501,
         n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511,
         n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521,
         n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531,
         n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541,
         n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551,
         n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561,
         n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571,
         n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581,
         n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591,
         n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601,
         n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611,
         n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621,
         n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631,
         n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641,
         n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651,
         n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661,
         n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671,
         n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681,
         n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691,
         n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701,
         n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711,
         n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721,
         n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731,
         n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741,
         n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751,
         n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761,
         n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771,
         n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781,
         n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791,
         n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801,
         n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811,
         n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821,
         n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831,
         n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841,
         n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851,
         n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861,
         n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871,
         n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881,
         n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891,
         n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901,
         n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911,
         n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921,
         n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931,
         n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941,
         n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951,
         n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961,
         n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971,
         n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981,
         n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991,
         n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001,
         n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011,
         n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021,
         n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031,
         n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041,
         n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051,
         n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061,
         n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071,
         n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081,
         n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091,
         n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101,
         n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111,
         n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121,
         n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131,
         n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141,
         n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151,
         n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161,
         n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171,
         n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181,
         n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191,
         n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201,
         n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211,
         n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221,
         n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231,
         n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241,
         n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251,
         n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261,
         n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271,
         n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281,
         n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291,
         n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301,
         n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311,
         n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321,
         n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331,
         n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341,
         n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351,
         n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361,
         n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371,
         n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381,
         n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391,
         n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401,
         n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411,
         n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421,
         n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431,
         n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441,
         n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451,
         n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461,
         n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471,
         n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481,
         n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491,
         n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501,
         n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511,
         n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521,
         n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531,
         n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541,
         n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551,
         n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561,
         n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571,
         n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581,
         n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591,
         n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601,
         n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611,
         n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621,
         n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631,
         n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641,
         n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651,
         n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661,
         n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671,
         n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681,
         n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691,
         n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701,
         n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711,
         n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721,
         n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731,
         n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741,
         n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751,
         n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761,
         n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771,
         n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781,
         n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791,
         n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801,
         n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811,
         n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821,
         n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831,
         n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841,
         n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851,
         n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861,
         n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871,
         n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881,
         n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891,
         n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901,
         n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911,
         n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920;

  CLKBUF_X2 U2424 ( .A(U4043), .Z(n2181) );
  INV_X2 U2425 ( .A(n2798), .ZN(n2767) );
  NAND3_X2 U2426 ( .A1(n4710), .A2(n4711), .A3(n3281), .ZN(n2417) );
  NAND4_X1 U2427 ( .A1(n2414), .A2(n2413), .A3(n2412), .A4(n2411), .ZN(n4091)
         );
  BUF_X1 U2428 ( .A(n2419), .Z(n2804) );
  NAND2_X1 U2429 ( .A1(n4071), .A2(n4005), .ZN(n3425) );
  OAI22_X1 U2430 ( .A1(n3616), .A2(n2864), .B1(n3621), .B2(n3676), .ZN(n3677)
         );
  CLKBUF_X2 U2431 ( .A(n2430), .Z(n3302) );
  NOR2_X1 U2432 ( .A1(n2375), .A2(n4708), .ZN(n2430) );
  INV_X1 U2433 ( .A(n3551), .ZN(n4879) );
  CLKBUF_X2 U2434 ( .A(n2415), .Z(n3929) );
  AND4_X1 U2436 ( .A1(n2434), .A2(n2433), .A3(n2432), .A4(n2431), .ZN(n2852)
         );
  OR2_X1 U2437 ( .A1(n4416), .A2(n4419), .ZN(n4417) );
  NOR2_X1 U2438 ( .A1(n2437), .A2(n2436), .ZN(n4719) );
  INV_X1 U2439 ( .A(n2751), .ZN(n2406) );
  OAI21_X2 U2440 ( .B1(n3502), .B2(n3497), .A(n4029), .ZN(n3617) );
  NAND2_X2 U2441 ( .A1(n2406), .A2(n2405), .ZN(n2755) );
  INV_X2 U2442 ( .A(n2802), .ZN(n2753) );
  XNOR2_X1 U2443 ( .A(n2393), .B(n2367), .ZN(n4071) );
  XNOR2_X1 U2444 ( .A(n2394), .B(IR_REG_21__SCAN_IN), .ZN(n4005) );
  XNOR2_X1 U2445 ( .A(n2386), .B(n2385), .ZN(n2774) );
  XNOR2_X1 U2446 ( .A(n2371), .B(IR_REG_29__SCAN_IN), .ZN(n4708) );
  OAI21_X1 U2447 ( .B1(n2387), .B2(n2348), .A(IR_REG_31__SCAN_IN), .ZN(n3243)
         );
  AND4_X1 U2448 ( .A1(n2480), .A2(n2603), .A3(n2464), .A4(n2363), .ZN(n2305)
         );
  AND2_X1 U2449 ( .A1(n2366), .A2(n2345), .ZN(n2344) );
  AND4_X1 U2450 ( .A1(n2222), .A2(n2223), .A3(n2221), .A4(n2224), .ZN(n2304)
         );
  INV_X1 U2451 ( .A(IR_REG_15__SCAN_IN), .ZN(n2642) );
  INV_X1 U2452 ( .A(IR_REG_20__SCAN_IN), .ZN(n2367) );
  INV_X1 U2453 ( .A(IR_REG_3__SCAN_IN), .ZN(n2464) );
  NOR2_X1 U2454 ( .A1(IR_REG_11__SCAN_IN), .A2(IR_REG_12__SCAN_IN), .ZN(n2224)
         );
  INV_X1 U2455 ( .A(IR_REG_0__SCAN_IN), .ZN(n2225) );
  AOI21_X1 U2456 ( .B1(n2320), .B2(n2884), .A(n2319), .ZN(n2318) );
  INV_X1 U2457 ( .A(n3966), .ZN(n2319) );
  INV_X1 U2458 ( .A(n2883), .ZN(n2320) );
  AOI21_X1 U2459 ( .B1(n4091), .B2(n2798), .A(n2416), .ZN(n2423) );
  INV_X1 U2460 ( .A(n3511), .ZN(n2405) );
  OR2_X1 U2461 ( .A1(n4374), .A2(n4572), .ZN(n2881) );
  NAND2_X1 U2462 ( .A1(n2871), .A2(n2870), .ZN(n3716) );
  INV_X1 U2463 ( .A(IR_REG_30__SCAN_IN), .ZN(n2372) );
  INV_X1 U2464 ( .A(n3284), .ZN(n2784) );
  NAND2_X1 U2465 ( .A1(n2309), .A2(n2313), .ZN(n2307) );
  OR2_X1 U2466 ( .A1(n3904), .A2(n3900), .ZN(n2299) );
  NAND2_X1 U2467 ( .A1(n3473), .A2(n3472), .ZN(n2276) );
  AOI21_X1 U2468 ( .B1(n2291), .B2(n2203), .A(n2651), .ZN(n2289) );
  INV_X1 U2469 ( .A(n2649), .ZN(n2293) );
  BUF_X1 U2470 ( .A(n2446), .Z(n2822) );
  NAND2_X1 U2471 ( .A1(n3290), .A2(n4708), .ZN(n2446) );
  NAND2_X1 U2472 ( .A1(n4739), .A2(n4740), .ZN(n4738) );
  XNOR2_X1 U2473 ( .A(n3584), .B(n2270), .ZN(n4751) );
  NAND2_X1 U2474 ( .A1(n2891), .A2(n2335), .ZN(n2334) );
  NOR2_X1 U2475 ( .A1(n2893), .A2(n2336), .ZN(n2335) );
  INV_X1 U2476 ( .A(n2890), .ZN(n2336) );
  NAND2_X1 U2477 ( .A1(n2229), .A2(n2228), .ZN(n2337) );
  AOI21_X1 U2478 ( .B1(n2230), .B2(n2232), .A(n2208), .ZN(n2228) );
  NAND2_X1 U2479 ( .A1(n4474), .A2(n2358), .ZN(n2340) );
  OAI21_X1 U2480 ( .B1(n4204), .B2(n2899), .A(n2898), .ZN(n3235) );
  AND2_X1 U2481 ( .A1(n2351), .A2(n2368), .ZN(n2258) );
  INV_X1 U2482 ( .A(IR_REG_22__SCAN_IN), .ZN(n2368) );
  INV_X1 U2483 ( .A(IR_REG_28__SCAN_IN), .ZN(n2824) );
  NAND2_X1 U2484 ( .A1(n2185), .A2(n2342), .ZN(n2341) );
  INV_X1 U2485 ( .A(IR_REG_21__SCAN_IN), .ZN(n2342) );
  INV_X1 U2486 ( .A(IR_REG_19__SCAN_IN), .ZN(n2401) );
  NOR2_X1 U2487 ( .A1(REG1_REG_16__SCAN_IN), .A2(n4805), .ZN(n4806) );
  XNOR2_X1 U2488 ( .A(n3235), .B(n3964), .ZN(n3753) );
  NAND2_X1 U2489 ( .A1(n3804), .A2(n3805), .ZN(n2279) );
  AND2_X1 U2490 ( .A1(n3861), .A2(n2284), .ZN(n2283) );
  INV_X1 U2491 ( .A(n3860), .ZN(n2284) );
  NOR2_X1 U2492 ( .A1(n2283), .A2(n2282), .ZN(n2281) );
  INV_X1 U2493 ( .A(n3805), .ZN(n2282) );
  XNOR2_X1 U2494 ( .A(n2454), .B(n2753), .ZN(n2455) );
  NAND2_X1 U2495 ( .A1(n2453), .A2(n2452), .ZN(n2454) );
  INV_X1 U2496 ( .A(n2892), .ZN(n2333) );
  NAND2_X1 U2497 ( .A1(n4580), .A2(n4593), .ZN(n2878) );
  NOR2_X1 U2498 ( .A1(n2330), .A2(n2326), .ZN(n2323) );
  NAND3_X1 U2499 ( .A1(n3443), .A2(n2851), .A3(n3521), .ZN(n3519) );
  NAND2_X1 U2500 ( .A1(n2350), .A2(n2349), .ZN(n2348) );
  INV_X1 U2501 ( .A(IR_REG_26__SCAN_IN), .ZN(n2350) );
  INV_X1 U2502 ( .A(IR_REG_25__SCAN_IN), .ZN(n2349) );
  OR2_X1 U2503 ( .A1(n2383), .A2(n3293), .ZN(n2788) );
  INV_X1 U2504 ( .A(IR_REG_23__SCAN_IN), .ZN(n2787) );
  NOR2_X1 U2505 ( .A1(IR_REG_8__SCAN_IN), .A2(IR_REG_7__SCAN_IN), .ZN(n2222)
         );
  NOR2_X1 U2506 ( .A1(IR_REG_10__SCAN_IN), .A2(IR_REG_9__SCAN_IN), .ZN(n2223)
         );
  NOR2_X1 U2507 ( .A1(IR_REG_6__SCAN_IN), .A2(IR_REG_5__SCAN_IN), .ZN(n2221)
         );
  OR3_X1 U2508 ( .A1(n2539), .A2(IR_REG_7__SCAN_IN), .A3(IR_REG_8__SCAN_IN), 
        .ZN(n2555) );
  AND2_X1 U2509 ( .A1(n2815), .A2(n3425), .ZN(n2802) );
  OAI22_X1 U2510 ( .A1(n4614), .A2(n2755), .B1(n2767), .B2(n4604), .ZN(n3860)
         );
  OAI21_X1 U2511 ( .B1(n3878), .B2(n3879), .A(n3880), .ZN(n2578) );
  INV_X1 U2512 ( .A(n3870), .ZN(n2310) );
  INV_X1 U2513 ( .A(n3464), .ZN(n2439) );
  INV_X1 U2514 ( .A(n3769), .ZN(n2624) );
  INV_X1 U2515 ( .A(n3833), .ZN(n2287) );
  NAND2_X1 U2516 ( .A1(n2649), .A2(n2634), .ZN(n2292) );
  NOR2_X1 U2517 ( .A1(n2744), .A2(n3818), .ZN(n2758) );
  NAND2_X1 U2518 ( .A1(n3354), .A2(n3353), .ZN(n3356) );
  NOR2_X1 U2519 ( .A1(n3395), .A2(n3394), .ZN(n3579) );
  XNOR2_X1 U2520 ( .A(n3582), .B(n4870), .ZN(n4730) );
  OR2_X1 U2521 ( .A1(n3579), .A2(n2271), .ZN(n3582) );
  NOR2_X1 U2522 ( .A1(n3580), .A2(n3679), .ZN(n2271) );
  NAND2_X1 U2523 ( .A1(n4738), .A2(n2204), .ZN(n3565) );
  NAND2_X1 U2524 ( .A1(n4741), .A2(n2206), .ZN(n3584) );
  NAND2_X1 U2525 ( .A1(n4140), .A2(n2253), .ZN(n4143) );
  NAND2_X1 U2526 ( .A1(n4155), .A2(REG1_REG_13__SCAN_IN), .ZN(n2253) );
  NOR2_X1 U2527 ( .A1(n4790), .A2(n2272), .ZN(n4163) );
  AND2_X1 U2528 ( .A1(n4161), .A2(REG2_REG_15__SCAN_IN), .ZN(n2272) );
  OAI21_X1 U2529 ( .B1(n4216), .B2(n2897), .A(n2896), .ZN(n4204) );
  NAND2_X1 U2530 ( .A1(n4294), .A2(n4278), .ZN(n2889) );
  AOI21_X1 U2531 ( .B1(n2211), .B2(n2318), .A(n2231), .ZN(n2230) );
  INV_X1 U2532 ( .A(n3967), .ZN(n2231) );
  INV_X1 U2533 ( .A(n2881), .ZN(n2316) );
  INV_X1 U2534 ( .A(n2318), .ZN(n2232) );
  AND2_X1 U2535 ( .A1(n4053), .A2(n4274), .ZN(n4312) );
  NAND2_X1 U2536 ( .A1(n4375), .A2(n2882), .ZN(n2883) );
  INV_X1 U2537 ( .A(n2884), .ZN(n2321) );
  NAND2_X1 U2538 ( .A1(n4366), .A2(n2881), .ZN(n4344) );
  AND2_X1 U2539 ( .A1(n4571), .A2(n4581), .ZN(n2879) );
  NAND2_X1 U2540 ( .A1(n2190), .A2(n2202), .ZN(n2327) );
  OR2_X1 U2541 ( .A1(n4423), .A2(n2876), .ZN(n2877) );
  AOI21_X1 U2542 ( .B1(n2340), .B2(n2191), .A(n2209), .ZN(n4435) );
  INV_X1 U2543 ( .A(n2875), .ZN(n2239) );
  NAND2_X1 U2544 ( .A1(n4435), .A2(n4434), .ZN(n4433) );
  NAND2_X1 U2545 ( .A1(n3686), .A2(n2874), .ZN(n4474) );
  OAI21_X1 U2546 ( .B1(n2236), .B2(n2235), .A(n2233), .ZN(n2338) );
  INV_X1 U2547 ( .A(n2234), .ZN(n2233) );
  OAI21_X1 U2548 ( .B1(n2865), .B2(n2235), .A(n2868), .ZN(n2234) );
  INV_X1 U2549 ( .A(n3456), .ZN(n3446) );
  AND2_X1 U2550 ( .A1(n2404), .A2(n3974), .ZN(n3416) );
  NAND2_X1 U2551 ( .A1(n3246), .A2(n3932), .ZN(n4502) );
  AND2_X1 U2552 ( .A1(n4205), .A2(n3233), .ZN(n3246) );
  AND2_X1 U2553 ( .A1(n3416), .A2(n4071), .ZN(n4585) );
  NAND2_X1 U2554 ( .A1(n4722), .A2(n3299), .ZN(n4878) );
  NAND2_X1 U2555 ( .A1(n2772), .A2(n4710), .ZN(n3284) );
  NOR2_X1 U2556 ( .A1(n2348), .A2(n2347), .ZN(n2346) );
  NAND2_X1 U2557 ( .A1(n2396), .A2(n2369), .ZN(n2347) );
  XNOR2_X1 U2558 ( .A(n2788), .B(n2787), .ZN(n3300) );
  AND2_X1 U2559 ( .A1(n2344), .A2(n2195), .ZN(n2185) );
  AND2_X1 U2560 ( .A1(n2436), .A2(n2464), .ZN(n2481) );
  INV_X1 U2561 ( .A(IR_REG_1__SCAN_IN), .ZN(n2226) );
  OR2_X1 U2562 ( .A1(n2353), .A2(n3898), .ZN(n2302) );
  NOR2_X1 U2563 ( .A1(n2201), .A2(n2298), .ZN(n2297) );
  INV_X1 U2564 ( .A(n3901), .ZN(n2298) );
  INV_X1 U2565 ( .A(n4354), .ZN(n4553) );
  AND4_X1 U2566 ( .A1(n2739), .A2(n2738), .A3(n2737), .A4(n2736), .ZN(n4279)
         );
  INV_X1 U2567 ( .A(n4327), .ZN(n3873) );
  OR2_X1 U2568 ( .A1(n2830), .A2(n2826), .ZN(n3923) );
  INV_X1 U2569 ( .A(n4395), .ZN(n4572) );
  INV_X1 U2570 ( .A(n4409), .ZN(n4581) );
  INV_X1 U2571 ( .A(n4605), .ZN(n4423) );
  XNOR2_X1 U2572 ( .A(n3356), .B(n4717), .ZN(n3405) );
  NAND2_X1 U2573 ( .A1(n4742), .A2(n4743), .ZN(n4741) );
  NAND2_X1 U2574 ( .A1(n4763), .A2(n4764), .ZN(n4762) );
  XNOR2_X1 U2575 ( .A(n4143), .B(n4861), .ZN(n4787) );
  NAND2_X1 U2576 ( .A1(n4787), .A2(REG1_REG_14__SCAN_IN), .ZN(n4786) );
  XNOR2_X1 U2577 ( .A(n4163), .B(n4162), .ZN(n4802) );
  NAND2_X1 U2578 ( .A1(n4802), .A2(n4800), .ZN(n4801) );
  XNOR2_X1 U2579 ( .A(n2268), .B(n4177), .ZN(n4178) );
  NOR2_X1 U2580 ( .A1(n4175), .A2(n2220), .ZN(n2268) );
  NAND2_X1 U2581 ( .A1(n2248), .A2(n2244), .ZN(n2251) );
  NOR2_X1 U2582 ( .A1(n2245), .A2(n2219), .ZN(n2244) );
  NAND2_X1 U2583 ( .A1(n4818), .A2(n2249), .ZN(n2248) );
  AOI21_X1 U2584 ( .B1(n3749), .B2(n4585), .A(n3750), .ZN(n2943) );
  OR2_X1 U2585 ( .A1(n3753), .A2(n2214), .ZN(n2240) );
  INV_X1 U2586 ( .A(IR_REG_31__SCAN_IN), .ZN(n3293) );
  NOR2_X1 U2587 ( .A1(n3778), .A2(n3777), .ZN(n2313) );
  AND2_X1 U2589 ( .A1(n4258), .A2(n3965), .ZN(n4056) );
  NAND2_X1 U2590 ( .A1(n4759), .A2(n3567), .ZN(n3568) );
  INV_X1 U2591 ( .A(n4173), .ZN(n2252) );
  AND2_X1 U2592 ( .A1(n3969), .A2(n4224), .ZN(n4001) );
  NOR2_X1 U2593 ( .A1(n4481), .A2(n4461), .ZN(n2339) );
  INV_X1 U2594 ( .A(n2867), .ZN(n2235) );
  OR3_X1 U2595 ( .A1(n4283), .A2(n4254), .A3(n2936), .ZN(n2264) );
  NAND2_X1 U2596 ( .A1(n4357), .A2(n2256), .ZN(n2255) );
  NOR2_X1 U2597 ( .A1(n4326), .A2(n4374), .ZN(n2256) );
  OR2_X1 U2598 ( .A1(n4421), .A2(n4580), .ZN(n4388) );
  NAND2_X1 U2599 ( .A1(n2261), .A2(n3883), .ZN(n2260) );
  INV_X1 U2600 ( .A(n2262), .ZN(n2261) );
  NAND2_X1 U2601 ( .A1(n3726), .A2(n3740), .ZN(n2262) );
  INV_X1 U2602 ( .A(n3700), .ZN(n2911) );
  NOR2_X1 U2603 ( .A1(n3621), .A2(n2266), .ZN(n2265) );
  INV_X1 U2604 ( .A(n2267), .ZN(n2266) );
  NOR2_X1 U2605 ( .A1(n2858), .A2(n3506), .ZN(n2267) );
  NOR2_X1 U2606 ( .A1(IR_REG_24__SCAN_IN), .A2(IR_REG_23__SCAN_IN), .ZN(n2369)
         );
  INV_X1 U2607 ( .A(IR_REG_18__SCAN_IN), .ZN(n2366) );
  INV_X1 U2608 ( .A(IR_REG_16__SCAN_IN), .ZN(n2365) );
  INV_X1 U2609 ( .A(IR_REG_14__SCAN_IN), .ZN(n2363) );
  OAI21_X1 U2610 ( .B1(n2575), .B2(IR_REG_10__SCAN_IN), .A(IR_REG_31__SCAN_IN), 
        .ZN(n2586) );
  OR2_X1 U2611 ( .A1(n2555), .A2(IR_REG_9__SCAN_IN), .ZN(n2575) );
  INV_X1 U2612 ( .A(IR_REG_6__SCAN_IN), .ZN(n2508) );
  INV_X1 U2613 ( .A(IR_REG_4__SCAN_IN), .ZN(n2480) );
  INV_X1 U2614 ( .A(n2278), .ZN(n2277) );
  OAI22_X1 U2615 ( .A1(n2283), .A2(n2279), .B1(n2284), .B2(n3861), .ZN(n2278)
         );
  INV_X1 U2616 ( .A(n3542), .ZN(n3475) );
  NAND2_X1 U2617 ( .A1(n3608), .A2(n2295), .ZN(n2294) );
  AOI21_X1 U2618 ( .B1(n3631), .B2(n3630), .A(n2296), .ZN(n2295) );
  INV_X1 U2619 ( .A(n2489), .ZN(n2296) );
  AND2_X1 U2620 ( .A1(n2635), .A2(REG3_REG_16__SCAN_IN), .ZN(n2652) );
  INV_X1 U2621 ( .A(n2818), .ZN(n2752) );
  NOR2_X1 U2622 ( .A1(n3261), .A2(n2275), .ZN(n2274) );
  INV_X1 U2623 ( .A(n2458), .ZN(n2275) );
  INV_X1 U2624 ( .A(REG3_REG_9__SCAN_IN), .ZN(n2532) );
  NOR2_X1 U2625 ( .A1(n2579), .A2(n3809), .ZN(n2594) );
  AOI21_X1 U2626 ( .B1(n2189), .B2(n3852), .A(n2210), .ZN(n2312) );
  INV_X1 U2627 ( .A(n3793), .ZN(n2711) );
  INV_X1 U2628 ( .A(n3794), .ZN(n2712) );
  NAND2_X1 U2629 ( .A1(n3792), .A2(n2189), .ZN(n2311) );
  OAI22_X1 U2630 ( .A1(n2850), .A2(n2755), .B1(n2672), .B2(n3446), .ZN(n2426)
         );
  XNOR2_X1 U2631 ( .A(n2273), .B(n2802), .ZN(n2425) );
  OAI22_X1 U2632 ( .A1(n3446), .A2(n2751), .B1(n2752), .B2(n2850), .ZN(n2273)
         );
  XNOR2_X1 U2633 ( .A(n2438), .B(n2753), .ZN(n2441) );
  OAI22_X1 U2634 ( .A1(n2852), .A2(n2752), .B1(n4877), .B2(n2751), .ZN(n2438)
         );
  AND3_X1 U2635 ( .A1(REG3_REG_4__SCAN_IN), .A2(REG3_REG_3__SCAN_IN), .A3(
        REG3_REG_5__SCAN_IN), .ZN(n2490) );
  INV_X1 U2636 ( .A(REG3_REG_15__SCAN_IN), .ZN(n2626) );
  NOR2_X1 U2637 ( .A1(n2627), .A2(n2626), .ZN(n2635) );
  NAND2_X1 U2638 ( .A1(n2650), .A2(n2649), .ZN(n3913) );
  NOR2_X1 U2639 ( .A1(n2650), .A2(n2649), .ZN(n3915) );
  AND4_X1 U2640 ( .A1(n2507), .A2(n2506), .A3(n2505), .A4(n2504), .ZN(n3657)
         );
  NAND2_X1 U2641 ( .A1(n4116), .A2(n3335), .ZN(n3352) );
  XNOR2_X1 U2642 ( .A(n3384), .B(n4716), .ZN(n3367) );
  NAND2_X1 U2643 ( .A1(n4128), .A2(n2241), .ZN(n3384) );
  NAND2_X1 U2644 ( .A1(n2242), .A2(REG1_REG_5__SCAN_IN), .ZN(n2241) );
  INV_X1 U2645 ( .A(n4131), .ZN(n2242) );
  NAND2_X1 U2646 ( .A1(n4734), .A2(n3564), .ZN(n4739) );
  NAND2_X1 U2647 ( .A1(n4755), .A2(n3566), .ZN(n4760) );
  NAND2_X1 U2648 ( .A1(n4760), .A2(n4761), .ZN(n4759) );
  XNOR2_X1 U2649 ( .A(n3568), .B(n4863), .ZN(n4771) );
  NAND2_X1 U2650 ( .A1(n4762), .A2(n2205), .ZN(n3587) );
  NAND2_X1 U2651 ( .A1(n4811), .A2(n2269), .ZN(n4166) );
  OR2_X1 U2652 ( .A1(n4165), .A2(REG2_REG_17__SCAN_IN), .ZN(n2269) );
  NOR2_X1 U2653 ( .A1(n4166), .A2(n4167), .ZN(n4175) );
  NOR2_X1 U2654 ( .A1(n2252), .A2(n4148), .ZN(n2249) );
  NOR2_X1 U2655 ( .A1(n2252), .A2(n2246), .ZN(n2245) );
  NAND2_X1 U2656 ( .A1(n4817), .A2(n2247), .ZN(n2246) );
  INV_X1 U2657 ( .A(n4148), .ZN(n2247) );
  OR3_X1 U2658 ( .A1(n2793), .A2(n2839), .A3(n2827), .ZN(n4192) );
  NOR2_X1 U2659 ( .A1(n2200), .A2(n2333), .ZN(n2332) );
  INV_X1 U2660 ( .A(n4518), .ZN(n4217) );
  INV_X1 U2661 ( .A(REG3_REG_18__SCAN_IN), .ZN(n3085) );
  INV_X1 U2662 ( .A(n2325), .ZN(n2324) );
  OAI21_X1 U2663 ( .B1(n2327), .B2(n2326), .A(n2878), .ZN(n2325) );
  INV_X1 U2664 ( .A(REG3_REG_14__SCAN_IN), .ZN(n2608) );
  OR2_X1 U2665 ( .A1(n2609), .A2(n2608), .ZN(n2627) );
  OAI22_X1 U2666 ( .A1(n3716), .A2(n2872), .B1(n3884), .B2(n3726), .ZN(n3684)
         );
  OR2_X1 U2667 ( .A1(n3684), .A2(n3979), .ZN(n3686) );
  OR2_X1 U2668 ( .A1(n2533), .A2(n2532), .ZN(n2569) );
  INV_X1 U2669 ( .A(n4019), .ZN(n2865) );
  INV_X1 U2670 ( .A(n3677), .ZN(n2236) );
  INV_X1 U2671 ( .A(REG3_REG_7__SCAN_IN), .ZN(n3387) );
  AND2_X1 U2672 ( .A1(n2908), .A2(n4028), .ZN(n4019) );
  AND2_X1 U2673 ( .A1(n4018), .A2(n4031), .ZN(n3991) );
  AND2_X1 U2674 ( .A1(n4013), .A2(n4017), .ZN(n3495) );
  NAND2_X1 U2675 ( .A1(n3519), .A2(n2853), .ZN(n3482) );
  AND2_X1 U2676 ( .A1(n4012), .A2(n4009), .ZN(n3992) );
  NAND2_X1 U2677 ( .A1(n4010), .A2(n4007), .ZN(n3521) );
  OAI21_X1 U2678 ( .B1(n3243), .B2(n2824), .A(IR_REG_27__SCAN_IN), .ZN(n2314)
         );
  NAND2_X1 U2679 ( .A1(n2397), .A2(n2396), .ZN(n2315) );
  NOR2_X1 U2680 ( .A1(n3454), .A2(n3447), .ZN(n3441) );
  NAND2_X1 U2681 ( .A1(n2902), .A2(n3441), .ZN(n3443) );
  AND2_X1 U2682 ( .A1(n4585), .A2(n4179), .ZN(n3511) );
  NOR2_X1 U2683 ( .A1(n4884), .A2(n4005), .ZN(n2945) );
  OAI21_X1 U2684 ( .B1(n2786), .B2(n2785), .A(n2784), .ZN(n3420) );
  AND2_X1 U2685 ( .A1(n4002), .A2(n4004), .ZN(n3985) );
  INV_X1 U2686 ( .A(n3376), .ZN(n3447) );
  INV_X1 U2687 ( .A(n4505), .ZN(n4503) );
  NOR2_X1 U2688 ( .A1(n4502), .A2(n4503), .ZN(n4501) );
  NOR2_X1 U2689 ( .A1(n2183), .A2(n4509), .ZN(n4205) );
  INV_X1 U2690 ( .A(n4209), .ZN(n4509) );
  NOR3_X1 U2691 ( .A1(n4300), .A2(n4283), .A3(n4254), .ZN(n4252) );
  NOR2_X1 U2692 ( .A1(n4300), .A2(n4283), .ZN(n4284) );
  INV_X1 U2693 ( .A(n4293), .ZN(n4298) );
  OR2_X1 U2694 ( .A1(n2184), .A2(n4298), .ZN(n4300) );
  NAND2_X1 U2695 ( .A1(n2337), .A2(n2207), .ZN(n4546) );
  NOR2_X1 U2696 ( .A1(n4389), .A2(n2255), .ZN(n4334) );
  NOR2_X1 U2697 ( .A1(n4389), .A2(n4374), .ZN(n4368) );
  NOR3_X1 U2698 ( .A1(n4389), .A2(n2882), .A3(n4374), .ZN(n4359) );
  OR2_X1 U2699 ( .A1(n4388), .A2(n4571), .ZN(n4389) );
  NAND2_X1 U2700 ( .A1(n4441), .A2(n4422), .ZN(n4421) );
  AND2_X1 U2701 ( .A1(n4459), .A2(n4443), .ZN(n4441) );
  NOR2_X1 U2702 ( .A1(n4477), .A2(n4461), .ZN(n4459) );
  INV_X1 U2703 ( .A(n4491), .ZN(n4637) );
  NOR2_X1 U2704 ( .A1(n3696), .A2(n2262), .ZN(n4903) );
  NOR2_X1 U2705 ( .A1(n3696), .A2(n3710), .ZN(n3727) );
  OR2_X1 U2706 ( .A1(n3695), .A2(n2911), .ZN(n3696) );
  AND2_X1 U2707 ( .A1(n3556), .A2(n2265), .ZN(n3670) );
  NAND2_X1 U2708 ( .A1(n3556), .A2(n3555), .ZN(n3554) );
  NAND2_X1 U2709 ( .A1(n3556), .A2(n2267), .ZN(n3622) );
  AND2_X1 U2710 ( .A1(n3527), .A2(n3475), .ZN(n3556) );
  INV_X1 U2711 ( .A(n4878), .ZN(n4592) );
  INV_X1 U2712 ( .A(n4627), .ZN(n4876) );
  INV_X1 U2713 ( .A(n4615), .ZN(n4881) );
  AND2_X1 U2714 ( .A1(n2417), .A2(n4853), .ZN(n3296) );
  INV_X1 U2715 ( .A(IR_REG_24__SCAN_IN), .ZN(n2385) );
  NAND2_X1 U2716 ( .A1(n2384), .A2(IR_REG_31__SCAN_IN), .ZN(n2386) );
  INV_X1 U2717 ( .A(n2658), .ZN(n2343) );
  INV_X1 U2718 ( .A(IR_REG_2__SCAN_IN), .ZN(n2364) );
  INV_X1 U2719 ( .A(n2866), .ZN(n3671) );
  AND4_X1 U2720 ( .A1(n2574), .A2(n2573), .A3(n2572), .A4(n2571), .ZN(n4616)
         );
  AND4_X1 U2721 ( .A1(n2522), .A2(n2521), .A3(n2520), .A4(n2519), .ZN(n3741)
         );
  OAI21_X1 U2722 ( .B1(n3803), .B2(n3804), .A(n3805), .ZN(n3863) );
  NAND2_X1 U2723 ( .A1(n3929), .A2(DATAI_22_), .ZN(n4293) );
  NAND2_X1 U2724 ( .A1(n2311), .A2(n2312), .ZN(n3869) );
  INV_X1 U2725 ( .A(n4628), .ZN(n3883) );
  INV_X1 U2726 ( .A(n3532), .ZN(n4877) );
  XNOR2_X1 U2727 ( .A(n2441), .B(n2442), .ZN(n3464) );
  AOI21_X1 U2729 ( .B1(n2285), .B2(n2182), .A(n2286), .ZN(n3892) );
  INV_X1 U2730 ( .A(n2650), .ZN(n2285) );
  OR2_X1 U2731 ( .A1(n2819), .A2(n3377), .ZN(n3895) );
  AND4_X1 U2732 ( .A1(n2479), .A2(n2478), .A3(n2477), .A4(n2476), .ZN(n2859)
         );
  NAND2_X1 U2733 ( .A1(n3608), .A2(n2489), .ZN(n3633) );
  NAND2_X1 U2734 ( .A1(n3929), .A2(DATAI_26_), .ZN(n4518) );
  INV_X1 U2735 ( .A(n3895), .ZN(n3928) );
  AND2_X1 U2736 ( .A1(n2818), .A2(n2817), .ZN(n4078) );
  NAND2_X1 U2737 ( .A1(n2380), .A2(n2379), .ZN(n4520) );
  NAND4_X1 U2738 ( .A1(n2693), .A2(n2692), .A3(n2691), .A4(n2690), .ZN(n4354)
         );
  INV_X1 U2739 ( .A(n3741), .ZN(n3667) );
  INV_X1 U2740 ( .A(n3657), .ZN(n4087) );
  INV_X1 U2741 ( .A(n2859), .ZN(n4088) );
  INV_X1 U2742 ( .A(n2857), .ZN(n4089) );
  NAND4_X1 U2743 ( .A1(n2451), .A2(n2450), .A3(n2449), .A4(n2448), .ZN(n3551)
         );
  INV_X1 U2744 ( .A(n2850), .ZN(n3375) );
  NAND2_X1 U2745 ( .A1(n4117), .A2(n4118), .ZN(n4116) );
  XNOR2_X1 U2746 ( .A(n3362), .B(n3343), .ZN(n3344) );
  NAND2_X1 U2747 ( .A1(n3406), .A2(n2243), .ZN(n4129) );
  NAND2_X1 U2748 ( .A1(n3365), .A2(n4717), .ZN(n2243) );
  NAND2_X1 U2749 ( .A1(n4129), .A2(n4130), .ZN(n4128) );
  OAI21_X1 U2750 ( .B1(n3405), .B2(n3355), .A(n3357), .ZN(n4135) );
  NAND2_X1 U2751 ( .A1(n4729), .A2(n3583), .ZN(n4742) );
  XNOR2_X1 U2752 ( .A(n3565), .B(n2270), .ZN(n4756) );
  NAND2_X1 U2753 ( .A1(n4750), .A2(n3585), .ZN(n4763) );
  XNOR2_X1 U2754 ( .A(n3587), .B(n4863), .ZN(n4774) );
  NAND2_X1 U2755 ( .A1(n4786), .A2(n4144), .ZN(n4796) );
  NAND2_X1 U2756 ( .A1(n4801), .A2(n4164), .ZN(n4810) );
  NOR2_X1 U2757 ( .A1(n4147), .A2(n4806), .ZN(n4818) );
  AND2_X1 U2758 ( .A1(n4094), .A2(n4093), .ZN(n4816) );
  NOR2_X1 U2759 ( .A1(n4818), .A2(n4817), .ZN(n4819) );
  AND2_X1 U2760 ( .A1(n4094), .A2(n4079), .ZN(n4773) );
  INV_X1 U2761 ( .A(n4174), .ZN(n2250) );
  AND2_X1 U2762 ( .A1(n3338), .A2(n3336), .ZN(n4815) );
  INV_X1 U2763 ( .A(n4510), .ZN(n4238) );
  NAND2_X1 U2764 ( .A1(n3929), .A2(DATAI_27_), .ZN(n4209) );
  NAND2_X1 U2765 ( .A1(n2334), .A2(n2892), .ZN(n4233) );
  NAND2_X1 U2766 ( .A1(n2891), .A2(n2890), .ZN(n4250) );
  AND3_X1 U2767 ( .A1(n2750), .A2(n2749), .A3(n2748), .ZN(n4531) );
  NAND2_X1 U2768 ( .A1(n2337), .A2(n2885), .ZN(n4304) );
  OR2_X1 U2769 ( .A1(n4366), .A2(n2232), .ZN(n2227) );
  INV_X1 U2770 ( .A(n2317), .ZN(n4323) );
  AOI21_X1 U2771 ( .B1(n4344), .B2(n2883), .A(n2321), .ZN(n2317) );
  AND4_X1 U2772 ( .A1(n2669), .A2(n2668), .A3(n2667), .A4(n2666), .ZN(n4395)
         );
  AND4_X1 U2773 ( .A1(n2657), .A2(n2656), .A3(n2655), .A4(n2654), .ZN(n4409)
         );
  NAND2_X1 U2774 ( .A1(n4402), .A2(n4401), .ZN(n4400) );
  NAND2_X1 U2775 ( .A1(n2328), .A2(n2327), .ZN(n4402) );
  NAND2_X1 U2776 ( .A1(n4433), .A2(n2329), .ZN(n2328) );
  NAND2_X1 U2777 ( .A1(n4433), .A2(n2877), .ZN(n4420) );
  NAND2_X1 U2778 ( .A1(n2340), .A2(n2875), .ZN(n4458) );
  NAND2_X1 U2779 ( .A1(n2236), .A2(n2865), .ZN(n4897) );
  NAND2_X1 U2780 ( .A1(n4727), .A2(n3594), .ZN(n4415) );
  INV_X1 U2781 ( .A(n4415), .ZN(n4496) );
  INV_X1 U2782 ( .A(n4179), .ZN(n4379) );
  INV_X1 U2783 ( .A(n4825), .ZN(n4727) );
  MUX2_X1 U2784 ( .A(n4719), .B(DATAI_2_), .S(n2415), .Z(n3532) );
  NAND2_X1 U2785 ( .A1(n3296), .A2(n2945), .ZN(n4478) );
  AND2_X1 U2786 ( .A1(n2775), .A2(n2774), .ZN(n3288) );
  NAND2_X1 U2787 ( .A1(n3284), .A2(n3296), .ZN(n4847) );
  XNOR2_X1 U2788 ( .A(n2373), .B(IR_REG_30__SCAN_IN), .ZN(n3290) );
  NAND2_X1 U2789 ( .A1(n2383), .A2(n2186), .ZN(n2370) );
  XNOR2_X1 U2790 ( .A(n2825), .B(n2824), .ZN(n4722) );
  AND2_X1 U2791 ( .A1(n2383), .A2(n2346), .ZN(n2823) );
  AND2_X1 U2792 ( .A1(n3300), .A2(STATE_REG_SCAN_IN), .ZN(n4853) );
  XNOR2_X1 U2793 ( .A(n2400), .B(IR_REG_22__SCAN_IN), .ZN(n4712) );
  XNOR2_X1 U2794 ( .A(n2402), .B(n2401), .ZN(n4179) );
  NOR2_X1 U2795 ( .A1(n2658), .A2(IR_REG_17__SCAN_IN), .ZN(n2670) );
  INV_X1 U2796 ( .A(n4165), .ZN(n4855) );
  INV_X1 U2797 ( .A(n3577), .ZN(n4865) );
  INV_X1 U2798 ( .A(n3578), .ZN(n4868) );
  OAI22_X1 U2799 ( .A1(n2435), .A2(n2254), .B1(IR_REG_31__SCAN_IN), .B2(
        IR_REG_2__SCAN_IN), .ZN(n2437) );
  NAND2_X1 U2800 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_2__SCAN_IN), .ZN(n2254)
         );
  XNOR2_X1 U2801 ( .A(n2410), .B(IR_REG_1__SCAN_IN), .ZN(n4720) );
  NAND2_X1 U2802 ( .A1(n2303), .A2(n2301), .ZN(n2300) );
  OR2_X1 U2803 ( .A1(n4193), .A2(n4640), .ZN(n3254) );
  OAI211_X1 U2804 ( .C1(n2943), .C2(n3250), .A(n2240), .B(n2217), .ZN(n2331)
         );
  AND2_X1 U2805 ( .A1(n2291), .A2(n3832), .ZN(n2182) );
  OR3_X1 U2806 ( .A1(n4300), .A2(n2264), .A3(n4217), .ZN(n2183) );
  OR3_X1 U2807 ( .A1(n4389), .A2(n2255), .A3(n4550), .ZN(n2184) );
  AND2_X1 U2808 ( .A1(n2346), .A2(n2824), .ZN(n2186) );
  NAND2_X1 U2809 ( .A1(n2343), .A2(n2344), .ZN(n2391) );
  NAND2_X1 U2810 ( .A1(n2343), .A2(n2185), .ZN(n2187) );
  AND2_X1 U2811 ( .A1(n2560), .A2(n2547), .ZN(n2188) );
  NOR2_X1 U2812 ( .A1(n2357), .A2(n2710), .ZN(n2189) );
  INV_X1 U2813 ( .A(n4401), .ZN(n2326) );
  OR2_X1 U2814 ( .A1(n4404), .A2(n4591), .ZN(n2190) );
  NAND2_X1 U2815 ( .A1(n2548), .A2(n2547), .ZN(n3267) );
  NOR2_X1 U2816 ( .A1(n2239), .A2(n2339), .ZN(n2191) );
  OAI21_X1 U2817 ( .B1(n2289), .B2(n2288), .A(n2287), .ZN(n2286) );
  NAND2_X1 U2818 ( .A1(n3929), .A2(DATAI_24_), .ZN(n4530) );
  NAND2_X1 U2819 ( .A1(n2276), .A2(n2458), .ZN(n3258) );
  OR2_X1 U2820 ( .A1(n3631), .A2(n3630), .ZN(n2192) );
  AND2_X1 U2821 ( .A1(n2311), .A2(n2308), .ZN(n2193) );
  AND4_X1 U2822 ( .A1(n2463), .A2(n2462), .A3(n2461), .A4(n2460), .ZN(n2857)
         );
  NAND2_X1 U2823 ( .A1(n2227), .A2(n2230), .ZN(n4309) );
  AOI21_X1 U2824 ( .B1(n3841), .B2(n3844), .A(n2743), .ZN(n3813) );
  NOR2_X1 U2825 ( .A1(n4819), .A2(n4148), .ZN(n2194) );
  NAND2_X2 U2826 ( .A1(n2417), .A2(n3425), .ZN(n2751) );
  AND2_X1 U2827 ( .A1(n2401), .A2(n2367), .ZN(n2195) );
  AND3_X1 U2828 ( .A1(n2436), .A2(n2305), .A3(n2351), .ZN(n2196) );
  OR2_X1 U2829 ( .A1(n2658), .A2(n2341), .ZN(n2197) );
  INV_X1 U2830 ( .A(IR_REG_27__SCAN_IN), .ZN(n2396) );
  AND2_X1 U2831 ( .A1(n3662), .A2(n2192), .ZN(n2198) );
  AND2_X1 U2832 ( .A1(n2869), .A2(n2359), .ZN(n2199) );
  AND2_X1 U2833 ( .A1(n4449), .A2(n4451), .ZN(n3979) );
  NAND4_X1 U2834 ( .A1(n2727), .A2(n2726), .A3(n2725), .A4(n2724), .ZN(n4533)
         );
  NOR2_X1 U2835 ( .A1(n4218), .A2(n2936), .ZN(n2200) );
  XOR2_X1 U2836 ( .A(n2810), .B(n2808), .Z(n2201) );
  OAI21_X1 U2837 ( .B1(n2650), .B2(n2290), .A(n2289), .ZN(n3831) );
  NAND2_X1 U2838 ( .A1(n3268), .A2(n2565), .ZN(n3878) );
  NAND2_X1 U2839 ( .A1(n2280), .A2(n2277), .ZN(n3768) );
  AND4_X1 U2840 ( .A1(n2599), .A2(n2598), .A3(n2597), .A4(n2596), .ZN(n4614)
         );
  INV_X1 U2841 ( .A(n4614), .ZN(n4481) );
  AND2_X1 U2842 ( .A1(n4404), .A2(n4591), .ZN(n2202) );
  INV_X1 U2843 ( .A(n4632), .ZN(n4607) );
  AND4_X1 U2844 ( .A1(n2584), .A2(n2583), .A3(n2582), .A4(n2581), .ZN(n4632)
         );
  AND2_X1 U2845 ( .A1(n2293), .A2(n3916), .ZN(n2203) );
  INV_X1 U2846 ( .A(n2858), .ZN(n3555) );
  OR2_X1 U2847 ( .A1(n4868), .A2(n3734), .ZN(n2204) );
  OR2_X1 U2848 ( .A1(n4865), .A2(n3688), .ZN(n2205) );
  OR2_X1 U2849 ( .A1(n4868), .A2(n3643), .ZN(n2206) );
  INV_X1 U2850 ( .A(n2263), .ZN(n4243) );
  NOR2_X1 U2851 ( .A1(n4300), .A2(n2264), .ZN(n2263) );
  INV_X1 U2852 ( .A(n4329), .ZN(n4375) );
  AND4_X1 U2853 ( .A1(n2680), .A2(n2679), .A3(n2678), .A4(n2677), .ZN(n4329)
         );
  AND2_X1 U2854 ( .A1(n2887), .A2(n2885), .ZN(n2207) );
  NOR2_X1 U2855 ( .A1(n3873), .A2(n4314), .ZN(n2208) );
  AND2_X1 U2856 ( .A1(n4461), .A2(n4481), .ZN(n2209) );
  INV_X1 U2857 ( .A(n2330), .ZN(n2329) );
  NAND2_X1 U2858 ( .A1(n2190), .A2(n2877), .ZN(n2330) );
  AND2_X1 U2859 ( .A1(n2712), .A2(n2711), .ZN(n2210) );
  OR2_X1 U2860 ( .A1(n2321), .A2(n2316), .ZN(n2211) );
  INV_X1 U2861 ( .A(n2291), .ZN(n2290) );
  AND2_X1 U2862 ( .A1(n3824), .A2(n2292), .ZN(n2291) );
  INV_X1 U2863 ( .A(n2309), .ZN(n2308) );
  NAND2_X1 U2864 ( .A1(n2312), .A2(n2310), .ZN(n2309) );
  AND2_X1 U2865 ( .A1(n2313), .A2(n2189), .ZN(n2212) );
  NAND2_X1 U2866 ( .A1(n2355), .A2(n3918), .ZN(n2213) );
  AND2_X2 U2867 ( .A1(n3252), .A2(n3423), .ZN(n4910) );
  NAND2_X1 U2868 ( .A1(n3929), .A2(DATAI_25_), .ZN(n4244) );
  NAND2_X1 U2869 ( .A1(n3929), .A2(DATAI_21_), .ZN(n4314) );
  INV_X1 U2870 ( .A(n4895), .ZN(n4589) );
  NAND2_X1 U2871 ( .A1(n3929), .A2(DATAI_20_), .ZN(n4336) );
  OAI21_X1 U2872 ( .B1(n3651), .B2(n3653), .A(n3652), .ZN(n3737) );
  XNOR2_X1 U2873 ( .A(n2455), .B(n2456), .ZN(n3472) );
  NAND2_X1 U2874 ( .A1(n4897), .A2(n2867), .ZN(n3698) );
  NAND2_X1 U2875 ( .A1(n2338), .A2(n2869), .ZN(n3648) );
  INV_X1 U2876 ( .A(n3832), .ZN(n2288) );
  NAND2_X1 U2877 ( .A1(n4910), .A2(n4895), .ZN(n2214) );
  NAND2_X1 U2878 ( .A1(n2196), .A2(n2304), .ZN(n2658) );
  NOR3_X1 U2879 ( .A1(n3696), .A2(n2260), .A3(n4475), .ZN(n2259) );
  OR2_X1 U2880 ( .A1(n3696), .A2(n2260), .ZN(n2215) );
  AND2_X1 U2881 ( .A1(n2294), .A2(n2192), .ZN(n2216) );
  AND2_X2 U2882 ( .A1(n3252), .A2(n3251), .ZN(n4920) );
  NAND2_X1 U2883 ( .A1(n3374), .A2(n3373), .ZN(n3372) );
  OR2_X1 U2884 ( .A1(n4910), .A2(n2948), .ZN(n2217) );
  AND2_X1 U2885 ( .A1(n3443), .A2(n2851), .ZN(n2218) );
  INV_X1 U2886 ( .A(n4749), .ZN(n2270) );
  INV_X1 U2887 ( .A(IR_REG_29__SCAN_IN), .ZN(n2237) );
  INV_X1 U2888 ( .A(IR_REG_17__SCAN_IN), .ZN(n2345) );
  AND2_X1 U2889 ( .A1(n4714), .A2(REG1_REG_18__SCAN_IN), .ZN(n2219) );
  AND2_X1 U2890 ( .A1(n4714), .A2(REG2_REG_18__SCAN_IN), .ZN(n2220) );
  NAND4_X1 U2891 ( .A1(n2304), .A2(n2305), .A3(n2258), .A4(n2436), .ZN(n2257)
         );
  INV_X1 U2892 ( .A(n2304), .ZN(n2600) );
  AND2_X4 U2893 ( .A1(n2435), .A2(n2364), .ZN(n2436) );
  AND2_X2 U2894 ( .A1(n2226), .A2(n2225), .ZN(n2435) );
  INV_X1 U2895 ( .A(IR_REG_13__SCAN_IN), .ZN(n2603) );
  NAND2_X1 U2896 ( .A1(n4366), .A2(n2230), .ZN(n2229) );
  NAND2_X2 U2897 ( .A1(n2238), .A2(IR_REG_31__SCAN_IN), .ZN(n2373) );
  NAND3_X1 U2898 ( .A1(n2383), .A2(n2237), .A3(n2186), .ZN(n2238) );
  XNOR2_X1 U2899 ( .A(n2251), .B(n2250), .ZN(n4185) );
  XNOR2_X1 U2900 ( .A(n4146), .B(n4162), .ZN(n4805) );
  NAND2_X1 U2901 ( .A1(n4145), .A2(n4795), .ZN(n4146) );
  NOR2_X2 U2902 ( .A1(n2257), .A2(n2341), .ZN(n2383) );
  INV_X1 U2903 ( .A(n2259), .ZN(n4477) );
  NAND3_X1 U2904 ( .A1(n3556), .A2(n2265), .A3(n3671), .ZN(n3695) );
  MUX2_X1 U2905 ( .A(REG2_REG_2__SCAN_IN), .B(n3526), .S(n4719), .Z(n4118) );
  XNOR2_X1 U2906 ( .A(n2425), .B(n2426), .ZN(n3451) );
  NAND2_X1 U2907 ( .A1(n2276), .A2(n2274), .ZN(n3259) );
  NAND2_X1 U2908 ( .A1(n3803), .A2(n2281), .ZN(n2280) );
  NAND2_X1 U2909 ( .A1(n2548), .A2(n2188), .ZN(n3268) );
  NAND2_X1 U2910 ( .A1(n2294), .A2(n2198), .ZN(n2515) );
  NAND2_X1 U2911 ( .A1(n2299), .A2(n3901), .ZN(n2838) );
  NAND2_X1 U2912 ( .A1(n2299), .A2(n2297), .ZN(n2303) );
  OAI211_X1 U2913 ( .C1(n2213), .C2(n2303), .A(n2300), .B(n2837), .ZN(U3217)
         );
  NOR2_X1 U2914 ( .A1(n2355), .A2(n2302), .ZN(n2301) );
  NAND3_X1 U2915 ( .A1(n2304), .A2(n2305), .A3(n2436), .ZN(n2615) );
  NAND2_X1 U2916 ( .A1(n3792), .A2(n2212), .ZN(n2306) );
  NAND2_X1 U2917 ( .A1(n2306), .A2(n2307), .ZN(n3776) );
  NAND2_X2 U2918 ( .A1(n2315), .A2(n2314), .ZN(n2415) );
  NAND2_X1 U2919 ( .A1(n4433), .A2(n2323), .ZN(n2322) );
  NAND2_X1 U2920 ( .A1(n2322), .A2(n2324), .ZN(n4386) );
  OAI21_X1 U2921 ( .B1(n3753), .B2(n4589), .A(n2943), .ZN(n4508) );
  XNOR2_X1 U2922 ( .A(n2331), .B(n3232), .ZN(U3514) );
  NAND2_X2 U2923 ( .A1(n4003), .A2(n2903), .ZN(n2902) );
  NAND2_X2 U2924 ( .A1(n2850), .A2(n3456), .ZN(n2903) );
  AND4_X2 U2925 ( .A1(n2845), .A2(n2846), .A3(n2847), .A4(n2844), .ZN(n2850)
         );
  NAND2_X1 U2926 ( .A1(n2334), .A2(n2332), .ZN(n2895) );
  NAND2_X1 U2927 ( .A1(n2338), .A2(n2199), .ZN(n2871) );
  NAND2_X1 U2928 ( .A1(n2383), .A2(n2369), .ZN(n2387) );
  NOR2_X1 U2929 ( .A1(n2387), .A2(IR_REG_25__SCAN_IN), .ZN(n2381) );
  OAI21_X1 U2930 ( .B1(n3776), .B2(n2742), .A(n2741), .ZN(n3842) );
  AOI21_X2 U2931 ( .B1(n3786), .B2(n3785), .A(n2352), .ZN(n3792) );
  AOI21_X2 U2932 ( .B1(n2625), .B2(n2356), .A(n2624), .ZN(n2650) );
  AOI21_X1 U2933 ( .B1(n3235), .B2(n3964), .A(n3234), .ZN(n3236) );
  NAND2_X1 U2934 ( .A1(n3424), .A2(n4478), .ZN(n4724) );
  NAND2_X1 U2935 ( .A1(n2578), .A2(n2577), .ZN(n3803) );
  INV_X1 U2936 ( .A(n4583), .ZN(n4404) );
  AND2_X1 U2937 ( .A1(n2642), .A2(n2365), .ZN(n2351) );
  AND2_X1 U2938 ( .A1(n2686), .A2(n2685), .ZN(n2352) );
  AND2_X1 U2939 ( .A1(n2810), .A2(n2809), .ZN(n2353) );
  INV_X1 U2940 ( .A(n4580), .ZN(n3827) );
  NAND2_X1 U2941 ( .A1(n2856), .A2(n2855), .ZN(n3494) );
  AND4_X1 U2942 ( .A1(n2641), .A2(n2640), .A3(n2639), .A4(n2638), .ZN(n4575)
         );
  OR2_X1 U2943 ( .A1(n2675), .A2(n3889), .ZN(n2354) );
  INV_X1 U2944 ( .A(n4613), .ZN(n4475) );
  XOR2_X1 U2945 ( .A(n2807), .B(n2806), .Z(n2355) );
  NAND2_X1 U2946 ( .A1(n3929), .A2(DATAI_23_), .ZN(n4278) );
  INV_X1 U2947 ( .A(n2446), .ZN(n2409) );
  NAND2_X1 U2948 ( .A1(n2620), .A2(n2621), .ZN(n2356) );
  INV_X1 U2949 ( .A(n4357), .ZN(n2882) );
  INV_X1 U2950 ( .A(n4591), .ZN(n4422) );
  OAI22_X1 U2951 ( .A1(n3494), .A2(n2863), .B1(n2862), .B2(n2861), .ZN(n3616)
         );
  AND2_X1 U2952 ( .A1(n3794), .A2(n3793), .ZN(n2357) );
  OR2_X1 U2953 ( .A1(n4632), .A2(n4613), .ZN(n2358) );
  INV_X1 U2954 ( .A(n3851), .ZN(n2710) );
  NAND2_X1 U2955 ( .A1(n4086), .A2(n3710), .ZN(n2359) );
  AND2_X1 U2956 ( .A1(n4269), .A2(n4272), .ZN(n3948) );
  NAND2_X1 U2957 ( .A1(n2430), .A2(REG2_REG_1__SCAN_IN), .ZN(n2844) );
  INV_X1 U2958 ( .A(n2847), .ZN(n2848) );
  OR2_X1 U2959 ( .A1(n2425), .A2(n2427), .ZN(n2428) );
  AND2_X1 U2960 ( .A1(n3976), .A2(n4234), .ZN(n4062) );
  NAND2_X1 U2961 ( .A1(n4329), .A2(n4357), .ZN(n2884) );
  INV_X1 U2962 ( .A(n2755), .ZN(n2419) );
  OR2_X1 U2963 ( .A1(n2734), .A2(n3846), .ZN(n2744) );
  OR2_X1 U2964 ( .A1(n4520), .A2(n4209), .ZN(n3953) );
  NOR2_X1 U2965 ( .A1(n2886), .A2(n4275), .ZN(n4303) );
  NOR2_X1 U2966 ( .A1(n2687), .A2(n2361), .ZN(n2698) );
  NAND2_X1 U2967 ( .A1(n4613), .A2(n4632), .ZN(n2875) );
  INV_X1 U2968 ( .A(n3979), .ZN(n2873) );
  OR2_X1 U2969 ( .A1(n3495), .A2(n2861), .ZN(n2863) );
  INV_X1 U2970 ( .A(n4303), .ZN(n2887) );
  AND2_X1 U2971 ( .A1(n3416), .A2(n4713), .ZN(n4627) );
  INV_X1 U2972 ( .A(n2938), .ZN(n3299) );
  XNOR2_X1 U2973 ( .A(n2511), .B(n2512), .ZN(n3662) );
  AND2_X1 U2974 ( .A1(n2698), .A2(REG3_REG_21__SCAN_IN), .ZN(n2720) );
  INV_X1 U2975 ( .A(n4086), .ZN(n3721) );
  OAI21_X1 U2976 ( .B1(n3813), .B2(n3814), .A(n3815), .ZN(n3904) );
  AND2_X1 U2977 ( .A1(n2761), .A2(n2760), .ZN(n2762) );
  AND4_X1 U2978 ( .A1(n2632), .A2(n2631), .A3(n2630), .A4(n2629), .ZN(n4583)
         );
  INV_X1 U2979 ( .A(n4722), .ZN(n3402) );
  INV_X1 U2980 ( .A(REG3_REG_12__SCAN_IN), .ZN(n3809) );
  INV_X1 U2981 ( .A(n4709), .ZN(n4093) );
  INV_X1 U2982 ( .A(n4551), .ZN(n4318) );
  AND2_X1 U2983 ( .A1(n4022), .A2(n4032), .ZN(n3989) );
  INV_X1 U2984 ( .A(n3611), .ZN(n3506) );
  INV_X1 U2985 ( .A(n3348), .ZN(n4513) );
  INV_X1 U2986 ( .A(n4278), .ZN(n4283) );
  INV_X1 U2987 ( .A(n4390), .ZN(n4571) );
  INV_X1 U2988 ( .A(n4604), .ZN(n4461) );
  NAND2_X1 U2989 ( .A1(n3402), .A2(n3299), .ZN(n4615) );
  NOR2_X1 U2990 ( .A1(n2601), .A2(IR_REG_5__SCAN_IN), .ZN(n2509) );
  INV_X1 U2991 ( .A(n3718), .ZN(n3726) );
  OR2_X1 U2992 ( .A1(n2664), .A2(n3085), .ZN(n2687) );
  NAND2_X1 U2993 ( .A1(n2652), .A2(REG3_REG_17__SCAN_IN), .ZN(n2664) );
  OR2_X1 U2994 ( .A1(n2569), .A2(n2360), .ZN(n2579) );
  INV_X1 U2995 ( .A(n3898), .ZN(n3918) );
  NAND4_X1 U2996 ( .A1(n2703), .A2(n2702), .A3(n2701), .A4(n2700), .ZN(n4327)
         );
  AND4_X1 U2997 ( .A1(n2614), .A2(n2613), .A3(n2612), .A4(n2611), .ZN(n4605)
         );
  AND2_X1 U2998 ( .A1(n3338), .A2(n3337), .ZN(n4094) );
  NAND2_X1 U2999 ( .A1(n2937), .A2(n4075), .ZN(n4491) );
  INV_X1 U3000 ( .A(n4488), .ZN(n4828) );
  INV_X1 U3001 ( .A(n4483), .ZN(n4462) );
  OR2_X1 U3002 ( .A1(n4920), .A2(n3082), .ZN(n3253) );
  AOI21_X1 U3003 ( .B1(n2784), .B2(n3289), .A(n3288), .ZN(n3251) );
  NAND2_X1 U3004 ( .A1(n4333), .A2(n4884), .ZN(n4895) );
  INV_X1 U3005 ( .A(n2876), .ZN(n4443) );
  AND3_X1 U3006 ( .A1(n2947), .A2(n3420), .A3(n2946), .ZN(n3252) );
  AND2_X1 U3007 ( .A1(n2836), .A2(n2835), .ZN(n2837) );
  OR2_X1 U3008 ( .A1(n2830), .A2(n2792), .ZN(n3898) );
  INV_X1 U3009 ( .A(n4531), .ZN(n4218) );
  INV_X1 U3010 ( .A(n4575), .ZN(n4593) );
  INV_X1 U3011 ( .A(n4773), .ZN(n4809) );
  NAND2_X1 U3012 ( .A1(n4094), .A2(n4722), .ZN(n4822) );
  INV_X1 U3013 ( .A(n4724), .ZN(n4825) );
  INV_X1 U3014 ( .A(n4724), .ZN(n4493) );
  AND2_X1 U3015 ( .A1(n3254), .A2(n3253), .ZN(n3255) );
  NAND2_X1 U3016 ( .A1(n4920), .A2(n4585), .ZN(n4640) );
  AND2_X1 U3017 ( .A1(n3248), .A2(n3247), .ZN(n3249) );
  NAND2_X1 U3018 ( .A1(n4910), .A2(n4585), .ZN(n4706) );
  INV_X1 U3019 ( .A(n4847), .ZN(n4852) );
  NOR2_X1 U3020 ( .A1(n2417), .A2(n3257), .ZN(U4043) );
  OAI21_X1 U3021 ( .B1(n3256), .B2(n4918), .A(n3255), .ZN(U3547) );
  OAI21_X1 U3022 ( .B1(n3256), .B2(n3250), .A(n3249), .ZN(U3515) );
  INV_X2 U3023 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  NAND2_X1 U3024 ( .A1(n2490), .A2(REG3_REG_6__SCAN_IN), .ZN(n2502) );
  NOR2_X1 U3025 ( .A1(n2502), .A2(n3387), .ZN(n2517) );
  NAND2_X1 U3026 ( .A1(n2517), .A2(REG3_REG_8__SCAN_IN), .ZN(n2533) );
  NAND2_X1 U3027 ( .A1(REG3_REG_10__SCAN_IN), .A2(REG3_REG_11__SCAN_IN), .ZN(
        n2360) );
  NAND2_X1 U3028 ( .A1(n2594), .A2(REG3_REG_13__SCAN_IN), .ZN(n2609) );
  NAND2_X1 U3029 ( .A1(REG3_REG_19__SCAN_IN), .A2(REG3_REG_20__SCAN_IN), .ZN(
        n2361) );
  AND2_X1 U3030 ( .A1(REG3_REG_22__SCAN_IN), .A2(REG3_REG_23__SCAN_IN), .ZN(
        n2362) );
  NAND2_X1 U3031 ( .A1(n2720), .A2(n2362), .ZN(n2734) );
  INV_X1 U3032 ( .A(REG3_REG_24__SCAN_IN), .ZN(n3846) );
  INV_X1 U3033 ( .A(REG3_REG_25__SCAN_IN), .ZN(n3818) );
  NAND2_X1 U3034 ( .A1(n2758), .A2(REG3_REG_26__SCAN_IN), .ZN(n2793) );
  XNOR2_X1 U3035 ( .A(n2793), .B(REG3_REG_27__SCAN_IN), .ZN(n4207) );
  NAND2_X1 U3036 ( .A1(n2370), .A2(IR_REG_31__SCAN_IN), .ZN(n2371) );
  NAND2_X1 U3037 ( .A1(n4207), .A2(n2409), .ZN(n2380) );
  INV_X1 U3038 ( .A(REG1_REG_27__SCAN_IN), .ZN(n4516) );
  XNOR2_X2 U3039 ( .A(n2373), .B(n2372), .ZN(n2375) );
  NAND2_X1 U3040 ( .A1(n2375), .A2(n4708), .ZN(n2549) );
  NAND2_X1 U3041 ( .A1(n3302), .A2(REG2_REG_27__SCAN_IN), .ZN(n2377) );
  INV_X1 U3042 ( .A(n4708), .ZN(n2374) );
  AND2_X4 U3043 ( .A1(n2375), .A2(n2374), .ZN(n2429) );
  NAND2_X1 U3044 ( .A1(n2429), .A2(REG0_REG_27__SCAN_IN), .ZN(n2376) );
  OAI211_X1 U3045 ( .C1(n4516), .C2(n3305), .A(n2377), .B(n2376), .ZN(n2378)
         );
  INV_X1 U3046 ( .A(n2378), .ZN(n2379) );
  INV_X1 U3047 ( .A(n2381), .ZN(n2389) );
  NAND2_X1 U3048 ( .A1(n2389), .A2(IR_REG_31__SCAN_IN), .ZN(n2382) );
  XNOR2_X2 U3049 ( .A(n2382), .B(IR_REG_26__SCAN_IN), .ZN(n4710) );
  NAND2_X1 U3050 ( .A1(n2788), .A2(n2787), .ZN(n2384) );
  INV_X1 U3051 ( .A(n2774), .ZN(n4711) );
  NAND2_X1 U3052 ( .A1(n2387), .A2(IR_REG_31__SCAN_IN), .ZN(n2388) );
  MUX2_X1 U3053 ( .A(IR_REG_31__SCAN_IN), .B(n2388), .S(IR_REG_25__SCAN_IN), 
        .Z(n2390) );
  NAND2_X1 U3054 ( .A1(n2390), .A2(n2389), .ZN(n2773) );
  INV_X1 U3055 ( .A(n2773), .ZN(n3281) );
  NAND2_X1 U3056 ( .A1(n2391), .A2(IR_REG_31__SCAN_IN), .ZN(n2402) );
  NAND2_X1 U3057 ( .A1(n2402), .A2(n2401), .ZN(n2392) );
  NAND2_X1 U3058 ( .A1(n2392), .A2(IR_REG_31__SCAN_IN), .ZN(n2393) );
  NAND2_X1 U3059 ( .A1(n2187), .A2(IR_REG_31__SCAN_IN), .ZN(n2394) );
  INV_X1 U3060 ( .A(n3425), .ZN(n2395) );
  NAND2_X2 U3061 ( .A1(n2417), .A2(n2395), .ZN(n2672) );
  INV_X2 U3062 ( .A(n2672), .ZN(n2798) );
  NAND2_X1 U3063 ( .A1(n4520), .A2(n2798), .ZN(n2399) );
  NAND2_X1 U3064 ( .A1(n3243), .A2(n2824), .ZN(n2397) );
  NAND2_X1 U3065 ( .A1(n4509), .A2(n2799), .ZN(n2398) );
  NAND2_X1 U3066 ( .A1(n2399), .A2(n2398), .ZN(n2403) );
  NAND2_X1 U3067 ( .A1(n2197), .A2(IR_REG_31__SCAN_IN), .ZN(n2400) );
  NAND2_X1 U3068 ( .A1(n4712), .A2(n4179), .ZN(n2815) );
  XNOR2_X1 U3069 ( .A(n2403), .B(n2753), .ZN(n2810) );
  INV_X1 U3070 ( .A(n4712), .ZN(n2404) );
  INV_X1 U3071 ( .A(n4005), .ZN(n3974) );
  NOR2_X1 U3072 ( .A1(n4209), .A2(n2767), .ZN(n2407) );
  AOI21_X1 U3073 ( .B1(n4520), .B2(n2804), .A(n2407), .ZN(n2808) );
  NAND2_X1 U3074 ( .A1(n2429), .A2(REG0_REG_1__SCAN_IN), .ZN(n2845) );
  INV_X1 U3075 ( .A(n2549), .ZN(n2408) );
  INV_X1 U3076 ( .A(REG1_REG_1__SCAN_IN), .ZN(n3340) );
  NAND2_X1 U3077 ( .A1(n2408), .A2(REG1_REG_1__SCAN_IN), .ZN(n2846) );
  INV_X1 U3078 ( .A(REG3_REG_1__SCAN_IN), .ZN(n3512) );
  NAND2_X1 U3079 ( .A1(n2409), .A2(REG3_REG_1__SCAN_IN), .ZN(n2847) );
  INV_X1 U3080 ( .A(n2672), .ZN(n2818) );
  NAND2_X1 U3081 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n2410)
         );
  MUX2_X1 U3082 ( .A(n4720), .B(DATAI_1_), .S(n2415), .Z(n3456) );
  NAND2_X1 U3083 ( .A1(n2408), .A2(REG1_REG_0__SCAN_IN), .ZN(n2414) );
  INV_X1 U3084 ( .A(REG3_REG_0__SCAN_IN), .ZN(n3427) );
  OR2_X1 U3085 ( .A1(n2446), .A2(n3427), .ZN(n2413) );
  NAND2_X1 U3086 ( .A1(n2429), .A2(REG0_REG_0__SCAN_IN), .ZN(n2412) );
  NAND2_X1 U3087 ( .A1(n2430), .A2(REG2_REG_0__SCAN_IN), .ZN(n2411) );
  MUX2_X1 U3088 ( .A(IR_REG_0__SCAN_IN), .B(DATAI_0_), .S(n2415), .Z(n3376) );
  AND2_X1 U3089 ( .A1(n3376), .A2(n2406), .ZN(n2416) );
  INV_X1 U3090 ( .A(n2417), .ZN(n2420) );
  NAND2_X1 U3091 ( .A1(n2420), .A2(REG1_REG_0__SCAN_IN), .ZN(n2418) );
  NAND2_X1 U3092 ( .A1(n2423), .A2(n2418), .ZN(n3374) );
  NAND2_X1 U3093 ( .A1(n4091), .A2(n2419), .ZN(n2422) );
  AOI22_X1 U3094 ( .A1(n3376), .A2(n2798), .B1(IR_REG_0__SCAN_IN), .B2(n2420), 
        .ZN(n2421) );
  NAND2_X1 U3095 ( .A1(n2422), .A2(n2421), .ZN(n3373) );
  NAND2_X1 U3096 ( .A1(n2423), .A2(n2802), .ZN(n2424) );
  NAND2_X1 U3097 ( .A1(n3372), .A2(n2424), .ZN(n3452) );
  NAND2_X1 U3098 ( .A1(n3451), .A2(n3452), .ZN(n3453) );
  INV_X1 U3099 ( .A(n2426), .ZN(n2427) );
  NAND2_X1 U3100 ( .A1(n3453), .A2(n2428), .ZN(n3460) );
  INV_X1 U3101 ( .A(n3460), .ZN(n2440) );
  NAND2_X1 U3102 ( .A1(n2408), .A2(REG1_REG_2__SCAN_IN), .ZN(n2434) );
  NAND2_X1 U3103 ( .A1(n2429), .A2(REG0_REG_2__SCAN_IN), .ZN(n2433) );
  INV_X1 U3104 ( .A(REG3_REG_2__SCAN_IN), .ZN(n4111) );
  OR2_X1 U3105 ( .A1(n2446), .A2(n4111), .ZN(n2432) );
  NAND2_X1 U3106 ( .A1(n2430), .A2(REG2_REG_2__SCAN_IN), .ZN(n2431) );
  OAI22_X1 U3107 ( .A1(n2852), .A2(n2755), .B1(n4877), .B2(n2767), .ZN(n2442)
         );
  NAND2_X1 U3108 ( .A1(n2440), .A2(n2439), .ZN(n3461) );
  INV_X1 U3109 ( .A(n2441), .ZN(n2444) );
  INV_X1 U3110 ( .A(n2442), .ZN(n2443) );
  NAND2_X1 U3111 ( .A1(n2444), .A2(n2443), .ZN(n2445) );
  NAND2_X1 U3112 ( .A1(n3461), .A2(n2445), .ZN(n3473) );
  OR2_X1 U3113 ( .A1(n2446), .A2(REG3_REG_3__SCAN_IN), .ZN(n2451) );
  INV_X1 U3114 ( .A(REG1_REG_3__SCAN_IN), .ZN(n2447) );
  OR2_X1 U3115 ( .A1(n2549), .A2(n2447), .ZN(n2450) );
  NAND2_X1 U3116 ( .A1(n2429), .A2(REG0_REG_3__SCAN_IN), .ZN(n2449) );
  NAND2_X1 U3117 ( .A1(n2430), .A2(REG2_REG_3__SCAN_IN), .ZN(n2448) );
  NAND2_X1 U3118 ( .A1(n3551), .A2(n2798), .ZN(n2453) );
  OR2_X1 U3119 ( .A1(n2436), .A2(n3293), .ZN(n2465) );
  XNOR2_X1 U3120 ( .A(n2465), .B(IR_REG_3__SCAN_IN), .ZN(n4718) );
  MUX2_X1 U3121 ( .A(n4718), .B(DATAI_3_), .S(n2415), .Z(n3542) );
  NAND2_X1 U3122 ( .A1(n3542), .A2(n2799), .ZN(n2452) );
  AOI22_X1 U3123 ( .A1(n3551), .A2(n2804), .B1(n2798), .B2(n3542), .ZN(n2456)
         );
  INV_X1 U3124 ( .A(n2455), .ZN(n2457) );
  NAND2_X1 U3125 ( .A1(n2457), .A2(n2456), .ZN(n2458) );
  NAND2_X1 U3126 ( .A1(n2430), .A2(REG2_REG_4__SCAN_IN), .ZN(n2463) );
  NAND2_X1 U3127 ( .A1(n2429), .A2(REG0_REG_4__SCAN_IN), .ZN(n2462) );
  XNOR2_X1 U3128 ( .A(REG3_REG_4__SCAN_IN), .B(REG3_REG_3__SCAN_IN), .ZN(n3557) );
  OR2_X1 U3129 ( .A1(n2822), .A2(n3557), .ZN(n2461) );
  INV_X1 U3130 ( .A(REG1_REG_4__SCAN_IN), .ZN(n2459) );
  OR2_X1 U3131 ( .A1(n2549), .A2(n2459), .ZN(n2460) );
  NAND2_X1 U3132 ( .A1(n2465), .A2(n2464), .ZN(n2466) );
  NAND2_X1 U3133 ( .A1(n2466), .A2(IR_REG_31__SCAN_IN), .ZN(n2467) );
  XNOR2_X1 U3134 ( .A(n2467), .B(IR_REG_4__SCAN_IN), .ZN(n4717) );
  MUX2_X1 U3135 ( .A(n4717), .B(DATAI_4_), .S(n2415), .Z(n2858) );
  OAI22_X1 U3136 ( .A1(n2857), .A2(n2752), .B1(n2751), .B2(n3555), .ZN(n2468)
         );
  XNOR2_X1 U3137 ( .A(n2468), .B(n2753), .ZN(n2470) );
  OAI22_X1 U3138 ( .A1(n2857), .A2(n2755), .B1(n2767), .B2(n3555), .ZN(n2469)
         );
  XNOR2_X1 U3139 ( .A(n2470), .B(n2469), .ZN(n3261) );
  NAND2_X1 U3140 ( .A1(n2470), .A2(n2469), .ZN(n2471) );
  NAND2_X1 U3141 ( .A1(n3259), .A2(n2471), .ZN(n3610) );
  NAND2_X1 U3142 ( .A1(n2429), .A2(REG0_REG_5__SCAN_IN), .ZN(n2479) );
  NAND2_X1 U3143 ( .A1(n2430), .A2(REG2_REG_5__SCAN_IN), .ZN(n2478) );
  INV_X1 U3144 ( .A(REG1_REG_5__SCAN_IN), .ZN(n3366) );
  OR2_X1 U3145 ( .A1(n3305), .A2(n3366), .ZN(n2477) );
  INV_X1 U3146 ( .A(n2490), .ZN(n2475) );
  INV_X1 U3147 ( .A(REG3_REG_5__SCAN_IN), .ZN(n2473) );
  NAND2_X1 U31480 ( .A1(REG3_REG_4__SCAN_IN), .A2(REG3_REG_3__SCAN_IN), .ZN(
        n2472) );
  NAND2_X1 U31490 ( .A1(n2473), .A2(n2472), .ZN(n2474) );
  NAND2_X1 U3150 ( .A1(n2475), .A2(n2474), .ZN(n3615) );
  OR2_X1 U3151 ( .A1(n2822), .A2(n3615), .ZN(n2476) );
  NAND2_X1 U3152 ( .A1(n2481), .A2(n2480), .ZN(n2601) );
  NAND2_X1 U3153 ( .A1(n2601), .A2(IR_REG_31__SCAN_IN), .ZN(n2483) );
  INV_X1 U3154 ( .A(IR_REG_5__SCAN_IN), .ZN(n2482) );
  XNOR2_X1 U3155 ( .A(n2483), .B(n2482), .ZN(n4131) );
  INV_X1 U3156 ( .A(DATAI_5_), .ZN(n2484) );
  MUX2_X1 U3157 ( .A(n4131), .B(n2484), .S(n2415), .Z(n3611) );
  OAI22_X1 U3158 ( .A1(n2859), .A2(n2752), .B1(n2751), .B2(n3611), .ZN(n2485)
         );
  XNOR2_X1 U3159 ( .A(n2485), .B(n2802), .ZN(n2486) );
  OAI22_X1 U3160 ( .A1(n2859), .A2(n2755), .B1(n2767), .B2(n3611), .ZN(n2487)
         );
  XNOR2_X1 U3161 ( .A(n2486), .B(n2487), .ZN(n3609) );
  NAND2_X1 U3162 ( .A1(n3610), .A2(n3609), .ZN(n3608) );
  INV_X1 U3163 ( .A(n2486), .ZN(n2488) );
  NAND2_X1 U3164 ( .A1(n2488), .A2(n2487), .ZN(n2489) );
  OAI21_X1 U3165 ( .B1(n2490), .B2(REG3_REG_6__SCAN_IN), .A(n2502), .ZN(n3755)
         );
  OR2_X1 U3166 ( .A1(n2822), .A2(n3755), .ZN(n2495) );
  INV_X1 U3167 ( .A(REG1_REG_6__SCAN_IN), .ZN(n2491) );
  OR2_X1 U3168 ( .A1(n3305), .A2(n2491), .ZN(n2494) );
  NAND2_X1 U3169 ( .A1(n3302), .A2(REG2_REG_6__SCAN_IN), .ZN(n2493) );
  NAND2_X1 U3170 ( .A1(n2429), .A2(REG0_REG_6__SCAN_IN), .ZN(n2492) );
  NAND4_X1 U3171 ( .A1(n2495), .A2(n2494), .A3(n2493), .A4(n2492), .ZN(n3676)
         );
  NAND2_X1 U3172 ( .A1(n3676), .A2(n2804), .ZN(n2498) );
  OR2_X1 U3173 ( .A1(n2509), .A2(n3293), .ZN(n2496) );
  XNOR2_X1 U3174 ( .A(n2496), .B(IR_REG_6__SCAN_IN), .ZN(n4716) );
  MUX2_X1 U3175 ( .A(n4716), .B(DATAI_6_), .S(n3929), .Z(n3621) );
  NAND2_X1 U3176 ( .A1(n3621), .A2(n2798), .ZN(n2497) );
  NAND2_X1 U3177 ( .A1(n2498), .A2(n2497), .ZN(n3630) );
  NAND2_X1 U3178 ( .A1(n3676), .A2(n2798), .ZN(n2500) );
  NAND2_X1 U3179 ( .A1(n3621), .A2(n2799), .ZN(n2499) );
  NAND2_X1 U3180 ( .A1(n2500), .A2(n2499), .ZN(n2501) );
  XNOR2_X1 U3181 ( .A(n2501), .B(n2753), .ZN(n3631) );
  NAND2_X1 U3182 ( .A1(n3302), .A2(REG2_REG_7__SCAN_IN), .ZN(n2507) );
  NAND2_X1 U3183 ( .A1(n2429), .A2(REG0_REG_7__SCAN_IN), .ZN(n2506) );
  AND2_X1 U3184 ( .A1(n2502), .A2(n3387), .ZN(n2503) );
  OR2_X1 U3185 ( .A1(n2503), .A2(n2517), .ZN(n3678) );
  OR2_X1 U3186 ( .A1(n2822), .A2(n3678), .ZN(n2505) );
  INV_X1 U3187 ( .A(REG1_REG_7__SCAN_IN), .ZN(n3385) );
  OR2_X1 U3188 ( .A1(n3305), .A2(n3385), .ZN(n2504) );
  NAND2_X1 U3189 ( .A1(n2509), .A2(n2508), .ZN(n2539) );
  NAND2_X1 U3190 ( .A1(n2539), .A2(IR_REG_31__SCAN_IN), .ZN(n2524) );
  XNOR2_X1 U3191 ( .A(n2524), .B(IR_REG_7__SCAN_IN), .ZN(n4715) );
  MUX2_X1 U3192 ( .A(n4715), .B(DATAI_7_), .S(n3929), .Z(n2866) );
  OAI22_X1 U3193 ( .A1(n3657), .A2(n2752), .B1(n2751), .B2(n3671), .ZN(n2510)
         );
  XNOR2_X1 U3194 ( .A(n2510), .B(n2802), .ZN(n2511) );
  OAI22_X1 U3195 ( .A1(n3657), .A2(n2755), .B1(n2767), .B2(n3671), .ZN(n2512)
         );
  INV_X1 U3196 ( .A(n2511), .ZN(n2513) );
  NAND2_X1 U3197 ( .A1(n2513), .A2(n2512), .ZN(n2514) );
  NAND2_X1 U3198 ( .A1(n2515), .A2(n2514), .ZN(n3651) );
  NAND2_X1 U3199 ( .A1(n2429), .A2(REG0_REG_8__SCAN_IN), .ZN(n2522) );
  NAND2_X1 U3200 ( .A1(n3302), .A2(REG2_REG_8__SCAN_IN), .ZN(n2521) );
  INV_X1 U3201 ( .A(REG1_REG_8__SCAN_IN), .ZN(n2516) );
  OR2_X1 U3202 ( .A1(n3305), .A2(n2516), .ZN(n2520) );
  OR2_X1 U3203 ( .A1(n2517), .A2(REG3_REG_8__SCAN_IN), .ZN(n2518) );
  NAND2_X1 U3204 ( .A1(n2533), .A2(n2518), .ZN(n3656) );
  OR2_X1 U3205 ( .A1(n2822), .A2(n3656), .ZN(n2519) );
  INV_X1 U3206 ( .A(IR_REG_7__SCAN_IN), .ZN(n2523) );
  NAND2_X1 U3207 ( .A1(n2524), .A2(n2523), .ZN(n2525) );
  NAND2_X1 U3208 ( .A1(n2525), .A2(IR_REG_31__SCAN_IN), .ZN(n2526) );
  XNOR2_X1 U3209 ( .A(n2526), .B(IR_REG_8__SCAN_IN), .ZN(n3581) );
  INV_X1 U32100 ( .A(n3581), .ZN(n4870) );
  INV_X1 U32110 ( .A(DATAI_8_), .ZN(n4869) );
  MUX2_X1 U32120 ( .A(n4870), .B(n4869), .S(n3929), .Z(n3700) );
  OAI22_X1 U32130 ( .A1(n3741), .A2(n2672), .B1(n2751), .B2(n3700), .ZN(n2527)
         );
  XNOR2_X1 U32140 ( .A(n2527), .B(n2753), .ZN(n2528) );
  OAI22_X1 U32150 ( .A1(n3741), .A2(n2755), .B1(n2767), .B2(n3700), .ZN(n2529)
         );
  AND2_X1 U32160 ( .A1(n2528), .A2(n2529), .ZN(n3653) );
  INV_X1 U32170 ( .A(n2528), .ZN(n2531) );
  INV_X1 U32180 ( .A(n2529), .ZN(n2530) );
  NAND2_X1 U32190 ( .A1(n2531), .A2(n2530), .ZN(n3652) );
  NAND2_X1 U32200 ( .A1(n2533), .A2(n2532), .ZN(n2534) );
  NAND2_X1 U32210 ( .A1(n2569), .A2(n2534), .ZN(n3745) );
  OR2_X1 U32220 ( .A1(n2822), .A2(n3745), .ZN(n2538) );
  INV_X1 U32230 ( .A(REG1_REG_9__SCAN_IN), .ZN(n3734) );
  OR2_X1 U32240 ( .A1(n3305), .A2(n3734), .ZN(n2537) );
  NAND2_X1 U32250 ( .A1(n2429), .A2(REG0_REG_9__SCAN_IN), .ZN(n2536) );
  NAND2_X1 U32260 ( .A1(n3302), .A2(REG2_REG_9__SCAN_IN), .ZN(n2535) );
  NAND4_X1 U32270 ( .A1(n2538), .A2(n2537), .A3(n2536), .A4(n2535), .ZN(n4086)
         );
  NAND2_X1 U32280 ( .A1(n4086), .A2(n2798), .ZN(n2542) );
  NAND2_X1 U32290 ( .A1(n2555), .A2(IR_REG_31__SCAN_IN), .ZN(n2540) );
  XNOR2_X1 U32300 ( .A(n2540), .B(IR_REG_9__SCAN_IN), .ZN(n3578) );
  MUX2_X1 U32310 ( .A(n3578), .B(DATAI_9_), .S(n3929), .Z(n3710) );
  NAND2_X1 U32320 ( .A1(n3710), .A2(n2799), .ZN(n2541) );
  NAND2_X1 U32330 ( .A1(n2542), .A2(n2541), .ZN(n2543) );
  XNOR2_X1 U32340 ( .A(n2543), .B(n2753), .ZN(n2544) );
  AOI22_X1 U32350 ( .A1(n4086), .A2(n2804), .B1(n2798), .B2(n3710), .ZN(n2545)
         );
  XNOR2_X1 U32360 ( .A(n2544), .B(n2545), .ZN(n3738) );
  NAND2_X1 U32370 ( .A1(n3737), .A2(n3738), .ZN(n2548) );
  INV_X1 U32380 ( .A(n2544), .ZN(n2546) );
  NAND2_X1 U32390 ( .A1(n2546), .A2(n2545), .ZN(n2547) );
  INV_X1 U32400 ( .A(REG1_REG_10__SCAN_IN), .ZN(n2550) );
  OR2_X1 U32410 ( .A1(n3305), .A2(n2550), .ZN(n2554) );
  INV_X1 U32420 ( .A(REG3_REG_10__SCAN_IN), .ZN(n2568) );
  XNOR2_X1 U32430 ( .A(n2569), .B(n2568), .ZN(n3728) );
  OR2_X1 U32440 ( .A1(n2822), .A2(n3728), .ZN(n2553) );
  NAND2_X1 U32450 ( .A1(n2429), .A2(REG0_REG_10__SCAN_IN), .ZN(n2552) );
  NAND2_X1 U32460 ( .A1(n3302), .A2(REG2_REG_10__SCAN_IN), .ZN(n2551) );
  NAND4_X1 U32470 ( .A1(n2554), .A2(n2553), .A3(n2552), .A4(n2551), .ZN(n4629)
         );
  NAND2_X1 U32480 ( .A1(n4629), .A2(n2818), .ZN(n2558) );
  NAND2_X1 U32490 ( .A1(n2575), .A2(IR_REG_31__SCAN_IN), .ZN(n2556) );
  XNOR2_X1 U32500 ( .A(n2556), .B(IR_REG_10__SCAN_IN), .ZN(n4749) );
  MUX2_X1 U32510 ( .A(n4749), .B(DATAI_10_), .S(n3929), .Z(n3718) );
  NAND2_X1 U32520 ( .A1(n3718), .A2(n2799), .ZN(n2557) );
  NAND2_X1 U32530 ( .A1(n2558), .A2(n2557), .ZN(n2559) );
  XNOR2_X1 U32540 ( .A(n2559), .B(n2802), .ZN(n2561) );
  AOI22_X1 U32550 ( .A1(n4629), .A2(n2804), .B1(n2798), .B2(n3718), .ZN(n2562)
         );
  XNOR2_X1 U32560 ( .A(n2561), .B(n2562), .ZN(n3270) );
  INV_X1 U32570 ( .A(n3270), .ZN(n2560) );
  INV_X1 U32580 ( .A(n2561), .ZN(n2564) );
  INV_X1 U32590 ( .A(n2562), .ZN(n2563) );
  NAND2_X1 U32600 ( .A1(n2564), .A2(n2563), .ZN(n2565) );
  NAND2_X1 U32610 ( .A1(n2429), .A2(REG0_REG_11__SCAN_IN), .ZN(n2574) );
  NAND2_X1 U32620 ( .A1(n3302), .A2(REG2_REG_11__SCAN_IN), .ZN(n2573) );
  INV_X1 U32630 ( .A(REG1_REG_11__SCAN_IN), .ZN(n2566) );
  OR2_X1 U32640 ( .A1(n3305), .A2(n2566), .ZN(n2572) );
  INV_X1 U32650 ( .A(REG3_REG_11__SCAN_IN), .ZN(n2567) );
  OAI21_X1 U32660 ( .B1(n2569), .B2(n2568), .A(n2567), .ZN(n2570) );
  NAND2_X1 U32670 ( .A1(n2570), .A2(n2579), .ZN(n3888) );
  OR2_X1 U32680 ( .A1(n2822), .A2(n3888), .ZN(n2571) );
  XNOR2_X1 U32690 ( .A(n2586), .B(IR_REG_11__SCAN_IN), .ZN(n3577) );
  MUX2_X1 U32700 ( .A(n3577), .B(DATAI_11_), .S(n3929), .Z(n4628) );
  OAI22_X1 U32710 ( .A1(n4616), .A2(n2755), .B1(n2767), .B2(n3883), .ZN(n3879)
         );
  OAI22_X1 U32720 ( .A1(n4616), .A2(n2672), .B1(n2751), .B2(n3883), .ZN(n2576)
         );
  XNOR2_X1 U32730 ( .A(n2576), .B(n2753), .ZN(n3880) );
  NAND2_X1 U32740 ( .A1(n3878), .A2(n3879), .ZN(n2577) );
  NAND2_X1 U32750 ( .A1(n3302), .A2(REG2_REG_12__SCAN_IN), .ZN(n2584) );
  NAND2_X1 U32760 ( .A1(n2429), .A2(REG0_REG_12__SCAN_IN), .ZN(n2583) );
  AND2_X1 U32770 ( .A1(n2579), .A2(n3809), .ZN(n2580) );
  OR2_X1 U32780 ( .A1(n2580), .A2(n2594), .ZN(n4479) );
  OR2_X1 U32790 ( .A1(n2822), .A2(n4479), .ZN(n2582) );
  INV_X1 U32800 ( .A(REG1_REG_12__SCAN_IN), .ZN(n3084) );
  OR2_X1 U32810 ( .A1(n3305), .A2(n3084), .ZN(n2581) );
  INV_X1 U32820 ( .A(IR_REG_11__SCAN_IN), .ZN(n2585) );
  NAND2_X1 U32830 ( .A1(n2586), .A2(n2585), .ZN(n2587) );
  NAND2_X1 U32840 ( .A1(n2587), .A2(IR_REG_31__SCAN_IN), .ZN(n2588) );
  XNOR2_X1 U32850 ( .A(n2588), .B(IR_REG_12__SCAN_IN), .ZN(n3586) );
  INV_X1 U32860 ( .A(n3586), .ZN(n4863) );
  INV_X1 U32870 ( .A(DATAI_12_), .ZN(n4862) );
  MUX2_X1 U32880 ( .A(n4863), .B(n4862), .S(n3929), .Z(n4613) );
  OAI22_X1 U32890 ( .A1(n4632), .A2(n2672), .B1(n2751), .B2(n4613), .ZN(n2589)
         );
  XNOR2_X1 U32900 ( .A(n2589), .B(n2753), .ZN(n2590) );
  OAI22_X1 U32910 ( .A1(n4632), .A2(n2755), .B1(n2767), .B2(n4613), .ZN(n2591)
         );
  AND2_X1 U32920 ( .A1(n2590), .A2(n2591), .ZN(n3804) );
  INV_X1 U32930 ( .A(n2590), .ZN(n2593) );
  INV_X1 U32940 ( .A(n2591), .ZN(n2592) );
  NAND2_X1 U32950 ( .A1(n2593), .A2(n2592), .ZN(n3805) );
  NAND2_X1 U32960 ( .A1(n2429), .A2(REG0_REG_13__SCAN_IN), .ZN(n2599) );
  NAND2_X1 U32970 ( .A1(n3302), .A2(REG2_REG_13__SCAN_IN), .ZN(n2598) );
  OR2_X1 U32980 ( .A1(n3305), .A2(n4142), .ZN(n2597) );
  OR2_X1 U32990 ( .A1(n2594), .A2(REG3_REG_13__SCAN_IN), .ZN(n2595) );
  NAND2_X1 U33000 ( .A1(n2609), .A2(n2595), .ZN(n4464) );
  OR2_X1 U33010 ( .A1(n2822), .A2(n4464), .ZN(n2596) );
  NOR2_X1 U33020 ( .A1(n2601), .A2(n2600), .ZN(n2604) );
  OR2_X1 U33030 ( .A1(n2604), .A2(n3293), .ZN(n2602) );
  MUX2_X1 U33040 ( .A(n2602), .B(IR_REG_31__SCAN_IN), .S(n2603), .Z(n2605) );
  NAND2_X1 U33050 ( .A1(n2604), .A2(n2603), .ZN(n2616) );
  NAND2_X1 U33060 ( .A1(n2605), .A2(n2616), .ZN(n4141) );
  INV_X1 U33070 ( .A(DATAI_13_), .ZN(n2606) );
  MUX2_X1 U33080 ( .A(n4141), .B(n2606), .S(n3929), .Z(n4604) );
  OAI22_X1 U33090 ( .A1(n4614), .A2(n2672), .B1(n2751), .B2(n4604), .ZN(n2607)
         );
  XNOR2_X1 U33100 ( .A(n2607), .B(n2802), .ZN(n3861) );
  INV_X1 U33110 ( .A(n3768), .ZN(n2625) );
  NAND2_X1 U33120 ( .A1(n3302), .A2(REG2_REG_14__SCAN_IN), .ZN(n2614) );
  NAND2_X1 U33130 ( .A1(n2429), .A2(REG0_REG_14__SCAN_IN), .ZN(n2613) );
  NAND2_X1 U33140 ( .A1(n2609), .A2(n2608), .ZN(n2610) );
  NAND2_X1 U33150 ( .A1(n2627), .A2(n2610), .ZN(n4444) );
  OR2_X1 U33160 ( .A1(n2822), .A2(n4444), .ZN(n2612) );
  INV_X1 U33170 ( .A(REG1_REG_14__SCAN_IN), .ZN(n4602) );
  OR2_X1 U33180 ( .A1(n3305), .A2(n4602), .ZN(n2611) );
  NAND2_X1 U33190 ( .A1(n2616), .A2(IR_REG_31__SCAN_IN), .ZN(n2617) );
  MUX2_X1 U33200 ( .A(IR_REG_31__SCAN_IN), .B(n2617), .S(IR_REG_14__SCAN_IN), 
        .Z(n2618) );
  AND2_X1 U33210 ( .A1(n2615), .A2(n2618), .ZN(n4154) );
  MUX2_X1 U33220 ( .A(n4154), .B(DATAI_14_), .S(n3929), .Z(n2876) );
  OAI22_X1 U33230 ( .A1(n4605), .A2(n2672), .B1(n4443), .B2(n2751), .ZN(n2619)
         );
  XNOR2_X1 U33240 ( .A(n2619), .B(n2753), .ZN(n2620) );
  OAI22_X1 U33250 ( .A1(n4605), .A2(n2755), .B1(n4443), .B2(n2767), .ZN(n2621)
         );
  INV_X1 U33260 ( .A(n2620), .ZN(n2623) );
  INV_X1 U33270 ( .A(n2621), .ZN(n2622) );
  NAND2_X1 U33280 ( .A1(n2623), .A2(n2622), .ZN(n3769) );
  NAND2_X1 U33290 ( .A1(n3302), .A2(REG2_REG_15__SCAN_IN), .ZN(n2632) );
  NAND2_X1 U33300 ( .A1(n2429), .A2(REG0_REG_15__SCAN_IN), .ZN(n2631) );
  AND2_X1 U33310 ( .A1(n2627), .A2(n2626), .ZN(n2628) );
  OR2_X1 U33320 ( .A1(n2628), .A2(n2635), .ZN(n4424) );
  OR2_X1 U33330 ( .A1(n2822), .A2(n4424), .ZN(n2630) );
  INV_X1 U33340 ( .A(REG1_REG_15__SCAN_IN), .ZN(n4598) );
  OR2_X1 U33350 ( .A1(n3305), .A2(n4598), .ZN(n2629) );
  NAND2_X1 U33360 ( .A1(n2615), .A2(IR_REG_31__SCAN_IN), .ZN(n2643) );
  XNOR2_X1 U33370 ( .A(n2643), .B(IR_REG_15__SCAN_IN), .ZN(n4161) );
  MUX2_X1 U33380 ( .A(n4161), .B(DATAI_15_), .S(n3929), .Z(n4591) );
  OAI22_X1 U33390 ( .A1(n4583), .A2(n2672), .B1(n2751), .B2(n4422), .ZN(n2633)
         );
  XNOR2_X1 U33400 ( .A(n2633), .B(n2753), .ZN(n2649) );
  OAI22_X1 U33410 ( .A1(n4583), .A2(n2755), .B1(n2752), .B2(n4422), .ZN(n2634)
         );
  INV_X1 U33420 ( .A(n2634), .ZN(n3916) );
  NAND2_X1 U33430 ( .A1(n3302), .A2(REG2_REG_16__SCAN_IN), .ZN(n2641) );
  NAND2_X1 U33440 ( .A1(n2429), .A2(REG0_REG_16__SCAN_IN), .ZN(n2640) );
  NOR2_X1 U33450 ( .A1(n2635), .A2(REG3_REG_16__SCAN_IN), .ZN(n2636) );
  OR2_X1 U33460 ( .A1(n2652), .A2(n2636), .ZN(n4405) );
  OR2_X1 U33470 ( .A1(n2822), .A2(n4405), .ZN(n2639) );
  INV_X1 U33480 ( .A(REG1_REG_16__SCAN_IN), .ZN(n2637) );
  OR2_X1 U33490 ( .A1(n3305), .A2(n2637), .ZN(n2638) );
  NAND2_X1 U33500 ( .A1(n2643), .A2(n2642), .ZN(n2644) );
  NAND2_X1 U33510 ( .A1(n2644), .A2(IR_REG_31__SCAN_IN), .ZN(n2645) );
  XNOR2_X1 U33520 ( .A(n2645), .B(IR_REG_16__SCAN_IN), .ZN(n4162) );
  MUX2_X1 U3353 ( .A(n4162), .B(DATAI_16_), .S(n3929), .Z(n4580) );
  OAI22_X1 U33540 ( .A1(n4575), .A2(n2672), .B1(n3827), .B2(n2751), .ZN(n2646)
         );
  XNOR2_X1 U3355 ( .A(n2646), .B(n2753), .ZN(n2648) );
  OAI22_X1 U3356 ( .A1(n4575), .A2(n2755), .B1(n3827), .B2(n2767), .ZN(n2647)
         );
  NOR2_X1 U3357 ( .A1(n2648), .A2(n2647), .ZN(n2651) );
  AOI21_X1 U3358 ( .B1(n2648), .B2(n2647), .A(n2651), .ZN(n3824) );
  NAND2_X1 U3359 ( .A1(n2429), .A2(REG0_REG_17__SCAN_IN), .ZN(n2657) );
  NAND2_X1 U3360 ( .A1(n3302), .A2(REG2_REG_17__SCAN_IN), .ZN(n2656) );
  INV_X1 U3361 ( .A(REG1_REG_17__SCAN_IN), .ZN(n4578) );
  OR2_X1 U3362 ( .A1(n3305), .A2(n4578), .ZN(n2655) );
  OR2_X1 U3363 ( .A1(n2652), .A2(REG3_REG_17__SCAN_IN), .ZN(n2653) );
  NAND2_X1 U3364 ( .A1(n2664), .A2(n2653), .ZN(n4391) );
  OR2_X1 U3365 ( .A1(n2822), .A2(n4391), .ZN(n2654) );
  NAND2_X1 U3366 ( .A1(n2658), .A2(IR_REG_31__SCAN_IN), .ZN(n2659) );
  XNOR2_X1 U3367 ( .A(n2659), .B(IR_REG_17__SCAN_IN), .ZN(n4165) );
  INV_X1 U3368 ( .A(DATAI_17_), .ZN(n2660) );
  MUX2_X1 U3369 ( .A(n4855), .B(n2660), .S(n3929), .Z(n4390) );
  OAI22_X1 U3370 ( .A1(n4409), .A2(n2672), .B1(n2751), .B2(n4390), .ZN(n2661)
         );
  XNOR2_X1 U3371 ( .A(n2661), .B(n2753), .ZN(n2663) );
  OAI22_X1 U3372 ( .A1(n4409), .A2(n2755), .B1(n2767), .B2(n4390), .ZN(n2662)
         );
  NAND2_X1 U3373 ( .A1(n2663), .A2(n2662), .ZN(n3832) );
  NOR2_X1 U3374 ( .A1(n2663), .A2(n2662), .ZN(n3833) );
  NAND2_X1 U3375 ( .A1(n2429), .A2(REG0_REG_18__SCAN_IN), .ZN(n2669) );
  NAND2_X1 U3376 ( .A1(n3302), .A2(REG2_REG_18__SCAN_IN), .ZN(n2668) );
  INV_X1 U3377 ( .A(REG1_REG_18__SCAN_IN), .ZN(n3063) );
  OR2_X1 U3378 ( .A1(n3305), .A2(n3063), .ZN(n2667) );
  NAND2_X1 U3379 ( .A1(n2664), .A2(n3085), .ZN(n2665) );
  NAND2_X1 U3380 ( .A1(n2687), .A2(n2665), .ZN(n4380) );
  OR2_X1 U3381 ( .A1(n2822), .A2(n4380), .ZN(n2666) );
  OR2_X1 U3382 ( .A1(n2670), .A2(n3293), .ZN(n2671) );
  XNOR2_X1 U3383 ( .A(n2671), .B(IR_REG_18__SCAN_IN), .ZN(n4714) );
  MUX2_X1 U3384 ( .A(n4714), .B(DATAI_18_), .S(n3929), .Z(n4374) );
  INV_X1 U3385 ( .A(n4374), .ZN(n4370) );
  OAI22_X1 U3386 ( .A1(n4395), .A2(n2672), .B1(n2751), .B2(n4370), .ZN(n2673)
         );
  XOR2_X1 U3387 ( .A(n2753), .B(n2673), .Z(n3890) );
  OAI22_X1 U3388 ( .A1(n4395), .A2(n2755), .B1(n2672), .B2(n4370), .ZN(n3889)
         );
  INV_X1 U3389 ( .A(n3889), .ZN(n2674) );
  NOR2_X1 U3390 ( .A1(n3890), .A2(n2674), .ZN(n2676) );
  INV_X1 U3391 ( .A(n3890), .ZN(n2675) );
  OAI21_X2 U3392 ( .B1(n3892), .B2(n2676), .A(n2354), .ZN(n3786) );
  NAND2_X1 U3393 ( .A1(n3302), .A2(REG2_REG_19__SCAN_IN), .ZN(n2680) );
  NAND2_X1 U3394 ( .A1(n2429), .A2(REG0_REG_19__SCAN_IN), .ZN(n2679) );
  INV_X1 U3395 ( .A(REG3_REG_19__SCAN_IN), .ZN(n3788) );
  XNOR2_X1 U3396 ( .A(n2687), .B(n3788), .ZN(n4360) );
  OR2_X1 U3397 ( .A1(n2822), .A2(n4360), .ZN(n2678) );
  INV_X1 U3398 ( .A(REG1_REG_19__SCAN_IN), .ZN(n4566) );
  OR2_X1 U3399 ( .A1(n3305), .A2(n4566), .ZN(n2677) );
  INV_X1 U3400 ( .A(DATAI_19_), .ZN(n2681) );
  MUX2_X1 U3401 ( .A(n4179), .B(n2681), .S(n3929), .Z(n4357) );
  OAI22_X1 U3402 ( .A1(n4329), .A2(n2755), .B1(n2752), .B2(n4357), .ZN(n2684)
         );
  OAI22_X1 U3403 ( .A1(n4329), .A2(n2752), .B1(n2751), .B2(n4357), .ZN(n2682)
         );
  XNOR2_X1 U3404 ( .A(n2682), .B(n2753), .ZN(n2683) );
  XOR2_X1 U3405 ( .A(n2684), .B(n2683), .Z(n3785) );
  INV_X1 U3406 ( .A(n2683), .ZN(n2686) );
  INV_X1 U3407 ( .A(n2684), .ZN(n2685) );
  INV_X1 U3408 ( .A(n2687), .ZN(n2688) );
  AOI21_X1 U3409 ( .B1(n2688), .B2(REG3_REG_19__SCAN_IN), .A(
        REG3_REG_20__SCAN_IN), .ZN(n2689) );
  OR2_X1 U3410 ( .A1(n2689), .A2(n2698), .ZN(n4337) );
  OR2_X1 U3411 ( .A1(n2822), .A2(n4337), .ZN(n2693) );
  INV_X1 U3412 ( .A(REG1_REG_20__SCAN_IN), .ZN(n4562) );
  OR2_X1 U3413 ( .A1(n3305), .A2(n4562), .ZN(n2692) );
  NAND2_X1 U3414 ( .A1(n3302), .A2(REG2_REG_20__SCAN_IN), .ZN(n2691) );
  NAND2_X1 U3415 ( .A1(n2429), .A2(REG0_REG_20__SCAN_IN), .ZN(n2690) );
  NAND2_X1 U3416 ( .A1(n4354), .A2(n2798), .ZN(n2695) );
  INV_X1 U3417 ( .A(n4336), .ZN(n4326) );
  NAND2_X1 U3418 ( .A1(n4326), .A2(n2799), .ZN(n2694) );
  NAND2_X1 U3419 ( .A1(n2695), .A2(n2694), .ZN(n2696) );
  XNOR2_X1 U3420 ( .A(n2696), .B(n2802), .ZN(n2709) );
  NOR2_X1 U3421 ( .A1(n4336), .A2(n2767), .ZN(n2697) );
  AOI21_X1 U3422 ( .B1(n4354), .B2(n2804), .A(n2697), .ZN(n2708) );
  NOR2_X1 U3423 ( .A1(n2709), .A2(n2708), .ZN(n3852) );
  NOR2_X1 U3424 ( .A1(n2698), .A2(REG3_REG_21__SCAN_IN), .ZN(n2699) );
  OR2_X1 U3425 ( .A1(n2720), .A2(n2699), .ZN(n3797) );
  OR2_X1 U3426 ( .A1(n2822), .A2(n3797), .ZN(n2703) );
  INV_X1 U3427 ( .A(REG1_REG_21__SCAN_IN), .ZN(n4557) );
  OR2_X1 U3428 ( .A1(n3305), .A2(n4557), .ZN(n2702) );
  NAND2_X1 U3429 ( .A1(n2429), .A2(REG0_REG_21__SCAN_IN), .ZN(n2701) );
  NAND2_X1 U3430 ( .A1(n3302), .A2(REG2_REG_21__SCAN_IN), .ZN(n2700) );
  NAND2_X1 U3431 ( .A1(n4327), .A2(n2798), .ZN(n2705) );
  INV_X1 U3432 ( .A(n4314), .ZN(n4550) );
  NAND2_X1 U3433 ( .A1(n4550), .A2(n2799), .ZN(n2704) );
  NAND2_X1 U3434 ( .A1(n2705), .A2(n2704), .ZN(n2706) );
  XNOR2_X1 U3435 ( .A(n2706), .B(n2802), .ZN(n3794) );
  NOR2_X1 U3436 ( .A1(n4314), .A2(n2767), .ZN(n2707) );
  AOI21_X1 U3437 ( .B1(n4327), .B2(n2804), .A(n2707), .ZN(n3793) );
  NAND2_X1 U3438 ( .A1(n2709), .A2(n2708), .ZN(n3851) );
  INV_X1 U3439 ( .A(REG1_REG_22__SCAN_IN), .ZN(n4548) );
  OR2_X1 U3440 ( .A1(n3305), .A2(n4548), .ZN(n2716) );
  XNOR2_X1 U3441 ( .A(n2720), .B(REG3_REG_22__SCAN_IN), .ZN(n3871) );
  OR2_X1 U3442 ( .A1(n2822), .A2(n3871), .ZN(n2715) );
  NAND2_X1 U3443 ( .A1(n2429), .A2(REG0_REG_22__SCAN_IN), .ZN(n2714) );
  NAND2_X1 U3444 ( .A1(n3302), .A2(REG2_REG_22__SCAN_IN), .ZN(n2713) );
  NAND4_X1 U3445 ( .A1(n2716), .A2(n2715), .A3(n2714), .A4(n2713), .ZN(n4551)
         );
  OAI22_X1 U3446 ( .A1(n4318), .A2(n2752), .B1(n4293), .B2(n2751), .ZN(n2717)
         );
  XNOR2_X1 U3447 ( .A(n2717), .B(n2753), .ZN(n2719) );
  OAI22_X1 U3448 ( .A1(n4318), .A2(n2755), .B1(n4293), .B2(n2767), .ZN(n2718)
         );
  XNOR2_X1 U3449 ( .A(n2719), .B(n2718), .ZN(n3870) );
  NOR2_X1 U3450 ( .A1(n2719), .A2(n2718), .ZN(n3778) );
  INV_X1 U3451 ( .A(REG1_REG_23__SCAN_IN), .ZN(n4542) );
  OR2_X1 U3452 ( .A1(n3305), .A2(n4542), .ZN(n2727) );
  NAND2_X1 U3453 ( .A1(n2720), .A2(REG3_REG_22__SCAN_IN), .ZN(n2722) );
  INV_X1 U3454 ( .A(REG3_REG_23__SCAN_IN), .ZN(n2721) );
  NAND2_X1 U3455 ( .A1(n2722), .A2(n2721), .ZN(n2723) );
  NAND2_X1 U3456 ( .A1(n2723), .A2(n2734), .ZN(n4286) );
  OR2_X1 U3457 ( .A1(n2822), .A2(n4286), .ZN(n2726) );
  NAND2_X1 U34580 ( .A1(n2429), .A2(REG0_REG_23__SCAN_IN), .ZN(n2725) );
  NAND2_X1 U34590 ( .A1(n3302), .A2(REG2_REG_23__SCAN_IN), .ZN(n2724) );
  NAND2_X1 U3460 ( .A1(n4533), .A2(n2798), .ZN(n2729) );
  NAND2_X1 U3461 ( .A1(n4283), .A2(n2799), .ZN(n2728) );
  NAND2_X1 U3462 ( .A1(n2729), .A2(n2728), .ZN(n2730) );
  XNOR2_X1 U3463 ( .A(n2730), .B(n2802), .ZN(n2733) );
  NOR2_X1 U3464 ( .A1(n4278), .A2(n2767), .ZN(n2731) );
  AOI21_X1 U3465 ( .B1(n4533), .B2(n2804), .A(n2731), .ZN(n2732) );
  XNOR2_X1 U3466 ( .A(n2733), .B(n2732), .ZN(n3777) );
  NOR2_X1 U34670 ( .A1(n2733), .A2(n2732), .ZN(n2742) );
  NAND2_X1 U3468 ( .A1(n3302), .A2(REG2_REG_24__SCAN_IN), .ZN(n2739) );
  NAND2_X1 U34690 ( .A1(n2429), .A2(REG0_REG_24__SCAN_IN), .ZN(n2738) );
  NAND2_X1 U3470 ( .A1(n2734), .A2(n3846), .ZN(n2735) );
  NAND2_X1 U34710 ( .A1(n2744), .A2(n2735), .ZN(n3845) );
  OR2_X1 U3472 ( .A1(n2822), .A2(n3845), .ZN(n2737) );
  INV_X1 U34730 ( .A(REG1_REG_24__SCAN_IN), .ZN(n4538) );
  OR2_X1 U3474 ( .A1(n3305), .A2(n4538), .ZN(n2736) );
  OAI22_X1 U34750 ( .A1(n4279), .A2(n2755), .B1(n2767), .B2(n4530), .ZN(n2741)
         );
  OR3_X2 U3476 ( .A1(n3776), .A2(n2742), .A3(n2741), .ZN(n3841) );
  OAI22_X1 U34770 ( .A1(n4279), .A2(n2752), .B1(n2751), .B2(n4530), .ZN(n2740)
         );
  XNOR2_X1 U3478 ( .A(n2740), .B(n2753), .ZN(n3844) );
  INV_X1 U34790 ( .A(n3842), .ZN(n2743) );
  AND2_X1 U3480 ( .A1(n2744), .A2(n3818), .ZN(n2745) );
  NOR2_X1 U34810 ( .A1(n2758), .A2(n2745), .ZN(n4245) );
  NAND2_X1 U3482 ( .A1(n4245), .A2(n2409), .ZN(n2750) );
  INV_X1 U34830 ( .A(REG1_REG_25__SCAN_IN), .ZN(n4528) );
  OR2_X1 U3484 ( .A1(n3305), .A2(n4528), .ZN(n2747) );
  NAND2_X1 U34850 ( .A1(n2429), .A2(REG0_REG_25__SCAN_IN), .ZN(n2746) );
  AND2_X1 U3486 ( .A1(n2747), .A2(n2746), .ZN(n2749) );
  NAND2_X1 U34870 ( .A1(n3302), .A2(REG2_REG_25__SCAN_IN), .ZN(n2748) );
  OAI22_X1 U3488 ( .A1(n4531), .A2(n2752), .B1(n2751), .B2(n4244), .ZN(n2754)
         );
  XNOR2_X1 U34890 ( .A(n2754), .B(n2753), .ZN(n2757) );
  OAI22_X1 U3490 ( .A1(n4531), .A2(n2755), .B1(n2767), .B2(n4244), .ZN(n2756)
         );
  NOR2_X1 U34910 ( .A1(n2757), .A2(n2756), .ZN(n3814) );
  NAND2_X1 U3492 ( .A1(n2757), .A2(n2756), .ZN(n3815) );
  INV_X1 U34930 ( .A(REG1_REG_26__SCAN_IN), .ZN(n3131) );
  OR2_X1 U3494 ( .A1(n2758), .A2(REG3_REG_26__SCAN_IN), .ZN(n2759) );
  NAND2_X1 U34950 ( .A1(n2793), .A2(n2759), .ZN(n4219) );
  OR2_X1 U3496 ( .A1(n4219), .A2(n2822), .ZN(n2763) );
  NAND2_X1 U34970 ( .A1(n3302), .A2(REG2_REG_26__SCAN_IN), .ZN(n2761) );
  NAND2_X1 U3498 ( .A1(n2429), .A2(REG0_REG_26__SCAN_IN), .ZN(n2760) );
  OAI211_X1 U34990 ( .C1(n3305), .C2(n3131), .A(n2763), .B(n2762), .ZN(n4510)
         );
  NAND2_X1 U3500 ( .A1(n4510), .A2(n2798), .ZN(n2765) );
  NAND2_X1 U35010 ( .A1(n4217), .A2(n2799), .ZN(n2764) );
  NAND2_X1 U3502 ( .A1(n2765), .A2(n2764), .ZN(n2766) );
  XNOR2_X1 U35030 ( .A(n2766), .B(n2802), .ZN(n2770) );
  NOR2_X1 U3504 ( .A1(n4518), .A2(n2767), .ZN(n2768) );
  AOI21_X1 U35050 ( .B1(n4510), .B2(n2804), .A(n2768), .ZN(n2769) );
  NOR2_X1 U35060 ( .A1(n2770), .A2(n2769), .ZN(n3900) );
  NAND2_X1 U35070 ( .A1(n2770), .A2(n2769), .ZN(n3901) );
  NAND2_X1 U35080 ( .A1(n2774), .A2(n2773), .ZN(n2771) );
  MUX2_X1 U35090 ( .A(n2774), .B(n2771), .S(B_REG_SCAN_IN), .Z(n2772) );
  INV_X1 U35100 ( .A(n4710), .ZN(n2775) );
  NAND2_X1 U35110 ( .A1(n2775), .A2(n2773), .ZN(n3285) );
  OAI21_X1 U35120 ( .B1(n3284), .B2(D_REG_1__SCAN_IN), .A(n3285), .ZN(n2947)
         );
  INV_X1 U35130 ( .A(n2947), .ZN(n3422) );
  INV_X1 U35140 ( .A(D_REG_0__SCAN_IN), .ZN(n3289) );
  NOR2_X1 U35150 ( .A1(D_REG_30__SCAN_IN), .A2(D_REG_19__SCAN_IN), .ZN(n2779)
         );
  NOR4_X1 U35160 ( .A1(D_REG_28__SCAN_IN), .A2(D_REG_29__SCAN_IN), .A3(
        D_REG_5__SCAN_IN), .A4(D_REG_10__SCAN_IN), .ZN(n2778) );
  NOR4_X1 U35170 ( .A1(D_REG_20__SCAN_IN), .A2(D_REG_3__SCAN_IN), .A3(
        D_REG_2__SCAN_IN), .A4(D_REG_11__SCAN_IN), .ZN(n2777) );
  NOR4_X1 U35180 ( .A1(D_REG_16__SCAN_IN), .A2(D_REG_12__SCAN_IN), .A3(
        D_REG_15__SCAN_IN), .A4(D_REG_4__SCAN_IN), .ZN(n2776) );
  NAND4_X1 U35190 ( .A1(n2779), .A2(n2778), .A3(n2777), .A4(n2776), .ZN(n2786)
         );
  NOR4_X1 U35200 ( .A1(D_REG_23__SCAN_IN), .A2(D_REG_6__SCAN_IN), .A3(
        D_REG_7__SCAN_IN), .A4(D_REG_8__SCAN_IN), .ZN(n2783) );
  NOR4_X1 U35210 ( .A1(D_REG_26__SCAN_IN), .A2(D_REG_17__SCAN_IN), .A3(
        D_REG_14__SCAN_IN), .A4(D_REG_27__SCAN_IN), .ZN(n2782) );
  NOR4_X1 U35220 ( .A1(D_REG_22__SCAN_IN), .A2(D_REG_24__SCAN_IN), .A3(
        D_REG_25__SCAN_IN), .A4(D_REG_31__SCAN_IN), .ZN(n2781) );
  NOR4_X1 U35230 ( .A1(D_REG_9__SCAN_IN), .A2(D_REG_13__SCAN_IN), .A3(
        D_REG_18__SCAN_IN), .A4(D_REG_21__SCAN_IN), .ZN(n2780) );
  NAND4_X1 U35240 ( .A1(n2783), .A2(n2782), .A3(n2781), .A4(n2780), .ZN(n2785)
         );
  NAND3_X1 U35250 ( .A1(n3422), .A2(n3251), .A3(n3420), .ZN(n2830) );
  INV_X1 U35260 ( .A(n4071), .ZN(n4713) );
  NAND2_X1 U35270 ( .A1(n3416), .A2(n4379), .ZN(n2789) );
  NAND2_X1 U35280 ( .A1(n4712), .A2(n4005), .ZN(n2938) );
  NAND2_X1 U35290 ( .A1(n2789), .A2(n2938), .ZN(n2790) );
  OR2_X1 U35300 ( .A1(n4627), .A2(n2790), .ZN(n2811) );
  INV_X1 U35310 ( .A(n2811), .ZN(n2791) );
  NAND2_X1 U35320 ( .A1(n3296), .A2(n2791), .ZN(n2792) );
  INV_X1 U35330 ( .A(REG1_REG_28__SCAN_IN), .ZN(n2797) );
  INV_X1 U35340 ( .A(REG3_REG_27__SCAN_IN), .ZN(n2839) );
  INV_X1 U35350 ( .A(REG3_REG_28__SCAN_IN), .ZN(n2827) );
  OAI21_X1 U35360 ( .B1(n2793), .B2(n2839), .A(n2827), .ZN(n2794) );
  NAND2_X1 U35370 ( .A1(n2794), .A2(n4192), .ZN(n3747) );
  OR2_X1 U35380 ( .A1(n3747), .A2(n2822), .ZN(n2796) );
  AOI22_X1 U35390 ( .A1(n3302), .A2(REG2_REG_28__SCAN_IN), .B1(n2429), .B2(
        REG0_REG_28__SCAN_IN), .ZN(n2795) );
  OAI211_X1 U35400 ( .C1(n3305), .C2(n2797), .A(n2796), .B(n2795), .ZN(n3348)
         );
  NAND2_X1 U35410 ( .A1(n3348), .A2(n2798), .ZN(n2801) );
  NAND2_X1 U35420 ( .A1(n3929), .A2(DATAI_28_), .ZN(n3233) );
  INV_X1 U35430 ( .A(n3233), .ZN(n2939) );
  NAND2_X1 U35440 ( .A1(n2939), .A2(n2799), .ZN(n2800) );
  NAND2_X1 U35450 ( .A1(n2801), .A2(n2800), .ZN(n2803) );
  XNOR2_X1 U35460 ( .A(n2803), .B(n2802), .ZN(n2807) );
  NAND2_X1 U35470 ( .A1(n3348), .A2(n2804), .ZN(n2805) );
  OAI21_X1 U35480 ( .B1(n2767), .B2(n3233), .A(n2805), .ZN(n2806) );
  INV_X1 U35490 ( .A(n2808), .ZN(n2809) );
  NAND3_X1 U35500 ( .A1(n2353), .A2(n2355), .A3(n3918), .ZN(n2836) );
  INV_X1 U35510 ( .A(n3747), .ZN(n2834) );
  NAND2_X1 U35520 ( .A1(n2811), .A2(n4876), .ZN(n2812) );
  NAND2_X1 U35530 ( .A1(n2830), .A2(n2812), .ZN(n3379) );
  AND2_X1 U35540 ( .A1(n4071), .A2(n4179), .ZN(n2813) );
  OR2_X1 U35550 ( .A1(n2938), .A2(n2813), .ZN(n2944) );
  AND3_X1 U35560 ( .A1(n2417), .A2(n2944), .A3(n3300), .ZN(n2814) );
  AOI21_X1 U35570 ( .B1(n3379), .B2(n2814), .A(U3149), .ZN(n2819) );
  INV_X1 U35580 ( .A(n2815), .ZN(n2816) );
  AND2_X1 U35590 ( .A1(n4853), .A2(n2816), .ZN(n2817) );
  AND2_X1 U35600 ( .A1(n2830), .A2(n4078), .ZN(n3377) );
  AOI22_X1 U35610 ( .A1(n3302), .A2(REG2_REG_29__SCAN_IN), .B1(n2429), .B2(
        REG0_REG_29__SCAN_IN), .ZN(n2821) );
  NAND2_X1 U35620 ( .A1(n2408), .A2(REG1_REG_29__SCAN_IN), .ZN(n2820) );
  OAI211_X1 U35630 ( .C1(n4192), .C2(n2822), .A(n2821), .B(n2820), .ZN(n4085)
         );
  INV_X1 U35640 ( .A(n4085), .ZN(n3939) );
  OR2_X1 U35650 ( .A1(n2823), .A2(n3293), .ZN(n2825) );
  NAND2_X1 U35660 ( .A1(n4078), .A2(n4722), .ZN(n2826) );
  OAI22_X1 U35670 ( .A1(n3939), .A2(n3923), .B1(STATE_REG_SCAN_IN), .B2(n2827), 
        .ZN(n2833) );
  INV_X1 U35680 ( .A(n4520), .ZN(n4223) );
  NAND2_X1 U35690 ( .A1(n3402), .A2(n4078), .ZN(n2828) );
  OR2_X2 U35700 ( .A1(n2830), .A2(n2828), .ZN(n3921) );
  NAND2_X1 U35710 ( .A1(n3296), .A2(n4627), .ZN(n2829) );
  OR2_X1 U35720 ( .A1(n2830), .A2(n2829), .ZN(n2831) );
  NAND2_X1 U35730 ( .A1(n4071), .A2(n4379), .ZN(n3419) );
  OR2_X1 U35740 ( .A1(n3419), .A2(n4712), .ZN(n4884) );
  NAND2_X1 U35750 ( .A1(n2831), .A2(n4478), .ZN(n3465) );
  INV_X2 U35760 ( .A(n3465), .ZN(n3920) );
  OAI22_X1 U35770 ( .A1(n4223), .A2(n3921), .B1(n3920), .B2(n3233), .ZN(n2832)
         );
  AOI211_X1 U35780 ( .C1(n2834), .C2(n3895), .A(n2833), .B(n2832), .ZN(n2835)
         );
  XNOR2_X1 U35790 ( .A(n2838), .B(n2201), .ZN(n2843) );
  OAI22_X1 U35800 ( .A1(n4238), .A2(n3921), .B1(n3920), .B2(n4209), .ZN(n2841)
         );
  OAI22_X1 U35810 ( .A1(n4513), .A2(n3923), .B1(STATE_REG_SCAN_IN), .B2(n2839), 
        .ZN(n2840) );
  AOI211_X1 U3582 ( .C1(n4207), .C2(n3895), .A(n2841), .B(n2840), .ZN(n2842)
         );
  OAI21_X1 U3583 ( .B1(n2843), .B2(n3898), .A(n2842), .ZN(U3211) );
  NAND3_X1 U3584 ( .A1(n2846), .A2(n2844), .A3(n2845), .ZN(n2849) );
  OAI21_X2 U3585 ( .B1(n2849), .B2(n2848), .A(n3446), .ZN(n4003) );
  INV_X1 U3586 ( .A(n4091), .ZN(n3454) );
  NAND2_X1 U3587 ( .A1(n3375), .A2(n3456), .ZN(n2851) );
  INV_X1 U3588 ( .A(n2852), .ZN(n4090) );
  NAND2_X1 U3589 ( .A1(n4090), .A2(n4877), .ZN(n4010) );
  NAND2_X1 U3590 ( .A1(n2852), .A2(n3532), .ZN(n4007) );
  NAND2_X1 U3591 ( .A1(n2852), .A2(n4877), .ZN(n2853) );
  NAND2_X1 U3592 ( .A1(n3551), .A2(n3542), .ZN(n2854) );
  NAND2_X1 U3593 ( .A1(n3482), .A2(n2854), .ZN(n2856) );
  NAND2_X1 U3594 ( .A1(n4879), .A2(n3475), .ZN(n2855) );
  NAND2_X1 U3595 ( .A1(n2857), .A2(n2858), .ZN(n4013) );
  NAND2_X1 U3596 ( .A1(n4089), .A2(n3555), .ZN(n4017) );
  AND2_X1 U3597 ( .A1(n2859), .A2(n3611), .ZN(n2861) );
  NAND2_X1 U3598 ( .A1(n4089), .A2(n2858), .ZN(n3496) );
  NAND2_X1 U3599 ( .A1(n4088), .A2(n3506), .ZN(n2860) );
  AND2_X1 U3600 ( .A1(n3496), .A2(n2860), .ZN(n2862) );
  AND2_X1 U3601 ( .A1(n3676), .A2(n3621), .ZN(n2864) );
  NAND2_X1 U3602 ( .A1(n3657), .A2(n2866), .ZN(n2908) );
  NAND2_X1 U3603 ( .A1(n4087), .A2(n3671), .ZN(n4028) );
  NAND2_X1 U3604 ( .A1(n4087), .A2(n2866), .ZN(n2867) );
  NAND2_X1 U3605 ( .A1(n3741), .A2(n3700), .ZN(n2868) );
  NAND2_X1 U3606 ( .A1(n3667), .A2(n2911), .ZN(n2869) );
  INV_X1 U3607 ( .A(n3710), .ZN(n3740) );
  NAND2_X1 U3608 ( .A1(n3721), .A2(n3740), .ZN(n2870) );
  NOR2_X1 U3609 ( .A1(n4629), .A2(n3718), .ZN(n2872) );
  INV_X1 U3610 ( .A(n4629), .ZN(n3884) );
  NAND2_X1 U3611 ( .A1(n4616), .A2(n4628), .ZN(n4449) );
  INV_X1 U3612 ( .A(n4616), .ZN(n3719) );
  NAND2_X1 U3613 ( .A1(n3719), .A2(n3883), .ZN(n4451) );
  NAND2_X1 U3614 ( .A1(n4616), .A2(n3883), .ZN(n2874) );
  NAND2_X1 U3615 ( .A1(n4605), .A2(n2876), .ZN(n3942) );
  NAND2_X1 U3616 ( .A1(n4423), .A2(n4443), .ZN(n3943) );
  NAND2_X1 U3617 ( .A1(n3942), .A2(n3943), .ZN(n4434) );
  NAND2_X1 U3618 ( .A1(n4575), .A2(n4580), .ZN(n4050) );
  NAND2_X1 U3619 ( .A1(n4593), .A2(n3827), .ZN(n3946) );
  NAND2_X1 U3620 ( .A1(n4050), .A2(n3946), .ZN(n4401) );
  NAND2_X1 U3621 ( .A1(n4409), .A2(n4390), .ZN(n2880) );
  AOI21_X1 U3622 ( .B1(n4386), .B2(n2880), .A(n2879), .ZN(n4365) );
  NAND2_X1 U3623 ( .A1(n4572), .A2(n4370), .ZN(n4349) );
  NAND2_X1 U3624 ( .A1(n4395), .A2(n4374), .ZN(n4348) );
  NAND2_X1 U3625 ( .A1(n4349), .A2(n4348), .ZN(n4373) );
  NAND2_X1 U3626 ( .A1(n4365), .A2(n4373), .ZN(n4366) );
  NAND2_X1 U3627 ( .A1(n4354), .A2(n4326), .ZN(n3966) );
  NAND2_X1 U3628 ( .A1(n4553), .A2(n4336), .ZN(n3967) );
  NAND2_X1 U3629 ( .A1(n3873), .A2(n4314), .ZN(n2885) );
  NAND2_X1 U3630 ( .A1(n4551), .A2(n4293), .ZN(n2930) );
  INV_X1 U3631 ( .A(n2930), .ZN(n2886) );
  NAND2_X1 U3632 ( .A1(n4318), .A2(n4298), .ZN(n2931) );
  INV_X1 U3633 ( .A(n2931), .ZN(n4275) );
  NAND2_X1 U3634 ( .A1(n4551), .A2(n4298), .ZN(n2888) );
  NAND2_X1 U3635 ( .A1(n4546), .A2(n2888), .ZN(n4267) );
  NAND2_X1 U3636 ( .A1(n4267), .A2(n2889), .ZN(n2891) );
  NAND2_X1 U3637 ( .A1(n4533), .A2(n4283), .ZN(n2890) );
  NOR2_X1 U3638 ( .A1(n4279), .A2(n4530), .ZN(n2893) );
  NAND2_X1 U3639 ( .A1(n4279), .A2(n4530), .ZN(n2892) );
  INV_X1 U3640 ( .A(n4244), .ZN(n2936) );
  NAND2_X1 U3641 ( .A1(n4218), .A2(n2936), .ZN(n2894) );
  NAND2_X1 U3642 ( .A1(n2895), .A2(n2894), .ZN(n4216) );
  NOR2_X1 U3643 ( .A1(n4238), .A2(n4518), .ZN(n2897) );
  NAND2_X1 U3644 ( .A1(n4238), .A2(n4518), .ZN(n2896) );
  NOR2_X1 U3645 ( .A1(n4520), .A2(n4509), .ZN(n2899) );
  NAND2_X1 U3646 ( .A1(n4520), .A2(n4509), .ZN(n2898) );
  NAND2_X1 U3647 ( .A1(n4513), .A2(n2939), .ZN(n3954) );
  NAND2_X1 U3648 ( .A1(n3348), .A2(n3233), .ZN(n3933) );
  NAND2_X1 U3649 ( .A1(n3954), .A2(n3933), .ZN(n3964) );
  XNOR2_X1 U3650 ( .A(n4712), .B(n3425), .ZN(n2900) );
  NAND2_X1 U3651 ( .A1(n2900), .A2(n4179), .ZN(n4333) );
  NAND2_X1 U3652 ( .A1(n3446), .A2(n3447), .ZN(n3528) );
  NOR2_X1 U3653 ( .A1(n3528), .A2(n3532), .ZN(n3527) );
  INV_X1 U3654 ( .A(n4205), .ZN(n2901) );
  AOI21_X1 U3655 ( .B1(n2939), .B2(n2901), .A(n3246), .ZN(n3749) );
  NAND2_X1 U3656 ( .A1(n3454), .A2(n3376), .ZN(n4002) );
  OR2_X1 U3657 ( .A1(n2902), .A2(n4002), .ZN(n3520) );
  NAND2_X1 U3658 ( .A1(n3520), .A2(n2903), .ZN(n2904) );
  INV_X1 U3659 ( .A(n3521), .ZN(n3978) );
  NAND2_X1 U3660 ( .A1(n2904), .A2(n3978), .ZN(n3523) );
  NAND2_X1 U3661 ( .A1(n3523), .A2(n4007), .ZN(n3485) );
  NAND2_X1 U3662 ( .A1(n4879), .A2(n3542), .ZN(n4012) );
  NAND2_X1 U3663 ( .A1(n3551), .A2(n3475), .ZN(n4009) );
  NAND2_X1 U3664 ( .A1(n3485), .A2(n3992), .ZN(n3484) );
  NAND2_X1 U3665 ( .A1(n3484), .A2(n4012), .ZN(n3548) );
  INV_X1 U3666 ( .A(n4013), .ZN(n2905) );
  OR2_X1 U3667 ( .A1(n3548), .A2(n2905), .ZN(n2906) );
  NAND2_X1 U3668 ( .A1(n2906), .A2(n4017), .ZN(n3502) );
  AND2_X1 U3669 ( .A1(n4088), .A2(n3611), .ZN(n3497) );
  NAND2_X1 U3670 ( .A1(n2859), .A2(n3506), .ZN(n4029) );
  INV_X1 U3671 ( .A(n3621), .ZN(n3758) );
  NAND2_X1 U3672 ( .A1(n3676), .A2(n3758), .ZN(n4031) );
  NAND2_X1 U3673 ( .A1(n3617), .A2(n4031), .ZN(n2907) );
  INV_X1 U3674 ( .A(n3676), .ZN(n3664) );
  NAND2_X1 U3675 ( .A1(n3664), .A2(n3621), .ZN(n4018) );
  NAND2_X1 U3676 ( .A1(n2907), .A2(n4018), .ZN(n3672) );
  INV_X1 U3677 ( .A(n2908), .ZN(n2909) );
  OR2_X1 U3678 ( .A1(n3672), .A2(n2909), .ZN(n2910) );
  NAND2_X1 U3679 ( .A1(n2910), .A2(n4028), .ZN(n3699) );
  NAND2_X1 U3680 ( .A1(n3741), .A2(n2911), .ZN(n4022) );
  NAND2_X1 U3681 ( .A1(n3699), .A2(n4022), .ZN(n2912) );
  NAND2_X1 U3682 ( .A1(n3667), .A2(n3700), .ZN(n4032) );
  NAND2_X1 U3683 ( .A1(n2912), .A2(n4032), .ZN(n3639) );
  AND2_X1 U3684 ( .A1(n4086), .A2(n3740), .ZN(n4026) );
  OR2_X1 U3685 ( .A1(n3639), .A2(n4026), .ZN(n2913) );
  NAND2_X1 U3686 ( .A1(n3721), .A2(n3710), .ZN(n4023) );
  NAND2_X1 U3687 ( .A1(n2913), .A2(n4023), .ZN(n3717) );
  NAND2_X1 U3688 ( .A1(n4629), .A2(n3726), .ZN(n4038) );
  NAND2_X1 U3689 ( .A1(n3717), .A2(n4038), .ZN(n2914) );
  NAND2_X1 U3690 ( .A1(n3884), .A2(n3718), .ZN(n4037) );
  NAND2_X1 U3691 ( .A1(n2914), .A2(n4037), .ZN(n4452) );
  NAND2_X1 U3692 ( .A1(n4607), .A2(n4613), .ZN(n4453) );
  NAND2_X1 U3693 ( .A1(n4481), .A2(n4604), .ZN(n2915) );
  NAND2_X1 U3694 ( .A1(n4453), .A2(n2915), .ZN(n2917) );
  INV_X1 U3695 ( .A(n4451), .ZN(n2916) );
  NOR2_X1 U3696 ( .A1(n2917), .A2(n2916), .ZN(n4039) );
  NAND2_X1 U3697 ( .A1(n4452), .A2(n4039), .ZN(n2921) );
  NAND2_X1 U3698 ( .A1(n4632), .A2(n4475), .ZN(n4455) );
  NAND2_X1 U3699 ( .A1(n4449), .A2(n4455), .ZN(n2920) );
  INV_X1 U3700 ( .A(n2917), .ZN(n2919) );
  NOR2_X1 U3701 ( .A1(n4481), .A2(n4604), .ZN(n2918) );
  AOI21_X1 U3702 ( .B1(n2920), .B2(n2919), .A(n2918), .ZN(n4042) );
  NAND2_X1 U3703 ( .A1(n2921), .A2(n4042), .ZN(n4432) );
  INV_X1 U3704 ( .A(n4434), .ZN(n3980) );
  NAND2_X1 U3705 ( .A1(n4432), .A2(n3980), .ZN(n2922) );
  NAND2_X1 U3706 ( .A1(n2922), .A2(n3942), .ZN(n4416) );
  NAND2_X1 U3707 ( .A1(n4583), .A2(n4591), .ZN(n3945) );
  NAND2_X1 U3708 ( .A1(n4404), .A2(n4422), .ZN(n3944) );
  NAND2_X1 U3709 ( .A1(n3945), .A2(n3944), .ZN(n4419) );
  NAND2_X1 U3710 ( .A1(n4417), .A2(n3944), .ZN(n4411) );
  NAND2_X1 U3711 ( .A1(n4411), .A2(n2326), .ZN(n4410) );
  NAND2_X1 U3712 ( .A1(n4410), .A2(n3946), .ZN(n4384) );
  NAND2_X1 U3713 ( .A1(n4409), .A2(n4571), .ZN(n4346) );
  NAND2_X1 U3714 ( .A1(n4348), .A2(n4346), .ZN(n2925) );
  NAND2_X1 U3715 ( .A1(n4375), .A2(n4357), .ZN(n2923) );
  AND2_X1 U3716 ( .A1(n4349), .A2(n2923), .ZN(n2926) );
  NOR2_X1 U3717 ( .A1(n4375), .A2(n4357), .ZN(n2924) );
  AOI21_X1 U3718 ( .B1(n2925), .B2(n2926), .A(n2924), .ZN(n4269) );
  NAND2_X1 U3719 ( .A1(n4553), .A2(n4326), .ZN(n4272) );
  NAND2_X1 U3720 ( .A1(n4384), .A2(n3948), .ZN(n2927) );
  NAND2_X1 U3721 ( .A1(n4581), .A2(n4390), .ZN(n4345) );
  NAND2_X1 U3722 ( .A1(n2926), .A2(n4345), .ZN(n4268) );
  AND2_X1 U3723 ( .A1(n4354), .A2(n4336), .ZN(n4052) );
  AOI21_X1 U3724 ( .B1(n3948), .B2(n4268), .A(n4052), .ZN(n3949) );
  NAND2_X1 U3725 ( .A1(n2927), .A2(n3949), .ZN(n2928) );
  NAND2_X1 U3726 ( .A1(n3873), .A2(n4550), .ZN(n4274) );
  AND2_X1 U3727 ( .A1(n4274), .A2(n2931), .ZN(n4058) );
  NAND2_X1 U3728 ( .A1(n2928), .A2(n4058), .ZN(n2935) );
  NAND2_X1 U3729 ( .A1(n4533), .A2(n4278), .ZN(n2929) );
  NAND2_X1 U3730 ( .A1(n2930), .A2(n2929), .ZN(n4059) );
  INV_X1 U3731 ( .A(n4059), .ZN(n2933) );
  AND2_X1 U3732 ( .A1(n4327), .A2(n4314), .ZN(n3990) );
  NAND2_X1 U3733 ( .A1(n2931), .A2(n3990), .ZN(n2932) );
  NAND2_X1 U3734 ( .A1(n2933), .A2(n2932), .ZN(n3952) );
  INV_X1 U3735 ( .A(n3952), .ZN(n2934) );
  NAND2_X1 U3736 ( .A1(n2935), .A2(n2934), .ZN(n4259) );
  INV_X1 U3737 ( .A(n4533), .ZN(n4294) );
  NAND2_X1 U3738 ( .A1(n4294), .A2(n4283), .ZN(n4258) );
  INV_X1 U3739 ( .A(n4530), .ZN(n4254) );
  NAND2_X1 U3740 ( .A1(n4279), .A2(n4254), .ZN(n3965) );
  NAND2_X1 U3741 ( .A1(n4259), .A2(n4056), .ZN(n4235) );
  NAND2_X1 U3742 ( .A1(n4218), .A2(n4244), .ZN(n3976) );
  INV_X1 U3743 ( .A(n4279), .ZN(n4240) );
  NAND2_X1 U3744 ( .A1(n4240), .A2(n4530), .ZN(n4234) );
  NAND2_X1 U3745 ( .A1(n4235), .A2(n4062), .ZN(n4225) );
  NAND2_X1 U3746 ( .A1(n4238), .A2(n4217), .ZN(n3969) );
  NAND2_X1 U3747 ( .A1(n4531), .A2(n2936), .ZN(n4224) );
  AND2_X1 U3748 ( .A1(n4510), .A2(n4518), .ZN(n4066) );
  AOI21_X1 U3749 ( .B1(n4225), .B2(n4001), .A(n4066), .ZN(n4200) );
  NAND2_X1 U3750 ( .A1(n4520), .A2(n4209), .ZN(n4060) );
  NAND2_X1 U3751 ( .A1(n3953), .A2(n4060), .ZN(n4203) );
  INV_X1 U3752 ( .A(n4203), .ZN(n4201) );
  NAND2_X1 U3753 ( .A1(n4200), .A2(n4201), .ZN(n4199) );
  NAND2_X1 U3754 ( .A1(n4199), .A2(n3953), .ZN(n3237) );
  XNOR2_X1 U3755 ( .A(n3237), .B(n3964), .ZN(n2942) );
  NAND2_X1 U3756 ( .A1(n4712), .A2(n4379), .ZN(n2937) );
  NAND2_X1 U3757 ( .A1(n4713), .A2(n4005), .ZN(n4075) );
  AOI22_X1 U3758 ( .A1(n4085), .A2(n4592), .B1(n4627), .B2(n2939), .ZN(n2941)
         );
  NAND2_X1 U3759 ( .A1(n4520), .A2(n4881), .ZN(n2940) );
  OAI211_X1 U3760 ( .C1(n2942), .C2(n4637), .A(n2941), .B(n2940), .ZN(n3750)
         );
  NAND2_X1 U3761 ( .A1(n3296), .A2(n2944), .ZN(n3378) );
  NOR2_X1 U3762 ( .A1(n3378), .A2(n2945), .ZN(n2946) );
  INV_X1 U3763 ( .A(n3251), .ZN(n3423) );
  INV_X1 U3764 ( .A(REG0_REG_28__SCAN_IN), .ZN(n2948) );
  NAND2_X1 U3765 ( .A1(keyinput99), .A2(keyinput103), .ZN(n2949) );
  NOR3_X1 U3766 ( .A1(keyinput102), .A2(keyinput98), .A3(n2949), .ZN(n2956) );
  INV_X1 U3767 ( .A(keyinput110), .ZN(n2950) );
  NOR4_X1 U3768 ( .A1(keyinput111), .A2(keyinput106), .A3(keyinput107), .A4(
        n2950), .ZN(n2955) );
  NAND2_X1 U3769 ( .A1(keyinput66), .A2(keyinput70), .ZN(n2951) );
  NOR3_X1 U3770 ( .A1(keyinput71), .A2(keyinput67), .A3(n2951), .ZN(n2954) );
  INV_X1 U3771 ( .A(keyinput74), .ZN(n2952) );
  NOR4_X1 U3772 ( .A1(keyinput79), .A2(keyinput78), .A3(keyinput75), .A4(n2952), .ZN(n2953) );
  AND4_X1 U3773 ( .A1(n2956), .A2(n2955), .A3(n2954), .A4(n2953), .ZN(n2997)
         );
  NOR2_X1 U3774 ( .A1(keyinput119), .A2(keyinput115), .ZN(n2957) );
  NAND3_X1 U3775 ( .A1(keyinput118), .A2(keyinput114), .A3(n2957), .ZN(n2964)
         );
  INV_X1 U3776 ( .A(keyinput126), .ZN(n2958) );
  NAND4_X1 U3777 ( .A1(keyinput123), .A2(keyinput122), .A3(keyinput127), .A4(
        n2958), .ZN(n2963) );
  INV_X1 U3778 ( .A(keyinput87), .ZN(n2959) );
  NAND4_X1 U3779 ( .A1(keyinput86), .A2(keyinput82), .A3(keyinput83), .A4(
        n2959), .ZN(n2962) );
  NOR2_X1 U3780 ( .A1(keyinput95), .A2(keyinput91), .ZN(n2960) );
  NAND3_X1 U3781 ( .A1(keyinput94), .A2(keyinput90), .A3(n2960), .ZN(n2961) );
  NOR4_X1 U3782 ( .A1(n2964), .A2(n2963), .A3(n2962), .A4(n2961), .ZN(n2996)
         );
  NAND2_X1 U3783 ( .A1(keyinput64), .A2(keyinput33), .ZN(n2965) );
  NOR3_X1 U3784 ( .A1(keyinput77), .A2(keyinput32), .A3(n2965), .ZN(n2966) );
  NAND3_X1 U3785 ( .A1(keyinput8), .A2(keyinput85), .A3(n2966), .ZN(n2979) );
  NAND2_X1 U3786 ( .A1(keyinput124), .A2(keyinput9), .ZN(n2967) );
  NOR3_X1 U3787 ( .A1(keyinput13), .A2(keyinput24), .A3(n2967), .ZN(n2977) );
  NOR4_X1 U3788 ( .A1(keyinput96), .A2(keyinput12), .A3(keyinput1), .A4(
        keyinput49), .ZN(n2976) );
  NAND4_X1 U3789 ( .A1(keyinput81), .A2(keyinput120), .A3(keyinput108), .A4(
        keyinput100), .ZN(n2974) );
  NOR2_X1 U3790 ( .A1(keyinput117), .A2(keyinput112), .ZN(n2968) );
  NAND3_X1 U3791 ( .A1(keyinput29), .A2(keyinput72), .A3(n2968), .ZN(n2973) );
  NOR2_X1 U3792 ( .A1(keyinput68), .A2(keyinput37), .ZN(n2969) );
  NAND3_X1 U3793 ( .A1(keyinput53), .A2(keyinput101), .A3(n2969), .ZN(n2972)
         );
  NOR2_X1 U3794 ( .A1(keyinput57), .A2(keyinput109), .ZN(n2970) );
  NAND3_X1 U3795 ( .A1(keyinput80), .A2(keyinput41), .A3(n2970), .ZN(n2971) );
  NOR4_X1 U3796 ( .A1(n2974), .A2(n2973), .A3(n2972), .A4(n2971), .ZN(n2975)
         );
  NAND3_X1 U3797 ( .A1(n2977), .A2(n2976), .A3(n2975), .ZN(n2978) );
  NOR4_X1 U3798 ( .A1(keyinput97), .A2(keyinput116), .A3(n2979), .A4(n2978), 
        .ZN(n2995) );
  NAND2_X1 U3799 ( .A1(keyinput73), .A2(keyinput121), .ZN(n2980) );
  NOR3_X1 U3800 ( .A1(keyinput45), .A2(keyinput88), .A3(n2980), .ZN(n2981) );
  NAND3_X1 U3801 ( .A1(keyinput56), .A2(keyinput5), .A3(n2981), .ZN(n2993) );
  NAND2_X1 U3802 ( .A1(keyinput65), .A2(keyinput21), .ZN(n2982) );
  NOR3_X1 U3803 ( .A1(keyinput125), .A2(keyinput104), .A3(n2982), .ZN(n2991)
         );
  INV_X1 U3804 ( .A(keyinput28), .ZN(n2983) );
  NOR4_X1 U3805 ( .A1(keyinput69), .A2(keyinput0), .A3(keyinput76), .A4(n2983), 
        .ZN(n2990) );
  NAND4_X1 U3806 ( .A1(keyinput36), .A2(keyinput93), .A3(keyinput16), .A4(
        keyinput61), .ZN(n2988) );
  OR4_X1 U3807 ( .A1(keyinput60), .A2(keyinput25), .A3(keyinput40), .A4(
        keyinput44), .ZN(n2987) );
  NAND4_X1 U3808 ( .A1(keyinput48), .A2(keyinput52), .A3(keyinput20), .A4(
        keyinput17), .ZN(n2986) );
  NOR2_X1 U3809 ( .A1(keyinput84), .A2(keyinput89), .ZN(n2984) );
  NAND3_X1 U3810 ( .A1(keyinput92), .A2(keyinput105), .A3(n2984), .ZN(n2985)
         );
  NOR4_X1 U3811 ( .A1(n2988), .A2(n2987), .A3(n2986), .A4(n2985), .ZN(n2989)
         );
  NAND3_X1 U3812 ( .A1(n2991), .A2(n2990), .A3(n2989), .ZN(n2992) );
  NOR4_X1 U3813 ( .A1(keyinput113), .A2(keyinput4), .A3(n2993), .A4(n2992), 
        .ZN(n2994) );
  NAND4_X1 U3814 ( .A1(n2997), .A2(n2996), .A3(n2995), .A4(n2994), .ZN(n3231)
         );
  NOR4_X1 U3815 ( .A1(keyinput58), .A2(keyinput59), .A3(keyinput51), .A4(
        keyinput50), .ZN(n2998) );
  NAND3_X1 U3816 ( .A1(keyinput54), .A2(keyinput55), .A3(n2998), .ZN(n2999) );
  NOR3_X1 U3817 ( .A1(keyinput62), .A2(keyinput63), .A3(n2999), .ZN(n3011) );
  NOR4_X1 U3818 ( .A1(keyinput26), .A2(keyinput27), .A3(keyinput18), .A4(
        keyinput19), .ZN(n3010) );
  NAND2_X1 U3819 ( .A1(keyinput23), .A2(keyinput31), .ZN(n3000) );
  NOR3_X1 U3820 ( .A1(keyinput30), .A2(keyinput22), .A3(n3000), .ZN(n3009) );
  NOR2_X1 U3821 ( .A1(keyinput35), .A2(keyinput38), .ZN(n3001) );
  NAND3_X1 U3822 ( .A1(keyinput39), .A2(keyinput34), .A3(n3001), .ZN(n3007) );
  NAND4_X1 U3823 ( .A1(keyinput46), .A2(keyinput47), .A3(keyinput43), .A4(
        keyinput42), .ZN(n3006) );
  NOR2_X1 U3824 ( .A1(keyinput2), .A2(keyinput6), .ZN(n3002) );
  NAND3_X1 U3825 ( .A1(keyinput7), .A2(keyinput3), .A3(n3002), .ZN(n3005) );
  NOR2_X1 U3826 ( .A1(keyinput14), .A2(keyinput10), .ZN(n3003) );
  NAND3_X1 U3827 ( .A1(keyinput15), .A2(keyinput11), .A3(n3003), .ZN(n3004) );
  NOR4_X1 U3828 ( .A1(n3007), .A2(n3006), .A3(n3005), .A4(n3004), .ZN(n3008)
         );
  NAND4_X1 U3829 ( .A1(n3011), .A2(n3010), .A3(n3009), .A4(n3008), .ZN(n3230)
         );
  INV_X1 U3830 ( .A(REG2_REG_11__SCAN_IN), .ZN(n3688) );
  INV_X1 U3831 ( .A(keyinput26), .ZN(n3013) );
  AOI22_X1 U3832 ( .A1(n3688), .A2(keyinput27), .B1(ADDR_REG_18__SCAN_IN), 
        .B2(n3013), .ZN(n3012) );
  OAI221_X1 U3833 ( .B1(n3688), .B2(keyinput27), .C1(n3013), .C2(
        ADDR_REG_18__SCAN_IN), .A(n3012), .ZN(n3018) );
  INV_X1 U3834 ( .A(keyinput14), .ZN(n3016) );
  INV_X1 U3835 ( .A(keyinput15), .ZN(n3015) );
  AOI22_X1 U3836 ( .A1(n3016), .A2(DATAO_REG_8__SCAN_IN), .B1(
        DATAO_REG_11__SCAN_IN), .B2(n3015), .ZN(n3014) );
  OAI221_X1 U3837 ( .B1(n3016), .B2(DATAO_REG_8__SCAN_IN), .C1(n3015), .C2(
        DATAO_REG_11__SCAN_IN), .A(n3014), .ZN(n3017) );
  NOR2_X1 U3838 ( .A1(n3018), .A2(n3017), .ZN(n3039) );
  INV_X1 U3839 ( .A(REG0_REG_23__SCAN_IN), .ZN(n3020) );
  AOI22_X1 U3840 ( .A1(n3020), .A2(keyinput40), .B1(keyinput44), .B2(n4516), 
        .ZN(n3019) );
  OAI221_X1 U3841 ( .B1(n3020), .B2(keyinput40), .C1(n4516), .C2(keyinput44), 
        .A(n3019), .ZN(n3025) );
  INV_X1 U3842 ( .A(keyinput54), .ZN(n3023) );
  INV_X1 U3843 ( .A(keyinput55), .ZN(n3022) );
  AOI22_X1 U3844 ( .A1(n3023), .A2(DATAO_REG_13__SCAN_IN), .B1(
        DATAO_REG_19__SCAN_IN), .B2(n3022), .ZN(n3021) );
  OAI221_X1 U3845 ( .B1(n3023), .B2(DATAO_REG_13__SCAN_IN), .C1(n3022), .C2(
        DATAO_REG_19__SCAN_IN), .A(n3021), .ZN(n3024) );
  NOR2_X1 U3846 ( .A1(n3025), .A2(n3024), .ZN(n3038) );
  INV_X1 U3847 ( .A(REG0_REG_22__SCAN_IN), .ZN(n4667) );
  INV_X1 U3848 ( .A(D_REG_12__SCAN_IN), .ZN(n4844) );
  AOI22_X1 U3849 ( .A1(n4667), .A2(keyinput62), .B1(n4844), .B2(keyinput63), 
        .ZN(n3026) );
  OAI221_X1 U3850 ( .B1(n4667), .B2(keyinput62), .C1(n4844), .C2(keyinput63), 
        .A(n3026), .ZN(n3030) );
  INV_X1 U3851 ( .A(REG0_REG_25__SCAN_IN), .ZN(n3028) );
  INV_X1 U3852 ( .A(D_REG_15__SCAN_IN), .ZN(n4842) );
  AOI22_X1 U3853 ( .A1(n3028), .A2(keyinput58), .B1(n4842), .B2(keyinput59), 
        .ZN(n3027) );
  OAI221_X1 U3854 ( .B1(n3028), .B2(keyinput58), .C1(n4842), .C2(keyinput59), 
        .A(n3027), .ZN(n3029) );
  NOR2_X1 U3855 ( .A1(n3030), .A2(n3029), .ZN(n3037) );
  INV_X1 U3856 ( .A(DATAI_16_), .ZN(n4856) );
  AOI22_X1 U3857 ( .A1(n4856), .A2(keyinput28), .B1(n2660), .B2(keyinput76), 
        .ZN(n3031) );
  OAI221_X1 U3858 ( .B1(n4856), .B2(keyinput28), .C1(n2660), .C2(keyinput76), 
        .A(n3031), .ZN(n3035) );
  INV_X1 U3859 ( .A(REG2_REG_30__SCAN_IN), .ZN(n4728) );
  INV_X1 U3860 ( .A(REG2_REG_22__SCAN_IN), .ZN(n3033) );
  AOI22_X1 U3861 ( .A1(n4728), .A2(keyinput95), .B1(n3033), .B2(keyinput94), 
        .ZN(n3032) );
  OAI221_X1 U3862 ( .B1(n4728), .B2(keyinput95), .C1(n3033), .C2(keyinput94), 
        .A(n3032), .ZN(n3034) );
  NOR2_X1 U3863 ( .A1(n3035), .A2(n3034), .ZN(n3036) );
  NAND4_X1 U3864 ( .A1(n3039), .A2(n3038), .A3(n3037), .A4(n3036), .ZN(n3057)
         );
  INV_X1 U3865 ( .A(D_REG_10__SCAN_IN), .ZN(n4846) );
  XNOR2_X1 U3866 ( .A(n4846), .B(n2959), .ZN(n3055) );
  INV_X1 U3867 ( .A(D_REG_30__SCAN_IN), .ZN(n4834) );
  INV_X1 U3868 ( .A(keyinput123), .ZN(n3040) );
  XNOR2_X1 U3869 ( .A(n4834), .B(n3040), .ZN(n3054) );
  INV_X1 U3870 ( .A(D_REG_20__SCAN_IN), .ZN(n4838) );
  INV_X1 U3871 ( .A(keyinput125), .ZN(n3041) );
  XNOR2_X1 U3872 ( .A(n4838), .B(n3041), .ZN(n3053) );
  XNOR2_X1 U3873 ( .A(REG1_REG_0__SCAN_IN), .B(keyinput114), .ZN(n3045) );
  XNOR2_X1 U3874 ( .A(DATAI_2_), .B(keyinput122), .ZN(n3044) );
  XNOR2_X1 U3875 ( .A(REG1_REG_1__SCAN_IN), .B(keyinput90), .ZN(n3043) );
  XNOR2_X1 U3876 ( .A(IR_REG_3__SCAN_IN), .B(keyinput86), .ZN(n3042) );
  NAND4_X1 U3877 ( .A1(n3045), .A2(n3044), .A3(n3043), .A4(n3042), .ZN(n3051)
         );
  XNOR2_X1 U3878 ( .A(keyinput115), .B(REG1_REG_19__SCAN_IN), .ZN(n3049) );
  XNOR2_X1 U3879 ( .A(REG3_REG_2__SCAN_IN), .B(keyinput91), .ZN(n3048) );
  XNOR2_X1 U3880 ( .A(keyinput10), .B(DATAI_11_), .ZN(n3047) );
  XNOR2_X1 U3881 ( .A(keyinput16), .B(DATAI_7_), .ZN(n3046) );
  NAND4_X1 U3882 ( .A1(n3049), .A2(n3048), .A3(n3047), .A4(n3046), .ZN(n3050)
         );
  NOR2_X1 U3883 ( .A1(n3051), .A2(n3050), .ZN(n3052) );
  NAND4_X1 U3884 ( .A1(n3055), .A2(n3054), .A3(n3053), .A4(n3052), .ZN(n3056)
         );
  NOR2_X1 U3885 ( .A1(n3057), .A2(n3056), .ZN(n3127) );
  INV_X1 U3886 ( .A(REG3_REG_21__SCAN_IN), .ZN(n3798) );
  INV_X1 U3887 ( .A(REG0_REG_7__SCAN_IN), .ZN(n4901) );
  AOI22_X1 U3888 ( .A1(n3798), .A2(keyinput82), .B1(keyinput83), .B2(n4901), 
        .ZN(n3058) );
  OAI221_X1 U3889 ( .B1(n3798), .B2(keyinput82), .C1(n4901), .C2(keyinput83), 
        .A(n3058), .ZN(n3061) );
  INV_X1 U3890 ( .A(D_REG_19__SCAN_IN), .ZN(n4839) );
  INV_X1 U3891 ( .A(D_REG_5__SCAN_IN), .ZN(n4848) );
  AOI22_X1 U3892 ( .A1(n4839), .A2(keyinput119), .B1(keyinput118), .B2(n4848), 
        .ZN(n3059) );
  OAI221_X1 U3893 ( .B1(n4839), .B2(keyinput119), .C1(n4848), .C2(keyinput118), 
        .A(n3059), .ZN(n3060) );
  NOR2_X1 U3894 ( .A1(n3061), .A2(n3060), .ZN(n3069) );
  AOI22_X1 U3895 ( .A1(n3063), .A2(keyinput30), .B1(keyinput31), .B2(n2550), 
        .ZN(n3062) );
  OAI221_X1 U3896 ( .B1(n3063), .B2(keyinput30), .C1(n2550), .C2(keyinput31), 
        .A(n3062), .ZN(n3067) );
  INV_X1 U3897 ( .A(REG2_REG_3__SCAN_IN), .ZN(n3065) );
  AOI22_X1 U3898 ( .A1(n3065), .A2(keyinput22), .B1(keyinput23), .B2(n2484), 
        .ZN(n3064) );
  OAI221_X1 U3899 ( .B1(n3065), .B2(keyinput22), .C1(n2484), .C2(keyinput23), 
        .A(n3064), .ZN(n3066) );
  NOR2_X1 U3900 ( .A1(n3067), .A2(n3066), .ZN(n3068) );
  NAND2_X1 U3901 ( .A1(n3069), .A2(n3068), .ZN(n3080) );
  INV_X1 U3902 ( .A(D_REG_11__SCAN_IN), .ZN(n4845) );
  INV_X1 U3903 ( .A(D_REG_26__SCAN_IN), .ZN(n4836) );
  OAI22_X1 U3904 ( .A1(n4845), .A2(keyinput92), .B1(n4836), .B2(keyinput84), 
        .ZN(n3070) );
  AOI221_X1 U3905 ( .B1(n4845), .B2(keyinput92), .C1(keyinput84), .C2(n4836), 
        .A(n3070), .ZN(n3078) );
  INV_X1 U3906 ( .A(D_REG_17__SCAN_IN), .ZN(n4840) );
  INV_X1 U3907 ( .A(D_REG_14__SCAN_IN), .ZN(n4843) );
  OAI22_X1 U3908 ( .A1(n4840), .A2(keyinput48), .B1(n4843), .B2(keyinput52), 
        .ZN(n3071) );
  AOI221_X1 U3909 ( .B1(n4840), .B2(keyinput48), .C1(keyinput52), .C2(n4843), 
        .A(n3071), .ZN(n3077) );
  INV_X1 U3910 ( .A(D_REG_27__SCAN_IN), .ZN(n4835) );
  INV_X1 U3911 ( .A(D_REG_23__SCAN_IN), .ZN(n4837) );
  OAI22_X1 U3912 ( .A1(n4835), .A2(keyinput20), .B1(n4837), .B2(keyinput17), 
        .ZN(n3072) );
  AOI221_X1 U3913 ( .B1(n4835), .B2(keyinput20), .C1(keyinput17), .C2(n4837), 
        .A(n3072), .ZN(n3076) );
  INV_X1 U3914 ( .A(D_REG_1__SCAN_IN), .ZN(n3287) );
  INV_X1 U3915 ( .A(keyinput89), .ZN(n3074) );
  OAI22_X1 U3916 ( .A1(n3287), .A2(keyinput105), .B1(n3074), .B2(
        REG0_REG_31__SCAN_IN), .ZN(n3073) );
  AOI221_X1 U3917 ( .B1(n3287), .B2(keyinput105), .C1(REG0_REG_31__SCAN_IN), 
        .C2(n3074), .A(n3073), .ZN(n3075) );
  NAND4_X1 U3918 ( .A1(n3078), .A2(n3077), .A3(n3076), .A4(n3075), .ZN(n3079)
         );
  NOR2_X1 U3919 ( .A1(n3080), .A2(n3079), .ZN(n3126) );
  INV_X1 U3920 ( .A(REG1_REG_29__SCAN_IN), .ZN(n3082) );
  OAI22_X1 U3921 ( .A1(n3082), .A2(keyinput56), .B1(n4557), .B2(keyinput5), 
        .ZN(n3081) );
  AOI221_X1 U3922 ( .B1(n3082), .B2(keyinput56), .C1(keyinput5), .C2(n4557), 
        .A(n3081), .ZN(n3091) );
  OAI22_X1 U3923 ( .A1(n3085), .A2(keyinput113), .B1(n3084), .B2(keyinput4), 
        .ZN(n3083) );
  AOI221_X1 U3924 ( .B1(n3085), .B2(keyinput113), .C1(keyinput4), .C2(n3084), 
        .A(n3083), .ZN(n3090) );
  INV_X1 U3925 ( .A(REG0_REG_6__SCAN_IN), .ZN(n3626) );
  OAI22_X1 U3926 ( .A1(n3387), .A2(keyinput45), .B1(n3626), .B2(keyinput121), 
        .ZN(n3086) );
  AOI221_X1 U3927 ( .B1(n3387), .B2(keyinput45), .C1(keyinput121), .C2(n3626), 
        .A(n3086), .ZN(n3089) );
  INV_X1 U3928 ( .A(REG0_REG_2__SCAN_IN), .ZN(n4888) );
  OAI22_X1 U3929 ( .A1(n4888), .A2(keyinput88), .B1(n2516), .B2(keyinput73), 
        .ZN(n3087) );
  AOI221_X1 U3930 ( .B1(n4888), .B2(keyinput88), .C1(keyinput73), .C2(n2516), 
        .A(n3087), .ZN(n3088) );
  NAND4_X1 U3931 ( .A1(n3091), .A2(n3090), .A3(n3089), .A4(n3088), .ZN(n3124)
         );
  INV_X1 U3932 ( .A(DATAI_3_), .ZN(n3094) );
  INV_X1 U3933 ( .A(DATAI_6_), .ZN(n3093) );
  AOI22_X1 U3934 ( .A1(n3094), .A2(keyinput36), .B1(n3093), .B2(keyinput93), 
        .ZN(n3092) );
  OAI221_X1 U3935 ( .B1(n3094), .B2(keyinput36), .C1(n3093), .C2(keyinput93), 
        .A(n3092), .ZN(n3098) );
  INV_X1 U3936 ( .A(REG0_REG_16__SCAN_IN), .ZN(n3096) );
  AOI22_X1 U3937 ( .A1(n4602), .A2(keyinput60), .B1(n3096), .B2(keyinput25), 
        .ZN(n3095) );
  OAI221_X1 U3938 ( .B1(n4602), .B2(keyinput60), .C1(n3096), .C2(keyinput25), 
        .A(n3095), .ZN(n3097) );
  NOR2_X1 U3939 ( .A1(n3098), .A2(n3097), .ZN(n3122) );
  INV_X1 U3940 ( .A(DATAI_25_), .ZN(n3283) );
  INV_X1 U3941 ( .A(REG2_REG_21__SCAN_IN), .ZN(n3100) );
  AOI22_X1 U3942 ( .A1(n3283), .A2(keyinput126), .B1(keyinput127), .B2(n3100), 
        .ZN(n3099) );
  OAI221_X1 U3943 ( .B1(n3283), .B2(keyinput126), .C1(n3100), .C2(keyinput127), 
        .A(n3099), .ZN(n3103) );
  INV_X1 U3944 ( .A(keyinput2), .ZN(n3101) );
  XNOR2_X1 U3945 ( .A(n3101), .B(DATAO_REG_28__SCAN_IN), .ZN(n3102) );
  NOR2_X1 U3946 ( .A1(n3103), .A2(n3102), .ZN(n3121) );
  INV_X1 U3947 ( .A(keyinput7), .ZN(n3105) );
  INV_X1 U3948 ( .A(DATAO_REG_22__SCAN_IN), .ZN(n3104) );
  XNOR2_X1 U3949 ( .A(n3105), .B(n3104), .ZN(n3108) );
  INV_X1 U3950 ( .A(keyinput51), .ZN(n3106) );
  XNOR2_X1 U3951 ( .A(n3106), .B(n3295), .ZN(n3107) );
  AND2_X1 U3952 ( .A1(n3108), .A2(n3107), .ZN(n3120) );
  XNOR2_X1 U3953 ( .A(IR_REG_10__SCAN_IN), .B(keyinput61), .ZN(n3112) );
  XNOR2_X1 U3954 ( .A(IR_REG_22__SCAN_IN), .B(keyinput21), .ZN(n3111) );
  XNOR2_X1 U3955 ( .A(IR_REG_15__SCAN_IN), .B(keyinput11), .ZN(n3110) );
  XNOR2_X1 U3956 ( .A(DATAI_4_), .B(keyinput50), .ZN(n3109) );
  NAND4_X1 U3957 ( .A1(n3112), .A2(n3111), .A3(n3110), .A4(n3109), .ZN(n3118)
         );
  XNOR2_X1 U3958 ( .A(IR_REG_27__SCAN_IN), .B(keyinput3), .ZN(n3116) );
  XNOR2_X1 U3959 ( .A(DATAI_24_), .B(keyinput18), .ZN(n3115) );
  XNOR2_X1 U3960 ( .A(IR_REG_16__SCAN_IN), .B(keyinput6), .ZN(n3114) );
  XNOR2_X1 U3961 ( .A(IR_REG_21__SCAN_IN), .B(keyinput19), .ZN(n3113) );
  NAND4_X1 U3962 ( .A1(n3116), .A2(n3115), .A3(n3114), .A4(n3113), .ZN(n3117)
         );
  NOR2_X1 U3963 ( .A1(n3118), .A2(n3117), .ZN(n3119) );
  NAND4_X1 U3964 ( .A1(n3122), .A2(n3121), .A3(n3120), .A4(n3119), .ZN(n3123)
         );
  NOR2_X1 U3965 ( .A1(n3124), .A2(n3123), .ZN(n3125) );
  AND3_X1 U3966 ( .A1(n3127), .A2(n3126), .A3(n3125), .ZN(n3145) );
  INV_X1 U3967 ( .A(REG0_REG_29__SCAN_IN), .ZN(n3129) );
  AOI22_X1 U3968 ( .A1(n3129), .A2(keyinput75), .B1(keyinput74), .B2(n2237), 
        .ZN(n3128) );
  OAI221_X1 U3969 ( .B1(n3129), .B2(keyinput75), .C1(n2237), .C2(keyinput74), 
        .A(n3128), .ZN(n3138) );
  AOI22_X1 U3970 ( .A1(n3131), .A2(keyinput79), .B1(n2523), .B2(keyinput78), 
        .ZN(n3130) );
  OAI221_X1 U3971 ( .B1(n3131), .B2(keyinput79), .C1(n2523), .C2(keyinput78), 
        .A(n3130), .ZN(n3137) );
  INV_X1 U3972 ( .A(keyinput66), .ZN(n3133) );
  AOI22_X1 U3973 ( .A1(n2787), .A2(keyinput67), .B1(DATAO_REG_10__SCAN_IN), 
        .B2(n3133), .ZN(n3132) );
  OAI221_X1 U3974 ( .B1(n2787), .B2(keyinput67), .C1(n3133), .C2(
        DATAO_REG_10__SCAN_IN), .A(n3132), .ZN(n3136) );
  INV_X1 U3975 ( .A(D_REG_16__SCAN_IN), .ZN(n4841) );
  INV_X1 U3976 ( .A(REG3_REG_16__SCAN_IN), .ZN(n3826) );
  AOI22_X1 U3977 ( .A1(n4841), .A2(keyinput71), .B1(keyinput70), .B2(n3826), 
        .ZN(n3134) );
  OAI221_X1 U3978 ( .B1(n4841), .B2(keyinput71), .C1(n3826), .C2(keyinput70), 
        .A(n3134), .ZN(n3135) );
  NOR4_X1 U3979 ( .A1(n3138), .A2(n3137), .A3(n3136), .A4(n3135), .ZN(n3144)
         );
  INV_X1 U3980 ( .A(D_REG_3__SCAN_IN), .ZN(n4850) );
  INV_X1 U3981 ( .A(D_REG_2__SCAN_IN), .ZN(n4851) );
  OAI22_X1 U3982 ( .A1(n4850), .A2(keyinput65), .B1(n4851), .B2(keyinput104), 
        .ZN(n3139) );
  AOI221_X1 U3983 ( .B1(n4850), .B2(keyinput65), .C1(keyinput104), .C2(n4851), 
        .A(n3139), .ZN(n3143) );
  INV_X1 U3984 ( .A(IR_REG_12__SCAN_IN), .ZN(n3141) );
  OAI22_X1 U3985 ( .A1(n2585), .A2(keyinput69), .B1(n3141), .B2(keyinput0), 
        .ZN(n3140) );
  AOI221_X1 U3986 ( .B1(n2585), .B2(keyinput69), .C1(keyinput0), .C2(n3141), 
        .A(n3140), .ZN(n3142) );
  NAND4_X1 U3987 ( .A1(n3145), .A2(n3144), .A3(n3143), .A4(n3142), .ZN(n3228)
         );
  INV_X1 U3988 ( .A(REG0_REG_30__SCAN_IN), .ZN(n4647) );
  INV_X1 U3989 ( .A(keyinput33), .ZN(n3147) );
  AOI22_X1 U3990 ( .A1(n4647), .A2(keyinput77), .B1(DATAI_30_), .B2(n3147), 
        .ZN(n3146) );
  OAI221_X1 U3991 ( .B1(n4647), .B2(keyinput77), .C1(n3147), .C2(DATAI_30_), 
        .A(n3146), .ZN(n3159) );
  INV_X1 U3992 ( .A(keyinput32), .ZN(n3149) );
  AOI22_X1 U3993 ( .A1(n2567), .A2(keyinput64), .B1(ADDR_REG_0__SCAN_IN), .B2(
        n3149), .ZN(n3148) );
  OAI221_X1 U3994 ( .B1(n2567), .B2(keyinput64), .C1(n3149), .C2(
        ADDR_REG_0__SCAN_IN), .A(n3148), .ZN(n3158) );
  INV_X1 U3995 ( .A(keyinput8), .ZN(n3152) );
  INV_X1 U3996 ( .A(keyinput85), .ZN(n3151) );
  AOI22_X1 U3997 ( .A1(n3152), .A2(ADDR_REG_4__SCAN_IN), .B1(
        ADDR_REG_5__SCAN_IN), .B2(n3151), .ZN(n3150) );
  OAI221_X1 U3998 ( .B1(n3152), .B2(ADDR_REG_4__SCAN_IN), .C1(n3151), .C2(
        ADDR_REG_5__SCAN_IN), .A(n3150), .ZN(n3157) );
  INV_X1 U3999 ( .A(REG2_REG_8__SCAN_IN), .ZN(n3155) );
  INV_X1 U4000 ( .A(keyinput97), .ZN(n3154) );
  AOI22_X1 U4001 ( .A1(n3155), .A2(keyinput116), .B1(ADDR_REG_7__SCAN_IN), 
        .B2(n3154), .ZN(n3153) );
  OAI221_X1 U4002 ( .B1(n3155), .B2(keyinput116), .C1(n3154), .C2(
        ADDR_REG_7__SCAN_IN), .A(n3153), .ZN(n3156) );
  NOR4_X1 U4003 ( .A1(n3159), .A2(n3158), .A3(n3157), .A4(n3156), .ZN(n3173)
         );
  INV_X1 U4004 ( .A(REG0_REG_9__SCAN_IN), .ZN(n3162) );
  INV_X1 U4005 ( .A(keyinput43), .ZN(n3161) );
  AOI22_X1 U4006 ( .A1(n3162), .A2(keyinput42), .B1(DATAO_REG_21__SCAN_IN), 
        .B2(n3161), .ZN(n3160) );
  OAI221_X1 U4007 ( .B1(n3162), .B2(keyinput42), .C1(n3161), .C2(
        DATAO_REG_21__SCAN_IN), .A(n3160), .ZN(n3171) );
  INV_X1 U4008 ( .A(REG3_REG_26__SCAN_IN), .ZN(n3908) );
  AOI22_X1 U4009 ( .A1(n3908), .A2(keyinput46), .B1(keyinput47), .B2(n4528), 
        .ZN(n3163) );
  OAI221_X1 U4010 ( .B1(n3908), .B2(keyinput46), .C1(n4528), .C2(keyinput47), 
        .A(n3163), .ZN(n3170) );
  INV_X1 U4011 ( .A(REG0_REG_10__SCAN_IN), .ZN(n4909) );
  INV_X1 U4012 ( .A(keyinput35), .ZN(n3165) );
  AOI22_X1 U4013 ( .A1(n4909), .A2(keyinput34), .B1(DATAO_REG_6__SCAN_IN), 
        .B2(n3165), .ZN(n3164) );
  OAI221_X1 U4014 ( .B1(n4909), .B2(keyinput34), .C1(n3165), .C2(
        DATAO_REG_6__SCAN_IN), .A(n3164), .ZN(n3169) );
  INV_X1 U4015 ( .A(REG0_REG_13__SCAN_IN), .ZN(n3167) );
  INV_X1 U4016 ( .A(D_REG_4__SCAN_IN), .ZN(n4849) );
  AOI22_X1 U4017 ( .A1(n3167), .A2(keyinput39), .B1(n4849), .B2(keyinput38), 
        .ZN(n3166) );
  OAI221_X1 U4018 ( .B1(n3167), .B2(keyinput39), .C1(n4849), .C2(keyinput38), 
        .A(n3166), .ZN(n3168) );
  NOR4_X1 U4019 ( .A1(n3171), .A2(n3170), .A3(n3169), .A4(n3168), .ZN(n3172)
         );
  NAND2_X1 U4020 ( .A1(n3173), .A2(n3172), .ZN(n3227) );
  INV_X1 U4021 ( .A(keyinput29), .ZN(n3176) );
  INV_X1 U4022 ( .A(keyinput117), .ZN(n3175) );
  AOI22_X1 U4023 ( .A1(n3176), .A2(ADDR_REG_8__SCAN_IN), .B1(
        ADDR_REG_9__SCAN_IN), .B2(n3175), .ZN(n3174) );
  OAI221_X1 U4024 ( .B1(n3176), .B2(ADDR_REG_8__SCAN_IN), .C1(n3175), .C2(
        ADDR_REG_9__SCAN_IN), .A(n3174), .ZN(n3187) );
  INV_X1 U4025 ( .A(REG2_REG_10__SCAN_IN), .ZN(n3179) );
  INV_X1 U4026 ( .A(REG2_REG_12__SCAN_IN), .ZN(n3178) );
  AOI22_X1 U4027 ( .A1(n3179), .A2(keyinput81), .B1(keyinput120), .B2(n3178), 
        .ZN(n3177) );
  OAI221_X1 U4028 ( .B1(n3179), .B2(keyinput81), .C1(n3178), .C2(keyinput120), 
        .A(n3177), .ZN(n3186) );
  INV_X1 U4029 ( .A(keyinput72), .ZN(n3182) );
  INV_X1 U4030 ( .A(keyinput112), .ZN(n3181) );
  AOI22_X1 U4031 ( .A1(n3182), .A2(ADDR_REG_14__SCAN_IN), .B1(
        ADDR_REG_17__SCAN_IN), .B2(n3181), .ZN(n3180) );
  OAI221_X1 U4032 ( .B1(n3182), .B2(ADDR_REG_14__SCAN_IN), .C1(n3181), .C2(
        ADDR_REG_17__SCAN_IN), .A(n3180), .ZN(n3185) );
  INV_X1 U4033 ( .A(REG1_REG_13__SCAN_IN), .ZN(n4142) );
  AOI22_X1 U4034 ( .A1(n4142), .A2(keyinput108), .B1(keyinput100), .B2(n3385), 
        .ZN(n3183) );
  OAI221_X1 U4035 ( .B1(n4142), .B2(keyinput108), .C1(n3385), .C2(keyinput100), 
        .A(n3183), .ZN(n3184) );
  NOR4_X1 U4036 ( .A1(n3187), .A2(n3186), .A3(n3185), .A4(n3184), .ZN(n3225)
         );
  INV_X1 U4037 ( .A(keyinput96), .ZN(n3189) );
  AOI22_X1 U4038 ( .A1(n2447), .A2(keyinput12), .B1(ADDR_REG_19__SCAN_IN), 
        .B2(n3189), .ZN(n3188) );
  OAI221_X1 U4039 ( .B1(n2447), .B2(keyinput12), .C1(n3189), .C2(
        ADDR_REG_19__SCAN_IN), .A(n3188), .ZN(n3199) );
  INV_X1 U4040 ( .A(keyinput1), .ZN(n3192) );
  INV_X1 U4041 ( .A(keyinput49), .ZN(n3191) );
  AOI22_X1 U4042 ( .A1(n3192), .A2(DATAO_REG_12__SCAN_IN), .B1(
        DATAO_REG_3__SCAN_IN), .B2(n3191), .ZN(n3190) );
  OAI221_X1 U40430 ( .B1(n3192), .B2(DATAO_REG_12__SCAN_IN), .C1(n3191), .C2(
        DATAO_REG_3__SCAN_IN), .A(n3190), .ZN(n3198) );
  INV_X1 U4044 ( .A(keyinput13), .ZN(n3194) );
  AOI22_X1 U4045 ( .A1(n3846), .A2(keyinput9), .B1(DATAO_REG_15__SCAN_IN), 
        .B2(n3194), .ZN(n3193) );
  OAI221_X1 U4046 ( .B1(n3846), .B2(keyinput9), .C1(n3194), .C2(
        DATAO_REG_15__SCAN_IN), .A(n3193), .ZN(n3197) );
  INV_X1 U4047 ( .A(REG2_REG_20__SCAN_IN), .ZN(n4338) );
  INV_X1 U4048 ( .A(REG2_REG_16__SCAN_IN), .ZN(n4800) );
  AOI22_X1 U4049 ( .A1(n4338), .A2(keyinput24), .B1(keyinput124), .B2(n4800), 
        .ZN(n3195) );
  OAI221_X1 U4050 ( .B1(n4338), .B2(keyinput24), .C1(n4800), .C2(keyinput124), 
        .A(n3195), .ZN(n3196) );
  NOR4_X1 U4051 ( .A1(n3199), .A2(n3198), .A3(n3197), .A4(n3196), .ZN(n3224)
         );
  INV_X1 U4052 ( .A(REG2_REG_17__SCAN_IN), .ZN(n4153) );
  AOI22_X1 U4053 ( .A1(n3366), .A2(keyinput57), .B1(n4153), .B2(keyinput80), 
        .ZN(n3200) );
  OAI221_X1 U4054 ( .B1(n3366), .B2(keyinput57), .C1(n4153), .C2(keyinput80), 
        .A(n3200), .ZN(n3211) );
  INV_X1 U4055 ( .A(REG2_REG_5__SCAN_IN), .ZN(n4132) );
  INV_X1 U4056 ( .A(REG2_REG_9__SCAN_IN), .ZN(n3643) );
  AOI22_X1 U4057 ( .A1(n4132), .A2(keyinput109), .B1(n3643), .B2(keyinput41), 
        .ZN(n3201) );
  OAI221_X1 U4058 ( .B1(n4132), .B2(keyinput109), .C1(n3643), .C2(keyinput41), 
        .A(n3201), .ZN(n3210) );
  INV_X1 U4059 ( .A(keyinput53), .ZN(n3204) );
  INV_X1 U4060 ( .A(keyinput68), .ZN(n3203) );
  AOI22_X1 U4061 ( .A1(n3204), .A2(DATAO_REG_20__SCAN_IN), .B1(
        DATAO_REG_26__SCAN_IN), .B2(n3203), .ZN(n3202) );
  OAI221_X1 U4062 ( .B1(n3204), .B2(DATAO_REG_20__SCAN_IN), .C1(n3203), .C2(
        DATAO_REG_26__SCAN_IN), .A(n3202), .ZN(n3209) );
  INV_X1 U4063 ( .A(keyinput101), .ZN(n3207) );
  INV_X1 U4064 ( .A(keyinput37), .ZN(n3206) );
  AOI22_X1 U4065 ( .A1(n3207), .A2(DATAO_REG_27__SCAN_IN), .B1(
        DATAO_REG_31__SCAN_IN), .B2(n3206), .ZN(n3205) );
  OAI221_X1 U4066 ( .B1(n3207), .B2(DATAO_REG_27__SCAN_IN), .C1(n3206), .C2(
        DATAO_REG_31__SCAN_IN), .A(n3205), .ZN(n3208) );
  NOR4_X1 U4067 ( .A1(n3211), .A2(n3210), .A3(n3209), .A4(n3208), .ZN(n3223)
         );
  INV_X1 U4068 ( .A(DATAI_1_), .ZN(n3213) );
  AOI22_X1 U4069 ( .A1(n3213), .A2(keyinput106), .B1(n3809), .B2(keyinput107), 
        .ZN(n3212) );
  OAI221_X1 U4070 ( .B1(n3213), .B2(keyinput106), .C1(n3809), .C2(keyinput107), 
        .A(n3212), .ZN(n3221) );
  INV_X1 U4071 ( .A(DATAI_23_), .ZN(n4854) );
  AOI22_X1 U4072 ( .A1(n3734), .A2(keyinput111), .B1(keyinput110), .B2(n4854), 
        .ZN(n3214) );
  OAI221_X1 U4073 ( .B1(n3734), .B2(keyinput111), .C1(n4854), .C2(keyinput110), 
        .A(n3214), .ZN(n3220) );
  AOI22_X1 U4074 ( .A1(n3818), .A2(keyinput98), .B1(n2345), .B2(keyinput99), 
        .ZN(n3215) );
  OAI221_X1 U4075 ( .B1(n3818), .B2(keyinput98), .C1(n2345), .C2(keyinput99), 
        .A(n3215), .ZN(n3219) );
  INV_X1 U4076 ( .A(DATAI_28_), .ZN(n4721) );
  INV_X1 U4077 ( .A(keyinput102), .ZN(n3217) );
  AOI22_X1 U4078 ( .A1(n4721), .A2(keyinput103), .B1(ADDR_REG_2__SCAN_IN), 
        .B2(n3217), .ZN(n3216) );
  OAI221_X1 U4079 ( .B1(n4721), .B2(keyinput103), .C1(n3217), .C2(
        ADDR_REG_2__SCAN_IN), .A(n3216), .ZN(n3218) );
  NOR4_X1 U4080 ( .A1(n3221), .A2(n3220), .A3(n3219), .A4(n3218), .ZN(n3222)
         );
  NAND4_X1 U4081 ( .A1(n3225), .A2(n3224), .A3(n3223), .A4(n3222), .ZN(n3226)
         );
  NOR3_X1 U4082 ( .A1(n3228), .A2(n3227), .A3(n3226), .ZN(n3229) );
  OAI21_X1 U4083 ( .B1(n3231), .B2(n3230), .A(n3229), .ZN(n3232) );
  NOR2_X1 U4084 ( .A1(n4513), .A2(n3233), .ZN(n3234) );
  NAND2_X1 U4085 ( .A1(n3929), .A2(DATAI_29_), .ZN(n3932) );
  XNOR2_X1 U4086 ( .A(n4085), .B(n3932), .ZN(n3994) );
  XNOR2_X1 U4087 ( .A(n3236), .B(n3994), .ZN(n4191) );
  INV_X1 U4088 ( .A(n3954), .ZN(n3931) );
  AOI21_X1 U4089 ( .B1(n3237), .B2(n3933), .A(n3931), .ZN(n3238) );
  XNOR2_X1 U4090 ( .A(n3238), .B(n3994), .ZN(n3239) );
  NAND2_X1 U4091 ( .A1(n3239), .A2(n4491), .ZN(n3245) );
  INV_X1 U4092 ( .A(REG1_REG_30__SCAN_IN), .ZN(n3242) );
  NAND2_X1 U4093 ( .A1(n3302), .A2(REG2_REG_30__SCAN_IN), .ZN(n3241) );
  NAND2_X1 U4094 ( .A1(n2429), .A2(REG0_REG_30__SCAN_IN), .ZN(n3240) );
  OAI211_X1 U4095 ( .C1(n3305), .C2(n3242), .A(n3241), .B(n3240), .ZN(n4084)
         );
  XNOR2_X1 U4096 ( .A(n3243), .B(IR_REG_27__SCAN_IN), .ZN(n4709) );
  AOI21_X1 U4097 ( .B1(n4709), .B2(B_REG_SCAN_IN), .A(n4878), .ZN(n4186) );
  INV_X1 U4098 ( .A(n3932), .ZN(n3938) );
  AOI22_X1 U4099 ( .A1(n4084), .A2(n4186), .B1(n3938), .B2(n4627), .ZN(n3244)
         );
  OAI211_X1 U4100 ( .C1(n4513), .C2(n4615), .A(n3245), .B(n3244), .ZN(n4195)
         );
  AOI21_X1 U4101 ( .B1(n4191), .B2(n4895), .A(n4195), .ZN(n3256) );
  INV_X1 U4102 ( .A(n4910), .ZN(n3250) );
  OAI21_X1 U4103 ( .B1(n3246), .B2(n3932), .A(n4502), .ZN(n4193) );
  OR2_X1 U4104 ( .A1(n4193), .A2(n4706), .ZN(n3248) );
  NAND2_X1 U4105 ( .A1(n3250), .A2(REG0_REG_29__SCAN_IN), .ZN(n3247) );
  INV_X1 U4106 ( .A(n4853), .ZN(n3257) );
  INV_X1 U4107 ( .A(n3259), .ZN(n3260) );
  AOI211_X1 U4108 ( .C1(n3261), .C2(n3258), .A(n3898), .B(n3260), .ZN(n3266)
         );
  NOR2_X1 U4109 ( .A1(n3928), .A2(n3557), .ZN(n3265) );
  NAND2_X1 U4110 ( .A1(REG3_REG_4__SCAN_IN), .A2(U3149), .ZN(n3408) );
  OAI21_X1 U4111 ( .B1(n2859), .B2(n3923), .A(n3408), .ZN(n3264) );
  INV_X1 U4112 ( .A(n3921), .ZN(n3466) );
  NAND2_X1 U4113 ( .A1(n3466), .A2(n3551), .ZN(n3262) );
  OAI21_X1 U4114 ( .B1(n3920), .B2(n3555), .A(n3262), .ZN(n3263) );
  OR4_X1 U4115 ( .A1(n3266), .A2(n3265), .A3(n3264), .A4(n3263), .ZN(U3227) );
  INV_X1 U4116 ( .A(n3268), .ZN(n3269) );
  AOI211_X1 U4117 ( .C1(n3270), .C2(n3267), .A(n3898), .B(n3269), .ZN(n3275)
         );
  NOR2_X1 U4118 ( .A1(n3928), .A2(n3728), .ZN(n3274) );
  NAND2_X1 U4119 ( .A1(REG3_REG_10__SCAN_IN), .A2(U3149), .ZN(n4752) );
  OAI21_X1 U4120 ( .B1(n4616), .B2(n3923), .A(n4752), .ZN(n3273) );
  NAND2_X1 U4121 ( .A1(n3466), .A2(n4086), .ZN(n3271) );
  OAI21_X1 U4122 ( .B1(n3920), .B2(n3726), .A(n3271), .ZN(n3272) );
  OR4_X1 U4123 ( .A1(n3275), .A2(n3274), .A3(n3273), .A4(n3272), .ZN(U3214) );
  MUX2_X1 U4124 ( .A(n2484), .B(n4131), .S(STATE_REG_SCAN_IN), .Z(n3276) );
  INV_X1 U4125 ( .A(n3276), .ZN(U3347) );
  INV_X1 U4126 ( .A(n4141), .ZN(n4155) );
  NAND2_X1 U4127 ( .A1(n4155), .A2(STATE_REG_SCAN_IN), .ZN(n3277) );
  OAI21_X1 U4128 ( .B1(STATE_REG_SCAN_IN), .B2(n2606), .A(n3277), .ZN(U3339)
         );
  MUX2_X1 U4129 ( .A(n2681), .B(n4179), .S(STATE_REG_SCAN_IN), .Z(n3278) );
  INV_X1 U4130 ( .A(n3278), .ZN(U3333) );
  INV_X1 U4131 ( .A(DATAI_21_), .ZN(n3280) );
  NAND2_X1 U4132 ( .A1(n4005), .A2(STATE_REG_SCAN_IN), .ZN(n3279) );
  OAI21_X1 U4133 ( .B1(STATE_REG_SCAN_IN), .B2(n3280), .A(n3279), .ZN(U3331)
         );
  NAND2_X1 U4134 ( .A1(n3281), .A2(STATE_REG_SCAN_IN), .ZN(n3282) );
  OAI21_X1 U4135 ( .B1(STATE_REG_SCAN_IN), .B2(n3283), .A(n3282), .ZN(U3327)
         );
  INV_X1 U4136 ( .A(n3285), .ZN(n3286) );
  AOI22_X1 U4137 ( .A1(n4847), .A2(n3287), .B1(n3286), .B2(n4853), .ZN(U3459)
         );
  AOI22_X1 U4138 ( .A1(n4847), .A2(n3289), .B1(n3288), .B2(n4853), .ZN(U3458)
         );
  INV_X1 U4139 ( .A(DATAI_30_), .ZN(n3292) );
  NAND2_X1 U4140 ( .A1(n3290), .A2(STATE_REG_SCAN_IN), .ZN(n3291) );
  OAI21_X1 U4141 ( .B1(STATE_REG_SCAN_IN), .B2(n3292), .A(n3291), .ZN(U3322)
         );
  INV_X1 U4142 ( .A(DATAI_31_), .ZN(n3295) );
  OR4_X1 U4143 ( .A1(n2238), .A2(IR_REG_30__SCAN_IN), .A3(n3293), .A4(U3149), 
        .ZN(n3294) );
  OAI21_X1 U4144 ( .B1(STATE_REG_SCAN_IN), .B2(n3295), .A(n3294), .ZN(U3321)
         );
  INV_X1 U4145 ( .A(n3296), .ZN(n3298) );
  INV_X1 U4146 ( .A(n3300), .ZN(n3297) );
  NAND2_X1 U4147 ( .A1(n3297), .A2(STATE_REG_SCAN_IN), .ZN(n4082) );
  NAND2_X1 U4148 ( .A1(n3298), .A2(n4082), .ZN(n3338) );
  NAND2_X1 U4149 ( .A1(n3300), .A2(n3299), .ZN(n3301) );
  NAND2_X1 U4150 ( .A1(n3929), .A2(n3301), .ZN(n3336) );
  NOR2_X1 U4151 ( .A1(n4815), .A2(U4043), .ZN(U3148) );
  INV_X1 U4152 ( .A(DATAO_REG_31__SCAN_IN), .ZN(n3307) );
  INV_X1 U4153 ( .A(REG1_REG_31__SCAN_IN), .ZN(n4498) );
  NAND2_X1 U4154 ( .A1(n2429), .A2(REG0_REG_31__SCAN_IN), .ZN(n3304) );
  NAND2_X1 U4155 ( .A1(n3302), .A2(REG2_REG_31__SCAN_IN), .ZN(n3303) );
  OAI211_X1 U4156 ( .C1(n3305), .C2(n4498), .A(n3304), .B(n3303), .ZN(n4187)
         );
  NAND2_X1 U4157 ( .A1(n4187), .A2(n2181), .ZN(n3306) );
  OAI21_X1 U4158 ( .B1(U4043), .B2(n3307), .A(n3306), .ZN(U3581) );
  INV_X1 U4159 ( .A(DATAO_REG_20__SCAN_IN), .ZN(n3309) );
  NAND2_X1 U4160 ( .A1(n4354), .A2(U4043), .ZN(n3308) );
  OAI21_X1 U4161 ( .B1(n2181), .B2(n3309), .A(n3308), .ZN(U3570) );
  INV_X1 U4162 ( .A(DATAO_REG_10__SCAN_IN), .ZN(n3311) );
  NAND2_X1 U4163 ( .A1(n4629), .A2(n2181), .ZN(n3310) );
  OAI21_X1 U4164 ( .B1(U4043), .B2(n3311), .A(n3310), .ZN(U3560) );
  INV_X1 U4165 ( .A(DATAO_REG_3__SCAN_IN), .ZN(n3313) );
  NAND2_X1 U4166 ( .A1(n3551), .A2(n2181), .ZN(n3312) );
  OAI21_X1 U4167 ( .B1(U4043), .B2(n3313), .A(n3312), .ZN(U3553) );
  INV_X1 U4168 ( .A(DATAO_REG_6__SCAN_IN), .ZN(n3315) );
  NAND2_X1 U4169 ( .A1(n3676), .A2(n2181), .ZN(n3314) );
  OAI21_X1 U4170 ( .B1(n2181), .B2(n3315), .A(n3314), .ZN(U3556) );
  NAND2_X1 U4171 ( .A1(n4551), .A2(n2181), .ZN(n3316) );
  OAI21_X1 U4172 ( .B1(n2181), .B2(n3104), .A(n3316), .ZN(U3572) );
  INV_X1 U4173 ( .A(DATAO_REG_21__SCAN_IN), .ZN(n3318) );
  NAND2_X1 U4174 ( .A1(n4327), .A2(U4043), .ZN(n3317) );
  OAI21_X1 U4175 ( .B1(n2181), .B2(n3318), .A(n3317), .ZN(U3571) );
  INV_X1 U4176 ( .A(DATAO_REG_26__SCAN_IN), .ZN(n3320) );
  NAND2_X1 U4177 ( .A1(n4510), .A2(n2181), .ZN(n3319) );
  OAI21_X1 U4178 ( .B1(n2181), .B2(n3320), .A(n3319), .ZN(U3576) );
  INV_X1 U4179 ( .A(DATAO_REG_11__SCAN_IN), .ZN(n3322) );
  NAND2_X1 U4180 ( .A1(n3719), .A2(n2181), .ZN(n3321) );
  OAI21_X1 U4181 ( .B1(n2181), .B2(n3322), .A(n3321), .ZN(U3561) );
  INV_X1 U4182 ( .A(DATAO_REG_8__SCAN_IN), .ZN(n3324) );
  NAND2_X1 U4183 ( .A1(n3667), .A2(n2181), .ZN(n3323) );
  OAI21_X1 U4184 ( .B1(n2181), .B2(n3324), .A(n3323), .ZN(U3558) );
  INV_X1 U4185 ( .A(DATAO_REG_13__SCAN_IN), .ZN(n3326) );
  NAND2_X1 U4186 ( .A1(n4481), .A2(U4043), .ZN(n3325) );
  OAI21_X1 U4187 ( .B1(n2181), .B2(n3326), .A(n3325), .ZN(U3563) );
  INV_X1 U4188 ( .A(DATAO_REG_27__SCAN_IN), .ZN(n3328) );
  NAND2_X1 U4189 ( .A1(n4520), .A2(n2181), .ZN(n3327) );
  OAI21_X1 U4190 ( .B1(n2181), .B2(n3328), .A(n3327), .ZN(U3577) );
  INV_X1 U4191 ( .A(DATAO_REG_12__SCAN_IN), .ZN(n3330) );
  NAND2_X1 U4192 ( .A1(n4607), .A2(n2181), .ZN(n3329) );
  OAI21_X1 U4193 ( .B1(n2181), .B2(n3330), .A(n3329), .ZN(U3562) );
  INV_X1 U4194 ( .A(DATAO_REG_15__SCAN_IN), .ZN(n3332) );
  NAND2_X1 U4195 ( .A1(n4404), .A2(n2181), .ZN(n3331) );
  OAI21_X1 U4196 ( .B1(n2181), .B2(n3332), .A(n3331), .ZN(U3565) );
  INV_X1 U4197 ( .A(REG2_REG_2__SCAN_IN), .ZN(n3526) );
  INV_X1 U4198 ( .A(REG2_REG_1__SCAN_IN), .ZN(n3333) );
  MUX2_X1 U4199 ( .A(REG2_REG_1__SCAN_IN), .B(n3333), .S(n4720), .Z(n4105) );
  AND2_X1 U4200 ( .A1(IR_REG_0__SCAN_IN), .A2(REG2_REG_0__SCAN_IN), .ZN(n4106)
         );
  NAND2_X1 U4201 ( .A1(n4105), .A2(n4106), .ZN(n4104) );
  NAND2_X1 U4202 ( .A1(n4720), .A2(REG2_REG_1__SCAN_IN), .ZN(n3334) );
  NAND2_X1 U4203 ( .A1(n4104), .A2(n3334), .ZN(n4117) );
  NAND2_X1 U4204 ( .A1(n4719), .A2(REG2_REG_2__SCAN_IN), .ZN(n3335) );
  INV_X1 U4205 ( .A(n4718), .ZN(n3343) );
  XNOR2_X1 U4206 ( .A(n3352), .B(n3343), .ZN(n3351) );
  XNOR2_X1 U4207 ( .A(n3351), .B(REG2_REG_3__SCAN_IN), .ZN(n3347) );
  INV_X1 U4208 ( .A(n3336), .ZN(n3337) );
  NOR2_X1 U4209 ( .A1(n4722), .A2(n4093), .ZN(n4079) );
  INV_X1 U4210 ( .A(REG3_REG_3__SCAN_IN), .ZN(n3536) );
  NOR2_X1 U4211 ( .A1(STATE_REG_SCAN_IN), .A2(n3536), .ZN(n3476) );
  NOR2_X1 U4212 ( .A1(n4822), .A2(n3343), .ZN(n3339) );
  AOI211_X1 U4213 ( .C1(n4815), .C2(ADDR_REG_3__SCAN_IN), .A(n3476), .B(n3339), 
        .ZN(n3346) );
  INV_X1 U4214 ( .A(REG1_REG_2__SCAN_IN), .ZN(n4915) );
  MUX2_X1 U4215 ( .A(REG1_REG_2__SCAN_IN), .B(n4915), .S(n4719), .Z(n4121) );
  XNOR2_X1 U4216 ( .A(n4720), .B(n3340), .ZN(n4103) );
  AND2_X1 U4217 ( .A1(IR_REG_0__SCAN_IN), .A2(REG1_REG_0__SCAN_IN), .ZN(n4102)
         );
  NAND2_X1 U4218 ( .A1(n4103), .A2(n4102), .ZN(n4101) );
  NAND2_X1 U4219 ( .A1(n4720), .A2(REG1_REG_1__SCAN_IN), .ZN(n3341) );
  NAND2_X1 U4220 ( .A1(n4101), .A2(n3341), .ZN(n4120) );
  NAND2_X1 U4221 ( .A1(n4121), .A2(n4120), .ZN(n4119) );
  NAND2_X1 U4222 ( .A1(n4719), .A2(REG1_REG_2__SCAN_IN), .ZN(n3342) );
  NAND2_X1 U4223 ( .A1(n4119), .A2(n3342), .ZN(n3362) );
  NAND2_X1 U4224 ( .A1(n3344), .A2(REG1_REG_3__SCAN_IN), .ZN(n3364) );
  OAI211_X1 U4225 ( .C1(REG1_REG_3__SCAN_IN), .C2(n3344), .A(n4816), .B(n3364), 
        .ZN(n3345) );
  OAI211_X1 U4226 ( .C1(n3347), .C2(n4809), .A(n3346), .B(n3345), .ZN(U3243)
         );
  INV_X1 U4227 ( .A(DATAO_REG_28__SCAN_IN), .ZN(n3350) );
  NAND2_X1 U4228 ( .A1(n3348), .A2(n2181), .ZN(n3349) );
  OAI21_X1 U4229 ( .B1(n2181), .B2(n3350), .A(n3349), .ZN(U3578) );
  NAND2_X1 U4230 ( .A1(n3351), .A2(REG2_REG_3__SCAN_IN), .ZN(n3354) );
  NAND2_X1 U4231 ( .A1(n3352), .A2(n4718), .ZN(n3353) );
  INV_X1 U4232 ( .A(REG2_REG_4__SCAN_IN), .ZN(n3355) );
  NAND2_X1 U4233 ( .A1(n3356), .A2(n4717), .ZN(n3357) );
  MUX2_X1 U4234 ( .A(n4132), .B(REG2_REG_5__SCAN_IN), .S(n4131), .Z(n3358) );
  NAND2_X1 U4235 ( .A1(n4135), .A2(n3358), .ZN(n4134) );
  OR2_X1 U4236 ( .A1(n4131), .A2(n4132), .ZN(n3359) );
  NAND2_X1 U4237 ( .A1(n4134), .A2(n3359), .ZN(n3391) );
  INV_X1 U4238 ( .A(n4716), .ZN(n3361) );
  XNOR2_X1 U4239 ( .A(n3391), .B(n3361), .ZN(n3393) );
  XOR2_X1 U4240 ( .A(REG2_REG_6__SCAN_IN), .B(n3393), .Z(n3370) );
  AND2_X1 U4241 ( .A1(U3149), .A2(REG3_REG_6__SCAN_IN), .ZN(n3636) );
  AOI21_X1 U4242 ( .B1(n4815), .B2(ADDR_REG_6__SCAN_IN), .A(n3636), .ZN(n3360)
         );
  OAI21_X1 U4243 ( .B1(n4822), .B2(n3361), .A(n3360), .ZN(n3369) );
  NAND2_X1 U4244 ( .A1(n3362), .A2(n4718), .ZN(n3363) );
  NAND2_X1 U4245 ( .A1(n3364), .A2(n3363), .ZN(n3365) );
  INV_X1 U4246 ( .A(n4717), .ZN(n3412) );
  XNOR2_X1 U4247 ( .A(n3365), .B(n3412), .ZN(n3407) );
  NAND2_X1 U4248 ( .A1(n3407), .A2(REG1_REG_4__SCAN_IN), .ZN(n3406) );
  MUX2_X1 U4249 ( .A(n3366), .B(REG1_REG_5__SCAN_IN), .S(n4131), .Z(n4130) );
  NOR2_X1 U4250 ( .A1(n3367), .A2(n2491), .ZN(n3383) );
  INV_X1 U4251 ( .A(n4816), .ZN(n4184) );
  AOI211_X1 U4252 ( .C1(n2491), .C2(n3367), .A(n3383), .B(n4184), .ZN(n3368)
         );
  AOI211_X1 U4253 ( .C1(n4773), .C2(n3370), .A(n3369), .B(n3368), .ZN(n3371)
         );
  INV_X1 U4254 ( .A(n3371), .ZN(U3246) );
  OAI21_X1 U4255 ( .B1(n3374), .B2(n3373), .A(n3372), .ZN(n3400) );
  INV_X1 U4256 ( .A(n3923), .ZN(n3906) );
  AOI22_X1 U4257 ( .A1(n3906), .A2(n3375), .B1(n3465), .B2(n3376), .ZN(n3382)
         );
  INV_X1 U4258 ( .A(n3377), .ZN(n3380) );
  INV_X1 U4259 ( .A(n3378), .ZN(n3421) );
  NAND3_X1 U4260 ( .A1(n3380), .A2(n3421), .A3(n3379), .ZN(n3469) );
  INV_X1 U4261 ( .A(n3469), .ZN(n3459) );
  OR2_X1 U4262 ( .A1(n3459), .A2(n3427), .ZN(n3381) );
  OAI211_X1 U4263 ( .C1(n3400), .C2(n3898), .A(n3382), .B(n3381), .ZN(U3229)
         );
  AOI21_X1 U4264 ( .B1(n4716), .B2(n3384), .A(n3383), .ZN(n3562) );
  MUX2_X1 U4265 ( .A(n3385), .B(REG1_REG_7__SCAN_IN), .S(n4715), .Z(n3386) );
  XNOR2_X1 U4266 ( .A(n3562), .B(n3386), .ZN(n3399) );
  INV_X1 U4267 ( .A(n4822), .ZN(n4170) );
  INV_X1 U4268 ( .A(n4815), .ZN(n3390) );
  INV_X1 U4269 ( .A(ADDR_REG_7__SCAN_IN), .ZN(n3389) );
  NOR2_X1 U4270 ( .A1(STATE_REG_SCAN_IN), .A2(n3387), .ZN(n3666) );
  INV_X1 U4271 ( .A(n3666), .ZN(n3388) );
  OAI21_X1 U4272 ( .B1(n3390), .B2(n3389), .A(n3388), .ZN(n3397) );
  AND2_X1 U4273 ( .A1(n3391), .A2(n4716), .ZN(n3392) );
  AOI21_X1 U4274 ( .B1(n3393), .B2(REG2_REG_6__SCAN_IN), .A(n3392), .ZN(n3395)
         );
  INV_X1 U4275 ( .A(REG2_REG_7__SCAN_IN), .ZN(n3679) );
  MUX2_X1 U4276 ( .A(n3679), .B(REG2_REG_7__SCAN_IN), .S(n4715), .Z(n3394) );
  AOI211_X1 U4277 ( .C1(n3395), .C2(n3394), .A(n3579), .B(n4809), .ZN(n3396)
         );
  AOI211_X1 U4278 ( .C1(n4170), .C2(n4715), .A(n3397), .B(n3396), .ZN(n3398)
         );
  OAI21_X1 U4279 ( .B1(n3399), .B2(n4184), .A(n3398), .ZN(U3247) );
  NAND3_X1 U4280 ( .A1(n3400), .A2(n3402), .A3(n4093), .ZN(n3404) );
  INV_X1 U4281 ( .A(REG2_REG_0__SCAN_IN), .ZN(n3428) );
  NAND2_X1 U4282 ( .A1(n4709), .A2(n3428), .ZN(n3401) );
  NAND2_X1 U4283 ( .A1(n3402), .A2(n3401), .ZN(n4097) );
  NAND2_X1 U4284 ( .A1(n4097), .A2(n2225), .ZN(n4095) );
  NAND2_X1 U4285 ( .A1(n4079), .A2(n4106), .ZN(n3403) );
  NAND4_X1 U4286 ( .A1(n3404), .A2(n2181), .A3(n4095), .A4(n3403), .ZN(n4125)
         );
  XNOR2_X1 U4287 ( .A(n3405), .B(REG2_REG_4__SCAN_IN), .ZN(n3414) );
  OAI211_X1 U4288 ( .C1(REG1_REG_4__SCAN_IN), .C2(n3407), .A(n4816), .B(n3406), 
        .ZN(n3411) );
  INV_X1 U4289 ( .A(n3408), .ZN(n3409) );
  AOI21_X1 U4290 ( .B1(n4815), .B2(ADDR_REG_4__SCAN_IN), .A(n3409), .ZN(n3410)
         );
  OAI211_X1 U4291 ( .C1(n4822), .C2(n3412), .A(n3411), .B(n3410), .ZN(n3413)
         );
  AOI21_X1 U4292 ( .B1(n4773), .B2(n3414), .A(n3413), .ZN(n3415) );
  NAND2_X1 U4293 ( .A1(n4125), .A2(n3415), .ZN(U3244) );
  INV_X1 U4294 ( .A(n3416), .ZN(n3417) );
  NOR2_X1 U4295 ( .A1(n3447), .A2(n3417), .ZN(n3433) );
  NAND2_X1 U4296 ( .A1(n4091), .A2(n3447), .ZN(n4004) );
  INV_X1 U4297 ( .A(n4333), .ZN(n4436) );
  NOR2_X1 U4298 ( .A1(n4436), .A2(n4491), .ZN(n3418) );
  OAI22_X1 U4299 ( .A1(n3985), .A2(n3418), .B1(n2850), .B2(n4878), .ZN(n3432)
         );
  AOI21_X1 U4300 ( .B1(n3433), .B2(n3419), .A(n3432), .ZN(n3431) );
  NAND4_X1 U4301 ( .A1(n3423), .A2(n3422), .A3(n3421), .A4(n3420), .ZN(n3424)
         );
  INV_X1 U4302 ( .A(n3985), .ZN(n3434) );
  OR2_X1 U4303 ( .A1(n3425), .A2(n4179), .ZN(n3593) );
  INV_X1 U4304 ( .A(n3593), .ZN(n3426) );
  NAND2_X1 U4305 ( .A1(n4724), .A2(n3426), .ZN(n4343) );
  INV_X1 U4306 ( .A(n4343), .ZN(n4829) );
  OAI22_X1 U4307 ( .A1(n4724), .A2(n3428), .B1(n3427), .B2(n4478), .ZN(n3429)
         );
  AOI21_X1 U4308 ( .B1(n3434), .B2(n4829), .A(n3429), .ZN(n3430) );
  OAI21_X1 U4309 ( .B1(n3431), .B2(n4493), .A(n3430), .ZN(U3290) );
  INV_X1 U4310 ( .A(n4884), .ZN(n4908) );
  AOI211_X1 U4311 ( .C1(n4908), .C2(n3434), .A(n3433), .B(n3432), .ZN(n4873)
         );
  INV_X1 U4312 ( .A(n4920), .ZN(n4918) );
  NAND2_X1 U4313 ( .A1(n4918), .A2(REG1_REG_0__SCAN_IN), .ZN(n3435) );
  OAI21_X1 U4314 ( .B1(n4873), .B2(n4918), .A(n3435), .ZN(U3518) );
  NAND2_X1 U4315 ( .A1(n2902), .A2(n4002), .ZN(n3436) );
  NAND2_X1 U4316 ( .A1(n3520), .A2(n3436), .ZN(n3440) );
  NAND2_X1 U4317 ( .A1(n3456), .A2(n4627), .ZN(n3438) );
  NAND2_X1 U4318 ( .A1(n4091), .A2(n4881), .ZN(n3437) );
  OAI211_X1 U4319 ( .C1(n2852), .C2(n4878), .A(n3438), .B(n3437), .ZN(n3439)
         );
  AOI21_X1 U4320 ( .B1(n3440), .B2(n4491), .A(n3439), .ZN(n3445) );
  OR2_X1 U4321 ( .A1(n3441), .A2(n2902), .ZN(n3442) );
  AND2_X1 U4322 ( .A1(n3443), .A2(n3442), .ZN(n3517) );
  NAND2_X1 U4323 ( .A1(n3517), .A2(n4436), .ZN(n3444) );
  NAND2_X1 U4324 ( .A1(n3445), .A2(n3444), .ZN(n3514) );
  INV_X1 U4325 ( .A(n3517), .ZN(n3448) );
  INV_X1 U4326 ( .A(n4585), .ZN(n4902) );
  OAI21_X1 U4327 ( .B1(n3447), .B2(n3446), .A(n3528), .ZN(n3513) );
  OAI22_X1 U4328 ( .A1(n3448), .A2(n4884), .B1(n4902), .B2(n3513), .ZN(n3449)
         );
  NOR2_X1 U4329 ( .A1(n3514), .A2(n3449), .ZN(n4875) );
  NAND2_X1 U4330 ( .A1(n4918), .A2(REG1_REG_1__SCAN_IN), .ZN(n3450) );
  OAI21_X1 U4331 ( .B1(n4875), .B2(n4918), .A(n3450), .ZN(U3519) );
  OAI211_X1 U4332 ( .C1(n3451), .C2(n3452), .A(n3453), .B(n3918), .ZN(n3458)
         );
  OAI22_X1 U4333 ( .A1(n3454), .A2(n3921), .B1(n2852), .B2(n3923), .ZN(n3455)
         );
  AOI21_X1 U4334 ( .B1(n3456), .B2(n3465), .A(n3455), .ZN(n3457) );
  OAI211_X1 U4335 ( .C1(n3459), .C2(n3512), .A(n3458), .B(n3457), .ZN(U3219)
         );
  INV_X1 U4336 ( .A(n3461), .ZN(n3463) );
  AOI21_X1 U4337 ( .B1(n3464), .B2(n3460), .A(n3463), .ZN(n3471) );
  AOI22_X1 U4338 ( .A1(n3375), .A2(n3466), .B1(n3906), .B2(n3551), .ZN(n3467)
         );
  OAI21_X1 U4339 ( .B1(n3920), .B2(n4877), .A(n3467), .ZN(n3468) );
  AOI21_X1 U4340 ( .B1(REG3_REG_2__SCAN_IN), .B2(n3469), .A(n3468), .ZN(n3470)
         );
  OAI21_X1 U4341 ( .B1(n3471), .B2(n3898), .A(n3470), .ZN(U3234) );
  XNOR2_X1 U4342 ( .A(n3472), .B(n3473), .ZN(n3474) );
  NAND2_X1 U4343 ( .A1(n3474), .A2(n3918), .ZN(n3481) );
  OAI22_X1 U4344 ( .A1(n2852), .A2(n3921), .B1(n3920), .B2(n3475), .ZN(n3479)
         );
  INV_X1 U4345 ( .A(n3476), .ZN(n3477) );
  OAI21_X1 U4346 ( .B1(n2857), .B2(n3923), .A(n3477), .ZN(n3478) );
  NOR2_X1 U4347 ( .A1(n3479), .A2(n3478), .ZN(n3480) );
  OAI211_X1 U4348 ( .C1(REG3_REG_3__SCAN_IN), .C2(n3928), .A(n3481), .B(n3480), 
        .ZN(U3215) );
  XNOR2_X1 U4349 ( .A(n3482), .B(n3992), .ZN(n3545) );
  INV_X1 U4350 ( .A(n3545), .ZN(n3489) );
  AOI22_X1 U4351 ( .A1(n4089), .A2(n4592), .B1(n4627), .B2(n3542), .ZN(n3483)
         );
  OAI21_X1 U4352 ( .B1(n2852), .B2(n4615), .A(n3483), .ZN(n3488) );
  OAI21_X1 U4353 ( .B1(n3992), .B2(n3485), .A(n3484), .ZN(n3486) );
  NAND2_X1 U4354 ( .A1(n3486), .A2(n4491), .ZN(n3487) );
  OAI21_X1 U4355 ( .B1(n3545), .B2(n4333), .A(n3487), .ZN(n3535) );
  AOI211_X1 U4356 ( .C1(n4908), .C2(n3489), .A(n3488), .B(n3535), .ZN(n3493)
         );
  INV_X1 U4357 ( .A(n3527), .ZN(n3490) );
  AOI21_X1 U4358 ( .B1(n3542), .B2(n3490), .A(n3556), .ZN(n3538) );
  INV_X1 U4359 ( .A(n4640), .ZN(n4912) );
  AOI22_X1 U4360 ( .A1(n3538), .A2(n4912), .B1(REG1_REG_3__SCAN_IN), .B2(n4918), .ZN(n3491) );
  OAI21_X1 U4361 ( .B1(n3493), .B2(n4918), .A(n3491), .ZN(U3521) );
  INV_X1 U4362 ( .A(n4706), .ZN(n4886) );
  AOI22_X1 U4363 ( .A1(n3538), .A2(n4886), .B1(REG0_REG_3__SCAN_IN), .B2(n3250), .ZN(n3492) );
  OAI21_X1 U4364 ( .B1(n3493), .B2(n3250), .A(n3492), .ZN(U3473) );
  OR2_X1 U4365 ( .A1(n3494), .A2(n3495), .ZN(n3547) );
  NAND2_X1 U4366 ( .A1(n3547), .A2(n3496), .ZN(n3499) );
  INV_X1 U4367 ( .A(n3497), .ZN(n4015) );
  NAND2_X1 U4368 ( .A1(n4015), .A2(n4029), .ZN(n3977) );
  INV_X1 U4369 ( .A(n3977), .ZN(n3498) );
  XNOR2_X1 U4370 ( .A(n3499), .B(n3498), .ZN(n3602) );
  NAND2_X1 U4371 ( .A1(n3602), .A2(n4895), .ZN(n3505) );
  AOI22_X1 U4372 ( .A1(n3676), .A2(n4592), .B1(n4627), .B2(n3506), .ZN(n3500)
         );
  OAI21_X1 U4373 ( .B1(n2857), .B2(n4615), .A(n3500), .ZN(n3501) );
  INV_X1 U4374 ( .A(n3501), .ZN(n3504) );
  XNOR2_X1 U4375 ( .A(n3502), .B(n3977), .ZN(n3503) );
  NAND2_X1 U4376 ( .A1(n3503), .A2(n4491), .ZN(n3599) );
  NAND3_X1 U4377 ( .A1(n3505), .A2(n3504), .A3(n3599), .ZN(n3604) );
  INV_X1 U4378 ( .A(n3604), .ZN(n3510) );
  NAND2_X1 U4379 ( .A1(n3554), .A2(n3506), .ZN(n3507) );
  NAND2_X1 U4380 ( .A1(n3622), .A2(n3507), .ZN(n3607) );
  INV_X1 U4381 ( .A(n3607), .ZN(n3508) );
  AOI22_X1 U4382 ( .A1(n3508), .A2(n4886), .B1(REG0_REG_5__SCAN_IN), .B2(n3250), .ZN(n3509) );
  OAI21_X1 U4383 ( .B1(n3510), .B2(n3250), .A(n3509), .ZN(U3477) );
  NAND2_X1 U4384 ( .A1(n4727), .A2(n3511), .ZN(n4488) );
  OAI22_X1 U4385 ( .A1(n4488), .A2(n3513), .B1(n3512), .B2(n4478), .ZN(n3516)
         );
  MUX2_X1 U4386 ( .A(n3514), .B(REG2_REG_1__SCAN_IN), .S(n4493), .Z(n3515) );
  AOI211_X1 U4387 ( .C1(n3517), .C2(n4829), .A(n3516), .B(n3515), .ZN(n3518)
         );
  INV_X1 U4388 ( .A(n3518), .ZN(U3289) );
  OAI21_X1 U4389 ( .B1(n2218), .B2(n3521), .A(n3519), .ZN(n3525) );
  INV_X1 U4390 ( .A(n3525), .ZN(n4885) );
  NAND3_X1 U4391 ( .A1(n3521), .A2(n2903), .A3(n3520), .ZN(n3522) );
  AOI21_X1 U4392 ( .B1(n3523), .B2(n3522), .A(n4637), .ZN(n3524) );
  AOI21_X1 U4393 ( .B1(n3525), .B2(n4436), .A(n3524), .ZN(n4883) );
  MUX2_X1 U4394 ( .A(n3526), .B(n4883), .S(n4724), .Z(n3534) );
  NAND2_X1 U4395 ( .A1(n4727), .A2(n4627), .ZN(n4483) );
  NAND2_X1 U4396 ( .A1(n4727), .A2(n4592), .ZN(n4468) );
  OAI22_X1 U4397 ( .A1(n4879), .A2(n4468), .B1(n4111), .B2(n4478), .ZN(n3531)
         );
  AOI21_X1 U4398 ( .B1(n3532), .B2(n3528), .A(n3527), .ZN(n4911) );
  INV_X1 U4399 ( .A(n4911), .ZN(n3529) );
  NAND2_X1 U4400 ( .A1(n4727), .A2(n4881), .ZN(n4484) );
  OAI22_X1 U4401 ( .A1(n3529), .A2(n4488), .B1(n2850), .B2(n4484), .ZN(n3530)
         );
  AOI211_X1 U4402 ( .C1(n3532), .C2(n4462), .A(n3531), .B(n3530), .ZN(n3533)
         );
  OAI211_X1 U4403 ( .C1(n4885), .C2(n4343), .A(n3534), .B(n3533), .ZN(U3288)
         );
  NAND2_X1 U4404 ( .A1(n3535), .A2(n4727), .ZN(n3544) );
  INV_X1 U4405 ( .A(n4478), .ZN(n4823) );
  AOI22_X1 U4406 ( .A1(n4825), .A2(REG2_REG_3__SCAN_IN), .B1(n4823), .B2(n3536), .ZN(n3537) );
  OAI21_X1 U4407 ( .B1(n2857), .B2(n4468), .A(n3537), .ZN(n3541) );
  INV_X1 U4408 ( .A(n3538), .ZN(n3539) );
  OAI22_X1 U4409 ( .A1(n3539), .A2(n4488), .B1(n2852), .B2(n4484), .ZN(n3540)
         );
  AOI211_X1 U4410 ( .C1(n3542), .C2(n4462), .A(n3541), .B(n3540), .ZN(n3543)
         );
  OAI211_X1 U4411 ( .C1(n3545), .C2(n4343), .A(n3544), .B(n3543), .ZN(U3287)
         );
  NAND2_X1 U4412 ( .A1(n3494), .A2(n3495), .ZN(n3546) );
  NAND2_X1 U4413 ( .A1(n3547), .A2(n3546), .ZN(n4889) );
  XOR2_X1 U4414 ( .A(n3495), .B(n3548), .Z(n3553) );
  OAI22_X1 U4415 ( .A1(n2859), .A2(n4878), .B1(n3555), .B2(n4876), .ZN(n3550)
         );
  NOR2_X1 U4416 ( .A1(n4889), .A2(n4333), .ZN(n3549) );
  AOI211_X1 U4417 ( .C1(n4881), .C2(n3551), .A(n3550), .B(n3549), .ZN(n3552)
         );
  OAI21_X1 U4418 ( .B1(n4637), .B2(n3553), .A(n3552), .ZN(n4891) );
  OAI211_X1 U4419 ( .C1(n3556), .C2(n3555), .A(n4585), .B(n3554), .ZN(n4890)
         );
  OAI22_X1 U4420 ( .A1(n4890), .A2(n4379), .B1(n4478), .B2(n3557), .ZN(n3558)
         );
  OAI21_X1 U4421 ( .B1(n4891), .B2(n3558), .A(n4727), .ZN(n3560) );
  NAND2_X1 U4422 ( .A1(n4493), .A2(REG2_REG_4__SCAN_IN), .ZN(n3559) );
  OAI211_X1 U4423 ( .C1(n4889), .C2(n4343), .A(n3560), .B(n3559), .ZN(U3286)
         );
  NAND2_X1 U4424 ( .A1(n3577), .A2(REG1_REG_11__SCAN_IN), .ZN(n3567) );
  AOI22_X1 U4425 ( .A1(n3577), .A2(REG1_REG_11__SCAN_IN), .B1(n2566), .B2(
        n4865), .ZN(n4761) );
  AOI22_X1 U4426 ( .A1(REG1_REG_9__SCAN_IN), .A2(n3578), .B1(n4868), .B2(n3734), .ZN(n4740) );
  NOR2_X1 U4427 ( .A1(n4715), .A2(REG1_REG_7__SCAN_IN), .ZN(n3561) );
  INV_X1 U4428 ( .A(n4715), .ZN(n3580) );
  OAI22_X1 U4429 ( .A1(n3562), .A2(n3561), .B1(n3385), .B2(n3580), .ZN(n3563)
         );
  NAND2_X1 U4430 ( .A1(n3563), .A2(n3581), .ZN(n3564) );
  XNOR2_X1 U4431 ( .A(n3563), .B(n4870), .ZN(n4735) );
  NAND2_X1 U4432 ( .A1(REG1_REG_8__SCAN_IN), .A2(n4735), .ZN(n4734) );
  NAND2_X1 U4433 ( .A1(n4749), .A2(n3565), .ZN(n3566) );
  NAND2_X1 U4434 ( .A1(REG1_REG_10__SCAN_IN), .A2(n4756), .ZN(n4755) );
  NAND2_X1 U4435 ( .A1(n3586), .A2(n3568), .ZN(n3569) );
  NAND2_X1 U4436 ( .A1(REG1_REG_12__SCAN_IN), .A2(n4771), .ZN(n4770) );
  NAND2_X1 U4437 ( .A1(n3569), .A2(n4770), .ZN(n3573) );
  NAND2_X1 U4438 ( .A1(n4155), .A2(n4142), .ZN(n3570) );
  OAI21_X1 U4439 ( .B1(n4155), .B2(n4142), .A(n3570), .ZN(n3572) );
  NAND2_X1 U4440 ( .A1(n4141), .A2(n4142), .ZN(n3571) );
  OAI211_X1 U4441 ( .C1(n4141), .C2(n4142), .A(n3573), .B(n3571), .ZN(n4140)
         );
  OAI211_X1 U4442 ( .C1(n3573), .C2(n3572), .A(n4140), .B(n4816), .ZN(n3575)
         );
  AND2_X1 U4443 ( .A1(U3149), .A2(REG3_REG_13__SCAN_IN), .ZN(n3866) );
  AOI21_X1 U4444 ( .B1(n4815), .B2(ADDR_REG_13__SCAN_IN), .A(n3866), .ZN(n3574) );
  OAI211_X1 U4445 ( .C1(n4822), .C2(n4141), .A(n3575), .B(n3574), .ZN(n3592)
         );
  INV_X1 U4446 ( .A(REG2_REG_13__SCAN_IN), .ZN(n3576) );
  NOR2_X1 U4447 ( .A1(n4141), .A2(n3576), .ZN(n4156) );
  AOI21_X1 U4448 ( .B1(n3576), .B2(n4141), .A(n4156), .ZN(n3590) );
  AOI22_X1 U4449 ( .A1(n3577), .A2(REG2_REG_11__SCAN_IN), .B1(n3688), .B2(
        n4865), .ZN(n4764) );
  AOI22_X1 U4450 ( .A1(REG2_REG_9__SCAN_IN), .A2(n3578), .B1(n4868), .B2(n3643), .ZN(n4743) );
  NAND2_X1 U4451 ( .A1(n3581), .A2(n3582), .ZN(n3583) );
  NAND2_X1 U4452 ( .A1(REG2_REG_8__SCAN_IN), .A2(n4730), .ZN(n4729) );
  NAND2_X1 U4453 ( .A1(n4749), .A2(n3584), .ZN(n3585) );
  NAND2_X1 U4454 ( .A1(REG2_REG_10__SCAN_IN), .A2(n4751), .ZN(n4750) );
  NAND2_X1 U4455 ( .A1(n3586), .A2(n3587), .ZN(n3588) );
  NAND2_X1 U4456 ( .A1(REG2_REG_12__SCAN_IN), .A2(n4774), .ZN(n4772) );
  NAND2_X1 U4457 ( .A1(n3588), .A2(n4772), .ZN(n4157) );
  OAI21_X1 U4458 ( .B1(n3590), .B2(n4157), .A(n4773), .ZN(n3589) );
  AOI21_X1 U4459 ( .B1(n3590), .B2(n4157), .A(n3589), .ZN(n3591) );
  OR2_X1 U4460 ( .A1(n3592), .A2(n3591), .ZN(U3253) );
  NAND2_X1 U4461 ( .A1(n4333), .A2(n3593), .ZN(n3594) );
  INV_X1 U4462 ( .A(n4468), .ZN(n4482) );
  OAI22_X1 U4463 ( .A1(n4724), .A2(n4132), .B1(n3615), .B2(n4478), .ZN(n3595)
         );
  AOI21_X1 U4464 ( .B1(n4482), .B2(n3676), .A(n3595), .ZN(n3598) );
  OAI22_X1 U4465 ( .A1(n2857), .A2(n4484), .B1(n4483), .B2(n3611), .ZN(n3596)
         );
  INV_X1 U4466 ( .A(n3596), .ZN(n3597) );
  OAI211_X1 U4467 ( .C1(n3607), .C2(n4488), .A(n3598), .B(n3597), .ZN(n3601)
         );
  NOR2_X1 U4468 ( .A1(n3599), .A2(n4493), .ZN(n3600) );
  AOI211_X1 U4469 ( .C1(n3602), .C2(n4496), .A(n3601), .B(n3600), .ZN(n3603)
         );
  INV_X1 U4470 ( .A(n3603), .ZN(U3285) );
  MUX2_X1 U4471 ( .A(REG1_REG_5__SCAN_IN), .B(n3604), .S(n4920), .Z(n3605) );
  INV_X1 U4472 ( .A(n3605), .ZN(n3606) );
  OAI21_X1 U4473 ( .B1(n4640), .B2(n3607), .A(n3606), .ZN(U3523) );
  OAI211_X1 U4474 ( .C1(n3610), .C2(n3609), .A(n3608), .B(n3918), .ZN(n3614)
         );
  AND2_X1 U4475 ( .A1(U3149), .A2(REG3_REG_5__SCAN_IN), .ZN(n4127) );
  OAI22_X1 U4476 ( .A1(n2857), .A2(n3921), .B1(n3920), .B2(n3611), .ZN(n3612)
         );
  AOI211_X1 U4477 ( .C1(n3906), .C2(n3676), .A(n4127), .B(n3612), .ZN(n3613)
         );
  OAI211_X1 U4478 ( .C1(n3928), .C2(n3615), .A(n3614), .B(n3613), .ZN(U3224)
         );
  XOR2_X1 U4479 ( .A(n3991), .B(n3616), .Z(n3767) );
  XNOR2_X1 U4480 ( .A(n3617), .B(n3991), .ZN(n3765) );
  AOI22_X1 U4481 ( .A1(n4087), .A2(n4592), .B1(n4627), .B2(n3621), .ZN(n3618)
         );
  OAI21_X1 U4482 ( .B1(n2859), .B2(n4615), .A(n3618), .ZN(n3619) );
  AOI21_X1 U4483 ( .B1(n3765), .B2(n4491), .A(n3619), .ZN(n3620) );
  OAI21_X1 U4484 ( .B1(n3767), .B2(n4589), .A(n3620), .ZN(n3627) );
  NAND2_X1 U4485 ( .A1(n3627), .A2(n4910), .ZN(n3625) );
  AND2_X1 U4486 ( .A1(n3622), .A2(n3621), .ZN(n3623) );
  NOR2_X1 U4487 ( .A1(n3670), .A2(n3623), .ZN(n3754) );
  NAND2_X1 U4488 ( .A1(n3754), .A2(n4886), .ZN(n3624) );
  OAI211_X1 U4489 ( .C1(n4910), .C2(n3626), .A(n3625), .B(n3624), .ZN(U3479)
         );
  NAND2_X1 U4490 ( .A1(n3627), .A2(n4920), .ZN(n3629) );
  NAND2_X1 U4491 ( .A1(n3754), .A2(n4912), .ZN(n3628) );
  OAI211_X1 U4492 ( .C1(n4920), .C2(n2491), .A(n3629), .B(n3628), .ZN(U3524)
         );
  XNOR2_X1 U4493 ( .A(n3631), .B(n3630), .ZN(n3632) );
  XNOR2_X1 U4494 ( .A(n3633), .B(n3632), .ZN(n3634) );
  NAND2_X1 U4495 ( .A1(n3634), .A2(n3918), .ZN(n3638) );
  OAI22_X1 U4496 ( .A1(n2859), .A2(n3921), .B1(n3920), .B2(n3758), .ZN(n3635)
         );
  AOI211_X1 U4497 ( .C1(n3906), .C2(n4087), .A(n3636), .B(n3635), .ZN(n3637)
         );
  OAI211_X1 U4498 ( .C1(n3928), .C2(n3755), .A(n3638), .B(n3637), .ZN(U3236)
         );
  INV_X1 U4499 ( .A(n4026), .ZN(n4033) );
  AND2_X1 U4500 ( .A1(n4033), .A2(n4023), .ZN(n3993) );
  XOR2_X1 U4501 ( .A(n3993), .B(n3639), .Z(n3640) );
  NAND2_X1 U4502 ( .A1(n3640), .A2(n4491), .ZN(n3712) );
  INV_X1 U4503 ( .A(n3696), .ZN(n3642) );
  INV_X1 U4504 ( .A(n3727), .ZN(n3641) );
  OAI21_X1 U4505 ( .B1(n3642), .B2(n3740), .A(n3641), .ZN(n3736) );
  INV_X1 U4506 ( .A(n3736), .ZN(n3647) );
  OAI22_X1 U4507 ( .A1(n3745), .A2(n4478), .B1(n3643), .B2(n4727), .ZN(n3646)
         );
  INV_X1 U4508 ( .A(n4484), .ZN(n4463) );
  AOI22_X1 U4509 ( .A1(n4463), .A2(n3667), .B1(n4482), .B2(n4629), .ZN(n3644)
         );
  OAI21_X1 U4510 ( .B1(n3740), .B2(n4483), .A(n3644), .ZN(n3645) );
  AOI211_X1 U4511 ( .C1(n3647), .C2(n4828), .A(n3646), .B(n3645), .ZN(n3650)
         );
  XNOR2_X1 U4512 ( .A(n3648), .B(n3993), .ZN(n3714) );
  NAND2_X1 U4513 ( .A1(n3714), .A2(n4496), .ZN(n3649) );
  OAI211_X1 U4514 ( .C1(n3712), .C2(n4825), .A(n3650), .B(n3649), .ZN(U3281)
         );
  INV_X1 U4515 ( .A(n3652), .ZN(n3654) );
  NOR2_X1 U4516 ( .A1(n3654), .A2(n3653), .ZN(n3655) );
  XNOR2_X1 U4517 ( .A(n3651), .B(n3655), .ZN(n3661) );
  INV_X1 U4518 ( .A(n3656), .ZN(n4824) );
  NAND2_X1 U4519 ( .A1(REG3_REG_8__SCAN_IN), .A2(U3149), .ZN(n4732) );
  OAI21_X1 U4520 ( .B1(n3721), .B2(n3923), .A(n4732), .ZN(n3659) );
  OAI22_X1 U4521 ( .A1(n3657), .A2(n3921), .B1(n3920), .B2(n3700), .ZN(n3658)
         );
  AOI211_X1 U4522 ( .C1(n4824), .C2(n3895), .A(n3659), .B(n3658), .ZN(n3660)
         );
  OAI21_X1 U4523 ( .B1(n3661), .B2(n3898), .A(n3660), .ZN(U3218) );
  XOR2_X1 U4524 ( .A(n2216), .B(n3662), .Z(n3663) );
  NAND2_X1 U4525 ( .A1(n3663), .A2(n3918), .ZN(n3669) );
  OAI22_X1 U4526 ( .A1(n3664), .A2(n3921), .B1(n3920), .B2(n3671), .ZN(n3665)
         );
  AOI211_X1 U4527 ( .C1(n3906), .C2(n3667), .A(n3666), .B(n3665), .ZN(n3668)
         );
  OAI211_X1 U4528 ( .C1(n3928), .C2(n3678), .A(n3669), .B(n3668), .ZN(U3210)
         );
  OAI211_X1 U4529 ( .C1(n3670), .C2(n3671), .A(n3695), .B(n4585), .ZN(n4899)
         );
  OAI22_X1 U4530 ( .A1(n3741), .A2(n4878), .B1(n3671), .B2(n4876), .ZN(n3675)
         );
  XOR2_X1 U4531 ( .A(n4019), .B(n3672), .Z(n3673) );
  NOR2_X1 U4532 ( .A1(n3673), .A2(n4637), .ZN(n3674) );
  AOI211_X1 U4533 ( .C1(n4881), .C2(n3676), .A(n3675), .B(n3674), .ZN(n4900)
         );
  OAI21_X1 U4534 ( .B1(n4379), .B2(n4899), .A(n4900), .ZN(n3682) );
  NAND2_X1 U4535 ( .A1(n3677), .A2(n4019), .ZN(n4896) );
  AND3_X1 U4536 ( .A1(n4897), .A2(n4896), .A3(n4496), .ZN(n3681) );
  OAI22_X1 U4537 ( .A1(n4724), .A2(n3679), .B1(n3678), .B2(n4478), .ZN(n3680)
         );
  AOI211_X1 U4538 ( .C1(n3682), .C2(n4724), .A(n3681), .B(n3680), .ZN(n3683)
         );
  INV_X1 U4539 ( .A(n3683), .ZN(U3283) );
  XNOR2_X1 U4540 ( .A(n4452), .B(n2873), .ZN(n4636) );
  NAND2_X1 U4541 ( .A1(n4727), .A2(n4491), .ZN(n4473) );
  NAND2_X1 U4542 ( .A1(n3684), .A2(n3979), .ZN(n3685) );
  NAND2_X1 U4543 ( .A1(n3686), .A2(n3685), .ZN(n4626) );
  OR2_X1 U4544 ( .A1(n4903), .A2(n3883), .ZN(n3687) );
  NAND2_X1 U4545 ( .A1(n2215), .A2(n3687), .ZN(n4707) );
  OAI22_X1 U4546 ( .A1(n4724), .A2(n3688), .B1(n3888), .B2(n4478), .ZN(n3689)
         );
  AOI21_X1 U4547 ( .B1(n4482), .B2(n4607), .A(n3689), .ZN(n3692) );
  OAI22_X1 U4548 ( .A1(n3884), .A2(n4484), .B1(n4483), .B2(n3883), .ZN(n3690)
         );
  INV_X1 U4549 ( .A(n3690), .ZN(n3691) );
  OAI211_X1 U4550 ( .C1(n4707), .C2(n4488), .A(n3692), .B(n3691), .ZN(n3693)
         );
  AOI21_X1 U4551 ( .B1(n4626), .B2(n4496), .A(n3693), .ZN(n3694) );
  OAI21_X1 U4552 ( .B1(n4636), .B2(n4473), .A(n3694), .ZN(U3279) );
  INV_X1 U4553 ( .A(n3695), .ZN(n3697) );
  OAI21_X1 U4554 ( .B1(n3697), .B2(n3700), .A(n3696), .ZN(n4826) );
  INV_X1 U4555 ( .A(REG0_REG_8__SCAN_IN), .ZN(n3706) );
  XNOR2_X1 U4556 ( .A(n3698), .B(n3989), .ZN(n4830) );
  XNOR2_X1 U4557 ( .A(n3699), .B(n3989), .ZN(n3703) );
  OAI22_X1 U4558 ( .A1(n3721), .A2(n4878), .B1(n4876), .B2(n3700), .ZN(n3701)
         );
  AOI21_X1 U4559 ( .B1(n4881), .B2(n4087), .A(n3701), .ZN(n3702) );
  OAI21_X1 U4560 ( .B1(n3703), .B2(n4637), .A(n3702), .ZN(n3704) );
  AOI21_X1 U4561 ( .B1(n4436), .B2(n4830), .A(n3704), .ZN(n4833) );
  INV_X1 U4562 ( .A(n4833), .ZN(n3705) );
  AOI21_X1 U4563 ( .B1(n4908), .B2(n4830), .A(n3705), .ZN(n3708) );
  MUX2_X1 U4564 ( .A(n3706), .B(n3708), .S(n4910), .Z(n3707) );
  OAI21_X1 U4565 ( .B1(n4826), .B2(n4706), .A(n3707), .ZN(U3483) );
  MUX2_X1 U4566 ( .A(n2516), .B(n3708), .S(n4920), .Z(n3709) );
  OAI21_X1 U4567 ( .B1(n4826), .B2(n4640), .A(n3709), .ZN(U3526) );
  AOI22_X1 U4568 ( .A1(n4629), .A2(n4592), .B1(n4627), .B2(n3710), .ZN(n3711)
         );
  OAI211_X1 U4569 ( .C1(n3741), .C2(n4615), .A(n3712), .B(n3711), .ZN(n3713)
         );
  AOI21_X1 U4570 ( .B1(n3714), .B2(n4895), .A(n3713), .ZN(n3733) );
  MUX2_X1 U4571 ( .A(n3162), .B(n3733), .S(n4910), .Z(n3715) );
  OAI21_X1 U4572 ( .B1(n3736), .B2(n4706), .A(n3715), .ZN(U3485) );
  NAND2_X1 U4573 ( .A1(n4037), .A2(n4038), .ZN(n3973) );
  XOR2_X1 U4574 ( .A(n3973), .B(n3716), .Z(n3725) );
  XOR2_X1 U4575 ( .A(n3973), .B(n3717), .Z(n3723) );
  AOI22_X1 U4576 ( .A1(n3719), .A2(n4592), .B1(n4627), .B2(n3718), .ZN(n3720)
         );
  OAI21_X1 U4577 ( .B1(n3721), .B2(n4615), .A(n3720), .ZN(n3722) );
  AOI21_X1 U4578 ( .B1(n3723), .B2(n4491), .A(n3722), .ZN(n3724) );
  OAI21_X1 U4579 ( .B1(n3725), .B2(n4333), .A(n3724), .ZN(n4905) );
  INV_X1 U4580 ( .A(n4905), .ZN(n3732) );
  INV_X1 U4581 ( .A(n3725), .ZN(n4907) );
  NOR2_X1 U4582 ( .A1(n3727), .A2(n3726), .ZN(n4904) );
  NOR3_X1 U4583 ( .A1(n4904), .A2(n4903), .A3(n4488), .ZN(n3730) );
  OAI22_X1 U4584 ( .A1(n4724), .A2(n3179), .B1(n3728), .B2(n4478), .ZN(n3729)
         );
  AOI211_X1 U4585 ( .C1(n4907), .C2(n4829), .A(n3730), .B(n3729), .ZN(n3731)
         );
  OAI21_X1 U4586 ( .B1(n3732), .B2(n4493), .A(n3731), .ZN(U3280) );
  MUX2_X1 U4587 ( .A(n3734), .B(n3733), .S(n4920), .Z(n3735) );
  OAI21_X1 U4588 ( .B1(n4640), .B2(n3736), .A(n3735), .ZN(U3527) );
  XNOR2_X1 U4589 ( .A(n3737), .B(n3738), .ZN(n3739) );
  NAND2_X1 U4590 ( .A1(n3739), .A2(n3918), .ZN(n3744) );
  AND2_X1 U4591 ( .A1(U3149), .A2(REG3_REG_9__SCAN_IN), .ZN(n4747) );
  OAI22_X1 U4592 ( .A1(n3741), .A2(n3921), .B1(n3920), .B2(n3740), .ZN(n3742)
         );
  AOI211_X1 U4593 ( .C1(n3906), .C2(n4629), .A(n4747), .B(n3742), .ZN(n3743)
         );
  OAI211_X1 U4594 ( .C1(n3928), .C2(n3745), .A(n3744), .B(n3743), .ZN(U3228)
         );
  INV_X1 U4595 ( .A(REG2_REG_28__SCAN_IN), .ZN(n3746) );
  OAI22_X1 U4596 ( .A1(n3747), .A2(n4478), .B1(n4724), .B2(n3746), .ZN(n3748)
         );
  AOI21_X1 U4597 ( .B1(n3749), .B2(n4828), .A(n3748), .ZN(n3752) );
  NAND2_X1 U4598 ( .A1(n3750), .A2(n4727), .ZN(n3751) );
  OAI211_X1 U4599 ( .C1(n3753), .C2(n4415), .A(n3752), .B(n3751), .ZN(U3262)
         );
  INV_X1 U4600 ( .A(n4473), .ZN(n3764) );
  NAND2_X1 U4601 ( .A1(n3754), .A2(n4828), .ZN(n3762) );
  INV_X1 U4602 ( .A(REG2_REG_6__SCAN_IN), .ZN(n3756) );
  OAI22_X1 U4603 ( .A1(n4724), .A2(n3756), .B1(n3755), .B2(n4478), .ZN(n3757)
         );
  AOI21_X1 U4604 ( .B1(n4482), .B2(n4087), .A(n3757), .ZN(n3761) );
  OAI22_X1 U4605 ( .A1(n2859), .A2(n4484), .B1(n4483), .B2(n3758), .ZN(n3759)
         );
  INV_X1 U4606 ( .A(n3759), .ZN(n3760) );
  NAND3_X1 U4607 ( .A1(n3762), .A2(n3761), .A3(n3760), .ZN(n3763) );
  AOI21_X1 U4608 ( .B1(n3765), .B2(n3764), .A(n3763), .ZN(n3766) );
  OAI21_X1 U4609 ( .B1(n3767), .B2(n4415), .A(n3766), .ZN(U3284) );
  NAND2_X1 U4610 ( .A1(n2356), .A2(n3769), .ZN(n3770) );
  XNOR2_X1 U4611 ( .A(n3768), .B(n3770), .ZN(n3771) );
  NAND2_X1 U4612 ( .A1(n3771), .A2(n3918), .ZN(n3775) );
  OAI22_X1 U4613 ( .A1(n4614), .A2(n3921), .B1(n3920), .B2(n4443), .ZN(n3773)
         );
  NAND2_X1 U4614 ( .A1(REG3_REG_14__SCAN_IN), .A2(U3149), .ZN(n4780) );
  OAI21_X1 U4615 ( .B1(n4583), .B2(n3923), .A(n4780), .ZN(n3772) );
  NOR2_X1 U4616 ( .A1(n3773), .A2(n3772), .ZN(n3774) );
  OAI211_X1 U4617 ( .C1(n3928), .C2(n4444), .A(n3775), .B(n3774), .ZN(U3212)
         );
  INV_X1 U4618 ( .A(n3776), .ZN(n3780) );
  OAI21_X1 U4619 ( .B1(n2193), .B2(n3778), .A(n3777), .ZN(n3779) );
  NAND3_X1 U4620 ( .A1(n3780), .A2(n3918), .A3(n3779), .ZN(n3784) );
  NOR2_X1 U4621 ( .A1(n4279), .A2(n3923), .ZN(n3782) );
  OAI22_X1 U4622 ( .A1(n4318), .A2(n3921), .B1(n3920), .B2(n4278), .ZN(n3781)
         );
  AOI211_X1 U4623 ( .C1(REG3_REG_23__SCAN_IN), .C2(U3149), .A(n3782), .B(n3781), .ZN(n3783) );
  OAI211_X1 U4624 ( .C1(n3928), .C2(n4286), .A(n3784), .B(n3783), .ZN(U3213)
         );
  XNOR2_X1 U4625 ( .A(n3786), .B(n3785), .ZN(n3787) );
  NAND2_X1 U4626 ( .A1(n3787), .A2(n3918), .ZN(n3791) );
  NOR2_X1 U4627 ( .A1(n3788), .A2(STATE_REG_SCAN_IN), .ZN(n4181) );
  OAI22_X1 U4628 ( .A1(n4395), .A2(n3921), .B1(n3920), .B2(n4357), .ZN(n3789)
         );
  AOI211_X1 U4629 ( .C1(n3906), .C2(n4354), .A(n4181), .B(n3789), .ZN(n3790)
         );
  OAI211_X1 U4630 ( .C1(n3928), .C2(n4360), .A(n3791), .B(n3790), .ZN(U3216)
         );
  AOI21_X1 U4631 ( .B1(n3792), .B2(n3851), .A(n3852), .ZN(n3796) );
  XNOR2_X1 U4632 ( .A(n3794), .B(n3793), .ZN(n3795) );
  XNOR2_X1 U4633 ( .A(n3796), .B(n3795), .ZN(n3802) );
  INV_X1 U4634 ( .A(n3797), .ZN(n4315) );
  OAI22_X1 U4635 ( .A1(n4318), .A2(n3923), .B1(STATE_REG_SCAN_IN), .B2(n3798), 
        .ZN(n3800) );
  OAI22_X1 U4636 ( .A1(n4553), .A2(n3921), .B1(n3920), .B2(n4314), .ZN(n3799)
         );
  AOI211_X1 U4637 ( .C1(n4315), .C2(n3895), .A(n3800), .B(n3799), .ZN(n3801)
         );
  OAI21_X1 U4638 ( .B1(n3802), .B2(n3898), .A(n3801), .ZN(U3220) );
  INV_X1 U4639 ( .A(n3804), .ZN(n3806) );
  NAND2_X1 U4640 ( .A1(n3806), .A2(n3805), .ZN(n3807) );
  XNOR2_X1 U4641 ( .A(n3803), .B(n3807), .ZN(n3808) );
  NAND2_X1 U4642 ( .A1(n3808), .A2(n3918), .ZN(n3812) );
  NOR2_X1 U4643 ( .A1(STATE_REG_SCAN_IN), .A2(n3809), .ZN(n4778) );
  OAI22_X1 U4644 ( .A1(n4616), .A2(n3921), .B1(n3920), .B2(n4613), .ZN(n3810)
         );
  AOI211_X1 U4645 ( .C1(n3906), .C2(n4481), .A(n4778), .B(n3810), .ZN(n3811)
         );
  OAI211_X1 U4646 ( .C1(n3928), .C2(n4479), .A(n3812), .B(n3811), .ZN(U3221)
         );
  INV_X1 U4647 ( .A(n3814), .ZN(n3816) );
  NAND2_X1 U4648 ( .A1(n3816), .A2(n3815), .ZN(n3817) );
  XNOR2_X1 U4649 ( .A(n3813), .B(n3817), .ZN(n3822) );
  OAI22_X1 U4650 ( .A1(n4279), .A2(n3921), .B1(n3920), .B2(n4244), .ZN(n3820)
         );
  OAI22_X1 U4651 ( .A1(n4238), .A2(n3923), .B1(STATE_REG_SCAN_IN), .B2(n3818), 
        .ZN(n3819) );
  AOI211_X1 U4652 ( .C1(n4245), .C2(n3895), .A(n3820), .B(n3819), .ZN(n3821)
         );
  OAI21_X1 U4653 ( .B1(n3822), .B2(n3898), .A(n3821), .ZN(U3222) );
  AOI21_X1 U4654 ( .B1(n3916), .B2(n3913), .A(n3915), .ZN(n3823) );
  XOR2_X1 U4655 ( .A(n3824), .B(n3823), .Z(n3825) );
  NAND2_X1 U4656 ( .A1(n3825), .A2(n3918), .ZN(n3830) );
  NOR2_X1 U4657 ( .A1(STATE_REG_SCAN_IN), .A2(n3826), .ZN(n4804) );
  OAI22_X1 U4658 ( .A1(n4583), .A2(n3921), .B1(n3920), .B2(n3827), .ZN(n3828)
         );
  AOI211_X1 U4659 ( .C1(n3906), .C2(n4581), .A(n4804), .B(n3828), .ZN(n3829)
         );
  OAI211_X1 U4660 ( .C1(n3928), .C2(n4405), .A(n3830), .B(n3829), .ZN(U3223)
         );
  NOR2_X1 U4661 ( .A1(n3833), .A2(n2288), .ZN(n3834) );
  XNOR2_X1 U4662 ( .A(n3831), .B(n3834), .ZN(n3835) );
  NAND2_X1 U4663 ( .A1(n3835), .A2(n3918), .ZN(n3840) );
  OAI22_X1 U4664 ( .A1(n4575), .A2(n3921), .B1(n3920), .B2(n4390), .ZN(n3838)
         );
  AND2_X1 U4665 ( .A1(U3149), .A2(REG3_REG_17__SCAN_IN), .ZN(n4814) );
  INV_X1 U4666 ( .A(n4814), .ZN(n3836) );
  OAI21_X1 U4667 ( .B1(n4395), .B2(n3923), .A(n3836), .ZN(n3837) );
  NOR2_X1 U4668 ( .A1(n3838), .A2(n3837), .ZN(n3839) );
  OAI211_X1 U4669 ( .C1(n3928), .C2(n4391), .A(n3840), .B(n3839), .ZN(U3225)
         );
  NAND2_X1 U4670 ( .A1(n3842), .A2(n3841), .ZN(n3843) );
  XOR2_X1 U4671 ( .A(n3844), .B(n3843), .Z(n3850) );
  INV_X1 U4672 ( .A(n3845), .ZN(n4255) );
  OAI22_X1 U4673 ( .A1(n4294), .A2(n3921), .B1(n3920), .B2(n4530), .ZN(n3848)
         );
  OAI22_X1 U4674 ( .A1(n4531), .A2(n3923), .B1(STATE_REG_SCAN_IN), .B2(n3846), 
        .ZN(n3847) );
  AOI211_X1 U4675 ( .C1(n4255), .C2(n3895), .A(n3848), .B(n3847), .ZN(n3849)
         );
  OAI21_X1 U4676 ( .B1(n3850), .B2(n3898), .A(n3849), .ZN(U3226) );
  NOR2_X1 U4677 ( .A1(n3852), .A2(n2710), .ZN(n3853) );
  XNOR2_X1 U4678 ( .A(n3792), .B(n3853), .ZN(n3859) );
  INV_X1 U4679 ( .A(n4337), .ZN(n3857) );
  INV_X1 U4680 ( .A(REG3_REG_20__SCAN_IN), .ZN(n3854) );
  OAI22_X1 U4681 ( .A1(n3873), .A2(n3923), .B1(STATE_REG_SCAN_IN), .B2(n3854), 
        .ZN(n3856) );
  OAI22_X1 U4682 ( .A1(n4329), .A2(n3921), .B1(n3920), .B2(n4336), .ZN(n3855)
         );
  AOI211_X1 U4683 ( .C1(n3857), .C2(n3895), .A(n3856), .B(n3855), .ZN(n3858)
         );
  OAI21_X1 U4684 ( .B1(n3859), .B2(n3898), .A(n3858), .ZN(U3230) );
  XNOR2_X1 U4685 ( .A(n3861), .B(n3860), .ZN(n3862) );
  XNOR2_X1 U4686 ( .A(n3863), .B(n3862), .ZN(n3864) );
  NAND2_X1 U4687 ( .A1(n3864), .A2(n3918), .ZN(n3868) );
  OAI22_X1 U4688 ( .A1(n4632), .A2(n3921), .B1(n3920), .B2(n4604), .ZN(n3865)
         );
  AOI211_X1 U4689 ( .C1(n3906), .C2(n4423), .A(n3866), .B(n3865), .ZN(n3867)
         );
  OAI211_X1 U4690 ( .C1(n3928), .C2(n4464), .A(n3868), .B(n3867), .ZN(U3231)
         );
  AOI21_X1 U4691 ( .B1(n3870), .B2(n3869), .A(n2193), .ZN(n3877) );
  INV_X1 U4692 ( .A(n3871), .ZN(n4301) );
  INV_X1 U4693 ( .A(REG3_REG_22__SCAN_IN), .ZN(n3872) );
  OAI22_X1 U4694 ( .A1(n4294), .A2(n3923), .B1(STATE_REG_SCAN_IN), .B2(n3872), 
        .ZN(n3875) );
  OAI22_X1 U4695 ( .A1(n3873), .A2(n3921), .B1(n3920), .B2(n4293), .ZN(n3874)
         );
  AOI211_X1 U4696 ( .C1(n4301), .C2(n3895), .A(n3875), .B(n3874), .ZN(n3876)
         );
  OAI21_X1 U4697 ( .B1(n3877), .B2(n3898), .A(n3876), .ZN(U3232) );
  XNOR2_X1 U4698 ( .A(n3880), .B(n3879), .ZN(n3881) );
  XNOR2_X1 U4699 ( .A(n3878), .B(n3881), .ZN(n3882) );
  NAND2_X1 U4700 ( .A1(n3882), .A2(n3918), .ZN(n3887) );
  NOR2_X1 U4701 ( .A1(STATE_REG_SCAN_IN), .A2(n2567), .ZN(n4768) );
  OAI22_X1 U4702 ( .A1(n3884), .A2(n3921), .B1(n3920), .B2(n3883), .ZN(n3885)
         );
  AOI211_X1 U4703 ( .C1(n3906), .C2(n4607), .A(n4768), .B(n3885), .ZN(n3886)
         );
  OAI211_X1 U4704 ( .C1(n3928), .C2(n3888), .A(n3887), .B(n3886), .ZN(U3233)
         );
  XNOR2_X1 U4705 ( .A(n3890), .B(n3889), .ZN(n3891) );
  XNOR2_X1 U4706 ( .A(n3892), .B(n3891), .ZN(n3899) );
  INV_X1 U4707 ( .A(n4380), .ZN(n3896) );
  NAND2_X1 U4708 ( .A1(U3149), .A2(REG3_REG_18__SCAN_IN), .ZN(n4149) );
  OAI21_X1 U4709 ( .B1(n4329), .B2(n3923), .A(n4149), .ZN(n3894) );
  OAI22_X1 U4710 ( .A1(n4409), .A2(n3921), .B1(n3920), .B2(n4370), .ZN(n3893)
         );
  AOI211_X1 U4711 ( .C1(n3896), .C2(n3895), .A(n3894), .B(n3893), .ZN(n3897)
         );
  OAI21_X1 U4712 ( .B1(n3899), .B2(n3898), .A(n3897), .ZN(U3235) );
  INV_X1 U4713 ( .A(n3900), .ZN(n3902) );
  NAND2_X1 U4714 ( .A1(n3902), .A2(n3901), .ZN(n3903) );
  XNOR2_X1 U4715 ( .A(n3904), .B(n3903), .ZN(n3905) );
  NAND2_X1 U4716 ( .A1(n3905), .A2(n3918), .ZN(n3912) );
  NAND2_X1 U4717 ( .A1(n4520), .A2(n3906), .ZN(n3907) );
  OAI21_X1 U4718 ( .B1(STATE_REG_SCAN_IN), .B2(n3908), .A(n3907), .ZN(n3910)
         );
  OAI22_X1 U4719 ( .A1(n4531), .A2(n3921), .B1(n3920), .B2(n4518), .ZN(n3909)
         );
  NOR2_X1 U4720 ( .A1(n3910), .A2(n3909), .ZN(n3911) );
  OAI211_X1 U4721 ( .C1(n3928), .C2(n4219), .A(n3912), .B(n3911), .ZN(U3237)
         );
  INV_X1 U4722 ( .A(n3913), .ZN(n3914) );
  NOR2_X1 U4723 ( .A1(n3915), .A2(n3914), .ZN(n3917) );
  XNOR2_X1 U4724 ( .A(n3917), .B(n3916), .ZN(n3919) );
  NAND2_X1 U4725 ( .A1(n3919), .A2(n3918), .ZN(n3927) );
  OAI22_X1 U4726 ( .A1(n4605), .A2(n3921), .B1(n3920), .B2(n4422), .ZN(n3925)
         );
  AND2_X1 U4727 ( .A1(U3149), .A2(REG3_REG_15__SCAN_IN), .ZN(n4794) );
  INV_X1 U4728 ( .A(n4794), .ZN(n3922) );
  OAI21_X1 U4729 ( .B1(n4575), .B2(n3923), .A(n3922), .ZN(n3924) );
  NOR2_X1 U4730 ( .A1(n3925), .A2(n3924), .ZN(n3926) );
  OAI211_X1 U4731 ( .C1(n3928), .C2(n4424), .A(n3927), .B(n3926), .ZN(U3238)
         );
  NAND2_X1 U4732 ( .A1(n3929), .A2(DATAI_30_), .ZN(n4505) );
  NAND2_X1 U4733 ( .A1(n3929), .A2(DATAI_31_), .ZN(n4188) );
  INV_X1 U4734 ( .A(n3953), .ZN(n3930) );
  NOR2_X1 U4735 ( .A1(n3931), .A2(n3930), .ZN(n3940) );
  NAND2_X1 U4736 ( .A1(n4085), .A2(n3932), .ZN(n3934) );
  NAND2_X1 U4737 ( .A1(n3934), .A2(n3933), .ZN(n4065) );
  INV_X1 U4738 ( .A(n4084), .ZN(n3937) );
  INV_X1 U4739 ( .A(n4187), .ZN(n3936) );
  INV_X1 U4740 ( .A(n4188), .ZN(n3935) );
  NOR2_X1 U4741 ( .A1(n3936), .A2(n3935), .ZN(n4068) );
  AOI21_X1 U4742 ( .B1(n3937), .B2(n4503), .A(n4068), .ZN(n3988) );
  NAND2_X1 U4743 ( .A1(n3939), .A2(n3938), .ZN(n3955) );
  OAI211_X1 U4744 ( .C1(n3940), .C2(n4065), .A(n3988), .B(n3955), .ZN(n4069)
         );
  INV_X1 U4745 ( .A(n4069), .ZN(n3962) );
  INV_X1 U4746 ( .A(n4066), .ZN(n3970) );
  INV_X1 U4747 ( .A(n4065), .ZN(n3941) );
  NAND3_X1 U4748 ( .A1(n4201), .A2(n3970), .A3(n3941), .ZN(n3961) );
  NAND2_X1 U4749 ( .A1(n4084), .A2(n4505), .ZN(n3971) );
  AOI21_X1 U4750 ( .B1(n3971), .B2(n4187), .A(n4188), .ZN(n3960) );
  NAND2_X1 U4751 ( .A1(n3942), .A2(n3945), .ZN(n4044) );
  NAND2_X1 U4752 ( .A1(n3944), .A2(n3943), .ZN(n4025) );
  NAND2_X1 U4753 ( .A1(n4025), .A2(n3945), .ZN(n4043) );
  OAI21_X1 U4754 ( .B1(n4432), .B2(n4044), .A(n4043), .ZN(n3947) );
  INV_X1 U4755 ( .A(n3946), .ZN(n4046) );
  AOI21_X1 U4756 ( .B1(n4050), .B2(n3947), .A(n4046), .ZN(n3950) );
  INV_X1 U4757 ( .A(n3948), .ZN(n4054) );
  OAI21_X1 U4758 ( .B1(n3950), .B2(n4054), .A(n3949), .ZN(n3951) );
  OAI221_X1 U4759 ( .B1(n3952), .B2(n4058), .C1(n3952), .C2(n3951), .A(n4056), 
        .ZN(n3958) );
  NAND4_X1 U4760 ( .A1(n4001), .A2(n3955), .A3(n3954), .A4(n3953), .ZN(n3957)
         );
  INV_X1 U4761 ( .A(n3988), .ZN(n3956) );
  AOI211_X1 U4762 ( .C1(n3958), .C2(n4062), .A(n3957), .B(n3956), .ZN(n3959)
         );
  AOI211_X1 U4763 ( .C1(n3962), .C2(n3961), .A(n3960), .B(n3959), .ZN(n3963)
         );
  AOI21_X1 U4764 ( .B1(n4503), .B2(n4188), .A(n3963), .ZN(n4076) );
  INV_X1 U4765 ( .A(n3964), .ZN(n3968) );
  NAND2_X1 U4766 ( .A1(n4234), .A2(n3965), .ZN(n4251) );
  INV_X1 U4767 ( .A(n4251), .ZN(n4260) );
  NAND2_X1 U4768 ( .A1(n3967), .A2(n3966), .ZN(n4324) );
  NAND3_X1 U4769 ( .A1(n3968), .A2(n4260), .A3(n4324), .ZN(n3984) );
  NAND2_X1 U4770 ( .A1(n3970), .A2(n3969), .ZN(n4215) );
  INV_X1 U4771 ( .A(n4215), .ZN(n4226) );
  OR2_X1 U4772 ( .A1(n4187), .A2(n4188), .ZN(n3972) );
  AND2_X1 U4773 ( .A1(n3972), .A2(n3971), .ZN(n4067) );
  XNOR2_X1 U4774 ( .A(n4614), .B(n4461), .ZN(n4457) );
  NAND2_X1 U4775 ( .A1(n4455), .A2(n4453), .ZN(n4489) );
  NOR4_X1 U4776 ( .A1(n4203), .A2(n4457), .A3(n4489), .A4(n3973), .ZN(n3975)
         );
  NAND4_X1 U4777 ( .A1(n4226), .A2(n4067), .A3(n3975), .A4(n3974), .ZN(n3983)
         );
  NAND2_X1 U4778 ( .A1(n3976), .A2(n4224), .ZN(n4237) );
  NAND2_X1 U4779 ( .A1(n4346), .A2(n4345), .ZN(n4387) );
  OR4_X1 U4780 ( .A1(n4237), .A2(n3977), .A3(n4373), .A4(n4387), .ZN(n3982) );
  NAND4_X1 U4781 ( .A1(n3980), .A2(n3979), .A3(n3495), .A4(n3978), .ZN(n3981)
         );
  NOR4_X1 U4782 ( .A1(n3984), .A2(n3983), .A3(n3982), .A4(n3981), .ZN(n4000)
         );
  XNOR2_X1 U4783 ( .A(n4533), .B(n4283), .ZN(n4276) );
  XNOR2_X1 U4784 ( .A(n4329), .B(n2882), .ZN(n4351) );
  INV_X1 U4785 ( .A(n4351), .ZN(n3999) );
  INV_X1 U4786 ( .A(n2902), .ZN(n3987) );
  INV_X1 U4787 ( .A(n4419), .ZN(n3986) );
  NAND4_X1 U4788 ( .A1(n3988), .A2(n3987), .A3(n3986), .A4(n3985), .ZN(n3997)
         );
  NAND4_X1 U4789 ( .A1(n4303), .A2(n2326), .A3(n4019), .A4(n3989), .ZN(n3996)
         );
  INV_X1 U4790 ( .A(n3990), .ZN(n4053) );
  NAND4_X1 U4791 ( .A1(n3993), .A2(n4312), .A3(n3992), .A4(n3991), .ZN(n3995)
         );
  NOR4_X1 U4792 ( .A1(n3997), .A2(n3996), .A3(n3995), .A4(n3994), .ZN(n3998)
         );
  NAND4_X1 U4793 ( .A1(n4000), .A2(n4276), .A3(n3999), .A4(n3998), .ZN(n4073)
         );
  INV_X1 U4794 ( .A(n4001), .ZN(n4063) );
  INV_X1 U4795 ( .A(n4002), .ZN(n4006) );
  OAI211_X1 U4796 ( .C1(n4006), .C2(n4005), .A(n4004), .B(n4003), .ZN(n4008)
         );
  NAND3_X1 U4797 ( .A1(n4008), .A2(n4007), .A3(n2903), .ZN(n4011) );
  NAND3_X1 U4798 ( .A1(n4011), .A2(n4010), .A3(n4009), .ZN(n4014) );
  NAND3_X1 U4799 ( .A1(n4014), .A2(n4013), .A3(n4012), .ZN(n4016) );
  NAND4_X1 U4800 ( .A1(n4017), .A2(n4016), .A3(n4015), .A4(n4031), .ZN(n4020)
         );
  NAND3_X1 U4801 ( .A1(n4020), .A2(n4019), .A3(n4018), .ZN(n4021) );
  NAND3_X1 U4802 ( .A1(n4021), .A2(n4028), .A3(n4032), .ZN(n4024) );
  AND3_X1 U4803 ( .A1(n4024), .A2(n4023), .A3(n4022), .ZN(n4027) );
  NOR3_X1 U4804 ( .A1(n4027), .A2(n4026), .A3(n4025), .ZN(n4041) );
  INV_X1 U4805 ( .A(n4028), .ZN(n4030) );
  NOR2_X1 U4806 ( .A1(n4030), .A2(n4029), .ZN(n4034) );
  NAND4_X1 U4807 ( .A1(n4034), .A2(n4033), .A3(n4032), .A4(n4031), .ZN(n4036)
         );
  INV_X1 U4808 ( .A(n4043), .ZN(n4035) );
  AOI21_X1 U4809 ( .B1(n4037), .B2(n4036), .A(n4035), .ZN(n4040) );
  OAI211_X1 U4810 ( .C1(n4041), .C2(n4040), .A(n4039), .B(n4038), .ZN(n4048)
         );
  INV_X1 U4811 ( .A(n4042), .ZN(n4045) );
  OAI21_X1 U4812 ( .B1(n4045), .B2(n4044), .A(n4043), .ZN(n4047) );
  AOI21_X1 U4813 ( .B1(n4048), .B2(n4047), .A(n4046), .ZN(n4049) );
  INV_X1 U4814 ( .A(n4049), .ZN(n4051) );
  AOI21_X1 U4815 ( .B1(n4051), .B2(n4050), .A(n4268), .ZN(n4055) );
  INV_X1 U4816 ( .A(n4052), .ZN(n4271) );
  OAI211_X1 U4817 ( .C1(n4055), .C2(n4054), .A(n4053), .B(n4271), .ZN(n4057)
         );
  OAI221_X1 U4818 ( .B1(n4059), .B2(n4058), .C1(n4059), .C2(n4057), .A(n4056), 
        .ZN(n4061) );
  OAI221_X1 U4819 ( .B1(n4063), .B2(n4062), .C1(n4063), .C2(n4061), .A(n4060), 
        .ZN(n4064) );
  NOR3_X1 U4820 ( .A1(n4066), .A2(n4065), .A3(n4064), .ZN(n4070) );
  OAI22_X1 U4821 ( .A1(n4070), .A2(n4069), .B1(n4068), .B2(n4067), .ZN(n4072)
         );
  MUX2_X1 U4822 ( .A(n4073), .B(n4072), .S(n4071), .Z(n4074) );
  OAI21_X1 U4823 ( .B1(n4076), .B2(n4075), .A(n4074), .ZN(n4077) );
  XNOR2_X1 U4824 ( .A(n4077), .B(n4379), .ZN(n4083) );
  NAND2_X1 U4825 ( .A1(n4079), .A2(n4078), .ZN(n4080) );
  OAI211_X1 U4826 ( .C1(n4712), .C2(n4082), .A(n4080), .B(B_REG_SCAN_IN), .ZN(
        n4081) );
  OAI21_X1 U4827 ( .B1(n4083), .B2(n4082), .A(n4081), .ZN(U3239) );
  MUX2_X1 U4828 ( .A(DATAO_REG_30__SCAN_IN), .B(n4084), .S(n2181), .Z(U3580)
         );
  MUX2_X1 U4829 ( .A(DATAO_REG_29__SCAN_IN), .B(n4085), .S(n2181), .Z(U3579)
         );
  MUX2_X1 U4830 ( .A(DATAO_REG_25__SCAN_IN), .B(n4218), .S(n2181), .Z(U3575)
         );
  MUX2_X1 U4831 ( .A(DATAO_REG_24__SCAN_IN), .B(n4240), .S(U4043), .Z(U3574)
         );
  MUX2_X1 U4832 ( .A(DATAO_REG_23__SCAN_IN), .B(n4533), .S(n2181), .Z(U3573)
         );
  MUX2_X1 U4833 ( .A(DATAO_REG_19__SCAN_IN), .B(n4375), .S(n2181), .Z(U3569)
         );
  MUX2_X1 U4834 ( .A(DATAO_REG_18__SCAN_IN), .B(n4572), .S(n2181), .Z(U3568)
         );
  MUX2_X1 U4835 ( .A(DATAO_REG_17__SCAN_IN), .B(n4581), .S(n2181), .Z(U3567)
         );
  MUX2_X1 U4836 ( .A(DATAO_REG_16__SCAN_IN), .B(n4593), .S(n2181), .Z(U3566)
         );
  MUX2_X1 U4837 ( .A(DATAO_REG_14__SCAN_IN), .B(n4423), .S(n2181), .Z(U3564)
         );
  MUX2_X1 U4838 ( .A(DATAO_REG_9__SCAN_IN), .B(n4086), .S(n2181), .Z(U3559) );
  MUX2_X1 U4839 ( .A(DATAO_REG_7__SCAN_IN), .B(n4087), .S(n2181), .Z(U3557) );
  MUX2_X1 U4840 ( .A(DATAO_REG_5__SCAN_IN), .B(n4088), .S(U4043), .Z(U3555) );
  MUX2_X1 U4841 ( .A(DATAO_REG_4__SCAN_IN), .B(n4089), .S(n2181), .Z(U3554) );
  MUX2_X1 U4842 ( .A(DATAO_REG_2__SCAN_IN), .B(n4090), .S(n2181), .Z(U3552) );
  MUX2_X1 U4843 ( .A(DATAO_REG_1__SCAN_IN), .B(n3375), .S(n2181), .Z(U3551) );
  MUX2_X1 U4844 ( .A(DATAO_REG_0__SCAN_IN), .B(n4091), .S(n2181), .Z(U3550) );
  INV_X1 U4845 ( .A(REG1_REG_0__SCAN_IN), .ZN(n4092) );
  NAND3_X1 U4846 ( .A1(n4816), .A2(n4092), .A3(IR_REG_0__SCAN_IN), .ZN(n4100)
         );
  AOI22_X1 U4847 ( .A1(n4815), .A2(ADDR_REG_0__SCAN_IN), .B1(
        REG3_REG_0__SCAN_IN), .B2(U3149), .ZN(n4099) );
  AOI21_X1 U4848 ( .B1(n4093), .B2(n4092), .A(IR_REG_0__SCAN_IN), .ZN(n4096)
         );
  OAI211_X1 U4849 ( .C1(n4097), .C2(n4096), .A(n4095), .B(n4094), .ZN(n4098)
         );
  NAND3_X1 U4850 ( .A1(n4100), .A2(n4099), .A3(n4098), .ZN(U3240) );
  NAND2_X1 U4851 ( .A1(n4170), .A2(n4720), .ZN(n4110) );
  OAI211_X1 U4852 ( .C1(n4103), .C2(n4102), .A(n4816), .B(n4101), .ZN(n4109)
         );
  OAI211_X1 U4853 ( .C1(n4106), .C2(n4105), .A(n4773), .B(n4104), .ZN(n4108)
         );
  AOI22_X1 U4854 ( .A1(n4815), .A2(ADDR_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(U3149), .ZN(n4107) );
  NAND4_X1 U4855 ( .A1(n4110), .A2(n4109), .A3(n4108), .A4(n4107), .ZN(U3241)
         );
  INV_X1 U4856 ( .A(n4719), .ZN(n4114) );
  NOR2_X1 U4857 ( .A1(n4111), .A2(STATE_REG_SCAN_IN), .ZN(n4112) );
  AOI21_X1 U4858 ( .B1(n4815), .B2(ADDR_REG_2__SCAN_IN), .A(n4112), .ZN(n4113)
         );
  OAI21_X1 U4859 ( .B1(n4822), .B2(n4114), .A(n4113), .ZN(n4115) );
  INV_X1 U4860 ( .A(n4115), .ZN(n4124) );
  OAI211_X1 U4861 ( .C1(n4118), .C2(n4117), .A(n4773), .B(n4116), .ZN(n4123)
         );
  OAI211_X1 U4862 ( .C1(n4121), .C2(n4120), .A(n4816), .B(n4119), .ZN(n4122)
         );
  NAND4_X1 U4863 ( .A1(n4125), .A2(n4124), .A3(n4123), .A4(n4122), .ZN(U3242)
         );
  NOR2_X1 U4864 ( .A1(n4822), .A2(n4131), .ZN(n4126) );
  AOI211_X1 U4865 ( .C1(n4815), .C2(ADDR_REG_5__SCAN_IN), .A(n4127), .B(n4126), 
        .ZN(n4139) );
  OAI211_X1 U4866 ( .C1(n4130), .C2(n4129), .A(n4816), .B(n4128), .ZN(n4138)
         );
  MUX2_X1 U4867 ( .A(REG2_REG_5__SCAN_IN), .B(n4132), .S(n4131), .Z(n4133) );
  INV_X1 U4868 ( .A(n4133), .ZN(n4136) );
  OAI211_X1 U4869 ( .C1(n4136), .C2(n4135), .A(n4773), .B(n4134), .ZN(n4137)
         );
  NAND3_X1 U4870 ( .A1(n4139), .A2(n4138), .A3(n4137), .ZN(U3245) );
  NOR2_X1 U4871 ( .A1(n4165), .A2(REG1_REG_17__SCAN_IN), .ZN(n4148) );
  NAND2_X1 U4872 ( .A1(REG1_REG_15__SCAN_IN), .A2(n4161), .ZN(n4145) );
  INV_X1 U4873 ( .A(n4161), .ZN(n4859) );
  AOI22_X1 U4874 ( .A1(REG1_REG_15__SCAN_IN), .A2(n4161), .B1(n4859), .B2(
        n4598), .ZN(n4797) );
  NAND2_X1 U4875 ( .A1(n4154), .A2(n4143), .ZN(n4144) );
  NAND2_X1 U4876 ( .A1(n4797), .A2(n4796), .ZN(n4795) );
  NOR2_X1 U4877 ( .A1(n4162), .A2(n4146), .ZN(n4147) );
  AOI22_X1 U4878 ( .A1(n4165), .A2(n4578), .B1(REG1_REG_17__SCAN_IN), .B2(
        n4855), .ZN(n4817) );
  XOR2_X1 U4879 ( .A(REG1_REG_18__SCAN_IN), .B(n4714), .Z(n4173) );
  XNOR2_X1 U4880 ( .A(n2194), .B(n4173), .ZN(n4172) );
  NAND2_X1 U4881 ( .A1(n4815), .A2(ADDR_REG_18__SCAN_IN), .ZN(n4150) );
  NAND2_X1 U4882 ( .A1(n4150), .A2(n4149), .ZN(n4169) );
  INV_X1 U4883 ( .A(REG2_REG_18__SCAN_IN), .ZN(n4152) );
  NOR2_X1 U4884 ( .A1(n4714), .A2(n4152), .ZN(n4151) );
  AOI21_X1 U4885 ( .B1(n4714), .B2(n4152), .A(n4151), .ZN(n4167) );
  AOI22_X1 U4886 ( .A1(n4165), .A2(REG2_REG_17__SCAN_IN), .B1(n4153), .B2(
        n4855), .ZN(n4812) );
  INV_X1 U4887 ( .A(n4154), .ZN(n4861) );
  OAI22_X1 U4888 ( .A1(n4157), .A2(n4156), .B1(REG2_REG_13__SCAN_IN), .B2(
        n4155), .ZN(n4158) );
  NOR2_X1 U4889 ( .A1(n4861), .A2(n4158), .ZN(n4159) );
  INV_X1 U4890 ( .A(REG2_REG_14__SCAN_IN), .ZN(n4783) );
  XNOR2_X1 U4891 ( .A(n4861), .B(n4158), .ZN(n4782) );
  NOR2_X1 U4892 ( .A1(n4783), .A2(n4782), .ZN(n4781) );
  NOR2_X1 U4893 ( .A1(n4159), .A2(n4781), .ZN(n4792) );
  NAND2_X1 U4894 ( .A1(REG2_REG_15__SCAN_IN), .A2(n4161), .ZN(n4160) );
  OAI21_X1 U4895 ( .B1(REG2_REG_15__SCAN_IN), .B2(n4161), .A(n4160), .ZN(n4791) );
  NOR2_X1 U4896 ( .A1(n4792), .A2(n4791), .ZN(n4790) );
  INV_X1 U4897 ( .A(n4162), .ZN(n4857) );
  NAND2_X1 U4898 ( .A1(n4163), .A2(n4857), .ZN(n4164) );
  NAND2_X1 U4899 ( .A1(n4812), .A2(n4810), .ZN(n4811) );
  AOI211_X1 U4900 ( .C1(n4167), .C2(n4166), .A(n4175), .B(n4809), .ZN(n4168)
         );
  AOI211_X1 U4901 ( .C1(n4170), .C2(n4714), .A(n4169), .B(n4168), .ZN(n4171)
         );
  OAI21_X1 U4902 ( .B1(n4184), .B2(n4172), .A(n4171), .ZN(U3258) );
  MUX2_X1 U4903 ( .A(REG1_REG_19__SCAN_IN), .B(n4566), .S(n4179), .Z(n4174) );
  INV_X1 U4904 ( .A(REG2_REG_19__SCAN_IN), .ZN(n4176) );
  MUX2_X1 U4905 ( .A(n4176), .B(REG2_REG_19__SCAN_IN), .S(n4179), .Z(n4177) );
  NAND2_X1 U4906 ( .A1(n4178), .A2(n4773), .ZN(n4183) );
  NOR2_X1 U4907 ( .A1(n4822), .A2(n4179), .ZN(n4180) );
  AOI211_X1 U4908 ( .C1(n4815), .C2(ADDR_REG_19__SCAN_IN), .A(n4181), .B(n4180), .ZN(n4182) );
  OAI211_X1 U4909 ( .C1(n4185), .C2(n4184), .A(n4183), .B(n4182), .ZN(U3259)
         );
  XNOR2_X1 U4910 ( .A(n4501), .B(n4188), .ZN(n4644) );
  NAND2_X1 U4911 ( .A1(n4187), .A2(n4186), .ZN(n4504) );
  OAI21_X1 U4912 ( .B1(n4188), .B2(n4876), .A(n4504), .ZN(n4641) );
  NAND2_X1 U4913 ( .A1(n4641), .A2(n4727), .ZN(n4190) );
  NAND2_X1 U4914 ( .A1(n4493), .A2(REG2_REG_31__SCAN_IN), .ZN(n4189) );
  OAI211_X1 U4915 ( .C1(n4644), .C2(n4488), .A(n4190), .B(n4189), .ZN(U3260)
         );
  INV_X1 U4916 ( .A(n4191), .ZN(n4198) );
  OAI22_X1 U4917 ( .A1(n4193), .A2(n4488), .B1(n4192), .B2(n4478), .ZN(n4194)
         );
  OAI21_X1 U4918 ( .B1(n4195), .B2(n4194), .A(n4727), .ZN(n4197) );
  NAND2_X1 U4919 ( .A1(n4493), .A2(REG2_REG_29__SCAN_IN), .ZN(n4196) );
  OAI211_X1 U4920 ( .C1(n4198), .C2(n4415), .A(n4197), .B(n4196), .ZN(U3354)
         );
  OAI21_X1 U4921 ( .B1(n4201), .B2(n4200), .A(n4199), .ZN(n4202) );
  NAND2_X1 U4922 ( .A1(n4202), .A2(n4491), .ZN(n4512) );
  XNOR2_X1 U4923 ( .A(n4204), .B(n4203), .ZN(n4515) );
  NAND2_X1 U4924 ( .A1(n4515), .A2(n4496), .ZN(n4214) );
  AND2_X1 U4925 ( .A1(n2183), .A2(n4509), .ZN(n4206) );
  OR2_X1 U4926 ( .A1(n4206), .A2(n4205), .ZN(n4651) );
  INV_X1 U4927 ( .A(n4651), .ZN(n4212) );
  AOI22_X1 U4928 ( .A1(n4825), .A2(REG2_REG_27__SCAN_IN), .B1(n4207), .B2(
        n4823), .ZN(n4208) );
  OAI21_X1 U4929 ( .B1(n4513), .B2(n4468), .A(n4208), .ZN(n4211) );
  OAI22_X1 U4930 ( .A1(n4238), .A2(n4484), .B1(n4209), .B2(n4483), .ZN(n4210)
         );
  AOI211_X1 U4931 ( .C1(n4212), .C2(n4828), .A(n4211), .B(n4210), .ZN(n4213)
         );
  OAI211_X1 U4932 ( .C1(n4493), .C2(n4512), .A(n4214), .B(n4213), .ZN(U3263)
         );
  XNOR2_X1 U4933 ( .A(n4216), .B(n4215), .ZN(n4523) );
  OAI21_X1 U4934 ( .B1(n2263), .B2(n4518), .A(n2183), .ZN(n4655) );
  INV_X1 U4935 ( .A(n4655), .ZN(n4231) );
  AOI22_X1 U4936 ( .A1(n4218), .A2(n4463), .B1(n4462), .B2(n4217), .ZN(n4222)
         );
  INV_X1 U4937 ( .A(n4219), .ZN(n4220) );
  AOI22_X1 U4938 ( .A1(n4825), .A2(REG2_REG_26__SCAN_IN), .B1(n4220), .B2(
        n4823), .ZN(n4221) );
  OAI211_X1 U4939 ( .C1(n4223), .C2(n4468), .A(n4222), .B(n4221), .ZN(n4230)
         );
  NAND2_X1 U4940 ( .A1(n4225), .A2(n4224), .ZN(n4227) );
  XNOR2_X1 U4941 ( .A(n4227), .B(n4226), .ZN(n4228) );
  NAND2_X1 U4942 ( .A1(n4228), .A2(n4491), .ZN(n4521) );
  NOR2_X1 U4943 ( .A1(n4521), .A2(n4493), .ZN(n4229) );
  AOI211_X1 U4944 ( .C1(n4231), .C2(n4828), .A(n4230), .B(n4229), .ZN(n4232)
         );
  OAI21_X1 U4945 ( .B1(n4523), .B2(n4415), .A(n4232), .ZN(U3264) );
  XNOR2_X1 U4946 ( .A(n4233), .B(n4237), .ZN(n4527) );
  INV_X1 U4947 ( .A(n4527), .ZN(n4249) );
  NAND2_X1 U4948 ( .A1(n4235), .A2(n4234), .ZN(n4236) );
  XOR2_X1 U4949 ( .A(n4237), .B(n4236), .Z(n4242) );
  OAI22_X1 U4950 ( .A1(n4238), .A2(n4878), .B1(n4876), .B2(n4244), .ZN(n4239)
         );
  AOI21_X1 U4951 ( .B1(n4881), .B2(n4240), .A(n4239), .ZN(n4241) );
  OAI21_X1 U4952 ( .B1(n4242), .B2(n4637), .A(n4241), .ZN(n4526) );
  OAI21_X1 U4953 ( .B1(n4252), .B2(n4244), .A(n4243), .ZN(n4658) );
  AOI22_X1 U4954 ( .A1(n4825), .A2(REG2_REG_25__SCAN_IN), .B1(n4245), .B2(
        n4823), .ZN(n4246) );
  OAI21_X1 U4955 ( .B1(n4658), .B2(n4488), .A(n4246), .ZN(n4247) );
  AOI21_X1 U4956 ( .B1(n4526), .B2(n4724), .A(n4247), .ZN(n4248) );
  OAI21_X1 U4957 ( .B1(n4249), .B2(n4415), .A(n4248), .ZN(U3265) );
  XNOR2_X1 U4958 ( .A(n4250), .B(n4251), .ZN(n4536) );
  INV_X1 U4959 ( .A(n4252), .ZN(n4253) );
  OAI21_X1 U4960 ( .B1(n4284), .B2(n4530), .A(n4253), .ZN(n4662) );
  INV_X1 U4961 ( .A(n4662), .ZN(n4265) );
  AOI22_X1 U4962 ( .A1(n4254), .A2(n4462), .B1(n4463), .B2(n4533), .ZN(n4257)
         );
  AOI22_X1 U4963 ( .A1(n4825), .A2(REG2_REG_24__SCAN_IN), .B1(n4255), .B2(
        n4823), .ZN(n4256) );
  OAI211_X1 U4964 ( .C1(n4531), .C2(n4468), .A(n4257), .B(n4256), .ZN(n4264)
         );
  NAND2_X1 U4965 ( .A1(n4259), .A2(n4258), .ZN(n4261) );
  XNOR2_X1 U4966 ( .A(n4261), .B(n4260), .ZN(n4262) );
  NAND2_X1 U4967 ( .A1(n4262), .A2(n4491), .ZN(n4534) );
  NOR2_X1 U4968 ( .A1(n4534), .A2(n4493), .ZN(n4263) );
  AOI211_X1 U4969 ( .C1(n4265), .C2(n4828), .A(n4264), .B(n4263), .ZN(n4266)
         );
  OAI21_X1 U4970 ( .B1(n4536), .B2(n4415), .A(n4266), .ZN(U3266) );
  XNOR2_X1 U4971 ( .A(n4267), .B(n4276), .ZN(n4541) );
  INV_X1 U4972 ( .A(n4541), .ZN(n4291) );
  OR2_X1 U4973 ( .A1(n4384), .A2(n4268), .ZN(n4270) );
  NAND2_X1 U4974 ( .A1(n4270), .A2(n4269), .ZN(n4325) );
  NAND2_X1 U4975 ( .A1(n4325), .A2(n4271), .ZN(n4273) );
  NAND2_X1 U4976 ( .A1(n4273), .A2(n4272), .ZN(n4311) );
  NAND2_X1 U4977 ( .A1(n4311), .A2(n4312), .ZN(n4310) );
  NAND2_X1 U4978 ( .A1(n4310), .A2(n4274), .ZN(n4292) );
  AOI21_X1 U4979 ( .B1(n4292), .B2(n4303), .A(n4275), .ZN(n4277) );
  XNOR2_X1 U4980 ( .A(n4277), .B(n4276), .ZN(n4282) );
  OAI22_X1 U4981 ( .A1(n4279), .A2(n4878), .B1(n4876), .B2(n4278), .ZN(n4280)
         );
  AOI21_X1 U4982 ( .B1(n4881), .B2(n4551), .A(n4280), .ZN(n4281) );
  OAI21_X1 U4983 ( .B1(n4282), .B2(n4637), .A(n4281), .ZN(n4540) );
  AND2_X1 U4984 ( .A1(n4300), .A2(n4283), .ZN(n4285) );
  OR2_X1 U4985 ( .A1(n4285), .A2(n4284), .ZN(n4665) );
  INV_X1 U4986 ( .A(n4286), .ZN(n4287) );
  AOI22_X1 U4987 ( .A1(n4825), .A2(REG2_REG_23__SCAN_IN), .B1(n4287), .B2(
        n4823), .ZN(n4288) );
  OAI21_X1 U4988 ( .B1(n4665), .B2(n4488), .A(n4288), .ZN(n4289) );
  AOI21_X1 U4989 ( .B1(n4540), .B2(n4724), .A(n4289), .ZN(n4290) );
  OAI21_X1 U4990 ( .B1(n4291), .B2(n4415), .A(n4290), .ZN(U3267) );
  XOR2_X1 U4991 ( .A(n4303), .B(n4292), .Z(n4297) );
  OAI22_X1 U4992 ( .A1(n4294), .A2(n4878), .B1(n4293), .B2(n4876), .ZN(n4295)
         );
  AOI21_X1 U4993 ( .B1(n4881), .B2(n4327), .A(n4295), .ZN(n4296) );
  OAI21_X1 U4994 ( .B1(n4297), .B2(n4637), .A(n4296), .ZN(n4545) );
  NAND2_X1 U4995 ( .A1(n2184), .A2(n4298), .ZN(n4299) );
  NAND2_X1 U4996 ( .A1(n4300), .A2(n4299), .ZN(n4669) );
  AOI22_X1 U4997 ( .A1(n4825), .A2(REG2_REG_22__SCAN_IN), .B1(n4301), .B2(
        n4823), .ZN(n4302) );
  OAI21_X1 U4998 ( .B1(n4669), .B2(n4488), .A(n4302), .ZN(n4307) );
  INV_X1 U4999 ( .A(n4546), .ZN(n4305) );
  AND2_X1 U5000 ( .A1(n4304), .A2(n4303), .ZN(n4544) );
  NOR3_X1 U5001 ( .A1(n4305), .A2(n4544), .A3(n4415), .ZN(n4306) );
  AOI211_X1 U5002 ( .C1(n4727), .C2(n4545), .A(n4307), .B(n4306), .ZN(n4308)
         );
  INV_X1 U5003 ( .A(n4308), .ZN(U3268) );
  XOR2_X1 U5004 ( .A(n4312), .B(n4309), .Z(n4556) );
  INV_X1 U5005 ( .A(n4556), .ZN(n4322) );
  OAI21_X1 U5006 ( .B1(n4312), .B2(n4311), .A(n4310), .ZN(n4313) );
  AND2_X1 U5007 ( .A1(n4313), .A2(n4491), .ZN(n4555) );
  OAI21_X1 U5008 ( .B1(n4334), .B2(n4314), .A(n2184), .ZN(n4673) );
  NOR2_X1 U5009 ( .A1(n4673), .A2(n4488), .ZN(n4320) );
  AOI22_X1 U5010 ( .A1(n4462), .A2(n4550), .B1(n4463), .B2(n4354), .ZN(n4317)
         );
  AOI22_X1 U5011 ( .A1(n4825), .A2(REG2_REG_21__SCAN_IN), .B1(n4315), .B2(
        n4823), .ZN(n4316) );
  OAI211_X1 U5012 ( .C1(n4318), .C2(n4468), .A(n4317), .B(n4316), .ZN(n4319)
         );
  AOI211_X1 U5013 ( .C1(n4555), .C2(n4727), .A(n4320), .B(n4319), .ZN(n4321)
         );
  OAI21_X1 U5014 ( .B1(n4322), .B2(n4415), .A(n4321), .ZN(U3269) );
  XNOR2_X1 U5015 ( .A(n4323), .B(n4324), .ZN(n4559) );
  XNOR2_X1 U5016 ( .A(n4325), .B(n4324), .ZN(n4331) );
  AOI22_X1 U5017 ( .A1(n4327), .A2(n4592), .B1(n4326), .B2(n4627), .ZN(n4328)
         );
  OAI21_X1 U5018 ( .B1(n4329), .B2(n4615), .A(n4328), .ZN(n4330) );
  AOI21_X1 U5019 ( .B1(n4331), .B2(n4491), .A(n4330), .ZN(n4332) );
  OAI21_X1 U5020 ( .B1(n4559), .B2(n4333), .A(n4332), .ZN(n4560) );
  NAND2_X1 U5021 ( .A1(n4560), .A2(n4727), .ZN(n4342) );
  INV_X1 U5022 ( .A(n4334), .ZN(n4335) );
  OAI21_X1 U5023 ( .B1(n4359), .B2(n4336), .A(n4335), .ZN(n4677) );
  INV_X1 U5024 ( .A(n4677), .ZN(n4340) );
  OAI22_X1 U5025 ( .A1(n4724), .A2(n4338), .B1(n4337), .B2(n4478), .ZN(n4339)
         );
  AOI21_X1 U5026 ( .B1(n4340), .B2(n4828), .A(n4339), .ZN(n4341) );
  OAI211_X1 U5027 ( .C1(n4559), .C2(n4343), .A(n4342), .B(n4341), .ZN(U3270)
         );
  XNOR2_X1 U5028 ( .A(n4344), .B(n4351), .ZN(n4565) );
  INV_X1 U5029 ( .A(n4565), .ZN(n4364) );
  INV_X1 U5030 ( .A(n4345), .ZN(n4347) );
  OAI21_X1 U5031 ( .B1(n4384), .B2(n4347), .A(n4346), .ZN(n4372) );
  INV_X1 U5032 ( .A(n4348), .ZN(n4350) );
  OAI21_X1 U5033 ( .B1(n4372), .B2(n4350), .A(n4349), .ZN(n4352) );
  XNOR2_X1 U5034 ( .A(n4352), .B(n4351), .ZN(n4353) );
  NAND2_X1 U5035 ( .A1(n4353), .A2(n4491), .ZN(n4356) );
  AOI22_X1 U5036 ( .A1(n4354), .A2(n4592), .B1(n4627), .B2(n2882), .ZN(n4355)
         );
  OAI211_X1 U5037 ( .C1(n4395), .C2(n4615), .A(n4356), .B(n4355), .ZN(n4564)
         );
  NOR2_X1 U5038 ( .A1(n4368), .A2(n4357), .ZN(n4358) );
  OR2_X1 U5039 ( .A1(n4359), .A2(n4358), .ZN(n4681) );
  NOR2_X1 U5040 ( .A1(n4681), .A2(n4488), .ZN(n4362) );
  OAI22_X1 U5041 ( .A1(n4724), .A2(n4176), .B1(n4360), .B2(n4478), .ZN(n4361)
         );
  AOI211_X1 U5042 ( .C1(n4564), .C2(n4724), .A(n4362), .B(n4361), .ZN(n4363)
         );
  OAI21_X1 U5043 ( .B1(n4364), .B2(n4415), .A(n4363), .ZN(U3271) );
  OAI21_X1 U5044 ( .B1(n4365), .B2(n4373), .A(n4366), .ZN(n4367) );
  INV_X1 U5045 ( .A(n4367), .ZN(n4570) );
  INV_X1 U5046 ( .A(n4389), .ZN(n4371) );
  INV_X1 U5047 ( .A(n4368), .ZN(n4369) );
  OAI211_X1 U5048 ( .C1(n4371), .C2(n4370), .A(n4369), .B(n4585), .ZN(n4568)
         );
  XOR2_X1 U5049 ( .A(n4373), .B(n4372), .Z(n4378) );
  AOI22_X1 U5050 ( .A1(n4375), .A2(n4592), .B1(n4374), .B2(n4627), .ZN(n4376)
         );
  OAI21_X1 U5051 ( .B1(n4409), .B2(n4615), .A(n4376), .ZN(n4377) );
  AOI21_X1 U5052 ( .B1(n4378), .B2(n4491), .A(n4377), .ZN(n4569) );
  OAI21_X1 U5053 ( .B1(n4379), .B2(n4568), .A(n4569), .ZN(n4382) );
  OAI22_X1 U5054 ( .A1(n4724), .A2(n4152), .B1(n4380), .B2(n4478), .ZN(n4381)
         );
  AOI21_X1 U5055 ( .B1(n4382), .B2(n4724), .A(n4381), .ZN(n4383) );
  OAI21_X1 U5056 ( .B1(n4570), .B2(n4415), .A(n4383), .ZN(U3272) );
  XNOR2_X1 U5057 ( .A(n4384), .B(n4387), .ZN(n4385) );
  NAND2_X1 U5058 ( .A1(n4385), .A2(n4491), .ZN(n4574) );
  XOR2_X1 U5059 ( .A(n4387), .B(n4386), .Z(n4577) );
  NAND2_X1 U5060 ( .A1(n4577), .A2(n4496), .ZN(n4399) );
  INV_X1 U5061 ( .A(n4388), .ZN(n4403) );
  OAI21_X1 U5062 ( .B1(n4403), .B2(n4390), .A(n4389), .ZN(n4686) );
  INV_X1 U5063 ( .A(n4686), .ZN(n4397) );
  AOI22_X1 U5064 ( .A1(n4463), .A2(n4593), .B1(n4462), .B2(n4571), .ZN(n4394)
         );
  INV_X1 U5065 ( .A(n4391), .ZN(n4392) );
  AOI22_X1 U5066 ( .A1(n4825), .A2(REG2_REG_17__SCAN_IN), .B1(n4392), .B2(
        n4823), .ZN(n4393) );
  OAI211_X1 U5067 ( .C1(n4395), .C2(n4468), .A(n4394), .B(n4393), .ZN(n4396)
         );
  AOI21_X1 U5068 ( .B1(n4397), .B2(n4828), .A(n4396), .ZN(n4398) );
  OAI211_X1 U5069 ( .C1(n4493), .C2(n4574), .A(n4399), .B(n4398), .ZN(U3273)
         );
  OAI21_X1 U5070 ( .B1(n4402), .B2(n4401), .A(n4400), .ZN(n4590) );
  AOI21_X1 U5071 ( .B1(n4580), .B2(n4421), .A(n4403), .ZN(n4586) );
  AOI22_X1 U5072 ( .A1(n4463), .A2(n4404), .B1(n4462), .B2(n4580), .ZN(n4408)
         );
  INV_X1 U5073 ( .A(n4405), .ZN(n4406) );
  AOI22_X1 U5074 ( .A1(n4493), .A2(REG2_REG_16__SCAN_IN), .B1(n4406), .B2(
        n4823), .ZN(n4407) );
  OAI211_X1 U5075 ( .C1(n4409), .C2(n4468), .A(n4408), .B(n4407), .ZN(n4413)
         );
  OAI211_X1 U5076 ( .C1(n4411), .C2(n2326), .A(n4410), .B(n4491), .ZN(n4587)
         );
  NOR2_X1 U5077 ( .A1(n4587), .A2(n4493), .ZN(n4412) );
  AOI211_X1 U5078 ( .C1(n4586), .C2(n4828), .A(n4413), .B(n4412), .ZN(n4414)
         );
  OAI21_X1 U5079 ( .B1(n4590), .B2(n4415), .A(n4414), .ZN(U3274) );
  AOI21_X1 U5080 ( .B1(n4416), .B2(n4419), .A(n4637), .ZN(n4418) );
  NAND2_X1 U5081 ( .A1(n4418), .A2(n4417), .ZN(n4595) );
  XNOR2_X1 U5082 ( .A(n4420), .B(n4419), .ZN(n4597) );
  NAND2_X1 U5083 ( .A1(n4597), .A2(n4496), .ZN(n4431) );
  OAI21_X1 U5084 ( .B1(n4441), .B2(n4422), .A(n4421), .ZN(n4691) );
  INV_X1 U5085 ( .A(n4691), .ZN(n4429) );
  AOI22_X1 U5086 ( .A1(n4463), .A2(n4423), .B1(n4462), .B2(n4591), .ZN(n4427)
         );
  INV_X1 U5087 ( .A(n4424), .ZN(n4425) );
  AOI22_X1 U5088 ( .A1(n4493), .A2(REG2_REG_15__SCAN_IN), .B1(n4425), .B2(
        n4823), .ZN(n4426) );
  OAI211_X1 U5089 ( .C1(n4575), .C2(n4468), .A(n4427), .B(n4426), .ZN(n4428)
         );
  AOI21_X1 U5090 ( .B1(n4429), .B2(n4828), .A(n4428), .ZN(n4430) );
  OAI211_X1 U5091 ( .C1(n4493), .C2(n4595), .A(n4431), .B(n4430), .ZN(U3275)
         );
  XNOR2_X1 U5092 ( .A(n4432), .B(n4434), .ZN(n4440) );
  OAI21_X1 U5093 ( .B1(n4435), .B2(n4434), .A(n4433), .ZN(n4601) );
  NAND2_X1 U5094 ( .A1(n4601), .A2(n4436), .ZN(n4439) );
  OAI22_X1 U5095 ( .A1(n4583), .A2(n4878), .B1(n4443), .B2(n4876), .ZN(n4437)
         );
  AOI21_X1 U5096 ( .B1(n4881), .B2(n4481), .A(n4437), .ZN(n4438) );
  OAI211_X1 U5097 ( .C1(n4637), .C2(n4440), .A(n4439), .B(n4438), .ZN(n4600)
         );
  INV_X1 U5098 ( .A(n4600), .ZN(n4448) );
  INV_X1 U5099 ( .A(n4441), .ZN(n4442) );
  OAI21_X1 U5100 ( .B1(n4459), .B2(n4443), .A(n4442), .ZN(n4695) );
  NOR2_X1 U5101 ( .A1(n4695), .A2(n4488), .ZN(n4446) );
  OAI22_X1 U5102 ( .A1(n4724), .A2(n4783), .B1(n4444), .B2(n4478), .ZN(n4445)
         );
  AOI211_X1 U5103 ( .C1(n4601), .C2(n4829), .A(n4446), .B(n4445), .ZN(n4447)
         );
  OAI21_X1 U5104 ( .B1(n4448), .B2(n4493), .A(n4447), .ZN(U3276) );
  INV_X1 U5105 ( .A(n4449), .ZN(n4450) );
  AOI21_X1 U5106 ( .B1(n4452), .B2(n4451), .A(n4450), .ZN(n4490) );
  INV_X1 U5107 ( .A(n4453), .ZN(n4454) );
  AOI21_X1 U5108 ( .B1(n4490), .B2(n4455), .A(n4454), .ZN(n4456) );
  XNOR2_X1 U5109 ( .A(n4456), .B(n4457), .ZN(n4609) );
  XNOR2_X1 U5110 ( .A(n4458), .B(n4457), .ZN(n4611) );
  NAND2_X1 U5111 ( .A1(n4611), .A2(n4496), .ZN(n4472) );
  INV_X1 U5112 ( .A(n4459), .ZN(n4460) );
  OAI21_X1 U5113 ( .B1(n2259), .B2(n4604), .A(n4460), .ZN(n4698) );
  INV_X1 U5114 ( .A(n4698), .ZN(n4470) );
  AOI22_X1 U5115 ( .A1(n4463), .A2(n4607), .B1(n4462), .B2(n4461), .ZN(n4467)
         );
  INV_X1 U5116 ( .A(n4464), .ZN(n4465) );
  AOI22_X1 U5117 ( .A1(n4825), .A2(REG2_REG_13__SCAN_IN), .B1(n4465), .B2(
        n4823), .ZN(n4466) );
  OAI211_X1 U5118 ( .C1(n4605), .C2(n4468), .A(n4467), .B(n4466), .ZN(n4469)
         );
  AOI21_X1 U5119 ( .B1(n4470), .B2(n4828), .A(n4469), .ZN(n4471) );
  OAI211_X1 U5120 ( .C1(n4609), .C2(n4473), .A(n4472), .B(n4471), .ZN(U3277)
         );
  XNOR2_X1 U5121 ( .A(n4474), .B(n4489), .ZN(n4621) );
  NAND2_X1 U5122 ( .A1(n2215), .A2(n4475), .ZN(n4476) );
  NAND2_X1 U5123 ( .A1(n4477), .A2(n4476), .ZN(n4702) );
  OAI22_X1 U5124 ( .A1(n4727), .A2(n3178), .B1(n4479), .B2(n4478), .ZN(n4480)
         );
  AOI21_X1 U5125 ( .B1(n4482), .B2(n4481), .A(n4480), .ZN(n4487) );
  OAI22_X1 U5126 ( .A1(n4616), .A2(n4484), .B1(n4483), .B2(n4613), .ZN(n4485)
         );
  INV_X1 U5127 ( .A(n4485), .ZN(n4486) );
  OAI211_X1 U5128 ( .C1(n4702), .C2(n4488), .A(n4487), .B(n4486), .ZN(n4495)
         );
  XNOR2_X1 U5129 ( .A(n4490), .B(n4489), .ZN(n4492) );
  NAND2_X1 U5130 ( .A1(n4492), .A2(n4491), .ZN(n4620) );
  NOR2_X1 U5131 ( .A1(n4620), .A2(n4493), .ZN(n4494) );
  AOI211_X1 U5132 ( .C1(n4496), .C2(n4621), .A(n4495), .B(n4494), .ZN(n4497)
         );
  INV_X1 U5133 ( .A(n4497), .ZN(U3278) );
  NOR2_X1 U5134 ( .A1(n4920), .A2(n4498), .ZN(n4499) );
  AOI21_X1 U5135 ( .B1(n4641), .B2(n4920), .A(n4499), .ZN(n4500) );
  OAI21_X1 U5136 ( .B1(n4644), .B2(n4640), .A(n4500), .ZN(U3549) );
  AOI21_X1 U5137 ( .B1(n4503), .B2(n4502), .A(n4501), .ZN(n4725) );
  NAND2_X1 U5138 ( .A1(n4725), .A2(n4912), .ZN(n4507) );
  OAI21_X1 U5139 ( .B1(n4505), .B2(n4876), .A(n4504), .ZN(n4723) );
  NAND2_X1 U5140 ( .A1(n4723), .A2(n4920), .ZN(n4506) );
  OAI211_X1 U5141 ( .C1(n4920), .C2(n3242), .A(n4507), .B(n4506), .ZN(U3548)
         );
  MUX2_X1 U5142 ( .A(REG1_REG_28__SCAN_IN), .B(n4508), .S(n4920), .Z(U3546) );
  AOI22_X1 U5143 ( .A1(n4510), .A2(n4881), .B1(n4509), .B2(n4627), .ZN(n4511)
         );
  OAI211_X1 U5144 ( .C1(n4513), .C2(n4878), .A(n4512), .B(n4511), .ZN(n4514)
         );
  AOI21_X1 U5145 ( .B1(n4515), .B2(n4895), .A(n4514), .ZN(n4648) );
  MUX2_X1 U5146 ( .A(n4516), .B(n4648), .S(n4920), .Z(n4517) );
  OAI21_X1 U5147 ( .B1(n4640), .B2(n4651), .A(n4517), .ZN(U3545) );
  OAI22_X1 U5148 ( .A1(n4531), .A2(n4615), .B1(n4518), .B2(n4876), .ZN(n4519)
         );
  AOI21_X1 U5149 ( .B1(n4592), .B2(n4520), .A(n4519), .ZN(n4522) );
  OAI211_X1 U5150 ( .C1(n4523), .C2(n4589), .A(n4522), .B(n4521), .ZN(n4652)
         );
  MUX2_X1 U5151 ( .A(REG1_REG_26__SCAN_IN), .B(n4652), .S(n4920), .Z(n4524) );
  INV_X1 U5152 ( .A(n4524), .ZN(n4525) );
  OAI21_X1 U5153 ( .B1(n4640), .B2(n4655), .A(n4525), .ZN(U3544) );
  AOI21_X1 U5154 ( .B1(n4527), .B2(n4895), .A(n4526), .ZN(n4656) );
  MUX2_X1 U5155 ( .A(n4528), .B(n4656), .S(n4920), .Z(n4529) );
  OAI21_X1 U5156 ( .B1(n4640), .B2(n4658), .A(n4529), .ZN(U3543) );
  OAI22_X1 U5157 ( .A1(n4531), .A2(n4878), .B1(n4876), .B2(n4530), .ZN(n4532)
         );
  AOI21_X1 U5158 ( .B1(n4881), .B2(n4533), .A(n4532), .ZN(n4535) );
  OAI211_X1 U5159 ( .C1(n4536), .C2(n4589), .A(n4535), .B(n4534), .ZN(n4537)
         );
  INV_X1 U5160 ( .A(n4537), .ZN(n4659) );
  MUX2_X1 U5161 ( .A(n4538), .B(n4659), .S(n4920), .Z(n4539) );
  OAI21_X1 U5162 ( .B1(n4640), .B2(n4662), .A(n4539), .ZN(U3542) );
  AOI21_X1 U5163 ( .B1(n4541), .B2(n4895), .A(n4540), .ZN(n4663) );
  MUX2_X1 U5164 ( .A(n4542), .B(n4663), .S(n4920), .Z(n4543) );
  OAI21_X1 U5165 ( .B1(n4640), .B2(n4665), .A(n4543), .ZN(U3541) );
  NOR2_X1 U5166 ( .A1(n4544), .A2(n4589), .ZN(n4547) );
  AOI21_X1 U5167 ( .B1(n4547), .B2(n4546), .A(n4545), .ZN(n4666) );
  MUX2_X1 U5168 ( .A(n4548), .B(n4666), .S(n4920), .Z(n4549) );
  OAI21_X1 U5169 ( .B1(n4640), .B2(n4669), .A(n4549), .ZN(U3540) );
  AOI22_X1 U5170 ( .A1(n4551), .A2(n4592), .B1(n4627), .B2(n4550), .ZN(n4552)
         );
  OAI21_X1 U5171 ( .B1(n4553), .B2(n4615), .A(n4552), .ZN(n4554) );
  AOI211_X1 U5172 ( .C1(n4556), .C2(n4895), .A(n4555), .B(n4554), .ZN(n4670)
         );
  MUX2_X1 U5173 ( .A(n4557), .B(n4670), .S(n4920), .Z(n4558) );
  OAI21_X1 U5174 ( .B1(n4640), .B2(n4673), .A(n4558), .ZN(U3539) );
  INV_X1 U5175 ( .A(n4559), .ZN(n4561) );
  AOI21_X1 U5176 ( .B1(n4908), .B2(n4561), .A(n4560), .ZN(n4674) );
  MUX2_X1 U5177 ( .A(n4562), .B(n4674), .S(n4920), .Z(n4563) );
  OAI21_X1 U5178 ( .B1(n4640), .B2(n4677), .A(n4563), .ZN(U3538) );
  AOI21_X1 U5179 ( .B1(n4565), .B2(n4895), .A(n4564), .ZN(n4678) );
  MUX2_X1 U5180 ( .A(n4566), .B(n4678), .S(n4920), .Z(n4567) );
  OAI21_X1 U5181 ( .B1(n4640), .B2(n4681), .A(n4567), .ZN(U3537) );
  OAI211_X1 U5182 ( .C1(n4570), .C2(n4589), .A(n4569), .B(n4568), .ZN(n4682)
         );
  MUX2_X1 U5183 ( .A(REG1_REG_18__SCAN_IN), .B(n4682), .S(n4920), .Z(U3536) );
  AOI22_X1 U5184 ( .A1(n4572), .A2(n4592), .B1(n4627), .B2(n4571), .ZN(n4573)
         );
  OAI211_X1 U5185 ( .C1(n4575), .C2(n4615), .A(n4574), .B(n4573), .ZN(n4576)
         );
  AOI21_X1 U5186 ( .B1(n4577), .B2(n4895), .A(n4576), .ZN(n4683) );
  MUX2_X1 U5187 ( .A(n4578), .B(n4683), .S(n4920), .Z(n4579) );
  OAI21_X1 U5188 ( .B1(n4640), .B2(n4686), .A(n4579), .ZN(U3535) );
  AOI22_X1 U5189 ( .A1(n4581), .A2(n4592), .B1(n4580), .B2(n4627), .ZN(n4582)
         );
  OAI21_X1 U5190 ( .B1(n4583), .B2(n4615), .A(n4582), .ZN(n4584) );
  AOI21_X1 U5191 ( .B1(n4586), .B2(n4585), .A(n4584), .ZN(n4588) );
  OAI211_X1 U5192 ( .C1(n4590), .C2(n4589), .A(n4588), .B(n4587), .ZN(n4687)
         );
  MUX2_X1 U5193 ( .A(REG1_REG_16__SCAN_IN), .B(n4687), .S(n4920), .Z(U3534) );
  AOI22_X1 U5194 ( .A1(n4593), .A2(n4592), .B1(n4627), .B2(n4591), .ZN(n4594)
         );
  OAI211_X1 U5195 ( .C1(n4605), .C2(n4615), .A(n4595), .B(n4594), .ZN(n4596)
         );
  AOI21_X1 U5196 ( .B1(n4597), .B2(n4895), .A(n4596), .ZN(n4688) );
  MUX2_X1 U5197 ( .A(n4598), .B(n4688), .S(n4920), .Z(n4599) );
  OAI21_X1 U5198 ( .B1(n4640), .B2(n4691), .A(n4599), .ZN(U3533) );
  AOI21_X1 U5199 ( .B1(n4908), .B2(n4601), .A(n4600), .ZN(n4692) );
  MUX2_X1 U5200 ( .A(n4602), .B(n4692), .S(n4920), .Z(n4603) );
  OAI21_X1 U5201 ( .B1(n4640), .B2(n4695), .A(n4603), .ZN(U3532) );
  OAI22_X1 U5202 ( .A1(n4605), .A2(n4878), .B1(n4876), .B2(n4604), .ZN(n4606)
         );
  AOI21_X1 U5203 ( .B1(n4881), .B2(n4607), .A(n4606), .ZN(n4608) );
  OAI21_X1 U5204 ( .B1(n4609), .B2(n4637), .A(n4608), .ZN(n4610) );
  AOI21_X1 U5205 ( .B1(n4895), .B2(n4611), .A(n4610), .ZN(n4696) );
  MUX2_X1 U5206 ( .A(n4142), .B(n4696), .S(n4920), .Z(n4612) );
  OAI21_X1 U5207 ( .B1(n4640), .B2(n4698), .A(n4612), .ZN(U3531) );
  OAI22_X1 U5208 ( .A1(n4614), .A2(n4878), .B1(n4876), .B2(n4613), .ZN(n4618)
         );
  NOR2_X1 U5209 ( .A1(n4616), .A2(n4615), .ZN(n4617) );
  NOR2_X1 U5210 ( .A1(n4618), .A2(n4617), .ZN(n4619) );
  AND2_X1 U5211 ( .A1(n4620), .A2(n4619), .ZN(n4623) );
  NAND2_X1 U5212 ( .A1(n4621), .A2(n4895), .ZN(n4622) );
  NAND2_X1 U5213 ( .A1(n4623), .A2(n4622), .ZN(n4699) );
  MUX2_X1 U5214 ( .A(REG1_REG_12__SCAN_IN), .B(n4699), .S(n4920), .Z(n4624) );
  INV_X1 U5215 ( .A(n4624), .ZN(n4625) );
  OAI21_X1 U5216 ( .B1(n4640), .B2(n4702), .A(n4625), .ZN(U3530) );
  NAND2_X1 U5217 ( .A1(n4626), .A2(n4895), .ZN(n4635) );
  NAND2_X1 U5218 ( .A1(n4628), .A2(n4627), .ZN(n4631) );
  NAND2_X1 U5219 ( .A1(n4629), .A2(n4881), .ZN(n4630) );
  OAI211_X1 U5220 ( .C1(n4632), .C2(n4878), .A(n4631), .B(n4630), .ZN(n4633)
         );
  INV_X1 U5221 ( .A(n4633), .ZN(n4634) );
  OAI211_X1 U5222 ( .C1(n4637), .C2(n4636), .A(n4635), .B(n4634), .ZN(n4703)
         );
  MUX2_X1 U5223 ( .A(REG1_REG_11__SCAN_IN), .B(n4703), .S(n4920), .Z(n4638) );
  INV_X1 U5224 ( .A(n4638), .ZN(n4639) );
  OAI21_X1 U5225 ( .B1(n4640), .B2(n4707), .A(n4639), .ZN(U3529) );
  NAND2_X1 U5226 ( .A1(n4641), .A2(n4910), .ZN(n4643) );
  NAND2_X1 U5227 ( .A1(n3250), .A2(REG0_REG_31__SCAN_IN), .ZN(n4642) );
  OAI211_X1 U5228 ( .C1(n4644), .C2(n4706), .A(n4643), .B(n4642), .ZN(U3517)
         );
  NAND2_X1 U5229 ( .A1(n4725), .A2(n4886), .ZN(n4646) );
  NAND2_X1 U5230 ( .A1(n4723), .A2(n4910), .ZN(n4645) );
  OAI211_X1 U5231 ( .C1(n4910), .C2(n4647), .A(n4646), .B(n4645), .ZN(U3516)
         );
  INV_X1 U5232 ( .A(REG0_REG_27__SCAN_IN), .ZN(n4649) );
  MUX2_X1 U5233 ( .A(n4649), .B(n4648), .S(n4910), .Z(n4650) );
  OAI21_X1 U5234 ( .B1(n4651), .B2(n4706), .A(n4650), .ZN(U3513) );
  MUX2_X1 U5235 ( .A(REG0_REG_26__SCAN_IN), .B(n4652), .S(n4910), .Z(n4653) );
  INV_X1 U5236 ( .A(n4653), .ZN(n4654) );
  OAI21_X1 U5237 ( .B1(n4655), .B2(n4706), .A(n4654), .ZN(U3512) );
  MUX2_X1 U5238 ( .A(n3028), .B(n4656), .S(n4910), .Z(n4657) );
  OAI21_X1 U5239 ( .B1(n4658), .B2(n4706), .A(n4657), .ZN(U3511) );
  INV_X1 U5240 ( .A(REG0_REG_24__SCAN_IN), .ZN(n4660) );
  MUX2_X1 U5241 ( .A(n4660), .B(n4659), .S(n4910), .Z(n4661) );
  OAI21_X1 U5242 ( .B1(n4662), .B2(n4706), .A(n4661), .ZN(U3510) );
  MUX2_X1 U5243 ( .A(n3020), .B(n4663), .S(n4910), .Z(n4664) );
  OAI21_X1 U5244 ( .B1(n4665), .B2(n4706), .A(n4664), .ZN(U3509) );
  MUX2_X1 U5245 ( .A(n4667), .B(n4666), .S(n4910), .Z(n4668) );
  OAI21_X1 U5246 ( .B1(n4669), .B2(n4706), .A(n4668), .ZN(U3508) );
  INV_X1 U5247 ( .A(REG0_REG_21__SCAN_IN), .ZN(n4671) );
  MUX2_X1 U5248 ( .A(n4671), .B(n4670), .S(n4910), .Z(n4672) );
  OAI21_X1 U5249 ( .B1(n4673), .B2(n4706), .A(n4672), .ZN(U3507) );
  INV_X1 U5250 ( .A(REG0_REG_20__SCAN_IN), .ZN(n4675) );
  MUX2_X1 U5251 ( .A(n4675), .B(n4674), .S(n4910), .Z(n4676) );
  OAI21_X1 U5252 ( .B1(n4677), .B2(n4706), .A(n4676), .ZN(U3506) );
  INV_X1 U5253 ( .A(REG0_REG_19__SCAN_IN), .ZN(n4679) );
  MUX2_X1 U5254 ( .A(n4679), .B(n4678), .S(n4910), .Z(n4680) );
  OAI21_X1 U5255 ( .B1(n4681), .B2(n4706), .A(n4680), .ZN(U3505) );
  MUX2_X1 U5256 ( .A(REG0_REG_18__SCAN_IN), .B(n4682), .S(n4910), .Z(U3503) );
  INV_X1 U5257 ( .A(REG0_REG_17__SCAN_IN), .ZN(n4684) );
  MUX2_X1 U5258 ( .A(n4684), .B(n4683), .S(n4910), .Z(n4685) );
  OAI21_X1 U5259 ( .B1(n4686), .B2(n4706), .A(n4685), .ZN(U3501) );
  MUX2_X1 U5260 ( .A(REG0_REG_16__SCAN_IN), .B(n4687), .S(n4910), .Z(U3499) );
  INV_X1 U5261 ( .A(REG0_REG_15__SCAN_IN), .ZN(n4689) );
  MUX2_X1 U5262 ( .A(n4689), .B(n4688), .S(n4910), .Z(n4690) );
  OAI21_X1 U5263 ( .B1(n4691), .B2(n4706), .A(n4690), .ZN(U3497) );
  INV_X1 U5264 ( .A(REG0_REG_14__SCAN_IN), .ZN(n4693) );
  MUX2_X1 U5265 ( .A(n4693), .B(n4692), .S(n4910), .Z(n4694) );
  OAI21_X1 U5266 ( .B1(n4695), .B2(n4706), .A(n4694), .ZN(U3495) );
  MUX2_X1 U5267 ( .A(n3167), .B(n4696), .S(n4910), .Z(n4697) );
  OAI21_X1 U5268 ( .B1(n4698), .B2(n4706), .A(n4697), .ZN(U3493) );
  MUX2_X1 U5269 ( .A(REG0_REG_12__SCAN_IN), .B(n4699), .S(n4910), .Z(n4700) );
  INV_X1 U5270 ( .A(n4700), .ZN(n4701) );
  OAI21_X1 U5271 ( .B1(n4702), .B2(n4706), .A(n4701), .ZN(U3491) );
  MUX2_X1 U5272 ( .A(n4703), .B(REG0_REG_11__SCAN_IN), .S(n3250), .Z(n4704) );
  INV_X1 U5273 ( .A(n4704), .ZN(n4705) );
  OAI21_X1 U5274 ( .B1(n4707), .B2(n4706), .A(n4705), .ZN(U3489) );
  MUX2_X1 U5275 ( .A(n4708), .B(DATAI_29_), .S(U3149), .Z(U3323) );
  MUX2_X1 U5276 ( .A(n4709), .B(DATAI_27_), .S(U3149), .Z(U3325) );
  MUX2_X1 U5277 ( .A(n4710), .B(DATAI_26_), .S(U3149), .Z(U3326) );
  MUX2_X1 U5278 ( .A(n4711), .B(DATAI_24_), .S(U3149), .Z(U3328) );
  MUX2_X1 U5279 ( .A(n4712), .B(DATAI_22_), .S(U3149), .Z(U3330) );
  MUX2_X1 U5280 ( .A(DATAI_20_), .B(n4713), .S(STATE_REG_SCAN_IN), .Z(U3332)
         );
  MUX2_X1 U5281 ( .A(n4714), .B(DATAI_18_), .S(U3149), .Z(U3334) );
  MUX2_X1 U5282 ( .A(DATAI_7_), .B(n4715), .S(STATE_REG_SCAN_IN), .Z(U3345) );
  MUX2_X1 U5283 ( .A(DATAI_6_), .B(n4716), .S(STATE_REG_SCAN_IN), .Z(U3346) );
  MUX2_X1 U5284 ( .A(n4717), .B(DATAI_4_), .S(U3149), .Z(U3348) );
  MUX2_X1 U5285 ( .A(n4718), .B(DATAI_3_), .S(U3149), .Z(U3349) );
  MUX2_X1 U5286 ( .A(DATAI_2_), .B(n4719), .S(STATE_REG_SCAN_IN), .Z(U3350) );
  MUX2_X1 U5287 ( .A(n4720), .B(DATAI_1_), .S(U3149), .Z(U3351) );
  AOI22_X1 U5288 ( .A1(STATE_REG_SCAN_IN), .A2(n4722), .B1(n4721), .B2(U3149), 
        .ZN(U3324) );
  AOI22_X1 U5289 ( .A1(n4725), .A2(n4828), .B1(n4724), .B2(n4723), .ZN(n4726)
         );
  OAI21_X1 U5290 ( .B1(n4728), .B2(n4727), .A(n4726), .ZN(U3261) );
  OAI211_X1 U5291 ( .C1(REG2_REG_8__SCAN_IN), .C2(n4730), .A(n4773), .B(n4729), 
        .ZN(n4731) );
  NAND2_X1 U5292 ( .A1(n4732), .A2(n4731), .ZN(n4733) );
  AOI21_X1 U5293 ( .B1(n4815), .B2(ADDR_REG_8__SCAN_IN), .A(n4733), .ZN(n4737)
         );
  OAI211_X1 U5294 ( .C1(REG1_REG_8__SCAN_IN), .C2(n4735), .A(n4816), .B(n4734), 
        .ZN(n4736) );
  OAI211_X1 U5295 ( .C1(n4822), .C2(n4870), .A(n4737), .B(n4736), .ZN(U3248)
         );
  OAI211_X1 U5296 ( .C1(n4740), .C2(n4739), .A(n4816), .B(n4738), .ZN(n4745)
         );
  OAI211_X1 U5297 ( .C1(n4743), .C2(n4742), .A(n4773), .B(n4741), .ZN(n4744)
         );
  OAI211_X1 U5298 ( .C1(n4822), .C2(n4868), .A(n4745), .B(n4744), .ZN(n4746)
         );
  AOI211_X1 U5299 ( .C1(n4815), .C2(ADDR_REG_9__SCAN_IN), .A(n4747), .B(n4746), 
        .ZN(n4748) );
  INV_X1 U5300 ( .A(n4748), .ZN(U3249) );
  OAI211_X1 U5301 ( .C1(REG2_REG_10__SCAN_IN), .C2(n4751), .A(n4773), .B(n4750), .ZN(n4753) );
  NAND2_X1 U5302 ( .A1(n4753), .A2(n4752), .ZN(n4754) );
  AOI21_X1 U5303 ( .B1(n4815), .B2(ADDR_REG_10__SCAN_IN), .A(n4754), .ZN(n4758) );
  OAI211_X1 U5304 ( .C1(REG1_REG_10__SCAN_IN), .C2(n4756), .A(n4816), .B(n4755), .ZN(n4757) );
  OAI211_X1 U5305 ( .C1(n4822), .C2(n2270), .A(n4758), .B(n4757), .ZN(U3250)
         );
  OAI211_X1 U5306 ( .C1(n4761), .C2(n4760), .A(n4816), .B(n4759), .ZN(n4766)
         );
  OAI211_X1 U5307 ( .C1(n4764), .C2(n4763), .A(n4773), .B(n4762), .ZN(n4765)
         );
  OAI211_X1 U5308 ( .C1(n4822), .C2(n4865), .A(n4766), .B(n4765), .ZN(n4767)
         );
  AOI211_X1 U5309 ( .C1(n4815), .C2(ADDR_REG_11__SCAN_IN), .A(n4768), .B(n4767), .ZN(n4769) );
  INV_X1 U5310 ( .A(n4769), .ZN(U3251) );
  OAI211_X1 U5311 ( .C1(REG1_REG_12__SCAN_IN), .C2(n4771), .A(n4816), .B(n4770), .ZN(n4776) );
  OAI211_X1 U5312 ( .C1(REG2_REG_12__SCAN_IN), .C2(n4774), .A(n4773), .B(n4772), .ZN(n4775) );
  OAI211_X1 U5313 ( .C1(n4822), .C2(n4863), .A(n4776), .B(n4775), .ZN(n4777)
         );
  AOI211_X1 U5314 ( .C1(n4815), .C2(ADDR_REG_12__SCAN_IN), .A(n4778), .B(n4777), .ZN(n4779) );
  INV_X1 U5315 ( .A(n4779), .ZN(U3252) );
  INV_X1 U5316 ( .A(n4780), .ZN(n4785) );
  AOI211_X1 U5317 ( .C1(n4783), .C2(n4782), .A(n4781), .B(n4809), .ZN(n4784)
         );
  AOI211_X1 U5318 ( .C1(ADDR_REG_14__SCAN_IN), .C2(n4815), .A(n4785), .B(n4784), .ZN(n4789) );
  OAI211_X1 U5319 ( .C1(REG1_REG_14__SCAN_IN), .C2(n4787), .A(n4816), .B(n4786), .ZN(n4788) );
  OAI211_X1 U5320 ( .C1(n4822), .C2(n4861), .A(n4789), .B(n4788), .ZN(U3254)
         );
  AOI211_X1 U5321 ( .C1(n4792), .C2(n4791), .A(n4790), .B(n4809), .ZN(n4793)
         );
  AOI211_X1 U5322 ( .C1(n4815), .C2(ADDR_REG_15__SCAN_IN), .A(n4794), .B(n4793), .ZN(n4799) );
  OAI211_X1 U5323 ( .C1(n4797), .C2(n4796), .A(n4816), .B(n4795), .ZN(n4798)
         );
  OAI211_X1 U5324 ( .C1(n4822), .C2(n4859), .A(n4799), .B(n4798), .ZN(U3255)
         );
  AOI221_X1 U5325 ( .B1(n4802), .B2(n4801), .C1(n4800), .C2(n4801), .A(n4809), 
        .ZN(n4803) );
  AOI211_X1 U5326 ( .C1(n4815), .C2(ADDR_REG_16__SCAN_IN), .A(n4804), .B(n4803), .ZN(n4808) );
  OAI221_X1 U5327 ( .B1(n4806), .B2(REG1_REG_16__SCAN_IN), .C1(n4806), .C2(
        n4805), .A(n4816), .ZN(n4807) );
  OAI211_X1 U5328 ( .C1(n4822), .C2(n4857), .A(n4808), .B(n4807), .ZN(U3256)
         );
  AOI221_X1 U5329 ( .B1(n4812), .B2(n4811), .C1(n4810), .C2(n4811), .A(n4809), 
        .ZN(n4813) );
  AOI211_X1 U5330 ( .C1(ADDR_REG_17__SCAN_IN), .C2(n4815), .A(n4814), .B(n4813), .ZN(n4821) );
  OAI221_X1 U5331 ( .B1(n4819), .B2(n4818), .C1(n4819), .C2(n4817), .A(n4816), 
        .ZN(n4820) );
  OAI211_X1 U5332 ( .C1(n4822), .C2(n4855), .A(n4821), .B(n4820), .ZN(U3257)
         );
  AOI22_X1 U5333 ( .A1(n4825), .A2(REG2_REG_8__SCAN_IN), .B1(n4824), .B2(n4823), .ZN(n4832) );
  INV_X1 U5334 ( .A(n4826), .ZN(n4827) );
  AOI22_X1 U5335 ( .A1(n4830), .A2(n4829), .B1(n4828), .B2(n4827), .ZN(n4831)
         );
  OAI211_X1 U5336 ( .C1(n4493), .C2(n4833), .A(n4832), .B(n4831), .ZN(U3282)
         );
  AND2_X1 U5337 ( .A1(D_REG_31__SCAN_IN), .A2(n4847), .ZN(U3291) );
  NOR2_X1 U5338 ( .A1(n4852), .A2(n4834), .ZN(U3292) );
  AND2_X1 U5339 ( .A1(D_REG_29__SCAN_IN), .A2(n4847), .ZN(U3293) );
  AND2_X1 U5340 ( .A1(D_REG_28__SCAN_IN), .A2(n4847), .ZN(U3294) );
  NOR2_X1 U5341 ( .A1(n4852), .A2(n4835), .ZN(U3295) );
  NOR2_X1 U5342 ( .A1(n4852), .A2(n4836), .ZN(U3296) );
  AND2_X1 U5343 ( .A1(D_REG_25__SCAN_IN), .A2(n4847), .ZN(U3297) );
  AND2_X1 U5344 ( .A1(D_REG_24__SCAN_IN), .A2(n4847), .ZN(U3298) );
  NOR2_X1 U5345 ( .A1(n4852), .A2(n4837), .ZN(U3299) );
  AND2_X1 U5346 ( .A1(D_REG_22__SCAN_IN), .A2(n4847), .ZN(U3300) );
  AND2_X1 U5347 ( .A1(D_REG_21__SCAN_IN), .A2(n4847), .ZN(U3301) );
  NOR2_X1 U5348 ( .A1(n4852), .A2(n4838), .ZN(U3302) );
  NOR2_X1 U5349 ( .A1(n4852), .A2(n4839), .ZN(U3303) );
  AND2_X1 U5350 ( .A1(D_REG_18__SCAN_IN), .A2(n4847), .ZN(U3304) );
  NOR2_X1 U5351 ( .A1(n4852), .A2(n4840), .ZN(U3305) );
  NOR2_X1 U5352 ( .A1(n4852), .A2(n4841), .ZN(U3306) );
  NOR2_X1 U5353 ( .A1(n4852), .A2(n4842), .ZN(U3307) );
  NOR2_X1 U5354 ( .A1(n4852), .A2(n4843), .ZN(U3308) );
  AND2_X1 U5355 ( .A1(D_REG_13__SCAN_IN), .A2(n4847), .ZN(U3309) );
  NOR2_X1 U5356 ( .A1(n4852), .A2(n4844), .ZN(U3310) );
  NOR2_X1 U5357 ( .A1(n4852), .A2(n4845), .ZN(U3311) );
  NOR2_X1 U5358 ( .A1(n4852), .A2(n4846), .ZN(U3312) );
  AND2_X1 U5359 ( .A1(D_REG_9__SCAN_IN), .A2(n4847), .ZN(U3313) );
  AND2_X1 U5360 ( .A1(D_REG_8__SCAN_IN), .A2(n4847), .ZN(U3314) );
  AND2_X1 U5361 ( .A1(D_REG_7__SCAN_IN), .A2(n4847), .ZN(U3315) );
  AND2_X1 U5362 ( .A1(D_REG_6__SCAN_IN), .A2(n4847), .ZN(U3316) );
  NOR2_X1 U5363 ( .A1(n4852), .A2(n4848), .ZN(U3317) );
  NOR2_X1 U5364 ( .A1(n4852), .A2(n4849), .ZN(U3318) );
  NOR2_X1 U5365 ( .A1(n4852), .A2(n4850), .ZN(U3319) );
  NOR2_X1 U5366 ( .A1(n4852), .A2(n4851), .ZN(U3320) );
  AOI21_X1 U5367 ( .B1(U3149), .B2(n4854), .A(n4853), .ZN(U3329) );
  AOI22_X1 U5368 ( .A1(STATE_REG_SCAN_IN), .A2(n4855), .B1(n2660), .B2(U3149), 
        .ZN(U3335) );
  AOI22_X1 U5369 ( .A1(STATE_REG_SCAN_IN), .A2(n4857), .B1(n4856), .B2(U3149), 
        .ZN(U3336) );
  INV_X1 U5370 ( .A(DATAI_15_), .ZN(n4858) );
  AOI22_X1 U5371 ( .A1(STATE_REG_SCAN_IN), .A2(n4859), .B1(n4858), .B2(U3149), 
        .ZN(U3337) );
  INV_X1 U5372 ( .A(DATAI_14_), .ZN(n4860) );
  AOI22_X1 U5373 ( .A1(STATE_REG_SCAN_IN), .A2(n4861), .B1(n4860), .B2(U3149), 
        .ZN(U3338) );
  AOI22_X1 U5374 ( .A1(STATE_REG_SCAN_IN), .A2(n4863), .B1(n4862), .B2(U3149), 
        .ZN(U3340) );
  INV_X1 U5375 ( .A(DATAI_11_), .ZN(n4864) );
  AOI22_X1 U5376 ( .A1(STATE_REG_SCAN_IN), .A2(n4865), .B1(n4864), .B2(U3149), 
        .ZN(U3341) );
  INV_X1 U5377 ( .A(DATAI_10_), .ZN(n4866) );
  AOI22_X1 U5378 ( .A1(STATE_REG_SCAN_IN), .A2(n2270), .B1(n4866), .B2(U3149), 
        .ZN(U3342) );
  INV_X1 U5379 ( .A(DATAI_9_), .ZN(n4867) );
  AOI22_X1 U5380 ( .A1(STATE_REG_SCAN_IN), .A2(n4868), .B1(n4867), .B2(U3149), 
        .ZN(U3343) );
  AOI22_X1 U5381 ( .A1(STATE_REG_SCAN_IN), .A2(n4870), .B1(n4869), .B2(U3149), 
        .ZN(U3344) );
  INV_X1 U5382 ( .A(DATAI_0_), .ZN(n4871) );
  AOI22_X1 U5383 ( .A1(STATE_REG_SCAN_IN), .A2(n2225), .B1(n4871), .B2(U3149), 
        .ZN(U3352) );
  INV_X1 U5384 ( .A(REG0_REG_0__SCAN_IN), .ZN(n4872) );
  AOI22_X1 U5385 ( .A1(n4910), .A2(n4873), .B1(n4872), .B2(n3250), .ZN(U3467)
         );
  INV_X1 U5386 ( .A(REG0_REG_1__SCAN_IN), .ZN(n4874) );
  AOI22_X1 U5387 ( .A1(n4910), .A2(n4875), .B1(n4874), .B2(n3250), .ZN(U3469)
         );
  OAI22_X1 U5388 ( .A1(n4879), .A2(n4878), .B1(n4877), .B2(n4876), .ZN(n4880)
         );
  AOI21_X1 U5389 ( .B1(n4881), .B2(n3375), .A(n4880), .ZN(n4882) );
  OAI211_X1 U5390 ( .C1(n4885), .C2(n4884), .A(n4883), .B(n4882), .ZN(n4913)
         );
  AOI22_X1 U5391 ( .A1(n4913), .A2(n4910), .B1(n4886), .B2(n4911), .ZN(n4887)
         );
  OAI21_X1 U5392 ( .B1(n4910), .B2(n4888), .A(n4887), .ZN(U3471) );
  INV_X1 U5393 ( .A(n4889), .ZN(n4893) );
  INV_X1 U5394 ( .A(n4890), .ZN(n4892) );
  AOI211_X1 U5395 ( .C1(n4893), .C2(n4908), .A(n4892), .B(n4891), .ZN(n4916)
         );
  INV_X1 U5396 ( .A(REG0_REG_4__SCAN_IN), .ZN(n4894) );
  AOI22_X1 U5397 ( .A1(n4910), .A2(n4916), .B1(n4894), .B2(n3250), .ZN(U3475)
         );
  NAND3_X1 U5398 ( .A1(n4897), .A2(n4896), .A3(n4895), .ZN(n4898) );
  AND3_X1 U5399 ( .A1(n4900), .A2(n4899), .A3(n4898), .ZN(n4917) );
  AOI22_X1 U5400 ( .A1(n4910), .A2(n4917), .B1(n4901), .B2(n3250), .ZN(U3481)
         );
  NOR3_X1 U5401 ( .A1(n4904), .A2(n4903), .A3(n4902), .ZN(n4906) );
  AOI211_X1 U5402 ( .C1(n4908), .C2(n4907), .A(n4906), .B(n4905), .ZN(n4919)
         );
  AOI22_X1 U5403 ( .A1(n4910), .A2(n4919), .B1(n4909), .B2(n3250), .ZN(U3487)
         );
  AOI22_X1 U5404 ( .A1(n4913), .A2(n4920), .B1(n4912), .B2(n4911), .ZN(n4914)
         );
  OAI21_X1 U5405 ( .B1(n4920), .B2(n4915), .A(n4914), .ZN(U3520) );
  AOI22_X1 U5406 ( .A1(n4920), .A2(n4916), .B1(n2459), .B2(n4918), .ZN(U3522)
         );
  AOI22_X1 U5407 ( .A1(n4920), .A2(n4917), .B1(n3385), .B2(n4918), .ZN(U3525)
         );
  AOI22_X1 U5408 ( .A1(n4920), .A2(n4919), .B1(n2550), .B2(n4918), .ZN(U3528)
         );
  CLKBUF_X1 U2435 ( .A(n2406), .Z(n2799) );
  CLKBUF_X1 U2588 ( .A(n2549), .Z(n3305) );
endmodule

