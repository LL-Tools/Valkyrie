

module b22_C_AntiSAT_k_256_6 ( P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, 
        keyinput128, keyinput129, keyinput130, keyinput131, keyinput132, 
        keyinput133, keyinput134, keyinput135, keyinput136, keyinput137, 
        keyinput138, keyinput139, keyinput140, keyinput141, keyinput142, 
        keyinput143, keyinput144, keyinput145, keyinput146, keyinput147, 
        keyinput148, keyinput149, keyinput150, keyinput151, keyinput152, 
        keyinput153, keyinput154, keyinput155, keyinput156, keyinput157, 
        keyinput158, keyinput159, keyinput160, keyinput161, keyinput162, 
        keyinput163, keyinput164, keyinput165, keyinput166, keyinput167, 
        keyinput168, keyinput169, keyinput170, keyinput171, keyinput172, 
        keyinput173, keyinput174, keyinput175, keyinput176, keyinput177, 
        keyinput178, keyinput179, keyinput180, keyinput181, keyinput182, 
        keyinput183, keyinput184, keyinput185, keyinput186, keyinput187, 
        keyinput188, keyinput189, keyinput190, keyinput191, keyinput192, 
        keyinput193, keyinput194, keyinput195, keyinput196, keyinput197, 
        keyinput198, keyinput199, keyinput200, keyinput201, keyinput202, 
        keyinput203, keyinput204, keyinput205, keyinput206, keyinput207, 
        keyinput208, keyinput209, keyinput210, keyinput211, keyinput212, 
        keyinput213, keyinput214, keyinput215, keyinput216, keyinput217, 
        keyinput218, keyinput219, keyinput220, keyinput221, keyinput222, 
        keyinput223, keyinput224, keyinput225, keyinput226, keyinput227, 
        keyinput228, keyinput229, keyinput230, keyinput231, keyinput232, 
        keyinput233, keyinput234, keyinput235, keyinput236, keyinput237, 
        keyinput238, keyinput239, keyinput240, keyinput241, keyinput242, 
        keyinput243, keyinput244, keyinput245, keyinput246, keyinput247, 
        keyinput248, keyinput249, keyinput250, keyinput251, keyinput252, 
        keyinput253, keyinput254, keyinput255, SUB_1596_U4, SUB_1596_U62, 
        SUB_1596_U63, SUB_1596_U64, SUB_1596_U65, SUB_1596_U66, SUB_1596_U67, 
        SUB_1596_U68, SUB_1596_U69, SUB_1596_U70, SUB_1596_U54, SUB_1596_U55, 
        SUB_1596_U56, SUB_1596_U57, SUB_1596_U58, SUB_1596_U59, SUB_1596_U60, 
        SUB_1596_U61, SUB_1596_U5, SUB_1596_U53, U29, U28, P1_U3355, P1_U3354, 
        P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, P1_U3347, 
        P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, P1_U3340, 
        P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, P1_U3333, 
        P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, P1_U3326, 
        P1_U3325, P1_U3324, P1_U3445, P1_U3446, P1_U3323, P1_U3322, P1_U3321, 
        P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, P1_U3314, 
        P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, P1_U3307, 
        P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, P1_U3300, 
        P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, P1_U3459, 
        P1_U3462, P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, 
        P1_U3483, P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, 
        P1_U3504, P1_U3507, P1_U3510, P1_U3513, P1_U3515, P1_U3516, P1_U3517, 
        P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, P1_U3524, 
        P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, P1_U3531, 
        P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, P1_U3538, 
        P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, P1_U3545, 
        P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, P1_U3552, 
        P1_U3553, P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, 
        P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, P1_U3288, P1_U3287, 
        P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, P1_U3280, 
        P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, P1_U3273, 
        P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, P1_U3266, 
        P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, P1_U3261, P1_U3260, 
        P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, P1_U3253, 
        P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, P1_U3246, 
        P1_U3245, P1_U3244, P1_U3243, P1_U3560, P1_U3561, P1_U3562, P1_U3563, 
        P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, P1_U3570, 
        P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, P1_U3577, 
        P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, P1_U3584, 
        P1_U3585, P1_U3586, P1_U3587, P1_U3588, P1_U3589, P1_U3590, P1_U3591, 
        P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, P1_U3237, P1_U3236, 
        P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, P1_U3229, 
        P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, 
        P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, 
        P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U4016, P2_U3327, P2_U3326, 
        P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321, P2_U3320, P2_U3319, 
        P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314, P2_U3313, P2_U3312, 
        P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307, P2_U3306, P2_U3305, 
        P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300, P2_U3299, P2_U3298, 
        P2_U3297, P2_U3296, P2_U3416, P2_U3417, P2_U3295, P2_U3294, P2_U3293, 
        P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, 
        P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, 
        P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, 
        P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3430, 
        P2_U3433, P2_U3436, P2_U3439, P2_U3442, P2_U3445, P2_U3448, P2_U3451, 
        P2_U3454, P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, 
        P2_U3475, P2_U3478, P2_U3481, P2_U3484, P2_U3486, P2_U3487, P2_U3488, 
        P2_U3489, P2_U3490, P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, 
        P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, 
        P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, 
        P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, 
        P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, 
        P2_U3524, P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, 
        P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, 
        P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, 
        P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, 
        P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, 
        P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, 
        P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, 
        P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, 
        P2_U3216, P2_U3215, P2_U3214, P2_U3531, P2_U3532, P2_U3533, P2_U3534, 
        P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540, P2_U3541, 
        P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547, P2_U3548, 
        P2_U3549, P2_U3550, P2_U3551, P2_U3552, P2_U3553, P2_U3554, P2_U3555, 
        P2_U3556, P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, 
        P2_U3328, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3088, P2_U3087, P2_U3947, P3_U3295, P3_U3294, 
        P3_U3293, P3_U3292, P3_U3291, P3_U3290, P3_U3289, P3_U3288, P3_U3287, 
        P3_U3286, P3_U3285, P3_U3284, P3_U3283, P3_U3282, P3_U3281, P3_U3280, 
        P3_U3279, P3_U3278, P3_U3277, P3_U3276, P3_U3275, P3_U3274, P3_U3273, 
        P3_U3272, P3_U3271, P3_U3270, P3_U3269, P3_U3268, P3_U3267, P3_U3266, 
        P3_U3265, P3_U3264, P3_U3376, P3_U3377, P3_U3263, P3_U3262, P3_U3261, 
        P3_U3260, P3_U3259, P3_U3258, P3_U3257, P3_U3256, P3_U3255, P3_U3254, 
        P3_U3253, P3_U3252, P3_U3251, P3_U3250, P3_U3249, P3_U3248, P3_U3247, 
        P3_U3246, P3_U3245, P3_U3244, P3_U3243, P3_U3242, P3_U3241, P3_U3240, 
        P3_U3239, P3_U3238, P3_U3237, P3_U3236, P3_U3235, P3_U3234, P3_U3390, 
        P3_U3393, P3_U3396, P3_U3399, P3_U3402, P3_U3405, P3_U3408, P3_U3411, 
        P3_U3414, P3_U3417, P3_U3420, P3_U3423, P3_U3426, P3_U3429, P3_U3432, 
        P3_U3435, P3_U3438, P3_U3441, P3_U3444, P3_U3446, P3_U3447, P3_U3448, 
        P3_U3449, P3_U3450, P3_U3451, P3_U3452, P3_U3453, P3_U3454, P3_U3455, 
        P3_U3456, P3_U3457, P3_U3458, P3_U3459, P3_U3460, P3_U3461, P3_U3462, 
        P3_U3463, P3_U3464, P3_U3465, P3_U3466, P3_U3467, P3_U3468, P3_U3469, 
        P3_U3470, P3_U3471, P3_U3472, P3_U3473, P3_U3474, P3_U3475, P3_U3476, 
        P3_U3477, P3_U3478, P3_U3479, P3_U3480, P3_U3481, P3_U3482, P3_U3483, 
        P3_U3484, P3_U3485, P3_U3486, P3_U3487, P3_U3488, P3_U3489, P3_U3490, 
        P3_U3233, P3_U3232, P3_U3231, P3_U3230, P3_U3229, P3_U3228, P3_U3227, 
        P3_U3226, P3_U3225, P3_U3224, P3_U3223, P3_U3222, P3_U3221, P3_U3220, 
        P3_U3219, P3_U3218, P3_U3217, P3_U3216, P3_U3215, P3_U3214, P3_U3213, 
        P3_U3212, P3_U3211, P3_U3210, P3_U3209, P3_U3208, P3_U3207, P3_U3206, 
        P3_U3205, P3_U3204, P3_U3203, P3_U3202, P3_U3201, P3_U3200, P3_U3199, 
        P3_U3198, P3_U3197, P3_U3196, P3_U3195, P3_U3194, P3_U3193, P3_U3192, 
        P3_U3191, P3_U3190, P3_U3189, P3_U3188, P3_U3187, P3_U3186, P3_U3185, 
        P3_U3184, P3_U3183, P3_U3182, P3_U3491, P3_U3492, P3_U3493, P3_U3494, 
        P3_U3495, P3_U3496, P3_U3497, P3_U3498, P3_U3499, P3_U3500, P3_U3501, 
        P3_U3502, P3_U3503, P3_U3504, P3_U3505, P3_U3506, P3_U3507, P3_U3508, 
        P3_U3509, P3_U3510, P3_U3511, P3_U3512, P3_U3513, P3_U3514, P3_U3515, 
        P3_U3516, P3_U3517, P3_U3518, P3_U3519, P3_U3520, P3_U3521, P3_U3522, 
        P3_U3296, P3_U3181, P3_U3180, P3_U3179, P3_U3178, P3_U3177, P3_U3176, 
        P3_U3175, P3_U3174, P3_U3173, P3_U3172, P3_U3171, P3_U3170, P3_U3169, 
        P3_U3168, P3_U3167, P3_U3166, P3_U3165, P3_U3164, P3_U3163, P3_U3162, 
        P3_U3161, P3_U3160, P3_U3159, P3_U3158, P3_U3157, P3_U3156, P3_U3155, 
        P3_U3154, P3_U3153, P3_U3151, P3_U3150, P3_U3897 );
  input P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput0,
         keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6,
         keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12,
         keyinput13, keyinput14, keyinput15, keyinput16, keyinput17,
         keyinput18, keyinput19, keyinput20, keyinput21, keyinput22,
         keyinput23, keyinput24, keyinput25, keyinput26, keyinput27,
         keyinput28, keyinput29, keyinput30, keyinput31, keyinput32,
         keyinput33, keyinput34, keyinput35, keyinput36, keyinput37,
         keyinput38, keyinput39, keyinput40, keyinput41, keyinput42,
         keyinput43, keyinput44, keyinput45, keyinput46, keyinput47,
         keyinput48, keyinput49, keyinput50, keyinput51, keyinput52,
         keyinput53, keyinput54, keyinput55, keyinput56, keyinput57,
         keyinput58, keyinput59, keyinput60, keyinput61, keyinput62,
         keyinput63, keyinput64, keyinput65, keyinput66, keyinput67,
         keyinput68, keyinput69, keyinput70, keyinput71, keyinput72,
         keyinput73, keyinput74, keyinput75, keyinput76, keyinput77,
         keyinput78, keyinput79, keyinput80, keyinput81, keyinput82,
         keyinput83, keyinput84, keyinput85, keyinput86, keyinput87,
         keyinput88, keyinput89, keyinput90, keyinput91, keyinput92,
         keyinput93, keyinput94, keyinput95, keyinput96, keyinput97,
         keyinput98, keyinput99, keyinput100, keyinput101, keyinput102,
         keyinput103, keyinput104, keyinput105, keyinput106, keyinput107,
         keyinput108, keyinput109, keyinput110, keyinput111, keyinput112,
         keyinput113, keyinput114, keyinput115, keyinput116, keyinput117,
         keyinput118, keyinput119, keyinput120, keyinput121, keyinput122,
         keyinput123, keyinput124, keyinput125, keyinput126, keyinput127,
         keyinput128, keyinput129, keyinput130, keyinput131, keyinput132,
         keyinput133, keyinput134, keyinput135, keyinput136, keyinput137,
         keyinput138, keyinput139, keyinput140, keyinput141, keyinput142,
         keyinput143, keyinput144, keyinput145, keyinput146, keyinput147,
         keyinput148, keyinput149, keyinput150, keyinput151, keyinput152,
         keyinput153, keyinput154, keyinput155, keyinput156, keyinput157,
         keyinput158, keyinput159, keyinput160, keyinput161, keyinput162,
         keyinput163, keyinput164, keyinput165, keyinput166, keyinput167,
         keyinput168, keyinput169, keyinput170, keyinput171, keyinput172,
         keyinput173, keyinput174, keyinput175, keyinput176, keyinput177,
         keyinput178, keyinput179, keyinput180, keyinput181, keyinput182,
         keyinput183, keyinput184, keyinput185, keyinput186, keyinput187,
         keyinput188, keyinput189, keyinput190, keyinput191, keyinput192,
         keyinput193, keyinput194, keyinput195, keyinput196, keyinput197,
         keyinput198, keyinput199, keyinput200, keyinput201, keyinput202,
         keyinput203, keyinput204, keyinput205, keyinput206, keyinput207,
         keyinput208, keyinput209, keyinput210, keyinput211, keyinput212,
         keyinput213, keyinput214, keyinput215, keyinput216, keyinput217,
         keyinput218, keyinput219, keyinput220, keyinput221, keyinput222,
         keyinput223, keyinput224, keyinput225, keyinput226, keyinput227,
         keyinput228, keyinput229, keyinput230, keyinput231, keyinput232,
         keyinput233, keyinput234, keyinput235, keyinput236, keyinput237,
         keyinput238, keyinput239, keyinput240, keyinput241, keyinput242,
         keyinput243, keyinput244, keyinput245, keyinput246, keyinput247,
         keyinput248, keyinput249, keyinput250, keyinput251, keyinput252,
         keyinput253, keyinput254, keyinput255;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626,
         n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636,
         n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646,
         n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656,
         n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666,
         n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676,
         n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686,
         n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696,
         n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706,
         n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716,
         n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726,
         n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736,
         n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746,
         n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756,
         n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766,
         n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776,
         n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786,
         n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796,
         n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806,
         n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816,
         n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826,
         n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836,
         n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846,
         n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856,
         n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866,
         n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876,
         n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886,
         n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896,
         n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906,
         n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916,
         n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926,
         n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936,
         n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946,
         n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956,
         n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966,
         n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976,
         n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986,
         n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996,
         n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006,
         n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016,
         n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026,
         n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036,
         n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046,
         n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056,
         n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066,
         n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076,
         n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086,
         n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096,
         n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106,
         n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116,
         n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126,
         n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136,
         n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146,
         n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156,
         n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166,
         n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176,
         n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186,
         n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196,
         n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206,
         n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216,
         n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226,
         n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236,
         n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246,
         n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256,
         n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266,
         n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276,
         n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286,
         n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296,
         n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306,
         n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316,
         n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326,
         n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336,
         n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346,
         n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356,
         n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366,
         n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376,
         n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386,
         n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396,
         n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406,
         n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416,
         n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426,
         n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436,
         n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446,
         n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456,
         n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466,
         n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476,
         n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486,
         n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496,
         n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506,
         n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516,
         n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526,
         n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536,
         n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546,
         n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556,
         n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566,
         n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576,
         n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586,
         n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596,
         n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606,
         n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616,
         n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626,
         n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636,
         n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646,
         n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656,
         n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666,
         n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676,
         n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686,
         n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696,
         n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706,
         n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716,
         n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726,
         n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736,
         n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746,
         n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756,
         n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766,
         n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776,
         n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786,
         n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796,
         n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806,
         n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816,
         n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826,
         n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836,
         n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846,
         n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856,
         n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866,
         n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876,
         n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886,
         n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896,
         n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906,
         n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916,
         n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926,
         n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936,
         n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946,
         n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956,
         n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966,
         n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976,
         n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986,
         n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996,
         n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006,
         n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016,
         n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026,
         n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036,
         n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046,
         n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056,
         n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066,
         n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076,
         n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086,
         n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096,
         n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106,
         n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116,
         n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126,
         n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136,
         n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146,
         n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156,
         n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166,
         n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176,
         n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186,
         n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196,
         n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206,
         n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216,
         n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226,
         n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236,
         n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246,
         n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256,
         n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266,
         n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276,
         n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286,
         n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296,
         n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306,
         n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316,
         n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326,
         n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336,
         n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346,
         n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356,
         n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366,
         n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376,
         n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386,
         n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396,
         n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406,
         n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416,
         n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426,
         n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436,
         n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446,
         n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456,
         n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466,
         n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476,
         n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486,
         n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496,
         n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506,
         n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516,
         n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526,
         n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536,
         n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546,
         n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556,
         n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566,
         n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576,
         n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586,
         n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596,
         n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606,
         n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616,
         n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626,
         n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636,
         n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646,
         n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656,
         n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666,
         n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676,
         n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686,
         n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696,
         n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706,
         n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716,
         n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726,
         n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736,
         n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746,
         n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756,
         n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766,
         n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776,
         n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786,
         n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796,
         n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806,
         n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816,
         n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826,
         n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836,
         n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846,
         n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856,
         n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866,
         n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876,
         n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886,
         n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896,
         n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906,
         n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916,
         n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926,
         n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936,
         n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946,
         n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956,
         n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966,
         n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976,
         n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986,
         n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996,
         n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006,
         n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016,
         n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026,
         n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036,
         n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046,
         n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056,
         n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066,
         n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076,
         n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086,
         n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096,
         n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106,
         n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116,
         n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126,
         n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136,
         n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146,
         n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156,
         n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166,
         n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176,
         n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186,
         n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196,
         n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206,
         n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216,
         n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226,
         n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236,
         n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246,
         n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256,
         n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266,
         n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276,
         n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286,
         n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296,
         n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306,
         n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316,
         n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326,
         n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336,
         n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346,
         n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356,
         n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366,
         n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376,
         n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386,
         n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396,
         n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406,
         n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416,
         n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426,
         n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436,
         n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446,
         n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456,
         n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466,
         n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476,
         n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486,
         n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496,
         n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506,
         n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516,
         n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526,
         n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536,
         n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546,
         n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556,
         n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566,
         n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576,
         n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586,
         n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596,
         n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606,
         n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616,
         n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626,
         n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636,
         n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646,
         n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656,
         n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666,
         n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676,
         n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686,
         n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696,
         n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706,
         n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716,
         n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726,
         n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736,
         n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746,
         n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756,
         n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766,
         n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776,
         n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786,
         n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796,
         n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806,
         n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816,
         n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826,
         n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836,
         n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846,
         n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856,
         n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866,
         n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876,
         n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886,
         n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896,
         n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906,
         n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916,
         n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926,
         n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936,
         n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946,
         n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956,
         n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966,
         n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976,
         n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986,
         n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996,
         n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005,
         n10006, n10007, n10008, n10009, n10010, n10011, n10012, n10013,
         n10014, n10015, n10016, n10017, n10018, n10019, n10020, n10021,
         n10022, n10023, n10024, n10025, n10026, n10027, n10028, n10029,
         n10030, n10031, n10032, n10033, n10034, n10035, n10036, n10037,
         n10038, n10039, n10040, n10041, n10042, n10043, n10044, n10045,
         n10046, n10047, n10048, n10049, n10050, n10051, n10052, n10053,
         n10054, n10055, n10056, n10057, n10058, n10059, n10060, n10061,
         n10062, n10063, n10064, n10065, n10066, n10067, n10068, n10069,
         n10070, n10071, n10072, n10073, n10074, n10075, n10076, n10077,
         n10078, n10079, n10080, n10081, n10082, n10083, n10084, n10085,
         n10086, n10087, n10088, n10089, n10090, n10091, n10092, n10093,
         n10094, n10095, n10096, n10097, n10098, n10099, n10100, n10101,
         n10102, n10103, n10104, n10105, n10106, n10107, n10108, n10109,
         n10110, n10111, n10112, n10113, n10114, n10115, n10116, n10117,
         n10118, n10119, n10120, n10121, n10122, n10123, n10124, n10125,
         n10126, n10127, n10128, n10129, n10130, n10131, n10132, n10133,
         n10134, n10135, n10136, n10137, n10138, n10139, n10140, n10141,
         n10142, n10143, n10144, n10145, n10146, n10147, n10148, n10149,
         n10150, n10151, n10152, n10153, n10154, n10155, n10156, n10157,
         n10158, n10159, n10160, n10161, n10162, n10163, n10164, n10165,
         n10166, n10167, n10168, n10169, n10170, n10171, n10172, n10173,
         n10174, n10175, n10176, n10177, n10178, n10179, n10180, n10181,
         n10182, n10183, n10184, n10185, n10186, n10187, n10188, n10189,
         n10190, n10191, n10192, n10193, n10194, n10195, n10196, n10197,
         n10198, n10199, n10200, n10201, n10202, n10203, n10204, n10205,
         n10206, n10207, n10208, n10209, n10210, n10211, n10212, n10213,
         n10214, n10215, n10216, n10217, n10218, n10219, n10220, n10221,
         n10222, n10223, n10224, n10225, n10226, n10227, n10228, n10229,
         n10230, n10231, n10232, n10233, n10234, n10235, n10236, n10237,
         n10238, n10239, n10240, n10241, n10242, n10243, n10244, n10245,
         n10246, n10247, n10248, n10249, n10250, n10251, n10252, n10253,
         n10254, n10255, n10256, n10257, n10258, n10259, n10260, n10261,
         n10262, n10263, n10264, n10265, n10266, n10267, n10268, n10269,
         n10270, n10271, n10272, n10273, n10274, n10275, n10276, n10277,
         n10278, n10279, n10280, n10281, n10282, n10283, n10284, n10285,
         n10286, n10287, n10288, n10289, n10290, n10291, n10292, n10293,
         n10294, n10295, n10296, n10297, n10298, n10299, n10300, n10301,
         n10302, n10303, n10304, n10305, n10306, n10307, n10308, n10309,
         n10310, n10311, n10312, n10313, n10314, n10315, n10316, n10317,
         n10318, n10319, n10320, n10321, n10322, n10323, n10324, n10325,
         n10326, n10327, n10328, n10329, n10330, n10331, n10332, n10333,
         n10334, n10335, n10336, n10337, n10338, n10339, n10340, n10341,
         n10342, n10343, n10344, n10345, n10346, n10347, n10348, n10349,
         n10350, n10351, n10352, n10353, n10354, n10355, n10356, n10357,
         n10358, n10359, n10360, n10361, n10362, n10363, n10364, n10365,
         n10366, n10367, n10368, n10369, n10370, n10371, n10372, n10373,
         n10374, n10375, n10376, n10377, n10378, n10379, n10380, n10381,
         n10382, n10383, n10384, n10385, n10386, n10387, n10388, n10389,
         n10390, n10391, n10392, n10393, n10394, n10395, n10396, n10397,
         n10398, n10399, n10400, n10401, n10402, n10403, n10404, n10405,
         n10406, n10407, n10408, n10409, n10410, n10411, n10412, n10413,
         n10414, n10415, n10416, n10417, n10418, n10419, n10420, n10421,
         n10422, n10423, n10424, n10425, n10426, n10427, n10428, n10429,
         n10430, n10431, n10432, n10433, n10434, n10435, n10436, n10437,
         n10438, n10439, n10440, n10441, n10442, n10443, n10444, n10445,
         n10446, n10447, n10448, n10449, n10450, n10451, n10452, n10453,
         n10454, n10455, n10456, n10457, n10458, n10459, n10460, n10461,
         n10462, n10463, n10464, n10465, n10466, n10467, n10468, n10469,
         n10470, n10471, n10472, n10473, n10474, n10475, n10476, n10477,
         n10478, n10479, n10480, n10481, n10482, n10483, n10484, n10485,
         n10486, n10487, n10488, n10489, n10490, n10491, n10492, n10493,
         n10494, n10495, n10496, n10497, n10498, n10499, n10500, n10501,
         n10502, n10503, n10504, n10505, n10506, n10507, n10508, n10509,
         n10510, n10511, n10512, n10513, n10514, n10515, n10516, n10517,
         n10518, n10519, n10520, n10521, n10522, n10523, n10524, n10525,
         n10526, n10527, n10528, n10529, n10530, n10531, n10532, n10533,
         n10534, n10535, n10536, n10537, n10538, n10539, n10540, n10541,
         n10542, n10543, n10544, n10545, n10546, n10547, n10548, n10549,
         n10550, n10551, n10552, n10553, n10554, n10555, n10556, n10557,
         n10558, n10559, n10560, n10561, n10562, n10563, n10564, n10565,
         n10566, n10567, n10568, n10569, n10570, n10571, n10572, n10573,
         n10574, n10575, n10576, n10577, n10578, n10579, n10580, n10581,
         n10582, n10583, n10584, n10585, n10586, n10587, n10588, n10589,
         n10590, n10591, n10592, n10593, n10594, n10595, n10596, n10597,
         n10598, n10599, n10600, n10601, n10602, n10603, n10604, n10605,
         n10606, n10607, n10608, n10609, n10610, n10611, n10612, n10613,
         n10614, n10615, n10616, n10617, n10618, n10619, n10620, n10621,
         n10622, n10623, n10624, n10625, n10626, n10627, n10628, n10629,
         n10630, n10631, n10632, n10633, n10634, n10635, n10636, n10637,
         n10638, n10639, n10640, n10641, n10642, n10643, n10644, n10645,
         n10646, n10647, n10648, n10649, n10650, n10651, n10652, n10653,
         n10654, n10655, n10656, n10657, n10658, n10659, n10660, n10661,
         n10662, n10663, n10664, n10665, n10666, n10667, n10668, n10669,
         n10670, n10671, n10672, n10673, n10674, n10675, n10676, n10677,
         n10678, n10679, n10680, n10681, n10682, n10683, n10684, n10685,
         n10686, n10687, n10688, n10689, n10690, n10691, n10692, n10693,
         n10694, n10695, n10696, n10697, n10698, n10699, n10700, n10701,
         n10702, n10703, n10704, n10705, n10706, n10707, n10708, n10709,
         n10710, n10711, n10712, n10713, n10714, n10715, n10716, n10717,
         n10718, n10719, n10720, n10721, n10722, n10723, n10724, n10725,
         n10726, n10727, n10728, n10729, n10730, n10731, n10732, n10733,
         n10734, n10735, n10736, n10737, n10738, n10739, n10740, n10741,
         n10742, n10743, n10744, n10745, n10746, n10747, n10748, n10749,
         n10750, n10751, n10752, n10753, n10754, n10755, n10756, n10757,
         n10758, n10759, n10760, n10761, n10762, n10763, n10764, n10765,
         n10766, n10767, n10768, n10769, n10770, n10771, n10772, n10773,
         n10774, n10775, n10776, n10777, n10778, n10779, n10780, n10781,
         n10782, n10783, n10784, n10785, n10786, n10787, n10788, n10789,
         n10790, n10791, n10792, n10793, n10794, n10795, n10796, n10797,
         n10798, n10799, n10800, n10801, n10802, n10803, n10804, n10805,
         n10806, n10807, n10808, n10809, n10810, n10811, n10812, n10813,
         n10814, n10815, n10816, n10817, n10818, n10819, n10820, n10821,
         n10822, n10823, n10824, n10825, n10826, n10827, n10828, n10829,
         n10830, n10831, n10832, n10833, n10834, n10835, n10836, n10837,
         n10838, n10839, n10840, n10841, n10842, n10843, n10844, n10845,
         n10846, n10847, n10848, n10849, n10850, n10851, n10852, n10853,
         n10854, n10855, n10856, n10857, n10858, n10859, n10860, n10861,
         n10862, n10863, n10864, n10865, n10866, n10867, n10868, n10869,
         n10870, n10871, n10872, n10873, n10874, n10875, n10876, n10877,
         n10878, n10879, n10880, n10881, n10882, n10883, n10884, n10885,
         n10886, n10887, n10888, n10889, n10890, n10891, n10892, n10893,
         n10894, n10895, n10896, n10897, n10898, n10899, n10900, n10901,
         n10902, n10903, n10904, n10905, n10906, n10907, n10908, n10909,
         n10910, n10911, n10912, n10913, n10914, n10915, n10916, n10917,
         n10918, n10919, n10920, n10921, n10922, n10923, n10924, n10925,
         n10926, n10927, n10928, n10929, n10930, n10931, n10932, n10933,
         n10934, n10935, n10936, n10937, n10938, n10939, n10940, n10941,
         n10942, n10943, n10944, n10945, n10946, n10947, n10948, n10949,
         n10950, n10951, n10952, n10953, n10954, n10955, n10956, n10957,
         n10958, n10959, n10960, n10961, n10962, n10963, n10964, n10965,
         n10966, n10967, n10968, n10969, n10970, n10971, n10972, n10973,
         n10974, n10975, n10976, n10977, n10978, n10979, n10980, n10981,
         n10982, n10983, n10984, n10985, n10986, n10987, n10988, n10989,
         n10990, n10991, n10992, n10993, n10994, n10995, n10996, n10997,
         n10998, n10999, n11000, n11001, n11002, n11003, n11004, n11005,
         n11006, n11007, n11008, n11009, n11010, n11011, n11012, n11013,
         n11014, n11015, n11016, n11017, n11018, n11019, n11020, n11021,
         n11022, n11023, n11024, n11025, n11026, n11027, n11028, n11029,
         n11030, n11031, n11032, n11033, n11034, n11035, n11036, n11037,
         n11038, n11039, n11040, n11041, n11042, n11043, n11044, n11045,
         n11046, n11047, n11048, n11049, n11050, n11051, n11052, n11053,
         n11054, n11055, n11056, n11057, n11058, n11059, n11060, n11061,
         n11062, n11063, n11064, n11065, n11066, n11067, n11068, n11069,
         n11070, n11071, n11072, n11073, n11074, n11075, n11076, n11077,
         n11078, n11079, n11080, n11081, n11082, n11083, n11084, n11085,
         n11086, n11087, n11088, n11089, n11090, n11091, n11092, n11093,
         n11094, n11095, n11096, n11097, n11098, n11099, n11100, n11101,
         n11102, n11103, n11104, n11105, n11106, n11107, n11108, n11109,
         n11110, n11111, n11112, n11113, n11114, n11115, n11116, n11117,
         n11118, n11119, n11120, n11121, n11122, n11123, n11124, n11125,
         n11126, n11127, n11128, n11129, n11130, n11131, n11132, n11133,
         n11134, n11135, n11136, n11137, n11138, n11139, n11140, n11141,
         n11142, n11143, n11144, n11145, n11146, n11147, n11148, n11149,
         n11150, n11151, n11152, n11153, n11154, n11155, n11156, n11157,
         n11158, n11159, n11160, n11161, n11162, n11163, n11164, n11165,
         n11166, n11167, n11168, n11169, n11170, n11171, n11172, n11173,
         n11174, n11175, n11176, n11177, n11178, n11179, n11180, n11181,
         n11182, n11183, n11184, n11185, n11186, n11187, n11188, n11189,
         n11190, n11191, n11192, n11193, n11194, n11195, n11196, n11197,
         n11198, n11199, n11200, n11201, n11202, n11203, n11204, n11205,
         n11206, n11207, n11208, n11209, n11210, n11211, n11212, n11213,
         n11214, n11215, n11216, n11217, n11218, n11219, n11220, n11221,
         n11222, n11223, n11224, n11225, n11226, n11227, n11228, n11229,
         n11230, n11231, n11232, n11233, n11234, n11235, n11236, n11237,
         n11238, n11239, n11240, n11241, n11242, n11243, n11244, n11245,
         n11246, n11247, n11248, n11249, n11250, n11251, n11252, n11253,
         n11254, n11255, n11256, n11257, n11258, n11259, n11260, n11261,
         n11262, n11263, n11264, n11265, n11266, n11267, n11268, n11269,
         n11270, n11271, n11272, n11273, n11274, n11275, n11276, n11277,
         n11278, n11279, n11280, n11281, n11282, n11283, n11284, n11285,
         n11286, n11287, n11288, n11289, n11290, n11291, n11292, n11293,
         n11294, n11295, n11296, n11297, n11298, n11299, n11300, n11301,
         n11302, n11303, n11304, n11305, n11306, n11307, n11308, n11309,
         n11310, n11311, n11312, n11313, n11314, n11315, n11316, n11317,
         n11318, n11319, n11320, n11321, n11322, n11323, n11324, n11325,
         n11326, n11327, n11328, n11329, n11330, n11331, n11332, n11333,
         n11334, n11335, n11336, n11337, n11338, n11339, n11340, n11341,
         n11342, n11343, n11344, n11345, n11346, n11347, n11348, n11349,
         n11350, n11351, n11352, n11353, n11354, n11355, n11356, n11357,
         n11358, n11359, n11360, n11361, n11362, n11363, n11364, n11365,
         n11366, n11367, n11368, n11369, n11370, n11371, n11372, n11373,
         n11374, n11375, n11376, n11377, n11378, n11379, n11380, n11381,
         n11382, n11383, n11384, n11385, n11386, n11387, n11388, n11389,
         n11390, n11391, n11392, n11393, n11394, n11395, n11396, n11397,
         n11398, n11399, n11400, n11401, n11402, n11403, n11404, n11405,
         n11406, n11407, n11408, n11409, n11410, n11411, n11412, n11413,
         n11414, n11415, n11416, n11417, n11418, n11419, n11420, n11421,
         n11422, n11423, n11424, n11425, n11426, n11427, n11428, n11429,
         n11430, n11431, n11432, n11433, n11434, n11435, n11436, n11437,
         n11438, n11439, n11440, n11441, n11442, n11443, n11444, n11445,
         n11446, n11447, n11448, n11449, n11450, n11451, n11452, n11453,
         n11454, n11455, n11456, n11457, n11458, n11459, n11460, n11461,
         n11462, n11463, n11464, n11465, n11466, n11467, n11468, n11469,
         n11470, n11471, n11472, n11473, n11474, n11475, n11476, n11477,
         n11478, n11479, n11480, n11481, n11482, n11483, n11484, n11485,
         n11486, n11487, n11488, n11489, n11490, n11491, n11492, n11493,
         n11494, n11495, n11496, n11497, n11498, n11499, n11500, n11501,
         n11502, n11503, n11504, n11505, n11506, n11507, n11508, n11509,
         n11510, n11511, n11512, n11513, n11514, n11515, n11516, n11517,
         n11518, n11519, n11520, n11521, n11522, n11523, n11524, n11525,
         n11526, n11527, n11528, n11529, n11530, n11531, n11532, n11533,
         n11534, n11535, n11536, n11537, n11538, n11539, n11540, n11541,
         n11542, n11543, n11544, n11545, n11546, n11547, n11548, n11549,
         n11550, n11551, n11552, n11553, n11554, n11555, n11556, n11557,
         n11558, n11559, n11560, n11561, n11562, n11563, n11564, n11565,
         n11566, n11567, n11568, n11569, n11570, n11571, n11572, n11573,
         n11574, n11575, n11576, n11577, n11578, n11579, n11580, n11581,
         n11582, n11583, n11584, n11585, n11586, n11587, n11588, n11589,
         n11590, n11591, n11592, n11593, n11594, n11595, n11596, n11597,
         n11598, n11599, n11600, n11601, n11602, n11603, n11604, n11605,
         n11606, n11607, n11608, n11609, n11610, n11611, n11612, n11613,
         n11614, n11615, n11616, n11617, n11618, n11619, n11620, n11621,
         n11622, n11623, n11624, n11625, n11626, n11627, n11628, n11629,
         n11630, n11631, n11632, n11633, n11634, n11635, n11636, n11637,
         n11638, n11639, n11640, n11641, n11642, n11643, n11644, n11645,
         n11646, n11647, n11648, n11649, n11650, n11651, n11652, n11653,
         n11654, n11655, n11656, n11657, n11658, n11659, n11660, n11661,
         n11662, n11663, n11664, n11665, n11666, n11667, n11668, n11669,
         n11670, n11671, n11672, n11673, n11674, n11675, n11676, n11677,
         n11678, n11679, n11680, n11681, n11682, n11683, n11684, n11685,
         n11686, n11687, n11688, n11689, n11690, n11691, n11692, n11693,
         n11694, n11695, n11696, n11697, n11698, n11699, n11700, n11701,
         n11702, n11703, n11704, n11705, n11706, n11707, n11708, n11709,
         n11710, n11711, n11712, n11713, n11714, n11715, n11716, n11717,
         n11718, n11719, n11720, n11721, n11722, n11723, n11724, n11725,
         n11726, n11727, n11728, n11729, n11730, n11731, n11732, n11733,
         n11734, n11735, n11736, n11737, n11738, n11739, n11740, n11741,
         n11742, n11743, n11744, n11745, n11746, n11747, n11748, n11749,
         n11750, n11751, n11752, n11753, n11754, n11755, n11756, n11757,
         n11758, n11759, n11760, n11761, n11762, n11763, n11764, n11765,
         n11766, n11767, n11768, n11769, n11770, n11771, n11772, n11773,
         n11774, n11775, n11776, n11777, n11778, n11779, n11780, n11781,
         n11782, n11783, n11784, n11785, n11786, n11787, n11788, n11789,
         n11790, n11791, n11792, n11793, n11794, n11795, n11796, n11797,
         n11798, n11799, n11800, n11801, n11802, n11803, n11804, n11805,
         n11806, n11807, n11808, n11809, n11810, n11811, n11812, n11813,
         n11814, n11815, n11816, n11817, n11818, n11819, n11820, n11821,
         n11822, n11823, n11824, n11825, n11826, n11827, n11828, n11829,
         n11830, n11831, n11832, n11833, n11834, n11835, n11836, n11837,
         n11838, n11839, n11840, n11841, n11842, n11843, n11844, n11845,
         n11846, n11847, n11848, n11849, n11850, n11851, n11852, n11853,
         n11854, n11855, n11856, n11857, n11858, n11859, n11860, n11861,
         n11862, n11863, n11864, n11865, n11866, n11867, n11868, n11869,
         n11870, n11871, n11872, n11873, n11874, n11875, n11876, n11877,
         n11878, n11879, n11880, n11881, n11882, n11883, n11884, n11885,
         n11886, n11887, n11888, n11889, n11890, n11891, n11892, n11893,
         n11894, n11895, n11896, n11897, n11898, n11899, n11900, n11901,
         n11902, n11903, n11904, n11905, n11906, n11907, n11908, n11909,
         n11910, n11911, n11912, n11913, n11914, n11915, n11916, n11917,
         n11918, n11919, n11920, n11921, n11922, n11923, n11924, n11925,
         n11926, n11927, n11928, n11929, n11930, n11931, n11932, n11933,
         n11934, n11935, n11936, n11937, n11938, n11939, n11940, n11941,
         n11942, n11943, n11944, n11945, n11946, n11947, n11948, n11949,
         n11950, n11951, n11952, n11953, n11954, n11955, n11956, n11957,
         n11958, n11959, n11960, n11961, n11962, n11963, n11964, n11965,
         n11966, n11967, n11968, n11969, n11970, n11971, n11972, n11973,
         n11974, n11975, n11976, n11977, n11978, n11979, n11980, n11981,
         n11982, n11983, n11984, n11985, n11986, n11987, n11988, n11989,
         n11990, n11991, n11992, n11993, n11994, n11995, n11996, n11997,
         n11998, n11999, n12000, n12001, n12002, n12003, n12004, n12005,
         n12006, n12007, n12008, n12009, n12010, n12011, n12012, n12013,
         n12014, n12015, n12016, n12017, n12018, n12019, n12020, n12021,
         n12022, n12023, n12024, n12025, n12026, n12027, n12028, n12029,
         n12030, n12031, n12032, n12033, n12034, n12035, n12036, n12037,
         n12038, n12039, n12040, n12041, n12042, n12043, n12044, n12045,
         n12046, n12047, n12048, n12049, n12050, n12051, n12052, n12053,
         n12054, n12055, n12056, n12057, n12058, n12059, n12060, n12061,
         n12062, n12063, n12064, n12065, n12066, n12067, n12068, n12069,
         n12070, n12071, n12072, n12073, n12074, n12075, n12076, n12077,
         n12078, n12079, n12080, n12081, n12082, n12083, n12084, n12085,
         n12086, n12087, n12088, n12089, n12090, n12091, n12092, n12093,
         n12094, n12095, n12096, n12097, n12098, n12099, n12100, n12101,
         n12102, n12103, n12104, n12105, n12106, n12107, n12108, n12109,
         n12110, n12111, n12112, n12113, n12114, n12115, n12116, n12117,
         n12118, n12119, n12120, n12121, n12122, n12123, n12124, n12125,
         n12126, n12127, n12128, n12129, n12130, n12131, n12132, n12133,
         n12134, n12135, n12136, n12137, n12138, n12139, n12140, n12141,
         n12142, n12143, n12144, n12145, n12146, n12147, n12148, n12149,
         n12150, n12151, n12152, n12153, n12154, n12155, n12156, n12157,
         n12158, n12159, n12160, n12161, n12162, n12163, n12164, n12165,
         n12166, n12167, n12168, n12169, n12170, n12171, n12172, n12173,
         n12174, n12175, n12176, n12177, n12178, n12179, n12180, n12181,
         n12182, n12183, n12184, n12185, n12186, n12187, n12188, n12189,
         n12190, n12191, n12192, n12193, n12194, n12195, n12196, n12197,
         n12198, n12199, n12200, n12201, n12202, n12203, n12204, n12205,
         n12206, n12207, n12208, n12209, n12210, n12211, n12212, n12213,
         n12214, n12215, n12216, n12217, n12218, n12219, n12220, n12221,
         n12222, n12223, n12224, n12225, n12226, n12227, n12228, n12229,
         n12230, n12231, n12232, n12233, n12234, n12235, n12236, n12237,
         n12238, n12239, n12240, n12241, n12242, n12243, n12244, n12245,
         n12246, n12247, n12248, n12249, n12250, n12251, n12252, n12253,
         n12255, n12256, n12257, n12258, n12259, n12260, n12261, n12262,
         n12263, n12264, n12265, n12266, n12267, n12268, n12269, n12270,
         n12271, n12272, n12273, n12274, n12275, n12276, n12277, n12278,
         n12279, n12280, n12281, n12282, n12283, n12284, n12285, n12286,
         n12287, n12288, n12289, n12290, n12291, n12292, n12293, n12294,
         n12295, n12296, n12297, n12298, n12299, n12300, n12301, n12302,
         n12303, n12304, n12305, n12306, n12307, n12308, n12309, n12310,
         n12311, n12312, n12313, n12314, n12315, n12316, n12317, n12318,
         n12319, n12320, n12321, n12322, n12323, n12324, n12325, n12326,
         n12327, n12328, n12329, n12330, n12331, n12332, n12333, n12334,
         n12335, n12336, n12337, n12338, n12339, n12340, n12341, n12342,
         n12343, n12344, n12345, n12346, n12347, n12348, n12349, n12350,
         n12351, n12352, n12353, n12354, n12355, n12356, n12357, n12358,
         n12359, n12360, n12361, n12362, n12363, n12364, n12365, n12366,
         n12367, n12368, n12369, n12370, n12371, n12372, n12373, n12374,
         n12375, n12376, n12377, n12378, n12379, n12380, n12381, n12382,
         n12383, n12384, n12385, n12386, n12387, n12388, n12389, n12390,
         n12391, n12392, n12393, n12394, n12395, n12396, n12397, n12398,
         n12399, n12400, n12401, n12402, n12403, n12404, n12405, n12406,
         n12407, n12408, n12409, n12410, n12411, n12412, n12413, n12414,
         n12415, n12416, n12417, n12418, n12419, n12420, n12421, n12422,
         n12423, n12424, n12425, n12426, n12427, n12428, n12429, n12430,
         n12431, n12432, n12433, n12434, n12435, n12436, n12437, n12438,
         n12439, n12440, n12441, n12442, n12443, n12444, n12445, n12446,
         n12447, n12448, n12449, n12450, n12451, n12452, n12453, n12454,
         n12455, n12456, n12457, n12458, n12459, n12460, n12461, n12462,
         n12463, n12464, n12465, n12466, n12467, n12468, n12469, n12470,
         n12471, n12472, n12473, n12474, n12475, n12476, n12477, n12478,
         n12479, n12480, n12481, n12482, n12483, n12484, n12485, n12486,
         n12487, n12488, n12489, n12490, n12491, n12492, n12493, n12494,
         n12495, n12496, n12497, n12498, n12499, n12500, n12501, n12502,
         n12503, n12504, n12505, n12506, n12507, n12508, n12509, n12510,
         n12511, n12512, n12513, n12514, n12515, n12516, n12517, n12518,
         n12519, n12520, n12521, n12522, n12523, n12524, n12525, n12526,
         n12527, n12528, n12529, n12530, n12531, n12532, n12533, n12534,
         n12535, n12536, n12537, n12538, n12539, n12540, n12541, n12542,
         n12543, n12544, n12545, n12546, n12547, n12548, n12549, n12550,
         n12551, n12552, n12553, n12554, n12555, n12556, n12557, n12558,
         n12559, n12560, n12561, n12562, n12563, n12564, n12565, n12566,
         n12567, n12568, n12569, n12570, n12571, n12572, n12573, n12574,
         n12575, n12576, n12577, n12578, n12579, n12580, n12581, n12582,
         n12583, n12584, n12585, n12586, n12587, n12588, n12589, n12590,
         n12591, n12592, n12593, n12594, n12595, n12596, n12597, n12598,
         n12599, n12600, n12601, n12602, n12603, n12604, n12605, n12606,
         n12607, n12608, n12609, n12610, n12611, n12612, n12613, n12614,
         n12615, n12616, n12617, n12618, n12619, n12620, n12621, n12622,
         n12623, n12624, n12625, n12626, n12627, n12628, n12629, n12630,
         n12631, n12632, n12633, n12634, n12635, n12636, n12637, n12638,
         n12639, n12640, n12641, n12642, n12643, n12644, n12645, n12646,
         n12647, n12648, n12649, n12650, n12651, n12652, n12653, n12654,
         n12655, n12656, n12657, n12658, n12659, n12660, n12661, n12662,
         n12663, n12664, n12665, n12666, n12667, n12668, n12669, n12670,
         n12671, n12672, n12673, n12674, n12675, n12676, n12677, n12678,
         n12679, n12680, n12681, n12682, n12683, n12684, n12685, n12686,
         n12687, n12688, n12689, n12690, n12691, n12692, n12693, n12694,
         n12695, n12696, n12697, n12698, n12699, n12700, n12701, n12702,
         n12703, n12704, n12705, n12706, n12707, n12708, n12709, n12710,
         n12711, n12712, n12713, n12714, n12715, n12716, n12717, n12718,
         n12719, n12720, n12721, n12722, n12723, n12724, n12725, n12726,
         n12727, n12728, n12729, n12730, n12731, n12732, n12733, n12734,
         n12735, n12736, n12737, n12738, n12739, n12740, n12741, n12742,
         n12743, n12744, n12745, n12746, n12747, n12748, n12749, n12750,
         n12751, n12752, n12753, n12754, n12755, n12756, n12757, n12758,
         n12759, n12760, n12761, n12762, n12763, n12764, n12765, n12766,
         n12767, n12768, n12769, n12770, n12771, n12772, n12773, n12774,
         n12775, n12776, n12777, n12778, n12779, n12780, n12781, n12782,
         n12783, n12784, n12785, n12786, n12787, n12788, n12789, n12790,
         n12791, n12792, n12793, n12794, n12795, n12796, n12797, n12798,
         n12799, n12800, n12801, n12802, n12803, n12804, n12805, n12806,
         n12807, n12808, n12809, n12810, n12811, n12812, n12813, n12814,
         n12815, n12816, n12817, n12818, n12819, n12820, n12821, n12822,
         n12823, n12824, n12825, n12826, n12827, n12828, n12829, n12830,
         n12831, n12832, n12833, n12834, n12835, n12836, n12837, n12838,
         n12839, n12840, n12841, n12842, n12843, n12844, n12845, n12846,
         n12847, n12848, n12849, n12850, n12851, n12852, n12853, n12854,
         n12855, n12856, n12857, n12858, n12859, n12860, n12861, n12862,
         n12863, n12864, n12865, n12866, n12867, n12868, n12869, n12870,
         n12871, n12872, n12873, n12874, n12875, n12876, n12877, n12878,
         n12879, n12880, n12881, n12882, n12883, n12884, n12885, n12886,
         n12887, n12888, n12889, n12890, n12891, n12892, n12893, n12894,
         n12895, n12896, n12897, n12898, n12899, n12900, n12901, n12902,
         n12903, n12904, n12905, n12906, n12907, n12908, n12909, n12910,
         n12911, n12912, n12913, n12914, n12915, n12916, n12917, n12918,
         n12919, n12920, n12921, n12922, n12923, n12924, n12925, n12926,
         n12927, n12928, n12929, n12930, n12931, n12932, n12933, n12934,
         n12935, n12936, n12937, n12938, n12939, n12940, n12941, n12942,
         n12943, n12944, n12945, n12946, n12947, n12948, n12949, n12950,
         n12951, n12952, n12953, n12954, n12955, n12956, n12957, n12958,
         n12959, n12960, n12961, n12962, n12963, n12964, n12965, n12966,
         n12967, n12968, n12969, n12970, n12971, n12972, n12973, n12974,
         n12975, n12976, n12977, n12978, n12979, n12980, n12981, n12982,
         n12983, n12984, n12985, n12986, n12987, n12988, n12989, n12990,
         n12991, n12992, n12993, n12994, n12995, n12996, n12997, n12998,
         n12999, n13000, n13001, n13002, n13003, n13004, n13005, n13006,
         n13007, n13008, n13009, n13010, n13011, n13012, n13013, n13014,
         n13015, n13016, n13017, n13018, n13019, n13020, n13021, n13022,
         n13023, n13024, n13025, n13026, n13027, n13028, n13029, n13030,
         n13031, n13032, n13033, n13034, n13035, n13036, n13037, n13038,
         n13039, n13040, n13041, n13042, n13043, n13044, n13045, n13046,
         n13047, n13048, n13049, n13050, n13051, n13052, n13053, n13054,
         n13055, n13056, n13057, n13058, n13059, n13060, n13061, n13062,
         n13063, n13064, n13065, n13066, n13067, n13068, n13069, n13070,
         n13071, n13072, n13073, n13074, n13075, n13076, n13077, n13078,
         n13079, n13080, n13081, n13082, n13083, n13084, n13085, n13086,
         n13087, n13088, n13089, n13090, n13091, n13092, n13093, n13094,
         n13095, n13096, n13097, n13098, n13099, n13100, n13101, n13102,
         n13103, n13104, n13105, n13106, n13107, n13108, n13109, n13110,
         n13111, n13112, n13113, n13114, n13115, n13116, n13117, n13118,
         n13119, n13120, n13121, n13122, n13123, n13124, n13125, n13126,
         n13127, n13128, n13129, n13130, n13131, n13132, n13133, n13134,
         n13135, n13136, n13137, n13138, n13139, n13140, n13141, n13142,
         n13143, n13144, n13145, n13146, n13147, n13148, n13149, n13150,
         n13151, n13152, n13153, n13154, n13155, n13156, n13157, n13158,
         n13159, n13160, n13161, n13162, n13163, n13164, n13165, n13166,
         n13167, n13168, n13169, n13170, n13171, n13172, n13173, n13174,
         n13175, n13176, n13177, n13178, n13179, n13180, n13181, n13182,
         n13183, n13184, n13185, n13186, n13187, n13188, n13189, n13190,
         n13191, n13192, n13193, n13194, n13195, n13196, n13197, n13198,
         n13199, n13200, n13201, n13202, n13203, n13204, n13205, n13206,
         n13207, n13208, n13209, n13210, n13211, n13212, n13213, n13214,
         n13215, n13216, n13217, n13218, n13219, n13220, n13221, n13222,
         n13223, n13224, n13225, n13226, n13227, n13228, n13229, n13230,
         n13231, n13232, n13233, n13234, n13235, n13236, n13237, n13238,
         n13239, n13240, n13241, n13242, n13243, n13244, n13245, n13246,
         n13247, n13248, n13249, n13250, n13251, n13252, n13253, n13254,
         n13255, n13256, n13257, n13258, n13259, n13260, n13261, n13262,
         n13263, n13264, n13265, n13266, n13267, n13268, n13269, n13270,
         n13271, n13272, n13273, n13274, n13275, n13276, n13277, n13278,
         n13279, n13280, n13281, n13282, n13283, n13284, n13285, n13286,
         n13287, n13288, n13289, n13290, n13291, n13292, n13293, n13294,
         n13295, n13296, n13297, n13298, n13299, n13300, n13301, n13302,
         n13303, n13304, n13305, n13306, n13307, n13308, n13309, n13310,
         n13311, n13312, n13313, n13314, n13315, n13316, n13317, n13318,
         n13319, n13320, n13321, n13322, n13323, n13324, n13325, n13326,
         n13327, n13328, n13329, n13330, n13331, n13332, n13333, n13334,
         n13335, n13336, n13337, n13338, n13339, n13340, n13341, n13342,
         n13343, n13344, n13345, n13346, n13347, n13348, n13349, n13350,
         n13351, n13352, n13353, n13354, n13355, n13356, n13357, n13358,
         n13359, n13360, n13361, n13362, n13363, n13364, n13365, n13366,
         n13367, n13368, n13369, n13370, n13371, n13372, n13373, n13374,
         n13375, n13376, n13377, n13378, n13379, n13380, n13381, n13382,
         n13383, n13384, n13385, n13386, n13387, n13388, n13389, n13390,
         n13391, n13392, n13393, n13394, n13395, n13396, n13397, n13398,
         n13399, n13400, n13401, n13402, n13403, n13404, n13405, n13406,
         n13407, n13408, n13409, n13410, n13411, n13412, n13413, n13414,
         n13415, n13416, n13417, n13418, n13419, n13420, n13421, n13422,
         n13423, n13424, n13425, n13426, n13427, n13428, n13429, n13430,
         n13431, n13432, n13433, n13434, n13435, n13436, n13437, n13438,
         n13439, n13440, n13441, n13442, n13443, n13444, n13445, n13446,
         n13447, n13448, n13449, n13450, n13451, n13452, n13453, n13454,
         n13455, n13456, n13457, n13458, n13459, n13460, n13461, n13462,
         n13463, n13464, n13465, n13466, n13467, n13468, n13469, n13470,
         n13471, n13472, n13473, n13474, n13475, n13476, n13477, n13478,
         n13479, n13480, n13481, n13482, n13483, n13484, n13485, n13486,
         n13487, n13488, n13489, n13490, n13491, n13492, n13493, n13494,
         n13495, n13496, n13497, n13498, n13499, n13500, n13501, n13502,
         n13503, n13504, n13505, n13506, n13507, n13508, n13509, n13510,
         n13511, n13512, n13513, n13514, n13515, n13516, n13517, n13518,
         n13519, n13520, n13521, n13522, n13523, n13524, n13525, n13526,
         n13527, n13528, n13529, n13530, n13531, n13532, n13533, n13534,
         n13535, n13536, n13537, n13538, n13539, n13540, n13541, n13542,
         n13543, n13544, n13545, n13546, n13547, n13548, n13549, n13550,
         n13551, n13552, n13553, n13554, n13555, n13556, n13557, n13558,
         n13559, n13560, n13561, n13562, n13563, n13564, n13565, n13566,
         n13567, n13568, n13569, n13570, n13571, n13572, n13573, n13574,
         n13575, n13576, n13577, n13578, n13579, n13580, n13581, n13582,
         n13583, n13584, n13585, n13586, n13587, n13588, n13589, n13590,
         n13591, n13592, n13593, n13594, n13595, n13596, n13597, n13598,
         n13599, n13600, n13601, n13602, n13603, n13604, n13605, n13606,
         n13607, n13608, n13609, n13610, n13611, n13612, n13613, n13614,
         n13615, n13616, n13617, n13618, n13619, n13620, n13621, n13622,
         n13623, n13624, n13625, n13626, n13627, n13628, n13629, n13630,
         n13631, n13632, n13633, n13634, n13635, n13636, n13637, n13638,
         n13639, n13640, n13641, n13642, n13643, n13644, n13645, n13646,
         n13647, n13648, n13649, n13650, n13651, n13652, n13653, n13654,
         n13655, n13656, n13657, n13658, n13659, n13660, n13661, n13662,
         n13663, n13664, n13665, n13666, n13667, n13668, n13669, n13670,
         n13671, n13672, n13673, n13674, n13675, n13676, n13677, n13678,
         n13679, n13680, n13681, n13682, n13683, n13684, n13685, n13686,
         n13687, n13688, n13689, n13690, n13691, n13692, n13693, n13694,
         n13695, n13696, n13697, n13698, n13699, n13700, n13701, n13702,
         n13703, n13704, n13705, n13706, n13707, n13708, n13709, n13710,
         n13711, n13712, n13713, n13714, n13715, n13716, n13717, n13718,
         n13719, n13720, n13721, n13722, n13723, n13724, n13725, n13726,
         n13727, n13728, n13729, n13730, n13731, n13732, n13733, n13734,
         n13735, n13736, n13737, n13738, n13739, n13740, n13741, n13742,
         n13743, n13744, n13745, n13746, n13747, n13748, n13749, n13750,
         n13751, n13752, n13753, n13754, n13755, n13756, n13757, n13758,
         n13759, n13760, n13761, n13762, n13763, n13764, n13765, n13766,
         n13767, n13768, n13769, n13770, n13771, n13772, n13773, n13774,
         n13775, n13776, n13777, n13778, n13779, n13780, n13781, n13782,
         n13783, n13784, n13785, n13786, n13787, n13788, n13789, n13790,
         n13791, n13792, n13793, n13794, n13795, n13796, n13797, n13798,
         n13799, n13800, n13801, n13802, n13803, n13804, n13805, n13806,
         n13807, n13808, n13809, n13810, n13811, n13812, n13813, n13814,
         n13815, n13816, n13817, n13818, n13819, n13820, n13821, n13822,
         n13823, n13824, n13825, n13826, n13827, n13828, n13829, n13830,
         n13831, n13832, n13833, n13834, n13835, n13836, n13837, n13838,
         n13839, n13840, n13841, n13842, n13843, n13844, n13845, n13846,
         n13847, n13848, n13849, n13850, n13851, n13852, n13853, n13854,
         n13855, n13856, n13857, n13858, n13859, n13860, n13861, n13862,
         n13863, n13864, n13865, n13866, n13867, n13868, n13869, n13870,
         n13871, n13872, n13873, n13874, n13875, n13876, n13877, n13878,
         n13879, n13880, n13881, n13882, n13883, n13884, n13885, n13886,
         n13887, n13888, n13889, n13890, n13891, n13892, n13893, n13894,
         n13895, n13896, n13897, n13898, n13899, n13900, n13901, n13902,
         n13903, n13904, n13905, n13906, n13907, n13908, n13909, n13910,
         n13911, n13912, n13913, n13914, n13915, n13916, n13917, n13918,
         n13919, n13920, n13921, n13922, n13923, n13924, n13925, n13926,
         n13927, n13928, n13929, n13930, n13931, n13932, n13933, n13934,
         n13935, n13936, n13937, n13938, n13939, n13940, n13941, n13942,
         n13943, n13944, n13945, n13946, n13947, n13948, n13949, n13950,
         n13951, n13952, n13953, n13954, n13955, n13956, n13957, n13958,
         n13959, n13960, n13961, n13962, n13963, n13964, n13965, n13966,
         n13967, n13968, n13969, n13970, n13971, n13972, n13973, n13974,
         n13975, n13976, n13977, n13978, n13979, n13980, n13981, n13982,
         n13983, n13984, n13985, n13986, n13987, n13988, n13989, n13990,
         n13991, n13992, n13993, n13994, n13995, n13996, n13997, n13998,
         n13999, n14000, n14001, n14002, n14003, n14004, n14005, n14006,
         n14007, n14008, n14009, n14010, n14011, n14012, n14013, n14014,
         n14015, n14016, n14017, n14018, n14019, n14020, n14021, n14022,
         n14023, n14024, n14025, n14026, n14027, n14028, n14029, n14030,
         n14031, n14032, n14033, n14034, n14035, n14036, n14037, n14038,
         n14039, n14040, n14041, n14042, n14043, n14044, n14045, n14046,
         n14047, n14048, n14049, n14050, n14051, n14052, n14053, n14054,
         n14055, n14056, n14057, n14058, n14059, n14060, n14061, n14062,
         n14063, n14064, n14065, n14066, n14067, n14068, n14069, n14070,
         n14071, n14072, n14073, n14074, n14075, n14076, n14077, n14078,
         n14079, n14080, n14081, n14082, n14083, n14084, n14085, n14086,
         n14087, n14088, n14089, n14090, n14091, n14092, n14093, n14094,
         n14095, n14096, n14097, n14098, n14099, n14100, n14101, n14102,
         n14103, n14104, n14105, n14106, n14107, n14108, n14109, n14110,
         n14111, n14112, n14113, n14114, n14115, n14116, n14117, n14118,
         n14119, n14120, n14121, n14122, n14123, n14124, n14125, n14126,
         n14127, n14128, n14129, n14130, n14131, n14132, n14133, n14134,
         n14135, n14136, n14137, n14138, n14139, n14140, n14141, n14142,
         n14143, n14144, n14145, n14146, n14147, n14148, n14149, n14150,
         n14151, n14152, n14153, n14154, n14155, n14156, n14157, n14158,
         n14159, n14160, n14161, n14162, n14163, n14164, n14165, n14166,
         n14167, n14168, n14169, n14170, n14171, n14172, n14173, n14174,
         n14175, n14176, n14177, n14178, n14179, n14180, n14181, n14182,
         n14183, n14184, n14185, n14186, n14187, n14188, n14189, n14190,
         n14191, n14192, n14193, n14194, n14195, n14196, n14197, n14198,
         n14199, n14200, n14201, n14202, n14203, n14204, n14205, n14206,
         n14207, n14208, n14209, n14210, n14211, n14212, n14213, n14214,
         n14215, n14216, n14217, n14218, n14219, n14220, n14221, n14222,
         n14223, n14224, n14225, n14226, n14227, n14228, n14229, n14230,
         n14231, n14232, n14233, n14234, n14235, n14236, n14237, n14238,
         n14239, n14240, n14241, n14242, n14243, n14244, n14245, n14246,
         n14247, n14248, n14249, n14250, n14251, n14252, n14253, n14254,
         n14255, n14256, n14257, n14258, n14259, n14260, n14261, n14262,
         n14263, n14264, n14265, n14266, n14267, n14268, n14269, n14270,
         n14271, n14272, n14273, n14274, n14275, n14276, n14277, n14278,
         n14279, n14280, n14281, n14282, n14283, n14284, n14285, n14286,
         n14287, n14288, n14289, n14290, n14291, n14292, n14293, n14294,
         n14295, n14296, n14297, n14298, n14299, n14300, n14301, n14302,
         n14303, n14304, n14305, n14306, n14307, n14308, n14309, n14310,
         n14311, n14312, n14313, n14314, n14315, n14316, n14317, n14318,
         n14319, n14320, n14321, n14322, n14323, n14324, n14325, n14326,
         n14327, n14328, n14329, n14330, n14331, n14332, n14333, n14334,
         n14335, n14336, n14337, n14338, n14339, n14340, n14341, n14342,
         n14343, n14344, n14345, n14346, n14347, n14348, n14349, n14350,
         n14351, n14352, n14353, n14354, n14355, n14356, n14357, n14358,
         n14359, n14360, n14361, n14362, n14363, n14364, n14365, n14366,
         n14367, n14368, n14369, n14370, n14371, n14372, n14373, n14374,
         n14375, n14376, n14377, n14378, n14379, n14380, n14381, n14382,
         n14383, n14384, n14385, n14386, n14387, n14388, n14389, n14390,
         n14391, n14392, n14393, n14394, n14395, n14396, n14397, n14398,
         n14399, n14400, n14401, n14402, n14403, n14404, n14405, n14406,
         n14407, n14408, n14409, n14410, n14411, n14412, n14413, n14414,
         n14415, n14416, n14417, n14418, n14419, n14420, n14421, n14422,
         n14423, n14424, n14425, n14426, n14427, n14428, n14429, n14430,
         n14431, n14432, n14433, n14434, n14435, n14436, n14437, n14438,
         n14439, n14440, n14441, n14442, n14443, n14444, n14445, n14446,
         n14447, n14448, n14449, n14450, n14451, n14452, n14453, n14454,
         n14455, n14456, n14457, n14458, n14459, n14460, n14461, n14462,
         n14463, n14464, n14465, n14466, n14467, n14468, n14469, n14470,
         n14471, n14472, n14473, n14474, n14475, n14476, n14477, n14478,
         n14479, n14480, n14481, n14482, n14483, n14484, n14485, n14486,
         n14487, n14488, n14489, n14490, n14491, n14492, n14493, n14494,
         n14495, n14496, n14497, n14498, n14499, n14500, n14501, n14502,
         n14503, n14504, n14505, n14506, n14507, n14508, n14509, n14510,
         n14511, n14512, n14513, n14514, n14515, n14516, n14517, n14518,
         n14519, n14520, n14521, n14522, n14523, n14524, n14525, n14526,
         n14527, n14528, n14529, n14530, n14531, n14532, n14533, n14534,
         n14535, n14536, n14537, n14538, n14539, n14540, n14541, n14542,
         n14543, n14544, n14545, n14546, n14547, n14548, n14549, n14550,
         n14551, n14552, n14553, n14554, n14555, n14556, n14557, n14558,
         n14559, n14560, n14561, n14562, n14563, n14564, n14565, n14566,
         n14567, n14568, n14569, n14570, n14571, n14572, n14573, n14574,
         n14575, n14576, n14577, n14578, n14579, n14580, n14581, n14582,
         n14583, n14584, n14585, n14586, n14587, n14588, n14589, n14590,
         n14591, n14592, n14593, n14594, n14595, n14596, n14597, n14598,
         n14599, n14600, n14601, n14602, n14603, n14604, n14606, n14607,
         n14608, n14609, n14610, n14611, n14612, n14613, n14614, n14615,
         n14616, n14617, n14618, n14619, n14620, n14621, n14622, n14623,
         n14624, n14625, n14626, n14627, n14628, n14629, n14630, n14631,
         n14632, n14633, n14634, n14635, n14636, n14637, n14638, n14639,
         n14640, n14641, n14642, n14643, n14644, n14645, n14646, n14647,
         n14648, n14649, n14650, n14651, n14652, n14653, n14654, n14655,
         n14656, n14657, n14658, n14659, n14660, n14661, n14662, n14663,
         n14664, n14665, n14666, n14667, n14668, n14669, n14670, n14671,
         n14672, n14673, n14674, n14675, n14676, n14677, n14678, n14679,
         n14680, n14681, n14682, n14683, n14684, n14685, n14686, n14687,
         n14688, n14689, n14690, n14691, n14692, n14693, n14694, n14695,
         n14696, n14697, n14698, n14699, n14700, n14701, n14702, n14703,
         n14704, n14705, n14706, n14707, n14708, n14709, n14710, n14711,
         n14712, n14713, n14714, n14715, n14716, n14717, n14718, n14719,
         n14720, n14721, n14722, n14723, n14724, n14725, n14726, n14727,
         n14728, n14729, n14730, n14731, n14732, n14733, n14734, n14735,
         n14736, n14737, n14738, n14739, n14740, n14741, n14742, n14743,
         n14744, n14745, n14746, n14747, n14748, n14749, n14750, n14751,
         n14752, n14753, n14754, n14755, n14756, n14757, n14758, n14759,
         n14760, n14761, n14762, n14763, n14764, n14765, n14766, n14767,
         n14768, n14769, n14770, n14771, n14772, n14773, n14774, n14775,
         n14776, n14777, n14778, n14779, n14780, n14781, n14782, n14783,
         n14784, n14785, n14786, n14787, n14788, n14789, n14790, n14791,
         n14792, n14793, n14794, n14795, n14796, n14797, n14798, n14799,
         n14800, n14801, n14802, n14803, n14804, n14805, n14806, n14807,
         n14808, n14809, n14810, n14811, n14812, n14813, n14814, n14815,
         n14816, n14817, n14818, n14819, n14820, n14821, n14822, n14823,
         n14824, n14825, n14826, n14827, n14828, n14829, n14830, n14831,
         n14832, n14833, n14834, n14835, n14836, n14837, n14838, n14839,
         n14840, n14841, n14842, n14843, n14844, n14845, n14846, n14847,
         n14848, n14849, n14850, n14851, n14852, n14853, n14854, n14855,
         n14856, n14857, n14858, n14859, n14860, n14861, n14862, n14863,
         n14864, n14865, n14866, n14867, n14868, n14869, n14870, n14871,
         n14872, n14873, n14874, n14875, n14876, n14877, n14878, n14879,
         n14880, n14881, n14882, n14883, n14884, n14885, n14886, n14887,
         n14888, n14889, n14890, n14891, n14892, n14893, n14894, n14895,
         n14896, n14897, n14898, n14899, n14900, n14901, n14902, n14903,
         n14904, n14905, n14906, n14907, n14908, n14909, n14910, n14911,
         n14912, n14913, n14914, n14915, n14916, n14917, n14918, n14919,
         n14920, n14921, n14922, n14923, n14924, n14925, n14926, n14927,
         n14928, n14929, n14930, n14931, n14932, n14933, n14934, n14935,
         n14936, n14937, n14938, n14939, n14940, n14941, n14942, n14943,
         n14944, n14945, n14946, n14947, n14948, n14949, n14950, n14951,
         n14952, n14953, n14954, n14955, n14956, n14957, n14958, n14959,
         n14960, n14961, n14962, n14963, n14964, n14965, n14966, n14967,
         n14968, n14969, n14970, n14971, n14972, n14973, n14974, n14975,
         n14976, n14977, n14978, n14979, n14980, n14981, n14982, n14983,
         n14984, n14985, n14986, n14987, n14988, n14989, n14990, n14991,
         n14992, n14993, n14994, n14995, n14996, n14997, n14998, n14999,
         n15000, n15001, n15002, n15003, n15004, n15005, n15006, n15007,
         n15008, n15009, n15010, n15011, n15012, n15013, n15014, n15015,
         n15016, n15017, n15018, n15019, n15020, n15021, n15022, n15023,
         n15024, n15025, n15026, n15027, n15028, n15029, n15030, n15031,
         n15032, n15033, n15034, n15035, n15036, n15037, n15038, n15039,
         n15040, n15041, n15042, n15043, n15044, n15045, n15046, n15047,
         n15048, n15049, n15050, n15051, n15052, n15053, n15054, n15055,
         n15056, n15057, n15058, n15059, n15060, n15061, n15062, n15063,
         n15064, n15065, n15066, n15067, n15068, n15069, n15070, n15071,
         n15072, n15073, n15074, n15075, n15076, n15077, n15078, n15079,
         n15080, n15081, n15082, n15083, n15084, n15085, n15086, n15087,
         n15088, n15089, n15090, n15091, n15092, n15093, n15094, n15095,
         n15096, n15097, n15098, n15099, n15100, n15101, n15102, n15103,
         n15104, n15105, n15106, n15107, n15108, n15109, n15110, n15111,
         n15112, n15113, n15114, n15115, n15116, n15117, n15118, n15119,
         n15120, n15121, n15122, n15123, n15124, n15125, n15126, n15127,
         n15128, n15129, n15130, n15131, n15132, n15133, n15134, n15135,
         n15136, n15137, n15138, n15139, n15140, n15141, n15142, n15143,
         n15144, n15145, n15146, n15147, n15148, n15149, n15150, n15151,
         n15152, n15153, n15154, n15155, n15156, n15157, n15158, n15159,
         n15160, n15161, n15162, n15163, n15164, n15165, n15166, n15167,
         n15168, n15169, n15170, n15171, n15172, n15173, n15174, n15175,
         n15176, n15177, n15178, n15179, n15180, n15181, n15182, n15183,
         n15184, n15185, n15186, n15187, n15188, n15189, n15190, n15191,
         n15192, n15193, n15194, n15195, n15196, n15197, n15198, n15199,
         n15200, n15201, n15202, n15203, n15204, n15205, n15206, n15207,
         n15208, n15209, n15210, n15211, n15212, n15213, n15214, n15215,
         n15216, n15217, n15218, n15219, n15220, n15221, n15222, n15223,
         n15224, n15225, n15226, n15227, n15228, n15229, n15230, n15231,
         n15232, n15233, n15234, n15235, n15236, n15237, n15238, n15239,
         n15240, n15241, n15242, n15243, n15244, n15245, n15246, n15247,
         n15248, n15249, n15250, n15251, n15252, n15253, n15254, n15255,
         n15256, n15257, n15258, n15259, n15260, n15261, n15262, n15263,
         n15264, n15265, n15266, n15267, n15268, n15269, n15270, n15271,
         n15272, n15273, n15274, n15275, n15276, n15277, n15278, n15279,
         n15280, n15281, n15282, n15283, n15284, n15285, n15286, n15287,
         n15288, n15289, n15290, n15291, n15292, n15293, n15294, n15295,
         n15296, n15297, n15298, n15299, n15300, n15301, n15302, n15303,
         n15304, n15305, n15306, n15307, n15308, n15309, n15310, n15311,
         n15312, n15313, n15314, n15315, n15316, n15317, n15318, n15319,
         n15320, n15321, n15322, n15323, n15324, n15325, n15326, n15327,
         n15328, n15329, n15330, n15331, n15332, n15333, n15334, n15335,
         n15336, n15337, n15338, n15339, n15340, n15341, n15342, n15343,
         n15344, n15345, n15346, n15347, n15348, n15349, n15350, n15351,
         n15352, n15353, n15354, n15355, n15356, n15357, n15358, n15359,
         n15360, n15361, n15362, n15363, n15364, n15365, n15366, n15367,
         n15368, n15369, n15370, n15371, n15372, n15373, n15374, n15375,
         n15376, n15377, n15378, n15379, n15380, n15381, n15382, n15383,
         n15384, n15385, n15386, n15387, n15388, n15389, n15390, n15391,
         n15392, n15393, n15394, n15395, n15396, n15397, n15398, n15399,
         n15400, n15401, n15402, n15403, n15404, n15405, n15406, n15407,
         n15408, n15409, n15410, n15411, n15412, n15413, n15414, n15415,
         n15416, n15417, n15418, n15419, n15420, n15421, n15422, n15423,
         n15424, n15425, n15426, n15427, n15428, n15429, n15430, n15431,
         n15432, n15433, n15434, n15435, n15436, n15437, n15438, n15439,
         n15440, n15441, n15442, n15443, n15444, n15445, n15446, n15447,
         n15448, n15449, n15450, n15451, n15452, n15453, n15454, n15455,
         n15456, n15457, n15458, n15459, n15460, n15461, n15462, n15463,
         n15464, n15465, n15467, n15468, n15469, n15470, n15471, n15472,
         n15473, n15474, n15475, n15476, n15477, n15478, n15479, n15480,
         n15481, n15482, n15483, n15484, n15485, n15486, n15487, n15488,
         n15489, n15490, n15491, n15492, n15493, n15494, n15495, n15496,
         n15497, n15498, n15499, n15500, n15501, n15502, n15503, n15504,
         n15505, n15506, n15507, n15508, n15509, n15510, n15511, n15512,
         n15513, n15514, n15515, n15516, n15517, n15518;

  AND2_X1 U7365 ( .A1(n6954), .A2(n6952), .ZN(n14166) );
  INV_X2 U7366 ( .A(n15464), .ZN(n13024) );
  INV_X2 U7367 ( .A(n11299), .ZN(n6622) );
  INV_X1 U7369 ( .A(n6617), .ZN(n8243) );
  INV_X2 U7370 ( .A(n7794), .ZN(n13954) );
  CLKBUF_X2 U7371 ( .A(n8813), .Z(n9168) );
  CLKBUF_X2 U7372 ( .A(n8415), .Z(n6626) );
  INV_X2 U7373 ( .A(n14127), .ZN(n7767) );
  AND2_X2 U7374 ( .A1(n8370), .A2(n8369), .ZN(n8424) );
  NOR2_X1 U7376 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n7691) );
  INV_X2 U7377 ( .A(n12647), .ZN(n12653) );
  NAND2_X1 U7378 ( .A1(n8802), .A2(n7520), .ZN(n8801) );
  AOI22_X1 U7379 ( .A1(n8060), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(n8059), .B2(
        n10449), .ZN(n7759) );
  CLKBUF_X2 U7380 ( .A(n9257), .Z(n11245) );
  AND2_X1 U7382 ( .A1(n7191), .A2(n7190), .ZN(n12659) );
  CLKBUF_X2 U7383 ( .A(n8412), .Z(n6627) );
  NAND2_X1 U7384 ( .A1(n8801), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8800) );
  INV_X1 U7385 ( .A(n7705), .ZN(n7707) );
  OAI22_X1 U7386 ( .A1(n7644), .A2(n7594), .B1(P1_ADDR_REG_6__SCAN_IN), .B2(
        n7593), .ZN(n7595) );
  INV_X1 U7387 ( .A(n11470), .ZN(n12722) );
  INV_X1 U7388 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n12321) );
  NAND2_X1 U7389 ( .A1(n8365), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8364) );
  OR2_X1 U7390 ( .A1(n7054), .A2(n14973), .ZN(n7053) );
  INV_X1 U7391 ( .A(n12458), .ZN(n13122) );
  BUF_X1 U7392 ( .A(n8262), .Z(n13959) );
  INV_X1 U7393 ( .A(n10653), .ZN(n13588) );
  XNOR2_X2 U7394 ( .A(n7655), .B(n7654), .ZN(n14794) );
  OAI21_X2 U7395 ( .B1(P1_REG1_REG_11__SCAN_IN), .B2(n11276), .A(n11271), .ZN(
        n11272) );
  NOR2_X2 U7396 ( .A1(n10610), .A2(P1_ADDR_REG_0__SCAN_IN), .ZN(n7632) );
  NAND2_X2 U7397 ( .A1(n13975), .A2(n7761), .ZN(n14168) );
  AND2_X2 U7398 ( .A1(n8325), .A2(n8324), .ZN(n8326) );
  OAI21_X2 U7399 ( .B1(n6648), .B2(n14381), .A(n14380), .ZN(n14628) );
  INV_X1 U7400 ( .A(n7706), .ZN(n14762) );
  NOR2_X2 U7401 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n8382) );
  XNOR2_X2 U7402 ( .A(n9672), .B(n9656), .ZN(n13160) );
  OAI21_X2 U7403 ( .B1(n9672), .B2(n9671), .A(n9670), .ZN(n12314) );
  AOI21_X2 U7404 ( .B1(n9653), .B2(n9654), .A(n7159), .ZN(n9672) );
  NAND2_X2 U7405 ( .A1(n7703), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7704) );
  BUF_X4 U7406 ( .A(n7740), .Z(n6617) );
  NAND2_X1 U7407 ( .A1(n7705), .A2(n14762), .ZN(n7740) );
  XNOR2_X2 U7408 ( .A(n12052), .B(n12054), .ZN(n12056) );
  XNOR2_X2 U7409 ( .A(n9209), .B(n9208), .ZN(n13162) );
  OAI22_X1 U7410 ( .A1(n11092), .A2(n11091), .B1(n11090), .B2(n11089), .ZN(
        n11336) );
  NAND2_X2 U7411 ( .A1(n10548), .A2(n12326), .ZN(n10653) );
  INV_X4 U7412 ( .A(n9101), .ZN(n6619) );
  AND2_X1 U7413 ( .A1(n8368), .A2(n8369), .ZN(n8412) );
  INV_X1 U7414 ( .A(n8368), .ZN(n8370) );
  NAND2_X1 U7415 ( .A1(n13504), .A2(n13507), .ZN(n8857) );
  AND2_X4 U7416 ( .A1(n9199), .A2(n13158), .ZN(n9256) );
  XNOR2_X2 U7417 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .ZN(n9238) );
  AOI21_X2 U7418 ( .B1(n7062), .B2(n7632), .A(n7061), .ZN(n7630) );
  XNOR2_X2 U7419 ( .A(n11203), .B(n10650), .ZN(n10593) );
  AOI21_X2 U7420 ( .B1(n9626), .B2(n9625), .A(n7160), .ZN(n9642) );
  NAND2_X2 U7421 ( .A1(n9611), .A2(n9612), .ZN(n9626) );
  AOI21_X2 U7422 ( .B1(P1_REG1_REG_3__SCAN_IN), .B2(n14252), .A(n14245), .ZN(
        n10459) );
  AOI21_X2 U7423 ( .B1(n12881), .B2(n9665), .A(n9651), .ZN(n12891) );
  XNOR2_X1 U7424 ( .A(n7647), .B(n7646), .ZN(n14791) );
  NAND2_X1 U7425 ( .A1(n7643), .A2(n15505), .ZN(n7647) );
  NAND2_X4 U7426 ( .A1(n9203), .A2(n9202), .ZN(n9269) );
  NOR2_X2 U7427 ( .A1(n7592), .A2(n7591), .ZN(n7644) );
  NAND2_X2 U7428 ( .A1(n8854), .A2(n8853), .ZN(n13528) );
  NOR2_X2 U7429 ( .A1(n13348), .A2(n6641), .ZN(n14850) );
  NAND2_X2 U7430 ( .A1(n14960), .A2(n15288), .ZN(n14959) );
  XNOR2_X2 U7431 ( .A(n7662), .B(n7661), .ZN(n14960) );
  OAI21_X2 U7432 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(n7601), .A(n7600), .ZN(
        n7620) );
  XNOR2_X2 U7433 ( .A(n9212), .B(n9211), .ZN(n9689) );
  CLKBUF_X1 U7434 ( .A(n12463), .Z(n6784) );
  OAI21_X1 U7435 ( .B1(n13521), .B2(n7241), .A(n7240), .ZN(n8715) );
  AND2_X1 U7436 ( .A1(n14526), .A2(n14082), .ZN(n14508) );
  NAND2_X1 U7437 ( .A1(n12157), .A2(n8845), .ZN(n13619) );
  OAI21_X1 U7438 ( .B1(n14929), .B2(n7224), .A(n7222), .ZN(n14576) );
  NAND2_X1 U7439 ( .A1(n8146), .A2(n8145), .ZN(n14732) );
  NAND2_X1 U7440 ( .A1(n6794), .A2(n6793), .ZN(n9584) );
  CLKBUF_X1 U7441 ( .A(n11869), .Z(n6783) );
  NAND2_X1 U7442 ( .A1(n8638), .A2(n8637), .ZN(n13731) );
  NAND2_X1 U7443 ( .A1(n11834), .A2(n7568), .ZN(n12004) );
  NAND2_X1 U7444 ( .A1(n8466), .A2(n8465), .ZN(n15323) );
  NAND2_X2 U7445 ( .A1(n12523), .A2(n12530), .ZN(n11016) );
  INV_X1 U7446 ( .A(n12392), .ZN(n12360) );
  AND4_X1 U7447 ( .A1(n9261), .A2(n9260), .A3(n9259), .A4(n9258), .ZN(n10709)
         );
  CLKBUF_X1 U7448 ( .A(n14228), .Z(n6624) );
  INV_X1 U7449 ( .A(n10913), .ZN(n11527) );
  INV_X1 U7450 ( .A(n14227), .ZN(n11213) );
  CLKBUF_X2 U7451 ( .A(P2_U3947), .Z(n6623) );
  CLKBUF_X2 U7452 ( .A(n13973), .Z(n14136) );
  INV_X1 U7453 ( .A(n9270), .ZN(n9620) );
  INV_X1 U7454 ( .A(n13380), .ZN(n10599) );
  NAND4_X2 U7455 ( .A1(n7712), .A2(n7711), .A3(n7710), .A4(n7709), .ZN(n14231)
         );
  INV_X2 U7456 ( .A(n9126), .ZN(n6618) );
  INV_X1 U7457 ( .A(n13384), .ZN(n9798) );
  INV_X1 U7458 ( .A(n10639), .ZN(n10727) );
  INV_X2 U7459 ( .A(n7943), .ZN(n13953) );
  INV_X4 U7460 ( .A(n9213), .ZN(n7088) );
  NOR2_X1 U7461 ( .A1(n9721), .A2(P3_IR_REG_26__SCAN_IN), .ZN(n7422) );
  AOI21_X1 U7462 ( .B1(n7069), .B2(n13226), .A(n13349), .ZN(n13228) );
  AND2_X1 U7463 ( .A1(n8309), .A2(n8308), .ZN(n8889) );
  XNOR2_X1 U7464 ( .A(n12714), .B(n12832), .ZN(n12717) );
  AND2_X1 U7465 ( .A1(n7026), .A2(n7024), .ZN(n12714) );
  OR2_X1 U7466 ( .A1(n12873), .A2(n7027), .ZN(n7026) );
  NAND2_X1 U7467 ( .A1(n14393), .A2(n7212), .ZN(n14380) );
  NAND2_X1 U7468 ( .A1(n14393), .A2(n14392), .ZN(n14630) );
  NAND2_X1 U7469 ( .A1(n14818), .A2(n12665), .ZN(n12710) );
  OR2_X1 U7470 ( .A1(n12871), .A2(n12872), .ZN(n12869) );
  AOI21_X2 U7471 ( .B1(n12469), .B2(n12967), .A(n12359), .ZN(n12449) );
  NAND2_X1 U7472 ( .A1(n7508), .A2(n7507), .ZN(n12903) );
  INV_X1 U7473 ( .A(n14820), .ZN(n12857) );
  OAI21_X1 U7474 ( .B1(n13447), .B2(n13456), .A(n13448), .ZN(n13682) );
  NAND2_X1 U7475 ( .A1(n7188), .A2(n6770), .ZN(n14820) );
  OAI22_X1 U7476 ( .A1(n12915), .A2(n9608), .B1(n12458), .B2(n12941), .ZN(
        n12901) );
  NAND2_X1 U7477 ( .A1(n13686), .A2(n8742), .ZN(n13447) );
  OR2_X1 U7478 ( .A1(n12916), .A2(n12914), .ZN(n12917) );
  NAND2_X1 U7479 ( .A1(n14129), .A2(n14128), .ZN(n14715) );
  AND2_X1 U7480 ( .A1(n14474), .A2(n8141), .ZN(n14464) );
  NAND2_X1 U7481 ( .A1(n9617), .A2(n9616), .ZN(n12908) );
  AOI21_X1 U7482 ( .B1(n7242), .B2(n7244), .A(n6686), .ZN(n7240) );
  NAND2_X1 U7483 ( .A1(n8732), .A2(n8731), .ZN(n13688) );
  NAND2_X1 U7484 ( .A1(n8223), .A2(n8222), .ZN(n14627) );
  NAND2_X1 U7485 ( .A1(n8717), .A2(n8716), .ZN(n13694) );
  NAND2_X1 U7486 ( .A1(n8194), .A2(n8193), .ZN(n14419) );
  NAND2_X1 U7487 ( .A1(n7257), .A2(n7255), .ZN(n13544) );
  NAND2_X1 U7488 ( .A1(n14507), .A2(n8283), .ZN(n14495) );
  NAND2_X1 U7489 ( .A1(n8180), .A2(n8179), .ZN(n14724) );
  XNOR2_X1 U7490 ( .A(n8204), .B(n8203), .ZN(n13799) );
  OAI21_X1 U7491 ( .B1(n8191), .B2(n8190), .A(n8189), .ZN(n8204) );
  NAND2_X1 U7492 ( .A1(n8175), .A2(n8174), .ZN(n8191) );
  NAND2_X1 U7493 ( .A1(n8160), .A2(n8159), .ZN(n14728) );
  NAND2_X2 U7494 ( .A1(n8697), .A2(n8696), .ZN(n13703) );
  NOR2_X1 U7495 ( .A1(n13010), .A2(n9517), .ZN(n7003) );
  NAND2_X1 U7496 ( .A1(n8607), .A2(n8606), .ZN(n13629) );
  NAND2_X1 U7497 ( .A1(n12138), .A2(n7263), .ZN(n8607) );
  NAND2_X1 U7498 ( .A1(n8664), .A2(n8663), .ZN(n13557) );
  NAND2_X1 U7499 ( .A1(n6798), .A2(n14965), .ZN(n14971) );
  NAND2_X1 U7500 ( .A1(n8575), .A2(n7265), .ZN(n12138) );
  XNOR2_X1 U7501 ( .A(n8173), .B(SI_24_), .ZN(n8170) );
  XNOR2_X1 U7502 ( .A(n13726), .B(n13270), .ZN(n13573) );
  NAND2_X1 U7503 ( .A1(n8677), .A2(n8676), .ZN(n13716) );
  OR2_X1 U7504 ( .A1(n12018), .A2(n8573), .ZN(n8575) );
  NAND2_X1 U7505 ( .A1(n14591), .A2(n14057), .ZN(n14565) );
  NAND2_X1 U7506 ( .A1(n7034), .A2(n7032), .ZN(n13021) );
  OAI21_X1 U7507 ( .B1(n11757), .B2(n8530), .A(n8531), .ZN(n11810) );
  NAND2_X1 U7508 ( .A1(n7177), .A2(n7175), .ZN(n9554) );
  NAND2_X1 U7509 ( .A1(n11422), .A2(n11423), .ZN(n11484) );
  NOR2_X1 U7510 ( .A1(n12158), .A2(n7264), .ZN(n7263) );
  NAND2_X1 U7511 ( .A1(n8041), .A2(n8040), .ZN(n14698) );
  AOI21_X1 U7512 ( .B1(n11617), .B2(n7013), .A(n7011), .ZN(n7010) );
  NAND2_X1 U7513 ( .A1(n8616), .A2(n8615), .ZN(n13630) );
  NAND2_X1 U7514 ( .A1(n9522), .A2(n9521), .ZN(n9541) );
  NAND2_X1 U7515 ( .A1(n8021), .A2(n8020), .ZN(n14705) );
  NAND2_X1 U7516 ( .A1(n7338), .A2(n7337), .ZN(n12052) );
  AOI21_X1 U7517 ( .B1(n14993), .B2(P1_REG1_REG_13__SCAN_IN), .A(n14988), .ZN(
        n14998) );
  NAND2_X1 U7518 ( .A1(n7012), .A2(n12682), .ZN(n7011) );
  OAI21_X1 U7519 ( .B1(n11435), .B2(n7292), .A(n7289), .ZN(n11443) );
  NAND2_X1 U7520 ( .A1(n8564), .A2(n8563), .ZN(n14845) );
  NAND2_X1 U7521 ( .A1(n9492), .A2(n9491), .ZN(n9500) );
  CLKBUF_X1 U7522 ( .A(n8032), .Z(n6782) );
  OAI22_X1 U7523 ( .A1(n11258), .A2(n8828), .B1(n10928), .B2(n15323), .ZN(
        n11455) );
  OAI21_X1 U7524 ( .B1(n11207), .B2(n11209), .A(n11206), .ZN(n11295) );
  AOI21_X1 U7525 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(n7605), .A(n7604), .ZN(
        n7616) );
  NAND2_X1 U7526 ( .A1(n8524), .A2(n8523), .ZN(n11783) );
  OAI21_X1 U7527 ( .B1(n15074), .B2(n8269), .A(n8268), .ZN(n11159) );
  NAND2_X1 U7528 ( .A1(n7922), .A2(n7921), .ZN(n14910) );
  NAND2_X2 U7529 ( .A1(n8484), .A2(n8483), .ZN(n15364) );
  NAND2_X2 U7530 ( .A1(n11395), .A2(n11394), .ZN(n15442) );
  OR2_X1 U7531 ( .A1(n9659), .A2(n9648), .ZN(n12881) );
  AND2_X1 U7532 ( .A1(n7050), .A2(n6715), .ZN(n7655) );
  INV_X2 U7533 ( .A(n13643), .ZN(n6620) );
  OAI21_X1 U7534 ( .B1(n14789), .B2(n7648), .A(P2_ADDR_REG_7__SCAN_IN), .ZN(
        n7046) );
  AOI21_X1 U7535 ( .B1(n8266), .B2(n7094), .A(n6665), .ZN(n7093) );
  NOR2_X1 U7536 ( .A1(n7597), .A2(n7596), .ZN(n7652) );
  AND3_X1 U7537 ( .A1(n9237), .A2(n9236), .A3(n9235), .ZN(n9253) );
  NAND2_X1 U7538 ( .A1(n10679), .A2(n11242), .ZN(n7288) );
  INV_X1 U7539 ( .A(n13658), .ZN(n6621) );
  INV_X2 U7540 ( .A(n15354), .ZN(n10651) );
  AND4_X1 U7541 ( .A1(n9274), .A2(n9273), .A3(n9272), .A4(n9271), .ZN(n15451)
         );
  NAND4_X1 U7542 ( .A1(n9245), .A2(n9244), .A3(n9243), .A4(n9242), .ZN(n12741)
         );
  AND2_X1 U7543 ( .A1(n10641), .A2(n10640), .ZN(n10728) );
  AND2_X2 U7544 ( .A1(n12722), .A2(n12528), .ZN(n12647) );
  INV_X1 U7545 ( .A(n10429), .ZN(n12300) );
  OAI211_X1 U7546 ( .C1(n9265), .C2(n9830), .A(n9241), .B(n9240), .ZN(n11370)
         );
  NAND2_X1 U7547 ( .A1(n9529), .A2(n9687), .ZN(n12832) );
  AND2_X1 U7548 ( .A1(n13961), .A2(n14134), .ZN(n13973) );
  CLKBUF_X1 U7549 ( .A(n8438), .Z(n9107) );
  NAND2_X1 U7550 ( .A1(n7763), .A2(n7762), .ZN(n7779) );
  NAND2_X2 U7551 ( .A1(n9250), .A2(n7088), .ZN(n9265) );
  NAND2_X1 U7552 ( .A1(n7752), .A2(n7751), .ZN(n7763) );
  NOR2_X1 U7553 ( .A1(n9791), .A2(n8877), .ZN(n9136) );
  INV_X2 U7554 ( .A(n7732), .ZN(n7794) );
  OR2_X1 U7555 ( .A1(n12320), .A2(n12321), .ZN(n9195) );
  NOR2_X1 U7556 ( .A1(n7588), .A2(n7587), .ZN(n7589) );
  NAND2_X2 U7557 ( .A1(n13162), .A2(n9689), .ZN(n9250) );
  NOR2_X1 U7558 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(n7627), .ZN(n7587) );
  MUX2_X1 U7559 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8319), .S(
        P1_IR_REG_26__SCAN_IN), .Z(n8321) );
  AND2_X1 U7560 ( .A1(n8262), .A2(n8258), .ZN(n10390) );
  CLKBUF_X1 U7561 ( .A(n7943), .Z(n8224) );
  XNOR2_X1 U7562 ( .A(n7063), .B(P3_ADDR_REG_4__SCAN_IN), .ZN(n7627) );
  NOR2_X1 U7563 ( .A1(n9423), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n9438) );
  NAND2_X2 U7564 ( .A1(n8090), .A2(n8251), .ZN(n14917) );
  OR2_X1 U7565 ( .A1(n9494), .A2(P3_IR_REG_16__SCAN_IN), .ZN(n9523) );
  NAND2_X1 U7566 ( .A1(n9221), .A2(n9220), .ZN(n9290) );
  NAND2_X1 U7567 ( .A1(n8251), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8253) );
  INV_X2 U7568 ( .A(n13786), .ZN(n13798) );
  INV_X1 U7569 ( .A(n13791), .ZN(n8369) );
  XNOR2_X1 U7570 ( .A(n7702), .B(n14752), .ZN(n7705) );
  NAND2_X1 U7571 ( .A1(n8257), .A2(n8311), .ZN(n14155) );
  OAI21_X1 U7572 ( .B1(n7628), .B2(P1_ADDR_REG_3__SCAN_IN), .A(n6698), .ZN(
        n7063) );
  NAND2_X1 U7573 ( .A1(n8805), .A2(n8804), .ZN(n8807) );
  NAND2_X1 U7574 ( .A1(n7457), .A2(n7422), .ZN(n9720) );
  NAND2_X1 U7575 ( .A1(n14755), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7702) );
  OR2_X1 U7576 ( .A1(n9366), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n9398) );
  NAND2_X1 U7577 ( .A1(n8089), .A2(n8088), .ZN(n8251) );
  XNOR2_X1 U7578 ( .A(n8259), .B(P1_IR_REG_22__SCAN_IN), .ZN(n14776) );
  AND2_X1 U7579 ( .A1(n7031), .A2(n7458), .ZN(n6809) );
  BUF_X1 U7580 ( .A(n9341), .Z(n9342) );
  NAND2_X1 U7581 ( .A1(n8320), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7102) );
  AND2_X1 U7582 ( .A1(n7187), .A2(n9339), .ZN(n7186) );
  XNOR2_X1 U7583 ( .A(n6863), .B(n6862), .ZN(n10533) );
  CLKBUF_X1 U7584 ( .A(n7993), .Z(n7864) );
  NAND2_X1 U7585 ( .A1(n9748), .A2(n9181), .ZN(n9721) );
  AND2_X1 U7586 ( .A1(n9192), .A2(n9193), .ZN(n7458) );
  AND2_X1 U7587 ( .A1(n6891), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n9246) );
  NAND4_X1 U7588 ( .A1(n7693), .A2(n7692), .A3(n7691), .A4(n7690), .ZN(n7994)
         );
  NAND2_X1 U7589 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(n11832), .ZN(n6793) );
  NOR2_X1 U7590 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .ZN(
        n7687) );
  INV_X1 U7591 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n7690) );
  NOR2_X1 U7592 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n7685) );
  NOR2_X1 U7593 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n7692) );
  NOR2_X1 U7594 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n7689) );
  INV_X4 U7595 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X1 U7596 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n8788) );
  NOR2_X1 U7597 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n8350) );
  INV_X1 U7598 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n8594) );
  INV_X1 U7599 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n8532) );
  INV_X1 U7600 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n8480) );
  INV_X4 U7601 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  INV_X4 U7602 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  INV_X1 U7603 ( .A(P3_IR_REG_5__SCAN_IN), .ZN(n9309) );
  NOR2_X1 U7604 ( .A1(P3_IR_REG_14__SCAN_IN), .A2(P3_IR_REG_12__SCAN_IN), .ZN(
        n9183) );
  NOR2_X1 U7605 ( .A1(P3_IR_REG_11__SCAN_IN), .A2(P3_IR_REG_10__SCAN_IN), .ZN(
        n9184) );
  NOR2_X1 U7606 ( .A1(P3_IR_REG_17__SCAN_IN), .A2(P3_IR_REG_18__SCAN_IN), .ZN(
        n9524) );
  NAND4_X1 U7607 ( .A1(n7798), .A2(n7797), .A3(n7796), .A4(n7795), .ZN(n14228)
         );
  XNOR2_X1 U7608 ( .A(n8765), .B(n9163), .ZN(n13679) );
  CLKBUF_X1 U7609 ( .A(n14765), .Z(n6625) );
  XNOR2_X1 U7610 ( .A(n7102), .B(n7701), .ZN(n14765) );
  NAND2_X1 U7611 ( .A1(n8367), .A2(n8365), .ZN(n13791) );
  INV_X1 U7612 ( .A(n10593), .ZN(n10596) );
  NAND4_X2 U7613 ( .A1(n8402), .A2(n8401), .A3(n8400), .A4(n8399), .ZN(n13382)
         );
  NOR2_X2 U7614 ( .A1(n14791), .A2(n14790), .ZN(n14789) );
  AND2_X1 U7615 ( .A1(n10390), .A2(n10394), .ZN(n10428) );
  INV_X1 U7617 ( .A(n10429), .ZN(n6628) );
  INV_X1 U7618 ( .A(n10429), .ZN(n6629) );
  INV_X1 U7619 ( .A(n6629), .ZN(n12256) );
  INV_X2 U7620 ( .A(n13381), .ZN(n10650) );
  OAI21_X2 U7621 ( .B1(n11295), .B2(n11294), .A(n11293), .ZN(n11301) );
  AOI21_X2 U7622 ( .B1(n13824), .B2(n11179), .A(n11180), .ZN(n11207) );
  BUF_X2 U7623 ( .A(n8413), .Z(n8870) );
  INV_X2 U7624 ( .A(n8413), .ZN(n8389) );
  XNOR2_X2 U7625 ( .A(n8313), .B(P1_IR_REG_25__SCAN_IN), .ZN(n8325) );
  INV_X1 U7626 ( .A(n8424), .ZN(n6630) );
  NAND2_X1 U7627 ( .A1(n12366), .A2(n12920), .ZN(n7312) );
  NOR2_X1 U7628 ( .A1(n13553), .A2(n7260), .ZN(n7259) );
  INV_X1 U7629 ( .A(n8662), .ZN(n7260) );
  OAI21_X1 U7630 ( .B1(n7368), .B2(n6947), .A(n6945), .ZN(n7973) );
  INV_X1 U7631 ( .A(n6946), .ZN(n6945) );
  OAI21_X1 U7632 ( .B1(n7369), .B2(n6947), .A(n7972), .ZN(n6946) );
  NAND2_X1 U7633 ( .A1(n7917), .A2(n7371), .ZN(n7368) );
  NAND2_X1 U7634 ( .A1(n13574), .A2(n7259), .ZN(n7257) );
  NAND2_X1 U7635 ( .A1(n9905), .A2(n9213), .ZN(n14127) );
  INV_X1 U7636 ( .A(n8087), .ZN(n8089) );
  NAND2_X1 U7637 ( .A1(n6839), .A2(n7554), .ZN(n8947) );
  NAND2_X1 U7638 ( .A1(n6642), .A2(n8941), .ZN(n7554) );
  OAI211_X1 U7639 ( .C1(n6642), .C2(n8941), .A(n6840), .B(n6703), .ZN(n6839)
         );
  INV_X1 U7640 ( .A(n8980), .ZN(n6858) );
  OR2_X1 U7641 ( .A1(n7130), .A2(n14058), .ZN(n7129) );
  NOR2_X1 U7642 ( .A1(n14054), .A2(n14053), .ZN(n7130) );
  INV_X1 U7643 ( .A(n14092), .ZN(n7155) );
  NOR2_X1 U7644 ( .A1(n14095), .A2(n14092), .ZN(n7156) );
  OAI21_X1 U7645 ( .B1(n9060), .B2(n7540), .A(n7537), .ZN(n9063) );
  INV_X1 U7646 ( .A(n7541), .ZN(n7540) );
  XNOR2_X1 U7647 ( .A(n14917), .B(n14776), .ZN(n13960) );
  AND2_X1 U7648 ( .A1(n7178), .A2(n6895), .ZN(n6894) );
  NOR2_X1 U7649 ( .A1(n7183), .A2(n7179), .ZN(n7178) );
  NAND2_X1 U7650 ( .A1(n6896), .A2(n9372), .ZN(n6895) );
  INV_X1 U7651 ( .A(n9374), .ZN(n7179) );
  NOR2_X1 U7652 ( .A1(n13969), .A2(n14231), .ZN(n13970) );
  INV_X1 U7653 ( .A(n7936), .ZN(n7373) );
  INV_X1 U7654 ( .A(n7372), .ZN(n7371) );
  OAI21_X1 U7655 ( .B1(n7374), .B2(n7373), .A(n7953), .ZN(n7372) );
  INV_X1 U7656 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n7938) );
  INV_X1 U7657 ( .A(n9199), .ZN(n9203) );
  OR2_X1 U7658 ( .A1(n9758), .A2(n12859), .ZN(n12706) );
  AOI21_X1 U7659 ( .B1(n7019), .B2(n9709), .A(n7017), .ZN(n7016) );
  NAND2_X1 U7660 ( .A1(n6899), .A2(n12511), .ZN(n7017) );
  INV_X1 U7661 ( .A(n6699), .ZN(n7485) );
  NAND2_X1 U7662 ( .A1(n10719), .A2(n11023), .ZN(n12523) );
  INV_X1 U7663 ( .A(n6663), .ZN(n6904) );
  INV_X1 U7664 ( .A(n12872), .ZN(n12874) );
  OR2_X1 U7665 ( .A1(n12492), .A2(n12876), .ZN(n12641) );
  INV_X1 U7666 ( .A(n9453), .ZN(n9722) );
  AND4_X1 U7667 ( .A1(n9524), .A2(n9178), .A3(n9180), .A4(n9179), .ZN(n9748)
         );
  NOR2_X1 U7668 ( .A1(P3_IR_REG_22__SCAN_IN), .A2(P3_IR_REG_21__SCAN_IN), .ZN(
        n9178) );
  NOR2_X1 U7669 ( .A1(P3_IR_REG_20__SCAN_IN), .A2(P3_IR_REG_19__SCAN_IN), .ZN(
        n9180) );
  NOR2_X1 U7670 ( .A1(P3_IR_REG_16__SCAN_IN), .A2(P3_IR_REG_15__SCAN_IN), .ZN(
        n9179) );
  CLKBUF_X1 U7671 ( .A(n9451), .Z(n9452) );
  OAI21_X1 U7672 ( .B1(P2_DATAO_REG_12__SCAN_IN), .B2(n10488), .A(n9415), .ZN(
        n9430) );
  NAND2_X1 U7673 ( .A1(n9341), .A2(n9192), .ZN(n9453) );
  NOR2_X1 U7674 ( .A1(n13507), .A2(n7246), .ZN(n7245) );
  INV_X1 U7675 ( .A(n7249), .ZN(n7246) );
  NOR2_X1 U7676 ( .A1(n7445), .A2(n8851), .ZN(n7438) );
  INV_X1 U7677 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n8352) );
  NOR2_X1 U7678 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(P2_IR_REG_4__SCAN_IN), .ZN(
        n7267) );
  NOR2_X1 U7679 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n7266) );
  AOI21_X1 U7680 ( .B1(n7351), .B2(n13901), .A(n6683), .ZN(n7349) );
  INV_X1 U7681 ( .A(n7351), .ZN(n7350) );
  NOR2_X1 U7682 ( .A1(n14476), .A2(n14732), .ZN(n7092) );
  OR2_X1 U7683 ( .A1(n14518), .A2(n14085), .ZN(n8283) );
  NOR2_X1 U7684 ( .A1(n14590), .A2(n14946), .ZN(n6918) );
  NOR2_X1 U7685 ( .A1(n14592), .A2(n7226), .ZN(n7225) );
  INV_X1 U7686 ( .A(n7990), .ZN(n7226) );
  INV_X1 U7687 ( .A(n7220), .ZN(n7216) );
  NAND2_X1 U7688 ( .A1(n13969), .A2(n7330), .ZN(n13967) );
  NOR2_X1 U7689 ( .A1(n14403), .A2(n14627), .ZN(n14383) );
  NAND2_X1 U7690 ( .A1(n7114), .A2(n7112), .ZN(n14544) );
  AOI21_X1 U7691 ( .B1(n6632), .B2(n14577), .A(n7113), .ZN(n7112) );
  INV_X1 U7692 ( .A(n14071), .ZN(n7113) );
  NAND2_X1 U7693 ( .A1(n11856), .A2(n14185), .ZN(n8279) );
  AND2_X1 U7694 ( .A1(n8189), .A2(n8203), .ZN(n7401) );
  INV_X1 U7695 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n7698) );
  INV_X1 U7696 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n8330) );
  INV_X1 U7697 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n7694) );
  AOI21_X1 U7698 ( .B1(n7310), .B2(n7307), .A(n7306), .ZN(n7305) );
  NOR2_X1 U7699 ( .A1(n12368), .A2(n12904), .ZN(n7306) );
  NOR2_X1 U7700 ( .A1(n6661), .A2(n12484), .ZN(n7307) );
  OR2_X1 U7701 ( .A1(n7297), .A2(n7296), .ZN(n7295) );
  AND2_X1 U7702 ( .A1(n7009), .A2(n7008), .ZN(n10953) );
  AND2_X1 U7703 ( .A1(n9268), .A2(n9267), .ZN(n7008) );
  AND2_X1 U7704 ( .A1(n9203), .A2(n13158), .ZN(n9257) );
  NOR2_X1 U7705 ( .A1(n7470), .A2(n7469), .ZN(n7468) );
  INV_X1 U7706 ( .A(n9652), .ZN(n7469) );
  OR2_X1 U7707 ( .A1(n12958), .A2(n12967), .ZN(n12522) );
  NOR2_X1 U7708 ( .A1(n9481), .A2(n7467), .ZN(n7466) );
  INV_X1 U7709 ( .A(n9465), .ZN(n7467) );
  NAND2_X1 U7710 ( .A1(n11386), .A2(n12670), .ZN(n9699) );
  NAND2_X1 U7711 ( .A1(n14764), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n7190) );
  NAND2_X1 U7712 ( .A1(n12314), .A2(n12315), .ZN(n7191) );
  XNOR2_X1 U7713 ( .A(n9197), .B(P3_IR_REG_29__SCAN_IN), .ZN(n9202) );
  NAND2_X1 U7714 ( .A1(n11772), .A2(n11773), .ZN(n11939) );
  NOR2_X1 U7715 ( .A1(n11777), .A2(n7070), .ZN(n7535) );
  INV_X1 U7716 ( .A(n11769), .ZN(n7070) );
  AND2_X1 U7717 ( .A1(n8786), .A2(n7521), .ZN(n7520) );
  INV_X1 U7718 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n7521) );
  INV_X1 U7719 ( .A(n7258), .ZN(n7256) );
  NAND2_X1 U7720 ( .A1(n8626), .A2(n8625), .ZN(n13609) );
  NOR2_X1 U7721 ( .A1(n11453), .A2(n7237), .ZN(n7236) );
  INV_X1 U7722 ( .A(n8476), .ZN(n7237) );
  AND2_X1 U7723 ( .A1(n8792), .A2(n8791), .ZN(n15337) );
  NAND2_X1 U7724 ( .A1(n8609), .A2(n7573), .ZN(n8778) );
  INV_X1 U7725 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n8775) );
  INV_X1 U7726 ( .A(n14223), .ZN(n11990) );
  NAND2_X1 U7727 ( .A1(n10433), .A2(n10432), .ZN(n10494) );
  NAND2_X1 U7728 ( .A1(n11430), .A2(n7767), .ZN(n6944) );
  NAND2_X1 U7729 ( .A1(n6957), .A2(n14154), .ZN(n6956) );
  NAND2_X1 U7730 ( .A1(n14142), .A2(n6677), .ZN(n6957) );
  AOI22_X1 U7731 ( .A1(n14153), .A2(n14152), .B1(n14151), .B2(n14150), .ZN(
        n14154) );
  NOR2_X1 U7732 ( .A1(n14350), .A2(n14715), .ZN(n14342) );
  AOI21_X1 U7733 ( .B1(n7119), .B2(n7121), .A(n7117), .ZN(n7116) );
  INV_X1 U7734 ( .A(n7119), .ZN(n7118) );
  NAND2_X1 U7735 ( .A1(n14509), .A2(n8112), .ZN(n14493) );
  NAND2_X1 U7736 ( .A1(n7204), .A2(n7203), .ZN(n14509) );
  NOR2_X1 U7737 ( .A1(n14512), .A2(n7207), .ZN(n7203) );
  NAND2_X1 U7738 ( .A1(n6944), .A2(n6941), .ZN(n14067) );
  NOR2_X1 U7739 ( .A1(n14551), .A2(n6942), .ZN(n6941) );
  INV_X1 U7740 ( .A(n8061), .ZN(n6942) );
  NAND2_X1 U7741 ( .A1(n14544), .A2(n14543), .ZN(n14542) );
  NAND2_X1 U7742 ( .A1(n14549), .A2(n8047), .ZN(n8049) );
  NAND2_X1 U7743 ( .A1(n14576), .A2(n8030), .ZN(n14549) );
  INV_X1 U7744 ( .A(n14917), .ZN(n8345) );
  NAND2_X1 U7745 ( .A1(n6925), .A2(n6645), .ZN(n6924) );
  NAND2_X1 U7746 ( .A1(n14627), .A2(n15155), .ZN(n6925) );
  NAND2_X1 U7747 ( .A1(n8093), .A2(n8092), .ZN(n14528) );
  AOI21_X1 U7748 ( .B1(n6929), .B2(n6932), .A(n7902), .ZN(n6926) );
  OAI21_X1 U7749 ( .B1(n7858), .B2(n6934), .A(n7071), .ZN(n7883) );
  NAND2_X1 U7750 ( .A1(n7858), .A2(n7857), .ZN(n7862) );
  OAI21_X1 U7751 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(n7607), .A(n7606), .ZN(
        n7614) );
  AOI21_X1 U7752 ( .B1(n14974), .B2(n14975), .A(n7055), .ZN(n7054) );
  INV_X1 U7753 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n7055) );
  XNOR2_X1 U7754 ( .A(n12358), .B(n12356), .ZN(n12469) );
  AOI21_X1 U7755 ( .B1(n14334), .B2(n15012), .A(n14917), .ZN(n6813) );
  NAND2_X1 U7756 ( .A1(n14337), .A2(n14917), .ZN(n6815) );
  OAI21_X1 U7757 ( .B1(n14960), .B2(n7059), .A(n7057), .ZN(n14961) );
  AOI22_X1 U7758 ( .A1(n8909), .A2(n13382), .B1(n8910), .B2(n15354), .ZN(n8917) );
  NAND2_X1 U7759 ( .A1(n14009), .A2(n7144), .ZN(n7143) );
  INV_X1 U7760 ( .A(n14008), .ZN(n7144) );
  NAND2_X1 U7761 ( .A1(n14020), .A2(n7139), .ZN(n7138) );
  INV_X1 U7762 ( .A(n14019), .ZN(n7139) );
  AOI21_X1 U7763 ( .B1(n8947), .B2(n8946), .A(n8944), .ZN(n8945) );
  NAND2_X1 U7764 ( .A1(n14031), .A2(n7149), .ZN(n7148) );
  INV_X1 U7765 ( .A(n14030), .ZN(n7149) );
  OR2_X1 U7766 ( .A1(n8962), .A2(n8961), .ZN(n8968) );
  NAND2_X1 U7767 ( .A1(n14042), .A2(n7134), .ZN(n7133) );
  INV_X1 U7768 ( .A(n14041), .ZN(n7134) );
  NAND2_X1 U7769 ( .A1(n6854), .A2(n6853), .ZN(n8984) );
  NOR2_X1 U7770 ( .A1(n8972), .A2(n8977), .ZN(n7561) );
  INV_X1 U7771 ( .A(n7128), .ZN(n7127) );
  OAI21_X1 U7772 ( .B1(n7129), .B2(n7131), .A(n6637), .ZN(n7128) );
  AND2_X1 U7773 ( .A1(n14167), .A2(n14056), .ZN(n7131) );
  INV_X1 U7774 ( .A(n9027), .ZN(n7558) );
  AND2_X1 U7775 ( .A1(n6726), .A2(n6846), .ZN(n6845) );
  NAND2_X1 U7776 ( .A1(n9022), .A2(n6669), .ZN(n6846) );
  NAND2_X1 U7777 ( .A1(n6660), .A2(n6852), .ZN(n6850) );
  INV_X1 U7778 ( .A(n9047), .ZN(n7557) );
  INV_X1 U7779 ( .A(n9059), .ZN(n7545) );
  NAND2_X1 U7780 ( .A1(n6937), .A2(n6935), .ZN(n14103) );
  NAND2_X1 U7781 ( .A1(n14099), .A2(n6936), .ZN(n6935) );
  AND2_X1 U7782 ( .A1(n7542), .A2(n9065), .ZN(n7541) );
  NAND2_X1 U7783 ( .A1(n7544), .A2(n7543), .ZN(n7542) );
  NAND2_X1 U7784 ( .A1(n7545), .A2(n6670), .ZN(n7543) );
  INV_X1 U7785 ( .A(n14109), .ZN(n7157) );
  NOR2_X1 U7786 ( .A1(n14112), .A2(n14109), .ZN(n7158) );
  AND2_X1 U7787 ( .A1(n14115), .A2(n6965), .ZN(n6964) );
  INV_X1 U7788 ( .A(n14113), .ZN(n6965) );
  AND2_X1 U7789 ( .A1(n12857), .A2(n12727), .ZN(n12711) );
  INV_X1 U7790 ( .A(n7416), .ZN(n7415) );
  OAI21_X1 U7791 ( .B1(n12686), .B2(n7417), .A(n13033), .ZN(n7416) );
  NAND2_X1 U7792 ( .A1(n15458), .A2(n10781), .ZN(n12534) );
  INV_X1 U7793 ( .A(n7197), .ZN(n7195) );
  AOI21_X1 U7794 ( .B1(n9583), .B2(n7198), .A(n9600), .ZN(n7197) );
  INV_X1 U7795 ( .A(n7198), .ZN(n7194) );
  INV_X1 U7796 ( .A(P3_IR_REG_6__SCAN_IN), .ZN(n9188) );
  INV_X1 U7797 ( .A(n8909), .ZN(n9126) );
  INV_X1 U7798 ( .A(n8910), .ZN(n9101) );
  INV_X1 U7799 ( .A(n8858), .ZN(n7437) );
  OR2_X1 U7800 ( .A1(n13990), .A2(n11192), .ZN(n8266) );
  NAND2_X1 U7801 ( .A1(n7729), .A2(n9941), .ZN(n7228) );
  NAND2_X1 U7802 ( .A1(n8077), .A2(n10725), .ZN(n8098) );
  OAI22_X1 U7803 ( .A1(n8017), .A2(n8016), .B1(n8015), .B2(SI_15_), .ZN(n8032)
         );
  OAI21_X1 U7804 ( .B1(n9213), .B2(n9822), .A(n7077), .ZN(n7076) );
  NAND4_X1 U7805 ( .A1(n14341), .A2(n13434), .A3(n7359), .A4(
        P3_ADDR_REG_19__SCAN_IN), .ZN(n7357) );
  INV_X1 U7806 ( .A(P1_RD_REG_SCAN_IN), .ZN(n7359) );
  INV_X1 U7807 ( .A(n9765), .ZN(n7287) );
  NAND2_X1 U7808 ( .A1(n11322), .A2(n9765), .ZN(n12703) );
  AND2_X1 U7809 ( .A1(n12708), .A2(n6824), .ZN(n12713) );
  NOR2_X1 U7810 ( .A1(n12709), .A2(n6825), .ZN(n6824) );
  NOR2_X1 U7811 ( .A1(n12857), .A2(n12851), .ZN(n6825) );
  NAND2_X1 U7812 ( .A1(n11918), .A2(n11919), .ZN(n11920) );
  NAND2_X1 U7813 ( .A1(n11920), .A2(n11926), .ZN(n12744) );
  NAND2_X1 U7814 ( .A1(n12795), .A2(n12796), .ZN(n12818) );
  NOR2_X1 U7815 ( .A1(n9618), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n9631) );
  OR2_X1 U7816 ( .A1(n9603), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n9618) );
  NOR2_X1 U7817 ( .A1(n12995), .A2(n7502), .ZN(n7501) );
  INV_X1 U7818 ( .A(n9518), .ZN(n7502) );
  OR2_X1 U7819 ( .A1(n13139), .A2(n13003), .ZN(n12621) );
  NAND2_X1 U7820 ( .A1(n7464), .A2(n6649), .ZN(n7463) );
  INV_X1 U7821 ( .A(n7466), .ZN(n7464) );
  INV_X1 U7822 ( .A(n7412), .ZN(n7033) );
  AOI21_X1 U7823 ( .B1(n7415), .B2(n7417), .A(n7413), .ZN(n7412) );
  AND2_X1 U7824 ( .A1(n7415), .A2(n7037), .ZN(n7036) );
  NAND2_X1 U7825 ( .A1(n7040), .A2(n7038), .ZN(n7037) );
  INV_X1 U7826 ( .A(n7042), .ZN(n7038) );
  NOR2_X1 U7827 ( .A1(n12126), .A2(n7043), .ZN(n7042) );
  INV_X1 U7828 ( .A(n12591), .ZN(n7043) );
  AOI21_X1 U7829 ( .B1(n7042), .B2(n9704), .A(n7041), .ZN(n7040) );
  INV_X1 U7830 ( .A(n12596), .ZN(n7041) );
  AOI21_X1 U7831 ( .B1(n7483), .B2(n7482), .A(n7481), .ZN(n7480) );
  INV_X1 U7832 ( .A(n7486), .ZN(n7482) );
  AOI21_X1 U7833 ( .B1(n9701), .B2(n7410), .A(n7409), .ZN(n7408) );
  INV_X1 U7834 ( .A(n9700), .ZN(n7410) );
  INV_X1 U7835 ( .A(n9702), .ZN(n7409) );
  NAND2_X1 U7836 ( .A1(n12534), .A2(n12533), .ZN(n9698) );
  INV_X1 U7837 ( .A(n7182), .ZN(n7181) );
  NAND2_X1 U7838 ( .A1(n6894), .A2(n6897), .ZN(n6893) );
  OAI21_X1 U7839 ( .B1(n9385), .B2(n7183), .A(n9405), .ZN(n7182) );
  NOR2_X1 U7840 ( .A1(n13247), .A2(n13190), .ZN(n7528) );
  NAND2_X1 U7841 ( .A1(n6837), .A2(n7546), .ZN(n6836) );
  NOR2_X1 U7842 ( .A1(n9094), .A2(n7547), .ZN(n7546) );
  NAND2_X1 U7843 ( .A1(n6695), .A2(n7548), .ZN(n7547) );
  INV_X1 U7844 ( .A(n7245), .ZN(n7244) );
  XNOR2_X1 U7845 ( .A(n13703), .B(n13281), .ZN(n9158) );
  NOR2_X1 U7846 ( .A1(n7443), .A2(n8851), .ZN(n7440) );
  INV_X1 U7847 ( .A(n13573), .ZN(n7443) );
  OAI21_X1 U7848 ( .B1(n13573), .B2(n8849), .A(n6673), .ZN(n7445) );
  NOR2_X1 U7849 ( .A1(n8847), .A2(n7455), .ZN(n7454) );
  INV_X1 U7850 ( .A(n8846), .ZN(n7455) );
  NOR2_X1 U7851 ( .A1(n12020), .A2(n14845), .ZN(n7274) );
  NAND2_X1 U7852 ( .A1(n13784), .A2(n9085), .ZN(n7381) );
  INV_X1 U7853 ( .A(n10585), .ZN(n10548) );
  XNOR2_X1 U7854 ( .A(P2_IR_REG_21__SCAN_IN), .B(P2_IR_REG_31__SCAN_IN), .ZN(
        n7519) );
  CLKBUF_X1 U7855 ( .A(n8609), .Z(n8596) );
  INV_X1 U7856 ( .A(n7323), .ZN(n7321) );
  INV_X1 U7857 ( .A(n8291), .ZN(n7122) );
  AND2_X1 U7858 ( .A1(n8295), .A2(n8236), .ZN(n14372) );
  INV_X1 U7859 ( .A(n7098), .ZN(n7097) );
  OAI21_X1 U7860 ( .B1(n8285), .B2(n7099), .A(n14458), .ZN(n7098) );
  INV_X1 U7861 ( .A(n8286), .ZN(n7099) );
  NAND2_X1 U7862 ( .A1(n14674), .A2(n6915), .ZN(n6914) );
  OR2_X1 U7863 ( .A1(n14705), .A2(n14582), .ZN(n8030) );
  OR2_X1 U7864 ( .A1(n14590), .A2(n14920), .ZN(n14057) );
  AND2_X1 U7865 ( .A1(n14051), .A2(n14055), .ZN(n14167) );
  NOR2_X1 U7866 ( .A1(n7202), .A2(n15117), .ZN(n7201) );
  INV_X1 U7867 ( .A(n7776), .ZN(n7202) );
  INV_X1 U7868 ( .A(n7228), .ZN(n7227) );
  NAND2_X1 U7869 ( .A1(n7739), .A2(n7729), .ZN(n14169) );
  NOR2_X1 U7870 ( .A1(n14419), .A2(n14629), .ZN(n6921) );
  NOR2_X1 U7871 ( .A1(n13999), .A2(n15083), .ZN(n7090) );
  AND2_X1 U7872 ( .A1(n14155), .A2(n8305), .ZN(n8344) );
  INV_X1 U7873 ( .A(n14776), .ZN(n8305) );
  NAND2_X1 U7874 ( .A1(n8240), .A2(n8239), .ZN(n9077) );
  NAND2_X1 U7875 ( .A1(n8191), .A2(n7401), .ZN(n7399) );
  AOI21_X1 U7876 ( .B1(n8190), .B2(n7401), .A(n6763), .ZN(n7400) );
  NAND2_X1 U7877 ( .A1(n8099), .A2(n8098), .ZN(n8127) );
  XNOR2_X1 U7878 ( .A(n8127), .B(SI_20_), .ZN(n8113) );
  AND2_X1 U7879 ( .A1(n8051), .A2(n8034), .ZN(n7382) );
  AOI21_X1 U7880 ( .B1(n6950), .B2(n7382), .A(n6949), .ZN(n6948) );
  INV_X1 U7881 ( .A(n8070), .ZN(n6949) );
  INV_X1 U7882 ( .A(n8031), .ZN(n6950) );
  NAND2_X1 U7883 ( .A1(n8032), .A2(n8031), .ZN(n8035) );
  XNOR2_X1 U7884 ( .A(n8015), .B(SI_15_), .ZN(n8016) );
  AOI21_X1 U7885 ( .B1(n7371), .B2(n7373), .A(n6700), .ZN(n7369) );
  NOR2_X1 U7886 ( .A1(n7937), .A2(n7375), .ZN(n7374) );
  INV_X1 U7887 ( .A(n7916), .ZN(n7375) );
  NAND2_X1 U7888 ( .A1(n7076), .A2(SI_4_), .ZN(n7800) );
  INV_X1 U7889 ( .A(n7063), .ZN(n7586) );
  INV_X1 U7890 ( .A(P3_ADDR_REG_5__SCAN_IN), .ZN(n7590) );
  NOR2_X1 U7891 ( .A1(n7626), .A2(n10374), .ZN(n7596) );
  INV_X1 U7892 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n7621) );
  NOR2_X1 U7893 ( .A1(n7618), .A2(n7619), .ZN(n7604) );
  INV_X1 U7894 ( .A(n11520), .ZN(n7293) );
  AND2_X1 U7895 ( .A1(n12403), .A2(n7284), .ZN(n7283) );
  OR2_X1 U7896 ( .A1(n12462), .A2(n7285), .ZN(n7284) );
  INV_X1 U7897 ( .A(n12354), .ZN(n7285) );
  NAND2_X1 U7898 ( .A1(n12381), .A2(n12351), .ZN(n12463) );
  NAND2_X1 U7899 ( .A1(n6773), .A2(n6772), .ZN(n11869) );
  INV_X1 U7900 ( .A(n11793), .ZN(n6772) );
  INV_X1 U7901 ( .A(n11792), .ZN(n6773) );
  INV_X1 U7902 ( .A(n12031), .ZN(n7296) );
  NAND2_X1 U7903 ( .A1(n6712), .A2(n7312), .ZN(n7310) );
  NAND2_X1 U7904 ( .A1(n12365), .A2(n12364), .ZN(n7311) );
  XNOR2_X1 U7905 ( .A(n7164), .B(n12847), .ZN(n7163) );
  NOR2_X1 U7906 ( .A1(n12699), .A2(n12700), .ZN(n7165) );
  NAND2_X1 U7907 ( .A1(n9720), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9212) );
  NAND2_X1 U7908 ( .A1(n6777), .A2(n6776), .ZN(n10520) );
  OR2_X1 U7909 ( .A1(n13165), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n6777) );
  NAND2_X1 U7910 ( .A1(n13165), .A2(n10797), .ZN(n6776) );
  NAND2_X1 U7911 ( .A1(n10520), .A2(n10798), .ZN(n10788) );
  XNOR2_X1 U7912 ( .A(n6870), .B(n10874), .ZN(n10867) );
  NAND2_X1 U7913 ( .A1(n10904), .A2(n10905), .ZN(n11078) );
  NAND2_X1 U7914 ( .A1(n11075), .A2(n6982), .ZN(n6981) );
  NAND2_X1 U7915 ( .A1(n11076), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n6982) );
  XNOR2_X1 U7916 ( .A(n12764), .B(n6775), .ZN(n12747) );
  AOI21_X1 U7917 ( .B1(n12756), .B2(n12755), .A(n12754), .ZN(n12781) );
  NAND2_X1 U7918 ( .A1(n12791), .A2(n6868), .ZN(n6867) );
  OR2_X1 U7919 ( .A1(n12794), .A2(n12792), .ZN(n6868) );
  NAND2_X1 U7920 ( .A1(n6900), .A2(n6902), .ZN(n6905) );
  NOR2_X1 U7921 ( .A1(n12874), .A2(n6903), .ZN(n6902) );
  NOR2_X1 U7922 ( .A1(n6904), .A2(n12641), .ZN(n6903) );
  INV_X1 U7923 ( .A(n9666), .ZN(n7470) );
  INV_X1 U7924 ( .A(n6905), .ZN(n12873) );
  INV_X1 U7925 ( .A(n7504), .ZN(n7503) );
  OAI21_X1 U7926 ( .B1(n7505), .B2(n9624), .A(n9640), .ZN(n7504) );
  AND2_X1 U7927 ( .A1(n12652), .A2(n12646), .ZN(n12872) );
  NAND2_X1 U7928 ( .A1(n7016), .A2(n7018), .ZN(n12890) );
  NAND2_X1 U7929 ( .A1(n12917), .A2(n12517), .ZN(n12900) );
  AOI21_X1 U7930 ( .B1(n7418), .B2(n6671), .A(n7004), .ZN(n7007) );
  NAND2_X1 U7931 ( .A1(n7005), .A2(n6689), .ZN(n7004) );
  OAI21_X1 U7932 ( .B1(n13002), .B2(n7500), .A(n7497), .ZN(n9553) );
  INV_X1 U7933 ( .A(n9540), .ZN(n7500) );
  INV_X1 U7934 ( .A(n12984), .ZN(n7418) );
  OAI21_X1 U7935 ( .B1(n7003), .B2(n7002), .A(n12621), .ZN(n12984) );
  INV_X1 U7936 ( .A(n12612), .ZN(n7002) );
  NAND2_X1 U7937 ( .A1(n13002), .A2(n7501), .ZN(n12987) );
  NAND2_X1 U7938 ( .A1(n9705), .A2(n12608), .ZN(n13010) );
  NAND2_X1 U7939 ( .A1(n7035), .A2(n7040), .ZN(n12152) );
  NAND2_X1 U7940 ( .A1(n12078), .A2(n7042), .ZN(n7035) );
  NAND2_X1 U7941 ( .A1(n12071), .A2(n12587), .ZN(n12078) );
  NOR2_X1 U7942 ( .A1(n12681), .A2(n7487), .ZN(n7486) );
  INV_X1 U7943 ( .A(n9396), .ZN(n7487) );
  NAND2_X1 U7944 ( .A1(n12072), .A2(n12681), .ZN(n12071) );
  AND4_X1 U7945 ( .A1(n9403), .A2(n9402), .A3(n9401), .A4(n9400), .ZN(n12081)
         );
  INV_X1 U7946 ( .A(n7408), .ZN(n7015) );
  INV_X1 U7947 ( .A(n7014), .ZN(n7013) );
  OAI21_X1 U7948 ( .B1(n7015), .B2(n12567), .A(n7405), .ZN(n7014) );
  AOI21_X1 U7949 ( .B1(n7408), .B2(n7411), .A(n7406), .ZN(n7405) );
  INV_X1 U7950 ( .A(n9701), .ZN(n7411) );
  NAND2_X1 U7951 ( .A1(n11617), .A2(n12567), .ZN(n11731) );
  NOR2_X1 U7952 ( .A1(n12671), .A2(n7476), .ZN(n7475) );
  AND2_X1 U7953 ( .A1(n12567), .A2(n12566), .ZN(n12671) );
  AND2_X1 U7954 ( .A1(n12676), .A2(n9318), .ZN(n7496) );
  NAND2_X1 U7955 ( .A1(n9317), .A2(n9316), .ZN(n11310) );
  NOR2_X1 U7956 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(P3_REG3_REG_3__SCAN_IN), 
        .ZN(n9298) );
  AOI21_X1 U7957 ( .B1(n12677), .B2(n7404), .A(n7403), .ZN(n7402) );
  INV_X1 U7958 ( .A(n12533), .ZN(n7404) );
  INV_X1 U7959 ( .A(n12542), .ZN(n7403) );
  AND4_X1 U7960 ( .A1(n9303), .A2(n9302), .A3(n9301), .A4(n9300), .ZN(n11437)
         );
  NAND2_X1 U7961 ( .A1(n10953), .A2(n10709), .ZN(n12533) );
  INV_X1 U7962 ( .A(n9698), .ZN(n15448) );
  NAND2_X1 U7963 ( .A1(n9255), .A2(n9254), .ZN(n15446) );
  NAND2_X1 U7964 ( .A1(n12741), .A2(n10913), .ZN(n11366) );
  INV_X1 U7965 ( .A(n15452), .ZN(n13027) );
  NAND2_X1 U7966 ( .A1(n9752), .A2(n12715), .ZN(n13032) );
  NAND2_X1 U7967 ( .A1(n11365), .A2(n11364), .ZN(n11393) );
  AND2_X1 U7968 ( .A1(n11363), .A2(n11362), .ZN(n11364) );
  AOI21_X1 U7969 ( .B1(n12334), .B2(n15477), .A(n9696), .ZN(n7491) );
  NAND2_X1 U7970 ( .A1(n9675), .A2(n9674), .ZN(n9758) );
  NAND2_X1 U7971 ( .A1(n9474), .A2(n9473), .ZN(n13093) );
  NOR2_X1 U7972 ( .A1(n9755), .A2(n13150), .ZN(n10705) );
  AND2_X1 U7973 ( .A1(n10671), .A2(n13151), .ZN(n10702) );
  INV_X1 U7974 ( .A(n15486), .ZN(n15479) );
  AOI21_X1 U7975 ( .B1(n9730), .B2(n12092), .A(n6828), .ZN(n9846) );
  INV_X1 U7976 ( .A(n12659), .ZN(n6822) );
  AND2_X1 U7977 ( .A1(n14773), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n7160) );
  INV_X1 U7978 ( .A(n9721), .ZN(n7456) );
  AND2_X1 U7979 ( .A1(n9723), .A2(n9722), .ZN(n9724) );
  NAND2_X1 U7980 ( .A1(n12321), .A2(n9185), .ZN(n6819) );
  NOR2_X1 U7981 ( .A1(n9721), .A2(n9187), .ZN(n7459) );
  NAND2_X1 U7982 ( .A1(n7277), .A2(n7276), .ZN(n9684) );
  INV_X1 U7983 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n7276) );
  INV_X1 U7984 ( .A(n9687), .ZN(n7277) );
  NAND2_X1 U7985 ( .A1(n9502), .A2(n6805), .ZN(n9520) );
  NAND2_X1 U7986 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(n6806), .ZN(n6805) );
  NAND2_X1 U7987 ( .A1(n9749), .A2(n9455), .ZN(n9494) );
  NAND2_X1 U7988 ( .A1(n7169), .A2(n7168), .ZN(n9468) );
  INV_X1 U7989 ( .A(n7170), .ZN(n7169) );
  OAI21_X1 U7990 ( .B1(n9431), .B2(n7173), .A(n9449), .ZN(n7170) );
  NAND2_X1 U7991 ( .A1(n9375), .A2(n9374), .ZN(n9386) );
  NAND2_X1 U7992 ( .A1(n9373), .A2(n9372), .ZN(n9375) );
  XNOR2_X1 U7993 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .ZN(n9339) );
  NAND2_X1 U7994 ( .A1(n6890), .A2(n9222), .ZN(n9306) );
  NOR2_X1 U7995 ( .A1(n9266), .A2(n12321), .ZN(n6863) );
  OR2_X1 U7996 ( .A1(n13222), .A2(n13221), .ZN(n13223) );
  NAND2_X1 U7997 ( .A1(n7517), .A2(n6816), .ZN(n11421) );
  AND2_X1 U7998 ( .A1(n11346), .A2(n11340), .ZN(n6816) );
  INV_X1 U7999 ( .A(n13364), .ZN(n13270) );
  OR2_X1 U8000 ( .A1(n13237), .A2(n13236), .ZN(n13205) );
  INV_X1 U8001 ( .A(n7528), .ZN(n7527) );
  NAND2_X1 U8002 ( .A1(n13194), .A2(n13193), .ZN(n7529) );
  NAND2_X1 U8003 ( .A1(n13202), .A2(n13201), .ZN(n13234) );
  XNOR2_X1 U8004 ( .A(n13203), .B(n6664), .ZN(n13202) );
  XNOR2_X1 U8005 ( .A(n10652), .B(n10651), .ZN(n10654) );
  AND2_X1 U8006 ( .A1(n6640), .A2(n13325), .ZN(n7079) );
  INV_X1 U8007 ( .A(n8424), .ZN(n8748) );
  OAI22_X1 U8008 ( .A1(n6630), .A2(P2_REG3_REG_3__SCAN_IN), .B1(n6626), .B2(
        n10314), .ZN(n7235) );
  NAND2_X1 U8009 ( .A1(n8368), .A2(n13791), .ZN(n8413) );
  NAND2_X1 U8010 ( .A1(n8360), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8377) );
  AND2_X1 U8011 ( .A1(n8608), .A2(n7513), .ZN(n7512) );
  INV_X1 U8012 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n7513) );
  AND2_X1 U8013 ( .A1(n13479), .A2(n6721), .ZN(n13441) );
  OR2_X1 U8014 ( .A1(n13455), .A2(n13254), .ZN(n6788) );
  INV_X1 U8015 ( .A(n9161), .ZN(n13456) );
  AOI21_X1 U8016 ( .B1(n7245), .B2(n7243), .A(n6681), .ZN(n7242) );
  INV_X1 U8017 ( .A(n6655), .ZN(n7243) );
  NAND2_X1 U8018 ( .A1(n8857), .A2(n8856), .ZN(n13492) );
  INV_X1 U8019 ( .A(n7244), .ZN(n7239) );
  OR2_X1 U8020 ( .A1(n13524), .A2(n13361), .ZN(n7249) );
  NAND2_X1 U8021 ( .A1(n7248), .A2(n6655), .ZN(n7247) );
  INV_X1 U8022 ( .A(n13521), .ZN(n7248) );
  INV_X1 U8023 ( .A(n9158), .ZN(n13507) );
  AOI21_X1 U8024 ( .B1(n7259), .B2(n8661), .A(n6701), .ZN(n7258) );
  INV_X1 U8025 ( .A(n7445), .ZN(n7444) );
  OR2_X1 U8026 ( .A1(n8850), .A2(n13573), .ZN(n7442) );
  NAND2_X1 U8027 ( .A1(n8649), .A2(n8648), .ZN(n13574) );
  NOR2_X1 U8028 ( .A1(n13597), .A2(n7253), .ZN(n7252) );
  INV_X1 U8029 ( .A(n8623), .ZN(n7253) );
  NAND2_X1 U8030 ( .A1(n13629), .A2(n13620), .ZN(n7254) );
  AND2_X1 U8031 ( .A1(n12141), .A2(n8574), .ZN(n7265) );
  NAND2_X1 U8032 ( .A1(n8551), .A2(n8550), .ZN(n11973) );
  INV_X1 U8033 ( .A(n7447), .ZN(n7446) );
  OAI21_X1 U8034 ( .B1(n11811), .B2(n7448), .A(n6709), .ZN(n7447) );
  NAND2_X1 U8035 ( .A1(n11113), .A2(n8462), .ZN(n11255) );
  NOR2_X1 U8036 ( .A1(n13652), .A2(n15354), .ZN(n13650) );
  CLKBUF_X1 U8037 ( .A(n8815), .Z(n8816) );
  NAND2_X1 U8038 ( .A1(n7381), .A2(n9086), .ZN(n9128) );
  NAND2_X1 U8039 ( .A1(n8707), .A2(n8706), .ZN(n13698) );
  OAI21_X1 U8040 ( .B1(n8801), .B2(P2_IR_REG_22__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8796) );
  INV_X1 U8041 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n8349) );
  OR2_X1 U8042 ( .A1(n8535), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n8559) );
  AND2_X1 U8043 ( .A1(n13931), .A2(n7335), .ZN(n7334) );
  OR2_X1 U8044 ( .A1(n13864), .A2(n7336), .ZN(n7335) );
  INV_X1 U8045 ( .A(n12283), .ZN(n7336) );
  NAND2_X1 U8046 ( .A1(n13893), .A2(n6676), .ZN(n13843) );
  NOR2_X1 U8047 ( .A1(n7321), .A2(n7315), .ZN(n7314) );
  INV_X1 U8048 ( .A(n12055), .ZN(n7315) );
  NOR2_X1 U8049 ( .A1(n7321), .A2(n7317), .ZN(n7316) );
  AND2_X1 U8050 ( .A1(n12061), .A2(n7318), .ZN(n7317) );
  INV_X1 U8051 ( .A(n12054), .ZN(n7318) );
  INV_X1 U8052 ( .A(n12061), .ZN(n7319) );
  NOR2_X1 U8053 ( .A1(n13858), .A2(n13859), .ZN(n13857) );
  OR2_X1 U8054 ( .A1(n13911), .A2(n7328), .ZN(n7327) );
  INV_X1 U8055 ( .A(n12262), .ZN(n7328) );
  NAND2_X1 U8056 ( .A1(n7342), .A2(n7344), .ZN(n7337) );
  AOI21_X1 U8057 ( .B1(n14233), .B2(n12301), .A(n10398), .ZN(n10399) );
  INV_X1 U8058 ( .A(n10397), .ZN(n10398) );
  NAND2_X1 U8059 ( .A1(n14124), .A2(n14123), .ZN(n14141) );
  NOR2_X1 U8060 ( .A1(n14198), .A2(n14160), .ZN(n6955) );
  AND2_X1 U8061 ( .A1(n7705), .A2(n7706), .ZN(n7943) );
  OR2_X1 U8062 ( .A1(n7809), .A2(P1_IR_REG_5__SCAN_IN), .ZN(n7845) );
  NAND2_X1 U8063 ( .A1(n14383), .A2(n14365), .ZN(n14350) );
  NAND2_X1 U8064 ( .A1(n6639), .A2(n14639), .ZN(n14413) );
  OR2_X1 U8065 ( .A1(n14423), .A2(n14430), .ZN(n14425) );
  NOR2_X1 U8066 ( .A1(n14447), .A2(n7232), .ZN(n7231) );
  INV_X1 U8067 ( .A(n8153), .ZN(n7232) );
  NAND2_X1 U8068 ( .A1(n14464), .A2(n14463), .ZN(n14462) );
  NAND2_X1 U8069 ( .A1(n14494), .A2(n8285), .ZN(n14486) );
  NAND2_X1 U8070 ( .A1(n14495), .A2(n14496), .ZN(n14494) );
  NAND2_X1 U8071 ( .A1(n7211), .A2(n8068), .ZN(n7208) );
  INV_X1 U8072 ( .A(n8068), .ZN(n7209) );
  AND2_X1 U8073 ( .A1(n8283), .A2(n8111), .ZN(n14512) );
  NOR2_X1 U8074 ( .A1(n14523), .A2(n7101), .ZN(n7100) );
  INV_X1 U8075 ( .A(n14067), .ZN(n7101) );
  AND2_X1 U8076 ( .A1(n14078), .A2(n14067), .ZN(n14543) );
  INV_X1 U8077 ( .A(n7223), .ZN(n7222) );
  OAI21_X1 U8078 ( .B1(n7225), .B2(n7224), .A(n14577), .ZN(n7223) );
  INV_X1 U8079 ( .A(n8014), .ZN(n7224) );
  NAND2_X1 U8080 ( .A1(n7105), .A2(n7103), .ZN(n14591) );
  NOR2_X1 U8081 ( .A1(n8280), .A2(n7104), .ZN(n7103) );
  NAND2_X1 U8082 ( .A1(n8279), .A2(n7106), .ZN(n7105) );
  AND2_X1 U8083 ( .A1(n14051), .A2(n8278), .ZN(n7106) );
  NAND2_X1 U8084 ( .A1(n14929), .A2(n7225), .ZN(n14581) );
  NAND2_X1 U8085 ( .A1(n8277), .A2(n8276), .ZN(n11856) );
  NOR2_X1 U8086 ( .A1(n7933), .A2(n7221), .ZN(n7220) );
  INV_X1 U8087 ( .A(n7914), .ZN(n7221) );
  INV_X1 U8088 ( .A(n7932), .ZN(n7218) );
  NAND2_X1 U8089 ( .A1(n11634), .A2(n11636), .ZN(n7915) );
  INV_X1 U8090 ( .A(n8272), .ZN(n7109) );
  INV_X1 U8091 ( .A(n14181), .ZN(n11636) );
  NAND2_X1 U8092 ( .A1(n7111), .A2(n7110), .ZN(n14596) );
  NOR2_X1 U8093 ( .A1(n10974), .A2(n13990), .ZN(n11040) );
  NAND2_X1 U8094 ( .A1(n10749), .A2(n14170), .ZN(n10748) );
  INV_X1 U8095 ( .A(n14915), .ZN(n15086) );
  OR2_X1 U8096 ( .A1(n9819), .A2(n14127), .ZN(n7760) );
  OR2_X1 U8097 ( .A1(n9077), .A2(n7387), .ZN(n7383) );
  INV_X1 U8098 ( .A(n7388), .ZN(n7387) );
  AOI21_X1 U8099 ( .B1(n7388), .B2(n7386), .A(n7385), .ZN(n7384) );
  INV_X1 U8100 ( .A(n9081), .ZN(n7385) );
  INV_X1 U8101 ( .A(n9076), .ZN(n7386) );
  NOR2_X1 U8102 ( .A1(n9104), .A2(n7389), .ZN(n7388) );
  INV_X1 U8103 ( .A(n9079), .ZN(n7389) );
  XNOR2_X1 U8104 ( .A(n9077), .B(n9076), .ZN(n13789) );
  NOR2_X1 U8105 ( .A1(n7700), .A2(P1_IR_REG_27__SCAN_IN), .ZN(n7233) );
  INV_X1 U8106 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n7715) );
  NOR2_X1 U8107 ( .A1(n7700), .A2(n7695), .ZN(n6993) );
  XNOR2_X1 U8108 ( .A(n8191), .B(n8190), .ZN(n13802) );
  NAND2_X1 U8109 ( .A1(n6797), .A2(SI_14_), .ZN(n7991) );
  OR2_X1 U8110 ( .A1(n7939), .A2(P1_IR_REG_11__SCAN_IN), .ZN(n7956) );
  XNOR2_X1 U8111 ( .A(n7068), .B(n7937), .ZN(n10289) );
  NAND2_X1 U8112 ( .A1(n7917), .A2(n7916), .ZN(n7068) );
  AOI21_X1 U8113 ( .B1(n6933), .B2(n6931), .A(n6930), .ZN(n6929) );
  INV_X1 U8114 ( .A(n7899), .ZN(n6930) );
  INV_X1 U8115 ( .A(n7071), .ZN(n6931) );
  INV_X1 U8116 ( .A(n6933), .ZN(n6932) );
  AOI21_X1 U8117 ( .B1(n7861), .B2(n7073), .A(n7072), .ZN(n7071) );
  INV_X1 U8118 ( .A(n7878), .ZN(n7072) );
  INV_X1 U8119 ( .A(n7857), .ZN(n7073) );
  AOI21_X1 U8120 ( .B1(n6934), .B2(n7071), .A(n7881), .ZN(n6933) );
  NAND2_X2 U8121 ( .A1(n7362), .A2(n7361), .ZN(n7858) );
  AOI21_X1 U8122 ( .B1(n7363), .B2(n7824), .A(n7841), .ZN(n7361) );
  INV_X1 U8123 ( .A(n7364), .ZN(n7363) );
  OAI21_X1 U8124 ( .B1(n7821), .B2(n7824), .A(n7838), .ZN(n7364) );
  NAND2_X1 U8125 ( .A1(n7822), .A2(n7821), .ZN(n7826) );
  OAI21_X1 U8126 ( .B1(P3_ADDR_REG_14__SCAN_IN), .B2(n15010), .A(n7609), .ZN(
        n7664) );
  NAND2_X1 U8127 ( .A1(n9646), .A2(n9645), .ZN(n12372) );
  INV_X1 U8128 ( .A(n12941), .ZN(n12451) );
  AND4_X1 U8129 ( .A1(n9463), .A2(n9462), .A3(n9461), .A4(n9460), .ZN(n12599)
         );
  AND4_X1 U8130 ( .A1(n9325), .A2(n9324), .A3(n9323), .A4(n9322), .ZN(n11444)
         );
  AND4_X1 U8131 ( .A1(n9516), .A2(n9515), .A3(n9514), .A4(n9513), .ZN(n13017)
         );
  INV_X1 U8132 ( .A(n12982), .ZN(n13078) );
  NAND2_X1 U8133 ( .A1(n9575), .A2(n9574), .ZN(n12958) );
  AND4_X1 U8134 ( .A1(n9384), .A2(n9383), .A3(n9382), .A4(n9381), .ZN(n12113)
         );
  INV_X1 U8135 ( .A(n9689), .ZN(n12720) );
  AND2_X1 U8136 ( .A1(n11251), .A2(n9680), .ZN(n12859) );
  INV_X1 U8137 ( .A(n12954), .ZN(n12977) );
  INV_X1 U8138 ( .A(n12478), .ZN(n13030) );
  INV_X1 U8139 ( .A(n12599), .ZN(n13028) );
  INV_X1 U8140 ( .A(n12113), .ZN(n12416) );
  AOI22_X1 U8141 ( .A1(n10846), .A2(n10847), .B1(n10809), .B2(n10795), .ZN(
        n10894) );
  NAND2_X1 U8142 ( .A1(n11654), .A2(n11655), .ZN(n11895) );
  AOI21_X1 U8143 ( .B1(n11892), .B2(n11891), .A(n11890), .ZN(n11894) );
  NAND2_X1 U8144 ( .A1(n11894), .A2(n11893), .ZN(n11930) );
  XNOR2_X1 U8145 ( .A(n12781), .B(n6775), .ZN(n12760) );
  NOR2_X1 U8146 ( .A1(n12760), .A2(n12759), .ZN(n12782) );
  XNOR2_X1 U8147 ( .A(n6867), .B(n6866), .ZN(n12810) );
  AOI21_X1 U8148 ( .B1(n6976), .B2(n15426), .A(n6973), .ZN(n6972) );
  NAND2_X1 U8149 ( .A1(n12840), .A2(n6974), .ZN(n6973) );
  XNOR2_X1 U8150 ( .A(n12838), .B(n12837), .ZN(n6976) );
  NAND2_X1 U8151 ( .A1(n6970), .A2(n15429), .ZN(n6969) );
  XNOR2_X1 U8152 ( .A(n12846), .B(n6971), .ZN(n6970) );
  INV_X1 U8153 ( .A(n12845), .ZN(n6971) );
  OAI22_X1 U8154 ( .A1(n12844), .A2(n12843), .B1(n12842), .B2(n13006), .ZN(
        n12846) );
  AOI21_X1 U8155 ( .B1(n12664), .B2(n9615), .A(n6769), .ZN(n12854) );
  NAND2_X1 U8156 ( .A1(n7491), .A2(n6898), .ZN(n7490) );
  AND2_X1 U8157 ( .A1(n7492), .A2(n15493), .ZN(n6898) );
  AND2_X1 U8158 ( .A1(n9586), .A2(n9585), .ZN(n13126) );
  OR2_X1 U8159 ( .A1(n15491), .A2(n15486), .ZN(n13144) );
  AND2_X1 U8160 ( .A1(n7511), .A2(n7510), .ZN(n7509) );
  INV_X1 U8161 ( .A(P3_IR_REG_29__SCAN_IN), .ZN(n7510) );
  NAND2_X1 U8162 ( .A1(n7421), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9209) );
  NAND2_X1 U8163 ( .A1(n13174), .A2(n6675), .ZN(n14842) );
  INV_X1 U8164 ( .A(n14839), .ZN(n13175) );
  NAND2_X1 U8165 ( .A1(n8509), .A2(n8508), .ZN(n15370) );
  NAND2_X1 U8166 ( .A1(n11336), .A2(n11335), .ZN(n7517) );
  NAND2_X1 U8167 ( .A1(n7534), .A2(n11939), .ZN(n7533) );
  NAND2_X1 U8168 ( .A1(n7532), .A2(n11939), .ZN(n7531) );
  INV_X1 U8169 ( .A(n11770), .ZN(n7534) );
  NAND2_X1 U8170 ( .A1(n8599), .A2(n8598), .ZN(n14853) );
  NAND2_X1 U8171 ( .A1(n11951), .A2(n11950), .ZN(n13174) );
  OR3_X1 U8172 ( .A1(n10637), .A2(n10636), .A3(n15355), .ZN(n13349) );
  NAND2_X1 U8173 ( .A1(n9109), .A2(n9108), .ZN(n13445) );
  OR2_X1 U8174 ( .A1(n14760), .A2(n9107), .ZN(n9109) );
  NAND2_X1 U8175 ( .A1(n13617), .A2(n8846), .ZN(n13596) );
  NAND2_X1 U8176 ( .A1(n8495), .A2(n8494), .ZN(n11746) );
  NAND2_X1 U8177 ( .A1(n8810), .A2(n8809), .ZN(n15348) );
  INV_X1 U8178 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n10823) );
  OR2_X1 U8179 ( .A1(n10821), .A2(n14127), .ZN(n7981) );
  OAI21_X1 U8180 ( .B1(n6704), .B2(n7087), .A(n9905), .ZN(n7086) );
  NOR2_X1 U8181 ( .A1(n6833), .A2(n7718), .ZN(n7087) );
  NAND2_X1 U8182 ( .A1(n6944), .A2(n8061), .ZN(n14537) );
  INV_X1 U8183 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n14341) );
  INV_X1 U8184 ( .A(n14333), .ZN(n6814) );
  NAND2_X1 U8185 ( .A1(n14374), .A2(n14375), .ZN(n6985) );
  NAND2_X1 U8186 ( .A1(n7909), .A2(n7908), .ZN(n14029) );
  NAND2_X1 U8187 ( .A1(n7890), .A2(n7889), .ZN(n15156) );
  NAND2_X1 U8188 ( .A1(n7961), .A2(n7960), .ZN(n14043) );
  NAND2_X1 U8189 ( .A1(n13963), .A2(n13962), .ZN(n14711) );
  OR2_X1 U8190 ( .A1(n14760), .A2(n14127), .ZN(n14129) );
  OR2_X1 U8191 ( .A1(n14374), .A2(n15075), .ZN(n6986) );
  OR2_X1 U8192 ( .A1(n14626), .A2(n6924), .ZN(n6988) );
  MUX2_X1 U8193 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8086), .S(
        P1_IR_REG_19__SCAN_IN), .Z(n8090) );
  INV_X1 U8194 ( .A(n15510), .ZN(n7045) );
  OAI21_X1 U8195 ( .B1(n14966), .B2(n14967), .A(n6799), .ZN(n6798) );
  INV_X1 U8196 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n6799) );
  NAND2_X1 U8197 ( .A1(n14814), .A2(n7673), .ZN(n14781) );
  INV_X1 U8198 ( .A(n7053), .ZN(n7672) );
  NAND2_X1 U8199 ( .A1(n14781), .A2(n14780), .ZN(n14779) );
  OAI21_X1 U8200 ( .B1(n14781), .B2(n14780), .A(n7067), .ZN(n7066) );
  INV_X1 U8201 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n7067) );
  INV_X1 U8202 ( .A(n8936), .ZN(n6840) );
  NAND2_X1 U8203 ( .A1(n7146), .A2(n14008), .ZN(n7145) );
  NAND2_X1 U8204 ( .A1(n7141), .A2(n14019), .ZN(n7140) );
  NAND2_X1 U8205 ( .A1(n7552), .A2(n6678), .ZN(n8960) );
  INV_X1 U8206 ( .A(n8953), .ZN(n7553) );
  NAND2_X1 U8207 ( .A1(n7151), .A2(n14030), .ZN(n7150) );
  NAND2_X1 U8208 ( .A1(n8969), .A2(n6656), .ZN(n8974) );
  NOR2_X1 U8209 ( .A1(n6857), .A2(n6856), .ZN(n6855) );
  NOR2_X1 U8210 ( .A1(n7560), .A2(n8973), .ZN(n6856) );
  NOR2_X1 U8211 ( .A1(n6658), .A2(n6858), .ZN(n6857) );
  INV_X1 U8212 ( .A(n8977), .ZN(n7560) );
  NAND2_X1 U8213 ( .A1(n7136), .A2(n14041), .ZN(n7135) );
  NAND2_X1 U8214 ( .A1(n8992), .A2(n6740), .ZN(n6842) );
  NAND2_X1 U8215 ( .A1(n6659), .A2(n8996), .ZN(n7556) );
  AOI21_X1 U8216 ( .B1(n9003), .B2(n9013), .A(n9002), .ZN(n9016) );
  NAND2_X1 U8217 ( .A1(n7127), .A2(n7129), .ZN(n7126) );
  NAND2_X1 U8218 ( .A1(n6844), .A2(n6843), .ZN(n9034) );
  AOI21_X1 U8219 ( .B1(n6845), .B2(n6847), .A(n6708), .ZN(n6843) );
  NOR2_X1 U8220 ( .A1(n9022), .A2(n6669), .ZN(n6847) );
  NAND2_X1 U8221 ( .A1(n6940), .A2(n14096), .ZN(n6939) );
  NAND2_X1 U8222 ( .A1(n14097), .A2(n14098), .ZN(n6940) );
  AOI21_X1 U8223 ( .B1(n6635), .B2(n6851), .A(n6710), .ZN(n6849) );
  NOR2_X1 U8224 ( .A1(n6660), .A2(n6852), .ZN(n6851) );
  NOR2_X1 U8225 ( .A1(n7545), .A2(n6670), .ZN(n7544) );
  AOI21_X1 U8226 ( .B1(n7541), .B2(n7539), .A(n7538), .ZN(n7537) );
  INV_X1 U8227 ( .A(n7543), .ZN(n7539) );
  INV_X1 U8228 ( .A(n9062), .ZN(n7538) );
  NAND2_X1 U8229 ( .A1(n14103), .A2(n14104), .ZN(n14102) );
  INV_X1 U8230 ( .A(n9228), .ZN(n6896) );
  NAND2_X1 U8231 ( .A1(n8890), .A2(n9168), .ZN(n8910) );
  INV_X1 U8232 ( .A(P2_RD_REG_SCAN_IN), .ZN(n7358) );
  NAND2_X1 U8233 ( .A1(n12914), .A2(n12517), .ZN(n7420) );
  NOR2_X1 U8234 ( .A1(n7419), .A2(n7020), .ZN(n7019) );
  INV_X1 U8235 ( .A(n7022), .ZN(n7020) );
  NAND2_X1 U8236 ( .A1(n7420), .A2(n12902), .ZN(n7419) );
  INV_X1 U8237 ( .A(n12603), .ZN(n7417) );
  NAND2_X1 U8238 ( .A1(n12739), .A2(n10785), .ZN(n12541) );
  INV_X1 U8239 ( .A(P3_IR_REG_9__SCAN_IN), .ZN(n9182) );
  INV_X1 U8240 ( .A(n9387), .ZN(n7183) );
  INV_X1 U8241 ( .A(n9372), .ZN(n6897) );
  NAND2_X1 U8242 ( .A1(n7549), .A2(n9095), .ZN(n7548) );
  INV_X1 U8243 ( .A(n9100), .ZN(n7549) );
  INV_X1 U8244 ( .A(n9071), .ZN(n6838) );
  INV_X1 U8245 ( .A(n9095), .ZN(n7550) );
  INV_X1 U8246 ( .A(n9165), .ZN(n9141) );
  INV_X1 U8247 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n8419) );
  NAND2_X1 U8248 ( .A1(n14116), .A2(n14113), .ZN(n6963) );
  AOI21_X1 U8249 ( .B1(n14715), .B2(n14091), .A(n14133), .ZN(n14149) );
  NAND2_X1 U8250 ( .A1(n8155), .A2(n8674), .ZN(n7367) );
  NOR2_X1 U8251 ( .A1(n7394), .A2(n7393), .ZN(n7392) );
  INV_X1 U8252 ( .A(n8098), .ZN(n7393) );
  INV_X1 U8253 ( .A(n8069), .ZN(n8074) );
  INV_X1 U8254 ( .A(n7969), .ZN(n6947) );
  NAND2_X1 U8255 ( .A1(n6808), .A2(n6807), .ZN(n7719) );
  NAND2_X1 U8256 ( .A1(n6834), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n6807) );
  OR2_X1 U8257 ( .A1(n6834), .A2(n9820), .ZN(n6808) );
  OR2_X1 U8258 ( .A1(n12657), .A2(n12656), .ZN(n6795) );
  AND2_X1 U8259 ( .A1(n12695), .A2(n12694), .ZN(n12697) );
  NAND2_X1 U8260 ( .A1(n6872), .A2(n6871), .ZN(n6870) );
  NAND2_X1 U8261 ( .A1(n10807), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n6871) );
  INV_X1 U8262 ( .A(n15393), .ZN(n6872) );
  NAND2_X1 U8263 ( .A1(n11078), .A2(n6860), .ZN(n11648) );
  OR2_X1 U8264 ( .A1(n11080), .A2(n11079), .ZN(n6860) );
  NAND2_X1 U8265 ( .A1(n15423), .A2(n6980), .ZN(n6979) );
  NAND2_X1 U8266 ( .A1(n11661), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n6980) );
  NAND2_X1 U8267 ( .A1(n11895), .A2(n6859), .ZN(n11917) );
  OR2_X1 U8268 ( .A1(n11901), .A2(n11896), .ZN(n6859) );
  AND2_X1 U8269 ( .A1(n7018), .A2(n6663), .ZN(n6901) );
  NAND2_X1 U8270 ( .A1(n7506), .A2(n9639), .ZN(n7505) );
  NAND2_X1 U8271 ( .A1(n12902), .A2(n9624), .ZN(n7506) );
  AND2_X1 U8272 ( .A1(n6666), .A2(n9569), .ZN(n7488) );
  AOI21_X1 U8273 ( .B1(n12937), .B2(n7023), .A(n12514), .ZN(n7022) );
  INV_X1 U8274 ( .A(n12522), .ZN(n7023) );
  OR2_X1 U8275 ( .A1(n9587), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n9603) );
  NAND2_X1 U8276 ( .A1(n9577), .A2(n9576), .ZN(n9587) );
  NAND2_X1 U8277 ( .A1(n9707), .A2(n7006), .ZN(n7005) );
  INV_X1 U8278 ( .A(n9706), .ZN(n7006) );
  AND2_X1 U8279 ( .A1(n12983), .A2(n7498), .ZN(n7497) );
  NAND2_X1 U8280 ( .A1(n7499), .A2(n9540), .ZN(n7498) );
  INV_X1 U8281 ( .A(n7501), .ZN(n7499) );
  AND2_X1 U8282 ( .A1(n12993), .A2(n12615), .ZN(n12690) );
  NAND2_X1 U8283 ( .A1(n7013), .A2(n7015), .ZN(n7012) );
  INV_X1 U8284 ( .A(P3_REG3_REG_11__SCAN_IN), .ZN(n11708) );
  AOI21_X1 U8285 ( .B1(n15446), .B2(n9698), .A(n7565), .ZN(n10780) );
  AND2_X1 U8286 ( .A1(n9191), .A2(n9344), .ZN(n9192) );
  INV_X1 U8287 ( .A(P3_IR_REG_25__SCAN_IN), .ZN(n9193) );
  AOI21_X1 U8288 ( .B1(n7197), .B2(n7194), .A(n6771), .ZN(n7193) );
  NAND2_X1 U8289 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(n7176), .ZN(n7175) );
  INV_X1 U8290 ( .A(n9446), .ZN(n7173) );
  NOR2_X1 U8291 ( .A1(n7173), .A2(n7174), .ZN(n7171) );
  NAND2_X1 U8292 ( .A1(n6650), .A2(n9225), .ZN(n7187) );
  INV_X1 U8293 ( .A(P3_IR_REG_4__SCAN_IN), .ZN(n9190) );
  INV_X1 U8294 ( .A(P3_IR_REG_3__SCAN_IN), .ZN(n9189) );
  AND2_X2 U8295 ( .A1(n6864), .A2(n6865), .ZN(n9266) );
  INV_X1 U8296 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n6864) );
  INV_X1 U8297 ( .A(P3_IR_REG_1__SCAN_IN), .ZN(n6865) );
  NOR2_X1 U8298 ( .A1(n8639), .A2(n10119), .ZN(n8652) );
  INV_X1 U8299 ( .A(n13288), .ZN(n7083) );
  NAND2_X1 U8300 ( .A1(n13267), .A2(n7074), .ZN(n13203) );
  NAND2_X1 U8301 ( .A1(n13199), .A2(n7075), .ZN(n7074) );
  INV_X1 U8302 ( .A(n13200), .ZN(n7075) );
  INV_X1 U8303 ( .A(n9086), .ZN(n7379) );
  INV_X1 U8304 ( .A(n9090), .ZN(n8690) );
  NOR2_X1 U8305 ( .A1(n13688), .A2(n6882), .ZN(n6881) );
  NOR2_X1 U8306 ( .A1(n7437), .A2(n7435), .ZN(n7434) );
  INV_X1 U8307 ( .A(n8856), .ZN(n7435) );
  NOR2_X1 U8308 ( .A1(n13524), .A2(n6886), .ZN(n6885) );
  INV_X1 U8309 ( .A(n6887), .ZN(n6886) );
  NOR2_X1 U8310 ( .A1(n13716), .A2(n13557), .ZN(n6887) );
  INV_X1 U8311 ( .A(n8589), .ZN(n7264) );
  NOR2_X1 U8312 ( .A1(n13630), .A2(n6878), .ZN(n6877) );
  INV_X1 U8313 ( .A(n6879), .ZN(n6878) );
  NOR2_X1 U8314 ( .A1(n14853), .A2(n13642), .ZN(n6879) );
  NAND2_X1 U8315 ( .A1(n8837), .A2(n11756), .ZN(n7448) );
  NOR2_X1 U8316 ( .A1(n11811), .A2(n7450), .ZN(n7451) );
  INV_X1 U8317 ( .A(n11589), .ZN(n7269) );
  INV_X1 U8318 ( .A(n10648), .ZN(n8899) );
  NAND2_X1 U8319 ( .A1(n13479), .A2(n6636), .ZN(n13452) );
  INV_X1 U8320 ( .A(n9796), .ZN(n9794) );
  NAND2_X1 U8321 ( .A1(n9794), .A2(n9793), .ZN(n9792) );
  CLKBUF_X1 U8322 ( .A(n8477), .Z(n8478) );
  NAND2_X1 U8323 ( .A1(n13969), .A2(n6629), .ZN(n7329) );
  NOR2_X1 U8324 ( .A1(n11989), .A2(n7340), .ZN(n7339) );
  INV_X1 U8325 ( .A(n11548), .ZN(n7340) );
  INV_X1 U8326 ( .A(n10428), .ZN(n11299) );
  OR2_X1 U8327 ( .A1(n14155), .A2(n8305), .ZN(n13949) );
  NOR2_X1 U8328 ( .A1(n15044), .A2(n14328), .ZN(n14330) );
  INV_X1 U8329 ( .A(n14373), .ZN(n7117) );
  OR2_X1 U8330 ( .A1(n14419), .A2(n12285), .ZN(n7123) );
  NAND2_X1 U8331 ( .A1(n14425), .A2(n7120), .ZN(n7124) );
  AND2_X1 U8332 ( .A1(n14193), .A2(n7123), .ZN(n7119) );
  NAND2_X1 U8333 ( .A1(n6913), .A2(n6912), .ZN(n6911) );
  INV_X1 U8334 ( .A(n6914), .ZN(n6913) );
  NOR2_X1 U8335 ( .A1(n6917), .A2(n14705), .ZN(n6916) );
  INV_X1 U8336 ( .A(n6918), .ZN(n6917) );
  INV_X1 U8337 ( .A(n8265), .ZN(n7094) );
  NOR2_X1 U8338 ( .A1(n10745), .A2(n7095), .ZN(n7001) );
  OR2_X1 U8339 ( .A1(n6617), .A2(n7741), .ZN(n7742) );
  NOR2_X1 U8340 ( .A1(n14610), .A2(n15156), .ZN(n14613) );
  NAND2_X1 U8341 ( .A1(n7739), .A2(n7228), .ZN(n11051) );
  AND2_X1 U8342 ( .A1(n8098), .A2(n8079), .ZN(n8080) );
  OAI21_X1 U8343 ( .B1(n7088), .B2(n6811), .A(n6810), .ZN(n7802) );
  NAND2_X1 U8344 ( .A1(n7088), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n6810) );
  OAI21_X1 U8345 ( .B1(n7076), .B2(SI_4_), .A(n7800), .ZN(n7782) );
  NAND2_X1 U8346 ( .A1(n7719), .A2(SI_1_), .ZN(n7746) );
  OAI21_X1 U8347 ( .B1(SI_1_), .B2(n7719), .A(n7746), .ZN(n7723) );
  NAND2_X1 U8348 ( .A1(n8192), .A2(n9214), .ZN(n6831) );
  XNOR2_X1 U8349 ( .A(n10934), .B(P1_ADDR_REG_1__SCAN_IN), .ZN(n7631) );
  INV_X1 U8350 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10158) );
  NOR2_X1 U8351 ( .A1(n7583), .A2(n7582), .ZN(n7585) );
  INV_X1 U8352 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n7581) );
  INV_X1 U8353 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n7584) );
  NAND2_X1 U8355 ( .A1(n7310), .A2(n7309), .ZN(n7308) );
  INV_X1 U8356 ( .A(n12484), .ZN(n7309) );
  AND2_X1 U8357 ( .A1(n11870), .A2(n11868), .ZN(n7297) );
  OAI21_X1 U8358 ( .B1(n7305), .B2(n7301), .A(n6707), .ZN(n7300) );
  INV_X1 U8359 ( .A(n12390), .ZN(n7301) );
  INV_X1 U8360 ( .A(n7308), .ZN(n7303) );
  AND2_X1 U8361 ( .A1(n9562), .A2(n9561), .ZN(n9577) );
  INV_X1 U8362 ( .A(n12361), .ZN(n12448) );
  AOI21_X1 U8363 ( .B1(n7283), .B2(n7285), .A(n6741), .ZN(n7281) );
  NAND2_X1 U8364 ( .A1(n12032), .A2(n12031), .ZN(n12411) );
  XNOR2_X1 U8365 ( .A(n12392), .B(n11370), .ZN(n10681) );
  XNOR2_X1 U8366 ( .A(n12360), .B(n10953), .ZN(n10688) );
  INV_X1 U8367 ( .A(n12703), .ZN(n7162) );
  NAND2_X1 U8368 ( .A1(n12713), .A2(n7028), .ZN(n7027) );
  AND2_X1 U8369 ( .A1(n6720), .A2(n7025), .ZN(n7024) );
  NAND2_X1 U8370 ( .A1(n12713), .A2(n6696), .ZN(n7025) );
  AND2_X1 U8371 ( .A1(n9234), .A2(n9233), .ZN(n9236) );
  XNOR2_X1 U8372 ( .A(n10799), .B(n10798), .ZN(n10796) );
  OAI22_X1 U8373 ( .A1(n10796), .A2(n10797), .B1(n10799), .B2(n10798), .ZN(
        n15397) );
  NAND2_X1 U8374 ( .A1(n15397), .A2(n15398), .ZN(n15396) );
  NOR2_X1 U8375 ( .A1(n10790), .A2(n10789), .ZN(n15405) );
  NOR2_X1 U8376 ( .A1(n15405), .A2(n15404), .ZN(n15403) );
  NAND2_X1 U8377 ( .A1(n10856), .A2(n10855), .ZN(n10854) );
  OAI22_X1 U8378 ( .A1(n10867), .A2(n10067), .B1(n6869), .B2(n10808), .ZN(
        n10853) );
  INV_X1 U8379 ( .A(n6870), .ZN(n6869) );
  NAND2_X1 U8380 ( .A1(n10854), .A2(n6967), .ZN(n10895) );
  OR2_X1 U8381 ( .A1(n10809), .A2(n9319), .ZN(n6967) );
  NAND2_X1 U8382 ( .A1(n10902), .A2(n10903), .ZN(n10904) );
  XNOR2_X1 U8383 ( .A(n11648), .B(n11659), .ZN(n11081) );
  INV_X1 U8384 ( .A(n6981), .ZN(n11660) );
  XNOR2_X1 U8385 ( .A(n6979), .B(n11713), .ZN(n11709) );
  OAI22_X1 U8386 ( .A1(n11709), .A2(n11662), .B1(n11675), .B2(n6978), .ZN(
        n11665) );
  INV_X1 U8387 ( .A(n6979), .ZN(n6978) );
  XNOR2_X1 U8388 ( .A(n11911), .B(n11899), .ZN(n11902) );
  XNOR2_X1 U8389 ( .A(n11917), .B(n11899), .ZN(n11897) );
  NAND2_X1 U8390 ( .A1(n11900), .A2(n6977), .ZN(n11911) );
  OR2_X1 U8391 ( .A1(n11901), .A2(n11663), .ZN(n6977) );
  NAND2_X1 U8392 ( .A1(n11902), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n11912) );
  NAND2_X1 U8393 ( .A1(n12744), .A2(n6861), .ZN(n12764) );
  OR2_X1 U8394 ( .A1(n12746), .A2(n12745), .ZN(n6861) );
  OAI21_X1 U8395 ( .B1(n12816), .B2(n13090), .A(n12819), .ZN(n12836) );
  AOI21_X1 U8396 ( .B1(n15417), .B2(n12847), .A(n6975), .ZN(n6974) );
  INV_X1 U8397 ( .A(n12839), .ZN(n6975) );
  AND2_X1 U8398 ( .A1(n12706), .A2(n12660), .ZN(n12695) );
  NAND2_X1 U8399 ( .A1(n12903), .A2(n9624), .ZN(n12887) );
  NAND2_X1 U8400 ( .A1(n12517), .A2(n12515), .ZN(n12914) );
  INV_X1 U8401 ( .A(n12914), .ZN(n12918) );
  NAND2_X1 U8402 ( .A1(n7021), .A2(n7022), .ZN(n12916) );
  OR2_X1 U8403 ( .A1(n9708), .A2(n9709), .ZN(n7021) );
  AND2_X1 U8404 ( .A1(n12522), .A2(n12521), .ZN(n12956) );
  AND4_X1 U8405 ( .A1(n9551), .A2(n9550), .A3(n9549), .A4(n9548), .ZN(n12966)
         );
  OR2_X1 U8406 ( .A1(n9533), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n9546) );
  INV_X1 U8407 ( .A(SI_18_), .ZN(n9506) );
  AOI21_X1 U8408 ( .B1(n6633), .B2(n7465), .A(n6692), .ZN(n7461) );
  INV_X1 U8409 ( .A(n6649), .ZN(n7465) );
  INV_X1 U8410 ( .A(n13013), .ZN(n13020) );
  AOI21_X1 U8411 ( .B1(n7036), .B2(n7039), .A(n7033), .ZN(n7032) );
  INV_X1 U8412 ( .A(n7040), .ZN(n7039) );
  NOR2_X1 U8413 ( .A1(n9475), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n9483) );
  AOI21_X1 U8414 ( .B1(n7480), .B2(n7484), .A(n6746), .ZN(n7478) );
  AND4_X1 U8415 ( .A1(n9371), .A2(n9370), .A3(n9369), .A4(n9368), .ZN(n12006)
         );
  OAI21_X1 U8416 ( .B1(n9317), .B2(n7495), .A(n7494), .ZN(n11405) );
  AOI21_X1 U8417 ( .B1(n7496), .B2(n12672), .A(n6638), .ZN(n7494) );
  INV_X1 U8418 ( .A(n7496), .ZN(n7495) );
  OR2_X1 U8419 ( .A1(n9320), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n9333) );
  INV_X1 U8420 ( .A(n10953), .ZN(n15458) );
  NAND2_X1 U8421 ( .A1(n9716), .A2(n9764), .ZN(n15454) );
  CLKBUF_X1 U8422 ( .A(n9253), .Z(n10678) );
  INV_X1 U8423 ( .A(n12854), .ZN(n14818) );
  NAND2_X1 U8424 ( .A1(n13153), .A2(n9615), .ZN(n7188) );
  AOI21_X1 U8425 ( .B1(n12890), .B2(n12641), .A(n6904), .ZN(n12875) );
  AND3_X1 U8426 ( .A1(n9295), .A2(n9294), .A3(n9293), .ZN(n15480) );
  NOR2_X1 U8427 ( .A1(P3_IR_REG_28__SCAN_IN), .A2(P3_IR_REG_27__SCAN_IN), .ZN(
        n7511) );
  AND2_X1 U8428 ( .A1(n14767), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n7159) );
  XNOR2_X1 U8429 ( .A(n9751), .B(n9181), .ZN(n10670) );
  XNOR2_X1 U8430 ( .A(n9688), .B(P3_IR_REG_20__SCAN_IN), .ZN(n9765) );
  NAND2_X1 U8431 ( .A1(n9528), .A2(n9527), .ZN(n9687) );
  INV_X1 U8432 ( .A(P3_IR_REG_19__SCAN_IN), .ZN(n9527) );
  NOR2_X2 U8433 ( .A1(n9523), .A2(n7278), .ZN(n9528) );
  INV_X1 U8434 ( .A(n9524), .ZN(n7278) );
  NAND2_X1 U8435 ( .A1(n9490), .A2(n9489), .ZN(n9492) );
  NOR2_X2 U8436 ( .A1(n9453), .A2(n9452), .ZN(n9749) );
  INV_X1 U8437 ( .A(P3_IR_REG_15__SCAN_IN), .ZN(n9455) );
  INV_X1 U8438 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n9407) );
  OR2_X1 U8439 ( .A1(n9453), .A2(P3_IR_REG_9__SCAN_IN), .ZN(n9388) );
  XNOR2_X1 U8440 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(P2_DATAO_REG_9__SCAN_IN), 
        .ZN(n9372) );
  NAND2_X1 U8441 ( .A1(n9229), .A2(n9228), .ZN(n9373) );
  XNOR2_X1 U8442 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .ZN(n9359) );
  INV_X1 U8443 ( .A(P3_IR_REG_7__SCAN_IN), .ZN(n9344) );
  XNOR2_X1 U8444 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .ZN(n9304) );
  XNOR2_X1 U8445 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .ZN(n9288) );
  INV_X1 U8446 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n6891) );
  OR2_X1 U8447 ( .A1(n8566), .A2(n8565), .ZN(n8581) );
  INV_X1 U8448 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n10119) );
  INV_X1 U8449 ( .A(n13223), .ZN(n7523) );
  INV_X1 U8450 ( .A(n7535), .ZN(n7532) );
  NOR2_X1 U8451 ( .A1(n8581), .A2(n11503), .ZN(n8600) );
  AND2_X1 U8452 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n8445) );
  NAND2_X1 U8453 ( .A1(n7083), .A2(n7082), .ZN(n7081) );
  INV_X1 U8454 ( .A(n13287), .ZN(n7082) );
  INV_X1 U8455 ( .A(n8698), .ZN(n8699) );
  NAND2_X1 U8456 ( .A1(P2_REG3_REG_24__SCAN_IN), .A2(n8699), .ZN(n8719) );
  INV_X1 U8457 ( .A(n10843), .ZN(n6873) );
  NAND2_X1 U8458 ( .A1(n6830), .A2(n7528), .ZN(n7530) );
  AND2_X1 U8459 ( .A1(n8540), .A2(n8539), .ZN(n8552) );
  NAND2_X1 U8460 ( .A1(n8552), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n8566) );
  OR2_X1 U8461 ( .A1(n11771), .A2(n11770), .ZN(n7536) );
  OR2_X1 U8462 ( .A1(n10291), .A2(n10305), .ZN(n13301) );
  AND2_X1 U8463 ( .A1(n8445), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n8456) );
  OAI211_X1 U8464 ( .C1(n7381), .C2(n13436), .A(n7378), .B(n7376), .ZN(n9165)
         );
  NAND2_X1 U8465 ( .A1(n7380), .A2(n7379), .ZN(n7378) );
  NAND2_X1 U8466 ( .A1(n7381), .A2(n7377), .ZN(n7376) );
  NOR2_X1 U8467 ( .A1(n7380), .A2(n7379), .ZN(n7377) );
  AOI21_X1 U8468 ( .B1(n6835), .B2(n9132), .A(n9131), .ZN(n9169) );
  NAND2_X1 U8469 ( .A1(n6836), .A2(n9123), .ZN(n6835) );
  OR2_X1 U8470 ( .A1(n10291), .A2(n8867), .ZN(n13303) );
  AND2_X1 U8471 ( .A1(n15309), .A2(n15308), .ZN(n15310) );
  NAND2_X1 U8472 ( .A1(n8596), .A2(n8608), .ZN(n8610) );
  NAND2_X1 U8473 ( .A1(n13479), .A2(n8876), .ZN(n13480) );
  NAND3_X1 U8474 ( .A1(n7271), .A2(n6884), .A3(n6885), .ZN(n13514) );
  NOR2_X1 U8475 ( .A1(n13514), .A2(n13698), .ZN(n13479) );
  INV_X1 U8476 ( .A(n13301), .ZN(n13336) );
  NAND2_X1 U8477 ( .A1(n7271), .A2(n6885), .ZN(n13522) );
  NAND2_X1 U8478 ( .A1(n7271), .A2(n7270), .ZN(n13555) );
  AOI21_X1 U8479 ( .B1(n7444), .B2(n7440), .A(n6690), .ZN(n7439) );
  AOI21_X1 U8480 ( .B1(n7252), .B2(n13628), .A(n6688), .ZN(n7250) );
  INV_X1 U8481 ( .A(n7252), .ZN(n7251) );
  AOI21_X1 U8482 ( .B1(n7454), .B2(n13620), .A(n6691), .ZN(n7452) );
  AND2_X1 U8483 ( .A1(n7274), .A2(n6875), .ZN(n13606) );
  NOR2_X1 U8484 ( .A1(n13609), .A2(n6876), .ZN(n6875) );
  INV_X1 U8485 ( .A(n6877), .ZN(n6876) );
  OR2_X1 U8486 ( .A1(n13619), .A2(n13620), .ZN(n13617) );
  NAND2_X1 U8487 ( .A1(n7274), .A2(n6877), .ZN(n13632) );
  NAND2_X1 U8488 ( .A1(n7274), .A2(n7273), .ZN(n12162) );
  INV_X1 U8489 ( .A(n7274), .ZN(n12139) );
  NAND2_X1 U8490 ( .A1(n8840), .A2(n8839), .ZN(n12012) );
  OAI21_X1 U8491 ( .B1(n11810), .B2(n8548), .A(n8547), .ZN(n11968) );
  NAND2_X1 U8492 ( .A1(n7269), .A2(n6631), .ZN(n11820) );
  AND2_X1 U8493 ( .A1(n7269), .A2(n6643), .ZN(n11969) );
  NAND2_X1 U8494 ( .A1(n11750), .A2(n8837), .ZN(n11812) );
  NAND2_X1 U8495 ( .A1(n11750), .A2(n7451), .ZN(n11814) );
  NAND2_X1 U8496 ( .A1(n8835), .A2(n8834), .ZN(n11749) );
  OR2_X1 U8497 ( .A1(n11749), .A2(n11756), .ZN(n11750) );
  NOR2_X1 U8498 ( .A1(n8511), .A2(n8510), .ZN(n8540) );
  NAND2_X1 U8499 ( .A1(n7269), .A2(n7268), .ZN(n11759) );
  NAND2_X1 U8500 ( .A1(n8505), .A2(n8504), .ZN(n11582) );
  NOR2_X1 U8501 ( .A1(n11462), .A2(n15364), .ZN(n11564) );
  NAND2_X1 U8502 ( .A1(n11564), .A2(n11743), .ZN(n11589) );
  NOR2_X1 U8503 ( .A1(n10960), .A2(n10965), .ZN(n11115) );
  NAND2_X1 U8504 ( .A1(n6874), .A2(n11130), .ZN(n10960) );
  INV_X1 U8505 ( .A(n10768), .ZN(n6874) );
  NAND2_X1 U8506 ( .A1(n13650), .A2(n10736), .ZN(n10768) );
  NAND2_X1 U8507 ( .A1(n10648), .A2(n10639), .ZN(n13652) );
  AND2_X1 U8508 ( .A1(n12326), .A2(n13429), .ZN(n10916) );
  INV_X1 U8509 ( .A(n8876), .ZN(n6882) );
  AND2_X1 U8510 ( .A1(n8816), .A2(n15362), .ZN(n13734) );
  NOR2_X1 U8511 ( .A1(n9819), .A2(n8438), .ZN(n8409) );
  INV_X1 U8512 ( .A(n8438), .ZN(n6800) );
  NOR2_X1 U8513 ( .A1(n10544), .A2(n8808), .ZN(n10605) );
  XNOR2_X1 U8514 ( .A(n8796), .B(n8795), .ZN(n10630) );
  INV_X1 U8515 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n8784) );
  OR2_X1 U8516 ( .A1(n8433), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n8440) );
  INV_X1 U8517 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n8441) );
  CLKBUF_X1 U8518 ( .A(n8382), .Z(n8403) );
  INV_X1 U8519 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n9214) );
  AND2_X1 U8520 ( .A1(n12204), .A2(n7352), .ZN(n7351) );
  NAND2_X1 U8521 ( .A1(n7353), .A2(n12194), .ZN(n7352) );
  AND2_X1 U8522 ( .A1(n14888), .A2(n14889), .ZN(n12204) );
  NAND2_X1 U8523 ( .A1(n12053), .A2(n12054), .ZN(n7324) );
  NOR2_X1 U8524 ( .A1(n11172), .A2(n6817), .ZN(n13826) );
  NOR2_X1 U8525 ( .A1(n11170), .A2(n11171), .ZN(n6817) );
  AND2_X1 U8526 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(n8225), .ZN(n8226) );
  INV_X1 U8527 ( .A(n11721), .ZN(n7343) );
  INV_X1 U8528 ( .A(n8162), .ZN(n8163) );
  NAND2_X1 U8529 ( .A1(n8163), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n8182) );
  NOR2_X1 U8530 ( .A1(n8102), .A2(n13896), .ZN(n8120) );
  NOR2_X1 U8531 ( .A1(n6827), .A2(n12194), .ZN(n13900) );
  AND2_X1 U8532 ( .A1(n8120), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n8135) );
  NAND2_X1 U8533 ( .A1(n13910), .A2(n13911), .ZN(n13909) );
  AND2_X1 U8534 ( .A1(n14901), .A2(n14902), .ZN(n7323) );
  NOR2_X1 U8535 ( .A1(n10183), .A2(n8182), .ZN(n8197) );
  NOR2_X1 U8536 ( .A1(n10222), .A2(n8195), .ZN(n8225) );
  OR2_X1 U8537 ( .A1(n7983), .A2(n7982), .ZN(n8004) );
  AND2_X1 U8538 ( .A1(n14142), .A2(n6959), .ZN(n6958) );
  NAND2_X1 U8539 ( .A1(n14126), .A2(n6960), .ZN(n6959) );
  INV_X1 U8540 ( .A(n14140), .ZN(n6960) );
  AND4_X1 U8541 ( .A1(n8249), .A2(n8248), .A3(n8247), .A4(n8246), .ZN(n14138)
         );
  AND3_X1 U8542 ( .A1(n8046), .A2(n8045), .A3(n8044), .ZN(n14063) );
  OR2_X1 U8543 ( .A1(n6617), .A2(n6803), .ZN(n7775) );
  AOI21_X1 U8544 ( .B1(P1_REG1_REG_2__SCAN_IN), .B2(n10449), .A(n9915), .ZN(
        n14247) );
  AOI21_X1 U8545 ( .B1(n9917), .B2(P1_REG1_REG_4__SCAN_IN), .A(n10457), .ZN(
        n14261) );
  AOI21_X1 U8546 ( .B1(P1_REG1_REG_6__SCAN_IN), .B2(n10376), .A(n10375), .ZN(
        n10379) );
  AOI21_X1 U8547 ( .B1(n10989), .B2(P1_REG1_REG_7__SCAN_IN), .A(n10988), .ZN(
        n14275) );
  AOI21_X1 U8548 ( .B1(P1_REG1_REG_10__SCAN_IN), .B2(n11104), .A(n11099), .ZN(
        n11102) );
  NOR2_X1 U8549 ( .A1(n14372), .A2(n7213), .ZN(n7212) );
  INV_X1 U8550 ( .A(n8214), .ZN(n7213) );
  NAND2_X1 U8551 ( .A1(n7124), .A2(n7119), .ZN(n7567) );
  OR2_X1 U8552 ( .A1(n7231), .A2(n8169), .ZN(n7229) );
  NOR2_X1 U8553 ( .A1(n14724), .A2(n14728), .ZN(n6922) );
  AOI21_X1 U8554 ( .B1(n7097), .B2(n7099), .A(n6694), .ZN(n7096) );
  NAND2_X1 U8555 ( .A1(n7092), .A2(n7091), .ZN(n14450) );
  INV_X1 U8556 ( .A(n7092), .ZN(n14465) );
  NAND2_X1 U8557 ( .A1(n6910), .A2(n6909), .ZN(n14476) );
  NOR2_X1 U8558 ( .A1(n14481), .A2(n6911), .ZN(n6909) );
  OR2_X1 U8559 ( .A1(n8094), .A2(n13839), .ZN(n8102) );
  NOR2_X1 U8560 ( .A1(n14536), .A2(n14528), .ZN(n14527) );
  OR2_X1 U8561 ( .A1(n8063), .A2(n8062), .ZN(n8094) );
  OR2_X1 U8562 ( .A1(n6919), .A2(n14698), .ZN(n14555) );
  OR2_X1 U8563 ( .A1(n14565), .A2(n14577), .ZN(n7115) );
  NOR2_X1 U8564 ( .A1(n8004), .A2(n8003), .ZN(n8022) );
  NAND2_X1 U8565 ( .A1(n11858), .A2(n6918), .ZN(n14587) );
  AND4_X1 U8566 ( .A1(n7989), .A2(n7988), .A3(n7987), .A4(n7986), .ZN(n13904)
         );
  AOI21_X1 U8567 ( .B1(n7216), .B2(n7217), .A(n6685), .ZN(n7215) );
  NAND2_X1 U8568 ( .A1(n7085), .A2(n7084), .ZN(n11859) );
  INV_X1 U8569 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n7944) );
  NOR2_X1 U8570 ( .A1(n7945), .A2(n7944), .ZN(n7962) );
  AOI21_X1 U8571 ( .B1(n7108), .B2(n14607), .A(n6687), .ZN(n7107) );
  AND2_X1 U8572 ( .A1(n7090), .A2(n11040), .ZN(n15085) );
  AND3_X1 U8573 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n7831) );
  INV_X1 U8574 ( .A(n14175), .ZN(n15073) );
  NAND2_X1 U8575 ( .A1(n7200), .A2(n11192), .ZN(n7199) );
  NAND2_X1 U8576 ( .A1(n11040), .A2(n15123), .ZN(n15084) );
  NAND2_X1 U8577 ( .A1(n7093), .A2(n6998), .ZN(n11043) );
  NAND2_X1 U8578 ( .A1(n10749), .A2(n7001), .ZN(n6998) );
  INV_X1 U8579 ( .A(n14601), .ZN(n14921) );
  NAND2_X1 U8580 ( .A1(n7227), .A2(n7739), .ZN(n9775) );
  NAND2_X1 U8581 ( .A1(n8279), .A2(n8278), .ZN(n14930) );
  AND2_X1 U8582 ( .A1(n11040), .A2(n11557), .ZN(n7089) );
  NAND2_X1 U8583 ( .A1(n8261), .A2(n12288), .ZN(n15129) );
  NAND2_X1 U8584 ( .A1(n14928), .A2(n8346), .ZN(n15155) );
  OAI21_X1 U8585 ( .B1(n8191), .B2(n7398), .A(n7395), .ZN(n8220) );
  AOI21_X1 U8586 ( .B1(n7397), .B2(n7396), .A(n6647), .ZN(n7395) );
  INV_X1 U8587 ( .A(n7401), .ZN(n7396) );
  XNOR2_X1 U8588 ( .A(n8217), .B(n8207), .ZN(n13796) );
  NAND2_X1 U8589 ( .A1(n7399), .A2(n7400), .ZN(n8217) );
  XNOR2_X1 U8590 ( .A(n8331), .B(n8330), .ZN(n10413) );
  NOR2_X1 U8591 ( .A1(n8254), .A2(n7695), .ZN(n6991) );
  XNOR2_X1 U8592 ( .A(n8117), .B(n8116), .ZN(n11828) );
  AND3_X1 U8593 ( .A1(n7996), .A2(n7995), .A3(n6717), .ZN(n8085) );
  XNOR2_X1 U8594 ( .A(n8055), .B(n8054), .ZN(n11430) );
  INV_X1 U8595 ( .A(n7382), .ZN(n6951) );
  INV_X1 U8596 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n8037) );
  NAND2_X1 U8597 ( .A1(n8035), .A2(n8034), .ZN(n8050) );
  NAND2_X1 U8598 ( .A1(n7996), .A2(n7995), .ZN(n7999) );
  NAND2_X1 U8599 ( .A1(n7368), .A2(n7369), .ZN(n7970) );
  NAND2_X1 U8600 ( .A1(n7370), .A2(n7936), .ZN(n7954) );
  NAND2_X1 U8601 ( .A1(n7917), .A2(n7374), .ZN(n7370) );
  OR2_X1 U8602 ( .A1(n7786), .A2(P1_IR_REG_3__SCAN_IN), .ZN(n7788) );
  AND2_X1 U8603 ( .A1(n10158), .A2(P3_ADDR_REG_1__SCAN_IN), .ZN(n7061) );
  INV_X1 U8604 ( .A(n7631), .ZN(n7062) );
  NOR2_X1 U8605 ( .A1(n15502), .A2(n7638), .ZN(n7640) );
  NOR2_X1 U8606 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n7639), .ZN(n7591) );
  AOI21_X1 U8607 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(n7599), .A(n7598), .ZN(
        n7625) );
  NOR2_X1 U8608 ( .A1(n7652), .A2(n7651), .ZN(n7598) );
  AND2_X1 U8609 ( .A1(n7051), .A2(n14800), .ZN(n7658) );
  OAI21_X1 U8610 ( .B1(n14802), .B2(n14801), .A(n7052), .ZN(n7051) );
  AOI21_X1 U8611 ( .B1(n7622), .B2(n7603), .A(n7602), .ZN(n7618) );
  AOI22_X1 U8612 ( .A1(P3_ADDR_REG_13__SCAN_IN), .A2(n14996), .B1(n7614), .B2(
        n7608), .ZN(n7612) );
  AND4_X1 U8613 ( .A1(n9358), .A2(n9357), .A3(n9356), .A4(n9355), .ZN(n11794)
         );
  AOI21_X1 U8614 ( .B1(n7291), .B2(n7290), .A(n6697), .ZN(n7289) );
  INV_X1 U8615 ( .A(n11434), .ZN(n7290) );
  XNOR2_X1 U8616 ( .A(n12449), .B(n12448), .ZN(n12450) );
  NAND2_X1 U8617 ( .A1(n6783), .A2(n7297), .ZN(n12032) );
  AND3_X1 U8618 ( .A1(n9380), .A2(n9379), .A3(n9378), .ZN(n11874) );
  NAND2_X1 U8619 ( .A1(n10691), .A2(n10690), .ZN(n7280) );
  NAND2_X1 U8620 ( .A1(n10691), .A2(n6672), .ZN(n11005) );
  NAND2_X1 U8621 ( .A1(n12383), .A2(n12382), .ZN(n12381) );
  INV_X1 U8622 ( .A(n7298), .ZN(n12394) );
  OAI21_X1 U8623 ( .B1(n12449), .B2(n7302), .A(n7299), .ZN(n7298) );
  NAND2_X1 U8624 ( .A1(n7303), .A2(n12390), .ZN(n7302) );
  INV_X1 U8625 ( .A(n7300), .ZN(n7299) );
  NAND2_X1 U8626 ( .A1(n12461), .A2(n12354), .ZN(n12404) );
  OAI21_X1 U8627 ( .B1(n6784), .B2(n7285), .A(n7283), .ZN(n12402) );
  AND4_X1 U8628 ( .A1(n9287), .A2(n9286), .A3(n9285), .A4(n9284), .ZN(n11314)
         );
  AND3_X1 U8629 ( .A1(n9315), .A2(n9314), .A3(n9313), .ZN(n11155) );
  AND3_X1 U8630 ( .A1(n9623), .A2(n9622), .A3(n9621), .ZN(n12920) );
  NAND2_X1 U8631 ( .A1(n6906), .A2(n9602), .ZN(n12458) );
  NAND2_X1 U8632 ( .A1(n6784), .A2(n12462), .ZN(n12461) );
  OAI21_X1 U8633 ( .B1(n11869), .B2(n7296), .A(n6693), .ZN(n12040) );
  NAND2_X1 U8634 ( .A1(n7294), .A2(n11439), .ZN(n11519) );
  NAND2_X1 U8635 ( .A1(n11435), .A2(n11434), .ZN(n7294) );
  OR2_X1 U8636 ( .A1(n10708), .A2(n10707), .ZN(n12489) );
  NAND2_X1 U8637 ( .A1(n7304), .A2(n7310), .ZN(n12483) );
  NAND2_X1 U8638 ( .A1(n9629), .A2(n9628), .ZN(n12492) );
  NAND2_X1 U8639 ( .A1(n10703), .A2(n15440), .ZN(n12491) );
  OR2_X1 U8640 ( .A1(n10708), .A2(n10706), .ZN(n12500) );
  INV_X1 U8641 ( .A(n12494), .ZN(n12496) );
  NAND2_X1 U8642 ( .A1(n7163), .A2(n7162), .ZN(n7161) );
  INV_X1 U8643 ( .A(n12920), .ZN(n12728) );
  OAI211_X1 U8644 ( .C1(n9607), .C2(n13120), .A(n9606), .B(n9605), .ZN(n12941)
         );
  INV_X1 U8645 ( .A(n12081), .ZN(n12732) );
  INV_X1 U8646 ( .A(n12006), .ZN(n12733) );
  OR2_X1 U8647 ( .A1(n9270), .A2(n10513), .ZN(n9245) );
  INV_X1 U8648 ( .A(P3_ADDR_REG_1__SCAN_IN), .ZN(n10934) );
  AND2_X1 U8649 ( .A1(n10524), .A2(n10519), .ZN(n10578) );
  AOI21_X1 U8650 ( .B1(n10577), .B2(n10524), .A(n10523), .ZN(n10790) );
  INV_X1 U8651 ( .A(P3_ADDR_REG_4__SCAN_IN), .ZN(n15414) );
  OAI21_X1 U8652 ( .B1(n10866), .B2(n10862), .A(n10863), .ZN(n10846) );
  XNOR2_X1 U8653 ( .A(n10895), .B(n10810), .ZN(n10803) );
  NAND2_X1 U8654 ( .A1(n10803), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n10896) );
  AOI21_X1 U8655 ( .B1(n11074), .B2(n11073), .A(n6774), .ZN(n11672) );
  AND2_X1 U8656 ( .A1(n11072), .A2(n11080), .ZN(n6774) );
  XNOR2_X1 U8657 ( .A(n6981), .B(n11659), .ZN(n11077) );
  NAND2_X1 U8658 ( .A1(n11077), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n11658) );
  OAI22_X1 U8659 ( .A1(n11672), .A2(n11671), .B1(n11670), .B2(n11669), .ZN(
        n15419) );
  NAND2_X1 U8660 ( .A1(n11706), .A2(n11653), .ZN(n11654) );
  NAND2_X1 U8661 ( .A1(n11930), .A2(n6755), .ZN(n11933) );
  AOI21_X1 U8662 ( .B1(n12784), .B2(n12783), .A(n12782), .ZN(n12786) );
  AOI21_X1 U8663 ( .B1(n12803), .B2(n12802), .A(n12801), .ZN(n12805) );
  AOI21_X1 U8664 ( .B1(n12810), .B2(P3_REG2_REG_17__SCAN_IN), .A(n6662), .ZN(
        n12844) );
  XNOR2_X1 U8665 ( .A(n12707), .B(n12695), .ZN(n12334) );
  AND2_X1 U8666 ( .A1(n7029), .A2(n12648), .ZN(n12707) );
  NAND2_X1 U8667 ( .A1(n6905), .A2(n7028), .ZN(n7029) );
  NAND2_X1 U8668 ( .A1(n12869), .A2(n9652), .ZN(n12858) );
  XNOR2_X1 U8669 ( .A(n6789), .B(n9666), .ZN(n13042) );
  NAND2_X1 U8670 ( .A1(n6790), .A2(n12646), .ZN(n6789) );
  NAND2_X1 U8671 ( .A1(n12930), .A2(n12937), .ZN(n12932) );
  NAND2_X1 U8672 ( .A1(n9708), .A2(n12522), .ZN(n12930) );
  INV_X1 U8673 ( .A(n13126), .ZN(n12949) );
  NAND2_X1 U8674 ( .A1(n13075), .A2(n9706), .ZN(n12969) );
  NAND2_X1 U8675 ( .A1(n7418), .A2(n12976), .ZN(n13075) );
  NAND2_X1 U8676 ( .A1(n9544), .A2(n9543), .ZN(n12982) );
  NAND2_X1 U8677 ( .A1(n12987), .A2(n9540), .ZN(n12975) );
  INV_X1 U8678 ( .A(n7003), .ZN(n13084) );
  NAND2_X1 U8679 ( .A1(n7462), .A2(n6649), .ZN(n13014) );
  NAND2_X1 U8680 ( .A1(n9466), .A2(n7466), .ZN(n7462) );
  NAND2_X1 U8681 ( .A1(n7414), .A2(n12603), .ZN(n13034) );
  NAND2_X1 U8682 ( .A1(n12152), .A2(n12686), .ZN(n7414) );
  NAND2_X1 U8683 ( .A1(n9466), .A2(n9465), .ZN(n13026) );
  AOI21_X1 U8684 ( .B1(n10369), .B2(n9615), .A(n9457), .ZN(n12510) );
  NAND2_X1 U8685 ( .A1(n7044), .A2(n12591), .ZN(n12127) );
  OR2_X1 U8686 ( .A1(n12078), .A2(n9704), .ZN(n7044) );
  NAND2_X1 U8687 ( .A1(n7479), .A2(n7483), .ZN(n12079) );
  NAND2_X1 U8688 ( .A1(n12004), .A2(n7486), .ZN(n7479) );
  AOI21_X1 U8689 ( .B1(n12004), .B2(n9396), .A(n6699), .ZN(n12068) );
  OAI21_X1 U8690 ( .B1(n11617), .B2(n7015), .A(n7013), .ZN(n12003) );
  NAND2_X1 U8691 ( .A1(n7407), .A2(n9701), .ZN(n11833) );
  NAND2_X1 U8692 ( .A1(n11731), .A2(n9700), .ZN(n7407) );
  NAND2_X1 U8693 ( .A1(n11310), .A2(n7496), .ZN(n11378) );
  NAND2_X1 U8694 ( .A1(n10777), .A2(n12677), .ZN(n10776) );
  NAND2_X1 U8695 ( .A1(n15447), .A2(n12533), .ZN(n10777) );
  AND2_X1 U8696 ( .A1(n10702), .A2(n10701), .ZN(n15463) );
  AND2_X1 U8697 ( .A1(n15464), .A2(n15460), .ZN(n12927) );
  INV_X1 U8698 ( .A(n15463), .ZN(n15440) );
  AND3_X1 U8699 ( .A1(n9281), .A2(n9280), .A3(n9279), .ZN(n11479) );
  INV_X1 U8700 ( .A(n12398), .ZN(n13107) );
  INV_X1 U8701 ( .A(n12372), .ZN(n13111) );
  INV_X1 U8702 ( .A(n12492), .ZN(n9638) );
  AND2_X1 U8703 ( .A1(n9560), .A2(n9559), .ZN(n13134) );
  NAND2_X1 U8704 ( .A1(n9532), .A2(n9531), .ZN(n13139) );
  AND2_X1 U8705 ( .A1(n9735), .A2(n9734), .ZN(n13150) );
  AND2_X1 U8706 ( .A1(n10670), .A2(P3_STATE_REG_SCAN_IN), .ZN(n13151) );
  AOI21_X1 U8707 ( .B1(n6822), .B2(n7189), .A(n6821), .ZN(n12319) );
  AND2_X1 U8708 ( .A1(n14759), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n6821) );
  INV_X1 U8709 ( .A(P3_IR_REG_30__SCAN_IN), .ZN(n9194) );
  INV_X1 U8710 ( .A(n9202), .ZN(n13158) );
  OR2_X1 U8711 ( .A1(n9727), .A2(n9726), .ZN(n12051) );
  OAI21_X1 U8712 ( .B1(n9724), .B2(n6820), .A(n6819), .ZN(n9727) );
  NAND2_X1 U8713 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_24__SCAN_IN), 
        .ZN(n6820) );
  AND2_X1 U8714 ( .A1(n7196), .A2(n7198), .ZN(n9601) );
  OR2_X1 U8715 ( .A1(n9584), .A2(n9583), .ZN(n7196) );
  XNOR2_X1 U8716 ( .A(n9683), .B(n9682), .ZN(n11470) );
  OAI21_X1 U8717 ( .B1(n9684), .B2(P3_IR_REG_21__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n9683) );
  NAND2_X1 U8718 ( .A1(n9684), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9686) );
  INV_X1 U8719 ( .A(n9765), .ZN(n11242) );
  NAND2_X1 U8720 ( .A1(n7172), .A2(n9431), .ZN(n9447) );
  NAND2_X1 U8721 ( .A1(n9429), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n7172) );
  INV_X1 U8722 ( .A(SI_13_), .ZN(n9897) );
  INV_X1 U8723 ( .A(SI_12_), .ZN(n9877) );
  INV_X1 U8724 ( .A(SI_11_), .ZN(n9838) );
  NAND2_X1 U8725 ( .A1(n7180), .A2(n9387), .ZN(n9406) );
  NAND2_X1 U8726 ( .A1(n9386), .A2(n9385), .ZN(n7180) );
  NAND2_X1 U8727 ( .A1(n7185), .A2(n9225), .ZN(n9340) );
  OR2_X1 U8728 ( .A1(n9327), .A2(n6650), .ZN(n7185) );
  INV_X1 U8729 ( .A(SI_5_), .ZN(n10076) );
  OR2_X1 U8730 ( .A1(n9312), .A2(n9311), .ZN(n10874) );
  NAND2_X1 U8731 ( .A1(n13333), .A2(n13223), .ZN(n7069) );
  NAND2_X1 U8732 ( .A1(n13174), .A2(n13173), .ZN(n14840) );
  INV_X1 U8733 ( .A(n7530), .ZN(n13245) );
  NAND2_X1 U8734 ( .A1(n6830), .A2(n13191), .ZN(n13246) );
  CLKBUF_X1 U8735 ( .A(n13277), .Z(n13278) );
  NAND2_X1 U8736 ( .A1(n14850), .A2(n14849), .ZN(n14848) );
  NAND2_X1 U8737 ( .A1(n7078), .A2(n7081), .ZN(n13290) );
  AND2_X1 U8738 ( .A1(n13235), .A2(n13205), .ZN(n13206) );
  CLKBUF_X1 U8739 ( .A(n13298), .Z(n13299) );
  OR2_X1 U8740 ( .A1(n13311), .A2(n7529), .ZN(n7524) );
  NOR2_X1 U8741 ( .A1(n13311), .A2(n7527), .ZN(n7526) );
  AND2_X1 U8742 ( .A1(n7530), .A2(n7529), .ZN(n13310) );
  NAND2_X1 U8743 ( .A1(n11944), .A2(n15188), .ZN(n11951) );
  INV_X1 U8744 ( .A(n13202), .ZN(n13317) );
  NAND2_X1 U8745 ( .A1(n11776), .A2(n11939), .ZN(n11777) );
  NAND2_X1 U8746 ( .A1(n7536), .A2(n11769), .ZN(n11778) );
  AND2_X1 U8747 ( .A1(n10624), .A2(n10623), .ZN(n15190) );
  AND2_X1 U8748 ( .A1(n10622), .A2(n13655), .ZN(n13331) );
  AND2_X1 U8750 ( .A1(n7078), .A2(n6640), .ZN(n13326) );
  INV_X1 U8751 ( .A(n13349), .ZN(n15193) );
  INV_X1 U8752 ( .A(n15198), .ZN(n13344) );
  OR2_X1 U8753 ( .A1(n8413), .A2(n8414), .ZN(n8416) );
  OR2_X1 U8754 ( .A1(n8413), .A2(n8398), .ZN(n8402) );
  CLKBUF_X1 U8755 ( .A(n8866), .Z(n8867) );
  AND2_X1 U8756 ( .A1(n8536), .A2(n8559), .ZN(n15285) );
  NOR2_X1 U8757 ( .A1(n13435), .A2(n13651), .ZN(n13668) );
  INV_X1 U8758 ( .A(n8873), .ZN(n8874) );
  AOI22_X1 U8759 ( .A1(n11029), .A2(n13337), .B1(n13437), .B2(n13355), .ZN(
        n8873) );
  NAND2_X1 U8760 ( .A1(n13448), .A2(n8754), .ZN(n8765) );
  NAND2_X1 U8761 ( .A1(n7436), .A2(n8858), .ZN(n13485) );
  NAND2_X1 U8762 ( .A1(n13492), .A2(n13491), .ZN(n7436) );
  NAND2_X1 U8763 ( .A1(n7238), .A2(n7242), .ZN(n13500) );
  NAND2_X1 U8764 ( .A1(n13521), .A2(n7239), .ZN(n7238) );
  NAND2_X1 U8765 ( .A1(n7247), .A2(n7239), .ZN(n13510) );
  NAND2_X1 U8766 ( .A1(n7247), .A2(n7249), .ZN(n13508) );
  NAND2_X1 U8767 ( .A1(n7257), .A2(n7258), .ZN(n13542) );
  NAND2_X1 U8768 ( .A1(n7442), .A2(n7444), .ZN(n13549) );
  NAND2_X1 U8769 ( .A1(n7261), .A2(n8662), .ZN(n13554) );
  OR2_X1 U8770 ( .A1(n13574), .A2(n8661), .ZN(n7261) );
  AND2_X1 U8771 ( .A1(n8850), .A2(n8849), .ZN(n13565) );
  NAND2_X1 U8772 ( .A1(n7254), .A2(n7252), .ZN(n13600) );
  NAND2_X1 U8773 ( .A1(n7254), .A2(n8623), .ZN(n13598) );
  NAND2_X1 U8774 ( .A1(n12138), .A2(n8589), .ZN(n12156) );
  NAND2_X1 U8775 ( .A1(n10289), .A2(n9085), .ZN(n8524) );
  NAND2_X1 U8776 ( .A1(n11254), .A2(n8476), .ZN(n11450) );
  OR3_X1 U8777 ( .A1(n6620), .A2(n13213), .A3(n8817), .ZN(n13592) );
  INV_X1 U8778 ( .A(n15330), .ZN(n13641) );
  INV_X1 U8779 ( .A(n13612), .ZN(n15324) );
  INV_X1 U8780 ( .A(n13592), .ZN(n15333) );
  OR2_X1 U8781 ( .A1(n6620), .A2(n13429), .ZN(n13612) );
  NAND2_X1 U8782 ( .A1(n15349), .A2(n8811), .ZN(n13655) );
  INV_X1 U8783 ( .A(n15392), .ZN(n15389) );
  INV_X1 U8784 ( .A(n9128), .ZN(n13753) );
  INV_X1 U8785 ( .A(n15383), .ZN(n15382) );
  AND2_X1 U8786 ( .A1(n10631), .A2(n9771), .ZN(n15349) );
  INV_X1 U8787 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n8361) );
  INV_X1 U8788 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n13800) );
  NAND2_X1 U8789 ( .A1(n8778), .A2(n8777), .ZN(n13801) );
  XNOR2_X1 U8790 ( .A(n8789), .B(n8788), .ZN(n12136) );
  NAND2_X1 U8791 ( .A1(n8787), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8789) );
  INV_X1 U8792 ( .A(n9168), .ZN(n11829) );
  INV_X1 U8793 ( .A(n13429), .ZN(n11531) );
  INV_X1 U8794 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n11269) );
  CLKBUF_X1 U8795 ( .A(n8591), .Z(n8592) );
  INV_X1 U8796 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n10488) );
  INV_X1 U8797 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n9828) );
  INV_X1 U8798 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n9821) );
  INV_X1 U8799 ( .A(n15141), .ZN(n11557) );
  NAND2_X1 U8800 ( .A1(n11542), .A2(n6786), .ZN(n11549) );
  NAND2_X1 U8801 ( .A1(n11541), .A2(n6787), .ZN(n6786) );
  INV_X1 U8802 ( .A(n11543), .ZN(n6787) );
  NAND2_X1 U8803 ( .A1(n11549), .A2(n11548), .ZN(n11722) );
  AOI21_X1 U8804 ( .B1(n7334), .B2(n7336), .A(n6706), .ZN(n7331) );
  NAND2_X1 U8805 ( .A1(n7348), .A2(n7351), .ZN(n14892) );
  NAND2_X1 U8806 ( .A1(n6827), .A2(n7353), .ZN(n7348) );
  AND2_X1 U8807 ( .A1(n7322), .A2(n7324), .ZN(n12062) );
  NOR2_X1 U8808 ( .A1(n13833), .A2(n7346), .ZN(n7345) );
  INV_X1 U8809 ( .A(n12236), .ZN(n7346) );
  NAND2_X1 U8810 ( .A1(n7347), .A2(n12236), .ZN(n13834) );
  NAND2_X1 U8811 ( .A1(n11722), .A2(n11721), .ZN(n11723) );
  NOR2_X1 U8812 ( .A1(n10426), .A2(n6657), .ZN(n10434) );
  NAND2_X1 U8813 ( .A1(n13893), .A2(n12248), .ZN(n13845) );
  OAI21_X1 U8814 ( .B1(n12053), .B2(n7319), .A(n7316), .ZN(n7320) );
  AOI21_X1 U8816 ( .B1(n6634), .B2(n7328), .A(n6679), .ZN(n7325) );
  AND2_X1 U8817 ( .A1(n8101), .A2(n8100), .ZN(n14674) );
  OR2_X1 U8818 ( .A1(n13900), .A2(n13901), .ZN(n14890) );
  NAND2_X1 U8819 ( .A1(n12182), .A2(n7323), .ZN(n14905) );
  NAND2_X1 U8820 ( .A1(n7333), .A2(n12283), .ZN(n13930) );
  NAND2_X1 U8821 ( .A1(n11190), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14914) );
  NAND2_X1 U8822 ( .A1(n10411), .A2(n14602), .ZN(n14909) );
  AND2_X1 U8823 ( .A1(n14164), .A2(n14163), .ZN(n14165) );
  OR2_X1 U8824 ( .A1(n8028), .A2(n8027), .ZN(n14582) );
  NAND2_X1 U8825 ( .A1(n7794), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n7710) );
  OR2_X1 U8826 ( .A1(n8244), .A2(n7730), .ZN(n7736) );
  AND2_X1 U8827 ( .A1(n7810), .A2(n7845), .ZN(n14266) );
  INV_X1 U8828 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n10374) );
  AND2_X1 U8829 ( .A1(n15043), .A2(n15042), .ZN(n15044) );
  INV_X1 U8830 ( .A(n14342), .ZN(n14352) );
  NAND2_X1 U8831 ( .A1(n14425), .A2(n8291), .ZN(n14410) );
  AOI21_X1 U8832 ( .B1(n14427), .B2(n14952), .A(n14426), .ZN(n14645) );
  NAND2_X1 U8833 ( .A1(n14462), .A2(n8153), .ZN(n14448) );
  NAND2_X1 U8834 ( .A1(n14486), .A2(n8286), .ZN(n14459) );
  INV_X1 U8835 ( .A(n14674), .ZN(n14518) );
  NAND2_X1 U8836 ( .A1(n7204), .A2(n7206), .ZN(n14511) );
  NAND2_X1 U8837 ( .A1(n7205), .A2(n8068), .ZN(n14522) );
  NAND2_X1 U8838 ( .A1(n8049), .A2(n7210), .ZN(n7205) );
  NAND2_X1 U8839 ( .A1(n14542), .A2(n14067), .ZN(n14524) );
  NAND2_X1 U8840 ( .A1(n8049), .A2(n8048), .ZN(n14535) );
  NAND2_X1 U8841 ( .A1(n7115), .A2(n6632), .ZN(n14694) );
  NAND2_X1 U8842 ( .A1(n14581), .A2(n8014), .ZN(n14578) );
  NAND2_X1 U8843 ( .A1(n8002), .A2(n8001), .ZN(n14590) );
  OR2_X1 U8844 ( .A1(n13959), .A2(n9942), .ZN(n14928) );
  NAND2_X1 U8845 ( .A1(n7219), .A2(n7932), .ZN(n11843) );
  NAND2_X1 U8846 ( .A1(n7915), .A2(n7220), .ZN(n7219) );
  NAND2_X1 U8847 ( .A1(n14596), .A2(n8272), .ZN(n11635) );
  NAND2_X1 U8848 ( .A1(n10748), .A2(n8265), .ZN(n10970) );
  INV_X1 U8849 ( .A(n14570), .ZN(n15081) );
  INV_X1 U8850 ( .A(n15111), .ZN(n13978) );
  NAND2_X1 U8851 ( .A1(n14539), .A2(n10409), .ZN(n14570) );
  AND2_X1 U8852 ( .A1(n8242), .A2(n8241), .ZN(n14365) );
  NAND2_X1 U8853 ( .A1(n14645), .A2(n6779), .ZN(n14722) );
  AND2_X1 U8854 ( .A1(n6780), .A2(n14644), .ZN(n6779) );
  OR2_X1 U8855 ( .A1(n14646), .A2(n14949), .ZN(n6780) );
  INV_X1 U8856 ( .A(n14043), .ZN(n14044) );
  AND2_X2 U8857 ( .A1(n8321), .A2(n8320), .ZN(n9815) );
  OAI21_X1 U8858 ( .B1(n8318), .B2(P1_IR_REG_25__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n8319) );
  AND2_X1 U8859 ( .A1(n7715), .A2(n7355), .ZN(n7354) );
  INV_X1 U8860 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n7355) );
  XNOR2_X1 U8861 ( .A(n9084), .B(n9083), .ZN(n13784) );
  NAND2_X1 U8862 ( .A1(n6796), .A2(n9106), .ZN(n14760) );
  NAND2_X1 U8863 ( .A1(n7390), .A2(n7388), .ZN(n9106) );
  NAND2_X1 U8864 ( .A1(n7390), .A2(n9079), .ZN(n9105) );
  INV_X1 U8865 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n14764) );
  NAND2_X1 U8866 ( .A1(n7714), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7716) );
  INV_X1 U8867 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n14767) );
  INV_X1 U8868 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n12313) );
  INV_X1 U8869 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n11238) );
  NAND2_X1 U8870 ( .A1(n7991), .A2(n7391), .ZN(n7976) );
  AND2_X1 U8871 ( .A1(n7978), .A2(n7959), .ZN(n14993) );
  INV_X1 U8872 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n10151) );
  OAI21_X1 U8873 ( .B1(n7858), .B2(n6932), .A(n6929), .ZN(n7904) );
  INV_X1 U8874 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n9902) );
  NAND2_X1 U8875 ( .A1(n6928), .A2(n6933), .ZN(n7900) );
  NAND2_X1 U8876 ( .A1(n7858), .A2(n7071), .ZN(n6928) );
  INV_X1 U8877 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n9896) );
  NAND2_X1 U8878 ( .A1(n7879), .A2(n6907), .ZN(n9895) );
  NAND2_X1 U8879 ( .A1(n7862), .A2(n7861), .ZN(n7879) );
  NAND2_X1 U8880 ( .A1(n6908), .A2(n6934), .ZN(n6907) );
  INV_X1 U8881 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n9893) );
  OAI21_X1 U8882 ( .B1(n7822), .B2(n7824), .A(n7363), .ZN(n7843) );
  INV_X1 U8883 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n9833) );
  NAND2_X1 U8884 ( .A1(n7826), .A2(n7825), .ZN(n7839) );
  NAND2_X1 U8885 ( .A1(n7822), .A2(n7807), .ZN(n9834) );
  NAND2_X1 U8886 ( .A1(n7786), .A2(n7758), .ZN(n9926) );
  NOR2_X1 U8887 ( .A1(n7658), .A2(n7657), .ZN(n14805) );
  NAND2_X1 U8888 ( .A1(n7060), .A2(n14961), .ZN(n14966) );
  NAND2_X1 U8889 ( .A1(n6778), .A2(n14969), .ZN(n14974) );
  NOR2_X1 U8890 ( .A1(n14974), .A2(n14975), .ZN(n14973) );
  XNOR2_X1 U8891 ( .A(n7053), .B(n7671), .ZN(n14816) );
  NAND2_X1 U8892 ( .A1(n14816), .A2(n14815), .ZN(n14814) );
  AND2_X1 U8893 ( .A1(n6972), .A2(n6969), .ZN(n6968) );
  NAND2_X1 U8894 ( .A1(n7423), .A2(n6756), .ZN(n9770) );
  NAND2_X1 U8895 ( .A1(n7490), .A2(n6757), .ZN(n9759) );
  CLKBUF_X1 U8896 ( .A(n11336), .Z(n11093) );
  NAND2_X1 U8897 ( .A1(n10735), .A2(n10734), .ZN(n10830) );
  NAND2_X1 U8898 ( .A1(n7517), .A2(n11340), .ZN(n11349) );
  NAND2_X1 U8899 ( .A1(n7514), .A2(n10828), .ZN(n10838) );
  NAND2_X1 U8900 ( .A1(n6815), .A2(n6812), .ZN(n14340) );
  NAND2_X1 U8901 ( .A1(n6985), .A2(n14952), .ZN(n6989) );
  NAND2_X1 U8902 ( .A1(n6990), .A2(n6754), .ZN(P1_U3524) );
  NAND2_X1 U8903 ( .A1(n14717), .A2(n15174), .ZN(n6990) );
  OAI222_X1 U8904 ( .A1(n14774), .A2(n14773), .B1(n14761), .B2(n14772), .C1(
        P1_U3086), .C2(n14771), .ZN(P1_U3330) );
  NAND2_X1 U8905 ( .A1(n7046), .A2(n7047), .ZN(n15509) );
  XNOR2_X1 U8906 ( .A(n7065), .B(n7064), .ZN(SUB_1596_U4) );
  XNOR2_X1 U8907 ( .A(n7684), .B(n7717), .ZN(n7064) );
  NAND2_X1 U8908 ( .A1(n14779), .A2(n7066), .ZN(n7065) );
  AND2_X1 U8909 ( .A1(n7268), .A2(n6889), .ZN(n6631) );
  INV_X1 U8910 ( .A(n6627), .ZN(n8467) );
  NAND2_X1 U8911 ( .A1(n12056), .A2(n12055), .ZN(n7322) );
  AND2_X1 U8912 ( .A1(n8281), .A2(n6654), .ZN(n6632) );
  NAND2_X1 U8913 ( .A1(n10292), .A2(n9213), .ZN(n8590) );
  NAND2_X1 U8914 ( .A1(n7322), .A2(n6737), .ZN(n12182) );
  INV_X1 U8915 ( .A(n12565), .ZN(n7472) );
  INV_X1 U8916 ( .A(n14963), .ZN(n7058) );
  INV_X1 U8917 ( .A(n12901), .ZN(n7508) );
  AND2_X1 U8918 ( .A1(n13013), .A2(n7463), .ZN(n6633) );
  AND2_X1 U8919 ( .A1(n7327), .A2(n13817), .ZN(n6634) );
  AND2_X1 U8920 ( .A1(n6684), .A2(n6850), .ZN(n6635) );
  INV_X1 U8921 ( .A(n14607), .ZN(n7110) );
  AND2_X1 U8922 ( .A1(n9136), .A2(n13429), .ZN(n8909) );
  AND2_X1 U8923 ( .A1(n6881), .A2(n13762), .ZN(n6636) );
  OR2_X1 U8924 ( .A1(n14057), .A2(n14091), .ZN(n6637) );
  AND2_X1 U8925 ( .A1(n12736), .A2(n11516), .ZN(n6638) );
  INV_X1 U8926 ( .A(n13901), .ZN(n7353) );
  AND2_X1 U8927 ( .A1(n7092), .A2(n6922), .ZN(n6639) );
  AND2_X1 U8928 ( .A1(n7081), .A2(n6680), .ZN(n6640) );
  INV_X1 U8929 ( .A(n7484), .ZN(n7483) );
  OAI22_X1 U8930 ( .A1(n12681), .A2(n7485), .B1(n12081), .B2(n14827), .ZN(
        n7484) );
  AND2_X1 U8931 ( .A1(n13182), .A2(n13181), .ZN(n6641) );
  AND2_X1 U8932 ( .A1(n8938), .A2(n8937), .ZN(n6642) );
  AND2_X1 U8933 ( .A1(n6631), .A2(n6888), .ZN(n6643) );
  OR2_X1 U8934 ( .A1(n9070), .A2(n9069), .ZN(n6644) );
  AND2_X1 U8935 ( .A1(n14379), .A2(n14378), .ZN(n6645) );
  AND2_X1 U8936 ( .A1(n7105), .A2(n14055), .ZN(n6646) );
  NAND2_X1 U8937 ( .A1(n7867), .A2(n7866), .ZN(n14018) );
  INV_X1 U8938 ( .A(n14018), .ZN(n6920) );
  NAND2_X1 U8939 ( .A1(n7942), .A2(n7941), .ZN(n14040) );
  INV_X1 U8940 ( .A(n14040), .ZN(n7084) );
  INV_X1 U8941 ( .A(n11783), .ZN(n6889) );
  AND2_X1 U8942 ( .A1(n8215), .A2(n13166), .ZN(n6647) );
  INV_X1 U8943 ( .A(n8244), .ZN(n8104) );
  AND2_X1 U8944 ( .A1(n14393), .A2(n8214), .ZN(n6648) );
  OR2_X1 U8945 ( .A1(n13035), .A2(n13016), .ZN(n6649) );
  AND2_X1 U8946 ( .A1(n9828), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n6650) );
  AND2_X1 U8947 ( .A1(n7460), .A2(n7461), .ZN(n6651) );
  AND2_X1 U8948 ( .A1(n11853), .A2(n7968), .ZN(n6652) );
  INV_X1 U8949 ( .A(n8192), .ZN(n6833) );
  INV_X1 U8950 ( .A(n14187), .ZN(n14577) );
  NAND2_X1 U8951 ( .A1(n7459), .A2(n9722), .ZN(n9725) );
  NAND2_X1 U8952 ( .A1(n9658), .A2(n9657), .ZN(n12398) );
  NAND2_X1 U8953 ( .A1(n9116), .A2(n9115), .ZN(n6653) );
  NAND2_X1 U8954 ( .A1(n14705), .A2(n14550), .ZN(n6654) );
  NAND2_X1 U8955 ( .A1(n13524), .A2(n13361), .ZN(n6655) );
  OR2_X1 U8956 ( .A1(n8968), .A2(n8967), .ZN(n6656) );
  INV_X1 U8957 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n9208) );
  AND2_X1 U8958 ( .A1(n10427), .A2(n12288), .ZN(n6657) );
  AND2_X1 U8959 ( .A1(n8979), .A2(n8978), .ZN(n6658) );
  AND2_X1 U8960 ( .A1(n8994), .A2(n8993), .ZN(n6659) );
  AND2_X1 U8961 ( .A1(n9041), .A2(n9040), .ZN(n6660) );
  NAND2_X1 U8962 ( .A1(n13909), .A2(n12262), .ZN(n13816) );
  INV_X1 U8963 ( .A(n9709), .ZN(n12937) );
  AND2_X1 U8964 ( .A1(n7312), .A2(n12364), .ZN(n6661) );
  AND2_X1 U8965 ( .A1(n6867), .A2(n12817), .ZN(n6662) );
  NAND2_X1 U8966 ( .A1(n12492), .A2(n12876), .ZN(n6663) );
  XOR2_X1 U8967 ( .A(n13716), .B(n13255), .Z(n6664) );
  OR2_X1 U8968 ( .A1(n12398), .A2(n12877), .ZN(n12648) );
  INV_X1 U8969 ( .A(n12685), .ZN(n7481) );
  AND2_X1 U8970 ( .A1(n12648), .A2(n12650), .ZN(n12863) );
  INV_X1 U8971 ( .A(n7861), .ZN(n6934) );
  AND2_X1 U8972 ( .A1(n13990), .A2(n11192), .ZN(n6665) );
  NAND2_X1 U8973 ( .A1(n12398), .A2(n12877), .ZN(n12650) );
  INV_X1 U8974 ( .A(n12650), .ZN(n7030) );
  NAND2_X1 U8975 ( .A1(n8687), .A2(n8686), .ZN(n13524) );
  INV_X1 U8976 ( .A(n12604), .ZN(n7413) );
  AND2_X1 U8977 ( .A1(n7492), .A2(n7493), .ZN(n12328) );
  NAND2_X1 U8978 ( .A1(n7457), .A2(n7456), .ZN(n9717) );
  INV_X1 U8979 ( .A(n14100), .ZN(n6936) );
  NAND2_X1 U8980 ( .A1(n8756), .A2(n8755), .ZN(n13676) );
  INV_X1 U8981 ( .A(n13676), .ZN(n6880) );
  NOR2_X1 U8982 ( .A1(n12934), .A2(n9597), .ZN(n6666) );
  AND3_X1 U8983 ( .A1(n7267), .A2(n7266), .A3(n8419), .ZN(n6667) );
  INV_X1 U8984 ( .A(n12902), .ZN(n7507) );
  AND2_X1 U8985 ( .A1(n7663), .A2(n7058), .ZN(n6668) );
  INV_X1 U8986 ( .A(n14698), .ZN(n14556) );
  INV_X1 U8987 ( .A(n12141), .ZN(n7424) );
  AND2_X1 U8988 ( .A1(n9020), .A2(n9019), .ZN(n6669) );
  INV_X1 U8989 ( .A(n12672), .ZN(n9316) );
  AND2_X1 U8990 ( .A1(n12549), .A2(n12554), .ZN(n12672) );
  AND2_X1 U8991 ( .A1(n9058), .A2(n9057), .ZN(n6670) );
  NAND2_X1 U8992 ( .A1(n7981), .A2(n7980), .ZN(n14946) );
  AND2_X1 U8993 ( .A1(n12976), .A2(n9707), .ZN(n6671) );
  AND2_X1 U8994 ( .A1(n10690), .A2(n7279), .ZN(n6672) );
  INV_X1 U8995 ( .A(n14728), .ZN(n7091) );
  INV_X1 U8996 ( .A(n13642), .ZN(n7273) );
  NAND2_X1 U8997 ( .A1(n8580), .A2(n8579), .ZN(n13642) );
  OR2_X1 U8998 ( .A1(n13572), .A2(n13364), .ZN(n6673) );
  AND2_X1 U8999 ( .A1(n10598), .A2(n15354), .ZN(n6674) );
  NOR2_X1 U9000 ( .A1(n7030), .A2(n9710), .ZN(n7028) );
  NAND2_X1 U9001 ( .A1(n13479), .A2(n6881), .ZN(n6883) );
  INV_X1 U9002 ( .A(n11447), .ZN(n11628) );
  AND3_X1 U9003 ( .A1(n9348), .A2(n9347), .A3(n9346), .ZN(n11447) );
  AND4_X1 U9004 ( .A1(n9338), .A2(n9337), .A3(n9336), .A4(n9335), .ZN(n11622)
         );
  AND2_X1 U9005 ( .A1(n14775), .A2(n9905), .ZN(n14481) );
  AND2_X1 U9006 ( .A1(n13175), .A2(n13173), .ZN(n6675) );
  INV_X1 U9007 ( .A(n7207), .ZN(n7206) );
  OAI22_X1 U9008 ( .A1(n8282), .A2(n7208), .B1(n14545), .B2(n14528), .ZN(n7207) );
  AND2_X1 U9009 ( .A1(n12250), .A2(n12248), .ZN(n6676) );
  AND2_X1 U9010 ( .A1(n6961), .A2(n14140), .ZN(n6677) );
  INV_X1 U9011 ( .A(n7121), .ZN(n7120) );
  OR2_X1 U9012 ( .A1(n8292), .A2(n7122), .ZN(n7121) );
  OR2_X1 U9013 ( .A1(n7553), .A2(n8954), .ZN(n6678) );
  AND2_X1 U9014 ( .A1(n12268), .A2(n12267), .ZN(n6679) );
  NAND2_X1 U9015 ( .A1(n13187), .A2(n13186), .ZN(n6680) );
  INV_X1 U9016 ( .A(n14419), .ZN(n14639) );
  AND2_X1 U9017 ( .A1(n13703), .A2(n13360), .ZN(n6681) );
  INV_X1 U9018 ( .A(n11989), .ZN(n7344) );
  OR2_X1 U9019 ( .A1(n6659), .A2(n8996), .ZN(n6682) );
  INV_X1 U9020 ( .A(n13455), .ZN(n13762) );
  NAND2_X1 U9021 ( .A1(n8744), .A2(n8743), .ZN(n13455) );
  AND2_X1 U9022 ( .A1(n12207), .A2(n12206), .ZN(n6683) );
  OR2_X1 U9023 ( .A1(n9047), .A2(n9049), .ZN(n6684) );
  NOR2_X1 U9024 ( .A1(n14040), .A2(n14220), .ZN(n6685) );
  NOR2_X1 U9025 ( .A1(n13698), .A2(n13359), .ZN(n6686) );
  NOR2_X1 U9026 ( .A1(n14029), .A2(n14899), .ZN(n6687) );
  NOR2_X1 U9027 ( .A1(n13609), .A2(n13366), .ZN(n6688) );
  NAND2_X1 U9028 ( .A1(n13134), .A2(n12977), .ZN(n6689) );
  NOR2_X1 U9029 ( .A1(n13557), .A2(n8852), .ZN(n6690) );
  NOR2_X1 U9030 ( .A1(n13609), .A2(n13292), .ZN(n6691) );
  NOR2_X1 U9031 ( .A1(n13145), .A2(n12478), .ZN(n6692) );
  AND2_X1 U9032 ( .A1(n7295), .A2(n12033), .ZN(n6693) );
  AND2_X1 U9033 ( .A1(n14732), .A2(n8287), .ZN(n6694) );
  OR2_X1 U9034 ( .A1(n9119), .A2(n9120), .ZN(n6695) );
  NAND2_X1 U9035 ( .A1(n12648), .A2(n12706), .ZN(n6696) );
  INV_X1 U9036 ( .A(n13969), .ZN(n10561) );
  NAND2_X1 U9037 ( .A1(n7728), .A2(n7086), .ZN(n13969) );
  AND2_X1 U9038 ( .A1(n12736), .A2(n11441), .ZN(n6697) );
  OR2_X1 U9039 ( .A1(n7585), .A2(n7584), .ZN(n6698) );
  INV_X1 U9040 ( .A(n14031), .ZN(n7151) );
  AND2_X1 U9041 ( .A1(n12416), .A2(n12117), .ZN(n6699) );
  AND2_X1 U9042 ( .A1(n7955), .A2(n9877), .ZN(n6700) );
  NOR2_X1 U9043 ( .A1(n13557), .A2(n13363), .ZN(n6701) );
  OR2_X1 U9044 ( .A1(n14537), .A2(n6943), .ZN(n6702) );
  OR2_X1 U9045 ( .A1(n8935), .A2(n8934), .ZN(n6703) );
  AND2_X1 U9046 ( .A1(n9811), .A2(n9213), .ZN(n6704) );
  INV_X1 U9047 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n7701) );
  INV_X1 U9048 ( .A(n7292), .ZN(n7291) );
  NAND2_X1 U9049 ( .A1(n11439), .A2(n7293), .ZN(n7292) );
  AND2_X1 U9050 ( .A1(n9720), .A2(n9719), .ZN(n9747) );
  INV_X1 U9051 ( .A(n9747), .ZN(n6828) );
  NAND2_X1 U9052 ( .A1(n14462), .A2(n7231), .ZN(n6705) );
  AND2_X1 U9053 ( .A1(n12293), .A2(n12292), .ZN(n6706) );
  NAND2_X1 U9054 ( .A1(n12389), .A2(n12891), .ZN(n6707) );
  AND2_X1 U9055 ( .A1(n7558), .A2(n7559), .ZN(n6708) );
  OR2_X1 U9056 ( .A1(n15194), .A2(n11952), .ZN(n6709) );
  INV_X1 U9057 ( .A(n8837), .ZN(n7450) );
  NOR2_X1 U9058 ( .A1(n7557), .A2(n9048), .ZN(n6710) );
  AND2_X1 U9059 ( .A1(n8168), .A2(n14463), .ZN(n6711) );
  NAND2_X1 U9060 ( .A1(n12428), .A2(n7311), .ZN(n6712) );
  INV_X1 U9061 ( .A(n14126), .ZN(n6961) );
  INV_X1 U9062 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n8360) );
  INV_X1 U9063 ( .A(n7211), .ZN(n7210) );
  NAND2_X1 U9064 ( .A1(n6702), .A2(n8048), .ZN(n7211) );
  INV_X1 U9065 ( .A(n7342), .ZN(n7341) );
  OR2_X1 U9066 ( .A1(n11724), .A2(n7343), .ZN(n7342) );
  INV_X1 U9067 ( .A(n14042), .ZN(n7136) );
  INV_X1 U9068 ( .A(n14020), .ZN(n7141) );
  INV_X1 U9069 ( .A(n14009), .ZN(n7146) );
  AND2_X1 U9070 ( .A1(n7492), .A2(n15498), .ZN(n6713) );
  INV_X1 U9071 ( .A(n14178), .ZN(n11222) );
  AND2_X1 U9072 ( .A1(n7083), .A2(n14849), .ZN(n6714) );
  OR2_X1 U9073 ( .A1(n7650), .A2(n7649), .ZN(n6715) );
  OR2_X1 U9074 ( .A1(n13731), .A2(n8848), .ZN(n6716) );
  AND3_X1 U9075 ( .A1(n8037), .A2(n7154), .A3(n7153), .ZN(n6717) );
  AND3_X1 U9076 ( .A1(n14543), .A2(n14061), .A3(n14075), .ZN(n6718) );
  NOR2_X1 U9077 ( .A1(n14183), .A2(n7218), .ZN(n7217) );
  AND2_X1 U9078 ( .A1(n8786), .A2(P2_IR_REG_21__SCAN_IN), .ZN(n6719) );
  AND2_X1 U9079 ( .A1(n12710), .A2(n12712), .ZN(n6720) );
  AND2_X1 U9080 ( .A1(n6636), .A2(n6880), .ZN(n6721) );
  OR2_X1 U9081 ( .A1(n6936), .A2(n14099), .ZN(n6722) );
  OR2_X1 U9082 ( .A1(n8953), .A2(n8955), .ZN(n6723) );
  AND2_X1 U9083 ( .A1(n6989), .A2(n6645), .ZN(n6724) );
  INV_X1 U9084 ( .A(n10779), .ZN(n12677) );
  NAND2_X1 U9085 ( .A1(n12541), .A2(n12542), .ZN(n10779) );
  AND2_X1 U9086 ( .A1(n9213), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n6725) );
  NAND2_X1 U9087 ( .A1(n9026), .A2(n9027), .ZN(n6726) );
  AND2_X1 U9088 ( .A1(n6658), .A2(n6858), .ZN(n6727) );
  AND2_X1 U9089 ( .A1(n7181), .A2(n6893), .ZN(n6728) );
  NOR2_X1 U9090 ( .A1(n8282), .A2(n7209), .ZN(n6729) );
  AND2_X1 U9091 ( .A1(n6682), .A2(n6842), .ZN(n6730) );
  INV_X1 U9092 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n9211) );
  INV_X1 U9093 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n6862) );
  AND2_X1 U9094 ( .A1(n14419), .A2(n14213), .ZN(n6731) );
  INV_X1 U9095 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n7551) );
  NAND2_X1 U9096 ( .A1(n7550), .A2(n9100), .ZN(n6732) );
  INV_X1 U9097 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n7153) );
  INV_X1 U9098 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n7154) );
  AND2_X1 U9099 ( .A1(n8360), .A2(n7551), .ZN(n6733) );
  INV_X1 U9100 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n9822) );
  NAND2_X1 U9101 ( .A1(n8209), .A2(n8208), .ZN(n14629) );
  INV_X1 U9102 ( .A(n14629), .ZN(n6923) );
  INV_X1 U9103 ( .A(n13557), .ZN(n7270) );
  AND2_X1 U9104 ( .A1(n7271), .A2(n6887), .ZN(n6734) );
  OR2_X1 U9105 ( .A1(n14536), .A2(n6911), .ZN(n6735) );
  AND2_X1 U9106 ( .A1(n11858), .A2(n8300), .ZN(n6736) );
  INV_X1 U9107 ( .A(n14536), .ZN(n6910) );
  INV_X1 U9108 ( .A(n8590), .ZN(n8730) );
  INV_X1 U9109 ( .A(n12578), .ZN(n7406) );
  AND2_X1 U9110 ( .A1(n7324), .A2(n12061), .ZN(n6737) );
  OR2_X1 U9111 ( .A1(n14536), .A2(n6914), .ZN(n6738) );
  INV_X1 U9112 ( .A(n7271), .ZN(n13569) );
  NOR2_X1 U9113 ( .A1(n13589), .A2(n13726), .ZN(n7271) );
  INV_X1 U9114 ( .A(n13703), .ZN(n6884) );
  NAND2_X1 U9115 ( .A1(n7274), .A2(n6879), .ZN(n6739) );
  AND2_X1 U9116 ( .A1(n8990), .A2(n8989), .ZN(n6740) );
  AND2_X1 U9117 ( .A1(n12355), .A2(n12977), .ZN(n6741) );
  AND2_X1 U9118 ( .A1(n14929), .A2(n7990), .ZN(n6742) );
  AND2_X1 U9119 ( .A1(n8575), .A2(n8574), .ZN(n6743) );
  AND2_X1 U9120 ( .A1(n7219), .A2(n7217), .ZN(n6744) );
  AND2_X1 U9121 ( .A1(n13002), .A2(n9518), .ZN(n6745) );
  AND3_X1 U9122 ( .A1(n8067), .A2(n8066), .A3(n8065), .ZN(n14551) );
  INV_X1 U9123 ( .A(n14551), .ZN(n6943) );
  INV_X1 U9124 ( .A(n9696), .ZN(n7493) );
  INV_X1 U9125 ( .A(SI_14_), .ZN(n10197) );
  NOR2_X1 U9126 ( .A1(n12070), .A2(n14822), .ZN(n6746) );
  NAND2_X1 U9127 ( .A1(n7115), .A2(n6654), .ZN(n6747) );
  INV_X1 U9128 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n7174) );
  OR2_X1 U9129 ( .A1(n13762), .A2(n13749), .ZN(n6748) );
  AND3_X1 U9130 ( .A1(n7996), .A2(n7995), .A3(n7154), .ZN(n8038) );
  OR2_X1 U9131 ( .A1(n6923), .A2(n14748), .ZN(n6749) );
  OR2_X1 U9132 ( .A1(n6923), .A2(n14686), .ZN(n6750) );
  AND2_X1 U9133 ( .A1(n6643), .A2(n14871), .ZN(n6751) );
  OR2_X1 U9134 ( .A1(n8992), .A2(n6740), .ZN(n6752) );
  AND2_X1 U9135 ( .A1(n6783), .A2(n11868), .ZN(n6753) );
  AND2_X2 U9136 ( .A1(n11365), .A2(n9769), .ZN(n15498) );
  INV_X1 U9137 ( .A(n15498), .ZN(n6791) );
  NAND2_X1 U9138 ( .A1(n11393), .A2(n15440), .ZN(n15464) );
  AND2_X1 U9139 ( .A1(n10916), .A2(n9110), .ZN(n8890) );
  AND2_X1 U9140 ( .A1(n14360), .A2(n14602), .ZN(n15105) );
  NAND2_X1 U9141 ( .A1(n14539), .A2(n14917), .ZN(n14557) );
  INV_X1 U9142 ( .A(n13630), .ZN(n7272) );
  INV_X1 U9143 ( .A(n14528), .ZN(n6915) );
  NOR2_X1 U9144 ( .A1(n11636), .A2(n7109), .ZN(n7108) );
  NOR2_X1 U9145 ( .A1(n11697), .A2(n14910), .ZN(n7085) );
  INV_X1 U9146 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7176) );
  NAND2_X1 U9147 ( .A1(n8538), .A2(n8537), .ZN(n15194) );
  INV_X1 U9148 ( .A(n15194), .ZN(n6888) );
  OR2_X1 U9149 ( .A1(n15174), .A2(n8230), .ZN(n6754) );
  NAND2_X1 U9150 ( .A1(n7915), .A2(n7914), .ZN(n11693) );
  OR2_X1 U9151 ( .A1(n11932), .A2(n11931), .ZN(n6755) );
  NAND2_X1 U9152 ( .A1(n8119), .A2(n8118), .ZN(n14739) );
  INV_X1 U9153 ( .A(n14739), .ZN(n6912) );
  OR2_X1 U9154 ( .A1(P3_REG1_REG_29__SCAN_IN), .A2(n15498), .ZN(n6756) );
  NOR2_X1 U9155 ( .A1(n11859), .A2(n14043), .ZN(n11858) );
  OR2_X1 U9156 ( .A1(n15493), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n6757) );
  AND2_X1 U9157 ( .A1(n14596), .A2(n7108), .ZN(n6758) );
  AND2_X1 U9158 ( .A1(n7294), .A2(n7291), .ZN(n6759) );
  OR2_X1 U9159 ( .A1(n8215), .A2(n13166), .ZN(n6760) );
  AND2_X1 U9160 ( .A1(n11722), .A2(n7341), .ZN(n6761) );
  AND2_X1 U9161 ( .A1(n7536), .A2(n7535), .ZN(n6762) );
  AND2_X1 U9162 ( .A1(n14057), .A2(n14056), .ZN(n14592) );
  INV_X1 U9163 ( .A(n14592), .ZN(n7104) );
  AND2_X1 U9164 ( .A1(n8206), .A2(SI_26_), .ZN(n6763) );
  INV_X1 U9165 ( .A(n7398), .ZN(n7397) );
  NAND2_X1 U9166 ( .A1(n7400), .A2(n6760), .ZN(n7398) );
  AND2_X1 U9167 ( .A1(n7089), .A2(n7090), .ZN(n6764) );
  INV_X1 U9168 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n11830) );
  INV_X1 U9169 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n11291) );
  INV_X1 U9170 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n11532) );
  OR2_X1 U9171 ( .A1(n15498), .A2(P3_REG1_REG_28__SCAN_IN), .ZN(n6765) );
  INV_X2 U9172 ( .A(n15491), .ZN(n15493) );
  OR2_X1 U9173 ( .A1(P3_REG0_REG_28__SCAN_IN), .A2(n15493), .ZN(n6766) );
  INV_X1 U9174 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n6806) );
  AND2_X1 U9175 ( .A1(n11310), .A2(n9318), .ZN(n6767) );
  AND2_X1 U9176 ( .A1(n7474), .A2(n7473), .ZN(n6768) );
  NAND2_X1 U9177 ( .A1(n8812), .A2(n13655), .ZN(n13643) );
  NAND2_X1 U9178 ( .A1(n8299), .A2(n8298), .ZN(n14952) );
  INV_X1 U9179 ( .A(n14952), .ZN(n15075) );
  INV_X1 U9180 ( .A(n12784), .ZN(n6775) );
  NOR2_X1 U9181 ( .A1(n9265), .A2(n12663), .ZN(n6769) );
  INV_X1 U9182 ( .A(n10709), .ZN(n10781) );
  INV_X1 U9183 ( .A(n15370), .ZN(n7268) );
  INV_X1 U9184 ( .A(n13436), .ZN(n7380) );
  XNOR2_X1 U9185 ( .A(n10659), .B(n10660), .ZN(n10643) );
  OR2_X1 U9186 ( .A1(n9265), .A2(n13155), .ZN(n6770) );
  AND2_X1 U9187 ( .A1(n12002), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n6771) );
  INV_X1 U9188 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n14752) );
  INV_X1 U9189 ( .A(n12658), .ZN(n7189) );
  AND2_X1 U9190 ( .A1(n9210), .A2(n7509), .ZN(n12320) );
  INV_X1 U9191 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n6803) );
  INV_X1 U9192 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n7052) );
  INV_X1 U9193 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6811) );
  INV_X1 U9194 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n7360) );
  INV_X1 U9195 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n6823) );
  OAI222_X1 U9196 ( .A1(n14774), .A2(n9808), .B1(n14761), .B2(n9807), .C1(
        P1_U3086), .C2(n9928), .ZN(P1_U3352) );
  OAI222_X1 U9197 ( .A1(n14774), .A2(n12135), .B1(n14761), .B2(n12137), .C1(
        P1_U3086), .C2(n12134), .ZN(P1_U3331) );
  OAI222_X1 U9198 ( .A1(n14774), .A2(n14767), .B1(n14761), .B2(n14766), .C1(
        P1_U3086), .C2(n6625), .ZN(P1_U3328) );
  NAND2_X2 U9199 ( .A1(n7088), .A2(P1_U3086), .ZN(n14774) );
  OAI222_X1 U9200 ( .A1(n14774), .A2(n14764), .B1(n14761), .B2(n14763), .C1(
        n14762), .C2(P1_U3086), .ZN(P1_U3326) );
  OAI222_X1 U9201 ( .A1(n14774), .A2(n12313), .B1(n14761), .B2(n12327), .C1(
        n13959), .C2(P1_U3086), .ZN(P1_U3335) );
  OAI222_X1 U9202 ( .A1(n14774), .A2(n11832), .B1(n14761), .B2(n11831), .C1(
        P1_U3086), .C2(n14155), .ZN(P1_U3334) );
  OAI222_X1 U9203 ( .A1(n14774), .A2(n11431), .B1(n14761), .B2(n11432), .C1(
        P1_U3086), .C2(n14329), .ZN(P1_U3337) );
  OAI222_X1 U9204 ( .A1(n14774), .A2(n7176), .B1(n14761), .B2(n11533), .C1(
        P1_U3086), .C2(n14917), .ZN(P1_U3336) );
  OAI222_X1 U9205 ( .A1(n14774), .A2(n10553), .B1(n14761), .B2(n10552), .C1(
        n10551), .C2(P1_U3086), .ZN(P1_U3342) );
  OAI222_X1 U9206 ( .A1(n14774), .A2(n11238), .B1(n14761), .B2(n11268), .C1(
        n15036), .C2(P1_U3086), .ZN(P1_U3339) );
  OAI222_X1 U9207 ( .A1(n14774), .A2(n9902), .B1(n14761), .B2(n9901), .C1(
        n10984), .C2(P1_U3086), .ZN(P1_U3346) );
  OAI222_X1 U9208 ( .A1(n14774), .A2(n10151), .B1(n14761), .B2(n9939), .C1(
        n10997), .C2(P1_U3086), .ZN(P1_U3345) );
  OAI222_X1 U9209 ( .A1(n14774), .A2(n9893), .B1(n14761), .B2(n9892), .C1(
        n10983), .C2(P1_U3086), .ZN(P1_U3348) );
  OAI222_X1 U9210 ( .A1(n14774), .A2(n9896), .B1(n14761), .B2(n9895), .C1(
        n10990), .C2(P1_U3086), .ZN(P1_U3347) );
  OAI222_X1 U9211 ( .A1(n14774), .A2(n9833), .B1(n14761), .B2(n9832), .C1(
        n10383), .C2(P1_U3086), .ZN(P1_U3349) );
  OAI222_X1 U9212 ( .A1(n14774), .A2(n6811), .B1(n14761), .B2(n9834), .C1(
        n9931), .C2(P1_U3086), .ZN(P1_U3350) );
  OAI222_X1 U9213 ( .A1(n14774), .A2(n9809), .B1(n14761), .B2(n9819), .C1(
        n9926), .C2(P1_U3086), .ZN(P1_U3353) );
  OAI222_X1 U9214 ( .A1(n14774), .A2(n7360), .B1(n14761), .B2(n9823), .C1(
        n10465), .C2(P1_U3086), .ZN(P1_U3351) );
  AOI21_X1 U9215 ( .B1(n12812), .B2(n12817), .A(n12811), .ZN(n12829) );
  INV_X1 U9216 ( .A(n12817), .ZN(n6866) );
  XNOR2_X1 U9217 ( .A(n12818), .B(n12817), .ZN(n12816) );
  NAND2_X2 U9218 ( .A1(n7088), .A2(P3_U3151), .ZN(n13167) );
  NAND2_X1 U9219 ( .A1(n6814), .A2(n6813), .ZN(n6812) );
  NOR2_X1 U9220 ( .A1(n15061), .A2(n14313), .ZN(n14314) );
  INV_X1 U9221 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n14979) );
  OR2_X1 U9222 ( .A1(n10749), .A2(n7000), .ZN(n6997) );
  NAND2_X1 U9223 ( .A1(n6781), .A2(n14447), .ZN(n14443) );
  NAND2_X1 U9224 ( .A1(n14598), .A2(n7108), .ZN(n6983) );
  NOR2_X1 U9225 ( .A1(n14634), .A2(n14633), .ZN(n14718) );
  INV_X1 U9226 ( .A(n9720), .ZN(n9210) );
  INV_X1 U9227 ( .A(n9187), .ZN(n7031) );
  INV_X1 U9228 ( .A(P3_IR_REG_13__SCAN_IN), .ZN(n9417) );
  NAND2_X1 U9229 ( .A1(n12861), .A2(n9668), .ZN(n9681) );
  NOR2_X1 U9230 ( .A1(n7569), .A2(n7472), .ZN(n7471) );
  NAND2_X1 U9231 ( .A1(n9568), .A2(n7579), .ZN(n7489) );
  NAND2_X1 U9232 ( .A1(n9599), .A2(n9598), .ZN(n12915) );
  NAND2_X1 U9233 ( .A1(n7491), .A2(n6713), .ZN(n7423) );
  OR2_X1 U9234 ( .A1(n7001), .A2(n7000), .ZN(n6999) );
  INV_X1 U9235 ( .A(n8266), .ZN(n7095) );
  INV_X1 U9236 ( .A(n14440), .ZN(n6781) );
  NAND2_X1 U9237 ( .A1(n11224), .A2(n8271), .ZN(n14598) );
  NAND2_X1 U9238 ( .A1(n6983), .A2(n7107), .ZN(n11695) );
  NAND2_X1 U9239 ( .A1(n14542), .A2(n7100), .ZN(n14526) );
  NAND2_X1 U9240 ( .A1(n14494), .A2(n7097), .ZN(n6995) );
  INV_X1 U9241 ( .A(n7569), .ZN(n7473) );
  NAND2_X1 U9242 ( .A1(n8820), .A2(n8819), .ZN(n10764) );
  NAND2_X1 U9243 ( .A1(n8863), .A2(n8862), .ZN(n13457) );
  NAND2_X1 U9244 ( .A1(n13684), .A2(n6748), .ZN(P2_U3527) );
  AOI21_X2 U9245 ( .B1(n13460), .B2(n13459), .A(n13458), .ZN(n13681) );
  INV_X2 U9246 ( .A(n11203), .ZN(n10736) );
  NAND2_X2 U9247 ( .A1(n8422), .A2(n8421), .ZN(n11203) );
  OAI22_X2 U9248 ( .A1(n13528), .A2(n8855), .B1(n13770), .B2(n13361), .ZN(
        n13504) );
  NAND2_X1 U9249 ( .A1(n13459), .A2(n6788), .ZN(n8864) );
  OAI21_X1 U9250 ( .B1(n14971), .B2(n14970), .A(n7666), .ZN(n6778) );
  NAND2_X1 U9251 ( .A1(n7049), .A2(n7048), .ZN(n7047) );
  NAND2_X1 U9252 ( .A1(n14792), .A2(n7656), .ZN(n14802) );
  NAND2_X1 U9253 ( .A1(n7662), .A2(n7660), .ZN(n7663) );
  NAND2_X1 U9254 ( .A1(n8081), .A2(n8080), .ZN(n8099) );
  NOR2_X1 U9255 ( .A1(n7256), .A2(n13541), .ZN(n7255) );
  OAI21_X1 U9256 ( .B1(n8675), .B2(n8144), .A(n8143), .ZN(n8156) );
  NOR2_X1 U9257 ( .A1(n14375), .A2(n15075), .ZN(n6984) );
  OAI211_X1 U9258 ( .C1(n14628), .C2(n14949), .A(n6987), .B(n6986), .ZN(n14717) );
  NAND2_X1 U9259 ( .A1(n7347), .A2(n7345), .ZN(n13835) );
  NOR2_X1 U9260 ( .A1(n10496), .A2(n10495), .ZN(n10499) );
  OR2_X2 U9261 ( .A1(n8410), .A2(n8409), .ZN(n15354) );
  NAND3_X1 U9262 ( .A1(n7515), .A2(n10734), .A3(n10735), .ZN(n7514) );
  NAND2_X2 U9263 ( .A1(n10664), .A2(n10665), .ZN(n10735) );
  NAND2_X1 U9264 ( .A1(n13269), .A2(n13268), .ZN(n13267) );
  NAND2_X1 U9265 ( .A1(n7525), .A2(n7524), .ZN(n13309) );
  NAND2_X1 U9266 ( .A1(n10926), .A2(n10925), .ZN(n11092) );
  OR2_X1 U9267 ( .A1(n12211), .A2(n12210), .ZN(n13939) );
  NAND2_X1 U9268 ( .A1(n13835), .A2(n12244), .ZN(n13895) );
  NAND2_X1 U9269 ( .A1(n13923), .A2(n13924), .ZN(n7347) );
  NAND2_X1 U9270 ( .A1(n11549), .A2(n7339), .ZN(n7338) );
  NOR2_X1 U9271 ( .A1(n10499), .A2(n10498), .ZN(n11172) );
  NAND2_X1 U9272 ( .A1(n6785), .A2(n7329), .ZN(n10431) );
  NAND2_X1 U9273 ( .A1(n10428), .A2(n14231), .ZN(n6785) );
  NAND2_X1 U9274 ( .A1(n7332), .A2(n7331), .ZN(n13808) );
  NAND2_X2 U9275 ( .A1(n7356), .A2(n7357), .ZN(n6834) );
  OAI21_X1 U9276 ( .B1(n7437), .B2(n13491), .A(n13486), .ZN(n7432) );
  INV_X1 U9277 ( .A(n7432), .ZN(n7431) );
  NAND2_X2 U9278 ( .A1(n9905), .A2(n7088), .ZN(n8083) );
  NAND2_X1 U9279 ( .A1(n6802), .A2(n6729), .ZN(n7204) );
  NAND2_X1 U9280 ( .A1(n14391), .A2(n14394), .ZN(n14393) );
  OR2_X1 U9281 ( .A1(n13976), .A2(n15111), .ZN(n7761) );
  NAND2_X1 U9282 ( .A1(n14475), .A2(n14484), .ZN(n14474) );
  NAND2_X1 U9283 ( .A1(n7230), .A2(n7229), .ZN(n14428) );
  NAND2_X1 U9284 ( .A1(n6801), .A2(n7217), .ZN(n7214) );
  NAND2_X1 U9285 ( .A1(n14720), .A2(n6749), .ZN(P1_U3523) );
  NAND2_X1 U9286 ( .A1(n14636), .A2(n6750), .ZN(P1_U3555) );
  INV_X1 U9287 ( .A(n8049), .ZN(n6802) );
  INV_X1 U9288 ( .A(n7915), .ZN(n6801) );
  INV_X1 U9289 ( .A(n14170), .ZN(n10745) );
  NAND2_X1 U9290 ( .A1(n7856), .A2(n7855), .ZN(n11219) );
  AOI21_X1 U9291 ( .B1(n14412), .B2(n14409), .A(n6731), .ZN(n14391) );
  OAI21_X1 U9292 ( .B1(n12012), .B2(n8841), .A(n8842), .ZN(n12142) );
  INV_X1 U9293 ( .A(n12873), .ZN(n6790) );
  NAND2_X1 U9294 ( .A1(n9224), .A2(n9223), .ZN(n9327) );
  NAND2_X1 U9295 ( .A1(n9361), .A2(n9359), .ZN(n9229) );
  NAND2_X1 U9296 ( .A1(n9570), .A2(n9571), .ZN(n6794) );
  NAND2_X1 U9297 ( .A1(n9218), .A2(n9217), .ZN(n9277) );
  OAI21_X1 U9298 ( .B1(n13105), .B2(n6791), .A(n6765), .ZN(n13043) );
  OAI21_X1 U9299 ( .B1(n13105), .B2(n15491), .A(n6766), .ZN(n13106) );
  NAND2_X1 U9300 ( .A1(n6792), .A2(n6716), .ZN(n8850) );
  AND2_X1 U9301 ( .A1(n8358), .A2(n6733), .ZN(n7262) );
  NAND2_X1 U9302 ( .A1(n8860), .A2(n8859), .ZN(n13463) );
  NAND2_X1 U9304 ( .A1(n9811), .A2(n6800), .ZN(n8386) );
  NAND2_X1 U9305 ( .A1(n7453), .A2(n7452), .ZN(n13578) );
  NAND2_X1 U9306 ( .A1(n7441), .A2(n7439), .ZN(n13534) );
  XNOR2_X2 U9307 ( .A(n10648), .B(n8388), .ZN(n9796) );
  INV_X1 U9308 ( .A(n13578), .ZN(n6792) );
  NAND3_X1 U9309 ( .A1(n12655), .A2(n6795), .A3(n12706), .ZN(n12662) );
  NAND3_X2 U9310 ( .A1(n8417), .A2(n8416), .A3(n7234), .ZN(n13381) );
  NAND2_X1 U9311 ( .A1(n9500), .A2(n9501), .ZN(n9502) );
  NAND2_X1 U9312 ( .A1(n9520), .A2(n9519), .ZN(n9522) );
  NAND2_X1 U9313 ( .A1(n8827), .A2(n8826), .ZN(n11258) );
  XNOR2_X1 U9314 ( .A(n9609), .B(n6823), .ZN(n9610) );
  NAND2_X1 U9315 ( .A1(n12704), .A2(n12705), .ZN(n7166) );
  NAND2_X1 U9316 ( .A1(n9105), .A2(n9104), .ZN(n6796) );
  NAND2_X1 U9317 ( .A1(n8133), .A2(n8132), .ZN(n8142) );
  AOI21_X1 U9318 ( .B1(n6833), .B2(n9247), .A(n9885), .ZN(n6832) );
  AOI21_X1 U9319 ( .B1(n14205), .B2(n14204), .A(n14203), .ZN(n14210) );
  NAND2_X1 U9320 ( .A1(n10887), .A2(n10888), .ZN(n10926) );
  XNOR2_X1 U9321 ( .A(n10638), .B(n10652), .ZN(n10659) );
  MUX2_X2 U9322 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8375), .S(
        P2_IR_REG_27__SCAN_IN), .Z(n7427) );
  AOI21_X2 U9323 ( .B1(n13198), .B2(n13197), .A(n13309), .ZN(n13269) );
  AND3_X4 U9324 ( .A1(n8387), .A2(n8386), .A3(n8385), .ZN(n10648) );
  NAND2_X1 U9325 ( .A1(n7366), .A2(n8155), .ZN(n7365) );
  NAND2_X1 U9326 ( .A1(n8076), .A2(n8075), .ZN(n8081) );
  INV_X1 U9327 ( .A(n7973), .ZN(n6797) );
  NAND2_X1 U9328 ( .A1(n10759), .A2(n8437), .ZN(n10959) );
  NAND2_X1 U9329 ( .A1(n13653), .A2(n8411), .ZN(n10594) );
  OAI22_X1 U9330 ( .A1(n13478), .A2(n8729), .B1(n6882), .B2(n13358), .ZN(
        n13475) );
  NAND2_X1 U9331 ( .A1(n11255), .A2(n11259), .ZN(n11254) );
  NAND2_X2 U9332 ( .A1(n13544), .A2(n8685), .ZN(n13521) );
  XNOR2_X1 U9333 ( .A(n7585), .B(n7584), .ZN(n7628) );
  NAND2_X1 U9334 ( .A1(n14802), .A2(n14801), .ZN(n14800) );
  XNOR2_X1 U9335 ( .A(n7642), .B(n7641), .ZN(n15507) );
  NAND2_X1 U9336 ( .A1(n15507), .A2(n15506), .ZN(n15505) );
  NOR2_X1 U9337 ( .A1(n13226), .A2(n7523), .ZN(n7522) );
  NAND2_X1 U9338 ( .A1(n13324), .A2(n7526), .ZN(n7525) );
  INV_X1 U9339 ( .A(n8801), .ZN(n8799) );
  INV_X1 U9340 ( .A(n10829), .ZN(n7515) );
  NAND2_X1 U9341 ( .A1(n12276), .A2(n12275), .ZN(n13863) );
  AND2_X1 U9342 ( .A1(n10399), .A2(n10400), .ZN(n10426) );
  NOR2_X1 U9343 ( .A1(n7993), .A2(n7994), .ZN(n6992) );
  NAND2_X1 U9344 ( .A1(n7286), .A2(n11322), .ZN(n6829) );
  NAND2_X2 U9345 ( .A1(n10292), .A2(n7088), .ZN(n8438) );
  OAI21_X2 U9346 ( .B1(n13629), .B2(n7251), .A(n7250), .ZN(n13582) );
  NAND2_X1 U9347 ( .A1(n8521), .A2(n8520), .ZN(n11757) );
  NAND2_X1 U9348 ( .A1(n11452), .A2(n8492), .ZN(n11558) );
  OAI21_X2 U9349 ( .B1(n14493), .B2(n14496), .A(n8126), .ZN(n14475) );
  NAND2_X1 U9350 ( .A1(n6804), .A2(n7567), .ZN(n14397) );
  NAND2_X1 U9351 ( .A1(n14395), .A2(n14394), .ZN(n6804) );
  NAND2_X1 U9352 ( .A1(n6826), .A2(n14178), .ZN(n11224) );
  NAND3_X1 U9353 ( .A1(n6999), .A2(n11042), .A3(n6997), .ZN(n6996) );
  AND2_X2 U9354 ( .A1(n12719), .A2(n12718), .ZN(n12726) );
  OR2_X2 U9355 ( .A1(n12700), .A2(n12645), .ZN(n12651) );
  XNOR2_X2 U9356 ( .A(n15354), .B(n13382), .ZN(n13658) );
  NAND2_X1 U9357 ( .A1(n7763), .A2(n7753), .ZN(n9819) );
  AOI21_X2 U9358 ( .B1(n12668), .B2(n12667), .A(n12701), .ZN(n12704) );
  INV_X4 U9359 ( .A(n6834), .ZN(n8192) );
  MUX2_X1 U9360 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .S(n6834), .Z(n7748) );
  NAND2_X1 U9361 ( .A1(n7430), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8376) );
  NAND2_X1 U9362 ( .A1(n7425), .A2(n7424), .ZN(n8844) );
  AND2_X2 U9363 ( .A1(n6809), .A2(n9342), .ZN(n7457) );
  OR2_X2 U9364 ( .A1(n11007), .A2(n11008), .ZN(n11151) );
  INV_X1 U9365 ( .A(n10697), .ZN(n7279) );
  NAND2_X1 U9366 ( .A1(n12814), .A2(n12813), .ZN(n12830) );
  NOR2_X1 U9367 ( .A1(n10936), .A2(n10937), .ZN(n10935) );
  INV_X1 U9368 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n7717) );
  NAND3_X1 U9369 ( .A1(n7991), .A2(n7391), .A3(n7974), .ZN(n7992) );
  NAND2_X1 U9370 ( .A1(n8035), .A2(n7382), .ZN(n8073) );
  NAND2_X1 U9371 ( .A1(n7449), .A2(n7446), .ZN(n11963) );
  INV_X1 U9372 ( .A(n12142), .ZN(n7425) );
  NAND2_X1 U9373 ( .A1(n10597), .A2(n10596), .ZN(n8820) );
  NAND3_X1 U9374 ( .A1(n7514), .A2(n7516), .A3(n10828), .ZN(n10886) );
  NAND2_X2 U9375 ( .A1(n13843), .A2(n12253), .ZN(n13910) );
  NAND2_X1 U9376 ( .A1(n8378), .A2(n8377), .ZN(n7426) );
  NOR2_X2 U9377 ( .A1(n13351), .A2(n13350), .ZN(n13348) );
  NAND2_X1 U9378 ( .A1(n7080), .A2(n7079), .ZN(n13324) );
  NAND2_X1 U9379 ( .A1(n12443), .A2(n12442), .ZN(n12441) );
  NAND2_X1 U9380 ( .A1(n12499), .A2(n12498), .ZN(n12497) );
  NOR2_X1 U9381 ( .A1(n10680), .A2(n7287), .ZN(n7286) );
  NAND2_X1 U9382 ( .A1(n7124), .A2(n7123), .ZN(n14395) );
  INV_X1 U9383 ( .A(n11223), .ZN(n6826) );
  NAND2_X1 U9384 ( .A1(n9541), .A2(n9542), .ZN(n7177) );
  XNOR2_X1 U9385 ( .A(n9554), .B(n12325), .ZN(n9555) );
  AND2_X2 U9386 ( .A1(n7192), .A2(n7193), .ZN(n9609) );
  NAND2_X1 U9387 ( .A1(n6995), .A2(n7096), .ZN(n14440) );
  NAND2_X1 U9388 ( .A1(n6996), .A2(n8267), .ZN(n15074) );
  INV_X1 U9389 ( .A(n7093), .ZN(n7000) );
  NAND2_X1 U9390 ( .A1(n7326), .A2(n7325), .ZN(n13885) );
  NAND2_X1 U9391 ( .A1(n6992), .A2(n6991), .ZN(n8311) );
  OR2_X1 U9392 ( .A1(n10429), .A2(n10389), .ZN(n10392) );
  NAND2_X1 U9393 ( .A1(n7282), .A2(n7281), .ZN(n12358) );
  NAND2_X2 U9394 ( .A1(n11151), .A2(n11150), .ZN(n11435) );
  NAND2_X4 U9395 ( .A1(n6829), .A2(n7288), .ZN(n12392) );
  NAND2_X1 U9396 ( .A1(n13219), .A2(n13218), .ZN(n13333) );
  AND2_X1 U9397 ( .A1(n6832), .A2(n6831), .ZN(n7721) );
  INV_X1 U9398 ( .A(n7862), .ZN(n6908) );
  OAI21_X1 U9399 ( .B1(n12848), .B2(n15406), .A(n6968), .ZN(P3_U3201) );
  NAND3_X1 U9400 ( .A1(n6838), .A2(n6644), .A3(n6732), .ZN(n6837) );
  NAND3_X1 U9401 ( .A1(n7571), .A2(n8988), .A3(n6752), .ZN(n6841) );
  NAND2_X1 U9402 ( .A1(n6841), .A2(n6730), .ZN(n7555) );
  NAND2_X1 U9403 ( .A1(n9023), .A2(n6845), .ZN(n6844) );
  NAND2_X1 U9404 ( .A1(n9043), .A2(n6635), .ZN(n6848) );
  NAND2_X1 U9405 ( .A1(n6848), .A2(n6849), .ZN(n9054) );
  INV_X1 U9406 ( .A(n9042), .ZN(n6852) );
  AOI21_X1 U9407 ( .B1(n6855), .B2(n7561), .A(n6727), .ZN(n6853) );
  NAND2_X1 U9408 ( .A1(n8974), .A2(n6855), .ZN(n6854) );
  OAI21_X2 U9409 ( .B1(n9834), .B2(n9107), .A(n8444), .ZN(n10965) );
  NAND2_X2 U9410 ( .A1(n7806), .A2(n7805), .ZN(n7822) );
  MUX2_X1 U9411 ( .A(n10532), .B(P3_REG2_REG_2__SCAN_IN), .S(n10533), .Z(
        n10567) );
  INV_X2 U9412 ( .A(n10292), .ZN(n8636) );
  NAND2_X2 U9413 ( .A1(n8868), .A2(n8866), .ZN(n10292) );
  NAND3_X1 U9414 ( .A1(n8867), .A2(n8868), .A3(n15208), .ZN(n8385) );
  NAND2_X1 U9415 ( .A1(n7426), .A2(n8379), .ZN(n8866) );
  INV_X1 U9416 ( .A(n6883), .ZN(n13468) );
  NAND2_X1 U9417 ( .A1(n7269), .A2(n6751), .ZN(n12020) );
  NAND2_X1 U9418 ( .A1(n9306), .A2(n9304), .ZN(n9224) );
  NAND2_X1 U9419 ( .A1(n9290), .A2(n9288), .ZN(n6890) );
  NAND2_X1 U9420 ( .A1(n9238), .A2(n9246), .ZN(n9216) );
  NAND2_X1 U9421 ( .A1(n6892), .A2(n6728), .ZN(n9409) );
  NAND2_X1 U9422 ( .A1(n9229), .A2(n6894), .ZN(n6892) );
  NAND3_X1 U9423 ( .A1(n12902), .A2(n12518), .A3(n7420), .ZN(n6899) );
  AND2_X2 U9424 ( .A1(n12512), .A2(n12511), .ZN(n12902) );
  NAND2_X1 U9425 ( .A1(n6901), .A2(n7016), .ZN(n6900) );
  NAND2_X1 U9426 ( .A1(n12048), .A2(n9615), .ZN(n6906) );
  XNOR2_X1 U9427 ( .A(n9610), .B(P2_DATAO_REG_24__SCAN_IN), .ZN(n12048) );
  NAND2_X1 U9428 ( .A1(n6916), .A2(n11858), .ZN(n6919) );
  INV_X1 U9429 ( .A(n6919), .ZN(n14569) );
  NAND4_X1 U9430 ( .A1(n6920), .A2(n11040), .A3(n11557), .A4(n7090), .ZN(
        n14610) );
  NAND2_X1 U9431 ( .A1(n6921), .A2(n6639), .ZN(n14403) );
  NAND2_X1 U9432 ( .A1(n7858), .A2(n6929), .ZN(n6927) );
  NAND2_X2 U9433 ( .A1(n6927), .A2(n6926), .ZN(n7917) );
  NAND3_X1 U9434 ( .A1(n6939), .A2(n6938), .A3(n6722), .ZN(n6937) );
  OR2_X2 U9435 ( .A1(n14097), .A2(n14098), .ZN(n6938) );
  NAND4_X1 U9436 ( .A1(n7717), .A2(n7358), .A3(P1_ADDR_REG_19__SCAN_IN), .A4(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n7356) );
  OAI21_X1 U9437 ( .B1(n6782), .B2(n6951), .A(n6948), .ZN(n8055) );
  OR2_X2 U9438 ( .A1(n14141), .A2(n6956), .ZN(n6954) );
  INV_X1 U9439 ( .A(n6953), .ZN(n6952) );
  OAI21_X1 U9440 ( .B1(n6956), .B2(n6958), .A(n6955), .ZN(n6953) );
  AOI21_X1 U9441 ( .B1(n14141), .B2(n6958), .A(n6956), .ZN(n14159) );
  INV_X1 U9442 ( .A(n14119), .ZN(n14122) );
  NAND2_X1 U9443 ( .A1(n6962), .A2(n6963), .ZN(n14119) );
  OR2_X1 U9444 ( .A1(n14114), .A2(n6964), .ZN(n6962) );
  NAND3_X1 U9445 ( .A1(n6966), .A2(n14079), .A3(n14080), .ZN(n14084) );
  NAND3_X1 U9446 ( .A1(n7125), .A2(n7126), .A3(n6718), .ZN(n6966) );
  NAND2_X1 U9447 ( .A1(n9266), .A2(n6862), .ZN(n9291) );
  NOR2_X1 U9448 ( .A1(n6984), .A2(n6988), .ZN(n6987) );
  NOR2_X1 U9449 ( .A1(n7994), .A2(n8254), .ZN(n6994) );
  NOR2_X1 U9450 ( .A1(n8254), .A2(n7993), .ZN(n7697) );
  NAND3_X1 U9451 ( .A1(n7996), .A2(n6994), .A3(n6993), .ZN(n8320) );
  NOR2_X1 U9452 ( .A1(n7994), .A2(n7695), .ZN(n7696) );
  NAND2_X2 U9453 ( .A1(n14765), .A2(n12173), .ZN(n9905) );
  INV_X1 U9454 ( .A(n7007), .ZN(n12957) );
  NAND2_X1 U9455 ( .A1(n9615), .A2(n9883), .ZN(n7009) );
  INV_X1 U9456 ( .A(n7010), .ZN(n9703) );
  NAND2_X1 U9457 ( .A1(n9708), .A2(n7019), .ZN(n7018) );
  NAND2_X1 U9458 ( .A1(n12078), .A2(n7036), .ZN(n7034) );
  NAND3_X1 U9459 ( .A1(n7047), .A2(n7046), .A3(n7045), .ZN(n7050) );
  NOR2_X1 U9460 ( .A1(n14789), .A2(n7648), .ZN(n7650) );
  NOR2_X1 U9461 ( .A1(n7648), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n7048) );
  INV_X1 U9462 ( .A(n14789), .ZN(n7049) );
  INV_X1 U9463 ( .A(n7050), .ZN(n15508) );
  NAND2_X1 U9464 ( .A1(n14959), .A2(n6668), .ZN(n7056) );
  NAND2_X1 U9465 ( .A1(n7056), .A2(n15305), .ZN(n7060) );
  AOI21_X1 U9466 ( .B1(n7663), .B2(P2_ADDR_REG_12__SCAN_IN), .A(n7058), .ZN(
        n7057) );
  INV_X1 U9467 ( .A(n7663), .ZN(n7059) );
  NAND2_X1 U9468 ( .A1(n14959), .A2(n7663), .ZN(n14962) );
  NAND2_X1 U9469 ( .A1(n9213), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n7077) );
  NAND2_X1 U9470 ( .A1(n14850), .A2(n6714), .ZN(n7080) );
  CLKBUF_X1 U9471 ( .A(n7080), .Z(n7078) );
  INV_X1 U9472 ( .A(n14598), .ZN(n7111) );
  NAND2_X1 U9473 ( .A1(n14565), .A2(n6632), .ZN(n7114) );
  OAI21_X1 U9474 ( .B1(n14425), .B2(n7118), .A(n7116), .ZN(n8294) );
  NAND2_X1 U9475 ( .A1(n14050), .A2(n7127), .ZN(n7125) );
  NAND2_X1 U9476 ( .A1(n7132), .A2(n7135), .ZN(n14047) );
  NAND3_X1 U9477 ( .A1(n14039), .A2(n7133), .A3(n14038), .ZN(n7132) );
  NAND2_X1 U9478 ( .A1(n7137), .A2(n7140), .ZN(n14023) );
  NAND3_X1 U9479 ( .A1(n14017), .A2(n7138), .A3(n14016), .ZN(n7137) );
  NAND2_X1 U9480 ( .A1(n7142), .A2(n7145), .ZN(n14012) );
  NAND3_X1 U9481 ( .A1(n14007), .A2(n7143), .A3(n14006), .ZN(n7142) );
  NAND2_X1 U9482 ( .A1(n7147), .A2(n7150), .ZN(n14034) );
  NAND3_X1 U9483 ( .A1(n14028), .A2(n7148), .A3(n14027), .ZN(n7147) );
  INV_X2 U9484 ( .A(n13973), .ZN(n14091) );
  OAI22_X2 U9485 ( .A1(n13971), .A2(n13972), .B1(n13970), .B2(n7152), .ZN(
        n13980) );
  MUX2_X1 U9486 ( .A(n13969), .B(n14231), .S(n13973), .Z(n7152) );
  NAND4_X1 U9487 ( .A1(n8037), .A2(n7995), .A3(n7996), .A4(n7154), .ZN(n8056)
         );
  OAI22_X1 U9488 ( .A1(n14093), .A2(n7156), .B1(n7155), .B2(n14094), .ZN(
        n14097) );
  OAI22_X1 U9489 ( .A1(n14110), .A2(n7158), .B1(n7157), .B2(n14111), .ZN(
        n14114) );
  OAI22_X2 U9490 ( .A1(n9642), .A2(n9641), .B1(P2_DATAO_REG_26__SCAN_IN), .B2(
        n13800), .ZN(n9653) );
  AND3_X2 U9491 ( .A1(n7167), .A2(n7166), .A3(n7161), .ZN(n12719) );
  NAND3_X1 U9492 ( .A1(n12710), .A2(n7165), .A3(n12708), .ZN(n7164) );
  OR2_X2 U9493 ( .A1(n12704), .A2(n12702), .ZN(n7167) );
  NAND2_X1 U9494 ( .A1(n9429), .A2(n7171), .ZN(n7168) );
  NAND2_X1 U9495 ( .A1(n7184), .A2(n7186), .ZN(n9227) );
  NAND2_X1 U9496 ( .A1(n9327), .A2(n9225), .ZN(n7184) );
  NAND2_X1 U9499 ( .A1(n12171), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n7198) );
  NAND2_X1 U9500 ( .A1(n9468), .A2(n9467), .ZN(n9469) );
  NAND2_X1 U9501 ( .A1(n7799), .A2(n7199), .ZN(n11039) );
  NAND2_X1 U9502 ( .A1(n10744), .A2(n7201), .ZN(n7200) );
  NAND2_X1 U9503 ( .A1(n10744), .A2(n7776), .ZN(n10972) );
  NAND2_X1 U9504 ( .A1(n11039), .A2(n14174), .ZN(n7820) );
  NAND2_X1 U9505 ( .A1(n7214), .A2(n7215), .ZN(n11855) );
  NAND2_X1 U9506 ( .A1(n11050), .A2(n11051), .ZN(n11052) );
  NAND2_X1 U9507 ( .A1(n14464), .A2(n6711), .ZN(n7230) );
  INV_X1 U9508 ( .A(n7714), .ZN(n7713) );
  NAND3_X1 U9509 ( .A1(n7697), .A2(n7696), .A3(n7233), .ZN(n7714) );
  INV_X1 U9510 ( .A(n7235), .ZN(n7234) );
  NAND2_X1 U9511 ( .A1(n11254), .A2(n7236), .ZN(n11452) );
  INV_X1 U9512 ( .A(n7242), .ZN(n7241) );
  AND2_X1 U9513 ( .A1(n8359), .A2(n8358), .ZN(n7573) );
  NAND4_X2 U9514 ( .A1(n8354), .A2(n7262), .A3(n8477), .A4(n8359), .ZN(n8379)
         );
  AND2_X2 U9515 ( .A1(n8354), .A2(n8477), .ZN(n8609) );
  NAND2_X1 U9516 ( .A1(n10292), .A2(n6725), .ZN(n8387) );
  NAND2_X1 U9517 ( .A1(n8778), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8375) );
  NOR2_X2 U9518 ( .A1(n9291), .A2(n7275), .ZN(n9341) );
  NAND4_X1 U9519 ( .A1(n9190), .A2(n9189), .A3(n9188), .A4(n9309), .ZN(n7275)
         );
  AOI21_X1 U9520 ( .B1(n7280), .B2(n10697), .A(n12494), .ZN(n10698) );
  NAND2_X1 U9521 ( .A1(n12463), .A2(n7283), .ZN(n7282) );
  OAI21_X1 U9522 ( .B1(n12449), .B2(n7308), .A(n7305), .ZN(n12391) );
  NAND2_X1 U9523 ( .A1(n12449), .A2(n6661), .ZN(n7304) );
  OAI21_X1 U9524 ( .B1(n12449), .B2(n12365), .A(n12364), .ZN(n12427) );
  NAND2_X1 U9525 ( .A1(n12056), .A2(n7314), .ZN(n7313) );
  NAND3_X1 U9526 ( .A1(n7313), .A2(n12186), .A3(n7320), .ZN(n13858) );
  NAND2_X1 U9527 ( .A1(n13910), .A2(n6634), .ZN(n7326) );
  AND2_X1 U9528 ( .A1(n14231), .A2(n14583), .ZN(n15095) );
  INV_X1 U9529 ( .A(n14231), .ZN(n7330) );
  NAND2_X1 U9530 ( .A1(n13863), .A2(n7334), .ZN(n7332) );
  NAND2_X1 U9531 ( .A1(n13863), .A2(n13864), .ZN(n7333) );
  NAND2_X2 U9532 ( .A1(n13895), .A2(n13894), .ZN(n13893) );
  OAI21_X1 U9533 ( .B1(n13857), .B2(n7350), .A(n7349), .ZN(n12211) );
  NAND2_X1 U9534 ( .A1(n7713), .A2(n7715), .ZN(n7703) );
  NAND2_X1 U9535 ( .A1(n7713), .A2(n7354), .ZN(n14755) );
  INV_X1 U9536 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n13434) );
  NAND2_X1 U9537 ( .A1(n7822), .A2(n7363), .ZN(n7362) );
  INV_X1 U9538 ( .A(n8143), .ZN(n7366) );
  OAI211_X2 U9539 ( .C1(n8675), .C2(n7367), .A(n8158), .B(n7365), .ZN(n8173)
         );
  XNOR2_X2 U9540 ( .A(n8142), .B(SI_22_), .ZN(n8675) );
  NAND2_X1 U9541 ( .A1(n8073), .A2(n8072), .ZN(n8076) );
  NAND2_X1 U9542 ( .A1(n7383), .A2(n7384), .ZN(n9084) );
  NAND2_X1 U9543 ( .A1(n9077), .A2(n9076), .ZN(n7390) );
  NAND2_X1 U9544 ( .A1(n7973), .A2(n10197), .ZN(n7391) );
  NAND2_X1 U9545 ( .A1(n8099), .A2(n7392), .ZN(n8133) );
  NAND2_X1 U9546 ( .A1(n7574), .A2(n7577), .ZN(n7394) );
  OAI21_X1 U9547 ( .B1(n15447), .B2(n10779), .A(n7402), .ZN(n11386) );
  NAND3_X1 U9548 ( .A1(n7422), .A2(n7457), .A3(n9211), .ZN(n7421) );
  NAND2_X2 U9549 ( .A1(n7427), .A2(n7430), .ZN(n8868) );
  OAI21_X2 U9550 ( .B1(n9795), .B2(n6621), .A(n7428), .ZN(n10597) );
  AOI21_X1 U9551 ( .B1(n7429), .B2(n13658), .A(n6674), .ZN(n7428) );
  INV_X1 U9552 ( .A(n8818), .ZN(n7429) );
  NAND2_X1 U9553 ( .A1(n9795), .A2(n8818), .ZN(n13659) );
  NAND3_X1 U9554 ( .A1(n8609), .A2(n7573), .A3(n7551), .ZN(n7430) );
  NAND2_X1 U9555 ( .A1(n7433), .A2(n7431), .ZN(n8860) );
  NAND2_X1 U9556 ( .A1(n8857), .A2(n7434), .ZN(n7433) );
  NAND2_X1 U9557 ( .A1(n8850), .A2(n7438), .ZN(n7441) );
  NAND2_X1 U9558 ( .A1(n11749), .A2(n7451), .ZN(n7449) );
  NAND2_X1 U9559 ( .A1(n13619), .A2(n7454), .ZN(n7453) );
  NAND2_X1 U9560 ( .A1(n9466), .A2(n6633), .ZN(n7460) );
  NAND2_X1 U9561 ( .A1(n12869), .A2(n7468), .ZN(n12861) );
  NAND2_X1 U9562 ( .A1(n11404), .A2(n7475), .ZN(n7474) );
  NAND2_X1 U9563 ( .A1(n7474), .A2(n7471), .ZN(n11732) );
  NAND2_X1 U9564 ( .A1(n11404), .A2(n9349), .ZN(n11620) );
  INV_X1 U9565 ( .A(n7474), .ZN(n11619) );
  INV_X1 U9566 ( .A(n9349), .ZN(n7476) );
  NAND2_X1 U9567 ( .A1(n12004), .A2(n7480), .ZN(n7477) );
  NAND2_X1 U9568 ( .A1(n7477), .A2(n7478), .ZN(n12124) );
  NAND2_X1 U9569 ( .A1(n7489), .A2(n7488), .ZN(n9599) );
  NAND2_X1 U9570 ( .A1(n7489), .A2(n9569), .ZN(n12933) );
  NAND2_X1 U9571 ( .A1(n9697), .A2(n13032), .ZN(n7492) );
  OAI21_X1 U9572 ( .B1(n12901), .B2(n7505), .A(n7503), .ZN(n12871) );
  NAND2_X1 U9573 ( .A1(n9210), .A2(n7511), .ZN(n9196) );
  AND2_X2 U9574 ( .A1(n8609), .A2(n7512), .ZN(n8785) );
  INV_X1 U9575 ( .A(n10837), .ZN(n7516) );
  NAND2_X1 U9576 ( .A1(n8802), .A2(n6719), .ZN(n7518) );
  NAND2_X1 U9577 ( .A1(n8802), .A2(n8786), .ZN(n8806) );
  AOI21_X2 U9578 ( .B1(n7518), .B2(n7519), .A(n8799), .ZN(n8813) );
  NAND2_X1 U9579 ( .A1(n13333), .A2(n7522), .ZN(n13253) );
  OAI21_X2 U9580 ( .B1(n11771), .B2(n7533), .A(n7531), .ZN(n15186) );
  OAI21_X1 U9581 ( .B1(n9060), .B2(n7544), .A(n7543), .ZN(n9064) );
  INV_X1 U9582 ( .A(n8379), .ZN(n8362) );
  NAND3_X1 U9583 ( .A1(n7564), .A2(n8948), .A3(n6723), .ZN(n7552) );
  NAND3_X1 U9584 ( .A1(n7572), .A2(n7556), .A3(n7555), .ZN(n9018) );
  INV_X1 U9585 ( .A(n9026), .ZN(n7559) );
  AND4_X2 U9586 ( .A1(n7745), .A2(n7744), .A3(n7743), .A4(n7742), .ZN(n13976)
         );
  NAND2_X1 U9587 ( .A1(n9557), .A2(n9556), .ZN(n9570) );
  NOR2_X2 U9588 ( .A1(n14233), .A2(n10389), .ZN(n13966) );
  NAND2_X1 U9589 ( .A1(n14005), .A2(n14004), .ZN(n14006) );
  NAND2_X1 U9590 ( .A1(n14122), .A2(n14121), .ZN(n14123) );
  OAI21_X1 U9591 ( .B1(n14233), .B2(n10417), .A(n9941), .ZN(n15098) );
  XNOR2_X1 U9592 ( .A(n12314), .B(n9673), .ZN(n13156) );
  NAND2_X1 U9593 ( .A1(n11470), .A2(n11322), .ZN(n15486) );
  INV_X1 U9594 ( .A(n8882), .ZN(n8883) );
  NAND2_X2 U9595 ( .A1(n8326), .A2(n9815), .ZN(n10394) );
  NAND2_X1 U9596 ( .A1(n8322), .A2(n9815), .ZN(n9813) );
  NAND2_X4 U9597 ( .A1(n7707), .A2(n7706), .ZN(n8244) );
  NAND2_X1 U9598 ( .A1(n7992), .A2(n7991), .ZN(n8017) );
  NAND2_X1 U9599 ( .A1(n10394), .A2(n9825), .ZN(n10406) );
  NOR2_X1 U9600 ( .A1(n10394), .A2(n9814), .ZN(n14232) );
  AND2_X1 U9601 ( .A1(n8327), .A2(n10394), .ZN(n10414) );
  NAND2_X1 U9602 ( .A1(n8085), .A2(n8084), .ZN(n8087) );
  INV_X1 U9603 ( .A(n8085), .ZN(n8057) );
  NAND2_X1 U9604 ( .A1(n8318), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8313) );
  INV_X1 U9605 ( .A(n7994), .ZN(n7995) );
  NAND4_X4 U9606 ( .A1(n7737), .A2(n7736), .A3(n7735), .A4(n7734), .ZN(n14233)
         );
  NAND4_X2 U9607 ( .A1(n8374), .A2(n8373), .A3(n8372), .A4(n8371), .ZN(n13383)
         );
  NAND2_X1 U9608 ( .A1(n8389), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n8372) );
  OAI21_X1 U9609 ( .B1(n13678), .B2(n6620), .A(n8881), .ZN(n8882) );
  INV_X1 U9610 ( .A(n13383), .ZN(n8388) );
  NAND2_X1 U9611 ( .A1(n11387), .A2(n9296), .ZN(n11312) );
  OAI21_X1 U9612 ( .B1(n8802), .B2(n8803), .A(P2_IR_REG_20__SCAN_IN), .ZN(
        n8805) );
  CLKBUF_X1 U9613 ( .A(n13253), .Z(n13227) );
  OR2_X2 U9614 ( .A1(n6617), .A2(n7708), .ZN(n7709) );
  OR2_X1 U9615 ( .A1(n12329), .A2(n9269), .ZN(n11251) );
  INV_X1 U9616 ( .A(n8877), .ZN(n9110) );
  INV_X2 U9617 ( .A(n8192), .ZN(n9213) );
  NAND2_X1 U9618 ( .A1(n9141), .A2(n6653), .ZN(n9094) );
  OR2_X1 U9619 ( .A1(n9056), .A2(n9055), .ZN(n9060) );
  AOI211_X1 U9620 ( .C1(n9169), .C2(n10916), .A(n9168), .B(n9167), .ZN(n9171)
         );
  OR2_X1 U9621 ( .A1(n12332), .A2(n13092), .ZN(n7562) );
  OR2_X1 U9622 ( .A1(n12332), .A2(n13144), .ZN(n7563) );
  NAND2_X1 U9623 ( .A1(n9445), .A2(n9444), .ZN(n12150) );
  OR2_X1 U9624 ( .A1(n8947), .A2(n8946), .ZN(n7564) );
  INV_X1 U9625 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n7718) );
  AND2_X1 U9626 ( .A1(n10709), .A2(n15458), .ZN(n7565) );
  AND2_X1 U9627 ( .A1(n7576), .A2(n8347), .ZN(n7566) );
  OR2_X1 U9628 ( .A1(n12006), .A2(n12574), .ZN(n7568) );
  INV_X1 U9629 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n8310) );
  AND2_X1 U9630 ( .A1(n11794), .A2(n11689), .ZN(n7569) );
  AND2_X1 U9631 ( .A1(n12299), .A2(n12298), .ZN(n7570) );
  OR2_X1 U9632 ( .A1(n8984), .A2(n8983), .ZN(n7571) );
  AND2_X1 U9633 ( .A1(n9016), .A2(n9007), .ZN(n7572) );
  INV_X1 U9634 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n11431) );
  INV_X1 U9635 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n8468) );
  INV_X1 U9636 ( .A(n14686), .ZN(n8887) );
  INV_X1 U9637 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n11433) );
  INV_X1 U9638 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n7923) );
  OR2_X1 U9639 ( .A1(n8884), .A2(n10404), .ZN(n15183) );
  OR2_X1 U9640 ( .A1(n8884), .A2(n9780), .ZN(n15172) );
  OR2_X1 U9641 ( .A1(n8128), .A2(SI_20_), .ZN(n7574) );
  OR2_X1 U9642 ( .A1(n13679), .A2(n13592), .ZN(n7575) );
  OR2_X1 U9643 ( .A1(n14365), .A2(n14748), .ZN(n7576) );
  INV_X1 U9644 ( .A(n13651), .ZN(n13604) );
  OR2_X1 U9645 ( .A1(n8130), .A2(SI_21_), .ZN(n7577) );
  INV_X1 U9646 ( .A(n13479), .ZN(n13495) );
  INV_X1 U9647 ( .A(n14167), .ZN(n14931) );
  NOR2_X1 U9648 ( .A1(n9354), .A2(n9353), .ZN(n7578) );
  NAND2_X1 U9649 ( .A1(n9637), .A2(n9636), .ZN(n12904) );
  OR2_X1 U9650 ( .A1(n13134), .A2(n12954), .ZN(n7579) );
  OR2_X1 U9651 ( .A1(n12510), .A2(n12599), .ZN(n7580) );
  INV_X1 U9652 ( .A(n12690), .ZN(n9517) );
  OR2_X1 U9653 ( .A1(n10727), .A2(n8893), .ZN(n8895) );
  NAND2_X1 U9654 ( .A1(n15354), .A2(n8909), .ZN(n8907) );
  NAND2_X1 U9655 ( .A1(n8908), .A2(n8907), .ZN(n8916) );
  AOI21_X1 U9656 ( .B1(n8935), .B2(n8934), .A(n8933), .ZN(n8936) );
  INV_X1 U9657 ( .A(n8954), .ZN(n8955) );
  AOI21_X1 U9658 ( .B1(n8960), .B2(n8959), .A(n8958), .ZN(n8962) );
  AOI21_X1 U9659 ( .B1(n9016), .B2(n9015), .A(n9014), .ZN(n9017) );
  NAND2_X1 U9660 ( .A1(n9039), .A2(n9038), .ZN(n9043) );
  AOI21_X1 U9661 ( .B1(n9070), .B2(n9069), .A(n9068), .ZN(n9071) );
  NOR2_X1 U9662 ( .A1(n12888), .A2(n12693), .ZN(n12694) );
  NAND2_X1 U9663 ( .A1(n14818), .A2(n12711), .ZN(n12712) );
  INV_X1 U9664 ( .A(n12877), .ZN(n9667) );
  INV_X1 U9665 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n9181) );
  INV_X1 U9666 ( .A(P3_IR_REG_8__SCAN_IN), .ZN(n9191) );
  NAND2_X1 U9667 ( .A1(n12398), .A2(n9667), .ZN(n9668) );
  NAND2_X1 U9668 ( .A1(n9638), .A2(n12876), .ZN(n9639) );
  AND2_X1 U9669 ( .A1(n9791), .A2(n8877), .ZN(n8814) );
  INV_X1 U9670 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n8608) );
  INV_X1 U9671 ( .A(n10394), .ZN(n10395) );
  INV_X1 U9672 ( .A(n8168), .ZN(n8169) );
  INV_X1 U9673 ( .A(P3_REG3_REG_14__SCAN_IN), .ZN(n9437) );
  INV_X1 U9674 ( .A(P3_REG3_REG_12__SCAN_IN), .ZN(n11656) );
  INV_X1 U9675 ( .A(P3_REG3_REG_18__SCAN_IN), .ZN(n9510) );
  OR2_X1 U9676 ( .A1(n9398), .A2(n9397), .ZN(n9423) );
  NAND2_X1 U9677 ( .A1(n11016), .A2(n11366), .ZN(n9255) );
  INV_X1 U9678 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n9669) );
  NAND2_X1 U9679 ( .A1(n13237), .A2(n13236), .ZN(n13207) );
  AND2_X1 U9680 ( .A1(n9122), .A2(n9121), .ZN(n9123) );
  AND2_X1 U9681 ( .A1(n8652), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n8665) );
  INV_X1 U9682 ( .A(n13694), .ZN(n8876) );
  INV_X1 U9683 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n8348) );
  AOI21_X1 U9684 ( .B1(n10428), .B2(n10417), .A(n10396), .ZN(n10397) );
  INV_X1 U9685 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n8003) );
  INV_X1 U9686 ( .A(n14946), .ZN(n8300) );
  INV_X1 U9687 ( .A(P1_B_REG_SCAN_IN), .ZN(n10211) );
  AND2_X1 U9688 ( .A1(n7581), .A2(P3_ADDR_REG_2__SCAN_IN), .ZN(n7582) );
  INV_X1 U9689 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n9200) );
  INV_X1 U9690 ( .A(P3_REG3_REG_8__SCAN_IN), .ZN(n9351) );
  INV_X1 U9691 ( .A(n12702), .ZN(n9763) );
  AND2_X1 U9692 ( .A1(n9631), .A2(n9630), .ZN(n9647) );
  NOR2_X1 U9693 ( .A1(n9546), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n9562) );
  NAND2_X1 U9694 ( .A1(n9511), .A2(n9510), .ZN(n9533) );
  OR2_X1 U9695 ( .A1(n9458), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n9475) );
  INV_X1 U9696 ( .A(n11322), .ZN(n12528) );
  OR2_X1 U9697 ( .A1(n12653), .A2(n9763), .ZN(n11359) );
  NAND2_X1 U9698 ( .A1(n10778), .A2(n9282), .ZN(n11389) );
  INV_X1 U9699 ( .A(P3_IR_REG_22__SCAN_IN), .ZN(n9682) );
  INV_X1 U9700 ( .A(n11348), .ZN(n11346) );
  AND2_X1 U9701 ( .A1(n8665), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n8678) );
  NOR2_X1 U9702 ( .A1(n8469), .A2(n8468), .ZN(n8485) );
  OR2_X1 U9703 ( .A1(n15293), .A2(n15294), .ZN(n15290) );
  INV_X1 U9704 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n11503) );
  OR2_X1 U9705 ( .A1(n8746), .A2(n13262), .ZN(n8757) );
  OR2_X1 U9706 ( .A1(n8497), .A2(n8496), .ZN(n8511) );
  INV_X1 U9707 ( .A(n13303), .ZN(n13337) );
  INV_X1 U9708 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n8786) );
  OR2_X1 U9709 ( .A1(n8506), .A2(P2_IR_REG_9__SCAN_IN), .ZN(n8593) );
  INV_X1 U9710 ( .A(n12208), .ZN(n10430) );
  AND2_X1 U9711 ( .A1(n11988), .A2(n11987), .ZN(n11989) );
  INV_X1 U9712 ( .A(n8197), .ZN(n8195) );
  INV_X1 U9713 ( .A(n14523), .ZN(n8282) );
  AND2_X1 U9714 ( .A1(n8022), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n8042) );
  INV_X1 U9715 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n8088) );
  INV_X1 U9716 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n9448) );
  INV_X1 U9717 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n8018) );
  INV_X1 U9718 ( .A(P3_ADDR_REG_6__SCAN_IN), .ZN(n7593) );
  INV_X1 U9719 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n7666) );
  NAND2_X1 U9720 ( .A1(n9354), .A2(n9200), .ZN(n9366) );
  AND2_X1 U9721 ( .A1(n9352), .A2(n9351), .ZN(n9354) );
  INV_X1 U9722 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n9297) );
  INV_X1 U9723 ( .A(n12500), .ZN(n12485) );
  INV_X1 U9724 ( .A(n12904), .ZN(n12876) );
  AND2_X1 U9725 ( .A1(n12647), .A2(n9763), .ZN(n10717) );
  AND2_X1 U9726 ( .A1(n9647), .A2(n12369), .ZN(n9659) );
  OR2_X1 U9727 ( .A1(n10535), .A2(n12720), .ZN(n12841) );
  INV_X1 U9728 ( .A(n12940), .ZN(n12967) );
  AND2_X1 U9729 ( .A1(n12621), .A2(n12620), .ZN(n12995) );
  AND2_X1 U9730 ( .A1(n12579), .A2(n12585), .ZN(n12682) );
  OR2_X1 U9731 ( .A1(n15454), .A2(n15460), .ZN(n15437) );
  AND2_X1 U9732 ( .A1(n12587), .A2(n12586), .ZN(n12681) );
  INV_X1 U9733 ( .A(n12734), .ZN(n11871) );
  NAND2_X1 U9734 ( .A1(n10707), .A2(n12647), .ZN(n15452) );
  INV_X1 U9735 ( .A(n13029), .ZN(n15450) );
  INV_X1 U9736 ( .A(n13032), .ZN(n15457) );
  AND2_X1 U9737 ( .A1(n11242), .A2(n12847), .ZN(n12705) );
  NAND2_X1 U9738 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(n11431), .ZN(n9521) );
  NAND2_X1 U9739 ( .A1(n9227), .A2(n9226), .ZN(n9361) );
  OR2_X1 U9740 ( .A1(n8628), .A2(n8627), .ZN(n8639) );
  INV_X1 U9741 ( .A(n15348), .ZN(n10619) );
  XNOR2_X1 U9742 ( .A(n13180), .B(n13179), .ZN(n13351) );
  AND2_X1 U9743 ( .A1(n8678), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n8688) );
  OR2_X1 U9744 ( .A1(n15273), .A2(n15272), .ZN(n15275) );
  INV_X1 U9745 ( .A(n11880), .ZN(n11883) );
  AND4_X1 U9746 ( .A1(n8752), .A2(n8751), .A3(n8750), .A4(n8749), .ZN(n13254)
         );
  INV_X1 U9747 ( .A(n9152), .ZN(n11811) );
  NAND2_X1 U9748 ( .A1(n13384), .A2(n10639), .ZN(n9142) );
  XNOR2_X1 U9749 ( .A(n8864), .B(n9163), .ZN(n8875) );
  AND2_X1 U9750 ( .A1(n8865), .A2(n9134), .ZN(n13623) );
  INV_X1 U9751 ( .A(n9173), .ZN(n10623) );
  INV_X1 U9752 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n8363) );
  INV_X1 U9753 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n8795) );
  NAND2_X1 U9754 ( .A1(n8042), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n8063) );
  AND2_X1 U9755 ( .A1(n8135), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n8147) );
  NAND2_X1 U9756 ( .A1(n14377), .A2(n14921), .ZN(n14378) );
  INV_X1 U9757 ( .A(n14928), .ZN(n10409) );
  OR2_X1 U9758 ( .A1(n14915), .A2(n14917), .ZN(n10412) );
  INV_X1 U9759 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n8252) );
  INV_X1 U9760 ( .A(n7975), .ZN(n7974) );
  NOR2_X1 U9761 ( .A1(n7887), .A2(P1_IR_REG_9__SCAN_IN), .ZN(n7919) );
  NAND2_X1 U9762 ( .A1(n7780), .A2(n7766), .ZN(n7777) );
  NOR2_X1 U9763 ( .A1(n9333), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n9352) );
  INV_X1 U9764 ( .A(n12729), .ZN(n12955) );
  AND2_X1 U9765 ( .A1(n9483), .A2(n9482), .ZN(n9511) );
  NOR2_X2 U9766 ( .A1(n12741), .A2(n11527), .ZN(n12529) );
  NAND2_X1 U9767 ( .A1(n10677), .A2(n10676), .ZN(n12486) );
  INV_X1 U9768 ( .A(n12489), .ZN(n12506) );
  INV_X1 U9769 ( .A(n9269), .ZN(n9665) );
  AND4_X1 U9770 ( .A1(n9567), .A2(n9566), .A3(n9565), .A4(n9564), .ZN(n12954)
         );
  AND4_X1 U9771 ( .A1(n9488), .A2(n9487), .A3(n9486), .A4(n9485), .ZN(n12478)
         );
  INV_X1 U9772 ( .A(n11661), .ZN(n15416) );
  INV_X1 U9773 ( .A(n12841), .ZN(n15426) );
  AND2_X1 U9774 ( .A1(n10706), .A2(n12647), .ZN(n13029) );
  AND2_X1 U9775 ( .A1(n15464), .A2(n15437), .ZN(n13039) );
  AND2_X1 U9776 ( .A1(n9762), .A2(n9761), .ZN(n11365) );
  OR2_X1 U9777 ( .A1(n15454), .A2(n15475), .ZN(n15477) );
  AND2_X1 U9778 ( .A1(n11470), .A2(n12705), .ZN(n15475) );
  NAND2_X1 U9779 ( .A1(n9733), .A2(n9732), .ZN(n10680) );
  INV_X1 U9780 ( .A(P3_IR_REG_21__SCAN_IN), .ZN(n9685) );
  INV_X1 U9781 ( .A(n13331), .ZN(n15195) );
  INV_X1 U9782 ( .A(n13254), .ZN(n11029) );
  AND2_X1 U9783 ( .A1(n15236), .A2(n10307), .ZN(n15307) );
  OR2_X1 U9784 ( .A1(n15300), .A2(n15299), .ZN(n15301) );
  INV_X1 U9785 ( .A(n15318), .ZN(n15224) );
  AND2_X1 U9786 ( .A1(n15236), .A2(n10296), .ZN(n15318) );
  INV_X1 U9787 ( .A(n9149), .ZN(n11559) );
  INV_X1 U9788 ( .A(n13623), .ZN(n13661) );
  NOR2_X1 U9789 ( .A1(n10632), .A2(n10545), .ZN(n10546) );
  INV_X1 U9790 ( .A(n13734), .ZN(n15381) );
  INV_X1 U9791 ( .A(n10632), .ZN(n10604) );
  AND2_X1 U9792 ( .A1(n10630), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9771) );
  AND2_X1 U9793 ( .A1(n7088), .A2(P2_U3088), .ZN(n13792) );
  INV_X1 U9794 ( .A(n13916), .ZN(n13934) );
  OR3_X1 U9795 ( .A1(n7925), .A2(n7924), .A3(n7923), .ZN(n7945) );
  AND2_X1 U9796 ( .A1(n14202), .A2(n14201), .ZN(n14203) );
  AND2_X1 U9797 ( .A1(n8110), .A2(n8109), .ZN(n14085) );
  AND4_X1 U9798 ( .A1(n8013), .A2(n8012), .A3(n8011), .A4(n8010), .ZN(n14920)
         );
  OR2_X1 U9799 ( .A1(n14983), .A2(n10441), .ZN(n15037) );
  INV_X1 U9800 ( .A(n15060), .ZN(n15012) );
  INV_X1 U9801 ( .A(n15037), .ZN(n15067) );
  XNOR2_X1 U9802 ( .A(n8250), .B(n8296), .ZN(n14357) );
  INV_X1 U9803 ( .A(n14919), .ZN(n14583) );
  INV_X1 U9805 ( .A(n15099), .ZN(n14609) );
  NAND2_X2 U9807 ( .A1(n9782), .A2(n9812), .ZN(n14602) );
  NAND2_X1 U9808 ( .A1(n8343), .A2(n9824), .ZN(n10404) );
  INV_X1 U9809 ( .A(n15170), .ZN(n14949) );
  INV_X1 U9810 ( .A(n15129), .ZN(n15162) );
  NAND2_X1 U9811 ( .A1(n15129), .A2(n15159), .ZN(n15170) );
  INV_X1 U9812 ( .A(n9825), .ZN(n9814) );
  XNOR2_X1 U9813 ( .A(n8315), .B(P1_IR_REG_24__SCAN_IN), .ZN(n8324) );
  INV_X1 U9814 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n8084) );
  INV_X1 U9815 ( .A(n7660), .ZN(n7661) );
  NAND2_X1 U9816 ( .A1(n9747), .A2(n9746), .ZN(n10671) );
  INV_X1 U9817 ( .A(n12486), .ZN(n12503) );
  NAND2_X1 U9818 ( .A1(n10696), .A2(n10702), .ZN(n12494) );
  AOI21_X1 U9819 ( .B1(n12864), .B2(n9665), .A(n9664), .ZN(n12877) );
  INV_X1 U9820 ( .A(n12966), .ZN(n12989) );
  INV_X1 U9821 ( .A(n15451), .ZN(n12739) );
  INV_X1 U9822 ( .A(n15417), .ZN(n11925) );
  OR2_X1 U9823 ( .A1(n10535), .A2(n10534), .ZN(n15401) );
  INV_X1 U9824 ( .A(n13039), .ZN(n12088) );
  NAND2_X1 U9825 ( .A1(n15498), .A2(n15479), .ZN(n13092) );
  INV_X1 U9826 ( .A(n11874), .ZN(n12574) );
  AND2_X1 U9827 ( .A1(n9757), .A2(n9756), .ZN(n15491) );
  INV_X1 U9828 ( .A(n13151), .ZN(n13149) );
  INV_X1 U9829 ( .A(SI_16_), .ZN(n10425) );
  INV_X1 U9830 ( .A(n11901), .ZN(n11891) );
  OR3_X1 U9831 ( .A1(n12136), .A2(n13803), .A3(n13801), .ZN(n10631) );
  NAND2_X1 U9832 ( .A1(n10737), .A2(P2_STATE_REG_SCAN_IN), .ZN(n15198) );
  INV_X1 U9833 ( .A(n15190), .ZN(n13347) );
  INV_X1 U9834 ( .A(n15314), .ZN(n15298) );
  OR2_X1 U9835 ( .A1(n6620), .A2(n10621), .ZN(n15330) );
  AND2_X2 U9836 ( .A1(n10620), .A2(n10546), .ZN(n15392) );
  INV_X1 U9837 ( .A(n13445), .ZN(n13757) );
  INV_X1 U9838 ( .A(n13524), .ZN(n13770) );
  NAND2_X1 U9839 ( .A1(n15383), .A2(n15355), .ZN(n13783) );
  AND2_X2 U9840 ( .A1(n10605), .A2(n10604), .ZN(n15383) );
  NOR2_X1 U9841 ( .A1(n15346), .A2(n15337), .ZN(n15342) );
  INV_X1 U9842 ( .A(n15342), .ZN(n15343) );
  INV_X1 U9843 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n12171) );
  INV_X1 U9844 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n11168) );
  INV_X1 U9845 ( .A(n14909), .ZN(n13922) );
  NAND2_X1 U9846 ( .A1(n10410), .A2(n10408), .ZN(n14904) );
  INV_X1 U9847 ( .A(n14981), .ZN(n15070) );
  INV_X1 U9848 ( .A(n14561), .ZN(n15100) );
  NAND2_X1 U9849 ( .A1(n14539), .A2(n10973), .ZN(n15099) );
  AOI21_X1 U9850 ( .B1(n14139), .B2(n8887), .A(n8886), .ZN(n8888) );
  INV_X2 U9851 ( .A(n15183), .ZN(n15185) );
  INV_X1 U9852 ( .A(n14481), .ZN(n14738) );
  INV_X2 U9853 ( .A(n15172), .ZN(n15174) );
  AND2_X1 U9854 ( .A1(n10413), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9825) );
  INV_X1 U9855 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n14773) );
  INV_X1 U9856 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n10553) );
  XNOR2_X1 U9857 ( .A(n7683), .B(n7682), .ZN(n7684) );
  NOR2_X2 U9858 ( .A1(n10671), .A2(n13149), .ZN(P3_U3897) );
  NAND2_X1 U9859 ( .A1(n7575), .A2(n8883), .ZN(P2_U3236) );
  CLKBUF_X2 U9860 ( .A(n14232), .Z(P1_U4016) );
  OAI21_X1 U9861 ( .B1(n8889), .B2(n15183), .A(n8888), .ZN(P1_U3557) );
  OAI21_X1 U9862 ( .B1(n8889), .B2(n15172), .A(n7566), .ZN(P1_U3525) );
  INV_X1 U9863 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n15041) );
  INV_X1 U9864 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n15023) );
  XNOR2_X1 U9865 ( .A(P1_ADDR_REG_15__SCAN_IN), .B(P3_ADDR_REG_15__SCAN_IN), 
        .ZN(n7665) );
  INV_X1 U9866 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n15010) );
  XNOR2_X1 U9867 ( .A(P1_ADDR_REG_14__SCAN_IN), .B(P3_ADDR_REG_14__SCAN_IN), 
        .ZN(n7613) );
  INV_X1 U9868 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n14996) );
  INV_X1 U9869 ( .A(P3_ADDR_REG_12__SCAN_IN), .ZN(n7607) );
  INV_X1 U9870 ( .A(P3_ADDR_REG_11__SCAN_IN), .ZN(n7605) );
  INV_X1 U9871 ( .A(P3_ADDR_REG_10__SCAN_IN), .ZN(n7622) );
  INV_X1 U9872 ( .A(P3_ADDR_REG_9__SCAN_IN), .ZN(n7601) );
  INV_X1 U9873 ( .A(P3_ADDR_REG_8__SCAN_IN), .ZN(n7599) );
  INV_X2 U9874 ( .A(P3_ADDR_REG_0__SCAN_IN), .ZN(n10610) );
  XOR2_X1 U9875 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(P3_ADDR_REG_2__SCAN_IN), .Z(
        n7629) );
  NOR2_X1 U9876 ( .A1(n7630), .A2(n7629), .ZN(n7583) );
  NOR2_X1 U9877 ( .A1(n7586), .A2(n15414), .ZN(n7588) );
  NOR2_X1 U9878 ( .A1(n7589), .A2(n7590), .ZN(n7592) );
  XNOR2_X1 U9879 ( .A(n7590), .B(n7589), .ZN(n7639) );
  INV_X1 U9880 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n9912) );
  NOR2_X1 U9881 ( .A1(P3_ADDR_REG_6__SCAN_IN), .A2(n9912), .ZN(n7594) );
  NOR2_X1 U9882 ( .A1(P3_ADDR_REG_7__SCAN_IN), .A2(n7595), .ZN(n7597) );
  XNOR2_X1 U9883 ( .A(P3_ADDR_REG_7__SCAN_IN), .B(n7595), .ZN(n7626) );
  XOR2_X1 U9884 ( .A(P3_ADDR_REG_8__SCAN_IN), .B(P1_ADDR_REG_8__SCAN_IN), .Z(
        n7651) );
  INV_X1 U9885 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n14292) );
  XOR2_X1 U9886 ( .A(P3_ADDR_REG_9__SCAN_IN), .B(n14292), .Z(n7624) );
  NAND2_X1 U9887 ( .A1(n7625), .A2(n7624), .ZN(n7600) );
  NAND2_X1 U9888 ( .A1(n7621), .A2(n7620), .ZN(n7603) );
  NOR2_X1 U9889 ( .A1(n7621), .A2(n7620), .ZN(n7602) );
  INV_X1 U9890 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n11108) );
  XOR2_X1 U9891 ( .A(n7605), .B(n11108), .Z(n7619) );
  XNOR2_X1 U9892 ( .A(P3_ADDR_REG_12__SCAN_IN), .B(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n7617) );
  NAND2_X1 U9893 ( .A1(n7616), .A2(n7617), .ZN(n7606) );
  OR2_X1 U9894 ( .A1(n14996), .A2(P3_ADDR_REG_13__SCAN_IN), .ZN(n7608) );
  NAND2_X1 U9895 ( .A1(n7613), .A2(n7612), .ZN(n7609) );
  NAND2_X1 U9896 ( .A1(n7665), .A2(n7664), .ZN(n7610) );
  OAI21_X1 U9897 ( .B1(P3_ADDR_REG_15__SCAN_IN), .B2(n15023), .A(n7610), .ZN(
        n7611) );
  INV_X1 U9898 ( .A(n7611), .ZN(n7667) );
  XOR2_X1 U9899 ( .A(n15041), .B(n7667), .Z(n7668) );
  XOR2_X1 U9900 ( .A(P3_ADDR_REG_16__SCAN_IN), .B(n7668), .Z(n14975) );
  XNOR2_X1 U9901 ( .A(n7613), .B(n7612), .ZN(n14967) );
  XNOR2_X1 U9902 ( .A(P3_ADDR_REG_13__SCAN_IN), .B(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n7615) );
  XOR2_X1 U9903 ( .A(n7615), .B(n7614), .Z(n14963) );
  XOR2_X1 U9904 ( .A(n7617), .B(n7616), .Z(n7660) );
  XNOR2_X1 U9905 ( .A(n7619), .B(n7618), .ZN(n14957) );
  XNOR2_X1 U9906 ( .A(n7621), .B(n7620), .ZN(n7623) );
  XNOR2_X1 U9907 ( .A(n7623), .B(n7622), .ZN(n7657) );
  XOR2_X1 U9908 ( .A(n7625), .B(n7624), .Z(n14801) );
  XNOR2_X1 U9909 ( .A(n7626), .B(n10374), .ZN(n15510) );
  XNOR2_X1 U9910 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(n7627), .ZN(n7637) );
  AND2_X1 U9911 ( .A1(n7637), .A2(P2_ADDR_REG_4__SCAN_IN), .ZN(n7638) );
  INV_X1 U9912 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n14250) );
  XNOR2_X1 U9913 ( .A(n7628), .B(n14250), .ZN(n15513) );
  XOR2_X1 U9914 ( .A(n7630), .B(n7629), .Z(n14787) );
  XNOR2_X1 U9915 ( .A(n7631), .B(n7632), .ZN(n7633) );
  INV_X1 U9916 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n15218) );
  NOR2_X1 U9917 ( .A1(n7633), .A2(n15218), .ZN(n7634) );
  INV_X1 U9918 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n15500) );
  AOI21_X1 U9919 ( .B1(n10610), .B2(P1_ADDR_REG_0__SCAN_IN), .A(n7632), .ZN(
        n15501) );
  NOR2_X1 U9920 ( .A1(n15500), .A2(n15501), .ZN(n15499) );
  INV_X1 U9921 ( .A(n15499), .ZN(n15518) );
  XNOR2_X1 U9922 ( .A(n15218), .B(n7633), .ZN(n15517) );
  NOR2_X1 U9923 ( .A1(n15518), .A2(n15517), .ZN(n15516) );
  NOR2_X1 U9924 ( .A1(n7634), .A2(n15516), .ZN(n14786) );
  NOR2_X1 U9925 ( .A1(n14787), .A2(n14786), .ZN(n7635) );
  NAND2_X1 U9926 ( .A1(n14787), .A2(n14786), .ZN(n14785) );
  OAI21_X1 U9927 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(n7635), .A(n14785), .ZN(
        n15512) );
  NAND2_X1 U9928 ( .A1(n15513), .A2(n15512), .ZN(n7636) );
  NOR2_X1 U9929 ( .A1(n15513), .A2(n15512), .ZN(n15511) );
  AOI21_X1 U9930 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(n7636), .A(n15511), .ZN(
        n15504) );
  XNOR2_X1 U9931 ( .A(P2_ADDR_REG_4__SCAN_IN), .B(n7637), .ZN(n15503) );
  NOR2_X1 U9932 ( .A1(n15504), .A2(n15503), .ZN(n15502) );
  INV_X1 U9933 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n14264) );
  XNOR2_X1 U9934 ( .A(n14264), .B(n7639), .ZN(n7641) );
  NAND2_X1 U9935 ( .A1(n7640), .A2(n7641), .ZN(n7643) );
  INV_X1 U9936 ( .A(n7640), .ZN(n7642) );
  INV_X1 U9937 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n15506) );
  INV_X1 U9938 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n7646) );
  XNOR2_X1 U9939 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(P3_ADDR_REG_6__SCAN_IN), 
        .ZN(n7645) );
  XNOR2_X1 U9940 ( .A(n7645), .B(n7644), .ZN(n14790) );
  NOR2_X1 U9941 ( .A1(n7647), .A2(n7646), .ZN(n7648) );
  INV_X1 U9942 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n7649) );
  XNOR2_X1 U9943 ( .A(n7652), .B(n7651), .ZN(n7653) );
  NAND2_X1 U9944 ( .A1(n7655), .A2(n7653), .ZN(n7656) );
  INV_X1 U9945 ( .A(n7653), .ZN(n7654) );
  INV_X1 U9946 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n14793) );
  NAND2_X1 U9947 ( .A1(n14794), .A2(n14793), .ZN(n14792) );
  INV_X1 U9948 ( .A(n14805), .ZN(n14806) );
  INV_X1 U9949 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n15271) );
  NAND2_X1 U9950 ( .A1(n7658), .A2(n7657), .ZN(n14807) );
  NAND2_X1 U9951 ( .A1(n15271), .A2(n14807), .ZN(n14804) );
  NAND2_X1 U9952 ( .A1(n14806), .A2(n14804), .ZN(n14956) );
  NOR2_X1 U9953 ( .A1(n14957), .A2(n14956), .ZN(n7659) );
  NAND2_X1 U9954 ( .A1(n14957), .A2(n14956), .ZN(n14955) );
  OAI21_X2 U9955 ( .B1(n7659), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n14955), .ZN(
        n7662) );
  INV_X1 U9956 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n15288) );
  NAND2_X1 U9957 ( .A1(n14967), .A2(n14966), .ZN(n14965) );
  XNOR2_X1 U9958 ( .A(n7665), .B(n7664), .ZN(n14970) );
  NAND2_X1 U9959 ( .A1(n14971), .A2(n14970), .ZN(n14969) );
  NAND2_X1 U9960 ( .A1(n7667), .A2(n15041), .ZN(n7670) );
  NAND2_X1 U9961 ( .A1(P3_ADDR_REG_16__SCAN_IN), .A2(n7668), .ZN(n7669) );
  NAND2_X1 U9962 ( .A1(n7670), .A2(n7669), .ZN(n7674) );
  XNOR2_X1 U9963 ( .A(P1_ADDR_REG_17__SCAN_IN), .B(n7674), .ZN(n7675) );
  XOR2_X1 U9964 ( .A(P3_ADDR_REG_17__SCAN_IN), .B(n7675), .Z(n7671) );
  INV_X1 U9965 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n14815) );
  NAND2_X1 U9966 ( .A1(n7672), .A2(n7671), .ZN(n7673) );
  XOR2_X1 U9967 ( .A(P3_ADDR_REG_18__SCAN_IN), .B(P1_ADDR_REG_18__SCAN_IN), 
        .Z(n7679) );
  INV_X1 U9968 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n15055) );
  NAND2_X1 U9969 ( .A1(n15055), .A2(n7674), .ZN(n7677) );
  NAND2_X1 U9970 ( .A1(P3_ADDR_REG_17__SCAN_IN), .A2(n7675), .ZN(n7676) );
  NAND2_X1 U9971 ( .A1(n7677), .A2(n7676), .ZN(n7678) );
  XNOR2_X1 U9972 ( .A(n7679), .B(n7678), .ZN(n14780) );
  INV_X1 U9973 ( .A(P3_ADDR_REG_18__SCAN_IN), .ZN(n7681) );
  NOR2_X1 U9974 ( .A1(n7679), .A2(n7678), .ZN(n7680) );
  AOI21_X1 U9975 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n7681), .A(n7680), .ZN(
        n7683) );
  XNOR2_X1 U9976 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(P1_ADDR_REG_19__SCAN_IN), 
        .ZN(n7682) );
  NOR2_X1 U9977 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n7688) );
  NOR2_X2 U9978 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n7686) );
  NAND4_X1 U9979 ( .A1(n7688), .A2(n7687), .A3(n7686), .A4(n7685), .ZN(n7993)
         );
  NAND4_X1 U9980 ( .A1(n7689), .A2(n8088), .A3(n7153), .A4(n8037), .ZN(n8254)
         );
  NOR2_X1 U9981 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n7693) );
  NAND2_X1 U9982 ( .A1(n7154), .A2(n7694), .ZN(n7695) );
  NOR2_X1 U9983 ( .A1(P1_IR_REG_25__SCAN_IN), .A2(P1_IR_REG_26__SCAN_IN), .ZN(
        n7699) );
  NAND4_X1 U9984 ( .A1(n7699), .A2(n8310), .A3(n7698), .A4(n8330), .ZN(n7700)
         );
  XNOR2_X2 U9985 ( .A(n7704), .B(P1_IR_REG_29__SCAN_IN), .ZN(n7706) );
  NAND2_X1 U9986 ( .A1(n7943), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n7712) );
  INV_X1 U9987 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n9783) );
  OR2_X1 U9988 ( .A1(n8244), .A2(n9783), .ZN(n7711) );
  NAND2_X1 U9989 ( .A1(n7707), .A2(n14762), .ZN(n7732) );
  INV_X1 U9990 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n7708) );
  XNOR2_X2 U9991 ( .A(n7716), .B(n7715), .ZN(n12173) );
  INV_X1 U9992 ( .A(n7723), .ZN(n7720) );
  INV_X1 U9993 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n9247) );
  INV_X1 U9994 ( .A(SI_0_), .ZN(n9885) );
  NAND2_X1 U9995 ( .A1(n7720), .A2(n7721), .ZN(n7747) );
  INV_X1 U9996 ( .A(n7721), .ZN(n7722) );
  NAND2_X1 U9997 ( .A1(n7723), .A2(n7722), .ZN(n7724) );
  AND2_X1 U9998 ( .A1(n7747), .A2(n7724), .ZN(n9811) );
  NAND2_X1 U9999 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n7725) );
  MUX2_X1 U10000 ( .A(P1_IR_REG_31__SCAN_IN), .B(n7725), .S(
        P1_IR_REG_1__SCAN_IN), .Z(n7727) );
  INV_X1 U10001 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n7726) );
  NAND2_X1 U10002 ( .A1(n14979), .A2(n7726), .ZN(n7755) );
  NAND2_X1 U10003 ( .A1(n7727), .A2(n7755), .ZN(n9923) );
  OR2_X1 U10004 ( .A1(n9905), .A2(n9923), .ZN(n7728) );
  INV_X1 U10005 ( .A(n13970), .ZN(n7739) );
  NAND2_X1 U10006 ( .A1(n14231), .A2(n13969), .ZN(n7729) );
  NAND2_X1 U10007 ( .A1(n7943), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n7737) );
  INV_X1 U10008 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n7730) );
  INV_X1 U10009 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n7731) );
  OR2_X1 U10010 ( .A1(n7732), .A2(n7731), .ZN(n7735) );
  INV_X1 U10011 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n7733) );
  OR2_X1 U10012 ( .A1(n6617), .A2(n7733), .ZN(n7734) );
  NOR2_X1 U10013 ( .A1(n7088), .A2(n9885), .ZN(n7738) );
  XNOR2_X1 U10014 ( .A(n7738), .B(P2_DATAO_REG_0__SCAN_IN), .ZN(n14777) );
  MUX2_X1 U10015 ( .A(n14979), .B(n14777), .S(n9905), .Z(n10389) );
  INV_X1 U10016 ( .A(n10389), .ZN(n10417) );
  NAND2_X1 U10017 ( .A1(n14233), .A2(n10417), .ZN(n9941) );
  INV_X1 U10018 ( .A(n9941), .ZN(n9773) );
  NAND2_X1 U10019 ( .A1(n7943), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n7745) );
  INV_X1 U10020 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n11062) );
  OR2_X1 U10021 ( .A1(n8244), .A2(n11062), .ZN(n7744) );
  INV_X1 U10022 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n9927) );
  OR2_X1 U10023 ( .A1(n7732), .A2(n9927), .ZN(n7743) );
  INV_X1 U10024 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n7741) );
  NAND2_X1 U10025 ( .A1(n7747), .A2(n7746), .ZN(n7752) );
  INV_X1 U10026 ( .A(n7752), .ZN(n7749) );
  NAND2_X1 U10027 ( .A1(n7748), .A2(SI_2_), .ZN(n7762) );
  OAI21_X1 U10028 ( .B1(n7748), .B2(SI_2_), .A(n7762), .ZN(n7750) );
  NAND2_X1 U10029 ( .A1(n7749), .A2(n7750), .ZN(n7753) );
  INV_X1 U10030 ( .A(n7750), .ZN(n7751) );
  INV_X2 U10031 ( .A(n8083), .ZN(n8060) );
  INV_X2 U10032 ( .A(n9905), .ZN(n8059) );
  NAND2_X1 U10033 ( .A1(n7755), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7754) );
  MUX2_X1 U10034 ( .A(P1_IR_REG_31__SCAN_IN), .B(n7754), .S(
        P1_IR_REG_2__SCAN_IN), .Z(n7758) );
  INV_X1 U10035 ( .A(n7755), .ZN(n7757) );
  INV_X1 U10036 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n7756) );
  NAND2_X1 U10037 ( .A1(n7757), .A2(n7756), .ZN(n7786) );
  INV_X1 U10038 ( .A(n9926), .ZN(n10449) );
  AND2_X2 U10039 ( .A1(n7760), .A2(n7759), .ZN(n15111) );
  NAND2_X1 U10040 ( .A1(n13976), .A2(n15111), .ZN(n13975) );
  INV_X1 U10041 ( .A(n13976), .ZN(n14230) );
  INV_X1 U10042 ( .A(n14168), .ZN(n11050) );
  NAND2_X1 U10043 ( .A1(n11052), .A2(n13975), .ZN(n10746) );
  MUX2_X1 U10044 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(P1_DATAO_REG_3__SCAN_IN), 
        .S(n8192), .Z(n7764) );
  NAND2_X1 U10045 ( .A1(n7764), .A2(SI_3_), .ZN(n7780) );
  INV_X1 U10046 ( .A(n7764), .ZN(n7765) );
  NAND2_X1 U10047 ( .A1(n7765), .A2(n10178), .ZN(n7766) );
  XNOR2_X1 U10048 ( .A(n7779), .B(n7777), .ZN(n9805) );
  NAND2_X1 U10049 ( .A1(n9805), .A2(n7767), .ZN(n7770) );
  NAND2_X1 U10050 ( .A1(n7786), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7768) );
  XNOR2_X1 U10051 ( .A(n7768), .B(P1_IR_REG_3__SCAN_IN), .ZN(n14252) );
  AOI22_X1 U10052 ( .A1(n8060), .A2(P2_DATAO_REG_3__SCAN_IN), .B1(n8059), .B2(
        n14252), .ZN(n7769) );
  NAND2_X1 U10053 ( .A1(n7770), .A2(n7769), .ZN(n13984) );
  OR2_X1 U10054 ( .A1(n8244), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n7774) );
  INV_X1 U10055 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n11032) );
  OR2_X1 U10056 ( .A1(n7732), .A2(n11032), .ZN(n7773) );
  INV_X1 U10057 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n7771) );
  OR2_X1 U10058 ( .A1(n13953), .A2(n7771), .ZN(n7772) );
  NAND4_X1 U10059 ( .A1(n7775), .A2(n7774), .A3(n7773), .A4(n7772), .ZN(n14229) );
  XNOR2_X1 U10060 ( .A(n13984), .B(n14229), .ZN(n14170) );
  NAND2_X1 U10061 ( .A1(n10746), .A2(n10745), .ZN(n10744) );
  OR2_X1 U10062 ( .A1(n14229), .A2(n13984), .ZN(n7776) );
  INV_X1 U10063 ( .A(n7777), .ZN(n7778) );
  NAND2_X1 U10064 ( .A1(n7779), .A2(n7778), .ZN(n7781) );
  NAND2_X1 U10065 ( .A1(n7781), .A2(n7780), .ZN(n7784) );
  INV_X1 U10066 ( .A(n7782), .ZN(n7783) );
  NAND2_X1 U10067 ( .A1(n7784), .A2(n7783), .ZN(n7801) );
  OR2_X1 U10068 ( .A1(n7784), .A2(n7783), .ZN(n7785) );
  AND2_X1 U10069 ( .A1(n7801), .A2(n7785), .ZN(n9810) );
  NAND2_X1 U10070 ( .A1(n9810), .A2(n7767), .ZN(n7793) );
  NAND2_X1 U10071 ( .A1(n7788), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7787) );
  MUX2_X1 U10072 ( .A(P1_IR_REG_31__SCAN_IN), .B(n7787), .S(
        P1_IR_REG_4__SCAN_IN), .Z(n7791) );
  INV_X1 U10073 ( .A(n7788), .ZN(n7790) );
  INV_X1 U10074 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n7789) );
  NAND2_X1 U10075 ( .A1(n7790), .A2(n7789), .ZN(n7809) );
  NAND2_X1 U10076 ( .A1(n7791), .A2(n7809), .ZN(n10465) );
  INV_X1 U10077 ( .A(n10465), .ZN(n9917) );
  AOI22_X1 U10078 ( .A1(n8060), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n8059), .B2(
        n9917), .ZN(n7792) );
  NAND2_X1 U10079 ( .A1(n7793), .A2(n7792), .ZN(n13990) );
  INV_X1 U10080 ( .A(n13990), .ZN(n15117) );
  NAND2_X1 U10081 ( .A1(n8243), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n7798) );
  INV_X1 U10082 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n9916) );
  OR2_X1 U10083 ( .A1(n13953), .A2(n9916), .ZN(n7797) );
  XNOR2_X1 U10084 ( .A(P1_REG3_REG_3__SCAN_IN), .B(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n11211) );
  OR2_X1 U10085 ( .A1(n8244), .A2(n11211), .ZN(n7796) );
  INV_X1 U10086 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n9929) );
  OR2_X1 U10087 ( .A1(n13954), .A2(n9929), .ZN(n7795) );
  INV_X1 U10088 ( .A(n14228), .ZN(n11192) );
  NAND2_X1 U10089 ( .A1(n10972), .A2(n15117), .ZN(n7799) );
  NAND2_X1 U10090 ( .A1(n7801), .A2(n7800), .ZN(n7806) );
  NAND2_X1 U10091 ( .A1(n7802), .A2(SI_5_), .ZN(n7821) );
  INV_X1 U10092 ( .A(n7802), .ZN(n7803) );
  NAND2_X1 U10093 ( .A1(n7803), .A2(n10076), .ZN(n7804) );
  AND2_X1 U10094 ( .A1(n7804), .A2(n7821), .ZN(n7805) );
  OR2_X1 U10095 ( .A1(n7806), .A2(n7805), .ZN(n7807) );
  OR2_X1 U10096 ( .A1(n9834), .A2(n14127), .ZN(n7812) );
  NAND2_X1 U10097 ( .A1(n7809), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7808) );
  MUX2_X1 U10098 ( .A(P1_IR_REG_31__SCAN_IN), .B(n7808), .S(
        P1_IR_REG_5__SCAN_IN), .Z(n7810) );
  AOI22_X1 U10099 ( .A1(n8060), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n8059), .B2(
        n14266), .ZN(n7811) );
  NAND2_X1 U10100 ( .A1(n7812), .A2(n7811), .ZN(n13999) );
  AOI21_X1 U10101 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(P1_REG3_REG_5__SCAN_IN), .ZN(n7813) );
  NOR2_X1 U10102 ( .A1(n7813), .A2(n7831), .ZN(n11195) );
  NAND2_X1 U10103 ( .A1(n8104), .A2(n11195), .ZN(n7818) );
  INV_X1 U10104 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n7814) );
  OR2_X1 U10105 ( .A1(n6617), .A2(n7814), .ZN(n7817) );
  INV_X1 U10106 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n9918) );
  OR2_X1 U10107 ( .A1(n13953), .A2(n9918), .ZN(n7816) );
  INV_X1 U10108 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n9930) );
  OR2_X1 U10109 ( .A1(n13954), .A2(n9930), .ZN(n7815) );
  NAND4_X1 U10110 ( .A1(n7818), .A2(n7817), .A3(n7816), .A4(n7815), .ZN(n14227) );
  XNOR2_X1 U10111 ( .A(n13999), .B(n11213), .ZN(n14174) );
  INV_X1 U10112 ( .A(n13999), .ZN(n15123) );
  NAND2_X1 U10113 ( .A1(n15123), .A2(n11213), .ZN(n7819) );
  NAND2_X1 U10114 ( .A1(n7820), .A2(n7819), .ZN(n15072) );
  MUX2_X1 U10115 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(P1_DATAO_REG_6__SCAN_IN), 
        .S(n8192), .Z(n7823) );
  NAND2_X1 U10116 ( .A1(n7823), .A2(SI_6_), .ZN(n7838) );
  OAI21_X1 U10117 ( .B1(SI_6_), .B2(n7823), .A(n7838), .ZN(n7824) );
  INV_X1 U10118 ( .A(n7824), .ZN(n7825) );
  OR2_X1 U10119 ( .A1(n7826), .A2(n7825), .ZN(n7827) );
  NAND2_X1 U10120 ( .A1(n7839), .A2(n7827), .ZN(n9832) );
  OR2_X1 U10121 ( .A1(n9832), .A2(n14127), .ZN(n7830) );
  NAND2_X1 U10122 ( .A1(n7845), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7828) );
  XNOR2_X1 U10123 ( .A(n7828), .B(P1_IR_REG_6__SCAN_IN), .ZN(n10376) );
  AOI22_X1 U10124 ( .A1(n8060), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n8059), .B2(
        n10376), .ZN(n7829) );
  NAND2_X1 U10125 ( .A1(n7830), .A2(n7829), .ZN(n15083) );
  NAND2_X1 U10126 ( .A1(n8243), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n7835) );
  INV_X1 U10127 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n9913) );
  OR2_X1 U10128 ( .A1(n13953), .A2(n9913), .ZN(n7834) );
  NAND2_X1 U10129 ( .A1(n7831), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n7870) );
  OAI21_X1 U10130 ( .B1(n7831), .B2(P1_REG3_REG_6__SCAN_IN), .A(n7870), .ZN(
        n15079) );
  OR2_X1 U10131 ( .A1(n8244), .A2(n15079), .ZN(n7833) );
  INV_X1 U10132 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n10384) );
  OR2_X1 U10133 ( .A1(n13954), .A2(n10384), .ZN(n7832) );
  NAND4_X1 U10134 ( .A1(n7835), .A2(n7834), .A3(n7833), .A4(n7832), .ZN(n14226) );
  XNOR2_X1 U10135 ( .A(n15083), .B(n14226), .ZN(n14175) );
  NAND2_X1 U10136 ( .A1(n15072), .A2(n15073), .ZN(n7837) );
  OR2_X1 U10137 ( .A1(n15083), .A2(n14226), .ZN(n7836) );
  NAND2_X1 U10138 ( .A1(n7837), .A2(n7836), .ZN(n11158) );
  MUX2_X1 U10139 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(P1_DATAO_REG_7__SCAN_IN), 
        .S(n8192), .Z(n7840) );
  NAND2_X1 U10140 ( .A1(n7840), .A2(SI_7_), .ZN(n7857) );
  OAI21_X1 U10141 ( .B1(n7840), .B2(SI_7_), .A(n7857), .ZN(n7841) );
  INV_X1 U10142 ( .A(n7841), .ZN(n7842) );
  OR2_X1 U10143 ( .A1(n7843), .A2(n7842), .ZN(n7844) );
  NAND2_X1 U10144 ( .A1(n7858), .A2(n7844), .ZN(n9892) );
  OR2_X1 U10145 ( .A1(n9892), .A2(n14127), .ZN(n7848) );
  OAI21_X1 U10146 ( .B1(n7845), .B2(P1_IR_REG_6__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n7846) );
  XNOR2_X1 U10147 ( .A(n7846), .B(P1_IR_REG_7__SCAN_IN), .ZN(n10989) );
  AOI22_X1 U10148 ( .A1(n8060), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n8059), .B2(
        n10989), .ZN(n7847) );
  NAND2_X1 U10149 ( .A1(n7848), .A2(n7847), .ZN(n15141) );
  NAND2_X1 U10150 ( .A1(n8243), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n7853) );
  INV_X1 U10151 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n10377) );
  OR2_X1 U10152 ( .A1(n13953), .A2(n10377), .ZN(n7852) );
  INV_X1 U10153 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n7849) );
  XNOR2_X1 U10154 ( .A(n7870), .B(n7849), .ZN(n11550) );
  OR2_X1 U10155 ( .A1(n8244), .A2(n11550), .ZN(n7851) );
  INV_X1 U10156 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n11162) );
  OR2_X1 U10157 ( .A1(n13954), .A2(n11162), .ZN(n7850) );
  NAND4_X1 U10158 ( .A1(n7853), .A2(n7852), .A3(n7851), .A4(n7850), .ZN(n14225) );
  XNOR2_X1 U10159 ( .A(n15141), .B(n14225), .ZN(n14176) );
  INV_X1 U10160 ( .A(n14176), .ZN(n7854) );
  NAND2_X1 U10161 ( .A1(n11158), .A2(n7854), .ZN(n7856) );
  OR2_X1 U10162 ( .A1(n15141), .A2(n14225), .ZN(n7855) );
  MUX2_X1 U10163 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(P1_DATAO_REG_8__SCAN_IN), 
        .S(n8192), .Z(n7859) );
  NAND2_X1 U10164 ( .A1(n7859), .A2(SI_8_), .ZN(n7878) );
  OAI21_X1 U10165 ( .B1(SI_8_), .B2(n7859), .A(n7878), .ZN(n7860) );
  INV_X1 U10166 ( .A(n7860), .ZN(n7861) );
  OR2_X1 U10167 ( .A1(n9895), .A2(n14127), .ZN(n7867) );
  NAND2_X1 U10168 ( .A1(n7864), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7863) );
  MUX2_X1 U10169 ( .A(P1_IR_REG_31__SCAN_IN), .B(n7863), .S(
        P1_IR_REG_8__SCAN_IN), .Z(n7865) );
  OR2_X1 U10170 ( .A1(n7864), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n7887) );
  NAND2_X1 U10171 ( .A1(n7865), .A2(n7887), .ZN(n10990) );
  INV_X1 U10172 ( .A(n10990), .ZN(n14280) );
  AOI22_X1 U10173 ( .A1(n8060), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n8059), .B2(
        n14280), .ZN(n7866) );
  NAND2_X1 U10174 ( .A1(n8243), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n7875) );
  INV_X1 U10175 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n10991) );
  OR2_X1 U10176 ( .A1(n13953), .A2(n10991), .ZN(n7874) );
  INV_X1 U10177 ( .A(n7870), .ZN(n7868) );
  AOI21_X1 U10178 ( .B1(n7868), .B2(P1_REG3_REG_7__SCAN_IN), .A(
        P1_REG3_REG_8__SCAN_IN), .ZN(n7871) );
  NAND2_X1 U10179 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_REG3_REG_7__SCAN_IN), 
        .ZN(n7869) );
  NOR2_X1 U10180 ( .A1(n7870), .A2(n7869), .ZN(n7891) );
  OR2_X1 U10181 ( .A1(n7871), .A2(n7891), .ZN(n11727) );
  OR2_X1 U10182 ( .A1(n8244), .A2(n11727), .ZN(n7873) );
  INV_X1 U10183 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n11230) );
  OR2_X1 U10184 ( .A1(n13954), .A2(n11230), .ZN(n7872) );
  NAND4_X1 U10185 ( .A1(n7875), .A2(n7874), .A3(n7873), .A4(n7872), .ZN(n14224) );
  XNOR2_X1 U10186 ( .A(n14018), .B(n14224), .ZN(n14178) );
  NAND2_X1 U10187 ( .A1(n11219), .A2(n11222), .ZN(n7877) );
  OR2_X1 U10188 ( .A1(n14018), .A2(n14224), .ZN(n7876) );
  NAND2_X1 U10189 ( .A1(n7877), .A2(n7876), .ZN(n14608) );
  MUX2_X1 U10190 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(P1_DATAO_REG_9__SCAN_IN), 
        .S(n8192), .Z(n7880) );
  NAND2_X1 U10191 ( .A1(n7880), .A2(SI_9_), .ZN(n7899) );
  OAI21_X1 U10192 ( .B1(n7880), .B2(SI_9_), .A(n7899), .ZN(n7881) );
  INV_X1 U10193 ( .A(n7881), .ZN(n7882) );
  OR2_X1 U10194 ( .A1(n7883), .A2(n7882), .ZN(n7884) );
  NAND2_X1 U10195 ( .A1(n7900), .A2(n7884), .ZN(n9901) );
  OR2_X1 U10196 ( .A1(n9901), .A2(n14127), .ZN(n7890) );
  NAND2_X1 U10197 ( .A1(n7887), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7885) );
  MUX2_X1 U10198 ( .A(P1_IR_REG_31__SCAN_IN), .B(n7885), .S(
        P1_IR_REG_9__SCAN_IN), .Z(n7886) );
  INV_X1 U10199 ( .A(n7886), .ZN(n7888) );
  NOR2_X1 U10200 ( .A1(n7888), .A2(n7919), .ZN(n14294) );
  AOI22_X1 U10201 ( .A1(n8060), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n8059), .B2(
        n14294), .ZN(n7889) );
  NAND2_X1 U10202 ( .A1(n8243), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n7896) );
  INV_X1 U10203 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n10992) );
  OR2_X1 U10204 ( .A1(n13953), .A2(n10992), .ZN(n7895) );
  NAND2_X1 U10205 ( .A1(n7891), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n7925) );
  OR2_X1 U10206 ( .A1(n7891), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n7892) );
  NAND2_X1 U10207 ( .A1(n7925), .A2(n7892), .ZN(n14603) );
  OR2_X1 U10208 ( .A1(n8244), .A2(n14603), .ZN(n7894) );
  INV_X1 U10209 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n14604) );
  OR2_X1 U10210 ( .A1(n13954), .A2(n14604), .ZN(n7893) );
  NAND4_X1 U10211 ( .A1(n7896), .A2(n7895), .A3(n7894), .A4(n7893), .ZN(n14223) );
  XNOR2_X1 U10212 ( .A(n15156), .B(n11990), .ZN(n14607) );
  NAND2_X1 U10213 ( .A1(n14608), .A2(n14607), .ZN(n7898) );
  OR2_X1 U10214 ( .A1(n15156), .A2(n14223), .ZN(n7897) );
  NAND2_X1 U10215 ( .A1(n7898), .A2(n7897), .ZN(n11634) );
  MUX2_X1 U10216 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(P1_DATAO_REG_10__SCAN_IN), 
        .S(n8192), .Z(n7901) );
  NAND2_X1 U10217 ( .A1(n7901), .A2(SI_10_), .ZN(n7916) );
  OAI21_X1 U10218 ( .B1(n7901), .B2(SI_10_), .A(n7916), .ZN(n7902) );
  INV_X1 U10219 ( .A(n7902), .ZN(n7903) );
  OR2_X1 U10220 ( .A1(n7904), .A2(n7903), .ZN(n7905) );
  NAND2_X1 U10221 ( .A1(n7917), .A2(n7905), .ZN(n9939) );
  OR2_X1 U10222 ( .A1(n9939), .A2(n14127), .ZN(n7909) );
  INV_X1 U10223 ( .A(n7919), .ZN(n7906) );
  NAND2_X1 U10224 ( .A1(n7906), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7907) );
  XNOR2_X1 U10225 ( .A(n7907), .B(P1_IR_REG_10__SCAN_IN), .ZN(n11104) );
  AOI22_X1 U10226 ( .A1(n8060), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n8059), 
        .B2(n11104), .ZN(n7908) );
  NAND2_X1 U10227 ( .A1(n8243), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n7913) );
  INV_X1 U10228 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n10987) );
  OR2_X1 U10229 ( .A1(n13953), .A2(n10987), .ZN(n7912) );
  XNOR2_X1 U10230 ( .A(n7925), .B(n7923), .ZN(n12063) );
  OR2_X1 U10231 ( .A1(n8244), .A2(n12063), .ZN(n7911) );
  INV_X1 U10232 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n11638) );
  OR2_X1 U10233 ( .A1(n13954), .A2(n11638), .ZN(n7910) );
  NAND4_X1 U10234 ( .A1(n7913), .A2(n7912), .A3(n7911), .A4(n7910), .ZN(n14222) );
  XNOR2_X1 U10235 ( .A(n14029), .B(n14222), .ZN(n14181) );
  OR2_X1 U10236 ( .A1(n14029), .A2(n14222), .ZN(n7914) );
  MUX2_X1 U10237 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(P1_DATAO_REG_11__SCAN_IN), 
        .S(n8192), .Z(n7934) );
  XNOR2_X1 U10238 ( .A(n7934), .B(SI_11_), .ZN(n7937) );
  NAND2_X1 U10239 ( .A1(n10289), .A2(n7767), .ZN(n7922) );
  INV_X1 U10240 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n7918) );
  NAND2_X1 U10241 ( .A1(n7919), .A2(n7918), .ZN(n7939) );
  NAND2_X1 U10242 ( .A1(n7939), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7920) );
  XNOR2_X1 U10243 ( .A(n7920), .B(P1_IR_REG_11__SCAN_IN), .ZN(n11276) );
  AOI22_X1 U10244 ( .A1(n8060), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n8059), 
        .B2(n11276), .ZN(n7921) );
  NAND2_X1 U10245 ( .A1(n7794), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n7931) );
  INV_X1 U10246 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n11100) );
  OR2_X1 U10247 ( .A1(n13953), .A2(n11100), .ZN(n7930) );
  INV_X1 U10248 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n7924) );
  OAI21_X1 U10249 ( .B1(n7925), .B2(n7923), .A(n7924), .ZN(n7926) );
  NAND2_X1 U10250 ( .A1(n7926), .A2(n7945), .ZN(n14913) );
  OR2_X1 U10251 ( .A1(n8244), .A2(n14913), .ZN(n7929) );
  INV_X1 U10252 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n7927) );
  OR2_X1 U10253 ( .A1(n6617), .A2(n7927), .ZN(n7928) );
  NAND4_X1 U10254 ( .A1(n7931), .A2(n7930), .A3(n7929), .A4(n7928), .ZN(n14221) );
  NOR2_X1 U10255 ( .A1(n14910), .A2(n14221), .ZN(n7933) );
  NAND2_X1 U10256 ( .A1(n14910), .A2(n14221), .ZN(n7932) );
  INV_X1 U10257 ( .A(n7934), .ZN(n7935) );
  NAND2_X1 U10258 ( .A1(n7935), .A2(n9838), .ZN(n7936) );
  MUX2_X1 U10259 ( .A(n7938), .B(n10488), .S(n8192), .Z(n7955) );
  XNOR2_X1 U10260 ( .A(n7955), .B(SI_12_), .ZN(n7953) );
  XNOR2_X1 U10261 ( .A(n7954), .B(n7953), .ZN(n10455) );
  NAND2_X1 U10262 ( .A1(n10455), .A2(n7767), .ZN(n7942) );
  NAND2_X1 U10263 ( .A1(n7956), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7940) );
  XNOR2_X1 U10264 ( .A(n7940), .B(P1_IR_REG_12__SCAN_IN), .ZN(n14319) );
  AOI22_X1 U10265 ( .A1(n8060), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n8059), 
        .B2(n14319), .ZN(n7941) );
  NAND2_X1 U10266 ( .A1(n8224), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n7952) );
  INV_X1 U10267 ( .A(n7962), .ZN(n7947) );
  NAND2_X1 U10268 ( .A1(n7945), .A2(n7944), .ZN(n7946) );
  NAND2_X1 U10269 ( .A1(n7947), .A2(n7946), .ZN(n13856) );
  OR2_X1 U10270 ( .A1(n8244), .A2(n13856), .ZN(n7951) );
  INV_X1 U10271 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n11848) );
  OR2_X1 U10272 ( .A1(n13954), .A2(n11848), .ZN(n7950) );
  INV_X1 U10273 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n7948) );
  OR2_X1 U10274 ( .A1(n6617), .A2(n7948), .ZN(n7949) );
  NAND4_X1 U10275 ( .A1(n7952), .A2(n7951), .A3(n7950), .A4(n7949), .ZN(n14220) );
  XNOR2_X1 U10276 ( .A(n14040), .B(n14220), .ZN(n14183) );
  MUX2_X1 U10277 ( .A(n10553), .B(n7174), .S(n8192), .Z(n7971) );
  XNOR2_X1 U10278 ( .A(n7971), .B(SI_13_), .ZN(n7969) );
  XNOR2_X1 U10279 ( .A(n7970), .B(n7969), .ZN(n10492) );
  NAND2_X1 U10280 ( .A1(n10492), .A2(n7767), .ZN(n7961) );
  OAI21_X1 U10281 ( .B1(n7956), .B2(P1_IR_REG_12__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n7958) );
  INV_X1 U10282 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n7957) );
  NAND2_X1 U10283 ( .A1(n7958), .A2(n7957), .ZN(n7978) );
  OR2_X1 U10284 ( .A1(n7958), .A2(n7957), .ZN(n7959) );
  AOI22_X1 U10285 ( .A1(n8060), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n8059), 
        .B2(n14993), .ZN(n7960) );
  NAND2_X1 U10286 ( .A1(n8243), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n7967) );
  INV_X1 U10287 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n14320) );
  OR2_X1 U10288 ( .A1(n13953), .A2(n14320), .ZN(n7966) );
  NAND2_X1 U10289 ( .A1(n7962), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n7983) );
  OR2_X1 U10290 ( .A1(n7962), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n7963) );
  NAND2_X1 U10291 ( .A1(n7983), .A2(n7963), .ZN(n13903) );
  OR2_X1 U10292 ( .A1(n8244), .A2(n13903), .ZN(n7965) );
  INV_X1 U10293 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n11860) );
  OR2_X1 U10294 ( .A1(n13954), .A2(n11860), .ZN(n7964) );
  NAND4_X1 U10295 ( .A1(n7967), .A2(n7966), .A3(n7965), .A4(n7964), .ZN(n14922) );
  XNOR2_X1 U10296 ( .A(n14043), .B(n14922), .ZN(n14185) );
  INV_X1 U10297 ( .A(n14185), .ZN(n11854) );
  NAND2_X1 U10298 ( .A1(n11855), .A2(n11854), .ZN(n11853) );
  OR2_X1 U10299 ( .A1(n14043), .A2(n14922), .ZN(n7968) );
  NAND2_X1 U10300 ( .A1(n7971), .A2(n9897), .ZN(n7972) );
  MUX2_X1 U10301 ( .A(n9448), .B(n10823), .S(n8192), .Z(n7975) );
  NAND2_X1 U10302 ( .A1(n7976), .A2(n7975), .ZN(n7977) );
  NAND2_X1 U10303 ( .A1(n7992), .A2(n7977), .ZN(n10821) );
  NAND2_X1 U10304 ( .A1(n7978), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7979) );
  XNOR2_X1 U10305 ( .A(n7979), .B(P1_IR_REG_14__SCAN_IN), .ZN(n15000) );
  AOI22_X1 U10306 ( .A1(n15000), .A2(n8059), .B1(n8060), .B2(
        P2_DATAO_REG_14__SCAN_IN), .ZN(n7980) );
  NAND2_X1 U10307 ( .A1(n7794), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n7989) );
  INV_X1 U10308 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n14317) );
  OR2_X1 U10309 ( .A1(n13953), .A2(n14317), .ZN(n7988) );
  INV_X1 U10310 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n7982) );
  NAND2_X1 U10311 ( .A1(n7983), .A2(n7982), .ZN(n7984) );
  NAND2_X1 U10312 ( .A1(n8004), .A2(n7984), .ZN(n14918) );
  OR2_X1 U10313 ( .A1(n8244), .A2(n14918), .ZN(n7987) );
  INV_X1 U10314 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n7985) );
  OR2_X1 U10315 ( .A1(n6617), .A2(n7985), .ZN(n7986) );
  OR2_X1 U10316 ( .A1(n14946), .A2(n13904), .ZN(n14051) );
  NAND2_X1 U10317 ( .A1(n14946), .A2(n13904), .ZN(n14055) );
  NAND2_X2 U10318 ( .A1(n6652), .A2(n14931), .ZN(n14929) );
  INV_X1 U10319 ( .A(n13904), .ZN(n14584) );
  NAND2_X1 U10320 ( .A1(n14946), .A2(n14584), .ZN(n7990) );
  MUX2_X1 U10321 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(P1_DATAO_REG_15__SCAN_IN), 
        .S(n7088), .Z(n8015) );
  XNOR2_X1 U10322 ( .A(n8017), .B(n8016), .ZN(n11069) );
  NAND2_X1 U10323 ( .A1(n11069), .A2(n7767), .ZN(n8002) );
  INV_X1 U10324 ( .A(n7993), .ZN(n7996) );
  NAND2_X1 U10325 ( .A1(n7999), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7997) );
  MUX2_X1 U10326 ( .A(P1_IR_REG_31__SCAN_IN), .B(n7997), .S(
        P1_IR_REG_15__SCAN_IN), .Z(n7998) );
  INV_X1 U10327 ( .A(n7998), .ZN(n8000) );
  NOR2_X1 U10328 ( .A1(n8000), .A2(n8038), .ZN(n14322) );
  AOI22_X1 U10329 ( .A1(n8060), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n8059), 
        .B2(n14322), .ZN(n8001) );
  AND2_X1 U10330 ( .A1(n8004), .A2(n8003), .ZN(n8005) );
  OR2_X1 U10331 ( .A1(n8005), .A2(n8022), .ZN(n14585) );
  INV_X1 U10332 ( .A(n14585), .ZN(n8006) );
  NAND2_X1 U10333 ( .A1(n8104), .A2(n8006), .ZN(n8013) );
  INV_X1 U10334 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n8007) );
  OR2_X1 U10335 ( .A1(n13953), .A2(n8007), .ZN(n8012) );
  INV_X1 U10336 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n8008) );
  OR2_X1 U10337 ( .A1(n13954), .A2(n8008), .ZN(n8011) );
  INV_X1 U10338 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n8009) );
  OR2_X1 U10339 ( .A1(n6617), .A2(n8009), .ZN(n8010) );
  AND2_X1 U10340 ( .A1(n14590), .A2(n14920), .ZN(n14053) );
  INV_X1 U10341 ( .A(n14053), .ZN(n14056) );
  INV_X1 U10342 ( .A(n14920), .ZN(n14567) );
  OR2_X1 U10343 ( .A1(n14590), .A2(n14567), .ZN(n8014) );
  MUX2_X1 U10344 ( .A(n11238), .B(n11269), .S(n8192), .Z(n8033) );
  XNOR2_X1 U10345 ( .A(n8033), .B(SI_16_), .ZN(n8031) );
  XNOR2_X1 U10346 ( .A(n6782), .B(n8031), .ZN(n11237) );
  NAND2_X1 U10347 ( .A1(n11237), .A2(n7767), .ZN(n8021) );
  OR2_X1 U10348 ( .A1(n8038), .A2(n8018), .ZN(n8019) );
  XNOR2_X1 U10349 ( .A(n8019), .B(P1_IR_REG_16__SCAN_IN), .ZN(n14316) );
  AOI22_X1 U10350 ( .A1(n8060), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n8059), 
        .B2(n14316), .ZN(n8020) );
  NOR2_X1 U10351 ( .A1(n8022), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n8023) );
  OR2_X1 U10352 ( .A1(n8042), .A2(n8023), .ZN(n14572) );
  NAND2_X1 U10353 ( .A1(n7794), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n8024) );
  OAI21_X1 U10354 ( .B1(n14572), .B2(n8244), .A(n8024), .ZN(n8028) );
  INV_X1 U10355 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n8026) );
  NAND2_X1 U10356 ( .A1(n8224), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n8025) );
  OAI21_X1 U10357 ( .B1(n8026), .B2(n6617), .A(n8025), .ZN(n8027) );
  NAND2_X1 U10358 ( .A1(n14705), .A2(n14582), .ZN(n8029) );
  NAND2_X1 U10359 ( .A1(n8030), .A2(n8029), .ZN(n14187) );
  NAND2_X1 U10360 ( .A1(n8033), .A2(n10425), .ZN(n8034) );
  MUX2_X1 U10361 ( .A(n6806), .B(n11291), .S(n8192), .Z(n8052) );
  XNOR2_X1 U10362 ( .A(n8052), .B(SI_17_), .ZN(n8036) );
  XNOR2_X1 U10363 ( .A(n8050), .B(n8036), .ZN(n11285) );
  NAND2_X1 U10364 ( .A1(n11285), .A2(n7767), .ZN(n8041) );
  NAND2_X1 U10365 ( .A1(n8056), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8039) );
  XNOR2_X1 U10366 ( .A(n8039), .B(P1_IR_REG_17__SCAN_IN), .ZN(n15052) );
  AOI22_X1 U10367 ( .A1(n8060), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n8059), 
        .B2(n15052), .ZN(n8040) );
  OR2_X1 U10368 ( .A1(n8042), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n8043) );
  AND2_X1 U10369 ( .A1(n8063), .A2(n8043), .ZN(n14552) );
  NAND2_X1 U10370 ( .A1(n14552), .A2(n8104), .ZN(n8046) );
  AOI22_X1 U10371 ( .A1(n8243), .A2(P1_REG0_REG_17__SCAN_IN), .B1(n8224), .B2(
        P1_REG1_REG_17__SCAN_IN), .ZN(n8045) );
  NAND2_X1 U10372 ( .A1(n7794), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n8044) );
  INV_X1 U10373 ( .A(n14063), .ZN(n14566) );
  NAND2_X1 U10374 ( .A1(n14698), .A2(n14566), .ZN(n8047) );
  OR2_X1 U10375 ( .A1(n14698), .A2(n14566), .ZN(n8048) );
  INV_X1 U10376 ( .A(SI_17_), .ZN(n9499) );
  NAND2_X1 U10377 ( .A1(n8052), .A2(n9499), .ZN(n8051) );
  INV_X1 U10378 ( .A(n8052), .ZN(n8053) );
  NAND2_X1 U10379 ( .A1(n8053), .A2(SI_17_), .ZN(n8070) );
  MUX2_X1 U10380 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(P1_DATAO_REG_18__SCAN_IN), 
        .S(n7088), .Z(n8069) );
  XNOR2_X1 U10381 ( .A(n8069), .B(SI_18_), .ZN(n8054) );
  NAND2_X1 U10382 ( .A1(n8057), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8058) );
  XNOR2_X1 U10383 ( .A(n8058), .B(n8084), .ZN(n14329) );
  INV_X1 U10384 ( .A(n14329), .ZN(n15066) );
  AOI22_X1 U10385 ( .A1(n8060), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n8059), 
        .B2(n15066), .ZN(n8061) );
  INV_X1 U10386 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n8062) );
  NAND2_X1 U10387 ( .A1(n8063), .A2(n8062), .ZN(n8064) );
  NAND2_X1 U10388 ( .A1(n8094), .A2(n8064), .ZN(n14538) );
  OR2_X1 U10389 ( .A1(n14538), .A2(n8244), .ZN(n8067) );
  AOI22_X1 U10390 ( .A1(n8243), .A2(P1_REG0_REG_18__SCAN_IN), .B1(n8224), .B2(
        P1_REG1_REG_18__SCAN_IN), .ZN(n8066) );
  INV_X1 U10391 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n15062) );
  OR2_X1 U10392 ( .A1(n13954), .A2(n15062), .ZN(n8065) );
  NAND2_X1 U10393 ( .A1(n14537), .A2(n6943), .ZN(n8068) );
  OAI21_X1 U10394 ( .B1(n8074), .B2(n9506), .A(n8070), .ZN(n8071) );
  INV_X1 U10395 ( .A(n8071), .ZN(n8072) );
  NAND2_X1 U10396 ( .A1(n8074), .A2(n9506), .ZN(n8075) );
  MUX2_X1 U10397 ( .A(n7176), .B(n11532), .S(n7088), .Z(n8077) );
  INV_X1 U10398 ( .A(SI_19_), .ZN(n10725) );
  INV_X1 U10399 ( .A(n8077), .ZN(n8078) );
  NAND2_X1 U10400 ( .A1(n8078), .A2(SI_19_), .ZN(n8079) );
  OR2_X1 U10401 ( .A1(n8081), .A2(n8080), .ZN(n8082) );
  NAND2_X1 U10402 ( .A1(n8099), .A2(n8082), .ZN(n11530) );
  NAND2_X1 U10403 ( .A1(n11530), .A2(n7767), .ZN(n8093) );
  NAND2_X1 U10404 ( .A1(n8087), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8086) );
  OAI22_X1 U10405 ( .A1(n8083), .A2(n7176), .B1(n14917), .B2(n9905), .ZN(n8091) );
  INV_X1 U10406 ( .A(n8091), .ZN(n8092) );
  INV_X1 U10407 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n13839) );
  NAND2_X1 U10408 ( .A1(n8094), .A2(n13839), .ZN(n8095) );
  NAND2_X1 U10409 ( .A1(n8102), .A2(n8095), .ZN(n14529) );
  AOI22_X1 U10410 ( .A1(n8243), .A2(P1_REG0_REG_19__SCAN_IN), .B1(n8224), .B2(
        P1_REG1_REG_19__SCAN_IN), .ZN(n8097) );
  INV_X1 U10411 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n14530) );
  OR2_X1 U10412 ( .A1(n13954), .A2(n14530), .ZN(n8096) );
  OAI211_X1 U10413 ( .C1(n14529), .C2(n8244), .A(n8097), .B(n8096), .ZN(n14545) );
  INV_X1 U10414 ( .A(n14545), .ZN(n14062) );
  XNOR2_X1 U10415 ( .A(n14528), .B(n14062), .ZN(n14523) );
  INV_X1 U10416 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n12325) );
  MUX2_X1 U10417 ( .A(n12313), .B(n12325), .S(n7088), .Z(n8129) );
  XNOR2_X1 U10418 ( .A(n8113), .B(n8129), .ZN(n12312) );
  NAND2_X1 U10419 ( .A1(n12312), .A2(n7767), .ZN(n8101) );
  OR2_X1 U10420 ( .A1(n8083), .A2(n12313), .ZN(n8100) );
  INV_X1 U10421 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n13896) );
  AND2_X1 U10422 ( .A1(n8102), .A2(n13896), .ZN(n8103) );
  NOR2_X1 U10423 ( .A1(n8120), .A2(n8103), .ZN(n14513) );
  NAND2_X1 U10424 ( .A1(n14513), .A2(n8104), .ZN(n8110) );
  INV_X1 U10425 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n8107) );
  NAND2_X1 U10426 ( .A1(n8243), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n8106) );
  INV_X1 U10427 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n14516) );
  OR2_X1 U10428 ( .A1(n13954), .A2(n14516), .ZN(n8105) );
  OAI211_X1 U10429 ( .C1(n13953), .C2(n8107), .A(n8106), .B(n8105), .ZN(n8108)
         );
  INV_X1 U10430 ( .A(n8108), .ZN(n8109) );
  NAND2_X1 U10431 ( .A1(n14518), .A2(n14085), .ZN(n8111) );
  OR2_X1 U10432 ( .A1(n14674), .A2(n14085), .ZN(n8112) );
  INV_X1 U10433 ( .A(n8129), .ZN(n8128) );
  NAND2_X1 U10434 ( .A1(n8113), .A2(n8128), .ZN(n8115) );
  INV_X1 U10435 ( .A(SI_20_), .ZN(n11240) );
  OR2_X1 U10436 ( .A1(n8127), .A2(n11240), .ZN(n8114) );
  NAND2_X1 U10437 ( .A1(n8115), .A2(n8114), .ZN(n8117) );
  MUX2_X1 U10438 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(P1_DATAO_REG_21__SCAN_IN), 
        .S(n7088), .Z(n8130) );
  XNOR2_X1 U10439 ( .A(n8130), .B(SI_21_), .ZN(n8116) );
  NAND2_X1 U10440 ( .A1(n11828), .A2(n7767), .ZN(n8119) );
  INV_X1 U10441 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n11832) );
  OR2_X1 U10442 ( .A1(n8083), .A2(n11832), .ZN(n8118) );
  NOR2_X1 U10443 ( .A1(n8120), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n8121) );
  OR2_X1 U10444 ( .A1(n8135), .A2(n8121), .ZN(n14501) );
  INV_X1 U10445 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n14741) );
  NAND2_X1 U10446 ( .A1(n7794), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n8123) );
  NAND2_X1 U10447 ( .A1(n8224), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n8122) );
  OAI211_X1 U10448 ( .C1(n6617), .C2(n14741), .A(n8123), .B(n8122), .ZN(n8124)
         );
  INV_X1 U10449 ( .A(n8124), .ZN(n8125) );
  OAI21_X1 U10450 ( .B1(n14501), .B2(n8244), .A(n8125), .ZN(n14218) );
  XNOR2_X1 U10451 ( .A(n14739), .B(n14218), .ZN(n14496) );
  OR2_X1 U10452 ( .A1(n14739), .A2(n14218), .ZN(n8126) );
  NOR2_X1 U10453 ( .A1(n8129), .A2(n11240), .ZN(n8131) );
  AOI22_X1 U10454 ( .A1(n8131), .A2(n7577), .B1(n8130), .B2(SI_21_), .ZN(n8132) );
  OR2_X1 U10455 ( .A1(n8675), .A2(n7088), .ZN(n8134) );
  XNOR2_X1 U10456 ( .A(n8134), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n14775) );
  NOR2_X1 U10457 ( .A1(n8135), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n8136) );
  OR2_X1 U10458 ( .A1(n8147), .A2(n8136), .ZN(n14479) );
  INV_X1 U10459 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n14478) );
  NAND2_X1 U10460 ( .A1(n8224), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n8138) );
  NAND2_X1 U10461 ( .A1(n8243), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n8137) );
  OAI211_X1 U10462 ( .C1(n14478), .C2(n13954), .A(n8138), .B(n8137), .ZN(n8139) );
  INV_X1 U10463 ( .A(n8139), .ZN(n8140) );
  OAI21_X1 U10464 ( .B1(n14479), .B2(n8244), .A(n8140), .ZN(n14217) );
  INV_X1 U10465 ( .A(n14217), .ZN(n12255) );
  XNOR2_X1 U10466 ( .A(n14738), .B(n12255), .ZN(n14191) );
  INV_X1 U10467 ( .A(n14191), .ZN(n14484) );
  OR2_X1 U10468 ( .A1(n14481), .A2(n14217), .ZN(n8141) );
  MUX2_X1 U10469 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(P1_DATAO_REG_22__SCAN_IN), 
        .S(n7088), .Z(n8674) );
  INV_X1 U10470 ( .A(n8674), .ZN(n8144) );
  NAND2_X1 U10471 ( .A1(n8142), .A2(SI_22_), .ZN(n8143) );
  MUX2_X1 U10472 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(P1_DATAO_REG_23__SCAN_IN), 
        .S(n7088), .Z(n8157) );
  XNOR2_X1 U10473 ( .A(n8157), .B(SI_23_), .ZN(n8154) );
  XNOR2_X1 U10474 ( .A(n8156), .B(n8154), .ZN(n11999) );
  NAND2_X1 U10475 ( .A1(n11999), .A2(n7767), .ZN(n8146) );
  INV_X1 U10476 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n11998) );
  OR2_X1 U10477 ( .A1(n8083), .A2(n11998), .ZN(n8145) );
  OR2_X1 U10478 ( .A1(n8147), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n8148) );
  NAND2_X1 U10479 ( .A1(n8147), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n8162) );
  NAND2_X1 U10480 ( .A1(n8148), .A2(n8162), .ZN(n14467) );
  INV_X1 U10481 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n10207) );
  NAND2_X1 U10482 ( .A1(n8224), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n8150) );
  NAND2_X1 U10483 ( .A1(n7794), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n8149) );
  OAI211_X1 U10484 ( .C1(n10207), .C2(n6617), .A(n8150), .B(n8149), .ZN(n8151)
         );
  INV_X1 U10485 ( .A(n8151), .ZN(n8152) );
  OAI21_X1 U10486 ( .B1(n14467), .B2(n8244), .A(n8152), .ZN(n14216) );
  INV_X1 U10487 ( .A(n14216), .ZN(n8287) );
  XNOR2_X1 U10488 ( .A(n14732), .B(n8287), .ZN(n14463) );
  NAND2_X1 U10489 ( .A1(n14732), .A2(n14216), .ZN(n8153) );
  INV_X1 U10490 ( .A(n8154), .ZN(n8155) );
  NAND2_X1 U10491 ( .A1(n8157), .A2(SI_23_), .ZN(n8158) );
  MUX2_X1 U10492 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(P1_DATAO_REG_24__SCAN_IN), 
        .S(n7088), .Z(n8171) );
  XNOR2_X1 U10493 ( .A(n8170), .B(n8171), .ZN(n12133) );
  NAND2_X1 U10494 ( .A1(n12133), .A2(n7767), .ZN(n8160) );
  INV_X1 U10495 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n12135) );
  OR2_X1 U10496 ( .A1(n8083), .A2(n12135), .ZN(n8159) );
  NAND2_X1 U10497 ( .A1(n8224), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n8167) );
  INV_X1 U10498 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n8161) );
  OR2_X1 U10499 ( .A1(n6617), .A2(n8161), .ZN(n8166) );
  OAI21_X1 U10500 ( .B1(P1_REG3_REG_24__SCAN_IN), .B2(n8163), .A(n8182), .ZN(
        n14452) );
  OR2_X1 U10501 ( .A1(n8244), .A2(n14452), .ZN(n8165) );
  INV_X1 U10502 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n14453) );
  OR2_X1 U10503 ( .A1(n13954), .A2(n14453), .ZN(n8164) );
  NAND4_X1 U10504 ( .A1(n8167), .A2(n8166), .A3(n8165), .A4(n8164), .ZN(n14215) );
  INV_X1 U10505 ( .A(n14215), .ZN(n8288) );
  XNOR2_X1 U10506 ( .A(n14728), .B(n8288), .ZN(n14441) );
  INV_X1 U10507 ( .A(n14441), .ZN(n14447) );
  OR2_X1 U10508 ( .A1(n14728), .A2(n14215), .ZN(n8168) );
  INV_X1 U10509 ( .A(n8170), .ZN(n8172) );
  NAND2_X1 U10510 ( .A1(n8172), .A2(n8171), .ZN(n8175) );
  NAND2_X1 U10511 ( .A1(n8173), .A2(SI_24_), .ZN(n8174) );
  INV_X1 U10512 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n13805) );
  MUX2_X1 U10513 ( .A(n14773), .B(n13805), .S(n7088), .Z(n8176) );
  INV_X1 U10514 ( .A(SI_25_), .ZN(n12091) );
  NAND2_X1 U10515 ( .A1(n8176), .A2(n12091), .ZN(n8189) );
  INV_X1 U10516 ( .A(n8176), .ZN(n8177) );
  NAND2_X1 U10517 ( .A1(n8177), .A2(SI_25_), .ZN(n8178) );
  NAND2_X1 U10518 ( .A1(n8189), .A2(n8178), .ZN(n8190) );
  NAND2_X1 U10519 ( .A1(n13802), .A2(n7767), .ZN(n8180) );
  OR2_X1 U10520 ( .A1(n8083), .A2(n14773), .ZN(n8179) );
  NAND2_X1 U10521 ( .A1(n8243), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n8187) );
  INV_X1 U10522 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n8181) );
  OR2_X1 U10523 ( .A1(n13953), .A2(n8181), .ZN(n8186) );
  INV_X1 U10524 ( .A(n8182), .ZN(n8183) );
  INV_X1 U10525 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n10183) );
  OAI21_X1 U10526 ( .B1(P1_REG3_REG_25__SCAN_IN), .B2(n8183), .A(n8195), .ZN(
        n14433) );
  OR2_X1 U10527 ( .A1(n8244), .A2(n14433), .ZN(n8185) );
  INV_X1 U10528 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n14434) );
  OR2_X1 U10529 ( .A1(n13954), .A2(n14434), .ZN(n8184) );
  NAND4_X1 U10530 ( .A1(n8187), .A2(n8186), .A3(n8185), .A4(n8184), .ZN(n14214) );
  INV_X1 U10531 ( .A(n14214), .ZN(n8290) );
  XNOR2_X1 U10532 ( .A(n14724), .B(n8290), .ZN(n14430) );
  NAND2_X1 U10533 ( .A1(n14428), .A2(n14430), .ZN(n14429) );
  NAND2_X1 U10534 ( .A1(n14724), .A2(n14214), .ZN(n8188) );
  NAND2_X1 U10535 ( .A1(n14429), .A2(n8188), .ZN(n14412) );
  INV_X1 U10536 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n14768) );
  MUX2_X1 U10537 ( .A(n14768), .B(n13800), .S(n8192), .Z(n8205) );
  XNOR2_X1 U10538 ( .A(n8205), .B(SI_26_), .ZN(n8203) );
  NAND2_X1 U10539 ( .A1(n13799), .A2(n7767), .ZN(n8194) );
  OR2_X1 U10540 ( .A1(n8083), .A2(n14768), .ZN(n8193) );
  NAND2_X1 U10541 ( .A1(n8224), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n8202) );
  INV_X1 U10542 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n14414) );
  OR2_X1 U10543 ( .A1(n13954), .A2(n14414), .ZN(n8201) );
  INV_X1 U10544 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n10222) );
  INV_X1 U10545 ( .A(n8225), .ZN(n8196) );
  OAI21_X1 U10546 ( .B1(P1_REG3_REG_26__SCAN_IN), .B2(n8197), .A(n8196), .ZN(
        n14416) );
  OR2_X1 U10547 ( .A1(n8244), .A2(n14416), .ZN(n8200) );
  INV_X1 U10548 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n8198) );
  OR2_X1 U10549 ( .A1(n6617), .A2(n8198), .ZN(n8199) );
  NAND4_X1 U10550 ( .A1(n8202), .A2(n8201), .A3(n8200), .A4(n8199), .ZN(n14213) );
  XNOR2_X1 U10551 ( .A(n14419), .B(n14213), .ZN(n14411) );
  INV_X1 U10552 ( .A(n14411), .ZN(n14409) );
  INV_X1 U10553 ( .A(n8205), .ZN(n8206) );
  INV_X1 U10554 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n13797) );
  MUX2_X1 U10555 ( .A(n14767), .B(n13797), .S(n7088), .Z(n8215) );
  INV_X1 U10556 ( .A(n8215), .ZN(n8216) );
  XNOR2_X1 U10557 ( .A(n8216), .B(SI_27_), .ZN(n8207) );
  NAND2_X1 U10558 ( .A1(n13796), .A2(n7767), .ZN(n8209) );
  OR2_X1 U10559 ( .A1(n8083), .A2(n14767), .ZN(n8208) );
  NAND2_X1 U10560 ( .A1(n8224), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n8213) );
  INV_X1 U10561 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n14719) );
  OR2_X1 U10562 ( .A1(n6617), .A2(n14719), .ZN(n8212) );
  XNOR2_X1 U10563 ( .A(P1_REG3_REG_27__SCAN_IN), .B(n8225), .ZN(n14400) );
  OR2_X1 U10564 ( .A1(n8244), .A2(n14400), .ZN(n8211) );
  INV_X1 U10565 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n14401) );
  OR2_X1 U10566 ( .A1(n13954), .A2(n14401), .ZN(n8210) );
  NAND4_X1 U10567 ( .A1(n8213), .A2(n8212), .A3(n8211), .A4(n8210), .ZN(n14377) );
  XNOR2_X1 U10568 ( .A(n14629), .B(n14377), .ZN(n14193) );
  INV_X1 U10569 ( .A(n14193), .ZN(n14394) );
  OR2_X1 U10570 ( .A1(n14629), .A2(n14377), .ZN(n8214) );
  INV_X1 U10571 ( .A(SI_27_), .ZN(n13166) );
  INV_X1 U10572 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n8218) );
  MUX2_X1 U10573 ( .A(n9669), .B(n8218), .S(n7088), .Z(n8238) );
  XNOR2_X1 U10574 ( .A(n8238), .B(SI_28_), .ZN(n8219) );
  OR2_X1 U10575 ( .A1(n8220), .A2(n8219), .ZN(n8221) );
  NAND2_X1 U10576 ( .A1(n8220), .A2(n8219), .ZN(n8240) );
  NAND2_X1 U10577 ( .A1(n8221), .A2(n8240), .ZN(n13793) );
  NAND2_X1 U10578 ( .A1(n13793), .A2(n7767), .ZN(n8223) );
  OR2_X1 U10579 ( .A1(n8083), .A2(n9669), .ZN(n8222) );
  NAND2_X1 U10580 ( .A1(n8224), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n8234) );
  INV_X1 U10581 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n14385) );
  OR2_X1 U10582 ( .A1(n13954), .A2(n14385), .ZN(n8233) );
  NAND2_X1 U10583 ( .A1(n8226), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n14358) );
  INV_X1 U10584 ( .A(n8226), .ZN(n8228) );
  INV_X1 U10585 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n8227) );
  NAND2_X1 U10586 ( .A1(n8228), .A2(n8227), .ZN(n8229) );
  NAND2_X1 U10587 ( .A1(n14358), .A2(n8229), .ZN(n14384) );
  OR2_X1 U10588 ( .A1(n8244), .A2(n14384), .ZN(n8232) );
  INV_X1 U10589 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n8230) );
  OR2_X1 U10590 ( .A1(n6617), .A2(n8230), .ZN(n8231) );
  NAND4_X1 U10591 ( .A1(n8234), .A2(n8233), .A3(n8232), .A4(n8231), .ZN(n14125) );
  INV_X1 U10592 ( .A(n14125), .ZN(n8235) );
  NAND2_X1 U10593 ( .A1(n14627), .A2(n8235), .ZN(n8295) );
  OR2_X1 U10594 ( .A1(n14627), .A2(n8235), .ZN(n8236) );
  NAND2_X1 U10595 ( .A1(n14627), .A2(n14125), .ZN(n8237) );
  NAND2_X1 U10596 ( .A1(n14380), .A2(n8237), .ZN(n8250) );
  INV_X1 U10597 ( .A(SI_28_), .ZN(n13163) );
  NAND2_X1 U10598 ( .A1(n8238), .A2(n13163), .ZN(n8239) );
  INV_X1 U10599 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n13790) );
  MUX2_X1 U10600 ( .A(n14764), .B(n13790), .S(n7088), .Z(n9078) );
  XNOR2_X1 U10601 ( .A(n9078), .B(SI_29_), .ZN(n9076) );
  NAND2_X1 U10602 ( .A1(n13789), .A2(n7767), .ZN(n8242) );
  OR2_X1 U10603 ( .A1(n8083), .A2(n14764), .ZN(n8241) );
  INV_X1 U10604 ( .A(n14365), .ZN(n14139) );
  NAND2_X1 U10605 ( .A1(n8243), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n8249) );
  INV_X1 U10606 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n8885) );
  OR2_X1 U10607 ( .A1(n13953), .A2(n8885), .ZN(n8248) );
  OR2_X1 U10608 ( .A1(n8244), .A2(n14358), .ZN(n8247) );
  INV_X1 U10609 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n8245) );
  OR2_X1 U10610 ( .A1(n13954), .A2(n8245), .ZN(n8246) );
  XNOR2_X1 U10611 ( .A(n14139), .B(n14138), .ZN(n14196) );
  INV_X1 U10612 ( .A(n14196), .ZN(n8296) );
  XNOR2_X1 U10613 ( .A(n8253), .B(n8252), .ZN(n8262) );
  INV_X1 U10614 ( .A(n8038), .ZN(n8255) );
  OAI21_X1 U10615 ( .B1(n8255), .B2(n8254), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n8256) );
  MUX2_X1 U10616 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8256), .S(
        P1_IR_REG_21__SCAN_IN), .Z(n8257) );
  INV_X1 U10617 ( .A(n14155), .ZN(n8258) );
  NAND2_X1 U10618 ( .A1(n8311), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8259) );
  AOI21_X1 U10619 ( .B1(n10390), .B2(n14776), .A(n8345), .ZN(n8261) );
  AND2_X1 U10620 ( .A1(n14917), .A2(n14776), .ZN(n8260) );
  OR2_X2 U10621 ( .A1(n8260), .A2(n10390), .ZN(n12208) );
  AND2_X1 U10622 ( .A1(n8345), .A2(n13959), .ZN(n15094) );
  NAND2_X1 U10623 ( .A1(n15094), .A2(n8305), .ZN(n15159) );
  NAND2_X1 U10624 ( .A1(n14357), .A2(n15170), .ZN(n8309) );
  NAND2_X1 U10625 ( .A1(n14231), .A2(n10561), .ZN(n8263) );
  NAND2_X1 U10626 ( .A1(n13966), .A2(n8263), .ZN(n13965) );
  NAND2_X1 U10627 ( .A1(n13965), .A2(n13967), .ZN(n11055) );
  NAND2_X1 U10628 ( .A1(n11055), .A2(n14168), .ZN(n11054) );
  NAND2_X1 U10629 ( .A1(n13976), .A2(n13978), .ZN(n8264) );
  NAND2_X1 U10630 ( .A1(n11054), .A2(n8264), .ZN(n10749) );
  INV_X1 U10631 ( .A(n14229), .ZN(n13985) );
  NAND2_X1 U10632 ( .A1(n13985), .A2(n13984), .ZN(n8265) );
  INV_X1 U10633 ( .A(n14174), .ZN(n11042) );
  NAND2_X1 U10634 ( .A1(n13999), .A2(n11213), .ZN(n8267) );
  INV_X1 U10635 ( .A(n14226), .ZN(n11191) );
  AND2_X1 U10636 ( .A1(n15083), .A2(n11191), .ZN(n8269) );
  OR2_X1 U10637 ( .A1(n15083), .A2(n11191), .ZN(n8268) );
  INV_X1 U10638 ( .A(n14225), .ZN(n11544) );
  NOR2_X1 U10639 ( .A1(n15141), .A2(n11544), .ZN(n8270) );
  OAI22_X1 U10640 ( .A1(n11159), .A2(n8270), .B1(n11557), .B2(n14225), .ZN(
        n11223) );
  INV_X1 U10641 ( .A(n14224), .ZN(n14600) );
  OR2_X1 U10642 ( .A1(n14018), .A2(n14600), .ZN(n8271) );
  NAND2_X1 U10643 ( .A1(n15156), .A2(n11990), .ZN(n8272) );
  INV_X1 U10644 ( .A(n14222), .ZN(n14899) );
  INV_X1 U10645 ( .A(n14221), .ZN(n12177) );
  NAND2_X1 U10646 ( .A1(n14910), .A2(n12177), .ZN(n8273) );
  NAND2_X1 U10647 ( .A1(n11695), .A2(n8273), .ZN(n8275) );
  OR2_X1 U10648 ( .A1(n14910), .A2(n12177), .ZN(n8274) );
  NAND2_X1 U10649 ( .A1(n8275), .A2(n8274), .ZN(n11844) );
  NAND2_X1 U10650 ( .A1(n11844), .A2(n14183), .ZN(n8277) );
  INV_X1 U10651 ( .A(n14220), .ZN(n14898) );
  OR2_X1 U10652 ( .A1(n14040), .A2(n14898), .ZN(n8276) );
  INV_X1 U10653 ( .A(n14922), .ZN(n14887) );
  OR2_X1 U10654 ( .A1(n14043), .A2(n14887), .ZN(n8278) );
  INV_X1 U10655 ( .A(n14055), .ZN(n8280) );
  INV_X1 U10656 ( .A(n14582), .ZN(n14550) );
  XNOR2_X1 U10657 ( .A(n14698), .B(n14063), .ZN(n14560) );
  INV_X1 U10658 ( .A(n14560), .ZN(n8281) );
  OR2_X1 U10659 ( .A1(n14698), .A2(n14063), .ZN(n14071) );
  NAND2_X1 U10660 ( .A1(n14537), .A2(n14551), .ZN(n14078) );
  NAND2_X1 U10661 ( .A1(n14528), .A2(n14062), .ZN(n14082) );
  NAND2_X1 U10662 ( .A1(n14508), .A2(n14512), .ZN(n14507) );
  INV_X1 U10663 ( .A(n14218), .ZN(n8284) );
  OR2_X1 U10664 ( .A1(n14739), .A2(n8284), .ZN(n14483) );
  AND2_X1 U10665 ( .A1(n14191), .A2(n14483), .ZN(n8285) );
  NAND2_X1 U10666 ( .A1(n14481), .A2(n12255), .ZN(n8286) );
  INV_X1 U10667 ( .A(n14463), .ZN(n14458) );
  OR2_X1 U10668 ( .A1(n14728), .A2(n8288), .ZN(n8289) );
  NAND2_X1 U10669 ( .A1(n14443), .A2(n8289), .ZN(n14423) );
  NAND2_X1 U10670 ( .A1(n14724), .A2(n8290), .ZN(n8291) );
  INV_X1 U10671 ( .A(n14213), .ZN(n12285) );
  AND2_X1 U10672 ( .A1(n14419), .A2(n12285), .ZN(n8292) );
  INV_X1 U10673 ( .A(n14377), .ZN(n8293) );
  NAND2_X1 U10674 ( .A1(n14629), .A2(n8293), .ZN(n14373) );
  NAND2_X1 U10675 ( .A1(n8294), .A2(n14372), .ZN(n14375) );
  NAND2_X1 U10676 ( .A1(n14375), .A2(n8295), .ZN(n8297) );
  XNOR2_X1 U10677 ( .A(n8297), .B(n8296), .ZN(n14369) );
  OR2_X1 U10678 ( .A1(n13959), .A2(n14155), .ZN(n8299) );
  NAND2_X1 U10679 ( .A1(n8345), .A2(n14776), .ZN(n8298) );
  INV_X1 U10680 ( .A(n14029), .ZN(n15167) );
  AND2_X1 U10681 ( .A1(n10561), .A2(n10389), .ZN(n11064) );
  NAND2_X1 U10682 ( .A1(n11064), .A2(n15111), .ZN(n11063) );
  OR2_X1 U10683 ( .A1(n11063), .A2(n13984), .ZN(n10974) );
  NAND2_X1 U10684 ( .A1(n15167), .A2(n14613), .ZN(n11697) );
  OR2_X1 U10685 ( .A1(n14555), .A2(n14537), .ZN(n14536) );
  NAND2_X2 U10686 ( .A1(n13959), .A2(n8344), .ZN(n14915) );
  OAI211_X1 U10687 ( .C1(n14365), .C2(n14383), .A(n15086), .B(n14350), .ZN(
        n14366) );
  INV_X1 U10688 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n8301) );
  NOR2_X1 U10689 ( .A1(n13953), .A2(n8301), .ZN(n8304) );
  INV_X1 U10690 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n14353) );
  NOR2_X1 U10691 ( .A1(n13954), .A2(n14353), .ZN(n8303) );
  INV_X1 U10692 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n10231) );
  NOR2_X1 U10693 ( .A1(n6617), .A2(n10231), .ZN(n8302) );
  OR3_X1 U10694 ( .A1(n8304), .A2(n8303), .A3(n8302), .ZN(n14212) );
  INV_X1 U10695 ( .A(n13949), .ZN(n10407) );
  NAND2_X1 U10696 ( .A1(n10407), .A2(n12173), .ZN(n14919) );
  NOR2_X1 U10697 ( .A1(n6625), .A2(n10211), .ZN(n8306) );
  NOR2_X1 U10698 ( .A1(n14919), .A2(n8306), .ZN(n14345) );
  NAND2_X1 U10699 ( .A1(n14212), .A2(n14345), .ZN(n14359) );
  INV_X1 U10700 ( .A(n12173), .ZN(n10441) );
  NAND2_X1 U10701 ( .A1(n10407), .A2(n10441), .ZN(n14601) );
  NAND2_X1 U10702 ( .A1(n14125), .A2(n14921), .ZN(n14361) );
  NAND3_X1 U10703 ( .A1(n14366), .A2(n14359), .A3(n14361), .ZN(n8307) );
  AOI21_X1 U10704 ( .B1(n14369), .B2(n14952), .A(n8307), .ZN(n8308) );
  NOR2_X2 U10705 ( .A1(n8311), .A2(P1_IR_REG_22__SCAN_IN), .ZN(n8328) );
  NAND2_X1 U10706 ( .A1(n8328), .A2(n8330), .ZN(n8314) );
  INV_X1 U10707 ( .A(n8314), .ZN(n8312) );
  NAND2_X1 U10708 ( .A1(n8312), .A2(n7698), .ZN(n8318) );
  NOR2_X1 U10709 ( .A1(n8325), .A2(n10211), .ZN(n8316) );
  NAND2_X1 U10710 ( .A1(n8314), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8315) );
  INV_X1 U10711 ( .A(n8324), .ZN(n12134) );
  MUX2_X1 U10712 ( .A(n10211), .B(n8316), .S(n12134), .Z(n8317) );
  INV_X1 U10713 ( .A(n8317), .ZN(n8322) );
  OAI22_X1 U10714 ( .A1(n9813), .A2(P1_D_REG_1__SCAN_IN), .B1(n9815), .B2(
        n8325), .ZN(n10405) );
  NAND2_X1 U10715 ( .A1(n13959), .A2(n14917), .ZN(n8323) );
  NAND2_X1 U10716 ( .A1(n8323), .A2(n10407), .ZN(n8327) );
  INV_X1 U10717 ( .A(n8328), .ZN(n8329) );
  NAND2_X1 U10718 ( .A1(n8329), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8331) );
  NAND2_X1 U10719 ( .A1(n10414), .A2(n9825), .ZN(n14206) );
  INV_X1 U10720 ( .A(n14206), .ZN(n10419) );
  INV_X1 U10721 ( .A(n9813), .ZN(n8342) );
  NOR4_X1 U10722 ( .A1(P1_D_REG_3__SCAN_IN), .A2(P1_D_REG_4__SCAN_IN), .A3(
        P1_D_REG_5__SCAN_IN), .A4(P1_D_REG_6__SCAN_IN), .ZN(n8340) );
  NOR4_X1 U10723 ( .A1(P1_D_REG_7__SCAN_IN), .A2(P1_D_REG_10__SCAN_IN), .A3(
        P1_D_REG_11__SCAN_IN), .A4(P1_D_REG_12__SCAN_IN), .ZN(n8339) );
  OR4_X1 U10724 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_9__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_2__SCAN_IN), .ZN(n8337) );
  NOR4_X1 U10725 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_18__SCAN_IN), .A3(
        P1_D_REG_19__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n8335) );
  NOR4_X1 U10726 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_13__SCAN_IN), .A3(
        P1_D_REG_14__SCAN_IN), .A4(P1_D_REG_16__SCAN_IN), .ZN(n8334) );
  NOR4_X1 U10727 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_27__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n8333) );
  NOR4_X1 U10728 ( .A1(P1_D_REG_21__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_23__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n8332) );
  NAND4_X1 U10729 ( .A1(n8335), .A2(n8334), .A3(n8333), .A4(n8332), .ZN(n8336)
         );
  NOR4_X1 U10730 ( .A1(P1_D_REG_28__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        n8337), .A4(n8336), .ZN(n8338) );
  NAND3_X1 U10731 ( .A1(n8340), .A2(n8339), .A3(n8338), .ZN(n8341) );
  NAND2_X1 U10732 ( .A1(n8342), .A2(n8341), .ZN(n10402) );
  NAND4_X1 U10733 ( .A1(n10405), .A2(n10419), .A3(n10402), .A4(n10412), .ZN(
        n8884) );
  INV_X1 U10734 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n9827) );
  NAND2_X1 U10735 ( .A1(n8342), .A2(n9827), .ZN(n8343) );
  INV_X1 U10736 ( .A(n9815), .ZN(n14770) );
  NAND2_X1 U10737 ( .A1(n14770), .A2(n12134), .ZN(n9824) );
  INV_X1 U10738 ( .A(n10404), .ZN(n9780) );
  INV_X1 U10739 ( .A(n8344), .ZN(n9942) );
  NAND2_X1 U10740 ( .A1(n8345), .A2(n8344), .ZN(n8346) );
  NAND2_X1 U10741 ( .A1(n15174), .A2(n15155), .ZN(n14748) );
  NAND2_X1 U10742 ( .A1(n15172), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n8347) );
  AND2_X2 U10743 ( .A1(n8382), .A2(n8348), .ZN(n8406) );
  AND2_X2 U10744 ( .A1(n6667), .A2(n8406), .ZN(n8477) );
  NOR2_X1 U10745 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), 
        .ZN(n8351) );
  NAND4_X1 U10746 ( .A1(n8351), .A2(n8350), .A3(n8349), .A4(n8532), .ZN(n8591)
         );
  NAND3_X1 U10747 ( .A1(n8480), .A2(n8352), .A3(n8594), .ZN(n8353) );
  NOR2_X2 U10748 ( .A1(n8591), .A2(n8353), .ZN(n8354) );
  NOR2_X1 U10749 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), 
        .ZN(n8357) );
  NOR2_X1 U10750 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), 
        .ZN(n8356) );
  NOR2_X1 U10751 ( .A1(P2_IR_REG_23__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), 
        .ZN(n8355) );
  NAND4_X1 U10752 ( .A1(n8357), .A2(n8356), .A3(n8355), .A4(n8788), .ZN(n8774)
         );
  INV_X1 U10753 ( .A(n8774), .ZN(n8359) );
  NOR3_X1 U10754 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_25__SCAN_IN), 
        .A3(P2_IR_REG_26__SCAN_IN), .ZN(n8358) );
  NAND2_X1 U10755 ( .A1(n8362), .A2(n8361), .ZN(n8365) );
  XNOR2_X2 U10756 ( .A(n8364), .B(n8363), .ZN(n8368) );
  NAND2_X1 U10757 ( .A1(n8379), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8366) );
  MUX2_X1 U10758 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8366), .S(
        P2_IR_REG_29__SCAN_IN), .Z(n8367) );
  NAND2_X1 U10759 ( .A1(n8424), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n8374) );
  NAND2_X1 U10760 ( .A1(n8412), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n8373) );
  NAND2_X2 U10761 ( .A1(n8370), .A2(n13791), .ZN(n8415) );
  INV_X1 U10762 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n10312) );
  OR2_X1 U10763 ( .A1(n8415), .A2(n10312), .ZN(n8371) );
  NAND2_X1 U10764 ( .A1(n8376), .A2(P2_IR_REG_28__SCAN_IN), .ZN(n8378) );
  INV_X1 U10765 ( .A(n9811), .ZN(n8380) );
  INV_X1 U10766 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n8396) );
  NAND2_X1 U10767 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), 
        .ZN(n8381) );
  MUX2_X1 U10768 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8381), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n8384) );
  INV_X1 U10769 ( .A(n8403), .ZN(n8383) );
  NAND2_X1 U10770 ( .A1(n8384), .A2(n8383), .ZN(n10313) );
  INV_X1 U10771 ( .A(n10313), .ZN(n15208) );
  NAND2_X1 U10772 ( .A1(n8389), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n8394) );
  NAND2_X1 U10773 ( .A1(n8424), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n8393) );
  NAND2_X1 U10774 ( .A1(n8412), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n8392) );
  INV_X1 U10775 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n8390) );
  OR2_X1 U10776 ( .A1(n8415), .A2(n8390), .ZN(n8391) );
  NAND4_X1 U10777 ( .A1(n8394), .A2(n8393), .A3(n8392), .A4(n8391), .ZN(n13384) );
  NAND2_X1 U10778 ( .A1(n7088), .A2(SI_0_), .ZN(n8395) );
  XNOR2_X1 U10779 ( .A(n8395), .B(n9214), .ZN(n13806) );
  MUX2_X1 U10780 ( .A(n8396), .B(n13806), .S(n10292), .Z(n10639) );
  NAND2_X1 U10781 ( .A1(n13384), .A2(n10727), .ZN(n9793) );
  INV_X1 U10782 ( .A(n13383), .ZN(n10649) );
  NAND2_X1 U10783 ( .A1(n10649), .A2(n10648), .ZN(n8397) );
  NAND2_X1 U10784 ( .A1(n9792), .A2(n8397), .ZN(n13654) );
  INV_X1 U10785 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n8398) );
  NAND2_X1 U10786 ( .A1(n8424), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n8401) );
  NAND2_X1 U10787 ( .A1(n8412), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n8400) );
  INV_X1 U10788 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n13663) );
  OR2_X1 U10789 ( .A1(n8415), .A2(n13663), .ZN(n8399) );
  INV_X1 U10790 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n9818) );
  NOR2_X1 U10791 ( .A1(n8403), .A2(n8803), .ZN(n8404) );
  MUX2_X1 U10792 ( .A(n8803), .B(n8404), .S(P2_IR_REG_2__SCAN_IN), .Z(n8405)
         );
  INV_X1 U10793 ( .A(n8405), .ZN(n8408) );
  INV_X1 U10794 ( .A(n8406), .ZN(n8407) );
  NAND2_X1 U10795 ( .A1(n8408), .A2(n8407), .ZN(n15223) );
  OAI22_X1 U10796 ( .A1(n8590), .A2(n9818), .B1(n10292), .B2(n15223), .ZN(
        n8410) );
  NAND2_X1 U10797 ( .A1(n13654), .A2(n6621), .ZN(n13653) );
  INV_X1 U10798 ( .A(n13382), .ZN(n10598) );
  NAND2_X1 U10799 ( .A1(n10598), .A2(n10651), .ZN(n8411) );
  NAND2_X1 U10800 ( .A1(n8412), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n8417) );
  INV_X1 U10801 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n8414) );
  INV_X1 U10802 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n10314) );
  INV_X4 U10803 ( .A(n8438), .ZN(n9085) );
  NAND2_X1 U10804 ( .A1(n9805), .A2(n9085), .ZN(n8422) );
  INV_X2 U10805 ( .A(n8590), .ZN(n8614) );
  NOR2_X1 U10806 ( .A1(n8406), .A2(n8803), .ZN(n8418) );
  MUX2_X1 U10807 ( .A(n8803), .B(n8418), .S(P2_IR_REG_3__SCAN_IN), .Z(n8420)
         );
  AND2_X1 U10808 ( .A1(n8406), .A2(n8419), .ZN(n8431) );
  NOR2_X1 U10809 ( .A1(n8420), .A2(n8431), .ZN(n10315) );
  AOI22_X1 U10810 ( .A1(n8614), .A2(P1_DATAO_REG_3__SCAN_IN), .B1(n8636), .B2(
        n10315), .ZN(n8421) );
  NAND2_X1 U10811 ( .A1(n10594), .A2(n10593), .ZN(n10592) );
  NAND2_X1 U10812 ( .A1(n10650), .A2(n10736), .ZN(n8423) );
  NAND2_X1 U10813 ( .A1(n10592), .A2(n8423), .ZN(n10761) );
  NAND2_X1 U10814 ( .A1(n8412), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n8430) );
  NOR2_X1 U10815 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n8425) );
  NOR2_X1 U10816 ( .A1(n8445), .A2(n8425), .ZN(n11128) );
  NAND2_X1 U10817 ( .A1(n8424), .A2(n11128), .ZN(n8429) );
  INV_X1 U10818 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n8426) );
  OR2_X1 U10819 ( .A1(n8870), .A2(n8426), .ZN(n8428) );
  INV_X1 U10820 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n11133) );
  OR2_X1 U10821 ( .A1(n9090), .A2(n11133), .ZN(n8427) );
  NAND4_X1 U10822 ( .A1(n8430), .A2(n8429), .A3(n8428), .A4(n8427), .ZN(n13380) );
  NAND2_X1 U10823 ( .A1(n9810), .A2(n9085), .ZN(n8436) );
  INV_X1 U10824 ( .A(n8431), .ZN(n8433) );
  NAND2_X1 U10825 ( .A1(n8433), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8432) );
  MUX2_X1 U10826 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8432), .S(
        P2_IR_REG_4__SCAN_IN), .Z(n8434) );
  AND2_X1 U10827 ( .A1(n8434), .A2(n8440), .ZN(n10316) );
  AOI22_X1 U10828 ( .A1(n8614), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n8636), .B2(
        n10316), .ZN(n8435) );
  NAND2_X1 U10829 ( .A1(n8436), .A2(n8435), .ZN(n10843) );
  XNOR2_X1 U10830 ( .A(n10599), .B(n10843), .ZN(n10760) );
  NAND2_X1 U10831 ( .A1(n10761), .A2(n10760), .ZN(n10759) );
  OR2_X1 U10832 ( .A1(n10843), .A2(n13380), .ZN(n8437) );
  NAND2_X1 U10833 ( .A1(n8440), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8439) );
  MUX2_X1 U10834 ( .A(n8439), .B(P2_IR_REG_31__SCAN_IN), .S(n8441), .Z(n8443)
         );
  INV_X1 U10835 ( .A(n8440), .ZN(n8442) );
  NAND2_X1 U10836 ( .A1(n8442), .A2(n8441), .ZN(n8463) );
  NAND2_X1 U10837 ( .A1(n8443), .A2(n8463), .ZN(n10359) );
  INV_X1 U10838 ( .A(n10359), .ZN(n10318) );
  AOI22_X1 U10839 ( .A1(n8614), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n8636), .B2(
        n10318), .ZN(n8444) );
  NAND2_X1 U10840 ( .A1(n6627), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n8451) );
  NOR2_X1 U10841 ( .A1(n8445), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n8446) );
  NOR2_X1 U10842 ( .A1(n8456), .A2(n8446), .ZN(n11327) );
  NAND2_X1 U10843 ( .A1(n8424), .A2(n11327), .ZN(n8450) );
  INV_X1 U10844 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n8447) );
  OR2_X1 U10845 ( .A1(n8870), .A2(n8447), .ZN(n8449) );
  INV_X1 U10846 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n10317) );
  OR2_X1 U10847 ( .A1(n9090), .A2(n10317), .ZN(n8448) );
  NAND4_X1 U10848 ( .A1(n8451), .A2(n8450), .A3(n8449), .A4(n8448), .ZN(n13379) );
  XNOR2_X1 U10849 ( .A(n10965), .B(n13379), .ZN(n9145) );
  INV_X1 U10850 ( .A(n9145), .ZN(n10961) );
  NAND2_X1 U10851 ( .A1(n10959), .A2(n10961), .ZN(n10958) );
  INV_X1 U10852 ( .A(n10965), .ZN(n11330) );
  INV_X1 U10853 ( .A(n13379), .ZN(n10927) );
  NAND2_X1 U10854 ( .A1(n11330), .A2(n10927), .ZN(n8452) );
  NAND2_X1 U10855 ( .A1(n10958), .A2(n8452), .ZN(n11114) );
  OR2_X1 U10856 ( .A1(n9832), .A2(n9107), .ZN(n8455) );
  NAND2_X1 U10857 ( .A1(n8463), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8453) );
  XNOR2_X1 U10858 ( .A(n8453), .B(P2_IR_REG_6__SCAN_IN), .ZN(n10344) );
  AOI22_X1 U10859 ( .A1(n8614), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n8636), .B2(
        n10344), .ZN(n8454) );
  NAND2_X1 U10860 ( .A1(n8455), .A2(n8454), .ZN(n11123) );
  NAND2_X1 U10861 ( .A1(n8456), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n8469) );
  OAI21_X1 U10862 ( .B1(n8456), .B2(P2_REG3_REG_6__SCAN_IN), .A(n8469), .ZN(
        n11142) );
  OR2_X1 U10863 ( .A1(n8748), .A2(n11142), .ZN(n8461) );
  NAND2_X1 U10864 ( .A1(n6627), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n8460) );
  INV_X1 U10865 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n8457) );
  OR2_X1 U10866 ( .A1(n8870), .A2(n8457), .ZN(n8459) );
  INV_X1 U10867 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n11141) );
  OR2_X1 U10868 ( .A1(n9090), .A2(n11141), .ZN(n8458) );
  NAND4_X1 U10869 ( .A1(n8461), .A2(n8460), .A3(n8459), .A4(n8458), .ZN(n13378) );
  XNOR2_X1 U10870 ( .A(n11123), .B(n13378), .ZN(n9147) );
  INV_X1 U10871 ( .A(n9147), .ZN(n11118) );
  NAND2_X1 U10872 ( .A1(n11114), .A2(n11118), .ZN(n11113) );
  OR2_X1 U10873 ( .A1(n11123), .A2(n13378), .ZN(n8462) );
  OR2_X1 U10874 ( .A1(n9892), .A2(n9107), .ZN(n8466) );
  OAI21_X1 U10875 ( .B1(n8463), .B2(P2_IR_REG_6__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8464) );
  XNOR2_X1 U10876 ( .A(n8464), .B(P2_IR_REG_7__SCAN_IN), .ZN(n13392) );
  AOI22_X1 U10877 ( .A1(n8614), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n8636), .B2(
        n13392), .ZN(n8465) );
  NAND2_X1 U10878 ( .A1(n6627), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n8475) );
  AND2_X1 U10879 ( .A1(n8469), .A2(n8468), .ZN(n8470) );
  NOR2_X1 U10880 ( .A1(n8485), .A2(n8470), .ZN(n15327) );
  NAND2_X1 U10881 ( .A1(n8424), .A2(n15327), .ZN(n8474) );
  INV_X1 U10882 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n8471) );
  OR2_X1 U10883 ( .A1(n8870), .A2(n8471), .ZN(n8473) );
  INV_X1 U10884 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n10337) );
  OR2_X1 U10885 ( .A1(n9090), .A2(n10337), .ZN(n8472) );
  NAND4_X1 U10886 ( .A1(n8475), .A2(n8474), .A3(n8473), .A4(n8472), .ZN(n13377) );
  INV_X1 U10887 ( .A(n13377), .ZN(n10928) );
  XNOR2_X1 U10888 ( .A(n15323), .B(n10928), .ZN(n11259) );
  OR2_X1 U10889 ( .A1(n15323), .A2(n13377), .ZN(n8476) );
  OR2_X1 U10890 ( .A1(n9895), .A2(n9107), .ZN(n8484) );
  NOR2_X1 U10891 ( .A1(n8478), .A2(n8803), .ZN(n8479) );
  MUX2_X1 U10892 ( .A(n8803), .B(n8479), .S(P2_IR_REG_8__SCAN_IN), .Z(n8482)
         );
  NAND2_X1 U10893 ( .A1(n8478), .A2(n8480), .ZN(n8506) );
  INV_X1 U10894 ( .A(n8506), .ZN(n8481) );
  NOR2_X1 U10895 ( .A1(n8482), .A2(n8481), .ZN(n10477) );
  AOI22_X1 U10896 ( .A1(n8614), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n8636), .B2(
        n10477), .ZN(n8483) );
  NAND2_X1 U10897 ( .A1(n8485), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n8497) );
  OR2_X1 U10898 ( .A1(n8485), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n8486) );
  NAND2_X1 U10899 ( .A1(n8497), .A2(n8486), .ZN(n11460) );
  OR2_X1 U10900 ( .A1(n8748), .A2(n11460), .ZN(n8491) );
  NAND2_X1 U10901 ( .A1(n6627), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n8490) );
  INV_X1 U10902 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n8487) );
  OR2_X1 U10903 ( .A1(n8870), .A2(n8487), .ZN(n8489) );
  INV_X1 U10904 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n11461) );
  OR2_X1 U10905 ( .A1(n9090), .A2(n11461), .ZN(n8488) );
  NAND4_X1 U10906 ( .A1(n8491), .A2(n8490), .A3(n8489), .A4(n8488), .ZN(n13376) );
  XNOR2_X1 U10907 ( .A(n15364), .B(n13376), .ZN(n11453) );
  NAND2_X1 U10908 ( .A1(n15364), .A2(n13376), .ZN(n8492) );
  OR2_X1 U10909 ( .A1(n9901), .A2(n9107), .ZN(n8495) );
  NAND2_X1 U10910 ( .A1(n8506), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8493) );
  XNOR2_X1 U10911 ( .A(n8493), .B(P2_IR_REG_9__SCAN_IN), .ZN(n15253) );
  AOI22_X1 U10912 ( .A1(n8614), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n8636), .B2(
        n15253), .ZN(n8494) );
  INV_X1 U10913 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n8496) );
  NAND2_X1 U10914 ( .A1(n8497), .A2(n8496), .ZN(n8498) );
  NAND2_X1 U10915 ( .A1(n8511), .A2(n8498), .ZN(n11567) );
  OR2_X1 U10916 ( .A1(n8748), .A2(n11567), .ZN(n8503) );
  NAND2_X1 U10917 ( .A1(n6627), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n8502) );
  INV_X1 U10918 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n8499) );
  OR2_X1 U10919 ( .A1(n8870), .A2(n8499), .ZN(n8501) );
  OR2_X1 U10920 ( .A1(n9090), .A2(n10471), .ZN(n8500) );
  NAND4_X1 U10921 ( .A1(n8503), .A2(n8502), .A3(n8501), .A4(n8500), .ZN(n13375) );
  XNOR2_X1 U10922 ( .A(n11746), .B(n13375), .ZN(n9149) );
  NAND2_X1 U10923 ( .A1(n11558), .A2(n11559), .ZN(n8505) );
  NAND2_X1 U10924 ( .A1(n11746), .A2(n13375), .ZN(n8504) );
  OR2_X1 U10925 ( .A1(n9939), .A2(n9107), .ZN(n8509) );
  NAND2_X1 U10926 ( .A1(n8593), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8507) );
  XNOR2_X1 U10927 ( .A(n8507), .B(P2_IR_REG_10__SCAN_IN), .ZN(n15264) );
  AOI22_X1 U10928 ( .A1(n8614), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n8636), 
        .B2(n15264), .ZN(n8508) );
  NAND2_X1 U10929 ( .A1(n6627), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n8518) );
  INV_X1 U10930 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n8510) );
  AND2_X1 U10931 ( .A1(n8511), .A2(n8510), .ZN(n8512) );
  NOR2_X1 U10932 ( .A1(n8540), .A2(n8512), .ZN(n11591) );
  NAND2_X1 U10933 ( .A1(n8424), .A2(n11591), .ZN(n8517) );
  INV_X1 U10934 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n8513) );
  OR2_X1 U10935 ( .A1(n8870), .A2(n8513), .ZN(n8516) );
  INV_X1 U10936 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n8514) );
  OR2_X1 U10937 ( .A1(n9090), .A2(n8514), .ZN(n8515) );
  NAND4_X1 U10938 ( .A1(n8518), .A2(n8517), .A3(n8516), .A4(n8515), .ZN(n13374) );
  XNOR2_X1 U10939 ( .A(n15370), .B(n13374), .ZN(n11583) );
  INV_X1 U10940 ( .A(n11583), .ZN(n8519) );
  NAND2_X1 U10941 ( .A1(n11582), .A2(n8519), .ZN(n8521) );
  NAND2_X1 U10942 ( .A1(n15370), .A2(n13374), .ZN(n8520) );
  NOR2_X1 U10943 ( .A1(n8593), .A2(P2_IR_REG_10__SCAN_IN), .ZN(n8533) );
  OR2_X1 U10944 ( .A1(n8533), .A2(n8803), .ZN(n8522) );
  XNOR2_X1 U10945 ( .A(n8522), .B(P2_IR_REG_11__SCAN_IN), .ZN(n11491) );
  AOI22_X1 U10946 ( .A1(n8614), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n8636), 
        .B2(n11491), .ZN(n8523) );
  XNOR2_X1 U10947 ( .A(n8540), .B(P2_REG3_REG_11__SCAN_IN), .ZN(n11779) );
  OR2_X1 U10948 ( .A1(n8748), .A2(n11779), .ZN(n8529) );
  NAND2_X1 U10949 ( .A1(n6627), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n8528) );
  INV_X1 U10950 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n8525) );
  OR2_X1 U10951 ( .A1(n8870), .A2(n8525), .ZN(n8527) );
  INV_X1 U10952 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n11758) );
  OR2_X1 U10953 ( .A1(n9090), .A2(n11758), .ZN(n8526) );
  NAND4_X1 U10954 ( .A1(n8529), .A2(n8528), .A3(n8527), .A4(n8526), .ZN(n13373) );
  AND2_X1 U10955 ( .A1(n11783), .A2(n13373), .ZN(n8530) );
  OR2_X1 U10956 ( .A1(n11783), .A2(n13373), .ZN(n8531) );
  NAND2_X1 U10957 ( .A1(n10455), .A2(n9085), .ZN(n8538) );
  NAND2_X1 U10958 ( .A1(n8533), .A2(n8532), .ZN(n8535) );
  NAND2_X1 U10959 ( .A1(n8535), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8534) );
  MUX2_X1 U10960 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8534), .S(
        P2_IR_REG_12__SCAN_IN), .Z(n8536) );
  AOI22_X1 U10961 ( .A1(n8614), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n8636), 
        .B2(n15285), .ZN(n8537) );
  AND2_X1 U10962 ( .A1(P2_REG3_REG_11__SCAN_IN), .A2(P2_REG3_REG_12__SCAN_IN), 
        .ZN(n8539) );
  AOI21_X1 U10963 ( .B1(n8540), .B2(P2_REG3_REG_11__SCAN_IN), .A(
        P2_REG3_REG_12__SCAN_IN), .ZN(n8541) );
  OR2_X1 U10964 ( .A1(n8552), .A2(n8541), .ZN(n15197) );
  OR2_X1 U10965 ( .A1(n8748), .A2(n15197), .ZN(n8546) );
  NAND2_X1 U10966 ( .A1(n6627), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n8545) );
  INV_X1 U10967 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n8542) );
  OR2_X1 U10968 ( .A1(n8870), .A2(n8542), .ZN(n8544) );
  INV_X1 U10969 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n11823) );
  OR2_X1 U10970 ( .A1(n9090), .A2(n11823), .ZN(n8543) );
  NAND4_X1 U10971 ( .A1(n8546), .A2(n8545), .A3(n8544), .A4(n8543), .ZN(n13372) );
  NOR2_X1 U10972 ( .A1(n15194), .A2(n13372), .ZN(n8548) );
  NAND2_X1 U10973 ( .A1(n15194), .A2(n13372), .ZN(n8547) );
  NAND2_X1 U10974 ( .A1(n10492), .A2(n9085), .ZN(n8551) );
  NAND2_X1 U10975 ( .A1(n8559), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8549) );
  XNOR2_X1 U10976 ( .A(n8549), .B(P2_IR_REG_13__SCAN_IN), .ZN(n15297) );
  AOI22_X1 U10977 ( .A1(n8614), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n15297), 
        .B2(n8636), .ZN(n8550) );
  OR2_X1 U10978 ( .A1(n8552), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n8553) );
  NAND2_X1 U10979 ( .A1(n8566), .A2(n8553), .ZN(n11970) );
  OR2_X1 U10980 ( .A1(n8748), .A2(n11970), .ZN(n8557) );
  NAND2_X1 U10981 ( .A1(n6627), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n8556) );
  OR2_X1 U10982 ( .A1(n8870), .A2(n14884), .ZN(n8555) );
  INV_X1 U10983 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n11971) );
  OR2_X1 U10984 ( .A1(n9090), .A2(n11971), .ZN(n8554) );
  NAND4_X1 U10985 ( .A1(n8557), .A2(n8556), .A3(n8555), .A4(n8554), .ZN(n13371) );
  AND2_X1 U10986 ( .A1(n11973), .A2(n13371), .ZN(n8558) );
  OAI22_X1 U10987 ( .A1(n11968), .A2(n8558), .B1(n13371), .B2(n11973), .ZN(
        n12018) );
  OR2_X1 U10988 ( .A1(n10821), .A2(n9107), .ZN(n8564) );
  INV_X1 U10989 ( .A(n8559), .ZN(n8561) );
  INV_X1 U10990 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n8560) );
  NAND2_X1 U10991 ( .A1(n8561), .A2(n8560), .ZN(n8576) );
  NAND2_X1 U10992 ( .A1(n8576), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8562) );
  XNOR2_X1 U10993 ( .A(n8562), .B(P2_IR_REG_14__SCAN_IN), .ZN(n15317) );
  AOI22_X1 U10994 ( .A1(n15317), .A2(n8636), .B1(n8730), .B2(
        P1_DATAO_REG_14__SCAN_IN), .ZN(n8563) );
  INV_X1 U10995 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n8565) );
  NAND2_X1 U10996 ( .A1(n8566), .A2(n8565), .ZN(n8567) );
  NAND2_X1 U10997 ( .A1(n8581), .A2(n8567), .ZN(n14847) );
  OR2_X1 U10998 ( .A1(n8748), .A2(n14847), .ZN(n8572) );
  NAND2_X1 U10999 ( .A1(n6627), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n8571) );
  INV_X1 U11000 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n8568) );
  OR2_X1 U11001 ( .A1(n8870), .A2(n8568), .ZN(n8570) );
  INV_X1 U11002 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n12022) );
  OR2_X1 U11003 ( .A1(n9090), .A2(n12022), .ZN(n8569) );
  NAND4_X1 U11004 ( .A1(n8572), .A2(n8571), .A3(n8570), .A4(n8569), .ZN(n13370) );
  NOR2_X1 U11005 ( .A1(n14845), .A2(n13370), .ZN(n8573) );
  NAND2_X1 U11006 ( .A1(n14845), .A2(n13370), .ZN(n8574) );
  NAND2_X1 U11007 ( .A1(n11069), .A2(n9085), .ZN(n8580) );
  OAI21_X1 U11008 ( .B1(n8576), .B2(P2_IR_REG_14__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8577) );
  XNOR2_X1 U11009 ( .A(n8577), .B(P2_IR_REG_15__SCAN_IN), .ZN(n11604) );
  NOR2_X1 U11010 ( .A1(n8590), .A2(n11168), .ZN(n8578) );
  AOI21_X1 U11011 ( .B1(n11604), .B2(n8636), .A(n8578), .ZN(n8579) );
  AND2_X1 U11012 ( .A1(n8581), .A2(n11503), .ZN(n8582) );
  OR2_X1 U11013 ( .A1(n8600), .A2(n8582), .ZN(n13639) );
  INV_X1 U11014 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n8583) );
  OR2_X1 U11015 ( .A1(n8870), .A2(n8583), .ZN(n8586) );
  INV_X1 U11016 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n8584) );
  OR2_X1 U11017 ( .A1(n9090), .A2(n8584), .ZN(n8585) );
  AND2_X1 U11018 ( .A1(n8586), .A2(n8585), .ZN(n8588) );
  NAND2_X1 U11019 ( .A1(n6627), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n8587) );
  OAI211_X1 U11020 ( .C1(n13639), .C2(n8748), .A(n8588), .B(n8587), .ZN(n13369) );
  INV_X1 U11021 ( .A(n13369), .ZN(n12160) );
  XNOR2_X1 U11022 ( .A(n13642), .B(n12160), .ZN(n12141) );
  OR2_X1 U11023 ( .A1(n13642), .A2(n13369), .ZN(n8589) );
  NAND2_X1 U11024 ( .A1(n11237), .A2(n9085), .ZN(n8599) );
  OAI21_X1 U11025 ( .B1(n8593), .B2(n8592), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n8595) );
  MUX2_X1 U11026 ( .A(n8595), .B(P2_IR_REG_31__SCAN_IN), .S(n8594), .Z(n8597)
         );
  INV_X1 U11027 ( .A(n8596), .ZN(n8611) );
  NAND2_X1 U11028 ( .A1(n8597), .A2(n8611), .ZN(n11880) );
  AOI22_X1 U11029 ( .A1(n8730), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n8636), 
        .B2(n11883), .ZN(n8598) );
  INV_X1 U11030 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n11607) );
  NAND2_X1 U11031 ( .A1(n8600), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8618) );
  INV_X1 U11032 ( .A(n8600), .ZN(n8602) );
  INV_X1 U11033 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n8601) );
  NAND2_X1 U11034 ( .A1(n8602), .A2(n8601), .ZN(n8603) );
  NAND2_X1 U11035 ( .A1(n8618), .A2(n8603), .ZN(n14856) );
  OR2_X1 U11036 ( .A1(n14856), .A2(n8748), .ZN(n8605) );
  AOI22_X1 U11037 ( .A1(n6627), .A2(P2_REG1_REG_16__SCAN_IN), .B1(n8389), .B2(
        P2_REG0_REG_16__SCAN_IN), .ZN(n8604) );
  OAI211_X1 U11038 ( .C1(n6626), .C2(n11607), .A(n8605), .B(n8604), .ZN(n13368) );
  XNOR2_X1 U11039 ( .A(n14853), .B(n13368), .ZN(n12158) );
  NAND2_X1 U11040 ( .A1(n14853), .A2(n13368), .ZN(n8606) );
  NAND2_X1 U11041 ( .A1(n11285), .A2(n9085), .ZN(n8616) );
  NAND2_X1 U11042 ( .A1(n8611), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8612) );
  MUX2_X1 U11043 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8612), .S(
        P2_IR_REG_17__SCAN_IN), .Z(n8613) );
  AND2_X1 U11044 ( .A1(n8610), .A2(n8613), .ZN(n13407) );
  AOI22_X1 U11045 ( .A1(n8614), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n8636), 
        .B2(n13407), .ZN(n8615) );
  INV_X1 U11046 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8622) );
  INV_X1 U11047 ( .A(n8618), .ZN(n8617) );
  NAND2_X1 U11048 ( .A1(n8617), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n8628) );
  INV_X1 U11049 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n13293) );
  NAND2_X1 U11050 ( .A1(n8618), .A2(n13293), .ZN(n8619) );
  NAND2_X1 U11051 ( .A1(n8628), .A2(n8619), .ZN(n13626) );
  OR2_X1 U11052 ( .A1(n13626), .A2(n8748), .ZN(n8621) );
  AOI22_X1 U11053 ( .A1(n6627), .A2(P2_REG1_REG_17__SCAN_IN), .B1(n8389), .B2(
        P2_REG0_REG_17__SCAN_IN), .ZN(n8620) );
  OAI211_X1 U11054 ( .C1(n6626), .C2(n8622), .A(n8621), .B(n8620), .ZN(n13367)
         );
  XNOR2_X1 U11055 ( .A(n13630), .B(n13367), .ZN(n13628) );
  INV_X1 U11056 ( .A(n13628), .ZN(n13620) );
  NAND2_X1 U11057 ( .A1(n13630), .A2(n13367), .ZN(n8623) );
  NAND2_X1 U11058 ( .A1(n11430), .A2(n9085), .ZN(n8626) );
  NAND2_X1 U11059 ( .A1(n8610), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8624) );
  XNOR2_X1 U11060 ( .A(n8624), .B(P2_IR_REG_18__SCAN_IN), .ZN(n13415) );
  AOI22_X1 U11061 ( .A1(n8730), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n8636), 
        .B2(n13415), .ZN(n8625) );
  INV_X1 U11062 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n8627) );
  NAND2_X1 U11063 ( .A1(n8628), .A2(n8627), .ZN(n8629) );
  AND2_X1 U11064 ( .A1(n8639), .A2(n8629), .ZN(n13608) );
  NAND2_X1 U11065 ( .A1(n13608), .A2(n8424), .ZN(n8634) );
  INV_X1 U11066 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n13742) );
  NAND2_X1 U11067 ( .A1(n8690), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n8631) );
  NAND2_X1 U11068 ( .A1(n8389), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n8630) );
  OAI211_X1 U11069 ( .C1(n8467), .C2(n13742), .A(n8631), .B(n8630), .ZN(n8632)
         );
  INV_X1 U11070 ( .A(n8632), .ZN(n8633) );
  NAND2_X1 U11071 ( .A1(n8634), .A2(n8633), .ZN(n13366) );
  INV_X1 U11072 ( .A(n13366), .ZN(n13292) );
  XNOR2_X1 U11073 ( .A(n13609), .B(n13292), .ZN(n13595) );
  INV_X1 U11074 ( .A(n13595), .ZN(n13597) );
  NAND2_X1 U11075 ( .A1(n11530), .A2(n9085), .ZN(n8638) );
  OR2_X1 U11076 ( .A1(n8785), .A2(n8803), .ZN(n8635) );
  XNOR2_X2 U11077 ( .A(n8635), .B(P2_IR_REG_19__SCAN_IN), .ZN(n13429) );
  AOI22_X1 U11078 ( .A1(n8730), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n13429), 
        .B2(n8636), .ZN(n8637) );
  INV_X1 U11079 ( .A(n8652), .ZN(n8654) );
  NAND2_X1 U11080 ( .A1(n8639), .A2(n10119), .ZN(n8640) );
  NAND2_X1 U11081 ( .A1(n8654), .A2(n8640), .ZN(n13584) );
  OR2_X1 U11082 ( .A1(n13584), .A2(n8748), .ZN(n8646) );
  INV_X1 U11083 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n8643) );
  NAND2_X1 U11084 ( .A1(n8389), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n8642) );
  NAND2_X1 U11085 ( .A1(n8690), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n8641) );
  OAI211_X1 U11086 ( .C1(n8643), .C2(n8467), .A(n8642), .B(n8641), .ZN(n8644)
         );
  INV_X1 U11087 ( .A(n8644), .ZN(n8645) );
  NAND2_X1 U11088 ( .A1(n8646), .A2(n8645), .ZN(n13365) );
  NAND2_X1 U11089 ( .A1(n13731), .A2(n13365), .ZN(n8647) );
  NAND2_X1 U11090 ( .A1(n13582), .A2(n8647), .ZN(n8649) );
  OR2_X1 U11091 ( .A1(n13731), .A2(n13365), .ZN(n8648) );
  NAND2_X1 U11092 ( .A1(n12312), .A2(n9085), .ZN(n8651) );
  NAND2_X1 U11093 ( .A1(n8730), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n8650) );
  NAND2_X2 U11094 ( .A1(n8651), .A2(n8650), .ZN(n13726) );
  INV_X1 U11095 ( .A(n8665), .ZN(n8666) );
  INV_X1 U11096 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n8653) );
  NAND2_X1 U11097 ( .A1(n8654), .A2(n8653), .ZN(n8655) );
  AND2_X1 U11098 ( .A1(n8666), .A2(n8655), .ZN(n13570) );
  NAND2_X1 U11099 ( .A1(n13570), .A2(n8424), .ZN(n8660) );
  INV_X1 U11100 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n10078) );
  NAND2_X1 U11101 ( .A1(n6627), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n8657) );
  NAND2_X1 U11102 ( .A1(n8690), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n8656) );
  OAI211_X1 U11103 ( .C1(n8870), .C2(n10078), .A(n8657), .B(n8656), .ZN(n8658)
         );
  INV_X1 U11104 ( .A(n8658), .ZN(n8659) );
  NAND2_X1 U11105 ( .A1(n8660), .A2(n8659), .ZN(n13364) );
  NOR2_X1 U11106 ( .A1(n13726), .A2(n13364), .ZN(n8661) );
  NAND2_X1 U11107 ( .A1(n13726), .A2(n13364), .ZN(n8662) );
  NAND2_X1 U11108 ( .A1(n11828), .A2(n9085), .ZN(n8664) );
  NAND2_X1 U11109 ( .A1(n8730), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n8663) );
  INV_X1 U11110 ( .A(n8678), .ZN(n8668) );
  INV_X1 U11111 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n13272) );
  NAND2_X1 U11112 ( .A1(n8666), .A2(n13272), .ZN(n8667) );
  NAND2_X1 U11113 ( .A1(n8668), .A2(n8667), .ZN(n13558) );
  OR2_X1 U11114 ( .A1(n13558), .A2(n8748), .ZN(n8673) );
  INV_X1 U11115 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n13723) );
  NAND2_X1 U11116 ( .A1(n8690), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n8670) );
  NAND2_X1 U11117 ( .A1(n8389), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n8669) );
  OAI211_X1 U11118 ( .C1(n8467), .C2(n13723), .A(n8670), .B(n8669), .ZN(n8671)
         );
  INV_X1 U11119 ( .A(n8671), .ZN(n8672) );
  NAND2_X1 U11120 ( .A1(n8673), .A2(n8672), .ZN(n13363) );
  INV_X1 U11121 ( .A(n13363), .ZN(n8852) );
  XNOR2_X1 U11122 ( .A(n13557), .B(n8852), .ZN(n13548) );
  INV_X1 U11123 ( .A(n13548), .ZN(n13553) );
  XNOR2_X1 U11124 ( .A(n8675), .B(n8674), .ZN(n12169) );
  NAND2_X1 U11125 ( .A1(n12169), .A2(n9085), .ZN(n8677) );
  NAND2_X1 U11126 ( .A1(n8730), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n8676) );
  NOR2_X1 U11127 ( .A1(n8678), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n8679) );
  OR2_X1 U11128 ( .A1(n8688), .A2(n8679), .ZN(n13319) );
  INV_X1 U11129 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n8682) );
  NAND2_X1 U11130 ( .A1(n8690), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n8681) );
  NAND2_X1 U11131 ( .A1(n8389), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n8680) );
  OAI211_X1 U11132 ( .C1(n8467), .C2(n8682), .A(n8681), .B(n8680), .ZN(n8683)
         );
  INV_X1 U11133 ( .A(n8683), .ZN(n8684) );
  OAI21_X1 U11134 ( .B1(n13319), .B2(n8748), .A(n8684), .ZN(n13362) );
  INV_X1 U11135 ( .A(n13362), .ZN(n13271) );
  XNOR2_X1 U11136 ( .A(n13716), .B(n13271), .ZN(n13533) );
  INV_X1 U11137 ( .A(n13533), .ZN(n13541) );
  NAND2_X1 U11138 ( .A1(n13716), .A2(n13362), .ZN(n8685) );
  NAND2_X1 U11139 ( .A1(n11999), .A2(n9085), .ZN(n8687) );
  NAND2_X1 U11140 ( .A1(n8730), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n8686) );
  OR2_X1 U11141 ( .A1(n8688), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n8689) );
  NAND2_X1 U11142 ( .A1(n8688), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n8698) );
  AND2_X1 U11143 ( .A1(n8689), .A2(n8698), .ZN(n13523) );
  NAND2_X1 U11144 ( .A1(n13523), .A2(n8424), .ZN(n8695) );
  INV_X1 U11145 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n10182) );
  NAND2_X1 U11146 ( .A1(n6627), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n8692) );
  NAND2_X1 U11147 ( .A1(n8690), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n8691) );
  OAI211_X1 U11148 ( .C1(n8870), .C2(n10182), .A(n8692), .B(n8691), .ZN(n8693)
         );
  INV_X1 U11149 ( .A(n8693), .ZN(n8694) );
  NAND2_X1 U11150 ( .A1(n8695), .A2(n8694), .ZN(n13361) );
  NAND2_X1 U11151 ( .A1(n12133), .A2(n9085), .ZN(n8697) );
  NAND2_X1 U11152 ( .A1(n8730), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n8696) );
  OAI21_X1 U11153 ( .B1(P2_REG3_REG_24__SCAN_IN), .B2(n8699), .A(n8719), .ZN(
        n13512) );
  OR2_X1 U11154 ( .A1(n8748), .A2(n13512), .ZN(n8705) );
  NAND2_X1 U11155 ( .A1(n6627), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n8704) );
  INV_X1 U11156 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n8700) );
  OR2_X1 U11157 ( .A1(n8870), .A2(n8700), .ZN(n8703) );
  INV_X1 U11158 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n8701) );
  OR2_X1 U11159 ( .A1(n9090), .A2(n8701), .ZN(n8702) );
  NAND4_X1 U11160 ( .A1(n8705), .A2(n8704), .A3(n8703), .A4(n8702), .ZN(n13360) );
  INV_X1 U11161 ( .A(n13360), .ZN(n13281) );
  NAND2_X1 U11162 ( .A1(n13802), .A2(n9085), .ZN(n8707) );
  NAND2_X1 U11163 ( .A1(n8730), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n8706) );
  NAND2_X1 U11164 ( .A1(n6627), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n8713) );
  XNOR2_X1 U11165 ( .A(n8719), .B(P2_REG3_REG_25__SCAN_IN), .ZN(n13496) );
  NAND2_X1 U11166 ( .A1(n8424), .A2(n13496), .ZN(n8712) );
  INV_X1 U11167 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n8708) );
  OR2_X1 U11168 ( .A1(n8870), .A2(n8708), .ZN(n8711) );
  INV_X1 U11169 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n8709) );
  OR2_X1 U11170 ( .A1(n9090), .A2(n8709), .ZN(n8710) );
  NAND4_X1 U11171 ( .A1(n8713), .A2(n8712), .A3(n8711), .A4(n8710), .ZN(n13359) );
  NAND2_X1 U11172 ( .A1(n13698), .A2(n13359), .ZN(n8714) );
  NAND2_X1 U11173 ( .A1(n8715), .A2(n8714), .ZN(n13478) );
  NAND2_X1 U11174 ( .A1(n13799), .A2(n9085), .ZN(n8717) );
  NAND2_X1 U11175 ( .A1(n8730), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n8716) );
  INV_X1 U11176 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n13282) );
  INV_X1 U11177 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n8718) );
  OAI21_X1 U11178 ( .B1(n8719), .B2(n13282), .A(n8718), .ZN(n8722) );
  INV_X1 U11179 ( .A(n8719), .ZN(n8721) );
  AND2_X1 U11180 ( .A1(P2_REG3_REG_26__SCAN_IN), .A2(P2_REG3_REG_25__SCAN_IN), 
        .ZN(n8720) );
  NAND2_X1 U11181 ( .A1(n8721), .A2(n8720), .ZN(n8734) );
  NAND2_X1 U11182 ( .A1(n8722), .A2(n8734), .ZN(n13338) );
  OR2_X1 U11183 ( .A1(n8748), .A2(n13338), .ZN(n8728) );
  NAND2_X1 U11184 ( .A1(n6627), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n8727) );
  INV_X1 U11185 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n8723) );
  OR2_X1 U11186 ( .A1(n8870), .A2(n8723), .ZN(n8726) );
  INV_X1 U11187 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n8724) );
  OR2_X1 U11188 ( .A1(n6626), .A2(n8724), .ZN(n8725) );
  NAND4_X1 U11189 ( .A1(n8728), .A2(n8727), .A3(n8726), .A4(n8725), .ZN(n13358) );
  AND2_X1 U11190 ( .A1(n13694), .A2(n13358), .ZN(n8729) );
  NAND2_X1 U11191 ( .A1(n13796), .A2(n9085), .ZN(n8732) );
  NAND2_X1 U11192 ( .A1(n8730), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n8731) );
  INV_X1 U11193 ( .A(n8734), .ZN(n8733) );
  NAND2_X1 U11194 ( .A1(n8733), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n8746) );
  INV_X1 U11195 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n13229) );
  NAND2_X1 U11196 ( .A1(n8734), .A2(n13229), .ZN(n8735) );
  NAND2_X1 U11197 ( .A1(n8746), .A2(n8735), .ZN(n13469) );
  OR2_X1 U11198 ( .A1(n8748), .A2(n13469), .ZN(n8741) );
  NAND2_X1 U11199 ( .A1(n6627), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n8740) );
  INV_X1 U11200 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n8736) );
  OR2_X1 U11201 ( .A1(n8870), .A2(n8736), .ZN(n8739) );
  INV_X1 U11202 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n8737) );
  OR2_X1 U11203 ( .A1(n6626), .A2(n8737), .ZN(n8738) );
  NAND4_X1 U11204 ( .A1(n8741), .A2(n8740), .A3(n8739), .A4(n8738), .ZN(n13357) );
  XNOR2_X1 U11205 ( .A(n13688), .B(n13357), .ZN(n13474) );
  OR2_X2 U11206 ( .A1(n13475), .A2(n13474), .ZN(n13686) );
  NAND2_X1 U11207 ( .A1(n13688), .A2(n13357), .ZN(n8742) );
  NAND2_X1 U11208 ( .A1(n13793), .A2(n9085), .ZN(n8744) );
  NAND2_X1 U11209 ( .A1(n8730), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n8743) );
  NAND2_X1 U11210 ( .A1(n6627), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n8752) );
  INV_X1 U11211 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n8745) );
  OR2_X1 U11212 ( .A1(n8870), .A2(n8745), .ZN(n8751) );
  INV_X1 U11213 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n13262) );
  NAND2_X1 U11214 ( .A1(n8746), .A2(n13262), .ZN(n8747) );
  NAND2_X1 U11215 ( .A1(n8757), .A2(n8747), .ZN(n13449) );
  OR2_X1 U11216 ( .A1(n8748), .A2(n13449), .ZN(n8750) );
  INV_X1 U11217 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n13450) );
  OR2_X1 U11218 ( .A1(n6626), .A2(n13450), .ZN(n8749) );
  NAND2_X1 U11219 ( .A1(n13455), .A2(n11029), .ZN(n8754) );
  OR2_X1 U11220 ( .A1(n13455), .A2(n11029), .ZN(n8753) );
  NAND2_X1 U11221 ( .A1(n8754), .A2(n8753), .ZN(n9161) );
  NAND2_X1 U11222 ( .A1(n13447), .A2(n13456), .ZN(n13448) );
  NAND2_X1 U11223 ( .A1(n13789), .A2(n9085), .ZN(n8756) );
  NAND2_X1 U11224 ( .A1(n8730), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n8755) );
  NAND2_X1 U11225 ( .A1(n6627), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n8763) );
  INV_X1 U11226 ( .A(n8757), .ZN(n8878) );
  NAND2_X1 U11227 ( .A1(n8424), .A2(n8878), .ZN(n8762) );
  INV_X1 U11228 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n8758) );
  OR2_X1 U11229 ( .A1(n8870), .A2(n8758), .ZN(n8761) );
  INV_X1 U11230 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n8759) );
  OR2_X1 U11231 ( .A1(n6626), .A2(n8759), .ZN(n8760) );
  NAND4_X1 U11232 ( .A1(n8763), .A2(n8762), .A3(n8761), .A4(n8760), .ZN(n13356) );
  INV_X1 U11233 ( .A(n13356), .ZN(n8764) );
  XNOR2_X1 U11234 ( .A(n13676), .B(n8764), .ZN(n9163) );
  NOR4_X1 U11235 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_16__SCAN_IN), .A3(
        P2_D_REG_17__SCAN_IN), .A4(P2_D_REG_18__SCAN_IN), .ZN(n8769) );
  NOR4_X1 U11236 ( .A1(P2_D_REG_12__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_11__SCAN_IN), .A4(P2_D_REG_13__SCAN_IN), .ZN(n8768) );
  NOR4_X1 U11237 ( .A1(P2_D_REG_24__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_27__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n8767) );
  NOR4_X1 U11238 ( .A1(P2_D_REG_19__SCAN_IN), .A2(P2_D_REG_20__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_22__SCAN_IN), .ZN(n8766) );
  NAND4_X1 U11239 ( .A1(n8769), .A2(n8768), .A3(n8767), .A4(n8766), .ZN(n8794)
         );
  NOR2_X1 U11240 ( .A1(P2_D_REG_14__SCAN_IN), .A2(P2_D_REG_28__SCAN_IN), .ZN(
        n8773) );
  NOR4_X1 U11241 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_23__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n8772) );
  NOR4_X1 U11242 ( .A1(P2_D_REG_6__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_8__SCAN_IN), .A4(P2_D_REG_9__SCAN_IN), .ZN(n8771) );
  NOR4_X1 U11243 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_4__SCAN_IN), .A4(P2_D_REG_5__SCAN_IN), .ZN(n8770) );
  NAND4_X1 U11244 ( .A1(n8773), .A2(n8772), .A3(n8771), .A4(n8770), .ZN(n8793)
         );
  NOR2_X1 U11245 ( .A1(n8610), .A2(n8774), .ZN(n8779) );
  NAND2_X1 U11246 ( .A1(n8779), .A2(n8775), .ZN(n8782) );
  NAND2_X1 U11247 ( .A1(n8782), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8776) );
  MUX2_X1 U11248 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8776), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n8777) );
  INV_X1 U11249 ( .A(n13801), .ZN(n8792) );
  INV_X1 U11250 ( .A(n8779), .ZN(n8780) );
  NAND2_X1 U11251 ( .A1(n8780), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8781) );
  MUX2_X1 U11252 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8781), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n8783) );
  NAND2_X1 U11253 ( .A1(n8783), .A2(n8782), .ZN(n13803) );
  AND2_X2 U11254 ( .A1(n8785), .A2(n8784), .ZN(n8802) );
  NAND2_X1 U11255 ( .A1(n8796), .A2(n8795), .ZN(n8787) );
  INV_X1 U11256 ( .A(P2_B_REG_SCAN_IN), .ZN(n10214) );
  XOR2_X1 U11257 ( .A(n12136), .B(n10214), .Z(n8790) );
  NAND2_X1 U11258 ( .A1(n13803), .A2(n8790), .ZN(n8791) );
  OAI21_X1 U11259 ( .B1(n8794), .B2(n8793), .A(n15337), .ZN(n10626) );
  NAND2_X1 U11260 ( .A1(n10626), .A2(n15349), .ZN(n10544) );
  NAND2_X1 U11261 ( .A1(n12136), .A2(n13801), .ZN(n8798) );
  INV_X1 U11262 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n15344) );
  NAND2_X1 U11263 ( .A1(n15337), .A2(n15344), .ZN(n8797) );
  NAND2_X1 U11264 ( .A1(n8798), .A2(n8797), .ZN(n15345) );
  XNOR2_X2 U11265 ( .A(n8800), .B(P2_IR_REG_22__SCAN_IN), .ZN(n8877) );
  NAND2_X1 U11266 ( .A1(n8877), .A2(n9168), .ZN(n10291) );
  NAND2_X1 U11267 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n8786), .ZN(n8804) );
  NAND2_X2 U11268 ( .A1(n8807), .A2(n8806), .ZN(n12326) );
  NAND2_X1 U11269 ( .A1(n12326), .A2(n11531), .ZN(n9173) );
  OR2_X1 U11270 ( .A1(n10291), .A2(n10623), .ZN(n10629) );
  NAND2_X1 U11271 ( .A1(n15345), .A2(n10629), .ZN(n8808) );
  INV_X1 U11272 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n15347) );
  NAND2_X1 U11273 ( .A1(n15337), .A2(n15347), .ZN(n8810) );
  NAND2_X1 U11274 ( .A1(n13801), .A2(n13803), .ZN(n8809) );
  NAND2_X1 U11275 ( .A1(n10605), .A2(n10619), .ZN(n8812) );
  NAND2_X1 U11276 ( .A1(n8890), .A2(n11829), .ZN(n10627) );
  INV_X1 U11277 ( .A(n10627), .ZN(n8811) );
  NAND2_X2 U11278 ( .A1(n8813), .A2(n12326), .ZN(n9791) );
  OAI21_X2 U11279 ( .B1(n9136), .B2(n8814), .A(n11531), .ZN(n8815) );
  NAND2_X2 U11280 ( .A1(n8815), .A2(n9791), .ZN(n10652) );
  BUF_X4 U11281 ( .A(n10652), .Z(n13255) );
  INV_X2 U11282 ( .A(n13255), .ZN(n13213) );
  AND2_X1 U11283 ( .A1(n8816), .A2(n11531), .ZN(n8817) );
  NAND2_X1 U11284 ( .A1(n9798), .A2(n10727), .ZN(n10641) );
  INV_X1 U11285 ( .A(n10641), .ZN(n9797) );
  NAND2_X1 U11286 ( .A1(n9797), .A2(n9796), .ZN(n9795) );
  NAND2_X1 U11287 ( .A1(n10649), .A2(n8899), .ZN(n8818) );
  NAND2_X1 U11288 ( .A1(n11203), .A2(n10650), .ZN(n8819) );
  INV_X1 U11289 ( .A(n10760), .ZN(n10763) );
  NAND2_X1 U11290 ( .A1(n10764), .A2(n10763), .ZN(n8822) );
  NAND2_X1 U11291 ( .A1(n10843), .A2(n10599), .ZN(n8821) );
  NAND2_X1 U11292 ( .A1(n8822), .A2(n8821), .ZN(n10962) );
  NAND2_X1 U11293 ( .A1(n10962), .A2(n9145), .ZN(n8824) );
  NAND2_X1 U11294 ( .A1(n10965), .A2(n10927), .ZN(n8823) );
  NAND2_X1 U11295 ( .A1(n8824), .A2(n8823), .ZN(n11119) );
  NAND2_X1 U11296 ( .A1(n11119), .A2(n9147), .ZN(n8827) );
  INV_X1 U11297 ( .A(n13378), .ZN(n8825) );
  NAND2_X1 U11298 ( .A1(n11123), .A2(n8825), .ZN(n8826) );
  AND2_X1 U11299 ( .A1(n15323), .A2(n10928), .ZN(n8828) );
  NAND2_X1 U11300 ( .A1(n11455), .A2(n11453), .ZN(n8830) );
  INV_X1 U11301 ( .A(n13376), .ZN(n11426) );
  OR2_X1 U11302 ( .A1(n15364), .A2(n11426), .ZN(n8829) );
  NAND2_X1 U11303 ( .A1(n8830), .A2(n8829), .ZN(n11560) );
  NAND2_X1 U11304 ( .A1(n11560), .A2(n9149), .ZN(n8833) );
  INV_X1 U11305 ( .A(n13375), .ZN(n8831) );
  OR2_X1 U11306 ( .A1(n11746), .A2(n8831), .ZN(n8832) );
  NAND2_X1 U11307 ( .A1(n8833), .A2(n8832), .ZN(n11584) );
  NAND2_X1 U11308 ( .A1(n11584), .A2(n11583), .ZN(n8835) );
  INV_X1 U11309 ( .A(n13374), .ZN(n11425) );
  OR2_X1 U11310 ( .A1(n15370), .A2(n11425), .ZN(n8834) );
  INV_X1 U11311 ( .A(n13373), .ZN(n8836) );
  XNOR2_X1 U11312 ( .A(n11783), .B(n8836), .ZN(n11756) );
  NAND2_X1 U11313 ( .A1(n11783), .A2(n8836), .ZN(n8837) );
  XNOR2_X1 U11314 ( .A(n15194), .B(n13372), .ZN(n9152) );
  INV_X1 U11315 ( .A(n13372), .ZN(n11952) );
  XNOR2_X1 U11316 ( .A(n11973), .B(n13371), .ZN(n11967) );
  NAND2_X1 U11317 ( .A1(n11963), .A2(n11967), .ZN(n8840) );
  INV_X1 U11318 ( .A(n13371), .ZN(n8838) );
  OR2_X1 U11319 ( .A1(n11973), .A2(n8838), .ZN(n8839) );
  INV_X1 U11320 ( .A(n13370), .ZN(n11953) );
  NOR2_X1 U11321 ( .A1(n14845), .A2(n11953), .ZN(n8841) );
  NAND2_X1 U11322 ( .A1(n14845), .A2(n11953), .ZN(n8842) );
  OR2_X1 U11323 ( .A1(n13642), .A2(n12160), .ZN(n8843) );
  NAND2_X1 U11324 ( .A1(n8844), .A2(n8843), .ZN(n12159) );
  NAND2_X1 U11325 ( .A1(n12159), .A2(n12158), .ZN(n12157) );
  INV_X1 U11326 ( .A(n13368), .ZN(n13291) );
  OR2_X1 U11327 ( .A1(n14853), .A2(n13291), .ZN(n8845) );
  INV_X1 U11328 ( .A(n13367), .ZN(n12161) );
  NAND2_X1 U11329 ( .A1(n13630), .A2(n12161), .ZN(n8846) );
  AND2_X1 U11330 ( .A1(n13609), .A2(n13292), .ZN(n8847) );
  INV_X1 U11331 ( .A(n13365), .ZN(n8848) );
  NAND2_X1 U11332 ( .A1(n13731), .A2(n8848), .ZN(n8849) );
  INV_X1 U11333 ( .A(n13726), .ZN(n13572) );
  AND2_X1 U11334 ( .A1(n13557), .A2(n8852), .ZN(n8851) );
  NAND2_X1 U11335 ( .A1(n13534), .A2(n13541), .ZN(n8854) );
  OR2_X1 U11336 ( .A1(n13716), .A2(n13271), .ZN(n8853) );
  INV_X1 U11337 ( .A(n13361), .ZN(n13304) );
  NOR2_X1 U11338 ( .A1(n13524), .A2(n13304), .ZN(n8855) );
  NAND2_X1 U11339 ( .A1(n13703), .A2(n13281), .ZN(n8856) );
  INV_X1 U11340 ( .A(n13359), .ZN(n13302) );
  XNOR2_X1 U11341 ( .A(n13698), .B(n13302), .ZN(n13499) );
  INV_X1 U11342 ( .A(n13499), .ZN(n13491) );
  NAND2_X1 U11343 ( .A1(n13698), .A2(n13302), .ZN(n8858) );
  XNOR2_X1 U11344 ( .A(n13694), .B(n13358), .ZN(n13486) );
  INV_X1 U11345 ( .A(n13358), .ZN(n13280) );
  NAND2_X1 U11346 ( .A1(n13694), .A2(n13280), .ZN(n8859) );
  NAND2_X1 U11347 ( .A1(n13463), .A2(n13474), .ZN(n8863) );
  INV_X1 U11348 ( .A(n13357), .ZN(n8861) );
  NAND2_X1 U11349 ( .A1(n13688), .A2(n8861), .ZN(n8862) );
  OR2_X2 U11350 ( .A1(n13457), .A2(n13456), .ZN(n13459) );
  NAND2_X1 U11351 ( .A1(n8877), .A2(n13429), .ZN(n8865) );
  INV_X1 U11352 ( .A(n12326), .ZN(n9143) );
  NAND2_X1 U11353 ( .A1(n9143), .A2(n9168), .ZN(n9134) );
  INV_X1 U11354 ( .A(n8867), .ZN(n10305) );
  NOR2_X1 U11355 ( .A1(n8868), .A2(n10214), .ZN(n8869) );
  NOR2_X1 U11356 ( .A1(n13301), .A2(n8869), .ZN(n13437) );
  INV_X1 U11357 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n13442) );
  NAND2_X1 U11358 ( .A1(n6627), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n8872) );
  INV_X1 U11359 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n13755) );
  OR2_X1 U11360 ( .A1(n8870), .A2(n13755), .ZN(n8871) );
  OAI211_X1 U11361 ( .C1(n6626), .C2(n13442), .A(n8872), .B(n8871), .ZN(n13355) );
  AOI21_X2 U11362 ( .B1(n8875), .B2(n13661), .A(n8874), .ZN(n13678) );
  INV_X1 U11363 ( .A(n11973), .ZN(n14871) );
  INV_X1 U11364 ( .A(n11746), .ZN(n11743) );
  INV_X1 U11365 ( .A(n11123), .ZN(n11143) );
  NAND2_X1 U11366 ( .A1(n11115), .A2(n11143), .ZN(n11257) );
  OR2_X1 U11367 ( .A1(n11257), .A2(n15323), .ZN(n11462) );
  INV_X1 U11368 ( .A(n13731), .ZN(n13586) );
  NAND2_X1 U11369 ( .A1(n13606), .A2(n13586), .ZN(n13589) );
  OR2_X2 U11370 ( .A1(n9168), .A2(n8877), .ZN(n10585) );
  INV_X2 U11371 ( .A(n13588), .ZN(n13651) );
  AOI211_X1 U11372 ( .C1(n13676), .C2(n13452), .A(n13651), .B(n13441), .ZN(
        n13675) );
  NAND2_X1 U11373 ( .A1(n10548), .A2(n9143), .ZN(n10621) );
  INV_X1 U11374 ( .A(n13655), .ZN(n15326) );
  AOI22_X1 U11375 ( .A1(n6620), .A2(P2_REG2_REG_29__SCAN_IN), .B1(n8878), .B2(
        n15326), .ZN(n8879) );
  OAI21_X1 U11376 ( .B1(n6880), .B2(n15330), .A(n8879), .ZN(n8880) );
  AOI21_X1 U11377 ( .B1(n13675), .B2(n15324), .A(n8880), .ZN(n8881) );
  NAND2_X1 U11378 ( .A1(n15185), .A2(n15155), .ZN(n14686) );
  NOR2_X1 U11379 ( .A1(n15185), .A2(n8885), .ZN(n8886) );
  NAND2_X1 U11380 ( .A1(n13698), .A2(n6618), .ZN(n8892) );
  NAND2_X1 U11381 ( .A1(n6619), .A2(n13359), .ZN(n8891) );
  NAND2_X1 U11382 ( .A1(n8892), .A2(n8891), .ZN(n9065) );
  NAND2_X1 U11383 ( .A1(n9142), .A2(n8909), .ZN(n8896) );
  INV_X1 U11384 ( .A(n9791), .ZN(n8893) );
  OAI211_X1 U11385 ( .C1(n9791), .C2(n10639), .A(n8910), .B(n13384), .ZN(n8894) );
  NAND3_X1 U11386 ( .A1(n8896), .A2(n8895), .A3(n8894), .ZN(n8903) );
  NAND2_X1 U11387 ( .A1(n8909), .A2(n8899), .ZN(n8898) );
  NAND2_X1 U11388 ( .A1(n8910), .A2(n13383), .ZN(n8897) );
  NAND2_X1 U11389 ( .A1(n8898), .A2(n8897), .ZN(n8904) );
  NAND2_X1 U11390 ( .A1(n8903), .A2(n8904), .ZN(n8902) );
  NAND2_X1 U11391 ( .A1(n8910), .A2(n8899), .ZN(n8900) );
  OAI21_X1 U11392 ( .B1(n9126), .B2(n10649), .A(n8900), .ZN(n8901) );
  NAND2_X1 U11393 ( .A1(n8902), .A2(n8901), .ZN(n8915) );
  INV_X1 U11394 ( .A(n8903), .ZN(n8906) );
  INV_X1 U11395 ( .A(n8904), .ZN(n8905) );
  NAND2_X1 U11396 ( .A1(n8906), .A2(n8905), .ZN(n8914) );
  NAND2_X1 U11397 ( .A1(n8910), .A2(n13382), .ZN(n8908) );
  INV_X1 U11398 ( .A(n8916), .ZN(n8912) );
  INV_X1 U11399 ( .A(n8917), .ZN(n8911) );
  NAND2_X1 U11400 ( .A1(n8912), .A2(n8911), .ZN(n8913) );
  NAND3_X1 U11401 ( .A1(n8915), .A2(n8914), .A3(n8913), .ZN(n8919) );
  NAND2_X1 U11402 ( .A1(n8917), .A2(n8916), .ZN(n8918) );
  NAND2_X1 U11403 ( .A1(n8919), .A2(n8918), .ZN(n8925) );
  OR2_X1 U11404 ( .A1(n9126), .A2(n10736), .ZN(n8921) );
  NAND2_X1 U11405 ( .A1(n6619), .A2(n13381), .ZN(n8920) );
  NAND2_X1 U11406 ( .A1(n8921), .A2(n8920), .ZN(n8926) );
  NAND2_X1 U11407 ( .A1(n8925), .A2(n8926), .ZN(n8924) );
  NAND2_X1 U11408 ( .A1(n6619), .A2(n11203), .ZN(n8922) );
  OAI21_X1 U11409 ( .B1(n9126), .B2(n10650), .A(n8922), .ZN(n8923) );
  NAND2_X1 U11410 ( .A1(n8924), .A2(n8923), .ZN(n8930) );
  INV_X1 U11411 ( .A(n8925), .ZN(n8928) );
  INV_X1 U11412 ( .A(n8926), .ZN(n8927) );
  NAND2_X1 U11413 ( .A1(n8928), .A2(n8927), .ZN(n8929) );
  NAND2_X1 U11414 ( .A1(n8930), .A2(n8929), .ZN(n8935) );
  NAND2_X1 U11415 ( .A1(n10843), .A2(n6619), .ZN(n8932) );
  NAND2_X1 U11416 ( .A1(n6618), .A2(n13380), .ZN(n8931) );
  NAND2_X1 U11417 ( .A1(n8932), .A2(n8931), .ZN(n8934) );
  AOI22_X1 U11418 ( .A1(n10843), .A2(n6618), .B1(n6619), .B2(n13380), .ZN(
        n8933) );
  NAND2_X1 U11419 ( .A1(n10965), .A2(n6618), .ZN(n8938) );
  NAND2_X1 U11420 ( .A1(n6619), .A2(n13379), .ZN(n8937) );
  NAND2_X1 U11421 ( .A1(n10965), .A2(n6619), .ZN(n8940) );
  NAND2_X1 U11422 ( .A1(n6618), .A2(n13379), .ZN(n8939) );
  NAND2_X1 U11423 ( .A1(n8940), .A2(n8939), .ZN(n8941) );
  NAND2_X1 U11424 ( .A1(n11123), .A2(n6619), .ZN(n8943) );
  NAND2_X1 U11425 ( .A1(n6618), .A2(n13378), .ZN(n8942) );
  NAND2_X1 U11426 ( .A1(n8943), .A2(n8942), .ZN(n8946) );
  AOI22_X1 U11427 ( .A1(n11123), .A2(n6618), .B1(n6619), .B2(n13378), .ZN(
        n8944) );
  INV_X1 U11428 ( .A(n8945), .ZN(n8948) );
  NAND2_X1 U11429 ( .A1(n15323), .A2(n6618), .ZN(n8950) );
  NAND2_X1 U11430 ( .A1(n6619), .A2(n13377), .ZN(n8949) );
  NAND2_X1 U11431 ( .A1(n8950), .A2(n8949), .ZN(n8954) );
  NAND2_X1 U11432 ( .A1(n15323), .A2(n6619), .ZN(n8952) );
  NAND2_X1 U11433 ( .A1(n6618), .A2(n13377), .ZN(n8951) );
  NAND2_X1 U11434 ( .A1(n8952), .A2(n8951), .ZN(n8953) );
  NAND2_X1 U11435 ( .A1(n15364), .A2(n6619), .ZN(n8957) );
  NAND2_X1 U11436 ( .A1(n6618), .A2(n13376), .ZN(n8956) );
  NAND2_X1 U11437 ( .A1(n8957), .A2(n8956), .ZN(n8959) );
  AOI22_X1 U11438 ( .A1(n15364), .A2(n9097), .B1(n6619), .B2(n13376), .ZN(
        n8958) );
  NOR2_X1 U11439 ( .A1(n8960), .A2(n8959), .ZN(n8961) );
  INV_X1 U11440 ( .A(n9126), .ZN(n9097) );
  NAND2_X1 U11441 ( .A1(n11746), .A2(n9097), .ZN(n8964) );
  NAND2_X1 U11442 ( .A1(n6619), .A2(n13375), .ZN(n8963) );
  NAND2_X1 U11443 ( .A1(n8964), .A2(n8963), .ZN(n8967) );
  AOI22_X1 U11444 ( .A1(n11746), .A2(n6619), .B1(n9097), .B2(n13375), .ZN(
        n8965) );
  AOI21_X1 U11445 ( .B1(n8968), .B2(n8967), .A(n8965), .ZN(n8966) );
  INV_X1 U11446 ( .A(n8966), .ZN(n8969) );
  NAND2_X1 U11447 ( .A1(n15370), .A2(n6619), .ZN(n8971) );
  NAND2_X1 U11448 ( .A1(n9097), .A2(n13374), .ZN(n8970) );
  NAND2_X1 U11449 ( .A1(n8971), .A2(n8970), .ZN(n8973) );
  INV_X1 U11450 ( .A(n8973), .ZN(n8972) );
  NAND2_X1 U11451 ( .A1(n15370), .A2(n6618), .ZN(n8976) );
  NAND2_X1 U11452 ( .A1(n6619), .A2(n13374), .ZN(n8975) );
  NAND2_X1 U11453 ( .A1(n8976), .A2(n8975), .ZN(n8977) );
  NAND2_X1 U11454 ( .A1(n11783), .A2(n9097), .ZN(n8979) );
  NAND2_X1 U11455 ( .A1(n6619), .A2(n13373), .ZN(n8978) );
  AOI22_X1 U11456 ( .A1(n11783), .A2(n6619), .B1(n9097), .B2(n13373), .ZN(
        n8980) );
  NAND2_X1 U11457 ( .A1(n15194), .A2(n6619), .ZN(n8982) );
  NAND2_X1 U11458 ( .A1(n6618), .A2(n13372), .ZN(n8981) );
  NAND2_X1 U11459 ( .A1(n8982), .A2(n8981), .ZN(n8983) );
  NAND2_X1 U11460 ( .A1(n8984), .A2(n8983), .ZN(n8987) );
  NAND2_X1 U11461 ( .A1(n15194), .A2(n6618), .ZN(n8985) );
  OAI21_X1 U11462 ( .B1(n9101), .B2(n11952), .A(n8985), .ZN(n8986) );
  NAND2_X1 U11463 ( .A1(n8987), .A2(n8986), .ZN(n8988) );
  NAND2_X1 U11464 ( .A1(n11973), .A2(n9097), .ZN(n8990) );
  NAND2_X1 U11465 ( .A1(n6619), .A2(n13371), .ZN(n8989) );
  AOI22_X1 U11466 ( .A1(n11973), .A2(n6619), .B1(n9097), .B2(n13371), .ZN(
        n8991) );
  INV_X1 U11467 ( .A(n8991), .ZN(n8992) );
  NAND2_X1 U11468 ( .A1(n14845), .A2(n6619), .ZN(n8994) );
  NAND2_X1 U11469 ( .A1(n6618), .A2(n13370), .ZN(n8993) );
  NAND2_X1 U11470 ( .A1(n14845), .A2(n9097), .ZN(n8995) );
  OAI21_X1 U11471 ( .B1(n9101), .B2(n11953), .A(n8995), .ZN(n8996) );
  AOI22_X1 U11472 ( .A1(n13630), .A2(n6619), .B1(n9097), .B2(n13367), .ZN(
        n9003) );
  NAND2_X1 U11473 ( .A1(n13630), .A2(n6618), .ZN(n8998) );
  NAND2_X1 U11474 ( .A1(n13367), .A2(n6619), .ZN(n8997) );
  NAND2_X1 U11475 ( .A1(n8998), .A2(n8997), .ZN(n9013) );
  AND2_X1 U11476 ( .A1(n13368), .A2(n9097), .ZN(n8999) );
  AOI21_X1 U11477 ( .B1(n14853), .B2(n6619), .A(n8999), .ZN(n9011) );
  NAND2_X1 U11478 ( .A1(n14853), .A2(n9097), .ZN(n9001) );
  NAND2_X1 U11479 ( .A1(n13368), .A2(n6619), .ZN(n9000) );
  NAND2_X1 U11480 ( .A1(n9001), .A2(n9000), .ZN(n9010) );
  AND2_X1 U11481 ( .A1(n9011), .A2(n9010), .ZN(n9002) );
  AND2_X1 U11482 ( .A1(n9097), .A2(n13369), .ZN(n9004) );
  AOI21_X1 U11483 ( .B1(n13642), .B2(n6619), .A(n9004), .ZN(n9009) );
  NAND2_X1 U11484 ( .A1(n13642), .A2(n6618), .ZN(n9006) );
  NAND2_X1 U11485 ( .A1(n13369), .A2(n6619), .ZN(n9005) );
  NAND2_X1 U11486 ( .A1(n9006), .A2(n9005), .ZN(n9008) );
  NAND2_X1 U11487 ( .A1(n9009), .A2(n9008), .ZN(n9007) );
  OAI22_X1 U11488 ( .A1(n9011), .A2(n9010), .B1(n9009), .B2(n9008), .ZN(n9015)
         );
  NOR2_X1 U11489 ( .A1(n13630), .A2(n13367), .ZN(n9012) );
  NOR2_X1 U11490 ( .A1(n9013), .A2(n9012), .ZN(n9014) );
  NAND2_X1 U11491 ( .A1(n9018), .A2(n9017), .ZN(n9023) );
  NAND2_X1 U11492 ( .A1(n13609), .A2(n6619), .ZN(n9020) );
  NAND2_X1 U11493 ( .A1(n13366), .A2(n9097), .ZN(n9019) );
  NAND2_X1 U11494 ( .A1(n13609), .A2(n6618), .ZN(n9021) );
  OAI21_X1 U11495 ( .B1(n9101), .B2(n13292), .A(n9021), .ZN(n9022) );
  NAND2_X1 U11496 ( .A1(n13731), .A2(n6618), .ZN(n9025) );
  NAND2_X1 U11497 ( .A1(n13365), .A2(n6619), .ZN(n9024) );
  NAND2_X1 U11498 ( .A1(n9025), .A2(n9024), .ZN(n9027) );
  AOI22_X1 U11499 ( .A1(n13731), .A2(n6619), .B1(n6618), .B2(n13365), .ZN(
        n9026) );
  NAND2_X1 U11500 ( .A1(n13726), .A2(n6619), .ZN(n9029) );
  NAND2_X1 U11501 ( .A1(n13364), .A2(n6618), .ZN(n9028) );
  NAND2_X1 U11502 ( .A1(n9029), .A2(n9028), .ZN(n9035) );
  NAND2_X1 U11503 ( .A1(n9034), .A2(n9035), .ZN(n9033) );
  NAND2_X1 U11504 ( .A1(n13726), .A2(n9097), .ZN(n9031) );
  NAND2_X1 U11505 ( .A1(n13364), .A2(n6619), .ZN(n9030) );
  NAND2_X1 U11506 ( .A1(n9031), .A2(n9030), .ZN(n9032) );
  NAND2_X1 U11507 ( .A1(n9033), .A2(n9032), .ZN(n9039) );
  INV_X1 U11508 ( .A(n9034), .ZN(n9037) );
  INV_X1 U11509 ( .A(n9035), .ZN(n9036) );
  NAND2_X1 U11510 ( .A1(n9037), .A2(n9036), .ZN(n9038) );
  NAND2_X1 U11511 ( .A1(n13557), .A2(n6618), .ZN(n9041) );
  NAND2_X1 U11512 ( .A1(n13363), .A2(n6619), .ZN(n9040) );
  AOI22_X1 U11513 ( .A1(n13557), .A2(n6619), .B1(n9097), .B2(n13363), .ZN(
        n9042) );
  NAND2_X1 U11514 ( .A1(n13716), .A2(n6619), .ZN(n9045) );
  NAND2_X1 U11515 ( .A1(n13362), .A2(n6618), .ZN(n9044) );
  NAND2_X1 U11516 ( .A1(n9045), .A2(n9044), .ZN(n9048) );
  NAND2_X1 U11517 ( .A1(n13716), .A2(n6618), .ZN(n9046) );
  OAI21_X1 U11518 ( .B1(n9101), .B2(n13271), .A(n9046), .ZN(n9047) );
  INV_X1 U11519 ( .A(n9048), .ZN(n9049) );
  NAND2_X1 U11520 ( .A1(n13524), .A2(n6618), .ZN(n9051) );
  NAND2_X1 U11521 ( .A1(n13361), .A2(n6619), .ZN(n9050) );
  NAND2_X1 U11522 ( .A1(n9051), .A2(n9050), .ZN(n9053) );
  AOI22_X1 U11523 ( .A1(n13524), .A2(n6619), .B1(n9097), .B2(n13361), .ZN(
        n9052) );
  AOI21_X1 U11524 ( .B1(n9054), .B2(n9053), .A(n9052), .ZN(n9056) );
  NOR2_X1 U11525 ( .A1(n9054), .A2(n9053), .ZN(n9055) );
  NAND2_X1 U11526 ( .A1(n13703), .A2(n6619), .ZN(n9058) );
  NAND2_X1 U11527 ( .A1(n9097), .A2(n13360), .ZN(n9057) );
  AOI22_X1 U11528 ( .A1(n13703), .A2(n6618), .B1(n6619), .B2(n13360), .ZN(
        n9059) );
  NAND2_X1 U11529 ( .A1(n13698), .A2(n6619), .ZN(n9061) );
  OAI21_X1 U11530 ( .B1(n13302), .B2(n9126), .A(n9061), .ZN(n9062) );
  OAI21_X1 U11531 ( .B1(n9065), .B2(n9064), .A(n9063), .ZN(n9070) );
  NAND2_X1 U11532 ( .A1(n13694), .A2(n6619), .ZN(n9067) );
  NAND2_X1 U11533 ( .A1(n9097), .A2(n13358), .ZN(n9066) );
  NAND2_X1 U11534 ( .A1(n9067), .A2(n9066), .ZN(n9069) );
  AOI22_X1 U11535 ( .A1(n13694), .A2(n9097), .B1(n6619), .B2(n13358), .ZN(
        n9068) );
  NAND2_X1 U11536 ( .A1(n13688), .A2(n9097), .ZN(n9073) );
  NAND2_X1 U11537 ( .A1(n6619), .A2(n13357), .ZN(n9072) );
  NAND2_X1 U11538 ( .A1(n9073), .A2(n9072), .ZN(n9100) );
  NAND2_X1 U11539 ( .A1(n13688), .A2(n6619), .ZN(n9075) );
  NAND2_X1 U11540 ( .A1(n9097), .A2(n13357), .ZN(n9074) );
  NAND2_X1 U11541 ( .A1(n9075), .A2(n9074), .ZN(n9095) );
  INV_X1 U11542 ( .A(SI_29_), .ZN(n13159) );
  NAND2_X1 U11543 ( .A1(n9078), .A2(n13159), .ZN(n9079) );
  MUX2_X1 U11544 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n7088), .Z(n9080) );
  NAND2_X1 U11545 ( .A1(n9080), .A2(SI_30_), .ZN(n9081) );
  OAI21_X1 U11546 ( .B1(n9080), .B2(SI_30_), .A(n9081), .ZN(n9104) );
  MUX2_X1 U11547 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n7088), .Z(n9082) );
  XNOR2_X1 U11548 ( .A(n9082), .B(SI_31_), .ZN(n9083) );
  NAND2_X1 U11549 ( .A1(n8730), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n9086) );
  INV_X1 U11550 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n9089) );
  NAND2_X1 U11551 ( .A1(n6627), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n9088) );
  NAND2_X1 U11552 ( .A1(n8389), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n9087) );
  OAI211_X1 U11553 ( .C1(n9090), .C2(n9089), .A(n9088), .B(n9087), .ZN(n13436)
         );
  AND2_X1 U11554 ( .A1(n6619), .A2(n13356), .ZN(n9091) );
  AOI21_X1 U11555 ( .B1(n13676), .B2(n9097), .A(n9091), .ZN(n9116) );
  NAND2_X1 U11556 ( .A1(n13676), .A2(n6619), .ZN(n9093) );
  NAND2_X1 U11557 ( .A1(n9097), .A2(n13356), .ZN(n9092) );
  NAND2_X1 U11558 ( .A1(n9093), .A2(n9092), .ZN(n9115) );
  NOR2_X1 U11559 ( .A1(n9126), .A2(n13254), .ZN(n9096) );
  AOI21_X1 U11560 ( .B1(n13455), .B2(n6619), .A(n9096), .ZN(n9120) );
  NAND2_X1 U11561 ( .A1(n13455), .A2(n9097), .ZN(n9099) );
  NAND2_X1 U11562 ( .A1(n6619), .A2(n11029), .ZN(n9098) );
  NAND2_X1 U11563 ( .A1(n9099), .A2(n9098), .ZN(n9119) );
  MUX2_X1 U11564 ( .A(n13436), .B(n9101), .S(n9128), .Z(n9103) );
  AND2_X1 U11565 ( .A1(n9101), .A2(n13436), .ZN(n9130) );
  INV_X1 U11566 ( .A(n9130), .ZN(n9102) );
  NAND2_X1 U11567 ( .A1(n9103), .A2(n9102), .ZN(n9118) );
  NAND2_X1 U11568 ( .A1(n8730), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n9108) );
  NAND2_X1 U11569 ( .A1(n6619), .A2(n13436), .ZN(n9127) );
  INV_X1 U11570 ( .A(n10916), .ZN(n9111) );
  OR2_X1 U11571 ( .A1(n9110), .A2(n9111), .ZN(n9133) );
  NAND4_X1 U11572 ( .A1(n9127), .A2(n9168), .A3(n9133), .A4(n9173), .ZN(n9112)
         );
  AOI22_X1 U11573 ( .A1(n13445), .A2(n6618), .B1(n13355), .B2(n9112), .ZN(
        n9125) );
  NAND2_X1 U11574 ( .A1(n13445), .A2(n6619), .ZN(n9114) );
  NAND2_X1 U11575 ( .A1(n6618), .A2(n13355), .ZN(n9113) );
  NAND2_X1 U11576 ( .A1(n9114), .A2(n9113), .ZN(n9124) );
  OAI22_X1 U11577 ( .A1(n9125), .A2(n9124), .B1(n9116), .B2(n9115), .ZN(n9117)
         );
  NAND2_X1 U11578 ( .A1(n9118), .A2(n9117), .ZN(n9122) );
  NAND4_X1 U11579 ( .A1(n9141), .A2(n9120), .A3(n9119), .A4(n6653), .ZN(n9121)
         );
  NAND2_X1 U11580 ( .A1(n9125), .A2(n9124), .ZN(n9132) );
  AND2_X1 U11581 ( .A1(n9127), .A2(n9126), .ZN(n9129) );
  MUX2_X1 U11582 ( .A(n9130), .B(n9129), .S(n9128), .Z(n9131) );
  OAI21_X1 U11583 ( .B1(n9134), .B2(n11531), .A(n9133), .ZN(n9135) );
  INV_X1 U11584 ( .A(n9135), .ZN(n9140) );
  INV_X1 U11585 ( .A(n9136), .ZN(n9137) );
  OAI211_X1 U11586 ( .C1(n13429), .C2(n11829), .A(n9137), .B(n9173), .ZN(n9138) );
  NAND2_X1 U11587 ( .A1(n9169), .A2(n9138), .ZN(n9139) );
  OAI21_X1 U11588 ( .B1(n9169), .B2(n9140), .A(n9139), .ZN(n9172) );
  XOR2_X1 U11589 ( .A(n13355), .B(n13445), .Z(n9164) );
  XNOR2_X1 U11590 ( .A(n13524), .B(n13304), .ZN(n13527) );
  XNOR2_X1 U11591 ( .A(n13731), .B(n13365), .ZN(n13581) );
  XNOR2_X1 U11592 ( .A(n14845), .B(n13370), .ZN(n12019) );
  AND2_X1 U11593 ( .A1(n10641), .A2(n9142), .ZN(n10924) );
  NAND4_X1 U11594 ( .A1(n10924), .A2(n9143), .A3(n13658), .A4(n9796), .ZN(
        n9144) );
  NOR2_X1 U11595 ( .A1(n9144), .A2(n10760), .ZN(n9146) );
  NAND4_X1 U11596 ( .A1(n9147), .A2(n9146), .A3(n9145), .A4(n10596), .ZN(n9148) );
  NOR2_X1 U11597 ( .A1(n11259), .A2(n9148), .ZN(n9150) );
  NAND4_X1 U11598 ( .A1(n11583), .A2(n9150), .A3(n9149), .A4(n11453), .ZN(
        n9151) );
  NOR2_X1 U11599 ( .A1(n11756), .A2(n9151), .ZN(n9153) );
  NAND4_X1 U11600 ( .A1(n12019), .A2(n9153), .A3(n11967), .A4(n9152), .ZN(
        n9154) );
  NOR2_X1 U11601 ( .A1(n12141), .A2(n9154), .ZN(n9155) );
  NAND4_X1 U11602 ( .A1(n13581), .A2(n9155), .A3(n13628), .A4(n12158), .ZN(
        n9156) );
  OR4_X1 U11603 ( .A1(n13548), .A2(n13573), .A3(n13595), .A4(n9156), .ZN(n9157) );
  OR4_X1 U11604 ( .A1(n9158), .A2(n13527), .A3(n13533), .A4(n9157), .ZN(n9159)
         );
  NOR2_X1 U11605 ( .A1(n13499), .A2(n9159), .ZN(n9160) );
  NAND4_X1 U11606 ( .A1(n9161), .A2(n9160), .A3(n13474), .A4(n13486), .ZN(
        n9162) );
  NOR4_X2 U11607 ( .A1(n9165), .A2(n9164), .A3(n9163), .A4(n9162), .ZN(n9166)
         );
  XNOR2_X1 U11608 ( .A(n9166), .B(n13429), .ZN(n9167) );
  OR2_X1 U11609 ( .A1(n10630), .A2(P2_U3088), .ZN(n12000) );
  INV_X1 U11610 ( .A(n12000), .ZN(n9170) );
  OAI21_X1 U11611 ( .B1(n9172), .B2(n9171), .A(n9170), .ZN(n9177) );
  INV_X1 U11612 ( .A(n15349), .ZN(n15346) );
  NOR4_X1 U11613 ( .A1(n15346), .A2(n13303), .A3(n8868), .A4(n9173), .ZN(n9175) );
  OAI21_X1 U11614 ( .B1(n12000), .B2(n8877), .A(P2_B_REG_SCAN_IN), .ZN(n9174)
         );
  OR2_X1 U11615 ( .A1(n9175), .A2(n9174), .ZN(n9176) );
  NAND2_X1 U11616 ( .A1(n9177), .A2(n9176), .ZN(P2_U3328) );
  NAND4_X1 U11617 ( .A1(n9184), .A2(n9183), .A3(n9182), .A4(n9417), .ZN(n9451)
         );
  INV_X1 U11618 ( .A(n9451), .ZN(n9186) );
  INV_X1 U11619 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n9185) );
  NAND2_X1 U11620 ( .A1(n9186), .A2(n9185), .ZN(n9187) );
  XNOR2_X2 U11621 ( .A(n9195), .B(n9194), .ZN(n9199) );
  NAND2_X1 U11622 ( .A1(n9196), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9197) );
  NAND2_X2 U11623 ( .A1(n9199), .A2(n9202), .ZN(n9270) );
  INV_X1 U11624 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n9198) );
  OR2_X1 U11625 ( .A1(n9270), .A2(n9198), .ZN(n9207) );
  NAND2_X1 U11626 ( .A1(n9298), .A2(n9297), .ZN(n9320) );
  OR2_X1 U11627 ( .A1(n9354), .A2(n9200), .ZN(n9201) );
  AND2_X1 U11628 ( .A1(n9366), .A2(n9201), .ZN(n11798) );
  OR2_X1 U11629 ( .A1(n9269), .A2(n11798), .ZN(n9206) );
  NAND2_X1 U11630 ( .A1(n11245), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n9205) );
  NAND2_X1 U11631 ( .A1(n9256), .A2(P3_REG0_REG_9__SCAN_IN), .ZN(n9204) );
  NAND4_X1 U11632 ( .A1(n9207), .A2(n9206), .A3(n9205), .A4(n9204), .ZN(n12734) );
  AND2_X2 U11633 ( .A1(n9250), .A2(n9213), .ZN(n9615) );
  INV_X1 U11634 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n9820) );
  NAND2_X1 U11635 ( .A1(n9820), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n9215) );
  NAND2_X1 U11636 ( .A1(n9216), .A2(n9215), .ZN(n9264) );
  XNOR2_X1 U11637 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .ZN(n9262) );
  NAND2_X1 U11638 ( .A1(n9264), .A2(n9262), .ZN(n9218) );
  NAND2_X1 U11639 ( .A1(n9818), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n9217) );
  XNOR2_X1 U11640 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .ZN(n9275) );
  NAND2_X1 U11641 ( .A1(n9277), .A2(n9275), .ZN(n9221) );
  INV_X1 U11642 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n9219) );
  NAND2_X1 U11643 ( .A1(n9219), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n9220) );
  NAND2_X1 U11644 ( .A1(n9822), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n9222) );
  NAND2_X1 U11645 ( .A1(n9821), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n9223) );
  NAND2_X1 U11646 ( .A1(n9833), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n9225) );
  NAND2_X1 U11647 ( .A1(n9893), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n9226) );
  NAND2_X1 U11648 ( .A1(n9896), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n9228) );
  XNOR2_X1 U11649 ( .A(n9373), .B(n9372), .ZN(n9835) );
  NAND2_X1 U11650 ( .A1(n9615), .A2(n9835), .ZN(n9232) );
  NAND2_X1 U11651 ( .A1(n9453), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9230) );
  XNOR2_X1 U11652 ( .A(n9230), .B(P3_IR_REG_9__SCAN_IN), .ZN(n11659) );
  OR2_X1 U11653 ( .A1(n10506), .A2(n11659), .ZN(n9231) );
  OAI211_X1 U11654 ( .C1(n9265), .C2(SI_9_), .A(n9232), .B(n9231), .ZN(n15485)
         );
  NAND2_X1 U11655 ( .A1(n9620), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n9237) );
  INV_X1 U11656 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n11027) );
  OR2_X1 U11657 ( .A1(n9269), .A2(n11027), .ZN(n9234) );
  NAND2_X1 U11658 ( .A1(n9257), .A2(P3_REG2_REG_1__SCAN_IN), .ZN(n9233) );
  NAND2_X1 U11659 ( .A1(n9256), .A2(P3_REG0_REG_1__SCAN_IN), .ZN(n9235) );
  INV_X1 U11660 ( .A(n9253), .ZN(n10719) );
  INV_X1 U11661 ( .A(SI_1_), .ZN(n9830) );
  XNOR2_X1 U11662 ( .A(n9238), .B(n9246), .ZN(n9829) );
  NAND2_X1 U11663 ( .A1(n9615), .A2(n9829), .ZN(n9241) );
  INV_X1 U11664 ( .A(P3_IR_REG_1__SCAN_IN), .ZN(n10528) );
  NAND2_X1 U11665 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), 
        .ZN(n9239) );
  XNOR2_X1 U11666 ( .A(n10528), .B(n9239), .ZN(n10511) );
  OR2_X1 U11667 ( .A1(n9250), .A2(n10511), .ZN(n9240) );
  INV_X1 U11668 ( .A(n11370), .ZN(n11023) );
  NAND2_X1 U11669 ( .A1(n9253), .A2(n11370), .ZN(n12530) );
  INV_X1 U11670 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n10513) );
  INV_X1 U11671 ( .A(P3_REG3_REG_0__SCAN_IN), .ZN(n11526) );
  OR2_X1 U11672 ( .A1(n9269), .A2(n11526), .ZN(n9244) );
  NAND2_X1 U11673 ( .A1(n9256), .A2(P3_REG0_REG_0__SCAN_IN), .ZN(n9243) );
  NAND2_X1 U11674 ( .A1(n9257), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n9242) );
  INV_X1 U11675 ( .A(n9246), .ZN(n9249) );
  NAND2_X1 U11676 ( .A1(n9247), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n9248) );
  NAND2_X1 U11677 ( .A1(n9249), .A2(n9248), .ZN(n9884) );
  NAND2_X1 U11678 ( .A1(n9615), .A2(n9884), .ZN(n9252) );
  INV_X1 U11679 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n10529) );
  OR2_X1 U11680 ( .A1(n9250), .A2(n10529), .ZN(n9251) );
  OAI211_X1 U11681 ( .C1(n9265), .C2(n9885), .A(n9252), .B(n9251), .ZN(n10913)
         );
  NAND2_X1 U11682 ( .A1(n10678), .A2(n11023), .ZN(n9254) );
  NAND2_X1 U11683 ( .A1(n9256), .A2(P3_REG0_REG_2__SCAN_IN), .ZN(n9261) );
  NAND2_X1 U11684 ( .A1(n9257), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n9260) );
  INV_X1 U11685 ( .A(P3_REG3_REG_2__SCAN_IN), .ZN(n10572) );
  OR2_X1 U11686 ( .A1(n9269), .A2(n10572), .ZN(n9259) );
  INV_X1 U11687 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n10516) );
  OR2_X1 U11688 ( .A1(n9270), .A2(n10516), .ZN(n9258) );
  INV_X1 U11689 ( .A(n9262), .ZN(n9263) );
  XNOR2_X1 U11690 ( .A(n9264), .B(n9263), .ZN(n9883) );
  OR2_X1 U11691 ( .A1(n9265), .A2(SI_2_), .ZN(n9268) );
  OR2_X1 U11692 ( .A1(n10506), .A2(n10533), .ZN(n9267) );
  NAND2_X1 U11693 ( .A1(n9256), .A2(P3_REG0_REG_3__SCAN_IN), .ZN(n9274) );
  NAND2_X1 U11694 ( .A1(n9257), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n9273) );
  OR2_X1 U11695 ( .A1(n9269), .A2(P3_REG3_REG_3__SCAN_IN), .ZN(n9272) );
  INV_X1 U11696 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n10797) );
  OR2_X1 U11697 ( .A1(n9270), .A2(n10797), .ZN(n9271) );
  INV_X1 U11698 ( .A(n9275), .ZN(n9276) );
  XNOR2_X1 U11699 ( .A(n9277), .B(n9276), .ZN(n9887) );
  NAND2_X1 U11700 ( .A1(n9615), .A2(n9887), .ZN(n9281) );
  OR2_X1 U11701 ( .A1(n9265), .A2(SI_3_), .ZN(n9280) );
  NAND2_X1 U11702 ( .A1(n9291), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9278) );
  XNOR2_X1 U11703 ( .A(n9278), .B(P3_IR_REG_3__SCAN_IN), .ZN(n10798) );
  OR2_X1 U11704 ( .A1(n10506), .A2(n10798), .ZN(n9279) );
  INV_X1 U11705 ( .A(n11479), .ZN(n10785) );
  NAND2_X1 U11706 ( .A1(n15451), .A2(n11479), .ZN(n12542) );
  NAND2_X1 U11707 ( .A1(n10780), .A2(n10779), .ZN(n10778) );
  NAND2_X1 U11708 ( .A1(n12739), .A2(n11479), .ZN(n9282) );
  NAND2_X1 U11709 ( .A1(n11245), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n9287) );
  NAND2_X1 U11710 ( .A1(n9256), .A2(P3_REG0_REG_4__SCAN_IN), .ZN(n9286) );
  INV_X1 U11711 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n10800) );
  OR2_X1 U11712 ( .A1(n9270), .A2(n10800), .ZN(n9285) );
  AND2_X1 U11713 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(P3_REG3_REG_3__SCAN_IN), 
        .ZN(n9283) );
  NOR2_X1 U11714 ( .A1(n9298), .A2(n9283), .ZN(n11009) );
  OR2_X1 U11715 ( .A1(n9269), .A2(n11009), .ZN(n9284) );
  INV_X1 U11716 ( .A(n9288), .ZN(n9289) );
  XNOR2_X1 U11717 ( .A(n9290), .B(n9289), .ZN(n9889) );
  NAND2_X1 U11718 ( .A1(n9615), .A2(n9889), .ZN(n9295) );
  OR2_X1 U11719 ( .A1(n9265), .A2(SI_4_), .ZN(n9294) );
  OR2_X1 U11720 ( .A1(n9291), .A2(P3_IR_REG_3__SCAN_IN), .ZN(n9307) );
  NAND2_X1 U11721 ( .A1(n9307), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9292) );
  XNOR2_X1 U11722 ( .A(n9292), .B(P3_IR_REG_4__SCAN_IN), .ZN(n15410) );
  OR2_X1 U11723 ( .A1(n10506), .A2(n15410), .ZN(n9293) );
  NAND2_X1 U11724 ( .A1(n11314), .A2(n15480), .ZN(n12546) );
  INV_X1 U11725 ( .A(n11314), .ZN(n12738) );
  INV_X1 U11726 ( .A(n15480), .ZN(n11010) );
  NAND2_X1 U11727 ( .A1(n12738), .A2(n11010), .ZN(n12545) );
  NAND2_X1 U11728 ( .A1(n12546), .A2(n12545), .ZN(n11388) );
  NAND2_X1 U11729 ( .A1(n11389), .A2(n11388), .ZN(n11387) );
  NAND2_X1 U11730 ( .A1(n12738), .A2(n15480), .ZN(n9296) );
  INV_X1 U11731 ( .A(n11312), .ZN(n9317) );
  NAND2_X1 U11732 ( .A1(n11245), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n9303) );
  NAND2_X1 U11733 ( .A1(n9256), .A2(P3_REG0_REG_5__SCAN_IN), .ZN(n9302) );
  INV_X1 U11734 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n10868) );
  OR2_X1 U11735 ( .A1(n9270), .A2(n10868), .ZN(n9301) );
  OR2_X1 U11736 ( .A1(n9298), .A2(n9297), .ZN(n9299) );
  AND2_X1 U11737 ( .A1(n9320), .A2(n9299), .ZN(n11534) );
  OR2_X1 U11738 ( .A1(n9269), .A2(n11534), .ZN(n9300) );
  INV_X1 U11739 ( .A(n9304), .ZN(n9305) );
  XNOR2_X1 U11740 ( .A(n9306), .B(n9305), .ZN(n9881) );
  NAND2_X1 U11741 ( .A1(n9615), .A2(n9881), .ZN(n9315) );
  OR2_X1 U11742 ( .A1(n9265), .A2(SI_5_), .ZN(n9314) );
  NOR2_X1 U11743 ( .A1(n9307), .A2(P3_IR_REG_4__SCAN_IN), .ZN(n9310) );
  NOR2_X1 U11744 ( .A1(n9310), .A2(n12321), .ZN(n9308) );
  MUX2_X1 U11745 ( .A(n12321), .B(n9308), .S(P3_IR_REG_5__SCAN_IN), .Z(n9312)
         );
  NAND2_X1 U11746 ( .A1(n9310), .A2(n9309), .ZN(n9328) );
  INV_X1 U11747 ( .A(n9328), .ZN(n9311) );
  INV_X1 U11748 ( .A(n10874), .ZN(n10808) );
  OR2_X1 U11749 ( .A1(n10506), .A2(n10808), .ZN(n9313) );
  NAND2_X1 U11750 ( .A1(n11437), .A2(n11155), .ZN(n12549) );
  INV_X1 U11751 ( .A(n11437), .ZN(n12737) );
  INV_X1 U11752 ( .A(n11155), .ZN(n11535) );
  NAND2_X1 U11753 ( .A1(n12737), .A2(n11535), .ZN(n12554) );
  NAND2_X1 U11754 ( .A1(n11437), .A2(n11535), .ZN(n9318) );
  NAND2_X1 U11755 ( .A1(n11245), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n9325) );
  NAND2_X1 U11756 ( .A1(n9256), .A2(P3_REG0_REG_6__SCAN_IN), .ZN(n9324) );
  INV_X1 U11757 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n9319) );
  OR2_X1 U11758 ( .A1(n9270), .A2(n9319), .ZN(n9323) );
  NAND2_X1 U11759 ( .A1(n9320), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n9321) );
  AND2_X1 U11760 ( .A1(n9333), .A2(n9321), .ZN(n15439) );
  OR2_X1 U11761 ( .A1(n9269), .A2(n15439), .ZN(n9322) );
  INV_X1 U11762 ( .A(SI_6_), .ZN(n9879) );
  XNOR2_X1 U11763 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .ZN(n9326) );
  XNOR2_X1 U11764 ( .A(n9327), .B(n9326), .ZN(n9878) );
  NAND2_X1 U11765 ( .A1(n9615), .A2(n9878), .ZN(n9331) );
  NAND2_X1 U11766 ( .A1(n9328), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9329) );
  XNOR2_X1 U11767 ( .A(n9329), .B(P3_IR_REG_6__SCAN_IN), .ZN(n10809) );
  INV_X1 U11768 ( .A(n10809), .ZN(n10849) );
  OR2_X1 U11769 ( .A1(n10506), .A2(n10849), .ZN(n9330) );
  OAI211_X1 U11770 ( .C1(n9265), .C2(n9879), .A(n9331), .B(n9330), .ZN(n11516)
         );
  NAND2_X1 U11771 ( .A1(n11444), .A2(n11516), .ZN(n12556) );
  INV_X1 U11772 ( .A(n11444), .ZN(n12736) );
  INV_X1 U11773 ( .A(n11516), .ZN(n15441) );
  NAND2_X1 U11774 ( .A1(n12736), .A2(n15441), .ZN(n12555) );
  NAND2_X1 U11775 ( .A1(n12556), .A2(n12555), .ZN(n12676) );
  NAND2_X1 U11776 ( .A1(n11245), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n9338) );
  NAND2_X1 U11777 ( .A1(n9256), .A2(P3_REG0_REG_7__SCAN_IN), .ZN(n9337) );
  INV_X1 U11778 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n9332) );
  OR2_X1 U11779 ( .A1(n9270), .A2(n9332), .ZN(n9336) );
  AND2_X1 U11780 ( .A1(n9333), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n9334) );
  NOR2_X1 U11781 ( .A1(n9352), .A2(n9334), .ZN(n11627) );
  OR2_X1 U11782 ( .A1(n9269), .A2(n11627), .ZN(n9335) );
  XNOR2_X1 U11783 ( .A(n9340), .B(n9339), .ZN(n9839) );
  NAND2_X1 U11784 ( .A1(n9615), .A2(n9839), .ZN(n9348) );
  OR2_X1 U11785 ( .A1(n9265), .A2(SI_7_), .ZN(n9347) );
  OR2_X1 U11786 ( .A1(n9342), .A2(n12321), .ZN(n9343) );
  MUX2_X1 U11787 ( .A(n9343), .B(P3_IR_REG_31__SCAN_IN), .S(n9344), .Z(n9345)
         );
  NAND2_X1 U11788 ( .A1(n9342), .A2(n9344), .ZN(n9362) );
  NAND2_X1 U11789 ( .A1(n9345), .A2(n9362), .ZN(n10900) );
  INV_X1 U11790 ( .A(n10900), .ZN(n10810) );
  OR2_X1 U11791 ( .A1(n10506), .A2(n10810), .ZN(n9346) );
  NAND2_X1 U11792 ( .A1(n11622), .A2(n11447), .ZN(n12561) );
  INV_X1 U11793 ( .A(n11622), .ZN(n12735) );
  NAND2_X1 U11794 ( .A1(n12735), .A2(n11628), .ZN(n12562) );
  NAND2_X1 U11795 ( .A1(n12561), .A2(n12562), .ZN(n11442) );
  NAND2_X1 U11796 ( .A1(n11405), .A2(n11442), .ZN(n11404) );
  NAND2_X1 U11797 ( .A1(n12735), .A2(n11447), .ZN(n9349) );
  NAND2_X1 U11798 ( .A1(n11245), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n9358) );
  NAND2_X1 U11799 ( .A1(n9256), .A2(P3_REG0_REG_8__SCAN_IN), .ZN(n9357) );
  INV_X1 U11800 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n9350) );
  OR2_X1 U11801 ( .A1(n9270), .A2(n9350), .ZN(n9356) );
  NOR2_X1 U11802 ( .A1(n9352), .A2(n9351), .ZN(n9353) );
  OR2_X1 U11803 ( .A1(n9269), .A2(n7578), .ZN(n9355) );
  INV_X1 U11804 ( .A(SI_8_), .ZN(n9842) );
  INV_X1 U11805 ( .A(n9359), .ZN(n9360) );
  XNOR2_X1 U11806 ( .A(n9361), .B(n9360), .ZN(n9841) );
  NAND2_X1 U11807 ( .A1(n9615), .A2(n9841), .ZN(n9365) );
  NAND2_X1 U11808 ( .A1(n9362), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9363) );
  XNOR2_X1 U11809 ( .A(n9363), .B(P3_IR_REG_8__SCAN_IN), .ZN(n11080) );
  INV_X1 U11810 ( .A(n11080), .ZN(n11076) );
  OR2_X1 U11811 ( .A1(n10506), .A2(n11076), .ZN(n9364) );
  OAI211_X1 U11812 ( .C1(n9265), .C2(n9842), .A(n9365), .B(n9364), .ZN(n11685)
         );
  NAND2_X1 U11813 ( .A1(n11794), .A2(n11685), .ZN(n12567) );
  INV_X1 U11814 ( .A(n11794), .ZN(n11788) );
  INV_X1 U11815 ( .A(n11685), .ZN(n11689) );
  NAND2_X1 U11816 ( .A1(n11788), .A2(n11689), .ZN(n12566) );
  XNOR2_X1 U11817 ( .A(n12734), .B(n15485), .ZN(n12565) );
  OAI21_X1 U11818 ( .B1(n11871), .B2(n15485), .A(n11732), .ZN(n11836) );
  NAND2_X1 U11819 ( .A1(n11245), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n9371) );
  NAND2_X1 U11820 ( .A1(n9256), .A2(P3_REG0_REG_10__SCAN_IN), .ZN(n9370) );
  INV_X1 U11821 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n11657) );
  OR2_X1 U11822 ( .A1(n9270), .A2(n11657), .ZN(n9369) );
  NAND2_X1 U11823 ( .A1(n9366), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n9367) );
  AND2_X1 U11824 ( .A1(n9398), .A2(n9367), .ZN(n11877) );
  OR2_X1 U11825 ( .A1(n9269), .A2(n11877), .ZN(n9368) );
  NAND2_X1 U11826 ( .A1(n9902), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n9374) );
  XNOR2_X1 U11827 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .ZN(n9385) );
  XNOR2_X1 U11828 ( .A(n9386), .B(n9385), .ZN(n9844) );
  NAND2_X1 U11829 ( .A1(n9615), .A2(n9844), .ZN(n9380) );
  OR2_X1 U11830 ( .A1(n9265), .A2(SI_10_), .ZN(n9379) );
  NAND2_X1 U11831 ( .A1(n9388), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9377) );
  INV_X1 U11832 ( .A(P3_IR_REG_10__SCAN_IN), .ZN(n9376) );
  XNOR2_X1 U11833 ( .A(n9377), .B(n9376), .ZN(n11661) );
  OR2_X1 U11834 ( .A1(n10506), .A2(n15416), .ZN(n9378) );
  NAND2_X1 U11835 ( .A1(n12006), .A2(n11874), .ZN(n12578) );
  NAND2_X1 U11836 ( .A1(n12733), .A2(n12574), .ZN(n9702) );
  NAND2_X1 U11837 ( .A1(n12578), .A2(n9702), .ZN(n11835) );
  NAND2_X1 U11838 ( .A1(n11836), .A2(n11835), .ZN(n11834) );
  NAND2_X1 U11839 ( .A1(n11245), .A2(P3_REG2_REG_11__SCAN_IN), .ZN(n9384) );
  NAND2_X1 U11840 ( .A1(n9256), .A2(P3_REG0_REG_11__SCAN_IN), .ZN(n9383) );
  INV_X1 U11841 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n11662) );
  OR2_X1 U11842 ( .A1(n9270), .A2(n11662), .ZN(n9382) );
  XNOR2_X1 U11843 ( .A(n9398), .B(n11708), .ZN(n12115) );
  OR2_X1 U11844 ( .A1(n9269), .A2(n12115), .ZN(n9381) );
  NAND2_X1 U11845 ( .A1(n10151), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n9387) );
  XNOR2_X1 U11846 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .ZN(n9405) );
  XNOR2_X1 U11847 ( .A(n9406), .B(n9405), .ZN(n9837) );
  NAND2_X1 U11848 ( .A1(n9615), .A2(n9837), .ZN(n9395) );
  NOR2_X1 U11849 ( .A1(n9388), .A2(P3_IR_REG_10__SCAN_IN), .ZN(n9391) );
  NOR2_X1 U11850 ( .A1(n9391), .A2(n12321), .ZN(n9389) );
  MUX2_X1 U11851 ( .A(n12321), .B(n9389), .S(P3_IR_REG_11__SCAN_IN), .Z(n9393)
         );
  INV_X1 U11852 ( .A(P3_IR_REG_11__SCAN_IN), .ZN(n9390) );
  NAND2_X1 U11853 ( .A1(n9391), .A2(n9390), .ZN(n9416) );
  INV_X1 U11854 ( .A(n9416), .ZN(n9392) );
  NOR2_X1 U11855 ( .A1(n9393), .A2(n9392), .ZN(n11675) );
  OR2_X1 U11856 ( .A1(n10506), .A2(n11675), .ZN(n9394) );
  OAI211_X1 U11857 ( .C1(n9265), .C2(SI_11_), .A(n9395), .B(n9394), .ZN(n12099) );
  NAND2_X1 U11858 ( .A1(n12113), .A2(n12099), .ZN(n9396) );
  INV_X1 U11859 ( .A(n12099), .ZN(n12117) );
  NAND2_X1 U11860 ( .A1(n11245), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n9403) );
  NAND2_X1 U11861 ( .A1(n9256), .A2(P3_REG0_REG_12__SCAN_IN), .ZN(n9402) );
  INV_X1 U11862 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n11663) );
  OR2_X1 U11863 ( .A1(n9270), .A2(n11663), .ZN(n9401) );
  NAND2_X1 U11864 ( .A1(n11656), .A2(n11708), .ZN(n9397) );
  OAI21_X1 U11865 ( .B1(n9398), .B2(P3_REG3_REG_11__SCAN_IN), .A(
        P3_REG3_REG_12__SCAN_IN), .ZN(n9399) );
  AND2_X1 U11866 ( .A1(n9423), .A2(n9399), .ZN(n12073) );
  OR2_X1 U11867 ( .A1(n9269), .A2(n12073), .ZN(n9400) );
  NAND2_X1 U11868 ( .A1(n9416), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9404) );
  XNOR2_X1 U11869 ( .A(n9404), .B(P3_IR_REG_12__SCAN_IN), .ZN(n11901) );
  NAND2_X1 U11870 ( .A1(n9407), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n9408) );
  NAND2_X1 U11871 ( .A1(n9409), .A2(n9408), .ZN(n9413) );
  XNOR2_X1 U11872 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .ZN(n9414) );
  INV_X1 U11873 ( .A(n9414), .ZN(n9410) );
  XNOR2_X1 U11874 ( .A(n9413), .B(n9410), .ZN(n9875) );
  NAND2_X1 U11875 ( .A1(n9615), .A2(n9875), .ZN(n9412) );
  OR2_X1 U11876 ( .A1(n9265), .A2(n9877), .ZN(n9411) );
  OAI211_X1 U11877 ( .C1(n10506), .C2(n11891), .A(n9412), .B(n9411), .ZN(
        n12417) );
  NAND2_X1 U11878 ( .A1(n12081), .A2(n12417), .ZN(n12587) );
  INV_X1 U11879 ( .A(n12417), .ZN(n14827) );
  NAND2_X1 U11880 ( .A1(n12732), .A2(n14827), .ZN(n12586) );
  NAND2_X1 U11881 ( .A1(n9414), .A2(n9413), .ZN(n9415) );
  XNOR2_X2 U11882 ( .A(n9430), .B(P2_DATAO_REG_13__SCAN_IN), .ZN(n9429) );
  XNOR2_X1 U11883 ( .A(n9429), .B(P1_DATAO_REG_13__SCAN_IN), .ZN(n9898) );
  NAND2_X1 U11884 ( .A1(n9898), .A2(n9615), .ZN(n9421) );
  OR2_X1 U11885 ( .A1(n9416), .A2(P3_IR_REG_12__SCAN_IN), .ZN(n9432) );
  NAND2_X1 U11886 ( .A1(n9432), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9418) );
  XNOR2_X1 U11887 ( .A(n9418), .B(n9417), .ZN(n11931) );
  INV_X1 U11888 ( .A(n11931), .ZN(n11899) );
  OAI22_X1 U11889 ( .A1(n9265), .A2(SI_13_), .B1(n11899), .B2(n10506), .ZN(
        n9419) );
  INV_X1 U11890 ( .A(n9419), .ZN(n9420) );
  NAND2_X1 U11891 ( .A1(n9421), .A2(n9420), .ZN(n14822) );
  INV_X1 U11892 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n9422) );
  OR2_X1 U11893 ( .A1(n9270), .A2(n9422), .ZN(n9428) );
  AND2_X1 U11894 ( .A1(n9423), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n9424) );
  NOR2_X1 U11895 ( .A1(n9438), .A2(n9424), .ZN(n12082) );
  OR2_X1 U11896 ( .A1(n9269), .A2(n12082), .ZN(n9427) );
  NAND2_X1 U11897 ( .A1(n11245), .A2(P3_REG2_REG_13__SCAN_IN), .ZN(n9426) );
  NAND2_X1 U11898 ( .A1(n9256), .A2(P3_REG0_REG_13__SCAN_IN), .ZN(n9425) );
  NAND4_X1 U11899 ( .A1(n9428), .A2(n9427), .A3(n9426), .A4(n9425), .ZN(n12419) );
  OR2_X1 U11900 ( .A1(n14822), .A2(n12419), .ZN(n12592) );
  NAND2_X1 U11901 ( .A1(n14822), .A2(n12419), .ZN(n12591) );
  NAND2_X1 U11902 ( .A1(n12592), .A2(n12591), .ZN(n12685) );
  INV_X1 U11903 ( .A(n12419), .ZN(n12070) );
  NAND2_X1 U11904 ( .A1(n10553), .A2(n9430), .ZN(n9431) );
  XNOR2_X1 U11905 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .ZN(n9446) );
  XNOR2_X1 U11906 ( .A(n9447), .B(n9446), .ZN(n9903) );
  NAND2_X1 U11907 ( .A1(n9903), .A2(n9615), .ZN(n9436) );
  OAI21_X1 U11908 ( .B1(n9432), .B2(P3_IR_REG_13__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n9433) );
  XNOR2_X1 U11909 ( .A(n9433), .B(P3_IR_REG_14__SCAN_IN), .ZN(n12746) );
  OAI22_X1 U11910 ( .A1(n9265), .A2(SI_14_), .B1(n12746), .B2(n10506), .ZN(
        n9434) );
  INV_X1 U11911 ( .A(n9434), .ZN(n9435) );
  NAND2_X1 U11912 ( .A1(n9436), .A2(n9435), .ZN(n12130) );
  INV_X1 U11913 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n11914) );
  OR2_X1 U11914 ( .A1(n9270), .A2(n11914), .ZN(n9443) );
  OR2_X1 U11915 ( .A1(n9438), .A2(n9437), .ZN(n9439) );
  NAND2_X1 U11916 ( .A1(n9438), .A2(n9437), .ZN(n9458) );
  AND2_X1 U11917 ( .A1(n9439), .A2(n9458), .ZN(n12106) );
  OR2_X1 U11918 ( .A1(n9269), .A2(n12106), .ZN(n9442) );
  NAND2_X1 U11919 ( .A1(n11245), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n9441) );
  NAND2_X1 U11920 ( .A1(n9256), .A2(P3_REG0_REG_14__SCAN_IN), .ZN(n9440) );
  NAND4_X1 U11921 ( .A1(n9443), .A2(n9442), .A3(n9441), .A4(n9440), .ZN(n12731) );
  OR2_X1 U11922 ( .A1(n12130), .A2(n12731), .ZN(n12596) );
  NAND2_X1 U11923 ( .A1(n12130), .A2(n12731), .ZN(n12595) );
  NAND2_X1 U11924 ( .A1(n12596), .A2(n12595), .ZN(n12126) );
  NAND2_X1 U11925 ( .A1(n12124), .A2(n12126), .ZN(n9445) );
  INV_X1 U11926 ( .A(n12130), .ZN(n13101) );
  NAND2_X1 U11927 ( .A1(n13101), .A2(n12731), .ZN(n9444) );
  INV_X1 U11928 ( .A(n12150), .ZN(n9464) );
  NAND2_X1 U11929 ( .A1(n9448), .A2(P1_DATAO_REG_14__SCAN_IN), .ZN(n9449) );
  XNOR2_X1 U11930 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .ZN(n9467) );
  INV_X1 U11931 ( .A(n9467), .ZN(n9450) );
  XNOR2_X1 U11932 ( .A(n9468), .B(n9450), .ZN(n10369) );
  INV_X1 U11933 ( .A(SI_15_), .ZN(n10371) );
  OR2_X1 U11934 ( .A1(n9749), .A2(n12321), .ZN(n9454) );
  MUX2_X1 U11935 ( .A(n9454), .B(P3_IR_REG_31__SCAN_IN), .S(n9455), .Z(n9456)
         );
  NAND2_X1 U11936 ( .A1(n9456), .A2(n9494), .ZN(n12784) );
  OAI22_X1 U11937 ( .A1(n9265), .A2(n10371), .B1(n10506), .B2(n12784), .ZN(
        n9457) );
  NAND2_X1 U11938 ( .A1(n9256), .A2(P3_REG0_REG_15__SCAN_IN), .ZN(n9463) );
  NAND2_X1 U11939 ( .A1(n11245), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n9462) );
  INV_X1 U11940 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n12757) );
  OR2_X1 U11941 ( .A1(n9270), .A2(n12757), .ZN(n9461) );
  NAND2_X1 U11942 ( .A1(n9458), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n9459) );
  AND2_X1 U11943 ( .A1(n9475), .A2(n9459), .ZN(n12502) );
  OR2_X1 U11944 ( .A1(n9269), .A2(n12502), .ZN(n9460) );
  NAND2_X1 U11945 ( .A1(n9464), .A2(n7580), .ZN(n9466) );
  NAND2_X1 U11946 ( .A1(n12510), .A2(n12599), .ZN(n9465) );
  OAI21_X2 U11947 ( .B1(P2_DATAO_REG_15__SCAN_IN), .B2(n11168), .A(n9469), 
        .ZN(n9490) );
  AOI22_X1 U11948 ( .A1(P2_DATAO_REG_16__SCAN_IN), .A2(n11269), .B1(
        P1_DATAO_REG_16__SCAN_IN), .B2(n11238), .ZN(n9489) );
  INV_X1 U11949 ( .A(n9489), .ZN(n9470) );
  XNOR2_X1 U11950 ( .A(n9490), .B(n9470), .ZN(n10423) );
  NAND2_X1 U11951 ( .A1(n10423), .A2(n9615), .ZN(n9474) );
  NAND2_X1 U11952 ( .A1(n9494), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9471) );
  XNOR2_X1 U11953 ( .A(n9471), .B(P3_IR_REG_16__SCAN_IN), .ZN(n12794) );
  INV_X1 U11954 ( .A(n12794), .ZN(n12802) );
  OAI22_X1 U11955 ( .A1(n9265), .A2(n10425), .B1(n10506), .B2(n12802), .ZN(
        n9472) );
  INV_X1 U11956 ( .A(n9472), .ZN(n9473) );
  INV_X1 U11957 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n12793) );
  OR2_X1 U11958 ( .A1(n9270), .A2(n12793), .ZN(n9480) );
  AND2_X1 U11959 ( .A1(n9475), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n9476) );
  NOR2_X1 U11960 ( .A1(n9483), .A2(n9476), .ZN(n13036) );
  OR2_X1 U11961 ( .A1(n9269), .A2(n13036), .ZN(n9479) );
  NAND2_X1 U11962 ( .A1(n11245), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n9478) );
  NAND2_X1 U11963 ( .A1(n9256), .A2(P3_REG0_REG_16__SCAN_IN), .ZN(n9477) );
  NAND4_X1 U11964 ( .A1(n9480), .A2(n9479), .A3(n9478), .A4(n9477), .ZN(n12730) );
  NOR2_X1 U11965 ( .A1(n13093), .A2(n12730), .ZN(n9481) );
  INV_X1 U11966 ( .A(n12730), .ZN(n13016) );
  INV_X1 U11967 ( .A(n13093), .ZN(n13035) );
  NAND2_X1 U11968 ( .A1(n11245), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n9488) );
  NAND2_X1 U11969 ( .A1(n9256), .A2(P3_REG0_REG_17__SCAN_IN), .ZN(n9487) );
  INV_X1 U11970 ( .A(P3_REG1_REG_17__SCAN_IN), .ZN(n13090) );
  OR2_X1 U11971 ( .A1(n9270), .A2(n13090), .ZN(n9486) );
  INV_X1 U11972 ( .A(P3_REG3_REG_17__SCAN_IN), .ZN(n9482) );
  NOR2_X1 U11973 ( .A1(n9483), .A2(n9482), .ZN(n9484) );
  NOR2_X1 U11974 ( .A1(n9511), .A2(n9484), .ZN(n13018) );
  OR2_X1 U11975 ( .A1(n9269), .A2(n13018), .ZN(n9485) );
  XNOR2_X1 U11976 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(P2_DATAO_REG_17__SCAN_IN), 
        .ZN(n9501) );
  INV_X1 U11977 ( .A(n9501), .ZN(n9493) );
  NAND2_X1 U11978 ( .A1(n11238), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n9491) );
  XNOR2_X1 U11979 ( .A(n9493), .B(n9500), .ZN(n10490) );
  NAND2_X1 U11980 ( .A1(n9615), .A2(n10490), .ZN(n9498) );
  NAND2_X1 U11981 ( .A1(n9523), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9496) );
  INV_X1 U11982 ( .A(P3_IR_REG_17__SCAN_IN), .ZN(n9495) );
  XNOR2_X1 U11983 ( .A(n9496), .B(n9495), .ZN(n12817) );
  OR2_X1 U11984 ( .A1(n10506), .A2(n12817), .ZN(n9497) );
  OAI211_X1 U11985 ( .C1(n9265), .C2(n9499), .A(n9498), .B(n9497), .ZN(n12445)
         );
  NAND2_X1 U11986 ( .A1(n12478), .A2(n12445), .ZN(n12608) );
  INV_X1 U11987 ( .A(n12445), .ZN(n13145) );
  NAND2_X1 U11988 ( .A1(n13030), .A2(n13145), .ZN(n12609) );
  NAND2_X1 U11989 ( .A1(n12608), .A2(n12609), .ZN(n13013) );
  AOI22_X1 U11990 ( .A1(P2_DATAO_REG_18__SCAN_IN), .A2(n11433), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(n11431), .ZN(n9519) );
  INV_X1 U11991 ( .A(n9519), .ZN(n9503) );
  XNOR2_X1 U11992 ( .A(n9520), .B(n9503), .ZN(n14797) );
  NAND2_X1 U11993 ( .A1(n14797), .A2(n9615), .ZN(n9509) );
  OAI21_X1 U11994 ( .B1(n9523), .B2(P3_IR_REG_17__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n9505) );
  INV_X1 U11995 ( .A(P3_IR_REG_18__SCAN_IN), .ZN(n9504) );
  XNOR2_X1 U11996 ( .A(n9505), .B(n9504), .ZN(n14799) );
  OAI22_X1 U11997 ( .A1(n9265), .A2(n9506), .B1(n10506), .B2(n14799), .ZN(
        n9507) );
  INV_X1 U11998 ( .A(n9507), .ZN(n9508) );
  NAND2_X1 U11999 ( .A1(n9509), .A2(n9508), .ZN(n13009) );
  NAND2_X1 U12000 ( .A1(n11245), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n9516) );
  NAND2_X1 U12001 ( .A1(n9256), .A2(P3_REG0_REG_18__SCAN_IN), .ZN(n9515) );
  INV_X1 U12002 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n12820) );
  OR2_X1 U12003 ( .A1(n9270), .A2(n12820), .ZN(n9514) );
  OR2_X1 U12004 ( .A1(n9511), .A2(n9510), .ZN(n9512) );
  AND2_X1 U12005 ( .A1(n9533), .A2(n9512), .ZN(n13005) );
  OR2_X1 U12006 ( .A1(n9269), .A2(n13005), .ZN(n9513) );
  OR2_X1 U12007 ( .A1(n13009), .A2(n13017), .ZN(n12993) );
  NAND2_X1 U12008 ( .A1(n13009), .A2(n13017), .ZN(n12615) );
  NAND2_X2 U12009 ( .A1(n6651), .A2(n9517), .ZN(n13002) );
  INV_X1 U12010 ( .A(n13009), .ZN(n13087) );
  NAND2_X1 U12011 ( .A1(n13087), .A2(n13017), .ZN(n9518) );
  AOI22_X1 U12012 ( .A1(P2_DATAO_REG_19__SCAN_IN), .A2(n11532), .B1(
        P1_DATAO_REG_19__SCAN_IN), .B2(n7176), .ZN(n9542) );
  XNOR2_X1 U12013 ( .A(n9541), .B(n9542), .ZN(n10726) );
  NAND2_X1 U12014 ( .A1(n10726), .A2(n9615), .ZN(n9532) );
  INV_X1 U12015 ( .A(n9528), .ZN(n9525) );
  NAND2_X1 U12016 ( .A1(n9525), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9526) );
  MUX2_X1 U12017 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9526), .S(
        P3_IR_REG_19__SCAN_IN), .Z(n9529) );
  INV_X2 U12018 ( .A(n12832), .ZN(n12847) );
  OAI22_X1 U12019 ( .A1(n9265), .A2(SI_19_), .B1(n12847), .B2(n10506), .ZN(
        n9530) );
  INV_X1 U12020 ( .A(n9530), .ZN(n9531) );
  INV_X1 U12021 ( .A(P3_REG1_REG_19__SCAN_IN), .ZN(n13081) );
  OR2_X1 U12022 ( .A1(n9270), .A2(n13081), .ZN(n9538) );
  NAND2_X1 U12023 ( .A1(n9533), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n9534) );
  AND2_X1 U12024 ( .A1(n9546), .A2(n9534), .ZN(n12996) );
  OR2_X1 U12025 ( .A1(n9269), .A2(n12996), .ZN(n9537) );
  NAND2_X1 U12026 ( .A1(n11245), .A2(P3_REG2_REG_19__SCAN_IN), .ZN(n9536) );
  NAND2_X1 U12027 ( .A1(n9256), .A2(P3_REG0_REG_19__SCAN_IN), .ZN(n9535) );
  NAND4_X1 U12028 ( .A1(n9538), .A2(n9537), .A3(n9536), .A4(n9535), .ZN(n13003) );
  NAND2_X1 U12029 ( .A1(n13139), .A2(n13003), .ZN(n12620) );
  INV_X1 U12030 ( .A(n13139), .ZN(n9539) );
  NAND2_X1 U12031 ( .A1(n9539), .A2(n13003), .ZN(n9540) );
  XNOR2_X1 U12032 ( .A(n9555), .B(P2_DATAO_REG_20__SCAN_IN), .ZN(n11239) );
  NAND2_X1 U12033 ( .A1(n11239), .A2(n9615), .ZN(n9544) );
  OR2_X1 U12034 ( .A1(n9265), .A2(n11240), .ZN(n9543) );
  NAND2_X1 U12035 ( .A1(n11245), .A2(P3_REG2_REG_20__SCAN_IN), .ZN(n9551) );
  NAND2_X1 U12036 ( .A1(n9256), .A2(P3_REG0_REG_20__SCAN_IN), .ZN(n9550) );
  INV_X1 U12037 ( .A(P3_REG1_REG_20__SCAN_IN), .ZN(n9545) );
  OR2_X1 U12038 ( .A1(n9270), .A2(n9545), .ZN(n9549) );
  AND2_X1 U12039 ( .A1(n9546), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n9547) );
  NOR2_X1 U12040 ( .A1(n9562), .A2(n9547), .ZN(n12979) );
  OR2_X1 U12041 ( .A1(n9269), .A2(n12979), .ZN(n9548) );
  XNOR2_X1 U12042 ( .A(n12982), .B(n12966), .ZN(n12983) );
  NAND2_X1 U12043 ( .A1(n12982), .A2(n12989), .ZN(n9552) );
  NAND2_X1 U12044 ( .A1(n9553), .A2(n9552), .ZN(n12964) );
  INV_X1 U12045 ( .A(n12964), .ZN(n9568) );
  NAND2_X1 U12046 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n9554), .ZN(n9557) );
  NAND2_X1 U12047 ( .A1(n9555), .A2(n12313), .ZN(n9556) );
  AOI22_X1 U12048 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(n11832), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(n11830), .ZN(n9571) );
  INV_X1 U12049 ( .A(n9571), .ZN(n9558) );
  XNOR2_X1 U12050 ( .A(n9570), .B(n9558), .ZN(n11321) );
  NAND2_X1 U12051 ( .A1(n11321), .A2(n9615), .ZN(n9560) );
  INV_X1 U12052 ( .A(SI_21_), .ZN(n11323) );
  OR2_X1 U12053 ( .A1(n9265), .A2(n11323), .ZN(n9559) );
  INV_X1 U12054 ( .A(P3_REG3_REG_21__SCAN_IN), .ZN(n9561) );
  NOR2_X1 U12055 ( .A1(n9562), .A2(n9561), .ZN(n9563) );
  OR2_X1 U12056 ( .A1(n9577), .A2(n9563), .ZN(n12970) );
  NAND2_X1 U12057 ( .A1(n9665), .A2(n12970), .ZN(n9567) );
  NAND2_X1 U12058 ( .A1(n11245), .A2(P3_REG2_REG_21__SCAN_IN), .ZN(n9566) );
  INV_X1 U12059 ( .A(P3_REG1_REG_21__SCAN_IN), .ZN(n13072) );
  OR2_X1 U12060 ( .A1(n9270), .A2(n13072), .ZN(n9565) );
  NAND2_X1 U12061 ( .A1(n9256), .A2(P3_REG0_REG_21__SCAN_IN), .ZN(n9564) );
  NAND2_X1 U12062 ( .A1(n13134), .A2(n12954), .ZN(n9569) );
  INV_X1 U12063 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n9572) );
  AOI22_X1 U12064 ( .A1(P2_DATAO_REG_22__SCAN_IN), .A2(
        P1_DATAO_REG_22__SCAN_IN), .B1(n12171), .B2(n9572), .ZN(n9583) );
  XNOR2_X1 U12065 ( .A(n9584), .B(n9583), .ZN(n11472) );
  NAND2_X1 U12066 ( .A1(n11472), .A2(n9615), .ZN(n9575) );
  INV_X1 U12067 ( .A(SI_22_), .ZN(n9573) );
  OR2_X1 U12068 ( .A1(n9265), .A2(n9573), .ZN(n9574) );
  INV_X1 U12069 ( .A(P3_REG1_REG_22__SCAN_IN), .ZN(n13068) );
  OR2_X1 U12070 ( .A1(n9270), .A2(n13068), .ZN(n9582) );
  INV_X1 U12071 ( .A(P3_REG3_REG_22__SCAN_IN), .ZN(n9576) );
  OR2_X1 U12072 ( .A1(n9577), .A2(n9576), .ZN(n9578) );
  NAND2_X1 U12073 ( .A1(n9587), .A2(n9578), .ZN(n12959) );
  NAND2_X1 U12074 ( .A1(n9665), .A2(n12959), .ZN(n9581) );
  NAND2_X1 U12075 ( .A1(n11245), .A2(P3_REG2_REG_22__SCAN_IN), .ZN(n9580) );
  NAND2_X1 U12076 ( .A1(n9256), .A2(P3_REG0_REG_22__SCAN_IN), .ZN(n9579) );
  NAND4_X1 U12077 ( .A1(n9582), .A2(n9581), .A3(n9580), .A4(n9579), .ZN(n12940) );
  NOR2_X1 U12078 ( .A1(n12958), .A2(n12940), .ZN(n12934) );
  INV_X1 U12079 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n12002) );
  AOI22_X1 U12080 ( .A1(P1_DATAO_REG_23__SCAN_IN), .A2(
        P2_DATAO_REG_23__SCAN_IN), .B1(n11998), .B2(n12002), .ZN(n9600) );
  XNOR2_X1 U12081 ( .A(n9601), .B(n9600), .ZN(n11645) );
  NAND2_X1 U12082 ( .A1(n11645), .A2(n9615), .ZN(n9586) );
  INV_X1 U12083 ( .A(SI_23_), .ZN(n11647) );
  OR2_X1 U12084 ( .A1(n9265), .A2(n11647), .ZN(n9585) );
  NAND2_X1 U12085 ( .A1(n9587), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n9588) );
  NAND2_X1 U12086 ( .A1(n9603), .A2(n9588), .ZN(n12945) );
  NAND2_X1 U12087 ( .A1(n12945), .A2(n9665), .ZN(n9592) );
  INV_X1 U12088 ( .A(P3_REG1_REG_23__SCAN_IN), .ZN(n13064) );
  OR2_X1 U12089 ( .A1(n9270), .A2(n13064), .ZN(n9591) );
  NAND2_X1 U12090 ( .A1(n9256), .A2(P3_REG0_REG_23__SCAN_IN), .ZN(n9590) );
  NAND2_X1 U12091 ( .A1(n11245), .A2(P3_REG2_REG_23__SCAN_IN), .ZN(n9589) );
  NAND4_X1 U12092 ( .A1(n9592), .A2(n9591), .A3(n9590), .A4(n9589), .ZN(n12729) );
  NAND2_X1 U12093 ( .A1(n12949), .A2(n12729), .ZN(n9595) );
  INV_X1 U12094 ( .A(n9595), .ZN(n9594) );
  NAND2_X1 U12095 ( .A1(n13126), .A2(n12729), .ZN(n12513) );
  NAND2_X1 U12096 ( .A1(n12949), .A2(n12955), .ZN(n9593) );
  NAND2_X1 U12097 ( .A1(n12513), .A2(n9593), .ZN(n9709) );
  NOR2_X1 U12098 ( .A1(n9594), .A2(n9709), .ZN(n9597) );
  NAND2_X1 U12099 ( .A1(n12958), .A2(n12940), .ZN(n12935) );
  AND2_X1 U12100 ( .A1(n12935), .A2(n9595), .ZN(n9596) );
  OR2_X1 U12101 ( .A1(n9597), .A2(n9596), .ZN(n9598) );
  INV_X1 U12102 ( .A(SI_24_), .ZN(n12050) );
  OR2_X1 U12103 ( .A1(n9265), .A2(n12050), .ZN(n9602) );
  INV_X1 U12104 ( .A(n9256), .ZN(n9607) );
  INV_X1 U12105 ( .A(P3_REG0_REG_24__SCAN_IN), .ZN(n13120) );
  NAND2_X1 U12106 ( .A1(n9603), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n9604) );
  NAND2_X1 U12107 ( .A1(n9618), .A2(n9604), .ZN(n12924) );
  NAND2_X1 U12108 ( .A1(n12924), .A2(n9665), .ZN(n9606) );
  AOI22_X1 U12109 ( .A1(n9620), .A2(P3_REG1_REG_24__SCAN_IN), .B1(n11245), 
        .B2(P3_REG2_REG_24__SCAN_IN), .ZN(n9605) );
  NOR2_X1 U12110 ( .A1(n13122), .A2(n12451), .ZN(n9608) );
  NAND2_X1 U12111 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n9609), .ZN(n9612) );
  NAND2_X1 U12112 ( .A1(n9610), .A2(n12135), .ZN(n9611) );
  AOI22_X1 U12113 ( .A1(P2_DATAO_REG_25__SCAN_IN), .A2(n13805), .B1(
        P1_DATAO_REG_25__SCAN_IN), .B2(n14773), .ZN(n9613) );
  INV_X1 U12114 ( .A(n9613), .ZN(n9614) );
  XNOR2_X1 U12115 ( .A(n9626), .B(n9614), .ZN(n12089) );
  NAND2_X1 U12116 ( .A1(n12089), .A2(n9615), .ZN(n9617) );
  OR2_X1 U12117 ( .A1(n9265), .A2(n12091), .ZN(n9616) );
  AND2_X1 U12118 ( .A1(n9618), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n9619) );
  OR2_X1 U12119 ( .A1(n9619), .A2(n9631), .ZN(n12909) );
  NAND2_X1 U12120 ( .A1(n12909), .A2(n9665), .ZN(n9623) );
  AOI22_X1 U12121 ( .A1(n9620), .A2(P3_REG1_REG_25__SCAN_IN), .B1(n11245), 
        .B2(P3_REG2_REG_25__SCAN_IN), .ZN(n9622) );
  NAND2_X1 U12122 ( .A1(n9256), .A2(P3_REG0_REG_25__SCAN_IN), .ZN(n9621) );
  OR2_X1 U12123 ( .A1(n12908), .A2(n12920), .ZN(n12512) );
  NAND2_X1 U12124 ( .A1(n12908), .A2(n12920), .ZN(n12511) );
  NAND2_X1 U12125 ( .A1(n12908), .A2(n12728), .ZN(n9624) );
  NAND2_X1 U12126 ( .A1(P2_DATAO_REG_25__SCAN_IN), .A2(n13805), .ZN(n9625) );
  AOI22_X1 U12127 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(n14768), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n13800), .ZN(n9627) );
  XNOR2_X1 U12128 ( .A(n9642), .B(n9627), .ZN(n13169) );
  NAND2_X1 U12129 ( .A1(n13169), .A2(n9615), .ZN(n9629) );
  INV_X1 U12130 ( .A(SI_26_), .ZN(n13170) );
  OR2_X1 U12131 ( .A1(n9265), .A2(n13170), .ZN(n9628) );
  INV_X1 U12132 ( .A(P3_REG3_REG_26__SCAN_IN), .ZN(n9630) );
  NOR2_X1 U12133 ( .A1(n9631), .A2(n9630), .ZN(n9632) );
  OR2_X1 U12134 ( .A1(n9647), .A2(n9632), .ZN(n12895) );
  NAND2_X1 U12135 ( .A1(n12895), .A2(n9665), .ZN(n9637) );
  INV_X1 U12136 ( .A(P3_REG1_REG_26__SCAN_IN), .ZN(n13051) );
  NAND2_X1 U12137 ( .A1(n11245), .A2(P3_REG2_REG_26__SCAN_IN), .ZN(n9634) );
  NAND2_X1 U12138 ( .A1(n9256), .A2(P3_REG0_REG_26__SCAN_IN), .ZN(n9633) );
  OAI211_X1 U12139 ( .C1(n9270), .C2(n13051), .A(n9634), .B(n9633), .ZN(n9635)
         );
  INV_X1 U12140 ( .A(n9635), .ZN(n9636) );
  NAND2_X1 U12141 ( .A1(n12492), .A2(n12904), .ZN(n9640) );
  NOR2_X1 U12142 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(n14768), .ZN(n9641) );
  AOI22_X1 U12143 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(n13797), .B1(
        P1_DATAO_REG_27__SCAN_IN), .B2(n14767), .ZN(n9643) );
  INV_X1 U12144 ( .A(n9643), .ZN(n9644) );
  XNOR2_X1 U12145 ( .A(n9653), .B(n9644), .ZN(n13164) );
  NAND2_X1 U12146 ( .A1(n13164), .A2(n9615), .ZN(n9646) );
  OR2_X1 U12147 ( .A1(n9265), .A2(n13166), .ZN(n9645) );
  INV_X1 U12148 ( .A(P3_REG3_REG_27__SCAN_IN), .ZN(n12369) );
  NOR2_X1 U12149 ( .A1(n9647), .A2(n12369), .ZN(n9648) );
  INV_X1 U12150 ( .A(P3_REG1_REG_27__SCAN_IN), .ZN(n13047) );
  NAND2_X1 U12151 ( .A1(n9256), .A2(P3_REG0_REG_27__SCAN_IN), .ZN(n9650) );
  NAND2_X1 U12152 ( .A1(n11245), .A2(P3_REG2_REG_27__SCAN_IN), .ZN(n9649) );
  OAI211_X1 U12153 ( .C1(n9270), .C2(n13047), .A(n9650), .B(n9649), .ZN(n9651)
         );
  OR2_X1 U12154 ( .A1(n12372), .A2(n12891), .ZN(n12652) );
  NAND2_X1 U12155 ( .A1(n12372), .A2(n12891), .ZN(n12646) );
  NAND2_X1 U12156 ( .A1(n13111), .A2(n12891), .ZN(n9652) );
  NAND2_X1 U12157 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(n13797), .ZN(n9654) );
  AOI22_X1 U12158 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(
        P2_DATAO_REG_28__SCAN_IN), .B1(n9669), .B2(n8218), .ZN(n9655) );
  INV_X1 U12159 ( .A(n9655), .ZN(n9656) );
  NAND2_X1 U12160 ( .A1(n13160), .A2(n9615), .ZN(n9658) );
  OR2_X1 U12161 ( .A1(n9265), .A2(n13163), .ZN(n9657) );
  INV_X1 U12162 ( .A(P3_REG3_REG_28__SCAN_IN), .ZN(n12395) );
  NAND2_X1 U12163 ( .A1(n9659), .A2(n12395), .ZN(n12329) );
  OR2_X1 U12164 ( .A1(n9659), .A2(n12395), .ZN(n9660) );
  NAND2_X1 U12165 ( .A1(n12329), .A2(n9660), .ZN(n12864) );
  INV_X1 U12166 ( .A(P3_REG1_REG_28__SCAN_IN), .ZN(n9663) );
  NAND2_X1 U12167 ( .A1(n11245), .A2(P3_REG2_REG_28__SCAN_IN), .ZN(n9662) );
  NAND2_X1 U12168 ( .A1(n9256), .A2(P3_REG0_REG_28__SCAN_IN), .ZN(n9661) );
  OAI211_X1 U12169 ( .C1(n9270), .C2(n9663), .A(n9662), .B(n9661), .ZN(n9664)
         );
  INV_X1 U12170 ( .A(n12863), .ZN(n9666) );
  NOR2_X1 U12171 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(n9669), .ZN(n9671) );
  NAND2_X1 U12172 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(n9669), .ZN(n9670) );
  OAI22_X1 U12173 ( .A1(n14764), .A2(n13790), .B1(P1_DATAO_REG_29__SCAN_IN), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n12315) );
  INV_X1 U12174 ( .A(n12315), .ZN(n9673) );
  NAND2_X1 U12175 ( .A1(n13156), .A2(n9615), .ZN(n9675) );
  OR2_X1 U12176 ( .A1(n9265), .A2(n13159), .ZN(n9674) );
  INV_X1 U12177 ( .A(P3_REG1_REG_29__SCAN_IN), .ZN(n9678) );
  NAND2_X1 U12178 ( .A1(n11245), .A2(P3_REG2_REG_29__SCAN_IN), .ZN(n9677) );
  NAND2_X1 U12179 ( .A1(n9256), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n9676) );
  OAI211_X1 U12180 ( .C1(n9678), .C2(n9270), .A(n9677), .B(n9676), .ZN(n9679)
         );
  INV_X1 U12181 ( .A(n9679), .ZN(n9680) );
  NAND2_X1 U12182 ( .A1(n9758), .A2(n12859), .ZN(n12660) );
  XNOR2_X1 U12183 ( .A(n9681), .B(n12695), .ZN(n9697) );
  NAND2_X1 U12184 ( .A1(n12722), .A2(n12847), .ZN(n9752) );
  XNOR2_X2 U12185 ( .A(n9686), .B(n9685), .ZN(n11322) );
  NAND2_X1 U12186 ( .A1(n9687), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9688) );
  NAND2_X1 U12187 ( .A1(n12528), .A2(n9765), .ZN(n12715) );
  INV_X4 U12188 ( .A(n12720), .ZN(n13165) );
  OR2_X1 U12189 ( .A1(n13162), .A2(n13165), .ZN(n10534) );
  NAND2_X1 U12190 ( .A1(n10506), .A2(n10534), .ZN(n10706) );
  INV_X1 U12191 ( .A(n10706), .ZN(n10707) );
  INV_X1 U12192 ( .A(P3_REG1_REG_30__SCAN_IN), .ZN(n14821) );
  NAND2_X1 U12193 ( .A1(n11245), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n9691) );
  NAND2_X1 U12194 ( .A1(n9256), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n9690) );
  OAI211_X1 U12195 ( .C1(n9270), .C2(n14821), .A(n9691), .B(n9690), .ZN(n9692)
         );
  INV_X1 U12196 ( .A(n9692), .ZN(n9693) );
  AND2_X1 U12197 ( .A1(n11251), .A2(n9693), .ZN(n12666) );
  INV_X1 U12198 ( .A(P3_B_REG_SCAN_IN), .ZN(n9694) );
  OR2_X1 U12199 ( .A1(n13162), .A2(n9694), .ZN(n9695) );
  NAND2_X1 U12200 ( .A1(n13029), .A2(n9695), .ZN(n12849) );
  OAI22_X1 U12201 ( .A1(n12877), .A2(n15452), .B1(n12666), .B2(n12849), .ZN(
        n9696) );
  NAND2_X1 U12202 ( .A1(n12529), .A2(n12523), .ZN(n10685) );
  NAND2_X1 U12203 ( .A1(n10685), .A2(n12530), .ZN(n15449) );
  NAND2_X1 U12204 ( .A1(n15449), .A2(n15448), .ZN(n15447) );
  INV_X1 U12205 ( .A(n11388), .ZN(n12670) );
  NAND2_X1 U12206 ( .A1(n9699), .A2(n12546), .ZN(n11309) );
  NAND2_X1 U12207 ( .A1(n11309), .A2(n12672), .ZN(n11308) );
  NAND2_X1 U12208 ( .A1(n11308), .A2(n12549), .ZN(n11377) );
  INV_X1 U12209 ( .A(n12676), .ZN(n11376) );
  NAND2_X1 U12210 ( .A1(n11377), .A2(n11376), .ZN(n11375) );
  NAND2_X1 U12211 ( .A1(n11375), .A2(n12556), .ZN(n11403) );
  INV_X1 U12212 ( .A(n11442), .ZN(n12673) );
  NAND2_X1 U12213 ( .A1(n11403), .A2(n12673), .ZN(n11402) );
  NAND2_X1 U12214 ( .A1(n11402), .A2(n12561), .ZN(n11618) );
  NAND2_X1 U12215 ( .A1(n11618), .A2(n12671), .ZN(n11617) );
  NAND2_X1 U12216 ( .A1(n12734), .A2(n15485), .ZN(n9700) );
  INV_X1 U12217 ( .A(n15485), .ZN(n11797) );
  NAND2_X1 U12218 ( .A1(n11871), .A2(n11797), .ZN(n9701) );
  NAND2_X1 U12219 ( .A1(n12113), .A2(n12117), .ZN(n12579) );
  NAND2_X1 U12220 ( .A1(n12416), .A2(n12099), .ZN(n12585) );
  NAND2_X1 U12221 ( .A1(n9703), .A2(n12579), .ZN(n12072) );
  INV_X1 U12222 ( .A(n12592), .ZN(n9704) );
  INV_X1 U12223 ( .A(n12510), .ZN(n13097) );
  XNOR2_X1 U12224 ( .A(n13097), .B(n13028), .ZN(n12686) );
  NAND2_X1 U12225 ( .A1(n13097), .A2(n12599), .ZN(n12603) );
  XNOR2_X1 U12226 ( .A(n13093), .B(n12730), .ZN(n13033) );
  NAND2_X1 U12227 ( .A1(n13093), .A2(n13016), .ZN(n12604) );
  NAND2_X1 U12228 ( .A1(n13021), .A2(n13020), .ZN(n9705) );
  AND2_X1 U12229 ( .A1(n12620), .A2(n12993), .ZN(n12612) );
  NAND2_X1 U12230 ( .A1(n13078), .A2(n12989), .ZN(n9706) );
  INV_X1 U12231 ( .A(n13134), .ZN(n12628) );
  NAND2_X1 U12232 ( .A1(n12628), .A2(n12954), .ZN(n9707) );
  NAND2_X1 U12233 ( .A1(n12958), .A2(n12967), .ZN(n12521) );
  NAND2_X1 U12234 ( .A1(n12957), .A2(n12521), .ZN(n9708) );
  NAND2_X1 U12235 ( .A1(n13122), .A2(n12941), .ZN(n12515) );
  NAND2_X1 U12236 ( .A1(n12458), .A2(n12451), .ZN(n12517) );
  INV_X1 U12237 ( .A(n12646), .ZN(n9710) );
  OAI21_X1 U12238 ( .B1(n11470), .B2(n9765), .A(n12847), .ZN(n9711) );
  NAND2_X1 U12239 ( .A1(n9711), .A2(n11322), .ZN(n9713) );
  OAI21_X1 U12240 ( .B1(n9765), .B2(n12528), .A(n11470), .ZN(n9712) );
  NAND2_X1 U12241 ( .A1(n9713), .A2(n9712), .ZN(n10692) );
  NAND2_X1 U12242 ( .A1(n11242), .A2(n12832), .ZN(n12702) );
  AND2_X1 U12243 ( .A1(n15486), .A2(n9763), .ZN(n9714) );
  NAND2_X1 U12244 ( .A1(n10692), .A2(n9714), .ZN(n9716) );
  AND2_X1 U12245 ( .A1(n9765), .A2(n12832), .ZN(n9715) );
  NAND2_X1 U12246 ( .A1(n12722), .A2(n9715), .ZN(n9764) );
  NAND2_X1 U12247 ( .A1(n9717), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9718) );
  MUX2_X1 U12248 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9718), .S(
        P3_IR_REG_26__SCAN_IN), .Z(n9719) );
  NOR2_X1 U12249 ( .A1(n9721), .A2(n9452), .ZN(n9723) );
  INV_X1 U12250 ( .A(n9725), .ZN(n9726) );
  XNOR2_X1 U12251 ( .A(n12051), .B(P3_B_REG_SCAN_IN), .ZN(n9730) );
  NAND2_X1 U12252 ( .A1(n9725), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9728) );
  MUX2_X1 U12253 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9728), .S(
        P3_IR_REG_25__SCAN_IN), .Z(n9729) );
  NAND2_X1 U12254 ( .A1(n9729), .A2(n9717), .ZN(n12092) );
  INV_X1 U12255 ( .A(P3_D_REG_0__SCAN_IN), .ZN(n9731) );
  NAND2_X1 U12256 ( .A1(n9846), .A2(n9731), .ZN(n9733) );
  NAND2_X1 U12257 ( .A1(n6828), .A2(n12051), .ZN(n9732) );
  INV_X1 U12258 ( .A(n10680), .ZN(n13152) );
  INV_X1 U12259 ( .A(P3_D_REG_1__SCAN_IN), .ZN(n10109) );
  NAND2_X1 U12260 ( .A1(n9846), .A2(n10109), .ZN(n9735) );
  NAND2_X1 U12261 ( .A1(n6828), .A2(n12092), .ZN(n9734) );
  NOR2_X1 U12262 ( .A1(P3_D_REG_5__SCAN_IN), .A2(P3_D_REG_20__SCAN_IN), .ZN(
        n9739) );
  NOR4_X1 U12263 ( .A1(P3_D_REG_2__SCAN_IN), .A2(P3_D_REG_8__SCAN_IN), .A3(
        P3_D_REG_24__SCAN_IN), .A4(P3_D_REG_19__SCAN_IN), .ZN(n9738) );
  NOR4_X1 U12264 ( .A1(P3_D_REG_27__SCAN_IN), .A2(P3_D_REG_29__SCAN_IN), .A3(
        P3_D_REG_10__SCAN_IN), .A4(P3_D_REG_31__SCAN_IN), .ZN(n9737) );
  NOR4_X1 U12265 ( .A1(P3_D_REG_17__SCAN_IN), .A2(P3_D_REG_22__SCAN_IN), .A3(
        P3_D_REG_25__SCAN_IN), .A4(P3_D_REG_18__SCAN_IN), .ZN(n9736) );
  NAND4_X1 U12266 ( .A1(n9739), .A2(n9738), .A3(n9737), .A4(n9736), .ZN(n9745)
         );
  NOR4_X1 U12267 ( .A1(P3_D_REG_26__SCAN_IN), .A2(P3_D_REG_9__SCAN_IN), .A3(
        P3_D_REG_16__SCAN_IN), .A4(P3_D_REG_15__SCAN_IN), .ZN(n9743) );
  NOR4_X1 U12268 ( .A1(P3_D_REG_12__SCAN_IN), .A2(P3_D_REG_14__SCAN_IN), .A3(
        P3_D_REG_21__SCAN_IN), .A4(P3_D_REG_11__SCAN_IN), .ZN(n9742) );
  NOR4_X1 U12269 ( .A1(P3_D_REG_6__SCAN_IN), .A2(P3_D_REG_3__SCAN_IN), .A3(
        P3_D_REG_4__SCAN_IN), .A4(P3_D_REG_7__SCAN_IN), .ZN(n9741) );
  NOR4_X1 U12270 ( .A1(P3_D_REG_30__SCAN_IN), .A2(P3_D_REG_13__SCAN_IN), .A3(
        P3_D_REG_28__SCAN_IN), .A4(P3_D_REG_23__SCAN_IN), .ZN(n9740) );
  NAND4_X1 U12271 ( .A1(n9743), .A2(n9742), .A3(n9741), .A4(n9740), .ZN(n9744)
         );
  OAI21_X1 U12272 ( .B1(n9745), .B2(n9744), .A(n9846), .ZN(n9760) );
  AND3_X1 U12273 ( .A1(n13152), .A2(n13150), .A3(n9760), .ZN(n10700) );
  NOR2_X1 U12274 ( .A1(n12092), .A2(n12051), .ZN(n9746) );
  NAND2_X1 U12275 ( .A1(n9749), .A2(n9748), .ZN(n9750) );
  NAND2_X1 U12276 ( .A1(n9750), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9751) );
  NAND2_X1 U12277 ( .A1(n10702), .A2(n10717), .ZN(n12721) );
  NOR2_X1 U12278 ( .A1(n9752), .A2(n12703), .ZN(n10693) );
  NAND2_X1 U12279 ( .A1(n10702), .A2(n10693), .ZN(n9753) );
  NAND2_X1 U12280 ( .A1(n12721), .A2(n9753), .ZN(n9754) );
  NAND2_X1 U12281 ( .A1(n10700), .A2(n9754), .ZN(n9757) );
  NAND2_X1 U12282 ( .A1(n10680), .A2(n9760), .ZN(n9755) );
  NAND3_X1 U12283 ( .A1(n10705), .A2(n10702), .A3(n10692), .ZN(n9756) );
  INV_X1 U12284 ( .A(n9758), .ZN(n12332) );
  NAND2_X1 U12285 ( .A1(n9759), .A2(n7563), .ZN(P3_U3456) );
  XNOR2_X1 U12286 ( .A(n13150), .B(n10680), .ZN(n9762) );
  AND2_X1 U12287 ( .A1(n9760), .A2(n10702), .ZN(n9761) );
  NAND2_X1 U12288 ( .A1(n12653), .A2(n9764), .ZN(n11360) );
  AND2_X1 U12289 ( .A1(n11359), .A2(n11360), .ZN(n9768) );
  OAI22_X1 U12290 ( .A1(n15486), .A2(n9765), .B1(n12847), .B2(n11470), .ZN(
        n9766) );
  AOI21_X1 U12291 ( .B1(n9766), .B2(n12702), .A(n12647), .ZN(n9767) );
  INV_X1 U12292 ( .A(n13150), .ZN(n11358) );
  MUX2_X1 U12293 ( .A(n9768), .B(n9767), .S(n11358), .Z(n9769) );
  NAND2_X1 U12294 ( .A1(n9770), .A2(n7562), .ZN(P3_U3488) );
  INV_X1 U12295 ( .A(n9771), .ZN(n9772) );
  NOR2_X1 U12296 ( .A1(n10631), .A2(n9772), .ZN(P2_U3947) );
  NAND2_X1 U12297 ( .A1(n14169), .A2(n9773), .ZN(n9774) );
  NAND2_X1 U12298 ( .A1(n9775), .A2(n9774), .ZN(n9784) );
  NAND2_X1 U12299 ( .A1(n9784), .A2(n15162), .ZN(n9779) );
  AOI22_X1 U12300 ( .A1(n14230), .A2(n14583), .B1(n14921), .B2(n14233), .ZN(
        n9778) );
  XNOR2_X1 U12301 ( .A(n14169), .B(n13966), .ZN(n9776) );
  NAND2_X1 U12302 ( .A1(n9776), .A2(n14952), .ZN(n9777) );
  NAND3_X1 U12303 ( .A1(n9779), .A2(n9778), .A3(n9777), .ZN(n10554) );
  NAND2_X1 U12304 ( .A1(n10419), .A2(n10402), .ZN(n9781) );
  OR3_X1 U12305 ( .A1(n9781), .A2(n9780), .A3(n10405), .ZN(n14360) );
  INV_X1 U12306 ( .A(n10412), .ZN(n9782) );
  INV_X1 U12307 ( .A(n10406), .ZN(n9812) );
  MUX2_X1 U12308 ( .A(n10554), .B(P1_REG2_REG_1__SCAN_IN), .S(n15105), .Z(
        n9790) );
  OAI22_X1 U12309 ( .A1(n14570), .A2(n10561), .B1(n9783), .B2(n14602), .ZN(
        n9789) );
  INV_X1 U12310 ( .A(n9784), .ZN(n10557) );
  INV_X1 U12311 ( .A(n10390), .ZN(n9785) );
  OR2_X1 U12312 ( .A1(n9785), .A2(n14917), .ZN(n13951) );
  INV_X1 U12313 ( .A(n13951), .ZN(n9786) );
  NAND2_X1 U12314 ( .A1(n14539), .A2(n9786), .ZN(n15082) );
  OAI21_X1 U12315 ( .B1(n10561), .B2(n10389), .A(n15086), .ZN(n9787) );
  OR2_X1 U12316 ( .A1(n11064), .A2(n9787), .ZN(n10555) );
  OAI22_X1 U12317 ( .A1(n10557), .A2(n15082), .B1(n14557), .B2(n10555), .ZN(
        n9788) );
  OR3_X1 U12318 ( .A1(n9790), .A2(n9789), .A3(n9788), .ZN(P1_U3292) );
  OAI211_X1 U12319 ( .C1(n10648), .C2(n10639), .A(n13604), .B(n13652), .ZN(
        n10586) );
  OR3_X1 U12320 ( .A1(n6620), .A2(n9791), .A3(n11531), .ZN(n11588) );
  OAI21_X1 U12321 ( .B1(n9794), .B2(n9793), .A(n9792), .ZN(n10589) );
  INV_X1 U12322 ( .A(n10589), .ZN(n9801) );
  OAI22_X1 U12323 ( .A1(n13612), .A2(n10586), .B1(n11588), .B2(n9801), .ZN(
        n9804) );
  OAI21_X1 U12324 ( .B1(n9797), .B2(n9796), .A(n9795), .ZN(n9799) );
  OAI22_X1 U12325 ( .A1(n10598), .A2(n13301), .B1(n9798), .B2(n13303), .ZN(
        n10635) );
  AOI21_X1 U12326 ( .B1(n9799), .B2(n13661), .A(n10635), .ZN(n9800) );
  OAI21_X1 U12327 ( .B1(n9801), .B2(n8816), .A(n9800), .ZN(n10587) );
  MUX2_X1 U12328 ( .A(n10587), .B(P2_REG2_REG_1__SCAN_IN), .S(n6620), .Z(n9803) );
  INV_X1 U12329 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n15211) );
  OAI22_X1 U12330 ( .A1(n15330), .A2(n10648), .B1(n15211), .B2(n13655), .ZN(
        n9802) );
  OR3_X1 U12331 ( .A1(n9804), .A2(n9803), .A3(n9802), .ZN(P2_U3264) );
  INV_X1 U12332 ( .A(n9805), .ZN(n9807) );
  INV_X2 U12333 ( .A(n13792), .ZN(n13804) );
  NOR2_X1 U12334 ( .A1(n7088), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13786) );
  AND2_X1 U12335 ( .A1(n10315), .A2(P2_STATE_REG_SCAN_IN), .ZN(n15235) );
  AOI21_X1 U12336 ( .B1(n13786), .B2(P1_DATAO_REG_3__SCAN_IN), .A(n15235), 
        .ZN(n9806) );
  OAI21_X1 U12337 ( .B1(n9807), .B2(n13804), .A(n9806), .ZN(P2_U3324) );
  INV_X1 U12338 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n9808) );
  NOR2_X1 U12339 ( .A1(n7088), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14757) );
  INV_X2 U12340 ( .A(n14757), .ZN(n14761) );
  INV_X1 U12341 ( .A(n14252), .ZN(n9928) );
  INV_X1 U12342 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n9809) );
  INV_X1 U12343 ( .A(n9810), .ZN(n9823) );
  OAI222_X1 U12344 ( .A1(P1_U3086), .A2(n9923), .B1(n14761), .B2(n8380), .C1(
        n7718), .C2(n14774), .ZN(P1_U3354) );
  NAND2_X1 U12345 ( .A1(n9813), .A2(n9812), .ZN(n15109) );
  INV_X1 U12346 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n9817) );
  NOR3_X1 U12347 ( .A1(n9815), .A2(n8325), .A3(n9814), .ZN(n9816) );
  AOI21_X1 U12348 ( .B1(n15109), .B2(n9817), .A(n9816), .ZN(P1_U3446) );
  OAI222_X1 U12349 ( .A1(n13804), .A2(n9819), .B1(n15223), .B2(P2_U3088), .C1(
        n9818), .C2(n13798), .ZN(P2_U3325) );
  OAI222_X1 U12350 ( .A1(n13804), .A2(n8380), .B1(n10313), .B2(P2_U3088), .C1(
        n9820), .C2(n13798), .ZN(P2_U3326) );
  OAI222_X1 U12351 ( .A1(n13804), .A2(n9834), .B1(n10359), .B2(P2_U3088), .C1(
        n9821), .C2(n13798), .ZN(P2_U3322) );
  INV_X1 U12352 ( .A(n10316), .ZN(n10329) );
  OAI222_X1 U12353 ( .A1(n13804), .A2(n9823), .B1(n10329), .B2(P2_U3088), .C1(
        n9822), .C2(n13798), .ZN(P2_U3323) );
  INV_X1 U12354 ( .A(n9824), .ZN(n9826) );
  AOI22_X1 U12355 ( .A1(n15109), .A2(n9827), .B1(n9826), .B2(n9825), .ZN(
        P1_U3445) );
  INV_X1 U12356 ( .A(n10344), .ZN(n10336) );
  OAI222_X1 U12357 ( .A1(n13804), .A2(n9832), .B1(n10336), .B2(P2_U3088), .C1(
        n9828), .C2(n13798), .ZN(P2_U3321) );
  NOR2_X1 U12358 ( .A1(n7088), .A2(P3_STATE_REG_SCAN_IN), .ZN(n14796) );
  INV_X2 U12359 ( .A(n14796), .ZN(n13172) );
  INV_X1 U12360 ( .A(n9829), .ZN(n9831) );
  OAI222_X1 U12361 ( .A1(n13172), .A2(n9831), .B1(n13167), .B2(n9830), .C1(
        P3_U3151), .C2(n10511), .ZN(P3_U3294) );
  INV_X1 U12362 ( .A(n10376), .ZN(n10383) );
  INV_X1 U12363 ( .A(n14266), .ZN(n9931) );
  INV_X1 U12364 ( .A(n11659), .ZN(n11669) );
  INV_X1 U12365 ( .A(SI_9_), .ZN(n9836) );
  OAI222_X1 U12366 ( .A1(P3_U3151), .A2(n11669), .B1(n13167), .B2(n9836), .C1(
        n13172), .C2(n9835), .ZN(P3_U3286) );
  INV_X1 U12367 ( .A(n11675), .ZN(n11713) );
  OAI222_X1 U12368 ( .A1(P3_U3151), .A2(n11713), .B1(n13167), .B2(n9838), .C1(
        n13172), .C2(n9837), .ZN(P3_U3284) );
  INV_X1 U12369 ( .A(SI_7_), .ZN(n9840) );
  OAI222_X1 U12370 ( .A1(P3_U3151), .A2(n10900), .B1(n13167), .B2(n9840), .C1(
        n13172), .C2(n9839), .ZN(P3_U3288) );
  INV_X1 U12371 ( .A(n9841), .ZN(n9843) );
  INV_X1 U12372 ( .A(n13167), .ZN(n14795) );
  OAI222_X1 U12373 ( .A1(n13172), .A2(n9843), .B1(n13167), .B2(n9842), .C1(
        P3_U3151), .C2(n11076), .ZN(P3_U3287) );
  INV_X1 U12374 ( .A(SI_10_), .ZN(n9845) );
  OAI222_X1 U12375 ( .A1(P3_U3151), .A2(n11661), .B1(n13167), .B2(n9845), .C1(
        n13172), .C2(n9844), .ZN(P3_U3285) );
  NOR2_X1 U12376 ( .A1(n9846), .A2(n13149), .ZN(n9854) );
  INV_X1 U12377 ( .A(P3_D_REG_26__SCAN_IN), .ZN(n9847) );
  NOR2_X1 U12378 ( .A1(n9874), .A2(n9847), .ZN(P3_U3239) );
  INV_X1 U12379 ( .A(P3_D_REG_29__SCAN_IN), .ZN(n9848) );
  NOR2_X1 U12380 ( .A1(n9854), .A2(n9848), .ZN(P3_U3236) );
  INV_X1 U12381 ( .A(P3_D_REG_30__SCAN_IN), .ZN(n9849) );
  NOR2_X1 U12382 ( .A1(n9854), .A2(n9849), .ZN(P3_U3235) );
  INV_X1 U12383 ( .A(P3_D_REG_28__SCAN_IN), .ZN(n9850) );
  NOR2_X1 U12384 ( .A1(n9854), .A2(n9850), .ZN(P3_U3237) );
  INV_X1 U12385 ( .A(P3_D_REG_24__SCAN_IN), .ZN(n10149) );
  NOR2_X1 U12386 ( .A1(n9854), .A2(n10149), .ZN(P3_U3241) );
  INV_X1 U12387 ( .A(P3_D_REG_25__SCAN_IN), .ZN(n9851) );
  NOR2_X1 U12388 ( .A1(n9854), .A2(n9851), .ZN(P3_U3240) );
  INV_X1 U12389 ( .A(P3_D_REG_21__SCAN_IN), .ZN(n9852) );
  NOR2_X1 U12390 ( .A1(n9854), .A2(n9852), .ZN(P3_U3244) );
  INV_X1 U12391 ( .A(P3_D_REG_27__SCAN_IN), .ZN(n9853) );
  NOR2_X1 U12392 ( .A1(n9854), .A2(n9853), .ZN(P3_U3238) );
  INV_X1 U12393 ( .A(P3_D_REG_20__SCAN_IN), .ZN(n10147) );
  NOR2_X1 U12394 ( .A1(n9854), .A2(n10147), .ZN(P3_U3245) );
  CLKBUF_X1 U12395 ( .A(n9854), .Z(n9874) );
  INV_X1 U12396 ( .A(P3_D_REG_19__SCAN_IN), .ZN(n10220) );
  NOR2_X1 U12397 ( .A1(n9874), .A2(n10220), .ZN(P3_U3246) );
  INV_X1 U12398 ( .A(P3_D_REG_18__SCAN_IN), .ZN(n9855) );
  NOR2_X1 U12399 ( .A1(n9874), .A2(n9855), .ZN(P3_U3247) );
  INV_X1 U12400 ( .A(P3_D_REG_31__SCAN_IN), .ZN(n9856) );
  NOR2_X1 U12401 ( .A1(n9854), .A2(n9856), .ZN(P3_U3234) );
  INV_X1 U12402 ( .A(P3_D_REG_23__SCAN_IN), .ZN(n9857) );
  NOR2_X1 U12403 ( .A1(n9854), .A2(n9857), .ZN(P3_U3242) );
  INV_X1 U12404 ( .A(P3_D_REG_15__SCAN_IN), .ZN(n9858) );
  NOR2_X1 U12405 ( .A1(n9874), .A2(n9858), .ZN(P3_U3250) );
  INV_X1 U12406 ( .A(P3_D_REG_14__SCAN_IN), .ZN(n9859) );
  NOR2_X1 U12407 ( .A1(n9874), .A2(n9859), .ZN(P3_U3251) );
  INV_X1 U12408 ( .A(P3_D_REG_13__SCAN_IN), .ZN(n9860) );
  NOR2_X1 U12409 ( .A1(n9874), .A2(n9860), .ZN(P3_U3252) );
  INV_X1 U12410 ( .A(P3_D_REG_12__SCAN_IN), .ZN(n9861) );
  NOR2_X1 U12411 ( .A1(n9874), .A2(n9861), .ZN(P3_U3253) );
  INV_X1 U12412 ( .A(P3_D_REG_11__SCAN_IN), .ZN(n9862) );
  NOR2_X1 U12413 ( .A1(n9874), .A2(n9862), .ZN(P3_U3254) );
  INV_X1 U12414 ( .A(P3_D_REG_10__SCAN_IN), .ZN(n9863) );
  NOR2_X1 U12415 ( .A1(n9874), .A2(n9863), .ZN(P3_U3255) );
  INV_X1 U12416 ( .A(P3_D_REG_9__SCAN_IN), .ZN(n9864) );
  NOR2_X1 U12417 ( .A1(n9874), .A2(n9864), .ZN(P3_U3256) );
  INV_X1 U12418 ( .A(P3_D_REG_8__SCAN_IN), .ZN(n9865) );
  NOR2_X1 U12419 ( .A1(n9874), .A2(n9865), .ZN(P3_U3257) );
  INV_X1 U12420 ( .A(P3_D_REG_7__SCAN_IN), .ZN(n9866) );
  NOR2_X1 U12421 ( .A1(n9854), .A2(n9866), .ZN(P3_U3258) );
  INV_X1 U12422 ( .A(P3_D_REG_6__SCAN_IN), .ZN(n9867) );
  NOR2_X1 U12423 ( .A1(n9874), .A2(n9867), .ZN(P3_U3259) );
  INV_X1 U12424 ( .A(P3_D_REG_22__SCAN_IN), .ZN(n9868) );
  NOR2_X1 U12425 ( .A1(n9874), .A2(n9868), .ZN(P3_U3243) );
  INV_X1 U12426 ( .A(P3_D_REG_5__SCAN_IN), .ZN(n10102) );
  NOR2_X1 U12427 ( .A1(n9874), .A2(n10102), .ZN(P3_U3260) );
  INV_X1 U12428 ( .A(P3_D_REG_4__SCAN_IN), .ZN(n9869) );
  NOR2_X1 U12429 ( .A1(n9874), .A2(n9869), .ZN(P3_U3261) );
  INV_X1 U12430 ( .A(P3_D_REG_3__SCAN_IN), .ZN(n9870) );
  NOR2_X1 U12431 ( .A1(n9874), .A2(n9870), .ZN(P3_U3262) );
  INV_X1 U12432 ( .A(P3_D_REG_2__SCAN_IN), .ZN(n9871) );
  NOR2_X1 U12433 ( .A1(n9874), .A2(n9871), .ZN(P3_U3263) );
  INV_X1 U12434 ( .A(P3_D_REG_17__SCAN_IN), .ZN(n9872) );
  NOR2_X1 U12435 ( .A1(n9874), .A2(n9872), .ZN(P3_U3248) );
  INV_X1 U12436 ( .A(P3_D_REG_16__SCAN_IN), .ZN(n9873) );
  NOR2_X1 U12437 ( .A1(n9874), .A2(n9873), .ZN(P3_U3249) );
  INV_X1 U12438 ( .A(n9875), .ZN(n9876) );
  OAI222_X1 U12439 ( .A1(n13167), .A2(n9877), .B1(n13172), .B2(n9876), .C1(
        n11891), .C2(P3_U3151), .ZN(P3_U3283) );
  INV_X1 U12440 ( .A(n9878), .ZN(n9880) );
  OAI222_X1 U12441 ( .A1(P3_U3151), .A2(n10849), .B1(n13172), .B2(n9880), .C1(
        n9879), .C2(n13167), .ZN(P3_U3289) );
  OAI222_X1 U12442 ( .A1(n10874), .A2(P3_U3151), .B1(n13172), .B2(n9881), .C1(
        n10076), .C2(n13167), .ZN(P3_U3290) );
  INV_X1 U12443 ( .A(n10533), .ZN(n10584) );
  INV_X1 U12444 ( .A(SI_2_), .ZN(n9882) );
  OAI222_X1 U12445 ( .A1(n10584), .A2(P3_U3151), .B1(n13172), .B2(n9883), .C1(
        n9882), .C2(n13167), .ZN(P3_U3293) );
  INV_X1 U12446 ( .A(n9884), .ZN(n9886) );
  OAI222_X1 U12447 ( .A1(P3_U3151), .A2(n10529), .B1(n13172), .B2(n9886), .C1(
        n9885), .C2(n13167), .ZN(P3_U3295) );
  INV_X1 U12448 ( .A(n10798), .ZN(n10805) );
  INV_X1 U12449 ( .A(SI_3_), .ZN(n10178) );
  OAI222_X1 U12450 ( .A1(n10805), .A2(P3_U3151), .B1(n13172), .B2(n9887), .C1(
        n10178), .C2(n13167), .ZN(P3_U3292) );
  INV_X1 U12451 ( .A(n15410), .ZN(n10807) );
  INV_X1 U12452 ( .A(SI_4_), .ZN(n9888) );
  OAI222_X1 U12453 ( .A1(n10807), .A2(P3_U3151), .B1(n13172), .B2(n9889), .C1(
        n9888), .C2(n13167), .ZN(P3_U3291) );
  INV_X1 U12454 ( .A(n13392), .ZN(n9891) );
  INV_X1 U12455 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n9890) );
  OAI222_X1 U12456 ( .A1(n13804), .A2(n9892), .B1(n9891), .B2(P2_U3088), .C1(
        n9890), .C2(n13798), .ZN(P2_U3320) );
  INV_X1 U12457 ( .A(n10989), .ZN(n10983) );
  INV_X1 U12458 ( .A(n10477), .ZN(n10341) );
  INV_X1 U12459 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n9894) );
  OAI222_X1 U12460 ( .A1(n13804), .A2(n9895), .B1(n10341), .B2(P2_U3088), .C1(
        n9894), .C2(n13798), .ZN(P2_U3319) );
  OAI222_X1 U12461 ( .A1(n11931), .A2(P3_U3151), .B1(n13172), .B2(n9898), .C1(
        n9897), .C2(n13167), .ZN(P3_U3282) );
  INV_X1 U12462 ( .A(n15253), .ZN(n9900) );
  INV_X1 U12463 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n9899) );
  OAI222_X1 U12464 ( .A1(n13804), .A2(n9901), .B1(n9900), .B2(P2_U3088), .C1(
        n9899), .C2(n13798), .ZN(P2_U3318) );
  INV_X1 U12465 ( .A(n14294), .ZN(n10984) );
  INV_X1 U12466 ( .A(n12746), .ZN(n12756) );
  OAI222_X1 U12467 ( .A1(P3_U3151), .A2(n12756), .B1(n13167), .B2(n10197), 
        .C1(n13172), .C2(n9903), .ZN(P3_U3281) );
  INV_X1 U12468 ( .A(n10413), .ZN(n9904) );
  NAND2_X1 U12469 ( .A1(n9904), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14209) );
  NAND2_X1 U12470 ( .A1(n10406), .A2(n14209), .ZN(n9910) );
  NAND2_X1 U12471 ( .A1(n10407), .A2(n10413), .ZN(n9906) );
  AND2_X1 U12472 ( .A1(n9906), .A2(n9905), .ZN(n9909) );
  INV_X1 U12473 ( .A(n9909), .ZN(n9907) );
  AND2_X1 U12474 ( .A1(n9910), .A2(n9907), .ZN(n14981) );
  NOR2_X1 U12475 ( .A1(n14981), .A2(P1_U4016), .ZN(P1_U3085) );
  INV_X1 U12476 ( .A(P3_DATAO_REG_13__SCAN_IN), .ZN(n10198) );
  NAND2_X1 U12477 ( .A1(n12419), .A2(P3_U3897), .ZN(n9908) );
  OAI21_X1 U12478 ( .B1(P3_U3897), .B2(n10198), .A(n9908), .ZN(P3_U3504) );
  NAND2_X1 U12479 ( .A1(n9910), .A2(n9909), .ZN(n14983) );
  NAND2_X1 U12480 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_U3086), .ZN(n9911) );
  OAI21_X1 U12481 ( .B1(n15070), .B2(n9912), .A(n9911), .ZN(n9922) );
  MUX2_X1 U12482 ( .A(n9913), .B(P1_REG1_REG_6__SCAN_IN), .S(n10376), .Z(n9920) );
  INV_X1 U12483 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n10560) );
  MUX2_X1 U12484 ( .A(n10560), .B(P1_REG1_REG_1__SCAN_IN), .S(n9923), .Z(
        n14239) );
  AND2_X1 U12485 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n14238) );
  NAND2_X1 U12486 ( .A1(n14239), .A2(n14238), .ZN(n14237) );
  INV_X1 U12487 ( .A(n9923), .ZN(n14240) );
  NAND2_X1 U12488 ( .A1(n14240), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n9914) );
  NAND2_X1 U12489 ( .A1(n14237), .A2(n9914), .ZN(n10444) );
  INV_X1 U12490 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n15175) );
  MUX2_X1 U12491 ( .A(n15175), .B(P1_REG1_REG_2__SCAN_IN), .S(n9926), .Z(
        n10445) );
  NAND2_X1 U12492 ( .A1(n10444), .A2(n10445), .ZN(n10443) );
  INV_X1 U12493 ( .A(n10443), .ZN(n9915) );
  XNOR2_X1 U12494 ( .A(n14252), .B(P1_REG1_REG_3__SCAN_IN), .ZN(n14246) );
  NOR2_X1 U12495 ( .A1(n14247), .A2(n14246), .ZN(n14245) );
  MUX2_X1 U12496 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n9916), .S(n10465), .Z(
        n10458) );
  NOR2_X1 U12497 ( .A1(n10459), .A2(n10458), .ZN(n10457) );
  MUX2_X1 U12498 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n9918), .S(n14266), .Z(
        n14260) );
  NAND2_X1 U12499 ( .A1(n14261), .A2(n14260), .ZN(n14259) );
  OAI21_X1 U12500 ( .B1(P1_REG1_REG_5__SCAN_IN), .B2(n14266), .A(n14259), .ZN(
        n9919) );
  INV_X1 U12501 ( .A(n6625), .ZN(n14978) );
  OR2_X1 U12502 ( .A1(n14983), .A2(n14978), .ZN(n15056) );
  NOR2_X1 U12503 ( .A1(n9919), .A2(n9920), .ZN(n10375) );
  AOI211_X1 U12504 ( .C1(n9920), .C2(n9919), .A(n15056), .B(n10375), .ZN(n9921) );
  AOI211_X1 U12505 ( .C1(n15067), .C2(n10376), .A(n9922), .B(n9921), .ZN(n9936) );
  MUX2_X1 U12506 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n10384), .S(n10376), .Z(
        n9934) );
  INV_X1 U12507 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n9924) );
  MUX2_X1 U12508 ( .A(n9924), .B(P1_REG2_REG_1__SCAN_IN), .S(n9923), .Z(n14236) );
  AND2_X1 U12509 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n14235) );
  NAND2_X1 U12510 ( .A1(n14236), .A2(n14235), .ZN(n14234) );
  NAND2_X1 U12511 ( .A1(n14240), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n9925) );
  NAND2_X1 U12512 ( .A1(n14234), .A2(n9925), .ZN(n10447) );
  MUX2_X1 U12513 ( .A(n9927), .B(P1_REG2_REG_2__SCAN_IN), .S(n9926), .Z(n10448) );
  NAND2_X1 U12514 ( .A1(n10447), .A2(n10448), .ZN(n10446) );
  OAI21_X1 U12515 ( .B1(n9927), .B2(n9926), .A(n10446), .ZN(n14254) );
  XOR2_X1 U12516 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n14252), .Z(n14255) );
  NAND2_X1 U12517 ( .A1(n14254), .A2(n14255), .ZN(n14253) );
  OAI21_X1 U12518 ( .B1(n11032), .B2(n9928), .A(n14253), .ZN(n10462) );
  MUX2_X1 U12519 ( .A(n9929), .B(P1_REG2_REG_4__SCAN_IN), .S(n10465), .Z(
        n10463) );
  NAND2_X1 U12520 ( .A1(n10462), .A2(n10463), .ZN(n10461) );
  OAI21_X1 U12521 ( .B1(n10465), .B2(n9929), .A(n10461), .ZN(n14268) );
  MUX2_X1 U12522 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n9930), .S(n14266), .Z(
        n14269) );
  NAND2_X1 U12523 ( .A1(n14268), .A2(n14269), .ZN(n14267) );
  OAI21_X1 U12524 ( .B1(n9931), .B2(n9930), .A(n14267), .ZN(n9933) );
  OR2_X1 U12525 ( .A1(n12173), .A2(n6625), .ZN(n9932) );
  OR2_X1 U12526 ( .A1(n14983), .A2(n9932), .ZN(n15060) );
  NAND2_X1 U12527 ( .A1(n9933), .A2(n9934), .ZN(n10382) );
  OAI211_X1 U12528 ( .C1(n9934), .C2(n9933), .A(n15012), .B(n10382), .ZN(n9935) );
  NAND2_X1 U12529 ( .A1(n9936), .A2(n9935), .ZN(P1_U3249) );
  INV_X1 U12530 ( .A(n15264), .ZN(n9938) );
  INV_X1 U12531 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n9937) );
  OAI222_X1 U12532 ( .A1(n13804), .A2(n9939), .B1(n9938), .B2(P2_U3088), .C1(
        n9937), .C2(n13798), .ZN(P2_U3317) );
  INV_X1 U12533 ( .A(n11104), .ZN(n10997) );
  INV_X1 U12534 ( .A(P3_DATAO_REG_11__SCAN_IN), .ZN(n10233) );
  NAND2_X1 U12535 ( .A1(n12416), .A2(P3_U3897), .ZN(n9940) );
  OAI21_X1 U12536 ( .B1(P3_U3897), .B2(n10233), .A(n9940), .ZN(P3_U3502) );
  AOI21_X1 U12537 ( .B1(n14949), .B2(n15075), .A(n15098), .ZN(n9943) );
  NOR2_X1 U12538 ( .A1(n10389), .A2(n9942), .ZN(n15097) );
  NOR3_X1 U12539 ( .A1(n9943), .A2(n15095), .A3(n15097), .ZN(n9946) );
  NAND2_X1 U12540 ( .A1(n15172), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n9944) );
  OAI21_X1 U12541 ( .B1(n9946), .B2(n15172), .A(n9944), .ZN(P1_U3459) );
  NAND2_X1 U12542 ( .A1(n15183), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n9945) );
  OAI21_X1 U12543 ( .B1(n9946), .B2(n15183), .A(n9945), .ZN(P1_U3528) );
  INV_X2 U12544 ( .A(P3_U3897), .ZN(n12740) );
  MUX2_X1 U12545 ( .A(n11788), .B(P3_DATAO_REG_8__SCAN_IN), .S(n12740), .Z(
        n10288) );
  OAI22_X1 U12546 ( .A1(P3_REG2_REG_18__SCAN_IN), .A2(keyinput92), .B1(
        P3_REG0_REG_13__SCAN_IN), .B2(keyinput69), .ZN(n9947) );
  AOI221_X1 U12547 ( .B1(P3_REG2_REG_18__SCAN_IN), .B2(keyinput92), .C1(
        keyinput69), .C2(P3_REG0_REG_13__SCAN_IN), .A(n9947), .ZN(n9954) );
  OAI22_X1 U12548 ( .A1(P3_REG1_REG_3__SCAN_IN), .A2(keyinput52), .B1(
        P2_REG2_REG_30__SCAN_IN), .B2(keyinput83), .ZN(n9948) );
  AOI221_X1 U12549 ( .B1(P3_REG1_REG_3__SCAN_IN), .B2(keyinput52), .C1(
        keyinput83), .C2(P2_REG2_REG_30__SCAN_IN), .A(n9948), .ZN(n9953) );
  OAI22_X1 U12550 ( .A1(P2_REG1_REG_0__SCAN_IN), .A2(keyinput116), .B1(
        P1_REG2_REG_19__SCAN_IN), .B2(keyinput126), .ZN(n9949) );
  AOI221_X1 U12551 ( .B1(P2_REG1_REG_0__SCAN_IN), .B2(keyinput116), .C1(
        keyinput126), .C2(P1_REG2_REG_19__SCAN_IN), .A(n9949), .ZN(n9952) );
  OAI22_X1 U12552 ( .A1(P2_REG0_REG_24__SCAN_IN), .A2(keyinput70), .B1(
        P1_REG2_REG_20__SCAN_IN), .B2(keyinput57), .ZN(n9950) );
  AOI221_X1 U12553 ( .B1(P2_REG0_REG_24__SCAN_IN), .B2(keyinput70), .C1(
        keyinput57), .C2(P1_REG2_REG_20__SCAN_IN), .A(n9950), .ZN(n9951) );
  NAND4_X1 U12554 ( .A1(n9954), .A2(n9953), .A3(n9952), .A4(n9951), .ZN(n9982)
         );
  OAI22_X1 U12555 ( .A1(P2_REG3_REG_28__SCAN_IN), .A2(keyinput15), .B1(
        keyinput4), .B2(P2_REG1_REG_19__SCAN_IN), .ZN(n9955) );
  AOI221_X1 U12556 ( .B1(P2_REG3_REG_28__SCAN_IN), .B2(keyinput15), .C1(
        P2_REG1_REG_19__SCAN_IN), .C2(keyinput4), .A(n9955), .ZN(n9962) );
  OAI22_X1 U12557 ( .A1(P3_REG3_REG_17__SCAN_IN), .A2(keyinput101), .B1(
        keyinput118), .B2(P2_IR_REG_11__SCAN_IN), .ZN(n9956) );
  AOI221_X1 U12558 ( .B1(P3_REG3_REG_17__SCAN_IN), .B2(keyinput101), .C1(
        P2_IR_REG_11__SCAN_IN), .C2(keyinput118), .A(n9956), .ZN(n9961) );
  OAI22_X1 U12559 ( .A1(P3_D_REG_1__SCAN_IN), .A2(keyinput18), .B1(
        P1_D_REG_0__SCAN_IN), .B2(keyinput68), .ZN(n9957) );
  AOI221_X1 U12560 ( .B1(P3_D_REG_1__SCAN_IN), .B2(keyinput18), .C1(keyinput68), .C2(P1_D_REG_0__SCAN_IN), .A(n9957), .ZN(n9960) );
  OAI22_X1 U12561 ( .A1(P3_REG2_REG_19__SCAN_IN), .A2(keyinput19), .B1(
        keyinput94), .B2(P2_REG1_REG_22__SCAN_IN), .ZN(n9958) );
  AOI221_X1 U12562 ( .B1(P3_REG2_REG_19__SCAN_IN), .B2(keyinput19), .C1(
        P2_REG1_REG_22__SCAN_IN), .C2(keyinput94), .A(n9958), .ZN(n9959) );
  NAND4_X1 U12563 ( .A1(n9962), .A2(n9961), .A3(n9960), .A4(n9959), .ZN(n9981)
         );
  OAI22_X1 U12564 ( .A1(P2_REG1_REG_8__SCAN_IN), .A2(keyinput27), .B1(
        P3_WR_REG_SCAN_IN), .B2(keyinput80), .ZN(n9963) );
  AOI221_X1 U12565 ( .B1(P2_REG1_REG_8__SCAN_IN), .B2(keyinput27), .C1(
        keyinput80), .C2(P3_WR_REG_SCAN_IN), .A(n9963), .ZN(n9970) );
  OAI22_X1 U12566 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(keyinput119), .B1(
        keyinput1), .B2(P1_REG1_REG_20__SCAN_IN), .ZN(n9964) );
  AOI221_X1 U12567 ( .B1(P1_REG3_REG_9__SCAN_IN), .B2(keyinput119), .C1(
        P1_REG1_REG_20__SCAN_IN), .C2(keyinput1), .A(n9964), .ZN(n9969) );
  OAI22_X1 U12568 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(keyinput74), .B1(
        keyinput49), .B2(P3_REG1_REG_8__SCAN_IN), .ZN(n9965) );
  AOI221_X1 U12569 ( .B1(P1_DATAO_REG_21__SCAN_IN), .B2(keyinput74), .C1(
        P3_REG1_REG_8__SCAN_IN), .C2(keyinput49), .A(n9965), .ZN(n9968) );
  OAI22_X1 U12570 ( .A1(P2_DATAO_REG_17__SCAN_IN), .A2(keyinput112), .B1(
        keyinput34), .B2(P1_IR_REG_12__SCAN_IN), .ZN(n9966) );
  AOI221_X1 U12571 ( .B1(P2_DATAO_REG_17__SCAN_IN), .B2(keyinput112), .C1(
        P1_IR_REG_12__SCAN_IN), .C2(keyinput34), .A(n9966), .ZN(n9967) );
  NAND4_X1 U12572 ( .A1(n9970), .A2(n9969), .A3(n9968), .A4(n9967), .ZN(n9980)
         );
  OAI22_X1 U12573 ( .A1(P3_REG2_REG_25__SCAN_IN), .A2(keyinput14), .B1(
        keyinput117), .B2(P2_REG2_REG_10__SCAN_IN), .ZN(n9971) );
  AOI221_X1 U12574 ( .B1(P3_REG2_REG_25__SCAN_IN), .B2(keyinput14), .C1(
        P2_REG2_REG_10__SCAN_IN), .C2(keyinput117), .A(n9971), .ZN(n9978) );
  OAI22_X1 U12575 ( .A1(SI_5_), .A2(keyinput42), .B1(P1_REG1_REG_5__SCAN_IN), 
        .B2(keyinput30), .ZN(n9972) );
  AOI221_X1 U12576 ( .B1(SI_5_), .B2(keyinput42), .C1(keyinput30), .C2(
        P1_REG1_REG_5__SCAN_IN), .A(n9972), .ZN(n9977) );
  OAI22_X1 U12577 ( .A1(P3_REG2_REG_5__SCAN_IN), .A2(keyinput76), .B1(
        keyinput51), .B2(P1_REG3_REG_27__SCAN_IN), .ZN(n9973) );
  AOI221_X1 U12578 ( .B1(P3_REG2_REG_5__SCAN_IN), .B2(keyinput76), .C1(
        P1_REG3_REG_27__SCAN_IN), .C2(keyinput51), .A(n9973), .ZN(n9976) );
  OAI22_X1 U12579 ( .A1(P2_D_REG_14__SCAN_IN), .A2(keyinput125), .B1(
        keyinput37), .B2(P1_REG1_REG_10__SCAN_IN), .ZN(n9974) );
  AOI221_X1 U12580 ( .B1(P2_D_REG_14__SCAN_IN), .B2(keyinput125), .C1(
        P1_REG1_REG_10__SCAN_IN), .C2(keyinput37), .A(n9974), .ZN(n9975) );
  NAND4_X1 U12581 ( .A1(n9978), .A2(n9977), .A3(n9976), .A4(n9975), .ZN(n9979)
         );
  NOR4_X1 U12582 ( .A1(n9982), .A2(n9981), .A3(n9980), .A4(n9979), .ZN(n10286)
         );
  AOI22_X1 U12583 ( .A1(P3_REG0_REG_13__SCAN_IN), .A2(keyinput197), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(keyinput218), .ZN(n9983) );
  OAI221_X1 U12584 ( .B1(P3_REG0_REG_13__SCAN_IN), .B2(keyinput197), .C1(
        P2_DATAO_REG_13__SCAN_IN), .C2(keyinput218), .A(n9983), .ZN(n9990) );
  AOI22_X1 U12585 ( .A1(P1_REG1_REG_11__SCAN_IN), .A2(keyinput138), .B1(
        P3_REG2_REG_10__SCAN_IN), .B2(keyinput231), .ZN(n9984) );
  OAI221_X1 U12586 ( .B1(P1_REG1_REG_11__SCAN_IN), .B2(keyinput138), .C1(
        P3_REG2_REG_10__SCAN_IN), .C2(keyinput231), .A(n9984), .ZN(n9989) );
  AOI22_X1 U12587 ( .A1(P1_REG0_REG_2__SCAN_IN), .A2(keyinput153), .B1(
        P2_D_REG_23__SCAN_IN), .B2(keyinput248), .ZN(n9985) );
  OAI221_X1 U12588 ( .B1(P1_REG0_REG_2__SCAN_IN), .B2(keyinput153), .C1(
        P2_D_REG_23__SCAN_IN), .C2(keyinput248), .A(n9985), .ZN(n9988) );
  AOI22_X1 U12589 ( .A1(P2_REG1_REG_8__SCAN_IN), .A2(keyinput155), .B1(
        P2_D_REG_28__SCAN_IN), .B2(keyinput201), .ZN(n9986) );
  OAI221_X1 U12590 ( .B1(P2_REG1_REG_8__SCAN_IN), .B2(keyinput155), .C1(
        P2_D_REG_28__SCAN_IN), .C2(keyinput201), .A(n9986), .ZN(n9987) );
  NOR4_X1 U12591 ( .A1(n9990), .A2(n9989), .A3(n9988), .A4(n9987), .ZN(n10018)
         );
  AOI22_X1 U12592 ( .A1(P1_REG1_REG_20__SCAN_IN), .A2(keyinput129), .B1(
        P1_REG3_REG_27__SCAN_IN), .B2(keyinput179), .ZN(n9991) );
  OAI221_X1 U12593 ( .B1(P1_REG1_REG_20__SCAN_IN), .B2(keyinput129), .C1(
        P1_REG3_REG_27__SCAN_IN), .C2(keyinput179), .A(n9991), .ZN(n9998) );
  AOI22_X1 U12594 ( .A1(P3_DATAO_REG_29__SCAN_IN), .A2(keyinput194), .B1(
        P1_REG3_REG_16__SCAN_IN), .B2(keyinput214), .ZN(n9992) );
  OAI221_X1 U12595 ( .B1(P3_DATAO_REG_29__SCAN_IN), .B2(keyinput194), .C1(
        P1_REG3_REG_16__SCAN_IN), .C2(keyinput214), .A(n9992), .ZN(n9997) );
  AOI22_X1 U12596 ( .A1(P1_DATAO_REG_0__SCAN_IN), .A2(keyinput195), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(keyinput228), .ZN(n9993) );
  OAI221_X1 U12597 ( .B1(P1_DATAO_REG_0__SCAN_IN), .B2(keyinput195), .C1(
        P2_DATAO_REG_27__SCAN_IN), .C2(keyinput228), .A(n9993), .ZN(n9996) );
  AOI22_X1 U12598 ( .A1(P3_DATAO_REG_31__SCAN_IN), .A2(keyinput212), .B1(
        P3_DATAO_REG_13__SCAN_IN), .B2(keyinput139), .ZN(n9994) );
  OAI221_X1 U12599 ( .B1(P3_DATAO_REG_31__SCAN_IN), .B2(keyinput212), .C1(
        P3_DATAO_REG_13__SCAN_IN), .C2(keyinput139), .A(n9994), .ZN(n9995) );
  NOR4_X1 U12600 ( .A1(n9998), .A2(n9997), .A3(n9996), .A4(n9995), .ZN(n10017)
         );
  AOI22_X1 U12601 ( .A1(P3_REG1_REG_8__SCAN_IN), .A2(keyinput177), .B1(
        P3_REG2_REG_19__SCAN_IN), .B2(keyinput147), .ZN(n9999) );
  OAI221_X1 U12602 ( .B1(P3_REG1_REG_8__SCAN_IN), .B2(keyinput177), .C1(
        P3_REG2_REG_19__SCAN_IN), .C2(keyinput147), .A(n9999), .ZN(n10006) );
  AOI22_X1 U12603 ( .A1(P1_B_REG_SCAN_IN), .A2(keyinput133), .B1(SI_14_), .B2(
        keyinput160), .ZN(n10000) );
  OAI221_X1 U12604 ( .B1(P1_B_REG_SCAN_IN), .B2(keyinput133), .C1(SI_14_), 
        .C2(keyinput160), .A(n10000), .ZN(n10005) );
  AOI22_X1 U12605 ( .A1(P1_REG2_REG_8__SCAN_IN), .A2(keyinput131), .B1(
        P1_REG3_REG_4__SCAN_IN), .B2(keyinput213), .ZN(n10001) );
  OAI221_X1 U12606 ( .B1(P1_REG2_REG_8__SCAN_IN), .B2(keyinput131), .C1(
        P1_REG3_REG_4__SCAN_IN), .C2(keyinput213), .A(n10001), .ZN(n10004) );
  AOI22_X1 U12607 ( .A1(P2_REG0_REG_24__SCAN_IN), .A2(keyinput198), .B1(
        P2_REG3_REG_3__SCAN_IN), .B2(keyinput167), .ZN(n10002) );
  OAI221_X1 U12608 ( .B1(P2_REG0_REG_24__SCAN_IN), .B2(keyinput198), .C1(
        P2_REG3_REG_3__SCAN_IN), .C2(keyinput167), .A(n10002), .ZN(n10003) );
  NOR4_X1 U12609 ( .A1(n10006), .A2(n10005), .A3(n10004), .A4(n10003), .ZN(
        n10016) );
  AOI22_X1 U12610 ( .A1(P1_REG3_REG_25__SCAN_IN), .A2(keyinput233), .B1(
        P2_REG1_REG_19__SCAN_IN), .B2(keyinput132), .ZN(n10007) );
  OAI221_X1 U12611 ( .B1(P1_REG3_REG_25__SCAN_IN), .B2(keyinput233), .C1(
        P2_REG1_REG_19__SCAN_IN), .C2(keyinput132), .A(n10007), .ZN(n10014) );
  AOI22_X1 U12612 ( .A1(P2_ADDR_REG_0__SCAN_IN), .A2(keyinput221), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(keyinput244), .ZN(n10008) );
  OAI221_X1 U12613 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(keyinput221), .C1(
        P2_REG1_REG_0__SCAN_IN), .C2(keyinput244), .A(n10008), .ZN(n10013) );
  AOI22_X1 U12614 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(keyinput162), .B1(
        P2_REG0_REG_23__SCAN_IN), .B2(keyinput241), .ZN(n10009) );
  OAI221_X1 U12615 ( .B1(P1_IR_REG_12__SCAN_IN), .B2(keyinput162), .C1(
        P2_REG0_REG_23__SCAN_IN), .C2(keyinput241), .A(n10009), .ZN(n10012) );
  AOI22_X1 U12616 ( .A1(P1_REG2_REG_19__SCAN_IN), .A2(keyinput254), .B1(
        P2_REG3_REG_28__SCAN_IN), .B2(keyinput143), .ZN(n10010) );
  OAI221_X1 U12617 ( .B1(P1_REG2_REG_19__SCAN_IN), .B2(keyinput254), .C1(
        P2_REG3_REG_28__SCAN_IN), .C2(keyinput143), .A(n10010), .ZN(n10011) );
  NOR4_X1 U12618 ( .A1(n10014), .A2(n10013), .A3(n10012), .A4(n10011), .ZN(
        n10015) );
  NAND4_X1 U12619 ( .A1(n10018), .A2(n10017), .A3(n10016), .A4(n10015), .ZN(
        n10144) );
  AOI22_X1 U12620 ( .A1(P3_REG1_REG_27__SCAN_IN), .A2(keyinput157), .B1(
        P3_REG3_REG_18__SCAN_IN), .B2(keyinput206), .ZN(n10019) );
  OAI221_X1 U12621 ( .B1(P3_REG1_REG_27__SCAN_IN), .B2(keyinput157), .C1(
        P3_REG3_REG_18__SCAN_IN), .C2(keyinput206), .A(n10019), .ZN(n10026) );
  AOI22_X1 U12622 ( .A1(P3_REG1_REG_23__SCAN_IN), .A2(keyinput200), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(keyinput223), .ZN(n10020) );
  OAI221_X1 U12623 ( .B1(P3_REG1_REG_23__SCAN_IN), .B2(keyinput200), .C1(
        P2_DATAO_REG_10__SCAN_IN), .C2(keyinput223), .A(n10020), .ZN(n10025)
         );
  AOI22_X1 U12624 ( .A1(P1_REG3_REG_15__SCAN_IN), .A2(keyinput215), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(keyinput240), .ZN(n10021) );
  OAI221_X1 U12625 ( .B1(P1_REG3_REG_15__SCAN_IN), .B2(keyinput215), .C1(
        P2_DATAO_REG_17__SCAN_IN), .C2(keyinput240), .A(n10021), .ZN(n10024)
         );
  AOI22_X1 U12626 ( .A1(P1_REG0_REG_0__SCAN_IN), .A2(keyinput252), .B1(
        P1_REG2_REG_11__SCAN_IN), .B2(keyinput250), .ZN(n10022) );
  OAI221_X1 U12627 ( .B1(P1_REG0_REG_0__SCAN_IN), .B2(keyinput252), .C1(
        P1_REG2_REG_11__SCAN_IN), .C2(keyinput250), .A(n10022), .ZN(n10023) );
  NOR4_X1 U12628 ( .A1(n10026), .A2(n10025), .A3(n10024), .A4(n10023), .ZN(
        n10054) );
  AOI22_X1 U12629 ( .A1(P1_REG0_REG_23__SCAN_IN), .A2(keyinput136), .B1(
        P3_IR_REG_13__SCAN_IN), .B2(keyinput144), .ZN(n10027) );
  OAI221_X1 U12630 ( .B1(P1_REG0_REG_23__SCAN_IN), .B2(keyinput136), .C1(
        P3_IR_REG_13__SCAN_IN), .C2(keyinput144), .A(n10027), .ZN(n10034) );
  AOI22_X1 U12631 ( .A1(P2_REG0_REG_30__SCAN_IN), .A2(keyinput234), .B1(
        P2_IR_REG_24__SCAN_IN), .B2(keyinput145), .ZN(n10028) );
  OAI221_X1 U12632 ( .B1(P2_REG0_REG_30__SCAN_IN), .B2(keyinput234), .C1(
        P2_IR_REG_24__SCAN_IN), .C2(keyinput145), .A(n10028), .ZN(n10033) );
  AOI22_X1 U12633 ( .A1(P2_REG0_REG_0__SCAN_IN), .A2(keyinput203), .B1(
        P3_REG2_REG_28__SCAN_IN), .B2(keyinput154), .ZN(n10029) );
  OAI221_X1 U12634 ( .B1(P2_REG0_REG_0__SCAN_IN), .B2(keyinput203), .C1(
        P3_REG2_REG_28__SCAN_IN), .C2(keyinput154), .A(n10029), .ZN(n10032) );
  AOI22_X1 U12635 ( .A1(P1_D_REG_9__SCAN_IN), .A2(keyinput232), .B1(
        P3_D_REG_24__SCAN_IN), .B2(keyinput238), .ZN(n10030) );
  OAI221_X1 U12636 ( .B1(P1_D_REG_9__SCAN_IN), .B2(keyinput232), .C1(
        P3_D_REG_24__SCAN_IN), .C2(keyinput238), .A(n10030), .ZN(n10031) );
  NOR4_X1 U12637 ( .A1(n10034), .A2(n10033), .A3(n10032), .A4(n10031), .ZN(
        n10053) );
  AOI22_X1 U12638 ( .A1(P1_REG0_REG_30__SCAN_IN), .A2(keyinput168), .B1(
        P1_REG1_REG_14__SCAN_IN), .B2(keyinput134), .ZN(n10035) );
  OAI221_X1 U12639 ( .B1(P1_REG0_REG_30__SCAN_IN), .B2(keyinput168), .C1(
        P1_REG1_REG_14__SCAN_IN), .C2(keyinput134), .A(n10035), .ZN(n10042) );
  AOI22_X1 U12640 ( .A1(P1_D_REG_0__SCAN_IN), .A2(keyinput196), .B1(
        P3_REG2_REG_25__SCAN_IN), .B2(keyinput142), .ZN(n10036) );
  OAI221_X1 U12641 ( .B1(P1_D_REG_0__SCAN_IN), .B2(keyinput196), .C1(
        P3_REG2_REG_25__SCAN_IN), .C2(keyinput142), .A(n10036), .ZN(n10041) );
  AOI22_X1 U12642 ( .A1(P1_REG2_REG_22__SCAN_IN), .A2(keyinput243), .B1(
        P2_REG1_REG_9__SCAN_IN), .B2(keyinput181), .ZN(n10037) );
  OAI221_X1 U12643 ( .B1(P1_REG2_REG_22__SCAN_IN), .B2(keyinput243), .C1(
        P2_REG1_REG_9__SCAN_IN), .C2(keyinput181), .A(n10037), .ZN(n10040) );
  AOI22_X1 U12644 ( .A1(P1_REG2_REG_20__SCAN_IN), .A2(keyinput185), .B1(
        P2_IR_REG_11__SCAN_IN), .B2(keyinput246), .ZN(n10038) );
  OAI221_X1 U12645 ( .B1(P1_REG2_REG_20__SCAN_IN), .B2(keyinput185), .C1(
        P2_IR_REG_11__SCAN_IN), .C2(keyinput246), .A(n10038), .ZN(n10039) );
  NOR4_X1 U12646 ( .A1(n10042), .A2(n10041), .A3(n10040), .A4(n10039), .ZN(
        n10052) );
  AOI22_X1 U12647 ( .A1(P3_ADDR_REG_1__SCAN_IN), .A2(keyinput242), .B1(
        P3_REG3_REG_17__SCAN_IN), .B2(keyinput229), .ZN(n10043) );
  OAI221_X1 U12648 ( .B1(P3_ADDR_REG_1__SCAN_IN), .B2(keyinput242), .C1(
        P3_REG3_REG_17__SCAN_IN), .C2(keyinput229), .A(n10043), .ZN(n10050) );
  AOI22_X1 U12649 ( .A1(P1_REG0_REG_12__SCAN_IN), .A2(keyinput159), .B1(
        P3_D_REG_20__SCAN_IN), .B2(keyinput173), .ZN(n10044) );
  OAI221_X1 U12650 ( .B1(P1_REG0_REG_12__SCAN_IN), .B2(keyinput159), .C1(
        P3_D_REG_20__SCAN_IN), .C2(keyinput173), .A(n10044), .ZN(n10049) );
  AOI22_X1 U12651 ( .A1(P3_DATAO_REG_11__SCAN_IN), .A2(keyinput224), .B1(
        P1_REG0_REG_31__SCAN_IN), .B2(keyinput175), .ZN(n10045) );
  OAI221_X1 U12652 ( .B1(P3_DATAO_REG_11__SCAN_IN), .B2(keyinput224), .C1(
        P1_REG0_REG_31__SCAN_IN), .C2(keyinput175), .A(n10045), .ZN(n10048) );
  AOI22_X1 U12653 ( .A1(P2_D_REG_25__SCAN_IN), .A2(keyinput152), .B1(n10220), 
        .B2(keyinput149), .ZN(n10046) );
  OAI221_X1 U12654 ( .B1(P2_D_REG_25__SCAN_IN), .B2(keyinput152), .C1(n10220), 
        .C2(keyinput149), .A(n10046), .ZN(n10047) );
  NOR4_X1 U12655 ( .A1(n10050), .A2(n10049), .A3(n10048), .A4(n10047), .ZN(
        n10051) );
  NAND4_X1 U12656 ( .A1(n10054), .A2(n10053), .A3(n10052), .A4(n10051), .ZN(
        n10143) );
  INV_X1 U12657 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n15305) );
  AOI22_X1 U12658 ( .A1(n15010), .A2(keyinput161), .B1(keyinput205), .B2(
        n15305), .ZN(n10055) );
  OAI221_X1 U12659 ( .B1(n15010), .B2(keyinput161), .C1(n15305), .C2(
        keyinput205), .A(n10055), .ZN(n10063) );
  INV_X1 U12660 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n13006) );
  AOI22_X1 U12661 ( .A1(n13006), .A2(keyinput220), .B1(n10488), .B2(
        keyinput137), .ZN(n10056) );
  OAI221_X1 U12662 ( .B1(n13006), .B2(keyinput220), .C1(n10488), .C2(
        keyinput137), .A(n10056), .ZN(n10062) );
  XNOR2_X1 U12663 ( .A(P3_REG3_REG_12__SCAN_IN), .B(keyinput217), .ZN(n10060)
         );
  XNOR2_X1 U12664 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(keyinput191), .ZN(n10059)
         );
  XNOR2_X1 U12665 ( .A(P3_IR_REG_4__SCAN_IN), .B(keyinput169), .ZN(n10058) );
  XNOR2_X1 U12666 ( .A(P1_IR_REG_22__SCAN_IN), .B(keyinput148), .ZN(n10057) );
  NAND4_X1 U12667 ( .A1(n10060), .A2(n10059), .A3(n10058), .A4(n10057), .ZN(
        n10061) );
  NOR3_X1 U12668 ( .A1(n10063), .A2(n10062), .A3(n10061), .ZN(n10097) );
  AOI22_X1 U12669 ( .A1(n10158), .A2(keyinput210), .B1(n14752), .B2(
        keyinput164), .ZN(n10064) );
  OAI221_X1 U12670 ( .B1(n10158), .B2(keyinput210), .C1(n14752), .C2(
        keyinput164), .A(n10064), .ZN(n10072) );
  INV_X1 U12671 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n12317) );
  AOI22_X1 U12672 ( .A1(n11830), .A2(keyinput202), .B1(keyinput156), .B2(
        n12317), .ZN(n10065) );
  OAI221_X1 U12673 ( .B1(n11830), .B2(keyinput202), .C1(n12317), .C2(
        keyinput156), .A(n10065), .ZN(n10071) );
  INV_X1 U12674 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n10067) );
  AOI22_X1 U12675 ( .A1(n10067), .A2(keyinput204), .B1(keyinput190), .B2(
        n10572), .ZN(n10066) );
  OAI221_X1 U12676 ( .B1(n10067), .B2(keyinput204), .C1(n10572), .C2(
        keyinput190), .A(n10066), .ZN(n10070) );
  INV_X1 U12677 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n14837) );
  AOI22_X1 U12678 ( .A1(n14837), .A2(keyinput199), .B1(keyinput174), .B2(
        n10178), .ZN(n10068) );
  OAI221_X1 U12679 ( .B1(n14837), .B2(keyinput199), .C1(n10178), .C2(
        keyinput174), .A(n10068), .ZN(n10069) );
  NOR4_X1 U12680 ( .A1(n10072), .A2(n10071), .A3(n10070), .A4(n10069), .ZN(
        n10096) );
  AOI22_X1 U12681 ( .A1(n9319), .A2(keyinput189), .B1(keyinput183), .B2(n10222), .ZN(n10073) );
  OAI221_X1 U12682 ( .B1(n9319), .B2(keyinput189), .C1(n10222), .C2(
        keyinput183), .A(n10073), .ZN(n10082) );
  INV_X1 U12683 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n15289) );
  AOI22_X1 U12684 ( .A1(n13800), .A2(keyinput192), .B1(keyinput150), .B2(
        n15289), .ZN(n10074) );
  OAI221_X1 U12685 ( .B1(n13800), .B2(keyinput192), .C1(n15289), .C2(
        keyinput150), .A(n10074), .ZN(n10081) );
  INV_X1 U12686 ( .A(P1_RD_REG_SCAN_IN), .ZN(n10195) );
  AOI22_X1 U12687 ( .A1(n10195), .A2(keyinput226), .B1(keyinput170), .B2(
        n10076), .ZN(n10075) );
  OAI221_X1 U12688 ( .B1(n10195), .B2(keyinput226), .C1(n10076), .C2(
        keyinput170), .A(n10075), .ZN(n10080) );
  INV_X1 U12689 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n14746) );
  AOI22_X1 U12690 ( .A1(n14746), .A2(keyinput225), .B1(n10078), .B2(
        keyinput249), .ZN(n10077) );
  OAI221_X1 U12691 ( .B1(n14746), .B2(keyinput225), .C1(n10078), .C2(
        keyinput249), .A(n10077), .ZN(n10079) );
  NOR4_X1 U12692 ( .A1(n10082), .A2(n10081), .A3(n10080), .A4(n10079), .ZN(
        n10095) );
  INV_X1 U12693 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n10084) );
  AOI22_X1 U12694 ( .A1(n10084), .A2(keyinput247), .B1(keyinput176), .B2(
        n14353), .ZN(n10083) );
  OAI221_X1 U12695 ( .B1(n10084), .B2(keyinput247), .C1(n14353), .C2(
        keyinput176), .A(n10083), .ZN(n10093) );
  INV_X1 U12696 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n10210) );
  INV_X1 U12697 ( .A(P2_D_REG_14__SCAN_IN), .ZN(n15341) );
  AOI22_X1 U12698 ( .A1(n10210), .A2(keyinput188), .B1(keyinput253), .B2(
        n15341), .ZN(n10085) );
  OAI221_X1 U12699 ( .B1(n10210), .B2(keyinput188), .C1(n15341), .C2(
        keyinput253), .A(n10085), .ZN(n10092) );
  AOI22_X1 U12700 ( .A1(n15023), .A2(keyinput171), .B1(n13442), .B2(
        keyinput211), .ZN(n10086) );
  OAI221_X1 U12701 ( .B1(n15023), .B2(keyinput171), .C1(n13442), .C2(
        keyinput211), .A(n10086), .ZN(n10091) );
  INV_X1 U12702 ( .A(P3_WR_REG_SCAN_IN), .ZN(n10087) );
  XOR2_X1 U12703 ( .A(keyinput208), .B(n10087), .Z(n10089) );
  XNOR2_X1 U12704 ( .A(P1_IR_REG_28__SCAN_IN), .B(keyinput251), .ZN(n10088) );
  NAND2_X1 U12705 ( .A1(n10089), .A2(n10088), .ZN(n10090) );
  NOR4_X1 U12706 ( .A1(n10093), .A2(n10092), .A3(n10091), .A4(n10090), .ZN(
        n10094) );
  NAND4_X1 U12707 ( .A1(n10097), .A2(n10096), .A3(n10095), .A4(n10094), .ZN(
        n10142) );
  INV_X1 U12708 ( .A(P3_REG2_REG_22__SCAN_IN), .ZN(n10099) );
  AOI22_X1 U12709 ( .A1(n10099), .A2(keyinput163), .B1(keyinput236), .B2(n8701), .ZN(n10098) );
  OAI221_X1 U12710 ( .B1(n10099), .B2(keyinput163), .C1(n8701), .C2(
        keyinput236), .A(n10098), .ZN(n10107) );
  AOI22_X1 U12711 ( .A1(n10516), .A2(keyinput230), .B1(keyinput245), .B2(n8514), .ZN(n10100) );
  OAI221_X1 U12712 ( .B1(n10516), .B2(keyinput230), .C1(n8514), .C2(
        keyinput245), .A(n10100), .ZN(n10106) );
  AOI22_X1 U12713 ( .A1(n15062), .A2(keyinput182), .B1(n10102), .B2(
        keyinput216), .ZN(n10101) );
  OAI221_X1 U12714 ( .B1(n15062), .B2(keyinput182), .C1(n10102), .C2(
        keyinput216), .A(n10101), .ZN(n10105) );
  INV_X1 U12715 ( .A(P3_REG2_REG_24__SCAN_IN), .ZN(n10167) );
  AOI22_X1 U12716 ( .A1(n12022), .A2(keyinput227), .B1(n10167), .B2(
        keyinput235), .ZN(n10103) );
  OAI221_X1 U12717 ( .B1(n12022), .B2(keyinput227), .C1(n10167), .C2(
        keyinput235), .A(n10103), .ZN(n10104) );
  NOR4_X1 U12718 ( .A1(n10107), .A2(n10106), .A3(n10105), .A4(n10104), .ZN(
        n10140) );
  AOI22_X1 U12719 ( .A1(n10109), .A2(keyinput146), .B1(keyinput128), .B2(
        n10610), .ZN(n10108) );
  OAI221_X1 U12720 ( .B1(n10109), .B2(keyinput146), .C1(n10610), .C2(
        keyinput128), .A(n10108), .ZN(n10117) );
  INV_X1 U12721 ( .A(P1_D_REG_29__SCAN_IN), .ZN(n15106) );
  AOI22_X1 U12722 ( .A1(n8363), .A2(keyinput209), .B1(keyinput186), .B2(n15106), .ZN(n10110) );
  OAI221_X1 U12723 ( .B1(n8363), .B2(keyinput209), .C1(n15106), .C2(
        keyinput186), .A(n10110), .ZN(n10116) );
  AOI22_X1 U12724 ( .A1(n14793), .A2(keyinput166), .B1(n10214), .B2(
        keyinput255), .ZN(n10111) );
  OAI221_X1 U12725 ( .B1(n14793), .B2(keyinput166), .C1(n10214), .C2(
        keyinput255), .A(n10111), .ZN(n10115) );
  XOR2_X1 U12726 ( .A(n9198), .B(keyinput135), .Z(n10113) );
  XNOR2_X1 U12727 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(keyinput193), .ZN(n10112)
         );
  NAND2_X1 U12728 ( .A1(n10113), .A2(n10112), .ZN(n10114) );
  NOR4_X1 U12729 ( .A1(n10117), .A2(n10116), .A3(n10115), .A4(n10114), .ZN(
        n10139) );
  INV_X1 U12730 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n10235) );
  AOI22_X1 U12731 ( .A1(n10119), .A2(keyinput219), .B1(keyinput184), .B2(
        n10235), .ZN(n10118) );
  OAI221_X1 U12732 ( .B1(n10119), .B2(keyinput219), .C1(n10235), .C2(
        keyinput184), .A(n10118), .ZN(n10127) );
  AOI22_X1 U12733 ( .A1(n15041), .A2(keyinput130), .B1(n9918), .B2(keyinput158), .ZN(n10120) );
  OAI221_X1 U12734 ( .B1(n15041), .B2(keyinput130), .C1(n9918), .C2(
        keyinput158), .A(n10120), .ZN(n10126) );
  AOI22_X1 U12735 ( .A1(n10987), .A2(keyinput165), .B1(n11848), .B2(
        keyinput207), .ZN(n10121) );
  OAI221_X1 U12736 ( .B1(n10987), .B2(keyinput165), .C1(n11848), .C2(
        keyinput207), .A(n10121), .ZN(n10125) );
  XNOR2_X1 U12737 ( .A(P3_IR_REG_31__SCAN_IN), .B(keyinput172), .ZN(n10123) );
  XNOR2_X1 U12738 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(keyinput237), .ZN(n10122)
         );
  NAND2_X1 U12739 ( .A1(n10123), .A2(n10122), .ZN(n10124) );
  NOR4_X1 U12740 ( .A1(n10127), .A2(n10126), .A3(n10125), .A4(n10124), .ZN(
        n10138) );
  AOI22_X1 U12741 ( .A1(n9089), .A2(keyinput141), .B1(n8218), .B2(keyinput178), 
        .ZN(n10128) );
  OAI221_X1 U12742 ( .B1(n9089), .B2(keyinput141), .C1(n8218), .C2(keyinput178), .A(n10128), .ZN(n10136) );
  INV_X1 U12743 ( .A(P1_D_REG_8__SCAN_IN), .ZN(n15107) );
  AOI22_X1 U12744 ( .A1(n10337), .A2(keyinput239), .B1(keyinput151), .B2(
        n15107), .ZN(n10129) );
  OAI221_X1 U12745 ( .B1(n10337), .B2(keyinput239), .C1(n15107), .C2(
        keyinput151), .A(n10129), .ZN(n10135) );
  AOI22_X1 U12746 ( .A1(n11607), .A2(keyinput187), .B1(n10797), .B2(
        keyinput180), .ZN(n10130) );
  OAI221_X1 U12747 ( .B1(n11607), .B2(keyinput187), .C1(n10797), .C2(
        keyinput180), .A(n10130), .ZN(n10134) );
  XNOR2_X1 U12748 ( .A(P2_REG1_REG_22__SCAN_IN), .B(keyinput222), .ZN(n10132)
         );
  XNOR2_X1 U12749 ( .A(P2_IR_REG_18__SCAN_IN), .B(keyinput140), .ZN(n10131) );
  NAND2_X1 U12750 ( .A1(n10132), .A2(n10131), .ZN(n10133) );
  NOR4_X1 U12751 ( .A1(n10136), .A2(n10135), .A3(n10134), .A4(n10133), .ZN(
        n10137) );
  NAND4_X1 U12752 ( .A1(n10140), .A2(n10139), .A3(n10138), .A4(n10137), .ZN(
        n10141) );
  NOR4_X1 U12753 ( .A1(n10144), .A2(n10143), .A3(n10142), .A4(n10141), .ZN(
        n10247) );
  AOI22_X1 U12754 ( .A1(P1_REG1_REG_11__SCAN_IN), .A2(keyinput10), .B1(n10488), 
        .B2(keyinput9), .ZN(n10145) );
  OAI221_X1 U12755 ( .B1(P1_REG1_REG_11__SCAN_IN), .B2(keyinput10), .C1(n10488), .C2(keyinput9), .A(n10145), .ZN(n10155) );
  AOI22_X1 U12756 ( .A1(n10147), .A2(keyinput45), .B1(keyinput93), .B2(n15500), 
        .ZN(n10146) );
  OAI221_X1 U12757 ( .B1(n10147), .B2(keyinput45), .C1(n15500), .C2(keyinput93), .A(n10146), .ZN(n10154) );
  INV_X1 U12758 ( .A(P2_D_REG_28__SCAN_IN), .ZN(n15338) );
  AOI22_X1 U12759 ( .A1(n15338), .A2(keyinput73), .B1(n10149), .B2(keyinput110), .ZN(n10148) );
  OAI221_X1 U12760 ( .B1(n15338), .B2(keyinput73), .C1(n10149), .C2(
        keyinput110), .A(n10148), .ZN(n10153) );
  AOI22_X1 U12761 ( .A1(n10151), .A2(keyinput95), .B1(keyinput99), .B2(n12022), 
        .ZN(n10150) );
  OAI221_X1 U12762 ( .B1(n10151), .B2(keyinput95), .C1(n12022), .C2(keyinput99), .A(n10150), .ZN(n10152) );
  NOR4_X1 U12763 ( .A1(n10155), .A2(n10154), .A3(n10153), .A4(n10152), .ZN(
        n10193) );
  INV_X1 U12764 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n10480) );
  AOI22_X1 U12765 ( .A1(n10337), .A2(keyinput111), .B1(n10480), .B2(keyinput53), .ZN(n10156) );
  OAI221_X1 U12766 ( .B1(n10337), .B2(keyinput111), .C1(n10480), .C2(
        keyinput53), .A(n10156), .ZN(n10165) );
  AOI22_X1 U12767 ( .A1(n14837), .A2(keyinput71), .B1(n12002), .B2(keyinput109), .ZN(n10157) );
  OAI221_X1 U12768 ( .B1(n14837), .B2(keyinput71), .C1(n12002), .C2(
        keyinput109), .A(n10157), .ZN(n10164) );
  XOR2_X1 U12769 ( .A(n10158), .B(keyinput82), .Z(n10161) );
  XNOR2_X1 U12770 ( .A(P2_IR_REG_18__SCAN_IN), .B(keyinput12), .ZN(n10160) );
  XNOR2_X1 U12771 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(keyinput65), .ZN(n10159)
         );
  NAND3_X1 U12772 ( .A1(n10161), .A2(n10160), .A3(n10159), .ZN(n10163) );
  XNOR2_X1 U12773 ( .A(n15010), .B(keyinput33), .ZN(n10162) );
  NOR4_X1 U12774 ( .A1(n10165), .A2(n10164), .A3(n10163), .A4(n10162), .ZN(
        n10192) );
  INV_X1 U12775 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n11651) );
  AOI22_X1 U12776 ( .A1(n11651), .A2(keyinput103), .B1(n10167), .B2(
        keyinput107), .ZN(n10166) );
  OAI221_X1 U12777 ( .B1(n11651), .B2(keyinput103), .C1(n10167), .C2(
        keyinput107), .A(n10166), .ZN(n10176) );
  AOI22_X1 U12778 ( .A1(n15023), .A2(keyinput43), .B1(n14752), .B2(keyinput36), 
        .ZN(n10168) );
  OAI221_X1 U12779 ( .B1(n15023), .B2(keyinput43), .C1(n14752), .C2(keyinput36), .A(n10168), .ZN(n10175) );
  INV_X1 U12780 ( .A(P2_D_REG_23__SCAN_IN), .ZN(n15340) );
  INV_X1 U12781 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n10170) );
  AOI22_X1 U12782 ( .A1(n15340), .A2(keyinput120), .B1(keyinput86), .B2(n10170), .ZN(n10169) );
  OAI221_X1 U12783 ( .B1(n15340), .B2(keyinput120), .C1(n10170), .C2(
        keyinput86), .A(n10169), .ZN(n10174) );
  XNOR2_X1 U12784 ( .A(P1_IR_REG_22__SCAN_IN), .B(keyinput20), .ZN(n10172) );
  XNOR2_X1 U12785 ( .A(keyinput61), .B(P3_REG1_REG_6__SCAN_IN), .ZN(n10171) );
  NAND2_X1 U12786 ( .A1(n10172), .A2(n10171), .ZN(n10173) );
  NOR4_X1 U12787 ( .A1(n10176), .A2(n10175), .A3(n10174), .A4(n10173), .ZN(
        n10191) );
  INV_X1 U12788 ( .A(P3_DATAO_REG_29__SCAN_IN), .ZN(n11290) );
  AOI22_X1 U12789 ( .A1(n10178), .A2(keyinput46), .B1(keyinput66), .B2(n11290), 
        .ZN(n10177) );
  OAI221_X1 U12790 ( .B1(n10178), .B2(keyinput46), .C1(n11290), .C2(keyinput66), .A(n10177), .ZN(n10189) );
  INV_X1 U12791 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n10180) );
  AOI22_X1 U12792 ( .A1(n7733), .A2(keyinput124), .B1(n10180), .B2(keyinput122), .ZN(n10179) );
  OAI221_X1 U12793 ( .B1(n7733), .B2(keyinput124), .C1(n10180), .C2(
        keyinput122), .A(n10179), .ZN(n10188) );
  AOI22_X1 U12794 ( .A1(n10183), .A2(keyinput105), .B1(n10182), .B2(
        keyinput113), .ZN(n10181) );
  OAI221_X1 U12795 ( .B1(n10183), .B2(keyinput105), .C1(n10182), .C2(
        keyinput113), .A(n10181), .ZN(n10187) );
  XNOR2_X1 U12796 ( .A(P2_REG3_REG_3__SCAN_IN), .B(keyinput39), .ZN(n10185) );
  XNOR2_X1 U12797 ( .A(P2_REG0_REG_20__SCAN_IN), .B(keyinput121), .ZN(n10184)
         );
  NAND2_X1 U12798 ( .A1(n10185), .A2(n10184), .ZN(n10186) );
  NOR4_X1 U12799 ( .A1(n10189), .A2(n10188), .A3(n10187), .A4(n10186), .ZN(
        n10190) );
  NAND4_X1 U12800 ( .A1(n10193), .A2(n10192), .A3(n10191), .A4(n10190), .ZN(
        n10246) );
  AOI22_X1 U12801 ( .A1(n10195), .A2(keyinput98), .B1(keyinput3), .B2(n11230), 
        .ZN(n10194) );
  OAI221_X1 U12802 ( .B1(n10195), .B2(keyinput98), .C1(n11230), .C2(keyinput3), 
        .A(n10194), .ZN(n10205) );
  AOI22_X1 U12803 ( .A1(n10198), .A2(keyinput11), .B1(n10197), .B2(keyinput32), 
        .ZN(n10196) );
  OAI221_X1 U12804 ( .B1(n10198), .B2(keyinput11), .C1(n10197), .C2(keyinput32), .A(n10196), .ZN(n10204) );
  XNOR2_X1 U12805 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(keyinput100), .ZN(n10202)
         );
  XNOR2_X1 U12806 ( .A(P3_IR_REG_13__SCAN_IN), .B(keyinput16), .ZN(n10201) );
  XNOR2_X1 U12807 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(keyinput63), .ZN(n10200)
         );
  XNOR2_X1 U12808 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(keyinput64), .ZN(n10199)
         );
  NAND4_X1 U12809 ( .A1(n10202), .A2(n10201), .A3(n10200), .A4(n10199), .ZN(
        n10203) );
  NOR3_X1 U12810 ( .A1(n10205), .A2(n10204), .A3(n10203), .ZN(n10244) );
  INV_X1 U12811 ( .A(P2_D_REG_25__SCAN_IN), .ZN(n15339) );
  AOI22_X1 U12812 ( .A1(n15339), .A2(keyinput24), .B1(keyinput8), .B2(n10207), 
        .ZN(n10206) );
  OAI221_X1 U12813 ( .B1(n15339), .B2(keyinput24), .C1(n10207), .C2(keyinput8), 
        .A(n10206), .ZN(n10218) );
  AOI22_X1 U12814 ( .A1(n10610), .A2(keyinput0), .B1(n14317), .B2(keyinput6), 
        .ZN(n10208) );
  OAI221_X1 U12815 ( .B1(n10610), .B2(keyinput0), .C1(n14317), .C2(keyinput6), 
        .A(n10208), .ZN(n10217) );
  AOI22_X1 U12816 ( .A1(n10211), .A2(keyinput5), .B1(n10210), .B2(keyinput60), 
        .ZN(n10209) );
  OAI221_X1 U12817 ( .B1(n10211), .B2(keyinput5), .C1(n10210), .C2(keyinput60), 
        .A(n10209), .ZN(n10216) );
  INV_X1 U12818 ( .A(P3_REG2_REG_28__SCAN_IN), .ZN(n10213) );
  AOI22_X1 U12819 ( .A1(n10214), .A2(keyinput127), .B1(n10213), .B2(keyinput26), .ZN(n10212) );
  OAI221_X1 U12820 ( .B1(n10214), .B2(keyinput127), .C1(n10213), .C2(
        keyinput26), .A(n10212), .ZN(n10215) );
  NOR4_X1 U12821 ( .A1(n10218), .A2(n10217), .A3(n10216), .A4(n10215), .ZN(
        n10243) );
  AOI22_X1 U12822 ( .A1(n9198), .A2(keyinput7), .B1(n10220), .B2(keyinput21), 
        .ZN(n10219) );
  OAI221_X1 U12823 ( .B1(n9198), .B2(keyinput7), .C1(n10220), .C2(keyinput21), 
        .A(n10219), .ZN(n10229) );
  AOI22_X1 U12824 ( .A1(n10222), .A2(keyinput55), .B1(n8218), .B2(keyinput50), 
        .ZN(n10221) );
  OAI221_X1 U12825 ( .B1(n10222), .B2(keyinput55), .C1(n8218), .C2(keyinput50), 
        .A(n10221), .ZN(n10228) );
  AOI22_X1 U12826 ( .A1(n14478), .A2(keyinput115), .B1(n10572), .B2(keyinput62), .ZN(n10223) );
  OAI221_X1 U12827 ( .B1(n14478), .B2(keyinput115), .C1(n10572), .C2(
        keyinput62), .A(n10223), .ZN(n10227) );
  XNOR2_X1 U12828 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(keyinput67), .ZN(n10225)
         );
  XNOR2_X1 U12829 ( .A(P1_REG2_REG_18__SCAN_IN), .B(keyinput54), .ZN(n10224)
         );
  NAND2_X1 U12830 ( .A1(n10225), .A2(n10224), .ZN(n10226) );
  NOR4_X1 U12831 ( .A1(n10229), .A2(n10228), .A3(n10227), .A4(n10226), .ZN(
        n10242) );
  AOI22_X1 U12832 ( .A1(n10231), .A2(keyinput40), .B1(n10553), .B2(keyinput90), 
        .ZN(n10230) );
  OAI221_X1 U12833 ( .B1(n10231), .B2(keyinput40), .C1(n10553), .C2(keyinput90), .A(n10230), .ZN(n10240) );
  AOI22_X1 U12834 ( .A1(n15107), .A2(keyinput23), .B1(keyinput96), .B2(n10233), 
        .ZN(n10232) );
  OAI221_X1 U12835 ( .B1(n15107), .B2(keyinput23), .C1(n10233), .C2(keyinput96), .A(n10232), .ZN(n10239) );
  AOI22_X1 U12836 ( .A1(n10235), .A2(keyinput56), .B1(keyinput59), .B2(n11607), 
        .ZN(n10234) );
  OAI221_X1 U12837 ( .B1(n10235), .B2(keyinput56), .C1(n11607), .C2(keyinput59), .A(n10234), .ZN(n10238) );
  INV_X1 U12838 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n13955) );
  AOI22_X1 U12839 ( .A1(n13955), .A2(keyinput47), .B1(n13047), .B2(keyinput29), 
        .ZN(n10236) );
  OAI221_X1 U12840 ( .B1(n13955), .B2(keyinput47), .C1(n13047), .C2(keyinput29), .A(n10236), .ZN(n10237) );
  NOR4_X1 U12841 ( .A1(n10240), .A2(n10239), .A3(n10238), .A4(n10237), .ZN(
        n10241) );
  NAND4_X1 U12842 ( .A1(n10244), .A2(n10243), .A3(n10242), .A4(n10241), .ZN(
        n10245) );
  NOR3_X1 U12843 ( .A1(n10247), .A2(n10246), .A3(n10245), .ZN(n10285) );
  OAI22_X1 U12844 ( .A1(P3_REG1_REG_23__SCAN_IN), .A2(keyinput72), .B1(
        keyinput77), .B2(P2_ADDR_REG_13__SCAN_IN), .ZN(n10248) );
  AOI221_X1 U12845 ( .B1(P3_REG1_REG_23__SCAN_IN), .B2(keyinput72), .C1(
        P2_ADDR_REG_13__SCAN_IN), .C2(keyinput77), .A(n10248), .ZN(n10255) );
  OAI22_X1 U12846 ( .A1(P3_IR_REG_4__SCAN_IN), .A2(keyinput41), .B1(
        P2_REG2_REG_31__SCAN_IN), .B2(keyinput13), .ZN(n10249) );
  AOI221_X1 U12847 ( .B1(P3_IR_REG_4__SCAN_IN), .B2(keyinput41), .C1(
        keyinput13), .C2(P2_REG2_REG_31__SCAN_IN), .A(n10249), .ZN(n10254) );
  OAI22_X1 U12848 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(keyinput91), .B1(
        P3_DATAO_REG_31__SCAN_IN), .B2(keyinput84), .ZN(n10250) );
  AOI221_X1 U12849 ( .B1(P2_REG3_REG_19__SCAN_IN), .B2(keyinput91), .C1(
        keyinput84), .C2(P3_DATAO_REG_31__SCAN_IN), .A(n10250), .ZN(n10253) );
  OAI22_X1 U12850 ( .A1(P3_REG3_REG_12__SCAN_IN), .A2(keyinput89), .B1(
        P1_REG2_REG_12__SCAN_IN), .B2(keyinput79), .ZN(n10251) );
  AOI221_X1 U12851 ( .B1(P3_REG3_REG_12__SCAN_IN), .B2(keyinput89), .C1(
        keyinput79), .C2(P1_REG2_REG_12__SCAN_IN), .A(n10251), .ZN(n10252) );
  NAND4_X1 U12852 ( .A1(n10255), .A2(n10254), .A3(n10253), .A4(n10252), .ZN(
        n10283) );
  OAI22_X1 U12853 ( .A1(P3_D_REG_5__SCAN_IN), .A2(keyinput88), .B1(keyinput123), .B2(P1_IR_REG_28__SCAN_IN), .ZN(n10256) );
  AOI221_X1 U12854 ( .B1(P3_D_REG_5__SCAN_IN), .B2(keyinput88), .C1(
        P1_IR_REG_28__SCAN_IN), .C2(keyinput123), .A(n10256), .ZN(n10263) );
  OAI22_X1 U12855 ( .A1(P1_REG0_REG_12__SCAN_IN), .A2(keyinput31), .B1(
        P3_ADDR_REG_1__SCAN_IN), .B2(keyinput114), .ZN(n10257) );
  AOI221_X1 U12856 ( .B1(P1_REG0_REG_12__SCAN_IN), .B2(keyinput31), .C1(
        keyinput114), .C2(P3_ADDR_REG_1__SCAN_IN), .A(n10257), .ZN(n10262) );
  OAI22_X1 U12857 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(keyinput22), .B1(
        P1_REG2_REG_30__SCAN_IN), .B2(keyinput48), .ZN(n10258) );
  AOI221_X1 U12858 ( .B1(P2_REG3_REG_13__SCAN_IN), .B2(keyinput22), .C1(
        keyinput48), .C2(P1_REG2_REG_30__SCAN_IN), .A(n10258), .ZN(n10261) );
  OAI22_X1 U12859 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(keyinput44), .B1(
        P1_DATAO_REG_31__SCAN_IN), .B2(keyinput28), .ZN(n10259) );
  AOI221_X1 U12860 ( .B1(P3_IR_REG_31__SCAN_IN), .B2(keyinput44), .C1(
        keyinput28), .C2(P1_DATAO_REG_31__SCAN_IN), .A(n10259), .ZN(n10260) );
  NAND4_X1 U12861 ( .A1(n10263), .A2(n10262), .A3(n10261), .A4(n10260), .ZN(
        n10282) );
  OAI22_X1 U12862 ( .A1(P2_REG0_REG_30__SCAN_IN), .A2(keyinput106), .B1(
        P1_D_REG_9__SCAN_IN), .B2(keyinput104), .ZN(n10264) );
  AOI221_X1 U12863 ( .B1(P2_REG0_REG_30__SCAN_IN), .B2(keyinput106), .C1(
        keyinput104), .C2(P1_D_REG_9__SCAN_IN), .A(n10264), .ZN(n10271) );
  OAI22_X1 U12864 ( .A1(P2_IR_REG_30__SCAN_IN), .A2(keyinput81), .B1(keyinput2), .B2(P1_ADDR_REG_16__SCAN_IN), .ZN(n10265) );
  AOI221_X1 U12865 ( .B1(P2_IR_REG_30__SCAN_IN), .B2(keyinput81), .C1(
        P1_ADDR_REG_16__SCAN_IN), .C2(keyinput2), .A(n10265), .ZN(n10270) );
  OAI22_X1 U12866 ( .A1(P3_REG3_REG_18__SCAN_IN), .A2(keyinput78), .B1(
        P1_REG0_REG_19__SCAN_IN), .B2(keyinput97), .ZN(n10266) );
  AOI221_X1 U12867 ( .B1(P3_REG3_REG_18__SCAN_IN), .B2(keyinput78), .C1(
        keyinput97), .C2(P1_REG0_REG_19__SCAN_IN), .A(n10266), .ZN(n10269) );
  OAI22_X1 U12868 ( .A1(P2_IR_REG_24__SCAN_IN), .A2(keyinput17), .B1(
        keyinput87), .B2(P1_REG3_REG_15__SCAN_IN), .ZN(n10267) );
  AOI221_X1 U12869 ( .B1(P2_IR_REG_24__SCAN_IN), .B2(keyinput17), .C1(
        P1_REG3_REG_15__SCAN_IN), .C2(keyinput87), .A(n10267), .ZN(n10268) );
  NAND4_X1 U12870 ( .A1(n10271), .A2(n10270), .A3(n10269), .A4(n10268), .ZN(
        n10281) );
  OAI22_X1 U12871 ( .A1(P2_REG0_REG_0__SCAN_IN), .A2(keyinput75), .B1(
        keyinput85), .B2(P1_REG3_REG_4__SCAN_IN), .ZN(n10272) );
  AOI221_X1 U12872 ( .B1(P2_REG0_REG_0__SCAN_IN), .B2(keyinput75), .C1(
        P1_REG3_REG_4__SCAN_IN), .C2(keyinput85), .A(n10272), .ZN(n10279) );
  OAI22_X1 U12873 ( .A1(P2_REG2_REG_24__SCAN_IN), .A2(keyinput108), .B1(
        keyinput58), .B2(P1_D_REG_29__SCAN_IN), .ZN(n10273) );
  AOI221_X1 U12874 ( .B1(P2_REG2_REG_24__SCAN_IN), .B2(keyinput108), .C1(
        P1_D_REG_29__SCAN_IN), .C2(keyinput58), .A(n10273), .ZN(n10278) );
  OAI22_X1 U12875 ( .A1(P1_REG0_REG_2__SCAN_IN), .A2(keyinput25), .B1(
        P2_ADDR_REG_8__SCAN_IN), .B2(keyinput38), .ZN(n10274) );
  AOI221_X1 U12876 ( .B1(P1_REG0_REG_2__SCAN_IN), .B2(keyinput25), .C1(
        keyinput38), .C2(P2_ADDR_REG_8__SCAN_IN), .A(n10274), .ZN(n10277) );
  OAI22_X1 U12877 ( .A1(P3_REG1_REG_2__SCAN_IN), .A2(keyinput102), .B1(
        P3_REG2_REG_22__SCAN_IN), .B2(keyinput35), .ZN(n10275) );
  AOI221_X1 U12878 ( .B1(P3_REG1_REG_2__SCAN_IN), .B2(keyinput102), .C1(
        keyinput35), .C2(P3_REG2_REG_22__SCAN_IN), .A(n10275), .ZN(n10276) );
  NAND4_X1 U12879 ( .A1(n10279), .A2(n10278), .A3(n10277), .A4(n10276), .ZN(
        n10280) );
  NOR4_X1 U12880 ( .A1(n10283), .A2(n10282), .A3(n10281), .A4(n10280), .ZN(
        n10284) );
  NAND3_X1 U12881 ( .A1(n10286), .A2(n10285), .A3(n10284), .ZN(n10287) );
  XNOR2_X1 U12882 ( .A(n10288), .B(n10287), .ZN(P3_U3499) );
  INV_X1 U12883 ( .A(n10289), .ZN(n10372) );
  INV_X1 U12884 ( .A(n14774), .ZN(n11286) );
  AOI22_X1 U12885 ( .A1(n11276), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n11286), .ZN(n10290) );
  OAI21_X1 U12886 ( .B1(n10372), .B2(n14761), .A(n10290), .ZN(P1_U3344) );
  INV_X1 U12887 ( .A(n10630), .ZN(n10295) );
  INV_X1 U12888 ( .A(n10291), .ZN(n10636) );
  NAND2_X1 U12889 ( .A1(n10636), .A2(n10630), .ZN(n10293) );
  NAND2_X1 U12890 ( .A1(n10293), .A2(n10292), .ZN(n10294) );
  OAI21_X1 U12891 ( .B1(n10631), .B2(n10295), .A(n10294), .ZN(n15236) );
  OR2_X1 U12892 ( .A1(n15236), .A2(P2_U3088), .ZN(n15306) );
  INV_X1 U12893 ( .A(n15306), .ZN(n15313) );
  AND2_X1 U12894 ( .A1(n8867), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10296) );
  NAND2_X1 U12895 ( .A1(P2_U3088), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n10929) );
  INV_X1 U12896 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n10297) );
  MUX2_X1 U12897 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n10297), .S(n10344), .Z(
        n10309) );
  INV_X1 U12898 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n15384) );
  MUX2_X1 U12899 ( .A(n15384), .B(P2_REG1_REG_2__SCAN_IN), .S(n15223), .Z(
        n15221) );
  INV_X1 U12900 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n10590) );
  MUX2_X1 U12901 ( .A(n10590), .B(P2_REG1_REG_1__SCAN_IN), .S(n10313), .Z(
        n15203) );
  NAND2_X1 U12902 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n15204) );
  INV_X1 U12903 ( .A(n15204), .ZN(n10298) );
  NAND2_X1 U12904 ( .A1(n15203), .A2(n10298), .ZN(n15207) );
  NAND2_X1 U12905 ( .A1(n15208), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n10299) );
  NAND2_X1 U12906 ( .A1(n15207), .A2(n10299), .ZN(n15220) );
  NAND2_X1 U12907 ( .A1(n15221), .A2(n15220), .ZN(n15219) );
  OR2_X1 U12908 ( .A1(n15223), .A2(n15384), .ZN(n10300) );
  NAND2_X1 U12909 ( .A1(n15219), .A2(n10300), .ZN(n15233) );
  INV_X1 U12910 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n10601) );
  MUX2_X1 U12911 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n10601), .S(n10315), .Z(
        n15234) );
  NAND2_X1 U12912 ( .A1(n15233), .A2(n15234), .ZN(n15232) );
  NAND2_X1 U12913 ( .A1(n10315), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n10301) );
  NAND2_X1 U12914 ( .A1(n15232), .A2(n10301), .ZN(n10326) );
  INV_X1 U12915 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n10772) );
  MUX2_X1 U12916 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n10772), .S(n10316), .Z(
        n10327) );
  NAND2_X1 U12917 ( .A1(n10326), .A2(n10327), .ZN(n10325) );
  NAND2_X1 U12918 ( .A1(n10316), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n10302) );
  NAND2_X1 U12919 ( .A1(n10325), .A2(n10302), .ZN(n10355) );
  INV_X1 U12920 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n10303) );
  MUX2_X1 U12921 ( .A(n10303), .B(P2_REG1_REG_5__SCAN_IN), .S(n10359), .Z(
        n10356) );
  NAND2_X1 U12922 ( .A1(n10355), .A2(n10356), .ZN(n10354) );
  NAND2_X1 U12923 ( .A1(n10318), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n10304) );
  NAND2_X1 U12924 ( .A1(n10354), .A2(n10304), .ZN(n10308) );
  NAND2_X1 U12925 ( .A1(n10305), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13794) );
  INV_X1 U12926 ( .A(n8868), .ZN(n10306) );
  NOR2_X1 U12927 ( .A1(n13794), .A2(n10306), .ZN(n10307) );
  NAND2_X1 U12928 ( .A1(n10308), .A2(n10309), .ZN(n10346) );
  OAI211_X1 U12929 ( .C1(n10309), .C2(n10308), .A(n15307), .B(n10346), .ZN(
        n10310) );
  OAI211_X1 U12930 ( .C1(n15224), .C2(n10336), .A(n10929), .B(n10310), .ZN(
        n10323) );
  NOR2_X1 U12931 ( .A1(n13794), .A2(n8868), .ZN(n10311) );
  AND2_X1 U12932 ( .A1(n15236), .A2(n10311), .ZN(n15314) );
  MUX2_X1 U12933 ( .A(n10312), .B(P2_REG2_REG_1__SCAN_IN), .S(n10313), .Z(
        n15214) );
  NAND3_X1 U12934 ( .A1(n15214), .A2(P2_IR_REG_0__SCAN_IN), .A3(
        P2_REG2_REG_0__SCAN_IN), .ZN(n15213) );
  OAI21_X1 U12935 ( .B1(n10312), .B2(n10313), .A(n15213), .ZN(n15228) );
  MUX2_X1 U12936 ( .A(n13663), .B(P2_REG2_REG_2__SCAN_IN), .S(n15223), .Z(
        n15227) );
  NAND2_X1 U12937 ( .A1(n15228), .A2(n15227), .ZN(n15226) );
  OAI21_X1 U12938 ( .B1(n13663), .B2(n15223), .A(n15226), .ZN(n15242) );
  MUX2_X1 U12939 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n10314), .S(n10315), .Z(
        n15241) );
  NAND2_X1 U12940 ( .A1(n15242), .A2(n15241), .ZN(n15240) );
  NAND2_X1 U12941 ( .A1(n10315), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n10331) );
  MUX2_X1 U12942 ( .A(n11133), .B(P2_REG2_REG_4__SCAN_IN), .S(n10316), .Z(
        n10330) );
  AOI21_X1 U12943 ( .B1(n15240), .B2(n10331), .A(n10330), .ZN(n10363) );
  NOR2_X1 U12944 ( .A1(n10329), .A2(n11133), .ZN(n10362) );
  MUX2_X1 U12945 ( .A(n10317), .B(P2_REG2_REG_5__SCAN_IN), .S(n10359), .Z(
        n10361) );
  OAI21_X1 U12946 ( .B1(n10363), .B2(n10362), .A(n10361), .ZN(n10360) );
  NAND2_X1 U12947 ( .A1(n10318), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n10320) );
  MUX2_X1 U12948 ( .A(n11141), .B(P2_REG2_REG_6__SCAN_IN), .S(n10344), .Z(
        n10319) );
  AOI21_X1 U12949 ( .B1(n10360), .B2(n10320), .A(n10319), .ZN(n13388) );
  AND3_X1 U12950 ( .A1(n10360), .A2(n10320), .A3(n10319), .ZN(n10321) );
  NOR3_X1 U12951 ( .A1(n15298), .A2(n13388), .A3(n10321), .ZN(n10322) );
  AOI211_X1 U12952 ( .C1(P2_ADDR_REG_6__SCAN_IN), .C2(n15313), .A(n10323), .B(
        n10322), .ZN(n10324) );
  INV_X1 U12953 ( .A(n10324), .ZN(P2_U3220) );
  NAND2_X1 U12954 ( .A1(P2_U3088), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n10840) );
  OAI211_X1 U12955 ( .C1(n10327), .C2(n10326), .A(n15307), .B(n10325), .ZN(
        n10328) );
  OAI211_X1 U12956 ( .C1(n15224), .C2(n10329), .A(n10840), .B(n10328), .ZN(
        n10334) );
  AND3_X1 U12957 ( .A1(n15240), .A2(n10331), .A3(n10330), .ZN(n10332) );
  NOR3_X1 U12958 ( .A1(n15298), .A2(n10363), .A3(n10332), .ZN(n10333) );
  AOI211_X1 U12959 ( .C1(P2_ADDR_REG_4__SCAN_IN), .C2(n15313), .A(n10334), .B(
        n10333), .ZN(n10335) );
  INV_X1 U12960 ( .A(n10335), .ZN(P2_U3218) );
  NOR2_X1 U12961 ( .A1(n10336), .A2(n11141), .ZN(n13387) );
  MUX2_X1 U12962 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n10337), .S(n13392), .Z(
        n13386) );
  OAI21_X1 U12963 ( .B1(n13388), .B2(n13387), .A(n13386), .ZN(n13385) );
  NAND2_X1 U12964 ( .A1(n13392), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n10339) );
  MUX2_X1 U12965 ( .A(n11461), .B(P2_REG2_REG_8__SCAN_IN), .S(n10477), .Z(
        n10338) );
  AOI21_X1 U12966 ( .B1(n13385), .B2(n10339), .A(n10338), .ZN(n10470) );
  NAND3_X1 U12967 ( .A1(n13385), .A2(n10339), .A3(n10338), .ZN(n10340) );
  NAND2_X1 U12968 ( .A1(n15314), .A2(n10340), .ZN(n10353) );
  NAND2_X1 U12969 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3088), .ZN(n11352) );
  INV_X1 U12970 ( .A(n11352), .ZN(n10343) );
  NOR2_X1 U12971 ( .A1(n15224), .A2(n10341), .ZN(n10342) );
  AOI211_X1 U12972 ( .C1(n15313), .C2(P2_ADDR_REG_8__SCAN_IN), .A(n10343), .B(
        n10342), .ZN(n10352) );
  INV_X1 U12973 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n15386) );
  MUX2_X1 U12974 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n15386), .S(n10477), .Z(
        n10350) );
  NAND2_X1 U12975 ( .A1(n10344), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n10345) );
  NAND2_X1 U12976 ( .A1(n10346), .A2(n10345), .ZN(n13395) );
  INV_X1 U12977 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n10347) );
  MUX2_X1 U12978 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n10347), .S(n13392), .Z(
        n13396) );
  NAND2_X1 U12979 ( .A1(n13395), .A2(n13396), .ZN(n13394) );
  NAND2_X1 U12980 ( .A1(n13392), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n10348) );
  NAND2_X1 U12981 ( .A1(n13394), .A2(n10348), .ZN(n10349) );
  NAND2_X1 U12982 ( .A1(n10349), .A2(n10350), .ZN(n10479) );
  OAI211_X1 U12983 ( .C1(n10350), .C2(n10349), .A(n15307), .B(n10479), .ZN(
        n10351) );
  OAI211_X1 U12984 ( .C1(n10470), .C2(n10353), .A(n10352), .B(n10351), .ZN(
        P2_U3222) );
  AND2_X1 U12985 ( .A1(P2_U3088), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n10879) );
  INV_X1 U12986 ( .A(n10879), .ZN(n10358) );
  OAI211_X1 U12987 ( .C1(n10356), .C2(n10355), .A(n15307), .B(n10354), .ZN(
        n10357) );
  OAI211_X1 U12988 ( .C1(n15224), .C2(n10359), .A(n10358), .B(n10357), .ZN(
        n10367) );
  INV_X1 U12989 ( .A(n10360), .ZN(n10365) );
  NOR3_X1 U12990 ( .A1(n10363), .A2(n10362), .A3(n10361), .ZN(n10364) );
  NOR3_X1 U12991 ( .A1(n15298), .A2(n10365), .A3(n10364), .ZN(n10366) );
  AOI211_X1 U12992 ( .C1(P2_ADDR_REG_5__SCAN_IN), .C2(n15313), .A(n10367), .B(
        n10366), .ZN(n10368) );
  INV_X1 U12993 ( .A(n10368), .ZN(P2_U3219) );
  INV_X1 U12994 ( .A(n10369), .ZN(n10370) );
  OAI222_X1 U12995 ( .A1(n13167), .A2(n10371), .B1(n13172), .B2(n10370), .C1(
        n12784), .C2(P3_U3151), .ZN(P3_U3280) );
  INV_X1 U12996 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n10373) );
  INV_X1 U12997 ( .A(n11491), .ZN(n11505) );
  OAI222_X1 U12998 ( .A1(n13798), .A2(n10373), .B1(n13804), .B2(n10372), .C1(
        P2_U3088), .C2(n11505), .ZN(P2_U3316) );
  NAND2_X1 U12999 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3086), .ZN(n11551) );
  OAI21_X1 U13000 ( .B1(n15070), .B2(n10374), .A(n11551), .ZN(n10381) );
  MUX2_X1 U13001 ( .A(n10377), .B(P1_REG1_REG_7__SCAN_IN), .S(n10989), .Z(
        n10378) );
  NOR2_X1 U13002 ( .A1(n10379), .A2(n10378), .ZN(n10988) );
  AOI211_X1 U13003 ( .C1(n10379), .C2(n10378), .A(n15056), .B(n10988), .ZN(
        n10380) );
  AOI211_X1 U13004 ( .C1(n15067), .C2(n10989), .A(n10381), .B(n10380), .ZN(
        n10388) );
  OAI21_X1 U13005 ( .B1(n10384), .B2(n10383), .A(n10382), .ZN(n10386) );
  MUX2_X1 U13006 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n11162), .S(n10989), .Z(
        n10385) );
  NAND2_X1 U13007 ( .A1(n10386), .A2(n10385), .ZN(n10982) );
  OAI211_X1 U13008 ( .C1(n10386), .C2(n10385), .A(n10982), .B(n15012), .ZN(
        n10387) );
  NAND2_X1 U13009 ( .A1(n10388), .A2(n10387), .ZN(P1_U3250) );
  INV_X1 U13010 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n10393) );
  OR2_X2 U13011 ( .A1(n10390), .A2(n10395), .ZN(n10429) );
  NAND2_X1 U13012 ( .A1(n14233), .A2(n10428), .ZN(n10391) );
  OAI211_X1 U13013 ( .C1(n10394), .C2(n10393), .A(n10392), .B(n10391), .ZN(
        n10400) );
  INV_X1 U13014 ( .A(n10400), .ZN(n10427) );
  AND2_X4 U13015 ( .A1(n6628), .A2(n14915), .ZN(n12301) );
  AND2_X1 U13016 ( .A1(n10395), .A2(P1_IR_REG_0__SCAN_IN), .ZN(n10396) );
  INV_X1 U13017 ( .A(n10399), .ZN(n10401) );
  AOI21_X1 U13018 ( .B1(n10427), .B2(n10401), .A(n10426), .ZN(n10439) );
  INV_X1 U13019 ( .A(n10402), .ZN(n10403) );
  OR3_X1 U13020 ( .A1(n10405), .A2(n10404), .A3(n10403), .ZN(n10418) );
  NOR2_X1 U13021 ( .A1(n10418), .A2(n10406), .ZN(n10410) );
  NOR2_X1 U13022 ( .A1(n15155), .A2(n10407), .ZN(n10408) );
  NAND2_X1 U13023 ( .A1(n10410), .A2(n10409), .ZN(n10411) );
  NAND2_X1 U13024 ( .A1(n10418), .A2(n10412), .ZN(n10416) );
  AND2_X1 U13025 ( .A1(n10414), .A2(n10413), .ZN(n10415) );
  NAND2_X1 U13026 ( .A1(n10416), .A2(n10415), .ZN(n11190) );
  OR2_X1 U13027 ( .A1(n11190), .A2(P1_U3086), .ZN(n10500) );
  AOI22_X1 U13028 ( .A1(n14909), .A2(n10417), .B1(P1_REG3_REG_0__SCAN_IN), 
        .B2(n10500), .ZN(n10422) );
  INV_X1 U13029 ( .A(n10418), .ZN(n10420) );
  NAND2_X1 U13030 ( .A1(n10420), .A2(n10419), .ZN(n13916) );
  NAND2_X1 U13031 ( .A1(n13934), .A2(n15095), .ZN(n10421) );
  OAI211_X1 U13032 ( .C1(n10439), .C2(n14904), .A(n10422), .B(n10421), .ZN(
        P1_U3232) );
  INV_X1 U13033 ( .A(n10423), .ZN(n10424) );
  OAI222_X1 U13034 ( .A1(n13167), .A2(n10425), .B1(n13172), .B2(n10424), .C1(
        n12802), .C2(P3_U3151), .ZN(P3_U3279) );
  XNOR2_X1 U13035 ( .A(n10431), .B(n10430), .ZN(n10433) );
  AOI22_X1 U13036 ( .A1(n12301), .A2(n14231), .B1(n10428), .B2(n13969), .ZN(
        n10432) );
  OAI21_X1 U13037 ( .B1(n10433), .B2(n10432), .A(n10494), .ZN(n10435) );
  NOR2_X1 U13038 ( .A1(n10434), .A2(n10435), .ZN(n10496) );
  AOI21_X1 U13039 ( .B1(n10434), .B2(n10435), .A(n10496), .ZN(n10438) );
  NAND2_X1 U13040 ( .A1(n13934), .A2(n14583), .ZN(n14897) );
  INV_X1 U13041 ( .A(n14897), .ZN(n13827) );
  NOR2_X2 U13042 ( .A1(n13916), .A2(n14601), .ZN(n13943) );
  AOI22_X1 U13043 ( .A1(n13827), .A2(n14230), .B1(n13943), .B2(n14233), .ZN(
        n10437) );
  AOI22_X1 U13044 ( .A1(n14909), .A2(n13969), .B1(P1_REG3_REG_1__SCAN_IN), 
        .B2(n10500), .ZN(n10436) );
  OAI211_X1 U13045 ( .C1(n10438), .C2(n14904), .A(n10437), .B(n10436), .ZN(
        P1_U3222) );
  MUX2_X1 U13046 ( .A(n14235), .B(n10439), .S(n6625), .Z(n10442) );
  AOI21_X1 U13047 ( .B1(n14978), .B2(n7731), .A(n12173), .ZN(n14977) );
  OAI21_X1 U13048 ( .B1(P1_IR_REG_0__SCAN_IN), .B2(n14977), .A(n14232), .ZN(
        n10440) );
  AOI21_X1 U13049 ( .B1(n10442), .B2(n10441), .A(n10440), .ZN(n10469) );
  INV_X1 U13050 ( .A(n15056), .ZN(n15015) );
  OAI211_X1 U13051 ( .C1(n10445), .C2(n10444), .A(n15015), .B(n10443), .ZN(
        n10453) );
  OAI211_X1 U13052 ( .C1(n10448), .C2(n10447), .A(n15012), .B(n10446), .ZN(
        n10452) );
  AOI22_X1 U13053 ( .A1(n14981), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n10451) );
  NAND2_X1 U13054 ( .A1(n15067), .A2(n10449), .ZN(n10450) );
  NAND4_X1 U13055 ( .A1(n10453), .A2(n10452), .A3(n10451), .A4(n10450), .ZN(
        n10454) );
  OR2_X1 U13056 ( .A1(n10469), .A2(n10454), .ZN(P1_U3245) );
  INV_X1 U13057 ( .A(n10455), .ZN(n10489) );
  AOI22_X1 U13058 ( .A1(n14319), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n11286), .ZN(n10456) );
  OAI21_X1 U13059 ( .B1(n10489), .B2(n14761), .A(n10456), .ZN(P1_U3343) );
  AOI211_X1 U13060 ( .C1(n10459), .C2(n10458), .A(n15056), .B(n10457), .ZN(
        n10468) );
  INV_X1 U13061 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n10460) );
  NAND2_X1 U13062 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_U3086), .ZN(n11212) );
  OAI21_X1 U13063 ( .B1(n15070), .B2(n10460), .A(n11212), .ZN(n10467) );
  OAI211_X1 U13064 ( .C1(n10463), .C2(n10462), .A(n15012), .B(n10461), .ZN(
        n10464) );
  OAI21_X1 U13065 ( .B1(n15037), .B2(n10465), .A(n10464), .ZN(n10466) );
  OR4_X1 U13066 ( .A1(n10469), .A2(n10468), .A3(n10467), .A4(n10466), .ZN(
        P1_U3247) );
  AOI21_X1 U13067 ( .B1(n10477), .B2(P2_REG2_REG_8__SCAN_IN), .A(n10470), .ZN(
        n15247) );
  INV_X1 U13068 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n10471) );
  MUX2_X1 U13069 ( .A(P2_REG2_REG_9__SCAN_IN), .B(n10471), .S(n15253), .Z(
        n15246) );
  NAND2_X1 U13070 ( .A1(n15247), .A2(n15246), .ZN(n15245) );
  OAI21_X1 U13071 ( .B1(P2_REG2_REG_9__SCAN_IN), .B2(n15253), .A(n15245), .ZN(
        n15266) );
  MUX2_X1 U13072 ( .A(n8514), .B(P2_REG2_REG_10__SCAN_IN), .S(n15264), .Z(
        n15267) );
  NOR2_X1 U13073 ( .A1(n15266), .A2(n15267), .ZN(n15265) );
  AOI21_X1 U13074 ( .B1(n15264), .B2(P2_REG2_REG_10__SCAN_IN), .A(n15265), 
        .ZN(n10473) );
  MUX2_X1 U13075 ( .A(P2_REG2_REG_11__SCAN_IN), .B(n11758), .S(n11491), .Z(
        n10472) );
  AND2_X1 U13076 ( .A1(n10473), .A2(n10472), .ZN(n11506) );
  INV_X1 U13077 ( .A(n11506), .ZN(n15280) );
  OAI21_X1 U13078 ( .B1(n10473), .B2(n10472), .A(n15280), .ZN(n10476) );
  AND2_X1 U13079 ( .A1(P2_U3088), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n11781) );
  AOI21_X1 U13080 ( .B1(n15313), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n11781), 
        .ZN(n10474) );
  OAI21_X1 U13081 ( .B1(n11505), .B2(n15224), .A(n10474), .ZN(n10475) );
  AOI21_X1 U13082 ( .B1(n10476), .B2(n15314), .A(n10475), .ZN(n10487) );
  NAND2_X1 U13083 ( .A1(n10477), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n10478) );
  NAND2_X1 U13084 ( .A1(n10479), .A2(n10478), .ZN(n15249) );
  MUX2_X1 U13085 ( .A(n10480), .B(P2_REG1_REG_9__SCAN_IN), .S(n15253), .Z(
        n15248) );
  OR2_X1 U13086 ( .A1(n15249), .A2(n15248), .ZN(n15251) );
  OR2_X1 U13087 ( .A1(n15253), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n10481) );
  NAND2_X1 U13088 ( .A1(n15251), .A2(n10481), .ZN(n15260) );
  INV_X1 U13089 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n10482) );
  MUX2_X1 U13090 ( .A(n10482), .B(P2_REG1_REG_10__SCAN_IN), .S(n15264), .Z(
        n15261) );
  OR2_X1 U13091 ( .A1(n15260), .A2(n15261), .ZN(n15258) );
  NAND2_X1 U13092 ( .A1(n15264), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n10483) );
  NAND2_X1 U13093 ( .A1(n15258), .A2(n10483), .ZN(n10485) );
  INV_X1 U13094 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n15390) );
  MUX2_X1 U13095 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n15390), .S(n11491), .Z(
        n10484) );
  NAND2_X1 U13096 ( .A1(n10485), .A2(n10484), .ZN(n11493) );
  OAI211_X1 U13097 ( .C1(n10485), .C2(n10484), .A(n11493), .B(n15307), .ZN(
        n10486) );
  NAND2_X1 U13098 ( .A1(n10487), .A2(n10486), .ZN(P2_U3225) );
  INV_X1 U13099 ( .A(n15285), .ZN(n11494) );
  OAI222_X1 U13100 ( .A1(n13804), .A2(n10489), .B1(n11494), .B2(P2_U3088), 
        .C1(n10488), .C2(n13798), .ZN(P2_U3315) );
  OAI22_X1 U13101 ( .A1(n13172), .A2(n10490), .B1(SI_17_), .B2(n13167), .ZN(
        n10491) );
  AOI21_X1 U13102 ( .B1(n12817), .B2(P3_STATE_REG_SCAN_IN), .A(n10491), .ZN(
        P3_U3278) );
  INV_X1 U13103 ( .A(n10492), .ZN(n10552) );
  INV_X1 U13104 ( .A(n15297), .ZN(n10493) );
  OAI222_X1 U13105 ( .A1(n13804), .A2(n10552), .B1(n10493), .B2(P2_U3088), 
        .C1(n7174), .C2(n13798), .ZN(P2_U3314) );
  INV_X1 U13106 ( .A(n10494), .ZN(n10495) );
  OAI22_X1 U13107 ( .A1(n13976), .A2(n11299), .B1(n10429), .B2(n15111), .ZN(
        n10497) );
  XNOR2_X1 U13108 ( .A(n10497), .B(n12208), .ZN(n11171) );
  INV_X2 U13109 ( .A(n12301), .ZN(n12284) );
  OAI22_X1 U13110 ( .A1(n12284), .A2(n13976), .B1(n15111), .B2(n11299), .ZN(
        n11170) );
  XNOR2_X1 U13111 ( .A(n11171), .B(n11170), .ZN(n10498) );
  AOI21_X1 U13112 ( .B1(n10499), .B2(n10498), .A(n11172), .ZN(n10503) );
  AOI22_X1 U13113 ( .A1(n13827), .A2(n14229), .B1(n13943), .B2(n14231), .ZN(
        n10502) );
  AOI22_X1 U13114 ( .A1(n14909), .A2(n13978), .B1(P1_REG3_REG_2__SCAN_IN), 
        .B2(n10500), .ZN(n10501) );
  OAI211_X1 U13115 ( .C1(n10503), .C2(n14904), .A(n10502), .B(n10501), .ZN(
        P1_U3237) );
  INV_X1 U13116 ( .A(n10702), .ZN(n10504) );
  OR2_X1 U13117 ( .A1(n10670), .A2(P3_U3151), .ZN(n12725) );
  NAND2_X1 U13118 ( .A1(n10504), .A2(n12725), .ZN(n10537) );
  NAND2_X1 U13119 ( .A1(n12647), .A2(n10670), .ZN(n10505) );
  NAND2_X1 U13120 ( .A1(n10506), .A2(n10505), .ZN(n10536) );
  INV_X1 U13121 ( .A(n10536), .ZN(n10507) );
  NAND2_X1 U13122 ( .A1(n10537), .A2(n10507), .ZN(n10535) );
  INV_X1 U13123 ( .A(n10535), .ZN(n10508) );
  MUX2_X1 U13124 ( .A(P3_U3897), .B(n10508), .S(n13162), .Z(n15417) );
  INV_X1 U13125 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n10510) );
  INV_X1 U13126 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n10509) );
  MUX2_X1 U13127 ( .A(n10510), .B(n10509), .S(n9689), .Z(n10512) );
  INV_X1 U13128 ( .A(n10511), .ZN(n10949) );
  NAND2_X1 U13129 ( .A1(n10512), .A2(n10949), .ZN(n10515) );
  OAI21_X1 U13130 ( .B1(n10512), .B2(n10949), .A(n10515), .ZN(n10936) );
  INV_X1 U13131 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n10514) );
  MUX2_X1 U13132 ( .A(n10514), .B(n10513), .S(n9689), .Z(n10614) );
  NAND2_X1 U13133 ( .A1(n10614), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n10937) );
  INV_X1 U13134 ( .A(n10515), .ZN(n10579) );
  INV_X1 U13135 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n10532) );
  MUX2_X1 U13136 ( .A(n10532), .B(n10516), .S(n9689), .Z(n10517) );
  NAND2_X1 U13137 ( .A1(n10517), .A2(n10533), .ZN(n10524) );
  INV_X1 U13138 ( .A(n10517), .ZN(n10518) );
  NAND2_X1 U13139 ( .A1(n10518), .A2(n10584), .ZN(n10519) );
  OAI21_X1 U13140 ( .B1(n10935), .B2(n10579), .A(n10578), .ZN(n10577) );
  INV_X1 U13141 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n11476) );
  INV_X1 U13142 ( .A(n10520), .ZN(n10521) );
  NAND2_X1 U13143 ( .A1(n10521), .A2(n10805), .ZN(n10522) );
  NAND2_X1 U13144 ( .A1(n10788), .A2(n10522), .ZN(n10523) );
  AND3_X1 U13145 ( .A1(n10577), .A2(n10524), .A3(n10523), .ZN(n10525) );
  NAND2_X1 U13146 ( .A1(P3_U3897), .A2(n13162), .ZN(n15406) );
  INV_X1 U13147 ( .A(n15406), .ZN(n15430) );
  OAI21_X1 U13148 ( .B1(n10790), .B2(n10525), .A(n15430), .ZN(n10543) );
  NAND2_X1 U13149 ( .A1(P3_REG1_REG_0__SCAN_IN), .A2(n10529), .ZN(n10527) );
  INV_X1 U13150 ( .A(n10527), .ZN(n10613) );
  NOR2_X1 U13151 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(n10527), .ZN(n10526) );
  AOI21_X1 U13152 ( .B1(n10949), .B2(n10527), .A(n10526), .ZN(n10942) );
  AND2_X1 U13153 ( .A1(n10942), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n10940) );
  AOI21_X1 U13154 ( .B1(n10528), .B2(n10613), .A(n10940), .ZN(n10569) );
  MUX2_X1 U13155 ( .A(P3_REG1_REG_2__SCAN_IN), .B(n10516), .S(n10533), .Z(
        n10570) );
  NOR2_X1 U13156 ( .A1(n10569), .A2(n10570), .ZN(n10568) );
  AOI21_X1 U13157 ( .B1(n10584), .B2(P3_REG1_REG_2__SCAN_IN), .A(n10568), .ZN(
        n10799) );
  XNOR2_X1 U13158 ( .A(n10796), .B(n10797), .ZN(n10541) );
  NAND2_X1 U13159 ( .A1(P3_REG2_REG_0__SCAN_IN), .A2(n10529), .ZN(n10609) );
  NAND2_X1 U13160 ( .A1(n9266), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n10531) );
  INV_X1 U13161 ( .A(n10531), .ZN(n10530) );
  AOI21_X1 U13162 ( .B1(n10949), .B2(n10609), .A(n10530), .ZN(n10939) );
  NAND2_X1 U13163 ( .A1(n10939), .A2(P3_REG2_REG_1__SCAN_IN), .ZN(n10938) );
  NAND2_X1 U13164 ( .A1(n10938), .A2(n10531), .ZN(n10566) );
  NAND2_X1 U13165 ( .A1(n10566), .A2(n10567), .ZN(n10565) );
  OAI21_X1 U13166 ( .B1(n10533), .B2(n10532), .A(n10565), .ZN(n10804) );
  XNOR2_X1 U13167 ( .A(n10804), .B(n10798), .ZN(n10806) );
  XNOR2_X1 U13168 ( .A(n10806), .B(n11476), .ZN(n10539) );
  AND2_X1 U13169 ( .A1(n10537), .A2(n10536), .ZN(n15415) );
  INV_X1 U13170 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n11478) );
  NOR2_X1 U13171 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11478), .ZN(n10711) );
  AOI21_X1 U13172 ( .B1(n15415), .B2(P3_ADDR_REG_3__SCAN_IN), .A(n10711), .ZN(
        n10538) );
  OAI21_X1 U13173 ( .B1(n10539), .B2(n15401), .A(n10538), .ZN(n10540) );
  AOI21_X1 U13174 ( .B1(n15426), .B2(n10541), .A(n10540), .ZN(n10542) );
  OAI211_X1 U13175 ( .C1(n11925), .C2(n10805), .A(n10543), .B(n10542), .ZN(
        P3_U3185) );
  NOR2_X1 U13176 ( .A1(n10544), .A2(n15345), .ZN(n10620) );
  NAND2_X1 U13177 ( .A1(n10627), .A2(n15348), .ZN(n10632) );
  INV_X1 U13178 ( .A(n10629), .ZN(n10545) );
  AND2_X1 U13179 ( .A1(n8816), .A2(n13623), .ZN(n10547) );
  NAND2_X1 U13180 ( .A1(n13336), .A2(n13383), .ZN(n10733) );
  OAI21_X1 U13181 ( .B1(n10924), .B2(n10547), .A(n10733), .ZN(n10919) );
  INV_X1 U13182 ( .A(n8890), .ZN(n15362) );
  NAND2_X1 U13183 ( .A1(n10548), .A2(n10727), .ZN(n10917) );
  OAI21_X1 U13184 ( .B1(n10924), .B2(n15362), .A(n10917), .ZN(n10549) );
  NOR2_X1 U13185 ( .A1(n10919), .A2(n10549), .ZN(n15351) );
  NAND2_X1 U13186 ( .A1(n15389), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n10550) );
  OAI21_X1 U13187 ( .B1(n15389), .B2(n15351), .A(n10550), .ZN(P2_U3499) );
  INV_X1 U13188 ( .A(n14993), .ZN(n10551) );
  INV_X1 U13189 ( .A(n10554), .ZN(n10556) );
  OAI211_X1 U13190 ( .C1(n10557), .C2(n15159), .A(n10556), .B(n10555), .ZN(
        n10563) );
  OAI22_X1 U13191 ( .A1(n14748), .A2(n10561), .B1(n15174), .B2(n7708), .ZN(
        n10558) );
  AOI21_X1 U13192 ( .B1(n10563), .B2(n15174), .A(n10558), .ZN(n10559) );
  INV_X1 U13193 ( .A(n10559), .ZN(P1_U3462) );
  OAI22_X1 U13194 ( .A1(n14686), .A2(n10561), .B1(n15185), .B2(n10560), .ZN(
        n10562) );
  AOI21_X1 U13195 ( .B1(n10563), .B2(n15185), .A(n10562), .ZN(n10564) );
  INV_X1 U13196 ( .A(n10564), .ZN(P1_U3529) );
  INV_X1 U13197 ( .A(n15401), .ZN(n15429) );
  OAI21_X1 U13198 ( .B1(n10567), .B2(n10566), .A(n10565), .ZN(n10576) );
  AOI21_X1 U13199 ( .B1(n10570), .B2(n10569), .A(n10568), .ZN(n10571) );
  NOR2_X1 U13200 ( .A1(n12841), .A2(n10571), .ZN(n10575) );
  INV_X1 U13201 ( .A(n15415), .ZN(n15413) );
  INV_X1 U13202 ( .A(P3_ADDR_REG_2__SCAN_IN), .ZN(n10573) );
  OAI22_X1 U13203 ( .A1(n15413), .A2(n10573), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n10572), .ZN(n10574) );
  AOI211_X1 U13204 ( .C1(n15429), .C2(n10576), .A(n10575), .B(n10574), .ZN(
        n10583) );
  INV_X1 U13205 ( .A(n10577), .ZN(n10581) );
  NOR3_X1 U13206 ( .A1(n10935), .A2(n10579), .A3(n10578), .ZN(n10580) );
  OAI21_X1 U13207 ( .B1(n10581), .B2(n10580), .A(n15430), .ZN(n10582) );
  OAI211_X1 U13208 ( .C1(n11925), .C2(n10584), .A(n10583), .B(n10582), .ZN(
        P3_U3184) );
  NOR2_X2 U13209 ( .A1(n10623), .A2(n10585), .ZN(n15355) );
  NAND2_X1 U13210 ( .A1(n15392), .A2(n15355), .ZN(n13749) );
  INV_X1 U13211 ( .A(n10586), .ZN(n10588) );
  AOI211_X1 U13212 ( .C1(n8890), .C2(n10589), .A(n10588), .B(n10587), .ZN(
        n10606) );
  MUX2_X1 U13213 ( .A(n10590), .B(n10606), .S(n15392), .Z(n10591) );
  OAI21_X1 U13214 ( .B1(n10648), .B2(n13749), .A(n10591), .ZN(P2_U3500) );
  OAI21_X1 U13215 ( .B1(n10594), .B2(n10593), .A(n10592), .ZN(n10595) );
  INV_X1 U13216 ( .A(n10595), .ZN(n11199) );
  XNOR2_X1 U13217 ( .A(n10597), .B(n10596), .ZN(n10600) );
  OAI22_X1 U13218 ( .A1(n10599), .A2(n13301), .B1(n10598), .B2(n13303), .ZN(
        n10738) );
  AOI21_X1 U13219 ( .B1(n10600), .B2(n13661), .A(n10738), .ZN(n11205) );
  OAI211_X1 U13220 ( .C1(n13650), .C2(n10736), .A(n10768), .B(n13604), .ZN(
        n11200) );
  OAI211_X1 U13221 ( .C1(n11199), .C2(n13734), .A(n11205), .B(n11200), .ZN(
        n10715) );
  OAI22_X1 U13222 ( .A1(n13749), .A2(n10736), .B1(n15392), .B2(n10601), .ZN(
        n10602) );
  AOI21_X1 U13223 ( .B1(n15392), .B2(n10715), .A(n10602), .ZN(n10603) );
  INV_X1 U13224 ( .A(n10603), .ZN(P2_U3502) );
  INV_X1 U13225 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n10607) );
  MUX2_X1 U13226 ( .A(n10607), .B(n10606), .S(n15383), .Z(n10608) );
  OAI21_X1 U13227 ( .B1(n10648), .B2(n13783), .A(n10608), .ZN(P2_U3433) );
  NOR3_X1 U13228 ( .A1(n15429), .A2(n15426), .A3(n15430), .ZN(n10618) );
  NOR2_X1 U13229 ( .A1(n15401), .A2(n10609), .ZN(n10612) );
  OAI22_X1 U13230 ( .A1(n15413), .A2(n10610), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n11526), .ZN(n10611) );
  AOI211_X1 U13231 ( .C1(n15426), .C2(n10613), .A(n10612), .B(n10611), .ZN(
        n10617) );
  OR2_X1 U13232 ( .A1(n10614), .A2(n15406), .ZN(n10615) );
  MUX2_X1 U13233 ( .A(n10615), .B(n11925), .S(P3_IR_REG_0__SCAN_IN), .Z(n10616) );
  OAI211_X1 U13234 ( .C1(n10618), .C2(n10937), .A(n10617), .B(n10616), .ZN(
        P3_U3182) );
  NAND2_X1 U13235 ( .A1(n10620), .A2(n10619), .ZN(n10637) );
  OR2_X1 U13236 ( .A1(n10637), .A2(n10621), .ZN(n10622) );
  INV_X1 U13237 ( .A(n10637), .ZN(n10624) );
  INV_X1 U13238 ( .A(n15345), .ZN(n10625) );
  NAND2_X1 U13239 ( .A1(n10626), .A2(n10625), .ZN(n10628) );
  NAND2_X1 U13240 ( .A1(n10628), .A2(n10627), .ZN(n10634) );
  AND4_X1 U13241 ( .A1(n10632), .A2(n10631), .A3(n10630), .A4(n10629), .ZN(
        n10633) );
  NAND2_X1 U13242 ( .A1(n10634), .A2(n10633), .ZN(n10737) );
  OR2_X1 U13243 ( .A1(n10737), .A2(P2_U3088), .ZN(n10729) );
  AOI22_X1 U13244 ( .A1(n15190), .A2(n10635), .B1(P2_REG3_REG_1__SCAN_IN), 
        .B2(n10729), .ZN(n10647) );
  INV_X1 U13245 ( .A(n10648), .ZN(n10638) );
  NAND2_X1 U13246 ( .A1(n10653), .A2(n13383), .ZN(n10660) );
  NAND2_X1 U13247 ( .A1(n13255), .A2(n10639), .ZN(n10642) );
  NAND2_X1 U13248 ( .A1(n13588), .A2(n10727), .ZN(n10640) );
  NAND2_X1 U13249 ( .A1(n10642), .A2(n10728), .ZN(n10644) );
  NAND2_X1 U13250 ( .A1(n10644), .A2(n10643), .ZN(n10663) );
  OAI21_X1 U13251 ( .B1(n10643), .B2(n10644), .A(n10663), .ZN(n10645) );
  NAND2_X1 U13252 ( .A1(n15193), .A2(n10645), .ZN(n10646) );
  OAI211_X1 U13253 ( .C1(n10648), .C2(n13331), .A(n10647), .B(n10646), .ZN(
        P2_U3194) );
  OAI22_X1 U13254 ( .A1(n10650), .A2(n13301), .B1(n10649), .B2(n13303), .ZN(
        n13660) );
  AOI22_X1 U13255 ( .A1(n15190), .A2(n13660), .B1(P2_REG3_REG_2__SCAN_IN), 
        .B2(n10729), .ZN(n10668) );
  NAND2_X1 U13256 ( .A1(n10653), .A2(n13382), .ZN(n10655) );
  NAND2_X1 U13257 ( .A1(n10654), .A2(n10655), .ZN(n10734) );
  INV_X1 U13258 ( .A(n10654), .ZN(n10657) );
  INV_X1 U13259 ( .A(n10655), .ZN(n10656) );
  NAND2_X1 U13260 ( .A1(n10657), .A2(n10656), .ZN(n10658) );
  AND2_X1 U13261 ( .A1(n10734), .A2(n10658), .ZN(n10665) );
  INV_X1 U13262 ( .A(n10659), .ZN(n10661) );
  NAND2_X1 U13263 ( .A1(n10661), .A2(n10660), .ZN(n10662) );
  NAND2_X1 U13264 ( .A1(n10663), .A2(n10662), .ZN(n10664) );
  OAI21_X1 U13265 ( .B1(n10665), .B2(n10664), .A(n10735), .ZN(n10666) );
  NAND2_X1 U13266 ( .A1(n15193), .A2(n10666), .ZN(n10667) );
  OAI211_X1 U13267 ( .C1(n10651), .C2(n13331), .A(n10668), .B(n10667), .ZN(
        P2_U3209) );
  INV_X1 U13268 ( .A(n10692), .ZN(n10674) );
  INV_X1 U13269 ( .A(n10693), .ZN(n10669) );
  OR2_X1 U13270 ( .A1(n10705), .A2(n10669), .ZN(n10673) );
  AND3_X1 U13271 ( .A1(n10671), .A2(n10670), .A3(n11359), .ZN(n10672) );
  OAI211_X1 U13272 ( .C1(n10700), .C2(n10674), .A(n10673), .B(n10672), .ZN(
        n10675) );
  NAND2_X1 U13273 ( .A1(n10675), .A2(P3_STATE_REG_SCAN_IN), .ZN(n10677) );
  OR2_X1 U13274 ( .A1(n10705), .A2(n12721), .ZN(n10676) );
  NAND2_X1 U13275 ( .A1(n11322), .A2(n12847), .ZN(n10679) );
  NAND2_X1 U13276 ( .A1(n12360), .A2(n11370), .ZN(n10682) );
  NAND2_X1 U13277 ( .A1(n10678), .A2(n10681), .ZN(n10687) );
  OAI21_X1 U13278 ( .B1(n10678), .B2(n10682), .A(n10687), .ZN(n10683) );
  INV_X1 U13279 ( .A(n10683), .ZN(n11020) );
  NAND2_X1 U13280 ( .A1(n11366), .A2(n12360), .ZN(n10684) );
  NAND2_X1 U13281 ( .A1(n10685), .A2(n10684), .ZN(n10686) );
  NAND2_X1 U13282 ( .A1(n11020), .A2(n10686), .ZN(n11019) );
  NAND2_X1 U13283 ( .A1(n11019), .A2(n10687), .ZN(n10951) );
  XNOR2_X1 U13284 ( .A(n10688), .B(n10709), .ZN(n10952) );
  NAND2_X1 U13285 ( .A1(n10951), .A2(n10952), .ZN(n10691) );
  INV_X1 U13286 ( .A(n10688), .ZN(n10689) );
  NAND2_X1 U13287 ( .A1(n10689), .A2(n10709), .ZN(n10690) );
  XNOR2_X1 U13288 ( .A(n11479), .B(n12392), .ZN(n11002) );
  XNOR2_X1 U13289 ( .A(n11002), .B(n15451), .ZN(n10697) );
  NAND3_X1 U13290 ( .A1(n10700), .A2(n10692), .A3(n15486), .ZN(n10695) );
  NAND2_X1 U13291 ( .A1(n10705), .A2(n10693), .ZN(n10694) );
  NAND2_X1 U13292 ( .A1(n10695), .A2(n10694), .ZN(n10696) );
  NAND2_X1 U13293 ( .A1(n10698), .A2(n11005), .ZN(n10713) );
  AND2_X1 U13294 ( .A1(n10702), .A2(n15479), .ZN(n10699) );
  NAND2_X1 U13295 ( .A1(n10700), .A2(n10699), .ZN(n10703) );
  INV_X1 U13296 ( .A(n12705), .ZN(n15459) );
  NOR2_X1 U13297 ( .A1(n15486), .A2(n15459), .ZN(n10701) );
  INV_X1 U13298 ( .A(n12721), .ZN(n10704) );
  NAND2_X1 U13299 ( .A1(n10705), .A2(n10704), .ZN(n10708) );
  OAI22_X1 U13300 ( .A1(n10709), .A2(n12500), .B1(n11314), .B2(n12489), .ZN(
        n10710) );
  AOI211_X1 U13301 ( .C1(n11479), .C2(n12491), .A(n10711), .B(n10710), .ZN(
        n10712) );
  OAI211_X1 U13302 ( .C1(P3_REG3_REG_3__SCAN_IN), .C2(n12503), .A(n10713), .B(
        n10712), .ZN(P3_U3158) );
  OAI22_X1 U13303 ( .A1(n13783), .A2(n10736), .B1(n15383), .B2(n8414), .ZN(
        n10714) );
  AOI21_X1 U13304 ( .B1(n15383), .B2(n10715), .A(n10714), .ZN(n10716) );
  INV_X1 U13305 ( .A(n10716), .ZN(P2_U3439) );
  AND2_X1 U13306 ( .A1(n12741), .A2(n11527), .ZN(n12526) );
  NOR2_X1 U13307 ( .A1(n12529), .A2(n12526), .ZN(n12678) );
  OR2_X1 U13308 ( .A1(n10717), .A2(n15479), .ZN(n10718) );
  OR2_X1 U13309 ( .A1(n12678), .A2(n10718), .ZN(n10721) );
  NAND2_X1 U13310 ( .A1(n10719), .A2(n13029), .ZN(n10720) );
  NAND2_X1 U13311 ( .A1(n10721), .A2(n10720), .ZN(n11525) );
  INV_X1 U13312 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n10722) );
  OAI22_X1 U13313 ( .A1(n11527), .A2(n13144), .B1(n15493), .B2(n10722), .ZN(
        n10723) );
  AOI21_X1 U13314 ( .B1(n11525), .B2(n15493), .A(n10723), .ZN(n10724) );
  INV_X1 U13315 ( .A(n10724), .ZN(P3_U3390) );
  OAI222_X1 U13316 ( .A1(n13172), .A2(n10726), .B1(n13167), .B2(n10725), .C1(
        P3_U3151), .C2(n12832), .ZN(P3_U3276) );
  NAND2_X1 U13317 ( .A1(n15195), .A2(n10727), .ZN(n10732) );
  OAI21_X1 U13318 ( .B1(n13604), .B2(n9142), .A(n10728), .ZN(n10730) );
  AOI22_X1 U13319 ( .A1(n15193), .A2(n10730), .B1(P2_REG3_REG_0__SCAN_IN), 
        .B2(n10729), .ZN(n10731) );
  OAI211_X1 U13320 ( .C1(n13347), .C2(n10733), .A(n10732), .B(n10731), .ZN(
        P2_U3204) );
  XNOR2_X1 U13321 ( .A(n10652), .B(n10736), .ZN(n10824) );
  NAND2_X1 U13322 ( .A1(n10653), .A2(n13381), .ZN(n10825) );
  XNOR2_X1 U13323 ( .A(n10824), .B(n10825), .ZN(n10829) );
  XNOR2_X1 U13324 ( .A(n10830), .B(n10829), .ZN(n10742) );
  NAND2_X1 U13325 ( .A1(n15190), .A2(n10738), .ZN(n10739) );
  NAND2_X1 U13326 ( .A1(P2_U3088), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n15238) );
  OAI211_X1 U13327 ( .C1(P2_REG3_REG_3__SCAN_IN), .C2(n15198), .A(n10739), .B(
        n15238), .ZN(n10740) );
  AOI21_X1 U13328 ( .B1(n11203), .B2(n15195), .A(n10740), .ZN(n10741) );
  OAI21_X1 U13329 ( .B1(n10742), .B2(n13349), .A(n10741), .ZN(P2_U3190) );
  AOI22_X1 U13330 ( .A1(n15000), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n11286), .ZN(n10743) );
  OAI21_X1 U13331 ( .B1(n10821), .B2(n14761), .A(n10743), .ZN(P1_U3341) );
  INV_X1 U13332 ( .A(n15159), .ZN(n15137) );
  OAI21_X1 U13333 ( .B1(n10746), .B2(n10745), .A(n10744), .ZN(n10753) );
  INV_X1 U13334 ( .A(n10974), .ZN(n10747) );
  AOI211_X1 U13335 ( .C1(n13984), .C2(n11063), .A(n14915), .B(n10747), .ZN(
        n11035) );
  INV_X1 U13336 ( .A(n10753), .ZN(n11038) );
  OAI21_X1 U13337 ( .B1(n10749), .B2(n14170), .A(n10748), .ZN(n10751) );
  OAI22_X1 U13338 ( .A1(n11192), .A2(n14919), .B1(n13976), .B2(n14601), .ZN(
        n10750) );
  AOI21_X1 U13339 ( .B1(n10751), .B2(n14952), .A(n10750), .ZN(n10752) );
  OAI21_X1 U13340 ( .B1(n11038), .B2(n15129), .A(n10752), .ZN(n11031) );
  AOI211_X1 U13341 ( .C1(n15137), .C2(n10753), .A(n11035), .B(n11031), .ZN(
        n10758) );
  INV_X1 U13342 ( .A(n13984), .ZN(n13983) );
  OAI22_X1 U13343 ( .A1(n14686), .A2(n13983), .B1(n15185), .B2(n7771), .ZN(
        n10754) );
  INV_X1 U13344 ( .A(n10754), .ZN(n10755) );
  OAI21_X1 U13345 ( .B1(n10758), .B2(n15183), .A(n10755), .ZN(P1_U3531) );
  OAI22_X1 U13346 ( .A1(n14748), .A2(n13983), .B1(n15174), .B2(n6803), .ZN(
        n10756) );
  INV_X1 U13347 ( .A(n10756), .ZN(n10757) );
  OAI21_X1 U13348 ( .B1(n10758), .B2(n15172), .A(n10757), .ZN(P1_U3468) );
  OAI21_X1 U13349 ( .B1(n10761), .B2(n10760), .A(n10759), .ZN(n10762) );
  INV_X1 U13350 ( .A(n10762), .ZN(n11137) );
  XNOR2_X1 U13351 ( .A(n10764), .B(n10763), .ZN(n10766) );
  AOI22_X1 U13352 ( .A1(n13337), .A2(n13381), .B1(n13336), .B2(n13379), .ZN(
        n10841) );
  INV_X1 U13353 ( .A(n10841), .ZN(n10765) );
  AOI21_X1 U13354 ( .B1(n10766), .B2(n13661), .A(n10765), .ZN(n11134) );
  INV_X1 U13355 ( .A(n10960), .ZN(n10767) );
  AOI211_X1 U13356 ( .C1(n10843), .C2(n10768), .A(n13651), .B(n10767), .ZN(
        n11132) );
  INV_X1 U13357 ( .A(n11132), .ZN(n10769) );
  OAI211_X1 U13358 ( .C1(n11137), .C2(n13734), .A(n11134), .B(n10769), .ZN(
        n10774) );
  INV_X1 U13359 ( .A(n10843), .ZN(n11130) );
  OAI22_X1 U13360 ( .A1(n13783), .A2(n11130), .B1(n15383), .B2(n8426), .ZN(
        n10770) );
  AOI21_X1 U13361 ( .B1(n10774), .B2(n15383), .A(n10770), .ZN(n10771) );
  INV_X1 U13362 ( .A(n10771), .ZN(P2_U3442) );
  OAI22_X1 U13363 ( .A1(n13749), .A2(n11130), .B1(n15392), .B2(n10772), .ZN(
        n10773) );
  AOI21_X1 U13364 ( .B1(n10774), .B2(n15392), .A(n10773), .ZN(n10775) );
  INV_X1 U13365 ( .A(n10775), .ZN(P2_U3503) );
  OAI21_X1 U13366 ( .B1(n10777), .B2(n12677), .A(n10776), .ZN(n11474) );
  OAI211_X1 U13367 ( .C1(n10780), .C2(n10779), .A(n13032), .B(n10778), .ZN(
        n10783) );
  AOI22_X1 U13368 ( .A1(n13027), .A2(n10781), .B1(n12738), .B2(n13029), .ZN(
        n10782) );
  NAND2_X1 U13369 ( .A1(n10783), .A2(n10782), .ZN(n11475) );
  AOI21_X1 U13370 ( .B1(n15477), .B2(n11474), .A(n11475), .ZN(n11244) );
  INV_X1 U13371 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n10784) );
  OAI22_X1 U13372 ( .A1(n10785), .A2(n13144), .B1(n15493), .B2(n10784), .ZN(
        n10786) );
  INV_X1 U13373 ( .A(n10786), .ZN(n10787) );
  OAI21_X1 U13374 ( .B1(n11244), .B2(n15491), .A(n10787), .ZN(P3_U3399) );
  MUX2_X1 U13375 ( .A(P3_REG2_REG_7__SCAN_IN), .B(P3_REG1_REG_7__SCAN_IN), .S(
        n13165), .Z(n10892) );
  XNOR2_X1 U13376 ( .A(n10892), .B(n10900), .ZN(n10893) );
  MUX2_X1 U13377 ( .A(P3_REG2_REG_4__SCAN_IN), .B(P3_REG1_REG_4__SCAN_IN), .S(
        n13165), .Z(n10791) );
  INV_X1 U13378 ( .A(n10791), .ZN(n10792) );
  INV_X1 U13379 ( .A(n10788), .ZN(n10789) );
  XOR2_X1 U13380 ( .A(n15410), .B(n10791), .Z(n15404) );
  AOI21_X1 U13381 ( .B1(n15410), .B2(n10792), .A(n15403), .ZN(n10866) );
  MUX2_X1 U13382 ( .A(n10067), .B(n10868), .S(n13165), .Z(n10793) );
  NOR2_X1 U13383 ( .A1(n10793), .A2(n10808), .ZN(n10862) );
  NAND2_X1 U13384 ( .A1(n10793), .A2(n10808), .ZN(n10863) );
  MUX2_X1 U13385 ( .A(P3_REG2_REG_6__SCAN_IN), .B(P3_REG1_REG_6__SCAN_IN), .S(
        n13165), .Z(n10794) );
  XNOR2_X1 U13386 ( .A(n10794), .B(n10809), .ZN(n10847) );
  INV_X1 U13387 ( .A(n10794), .ZN(n10795) );
  XOR2_X1 U13388 ( .A(n10894), .B(n10893), .Z(n10820) );
  AOI22_X1 U13389 ( .A1(n10809), .A2(n9319), .B1(P3_REG1_REG_6__SCAN_IN), .B2(
        n10849), .ZN(n10855) );
  MUX2_X1 U13390 ( .A(n10800), .B(P3_REG1_REG_4__SCAN_IN), .S(n15410), .Z(
        n15398) );
  OAI21_X1 U13391 ( .B1(n15410), .B2(n10800), .A(n15396), .ZN(n10801) );
  XNOR2_X1 U13392 ( .A(n10801), .B(n10874), .ZN(n10869) );
  INV_X1 U13393 ( .A(n10801), .ZN(n10802) );
  OAI22_X1 U13394 ( .A1(n10869), .A2(n10868), .B1(n10808), .B2(n10802), .ZN(
        n10856) );
  OAI21_X1 U13395 ( .B1(n10803), .B2(P3_REG1_REG_7__SCAN_IN), .A(n10896), .ZN(
        n10818) );
  INV_X1 U13396 ( .A(P3_ADDR_REG_7__SCAN_IN), .ZN(n10815) );
  INV_X1 U13397 ( .A(P3_REG2_REG_6__SCAN_IN), .ZN(n15445) );
  AOI22_X1 U13398 ( .A1(n10809), .A2(n15445), .B1(P3_REG2_REG_6__SCAN_IN), 
        .B2(n10849), .ZN(n10852) );
  AOI22_X1 U13399 ( .A1(n10806), .A2(P3_REG2_REG_3__SCAN_IN), .B1(n10805), 
        .B2(n10804), .ZN(n15395) );
  INV_X1 U13400 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n11398) );
  MUX2_X1 U13401 ( .A(P3_REG2_REG_4__SCAN_IN), .B(n11398), .S(n15410), .Z(
        n15394) );
  NOR2_X1 U13402 ( .A1(n15395), .A2(n15394), .ZN(n15393) );
  NAND2_X1 U13403 ( .A1(n10852), .A2(n10853), .ZN(n10851) );
  OAI21_X1 U13404 ( .B1(n10809), .B2(n15445), .A(n10851), .ZN(n10901) );
  XNOR2_X1 U13405 ( .A(n10901), .B(n10810), .ZN(n10811) );
  NAND2_X1 U13406 ( .A1(P3_REG2_REG_7__SCAN_IN), .A2(n10811), .ZN(n10902) );
  OAI21_X1 U13407 ( .B1(n10811), .B2(P3_REG2_REG_7__SCAN_IN), .A(n10902), .ZN(
        n10812) );
  NAND2_X1 U13408 ( .A1(n15429), .A2(n10812), .ZN(n10814) );
  AND2_X1 U13409 ( .A1(P3_U3151), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n11446) );
  INV_X1 U13410 ( .A(n11446), .ZN(n10813) );
  OAI211_X1 U13411 ( .C1(n15413), .C2(n10815), .A(n10814), .B(n10813), .ZN(
        n10817) );
  NOR2_X1 U13412 ( .A1(n11925), .A2(n10900), .ZN(n10816) );
  AOI211_X1 U13413 ( .C1(n15426), .C2(n10818), .A(n10817), .B(n10816), .ZN(
        n10819) );
  OAI21_X1 U13414 ( .B1(n10820), .B2(n15406), .A(n10819), .ZN(P3_U3189) );
  INV_X1 U13415 ( .A(n15317), .ZN(n10822) );
  OAI222_X1 U13416 ( .A1(n13798), .A2(n10823), .B1(n10822), .B2(P2_U3088), 
        .C1(n13804), .C2(n10821), .ZN(P2_U3313) );
  INV_X1 U13417 ( .A(n10824), .ZN(n10827) );
  INV_X1 U13418 ( .A(n10825), .ZN(n10826) );
  NAND2_X1 U13419 ( .A1(n10827), .A2(n10826), .ZN(n10828) );
  XNOR2_X1 U13420 ( .A(n13255), .B(n6873), .ZN(n10831) );
  NAND2_X1 U13421 ( .A1(n10653), .A2(n13380), .ZN(n10832) );
  NAND2_X1 U13422 ( .A1(n10831), .A2(n10832), .ZN(n10885) );
  INV_X1 U13423 ( .A(n10831), .ZN(n10834) );
  INV_X1 U13424 ( .A(n10832), .ZN(n10833) );
  NAND2_X1 U13425 ( .A1(n10834), .A2(n10833), .ZN(n10835) );
  NAND2_X1 U13426 ( .A1(n10885), .A2(n10835), .ZN(n10837) );
  INV_X1 U13427 ( .A(n10886), .ZN(n10836) );
  AOI21_X1 U13428 ( .B1(n10838), .B2(n10837), .A(n10836), .ZN(n10845) );
  NAND2_X1 U13429 ( .A1(n13344), .A2(n11128), .ZN(n10839) );
  OAI211_X1 U13430 ( .C1(n13347), .C2(n10841), .A(n10840), .B(n10839), .ZN(
        n10842) );
  AOI21_X1 U13431 ( .B1(n10843), .B2(n15195), .A(n10842), .ZN(n10844) );
  OAI21_X1 U13432 ( .B1(n10845), .B2(n13349), .A(n10844), .ZN(P2_U3202) );
  XOR2_X1 U13433 ( .A(n10846), .B(n10847), .Z(n10861) );
  INV_X1 U13434 ( .A(P3_REG3_REG_6__SCAN_IN), .ZN(n10848) );
  NOR2_X1 U13435 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10848), .ZN(n11515) );
  NOR2_X1 U13436 ( .A1(n11925), .A2(n10849), .ZN(n10850) );
  AOI211_X1 U13437 ( .C1(n15415), .C2(P3_ADDR_REG_6__SCAN_IN), .A(n11515), .B(
        n10850), .ZN(n10860) );
  OAI21_X1 U13438 ( .B1(n10853), .B2(n10852), .A(n10851), .ZN(n10858) );
  OAI21_X1 U13439 ( .B1(n10856), .B2(n10855), .A(n10854), .ZN(n10857) );
  AOI22_X1 U13440 ( .A1(n15429), .A2(n10858), .B1(n15426), .B2(n10857), .ZN(
        n10859) );
  OAI211_X1 U13441 ( .C1(n10861), .C2(n15406), .A(n10860), .B(n10859), .ZN(
        P3_U3188) );
  INV_X1 U13442 ( .A(n10862), .ZN(n10864) );
  NAND2_X1 U13443 ( .A1(n10864), .A2(n10863), .ZN(n10865) );
  XNOR2_X1 U13444 ( .A(n10866), .B(n10865), .ZN(n10876) );
  XNOR2_X1 U13445 ( .A(n10867), .B(n10067), .ZN(n10871) );
  XNOR2_X1 U13446 ( .A(n10869), .B(n10868), .ZN(n10870) );
  AOI22_X1 U13447 ( .A1(n15429), .A2(n10871), .B1(n15426), .B2(n10870), .ZN(
        n10873) );
  AND2_X1 U13448 ( .A1(P3_U3151), .A2(P3_REG3_REG_5__SCAN_IN), .ZN(n11154) );
  AOI21_X1 U13449 ( .B1(n15415), .B2(P3_ADDR_REG_5__SCAN_IN), .A(n11154), .ZN(
        n10872) );
  OAI211_X1 U13450 ( .C1(n11925), .C2(n10874), .A(n10873), .B(n10872), .ZN(
        n10875) );
  AOI21_X1 U13451 ( .B1(n10876), .B2(n15430), .A(n10875), .ZN(n10877) );
  INV_X1 U13452 ( .A(n10877), .ZN(P3_U3187) );
  AOI22_X1 U13453 ( .A1(n13337), .A2(n13380), .B1(n13336), .B2(n13378), .ZN(
        n10963) );
  NOR2_X1 U13454 ( .A1(n13347), .A2(n10963), .ZN(n10878) );
  AOI211_X1 U13455 ( .C1(n13344), .C2(n11327), .A(n10879), .B(n10878), .ZN(
        n10891) );
  XNOR2_X1 U13456 ( .A(n13213), .B(n10965), .ZN(n10880) );
  NAND2_X1 U13457 ( .A1(n13651), .A2(n13379), .ZN(n10881) );
  NAND2_X1 U13458 ( .A1(n10880), .A2(n10881), .ZN(n10925) );
  INV_X1 U13459 ( .A(n10880), .ZN(n10883) );
  INV_X1 U13460 ( .A(n10881), .ZN(n10882) );
  NAND2_X1 U13461 ( .A1(n10883), .A2(n10882), .ZN(n10884) );
  AND2_X1 U13462 ( .A1(n10925), .A2(n10884), .ZN(n10888) );
  NAND2_X1 U13463 ( .A1(n10886), .A2(n10885), .ZN(n10887) );
  OAI21_X1 U13464 ( .B1(n10888), .B2(n10887), .A(n10926), .ZN(n10889) );
  NAND2_X1 U13465 ( .A1(n10889), .A2(n15193), .ZN(n10890) );
  OAI211_X1 U13466 ( .C1(n11330), .C2(n13331), .A(n10891), .B(n10890), .ZN(
        P2_U3199) );
  MUX2_X1 U13467 ( .A(P3_REG2_REG_8__SCAN_IN), .B(P3_REG1_REG_8__SCAN_IN), .S(
        n13165), .Z(n11071) );
  XNOR2_X1 U13468 ( .A(n11071), .B(n11080), .ZN(n11073) );
  OAI22_X1 U13469 ( .A1(n10894), .A2(n10893), .B1(n10892), .B2(n10900), .ZN(
        n11074) );
  XOR2_X1 U13470 ( .A(n11073), .B(n11074), .Z(n10912) );
  AOI22_X1 U13471 ( .A1(P3_REG1_REG_8__SCAN_IN), .A2(n11076), .B1(n11080), 
        .B2(n9350), .ZN(n10899) );
  NAND2_X1 U13472 ( .A1(n10895), .A2(n10900), .ZN(n10897) );
  NAND2_X1 U13473 ( .A1(n10897), .A2(n10896), .ZN(n10898) );
  NAND2_X1 U13474 ( .A1(n10899), .A2(n10898), .ZN(n11075) );
  OAI21_X1 U13475 ( .B1(n10899), .B2(n10898), .A(n11075), .ZN(n10910) );
  INV_X1 U13476 ( .A(P3_REG2_REG_8__SCAN_IN), .ZN(n11079) );
  AOI22_X1 U13477 ( .A1(P3_REG2_REG_8__SCAN_IN), .A2(n11076), .B1(n11080), 
        .B2(n11079), .ZN(n10905) );
  NAND2_X1 U13478 ( .A1(n10901), .A2(n10900), .ZN(n10903) );
  OAI21_X1 U13479 ( .B1(n10905), .B2(n10904), .A(n11078), .ZN(n10906) );
  NAND2_X1 U13480 ( .A1(n10906), .A2(n15429), .ZN(n10908) );
  AND2_X1 U13481 ( .A1(P3_REG3_REG_8__SCAN_IN), .A2(P3_U3151), .ZN(n11579) );
  AOI21_X1 U13482 ( .B1(n15415), .B2(P3_ADDR_REG_8__SCAN_IN), .A(n11579), .ZN(
        n10907) );
  OAI211_X1 U13483 ( .C1(n11925), .C2(n11076), .A(n10908), .B(n10907), .ZN(
        n10909) );
  AOI21_X1 U13484 ( .B1(n15426), .B2(n10910), .A(n10909), .ZN(n10911) );
  OAI21_X1 U13485 ( .B1(n10912), .B2(n15406), .A(n10911), .ZN(P3_U3190) );
  AOI22_X1 U13486 ( .A1(n10719), .A2(n12506), .B1(n10913), .B2(n12491), .ZN(
        n10915) );
  NAND2_X1 U13487 ( .A1(n12503), .A2(P3_STATE_REG_SCAN_IN), .ZN(n11015) );
  NAND2_X1 U13488 ( .A1(n11015), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n10914) );
  OAI211_X1 U13489 ( .C1(n12678), .C2(n12494), .A(n10915), .B(n10914), .ZN(
        P3_U3172) );
  NOR2_X1 U13490 ( .A1(n10917), .A2(n10916), .ZN(n10918) );
  NOR2_X1 U13491 ( .A1(n10919), .A2(n10918), .ZN(n10921) );
  INV_X1 U13492 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n10920) );
  OAI22_X1 U13493 ( .A1(n6620), .A2(n10921), .B1(n10920), .B2(n13655), .ZN(
        n10922) );
  AOI21_X1 U13494 ( .B1(P2_REG2_REG_0__SCAN_IN), .B2(n6620), .A(n10922), .ZN(
        n10923) );
  OAI21_X1 U13495 ( .B1(n10924), .B2(n11588), .A(n10923), .ZN(P2_U3265) );
  XNOR2_X1 U13496 ( .A(n11123), .B(n13213), .ZN(n11090) );
  NAND2_X1 U13497 ( .A1(n13651), .A2(n13378), .ZN(n11089) );
  XNOR2_X1 U13498 ( .A(n11090), .B(n11089), .ZN(n11091) );
  XNOR2_X1 U13499 ( .A(n11092), .B(n11091), .ZN(n10933) );
  OAI22_X1 U13500 ( .A1(n10928), .A2(n13301), .B1(n10927), .B2(n13303), .ZN(
        n11120) );
  NAND2_X1 U13501 ( .A1(n15190), .A2(n11120), .ZN(n10930) );
  OAI211_X1 U13502 ( .C1(n15198), .C2(n11142), .A(n10930), .B(n10929), .ZN(
        n10931) );
  AOI21_X1 U13503 ( .B1(n11123), .B2(n15195), .A(n10931), .ZN(n10932) );
  OAI21_X1 U13504 ( .B1(n10933), .B2(n13349), .A(n10932), .ZN(P2_U3211) );
  OAI22_X1 U13505 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11027), .B1(n10934), .B2(
        n15413), .ZN(n10948) );
  AOI21_X1 U13506 ( .B1(n10937), .B2(n10936), .A(n10935), .ZN(n10946) );
  OAI21_X1 U13507 ( .B1(P3_REG2_REG_1__SCAN_IN), .B2(n10939), .A(n10938), .ZN(
        n10944) );
  INV_X1 U13508 ( .A(n10940), .ZN(n10941) );
  OAI21_X1 U13509 ( .B1(P3_REG1_REG_1__SCAN_IN), .B2(n10942), .A(n10941), .ZN(
        n10943) );
  AOI22_X1 U13510 ( .A1(n15429), .A2(n10944), .B1(n15426), .B2(n10943), .ZN(
        n10945) );
  OAI21_X1 U13511 ( .B1(n10946), .B2(n15406), .A(n10945), .ZN(n10947) );
  AOI211_X1 U13512 ( .C1(n15417), .C2(n10949), .A(n10948), .B(n10947), .ZN(
        n10950) );
  INV_X1 U13513 ( .A(n10950), .ZN(P3_U3183) );
  XOR2_X1 U13514 ( .A(n10951), .B(n10952), .Z(n10957) );
  AOI22_X1 U13515 ( .A1(n10719), .A2(n12485), .B1(n10953), .B2(n12491), .ZN(
        n10954) );
  OAI21_X1 U13516 ( .B1(n15451), .B2(n12489), .A(n10954), .ZN(n10955) );
  AOI21_X1 U13517 ( .B1(P3_REG3_REG_2__SCAN_IN), .B2(n11015), .A(n10955), .ZN(
        n10956) );
  OAI21_X1 U13518 ( .B1(n10957), .B2(n12494), .A(n10956), .ZN(P3_U3177) );
  OAI21_X1 U13519 ( .B1(n10959), .B2(n10961), .A(n10958), .ZN(n11332) );
  AOI211_X1 U13520 ( .C1(n10965), .C2(n10960), .A(n13651), .B(n11115), .ZN(
        n11326) );
  XNOR2_X1 U13521 ( .A(n10962), .B(n10961), .ZN(n10964) );
  OAI21_X1 U13522 ( .B1(n10964), .B2(n13623), .A(n10963), .ZN(n11325) );
  AOI211_X1 U13523 ( .C1(n15381), .C2(n11332), .A(n11326), .B(n11325), .ZN(
        n10969) );
  INV_X1 U13524 ( .A(n13749), .ZN(n12144) );
  AOI22_X1 U13525 ( .A1(n12144), .A2(n10965), .B1(n15389), .B2(
        P2_REG1_REG_5__SCAN_IN), .ZN(n10966) );
  OAI21_X1 U13526 ( .B1(n10969), .B2(n15389), .A(n10966), .ZN(P2_U3504) );
  OAI22_X1 U13527 ( .A1(n13783), .A2(n11330), .B1(n15383), .B2(n8447), .ZN(
        n10967) );
  INV_X1 U13528 ( .A(n10967), .ZN(n10968) );
  OAI21_X1 U13529 ( .B1(n10969), .B2(n15382), .A(n10968), .ZN(P2_U3445) );
  XNOR2_X1 U13530 ( .A(n13990), .B(n6624), .ZN(n14172) );
  XOR2_X1 U13531 ( .A(n14172), .B(n10970), .Z(n10971) );
  OAI222_X1 U13532 ( .A1(n14919), .A2(n11213), .B1(n14601), .B2(n13985), .C1(
        n15075), .C2(n10971), .ZN(n15118) );
  INV_X1 U13533 ( .A(n15118), .ZN(n10981) );
  XOR2_X1 U13534 ( .A(n10972), .B(n14172), .Z(n15120) );
  NAND2_X1 U13535 ( .A1(n15129), .A2(n13951), .ZN(n10973) );
  INV_X1 U13536 ( .A(n11040), .ZN(n10976) );
  AOI21_X1 U13537 ( .B1(n10974), .B2(n13990), .A(n14915), .ZN(n10975) );
  NAND2_X1 U13538 ( .A1(n10976), .A2(n10975), .ZN(n15116) );
  OAI22_X1 U13539 ( .A1(n14539), .A2(n9929), .B1(n11211), .B2(n14602), .ZN(
        n10977) );
  AOI21_X1 U13540 ( .B1(n15081), .B2(n13990), .A(n10977), .ZN(n10978) );
  OAI21_X1 U13541 ( .B1(n14557), .B2(n15116), .A(n10978), .ZN(n10979) );
  AOI21_X1 U13542 ( .B1(n15120), .B2(n14609), .A(n10979), .ZN(n10980) );
  OAI21_X1 U13543 ( .B1(n10981), .B2(n15105), .A(n10980), .ZN(P1_U3289) );
  OAI21_X1 U13544 ( .B1(n10983), .B2(n11162), .A(n10982), .ZN(n14283) );
  MUX2_X1 U13545 ( .A(n11230), .B(P1_REG2_REG_8__SCAN_IN), .S(n10990), .Z(
        n14282) );
  NAND2_X1 U13546 ( .A1(n14283), .A2(n14282), .ZN(n14281) );
  OAI21_X1 U13547 ( .B1(n11230), .B2(n10990), .A(n14281), .ZN(n14297) );
  MUX2_X1 U13548 ( .A(P1_REG2_REG_9__SCAN_IN), .B(n14604), .S(n14294), .Z(
        n14296) );
  NAND2_X1 U13549 ( .A1(n14297), .A2(n14296), .ZN(n14295) );
  OAI21_X1 U13550 ( .B1(n10984), .B2(n14604), .A(n14295), .ZN(n10986) );
  MUX2_X1 U13551 ( .A(P1_REG2_REG_10__SCAN_IN), .B(n11638), .S(n11104), .Z(
        n10985) );
  AND2_X1 U13552 ( .A1(n10986), .A2(n10985), .ZN(n11103) );
  OAI21_X1 U13553 ( .B1(n10986), .B2(n10985), .A(n15012), .ZN(n11001) );
  MUX2_X1 U13554 ( .A(n10987), .B(P1_REG1_REG_10__SCAN_IN), .S(n11104), .Z(
        n10994) );
  MUX2_X1 U13555 ( .A(n10991), .B(P1_REG1_REG_8__SCAN_IN), .S(n10990), .Z(
        n14274) );
  NAND2_X1 U13556 ( .A1(n14275), .A2(n14274), .ZN(n14273) );
  OAI21_X1 U13557 ( .B1(n14280), .B2(P1_REG1_REG_8__SCAN_IN), .A(n14273), .ZN(
        n14288) );
  MUX2_X1 U13558 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n10992), .S(n14294), .Z(
        n14289) );
  NAND2_X1 U13559 ( .A1(n14288), .A2(n14289), .ZN(n14287) );
  OAI21_X1 U13560 ( .B1(P1_REG1_REG_9__SCAN_IN), .B2(n14294), .A(n14287), .ZN(
        n10993) );
  NOR2_X1 U13561 ( .A1(n10993), .A2(n10994), .ZN(n11099) );
  AOI211_X1 U13562 ( .C1(n10994), .C2(n10993), .A(n15056), .B(n11099), .ZN(
        n10999) );
  NAND2_X1 U13563 ( .A1(P1_REG3_REG_10__SCAN_IN), .A2(P1_U3086), .ZN(n10996)
         );
  NAND2_X1 U13564 ( .A1(n14981), .A2(P1_ADDR_REG_10__SCAN_IN), .ZN(n10995) );
  OAI211_X1 U13565 ( .C1(n15037), .C2(n10997), .A(n10996), .B(n10995), .ZN(
        n10998) );
  NOR2_X1 U13566 ( .A1(n10999), .A2(n10998), .ZN(n11000) );
  OAI21_X1 U13567 ( .B1(n11103), .B2(n11001), .A(n11000), .ZN(P1_U3253) );
  XNOR2_X1 U13568 ( .A(n15480), .B(n12392), .ZN(n11149) );
  XNOR2_X1 U13569 ( .A(n11149), .B(n11314), .ZN(n11008) );
  INV_X1 U13570 ( .A(n11002), .ZN(n11003) );
  NAND2_X1 U13571 ( .A1(n12739), .A2(n11003), .ZN(n11004) );
  NAND2_X1 U13572 ( .A1(n11005), .A2(n11004), .ZN(n11007) );
  INV_X1 U13573 ( .A(n11151), .ZN(n11006) );
  AOI21_X1 U13574 ( .B1(n11008), .B2(n11007), .A(n11006), .ZN(n11014) );
  INV_X1 U13575 ( .A(n11009), .ZN(n11396) );
  INV_X1 U13576 ( .A(n12491), .ZN(n12509) );
  NAND2_X1 U13577 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(P3_U3151), .ZN(n15411) );
  OAI21_X1 U13578 ( .B1(n12509), .B2(n11010), .A(n15411), .ZN(n11012) );
  OAI22_X1 U13579 ( .A1(n15451), .A2(n12500), .B1(n11437), .B2(n12489), .ZN(
        n11011) );
  AOI211_X1 U13580 ( .C1(n11396), .C2(n12486), .A(n11012), .B(n11011), .ZN(
        n11013) );
  OAI21_X1 U13581 ( .B1(n11014), .B2(n12494), .A(n11013), .ZN(P3_U3170) );
  INV_X1 U13582 ( .A(n11015), .ZN(n11028) );
  INV_X1 U13583 ( .A(n12529), .ZN(n11017) );
  NAND3_X1 U13584 ( .A1(n11017), .A2(n11016), .A3(n12392), .ZN(n11018) );
  OAI211_X1 U13585 ( .C1(n11020), .C2(n11366), .A(n11019), .B(n11018), .ZN(
        n11021) );
  NAND2_X1 U13586 ( .A1(n11021), .A2(n12496), .ZN(n11026) );
  INV_X1 U13587 ( .A(n12741), .ZN(n11022) );
  OAI22_X1 U13588 ( .A1(n11023), .A2(n12509), .B1(n11022), .B2(n12500), .ZN(
        n11024) );
  AOI21_X1 U13589 ( .B1(n12506), .B2(n10781), .A(n11024), .ZN(n11025) );
  OAI211_X1 U13590 ( .C1(n11028), .C2(n11027), .A(n11026), .B(n11025), .ZN(
        P3_U3162) );
  NAND2_X1 U13591 ( .A1(n6623), .A2(n11029), .ZN(n11030) );
  OAI21_X1 U13592 ( .B1(n6623), .B2(n9669), .A(n11030), .ZN(P2_U3559) );
  NAND2_X1 U13593 ( .A1(n11031), .A2(n14539), .ZN(n11037) );
  INV_X1 U13594 ( .A(n14557), .ZN(n15090) );
  OAI22_X1 U13595 ( .A1(n14539), .A2(n11032), .B1(P1_REG3_REG_3__SCAN_IN), 
        .B2(n14602), .ZN(n11034) );
  NOR2_X1 U13596 ( .A1(n14570), .A2(n13983), .ZN(n11033) );
  AOI211_X1 U13597 ( .C1(n11035), .C2(n15090), .A(n11034), .B(n11033), .ZN(
        n11036) );
  OAI211_X1 U13598 ( .C1(n11038), .C2(n15082), .A(n11037), .B(n11036), .ZN(
        P1_U3290) );
  XNOR2_X1 U13599 ( .A(n11039), .B(n14174), .ZN(n15126) );
  OAI211_X1 U13600 ( .C1(n11040), .C2(n15123), .A(n15086), .B(n15084), .ZN(
        n15122) );
  INV_X1 U13601 ( .A(n14602), .ZN(n15102) );
  AOI22_X1 U13602 ( .A1(n15081), .A2(n13999), .B1(n11195), .B2(n15102), .ZN(
        n11041) );
  OAI21_X1 U13603 ( .B1(n14557), .B2(n15122), .A(n11041), .ZN(n11048) );
  XNOR2_X1 U13604 ( .A(n11043), .B(n11042), .ZN(n11044) );
  NAND2_X1 U13605 ( .A1(n11044), .A2(n14952), .ZN(n11046) );
  AOI22_X1 U13606 ( .A1(n14921), .A2(n6624), .B1(n14226), .B2(n14583), .ZN(
        n11045) );
  NAND2_X1 U13607 ( .A1(n11046), .A2(n11045), .ZN(n15124) );
  MUX2_X1 U13608 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n15124), .S(n14539), .Z(
        n11047) );
  AOI211_X1 U13609 ( .C1(n15126), .C2(n14609), .A(n11048), .B(n11047), .ZN(
        n11049) );
  INV_X1 U13610 ( .A(n11049), .ZN(P1_U3288) );
  OR2_X1 U13611 ( .A1(n11051), .A2(n11050), .ZN(n11053) );
  NAND2_X1 U13612 ( .A1(n11053), .A2(n11052), .ZN(n15113) );
  NAND2_X1 U13613 ( .A1(n15113), .A2(n15162), .ZN(n11061) );
  OAI21_X1 U13614 ( .B1(n11055), .B2(n14168), .A(n11054), .ZN(n11059) );
  NAND2_X1 U13615 ( .A1(n14231), .A2(n14921), .ZN(n11057) );
  NAND2_X1 U13616 ( .A1(n14229), .A2(n14583), .ZN(n11056) );
  NAND2_X1 U13617 ( .A1(n11057), .A2(n11056), .ZN(n11058) );
  AOI21_X1 U13618 ( .B1(n11059), .B2(n14952), .A(n11058), .ZN(n11060) );
  AND2_X1 U13619 ( .A1(n11061), .A2(n11060), .ZN(n15115) );
  OAI22_X1 U13620 ( .A1(n14539), .A2(n9927), .B1(n11062), .B2(n14602), .ZN(
        n11067) );
  INV_X1 U13621 ( .A(n15113), .ZN(n11065) );
  OAI211_X1 U13622 ( .C1(n11064), .C2(n15111), .A(n15086), .B(n11063), .ZN(
        n15110) );
  OAI22_X1 U13623 ( .A1(n11065), .A2(n15082), .B1(n14557), .B2(n15110), .ZN(
        n11066) );
  AOI211_X1 U13624 ( .C1(n15081), .C2(n13978), .A(n11067), .B(n11066), .ZN(
        n11068) );
  OAI21_X1 U13625 ( .B1(n15105), .B2(n15115), .A(n11068), .ZN(P1_U3291) );
  INV_X1 U13626 ( .A(n11069), .ZN(n11167) );
  AOI22_X1 U13627 ( .A1(n14322), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n11286), .ZN(n11070) );
  OAI21_X1 U13628 ( .B1(n11167), .B2(n14761), .A(n11070), .ZN(P1_U3340) );
  MUX2_X1 U13629 ( .A(P3_REG2_REG_9__SCAN_IN), .B(P3_REG1_REG_9__SCAN_IN), .S(
        n13165), .Z(n11670) );
  XOR2_X1 U13630 ( .A(n11659), .B(n11670), .Z(n11671) );
  INV_X1 U13631 ( .A(n11071), .ZN(n11072) );
  XOR2_X1 U13632 ( .A(n11671), .B(n11672), .Z(n11088) );
  OAI21_X1 U13633 ( .B1(n11077), .B2(P3_REG1_REG_9__SCAN_IN), .A(n11658), .ZN(
        n11086) );
  NAND2_X1 U13634 ( .A1(P3_REG2_REG_9__SCAN_IN), .A2(n11081), .ZN(n11649) );
  OAI21_X1 U13635 ( .B1(n11081), .B2(P3_REG2_REG_9__SCAN_IN), .A(n11649), .ZN(
        n11082) );
  NAND2_X1 U13636 ( .A1(n11082), .A2(n15429), .ZN(n11084) );
  AND2_X1 U13637 ( .A1(P3_U3151), .A2(P3_REG3_REG_9__SCAN_IN), .ZN(n11796) );
  AOI21_X1 U13638 ( .B1(n15415), .B2(P3_ADDR_REG_9__SCAN_IN), .A(n11796), .ZN(
        n11083) );
  OAI211_X1 U13639 ( .C1(n11925), .C2(n11669), .A(n11084), .B(n11083), .ZN(
        n11085) );
  AOI21_X1 U13640 ( .B1(n11086), .B2(n15426), .A(n11085), .ZN(n11087) );
  OAI21_X1 U13641 ( .B1(n11088), .B2(n15406), .A(n11087), .ZN(P3_U3191) );
  XNOR2_X1 U13642 ( .A(n15323), .B(n13255), .ZN(n11339) );
  NAND2_X1 U13643 ( .A1(n13651), .A2(n13377), .ZN(n11337) );
  XNOR2_X1 U13644 ( .A(n11339), .B(n11337), .ZN(n11335) );
  XNOR2_X1 U13645 ( .A(n11093), .B(n11335), .ZN(n11098) );
  INV_X1 U13646 ( .A(n15327), .ZN(n11094) );
  OAI22_X1 U13647 ( .A1(n15198), .A2(n11094), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8468), .ZN(n11096) );
  AOI22_X1 U13648 ( .A1(n13337), .A2(n13378), .B1(n13336), .B2(n13376), .ZN(
        n11260) );
  NOR2_X1 U13649 ( .A1(n13347), .A2(n11260), .ZN(n11095) );
  AOI211_X1 U13650 ( .C1(n15323), .C2(n15195), .A(n11096), .B(n11095), .ZN(
        n11097) );
  OAI21_X1 U13651 ( .B1(n11098), .B2(n13349), .A(n11097), .ZN(P2_U3185) );
  MUX2_X1 U13652 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n11100), .S(n11276), .Z(
        n11101) );
  NAND2_X1 U13653 ( .A1(n11102), .A2(n11101), .ZN(n11271) );
  OAI21_X1 U13654 ( .B1(n11102), .B2(n11101), .A(n11271), .ZN(n11111) );
  AOI21_X1 U13655 ( .B1(P1_REG2_REG_10__SCAN_IN), .B2(n11104), .A(n11103), 
        .ZN(n11106) );
  MUX2_X1 U13656 ( .A(n10180), .B(P1_REG2_REG_11__SCAN_IN), .S(n11276), .Z(
        n11105) );
  NOR2_X1 U13657 ( .A1(n11106), .A2(n11105), .ZN(n11275) );
  AOI211_X1 U13658 ( .C1(n11106), .C2(n11105), .A(n15060), .B(n11275), .ZN(
        n11110) );
  NAND2_X1 U13659 ( .A1(n15067), .A2(n11276), .ZN(n11107) );
  NAND2_X1 U13660 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n14911)
         );
  OAI211_X1 U13661 ( .C1(n11108), .C2(n15070), .A(n11107), .B(n14911), .ZN(
        n11109) );
  AOI211_X1 U13662 ( .C1(n11111), .C2(n15015), .A(n11110), .B(n11109), .ZN(
        n11112) );
  INV_X1 U13663 ( .A(n11112), .ZN(P1_U3254) );
  OAI21_X1 U13664 ( .B1(n11114), .B2(n11118), .A(n11113), .ZN(n11138) );
  INV_X1 U13665 ( .A(n11115), .ZN(n11117) );
  INV_X1 U13666 ( .A(n11257), .ZN(n11116) );
  AOI211_X1 U13667 ( .C1(n11123), .C2(n11117), .A(n13651), .B(n11116), .ZN(
        n11145) );
  XNOR2_X1 U13668 ( .A(n11119), .B(n11118), .ZN(n11122) );
  INV_X1 U13669 ( .A(n11120), .ZN(n11121) );
  OAI21_X1 U13670 ( .B1(n11122), .B2(n13623), .A(n11121), .ZN(n11139) );
  AOI211_X1 U13671 ( .C1(n15381), .C2(n11138), .A(n11145), .B(n11139), .ZN(
        n11127) );
  AOI22_X1 U13672 ( .A1(n12144), .A2(n11123), .B1(n15389), .B2(
        P2_REG1_REG_6__SCAN_IN), .ZN(n11124) );
  OAI21_X1 U13673 ( .B1(n11127), .B2(n15389), .A(n11124), .ZN(P2_U3505) );
  OAI22_X1 U13674 ( .A1(n13783), .A2(n11143), .B1(n15383), .B2(n8457), .ZN(
        n11125) );
  INV_X1 U13675 ( .A(n11125), .ZN(n11126) );
  OAI21_X1 U13676 ( .B1(n11127), .B2(n15382), .A(n11126), .ZN(P2_U3448) );
  INV_X1 U13677 ( .A(n11128), .ZN(n11129) );
  OAI22_X1 U13678 ( .A1(n15330), .A2(n11130), .B1(n13655), .B2(n11129), .ZN(
        n11131) );
  AOI21_X1 U13679 ( .B1(n15324), .B2(n11132), .A(n11131), .ZN(n11136) );
  MUX2_X1 U13680 ( .A(n11134), .B(n11133), .S(n6620), .Z(n11135) );
  OAI211_X1 U13681 ( .C1(n13592), .C2(n11137), .A(n11136), .B(n11135), .ZN(
        P2_U3261) );
  INV_X1 U13682 ( .A(n11138), .ZN(n11148) );
  INV_X1 U13683 ( .A(n11139), .ZN(n11140) );
  MUX2_X1 U13684 ( .A(n11141), .B(n11140), .S(n13643), .Z(n11147) );
  OAI22_X1 U13685 ( .A1(n15330), .A2(n11143), .B1(n13655), .B2(n11142), .ZN(
        n11144) );
  AOI21_X1 U13686 ( .B1(n15324), .B2(n11145), .A(n11144), .ZN(n11146) );
  OAI211_X1 U13687 ( .C1(n11148), .C2(n13592), .A(n11147), .B(n11146), .ZN(
        P2_U3259) );
  NAND2_X1 U13688 ( .A1(n11149), .A2(n11314), .ZN(n11150) );
  XNOR2_X1 U13689 ( .A(n11155), .B(n12360), .ZN(n11436) );
  XNOR2_X1 U13690 ( .A(n11436), .B(n11437), .ZN(n11434) );
  XNOR2_X1 U13691 ( .A(n11435), .B(n11434), .ZN(n11152) );
  NAND2_X1 U13692 ( .A1(n11152), .A2(n12496), .ZN(n11157) );
  OAI22_X1 U13693 ( .A1(n11314), .A2(n12500), .B1(n11444), .B2(n12489), .ZN(
        n11153) );
  AOI211_X1 U13694 ( .C1(n11155), .C2(n12491), .A(n11154), .B(n11153), .ZN(
        n11156) );
  OAI211_X1 U13695 ( .C1(n11534), .C2(n12503), .A(n11157), .B(n11156), .ZN(
        P3_U3167) );
  XNOR2_X1 U13696 ( .A(n11158), .B(n14176), .ZN(n15143) );
  XNOR2_X1 U13697 ( .A(n11159), .B(n14176), .ZN(n11160) );
  AOI22_X1 U13698 ( .A1(n14921), .A2(n14226), .B1(n14224), .B2(n14583), .ZN(
        n11552) );
  OAI21_X1 U13699 ( .B1(n11160), .B2(n15075), .A(n11552), .ZN(n15139) );
  INV_X1 U13700 ( .A(n15139), .ZN(n11161) );
  MUX2_X1 U13701 ( .A(n11162), .B(n11161), .S(n14539), .Z(n11166) );
  XNOR2_X1 U13702 ( .A(n11557), .B(n15085), .ZN(n11163) );
  NOR2_X1 U13703 ( .A1(n11163), .A2(n14915), .ZN(n15140) );
  OAI22_X1 U13704 ( .A1(n11557), .A2(n14570), .B1(n11550), .B2(n14602), .ZN(
        n11164) );
  AOI21_X1 U13705 ( .B1(n15140), .B2(n15090), .A(n11164), .ZN(n11165) );
  OAI211_X1 U13706 ( .C1(n15099), .C2(n15143), .A(n11166), .B(n11165), .ZN(
        P1_U3286) );
  INV_X1 U13707 ( .A(n11604), .ZN(n11596) );
  OAI222_X1 U13708 ( .A1(n13798), .A2(n11168), .B1(n13804), .B2(n11167), .C1(
        P2_U3088), .C2(n11596), .ZN(P2_U3312) );
  NAND2_X1 U13709 ( .A1(n12740), .A2(P3_DATAO_REG_27__SCAN_IN), .ZN(n11169) );
  OAI21_X1 U13710 ( .B1(n12891), .B2(n12740), .A(n11169), .ZN(P3_U3518) );
  OAI22_X1 U13711 ( .A1(n13983), .A2(n11299), .B1(n12284), .B2(n13985), .ZN(
        n11174) );
  OAI22_X1 U13712 ( .A1(n13983), .A2(n12256), .B1(n13985), .B2(n11299), .ZN(
        n11173) );
  XNOR2_X1 U13713 ( .A(n11173), .B(n12208), .ZN(n11175) );
  XOR2_X1 U13714 ( .A(n11174), .B(n11175), .Z(n13825) );
  NAND2_X1 U13715 ( .A1(n13826), .A2(n13825), .ZN(n13824) );
  NAND2_X1 U13716 ( .A1(n11175), .A2(n11174), .ZN(n11179) );
  NAND2_X1 U13717 ( .A1(n13990), .A2(n6622), .ZN(n11177) );
  NAND2_X1 U13718 ( .A1(n12301), .A2(n6624), .ZN(n11176) );
  AND2_X1 U13719 ( .A1(n11177), .A2(n11176), .ZN(n11180) );
  OAI22_X1 U13720 ( .A1(n15117), .A2(n12256), .B1(n11192), .B2(n11299), .ZN(
        n11178) );
  XNOR2_X1 U13721 ( .A(n11178), .B(n12208), .ZN(n11209) );
  NAND3_X1 U13722 ( .A1(n13824), .A2(n11180), .A3(n11179), .ZN(n11206) );
  NAND2_X1 U13723 ( .A1(n13999), .A2(n12300), .ZN(n11182) );
  NAND2_X1 U13724 ( .A1(n14227), .A2(n6622), .ZN(n11181) );
  NAND2_X1 U13725 ( .A1(n11182), .A2(n11181), .ZN(n11183) );
  XNOR2_X1 U13726 ( .A(n11183), .B(n12208), .ZN(n11187) );
  NAND2_X1 U13727 ( .A1(n13999), .A2(n6622), .ZN(n11185) );
  NAND2_X1 U13728 ( .A1(n12301), .A2(n14227), .ZN(n11184) );
  NAND2_X1 U13729 ( .A1(n11185), .A2(n11184), .ZN(n11186) );
  NOR2_X1 U13730 ( .A1(n11187), .A2(n11186), .ZN(n11294) );
  INV_X1 U13731 ( .A(n11294), .ZN(n11188) );
  NAND2_X1 U13732 ( .A1(n11187), .A2(n11186), .ZN(n11293) );
  NAND2_X1 U13733 ( .A1(n11188), .A2(n11293), .ZN(n11189) );
  XNOR2_X1 U13734 ( .A(n11295), .B(n11189), .ZN(n11197) );
  INV_X1 U13735 ( .A(n14914), .ZN(n13918) );
  NAND2_X1 U13736 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n14263) );
  OAI21_X1 U13737 ( .B1(n14897), .B2(n11191), .A(n14263), .ZN(n11194) );
  INV_X1 U13738 ( .A(n13943), .ZN(n14900) );
  OAI22_X1 U13739 ( .A1(n14900), .A2(n11192), .B1(n13922), .B2(n15123), .ZN(
        n11193) );
  AOI211_X1 U13740 ( .C1(n11195), .C2(n13918), .A(n11194), .B(n11193), .ZN(
        n11196) );
  OAI21_X1 U13741 ( .B1(n11197), .B2(n14904), .A(n11196), .ZN(P1_U3227) );
  NAND2_X1 U13742 ( .A1(n6620), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n11198) );
  OAI21_X1 U13743 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(n13655), .A(n11198), .ZN(
        n11202) );
  OAI22_X1 U13744 ( .A1(n13612), .A2(n11200), .B1(n13592), .B2(n11199), .ZN(
        n11201) );
  AOI211_X1 U13745 ( .C1(n13641), .C2(n11203), .A(n11202), .B(n11201), .ZN(
        n11204) );
  OAI21_X1 U13746 ( .B1(n6620), .B2(n11205), .A(n11204), .ZN(P2_U3262) );
  INV_X1 U13747 ( .A(n11206), .ZN(n11208) );
  NOR2_X1 U13748 ( .A1(n11208), .A2(n11207), .ZN(n11210) );
  XNOR2_X1 U13749 ( .A(n11210), .B(n11209), .ZN(n11218) );
  INV_X1 U13750 ( .A(n11211), .ZN(n11216) );
  OAI21_X1 U13751 ( .B1(n14897), .B2(n11213), .A(n11212), .ZN(n11215) );
  OAI22_X1 U13752 ( .A1(n14900), .A2(n13985), .B1(n13922), .B2(n15117), .ZN(
        n11214) );
  AOI211_X1 U13753 ( .C1(n11216), .C2(n13918), .A(n11215), .B(n11214), .ZN(
        n11217) );
  OAI21_X1 U13754 ( .B1(n11218), .B2(n14904), .A(n11217), .ZN(P1_U3230) );
  XNOR2_X1 U13755 ( .A(n11219), .B(n11222), .ZN(n15151) );
  OAI211_X1 U13756 ( .C1(n6920), .C2(n6764), .A(n15086), .B(n14610), .ZN(
        n15148) );
  NOR2_X1 U13757 ( .A1(n15148), .A2(n14557), .ZN(n11221) );
  OAI22_X1 U13758 ( .A1(n6920), .A2(n14570), .B1(n14602), .B2(n11727), .ZN(
        n11220) );
  AOI211_X1 U13759 ( .C1(n15151), .C2(n14609), .A(n11221), .B(n11220), .ZN(
        n11232) );
  AOI21_X1 U13760 ( .B1(n11223), .B2(n11222), .A(n15075), .ZN(n11225) );
  AND2_X1 U13761 ( .A1(n11225), .A2(n11224), .ZN(n15149) );
  NAND2_X1 U13762 ( .A1(n14225), .A2(n14921), .ZN(n11227) );
  NAND2_X1 U13763 ( .A1(n14223), .A2(n14583), .ZN(n11226) );
  AND2_X1 U13764 ( .A1(n11227), .A2(n11226), .ZN(n15147) );
  INV_X1 U13765 ( .A(n15147), .ZN(n11228) );
  NOR2_X1 U13766 ( .A1(n15149), .A2(n11228), .ZN(n11229) );
  MUX2_X1 U13767 ( .A(n11230), .B(n11229), .S(n14539), .Z(n11231) );
  NAND2_X1 U13768 ( .A1(n11232), .A2(n11231), .ZN(P1_U3285) );
  NAND2_X1 U13769 ( .A1(n12740), .A2(P3_DATAO_REG_28__SCAN_IN), .ZN(n11233) );
  OAI21_X1 U13770 ( .B1(n12877), .B2(n12740), .A(n11233), .ZN(P3_U3519) );
  NAND2_X1 U13771 ( .A1(n14125), .A2(n14232), .ZN(n11234) );
  OAI21_X1 U13772 ( .B1(n8218), .B2(P1_U4016), .A(n11234), .ZN(P1_U3588) );
  OAI22_X1 U13773 ( .A1(n13092), .A2(n11527), .B1(n15498), .B2(n10513), .ZN(
        n11235) );
  AOI21_X1 U13774 ( .B1(n11525), .B2(n15498), .A(n11235), .ZN(n11236) );
  INV_X1 U13775 ( .A(n11236), .ZN(P3_U3459) );
  INV_X1 U13776 ( .A(n11237), .ZN(n11268) );
  INV_X1 U13777 ( .A(n14316), .ZN(n15036) );
  INV_X1 U13778 ( .A(n11239), .ZN(n11241) );
  OAI222_X1 U13779 ( .A1(P3_U3151), .A2(n11242), .B1(n13172), .B2(n11241), 
        .C1(n11240), .C2(n13167), .ZN(P3_U3275) );
  INV_X1 U13780 ( .A(n13092), .ZN(n11686) );
  AOI22_X1 U13781 ( .A1(n11686), .A2(n11479), .B1(n6791), .B2(
        P3_REG1_REG_3__SCAN_IN), .ZN(n11243) );
  OAI21_X1 U13782 ( .B1(n11244), .B2(n6791), .A(n11243), .ZN(P3_U3462) );
  INV_X1 U13783 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n11253) );
  INV_X1 U13784 ( .A(P3_REG1_REG_31__SCAN_IN), .ZN(n11248) );
  NAND2_X1 U13785 ( .A1(n11245), .A2(P3_REG2_REG_31__SCAN_IN), .ZN(n11247) );
  NAND2_X1 U13786 ( .A1(n9256), .A2(P3_REG0_REG_31__SCAN_IN), .ZN(n11246) );
  OAI211_X1 U13787 ( .C1(n9270), .C2(n11248), .A(n11247), .B(n11246), .ZN(
        n11249) );
  INV_X1 U13788 ( .A(n11249), .ZN(n11250) );
  NAND2_X1 U13789 ( .A1(n11251), .A2(n11250), .ZN(n12851) );
  NAND2_X1 U13790 ( .A1(n12851), .A2(P3_U3897), .ZN(n11252) );
  OAI21_X1 U13791 ( .B1(P3_U3897), .B2(n11253), .A(n11252), .ZN(P3_U3522) );
  OAI21_X1 U13792 ( .B1(n11255), .B2(n11259), .A(n11254), .ZN(n15334) );
  INV_X1 U13793 ( .A(n11462), .ZN(n11256) );
  AOI211_X1 U13794 ( .C1(n15323), .C2(n11257), .A(n13651), .B(n11256), .ZN(
        n15325) );
  XOR2_X1 U13795 ( .A(n11258), .B(n11259), .Z(n11262) );
  INV_X1 U13796 ( .A(n11260), .ZN(n11261) );
  AOI21_X1 U13797 ( .B1(n11262), .B2(n13661), .A(n11261), .ZN(n15336) );
  INV_X1 U13798 ( .A(n15336), .ZN(n11263) );
  AOI211_X1 U13799 ( .C1(n15381), .C2(n15334), .A(n15325), .B(n11263), .ZN(
        n11267) );
  INV_X1 U13800 ( .A(n13783), .ZN(n12147) );
  NOR2_X1 U13801 ( .A1(n15383), .A2(n8471), .ZN(n11264) );
  AOI21_X1 U13802 ( .B1(n12147), .B2(n15323), .A(n11264), .ZN(n11265) );
  OAI21_X1 U13803 ( .B1(n11267), .B2(n15382), .A(n11265), .ZN(P2_U3451) );
  AOI22_X1 U13804 ( .A1(n12144), .A2(n15323), .B1(n15389), .B2(
        P2_REG1_REG_7__SCAN_IN), .ZN(n11266) );
  OAI21_X1 U13805 ( .B1(n11267), .B2(n15389), .A(n11266), .ZN(P2_U3506) );
  OAI222_X1 U13806 ( .A1(n13798), .A2(n11269), .B1(n11880), .B2(P2_U3088), 
        .C1(n13804), .C2(n11268), .ZN(P2_U3311) );
  INV_X1 U13807 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n11270) );
  MUX2_X1 U13808 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n11270), .S(n14319), .Z(
        n11273) );
  NAND2_X1 U13809 ( .A1(n11272), .A2(n11273), .ZN(n14318) );
  OAI21_X1 U13810 ( .B1(n11273), .B2(n11272), .A(n14318), .ZN(n11274) );
  NAND2_X1 U13811 ( .A1(n11274), .A2(n15015), .ZN(n11284) );
  AOI21_X1 U13812 ( .B1(n11276), .B2(P1_REG2_REG_11__SCAN_IN), .A(n11275), 
        .ZN(n11278) );
  MUX2_X1 U13813 ( .A(P1_REG2_REG_12__SCAN_IN), .B(n11848), .S(n14319), .Z(
        n11277) );
  NAND2_X1 U13814 ( .A1(n11278), .A2(n11277), .ZN(n14303) );
  OAI21_X1 U13815 ( .B1(n11278), .B2(n11277), .A(n14303), .ZN(n11282) );
  INV_X1 U13816 ( .A(n14319), .ZN(n11280) );
  NAND2_X1 U13817 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n13853)
         );
  NAND2_X1 U13818 ( .A1(n14981), .A2(P1_ADDR_REG_12__SCAN_IN), .ZN(n11279) );
  OAI211_X1 U13819 ( .C1(n15037), .C2(n11280), .A(n13853), .B(n11279), .ZN(
        n11281) );
  AOI21_X1 U13820 ( .B1(n11282), .B2(n15012), .A(n11281), .ZN(n11283) );
  NAND2_X1 U13821 ( .A1(n11284), .A2(n11283), .ZN(P1_U3255) );
  INV_X1 U13822 ( .A(n11285), .ZN(n11292) );
  AOI22_X1 U13823 ( .A1(n15052), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n11286), .ZN(n11287) );
  OAI21_X1 U13824 ( .B1(n11292), .B2(n14761), .A(n11287), .ZN(P1_U3338) );
  INV_X1 U13825 ( .A(n12859), .ZN(n11288) );
  NAND2_X1 U13826 ( .A1(n11288), .A2(P3_U3897), .ZN(n11289) );
  OAI21_X1 U13827 ( .B1(P3_U3897), .B2(n11290), .A(n11289), .ZN(P3_U3520) );
  INV_X1 U13828 ( .A(n13407), .ZN(n13404) );
  OAI222_X1 U13829 ( .A1(n13804), .A2(n11292), .B1(n13404), .B2(P2_U3088), 
        .C1(n11291), .C2(n13798), .ZN(P2_U3310) );
  NAND2_X1 U13830 ( .A1(n15083), .A2(n12300), .ZN(n11297) );
  NAND2_X1 U13831 ( .A1(n14226), .A2(n6622), .ZN(n11296) );
  NAND2_X1 U13832 ( .A1(n11297), .A2(n11296), .ZN(n11298) );
  XNOR2_X1 U13833 ( .A(n11298), .B(n12208), .ZN(n11541) );
  AOI22_X1 U13834 ( .A1(n15083), .A2(n6622), .B1(n12301), .B2(n14226), .ZN(
        n11543) );
  XNOR2_X1 U13835 ( .A(n11541), .B(n11543), .ZN(n11300) );
  NAND2_X1 U13836 ( .A1(n11301), .A2(n11300), .ZN(n11542) );
  INV_X1 U13837 ( .A(n14904), .ZN(n13912) );
  OAI211_X1 U13838 ( .C1(n11301), .C2(n11300), .A(n11542), .B(n13912), .ZN(
        n11307) );
  NAND2_X1 U13839 ( .A1(n14227), .A2(n14921), .ZN(n11303) );
  NAND2_X1 U13840 ( .A1(n14225), .A2(n14583), .ZN(n11302) );
  NAND2_X1 U13841 ( .A1(n11303), .A2(n11302), .ZN(n15078) );
  AOI22_X1 U13842 ( .A1(n13934), .A2(n15078), .B1(P1_REG3_REG_6__SCAN_IN), 
        .B2(P1_U3086), .ZN(n11304) );
  OAI21_X1 U13843 ( .B1(n15079), .B2(n14914), .A(n11304), .ZN(n11305) );
  AOI21_X1 U13844 ( .B1(n15083), .B2(n14909), .A(n11305), .ZN(n11306) );
  NAND2_X1 U13845 ( .A1(n11307), .A2(n11306), .ZN(P1_U3239) );
  OAI21_X1 U13846 ( .B1(n11309), .B2(n12672), .A(n11308), .ZN(n11539) );
  INV_X1 U13847 ( .A(n11310), .ZN(n11311) );
  AOI21_X1 U13848 ( .B1(n12672), .B2(n11312), .A(n11311), .ZN(n11313) );
  OAI222_X1 U13849 ( .A1(n15450), .A2(n11444), .B1(n15452), .B2(n11314), .C1(
        n15457), .C2(n11313), .ZN(n11536) );
  AOI21_X1 U13850 ( .B1(n15477), .B2(n11539), .A(n11536), .ZN(n11320) );
  INV_X1 U13851 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n11315) );
  OAI22_X1 U13852 ( .A1(n11535), .A2(n13144), .B1(n15493), .B2(n11315), .ZN(
        n11316) );
  INV_X1 U13853 ( .A(n11316), .ZN(n11317) );
  OAI21_X1 U13854 ( .B1(n11320), .B2(n15491), .A(n11317), .ZN(P3_U3405) );
  OAI22_X1 U13855 ( .A1(n13092), .A2(n11535), .B1(n15498), .B2(n10868), .ZN(
        n11318) );
  INV_X1 U13856 ( .A(n11318), .ZN(n11319) );
  OAI21_X1 U13857 ( .B1(n11320), .B2(n6791), .A(n11319), .ZN(P3_U3464) );
  INV_X1 U13858 ( .A(n11321), .ZN(n11324) );
  OAI222_X1 U13859 ( .A1(n13172), .A2(n11324), .B1(n13167), .B2(n11323), .C1(
        P3_U3151), .C2(n11322), .ZN(P3_U3274) );
  INV_X1 U13860 ( .A(n11325), .ZN(n11334) );
  NAND2_X1 U13861 ( .A1(n15324), .A2(n11326), .ZN(n11329) );
  AOI22_X1 U13862 ( .A1(n6620), .A2(P2_REG2_REG_5__SCAN_IN), .B1(n11327), .B2(
        n15326), .ZN(n11328) );
  OAI211_X1 U13863 ( .C1(n11330), .C2(n15330), .A(n11329), .B(n11328), .ZN(
        n11331) );
  AOI21_X1 U13864 ( .B1(n15333), .B2(n11332), .A(n11331), .ZN(n11333) );
  OAI21_X1 U13865 ( .B1(n6620), .B2(n11334), .A(n11333), .ZN(P2_U3260) );
  INV_X1 U13866 ( .A(n11337), .ZN(n11338) );
  NAND2_X1 U13867 ( .A1(n11339), .A2(n11338), .ZN(n11340) );
  XNOR2_X1 U13868 ( .A(n15364), .B(n13213), .ZN(n11341) );
  NAND2_X1 U13869 ( .A1(n13651), .A2(n13376), .ZN(n11342) );
  NAND2_X1 U13870 ( .A1(n11341), .A2(n11342), .ZN(n11420) );
  INV_X1 U13871 ( .A(n11341), .ZN(n11344) );
  INV_X1 U13872 ( .A(n11342), .ZN(n11343) );
  NAND2_X1 U13873 ( .A1(n11344), .A2(n11343), .ZN(n11345) );
  NAND2_X1 U13874 ( .A1(n11420), .A2(n11345), .ZN(n11348) );
  INV_X1 U13875 ( .A(n11421), .ZN(n11347) );
  AOI21_X1 U13876 ( .B1(n11349), .B2(n11348), .A(n11347), .ZN(n11356) );
  NAND2_X1 U13877 ( .A1(n13336), .A2(n13375), .ZN(n11351) );
  NAND2_X1 U13878 ( .A1(n13337), .A2(n13377), .ZN(n11350) );
  NAND2_X1 U13879 ( .A1(n11351), .A2(n11350), .ZN(n11456) );
  NAND2_X1 U13880 ( .A1(n15190), .A2(n11456), .ZN(n11353) );
  OAI211_X1 U13881 ( .C1(n15198), .C2(n11460), .A(n11353), .B(n11352), .ZN(
        n11354) );
  AOI21_X1 U13882 ( .B1(n15364), .B2(n15195), .A(n11354), .ZN(n11355) );
  OAI21_X1 U13883 ( .B1(n11356), .B2(n13349), .A(n11355), .ZN(P2_U3193) );
  INV_X1 U13884 ( .A(n11360), .ZN(n11357) );
  NAND2_X1 U13885 ( .A1(n11358), .A2(n11357), .ZN(n11363) );
  INV_X1 U13886 ( .A(n11359), .ZN(n11361) );
  OAI21_X1 U13887 ( .B1(n13150), .B2(n11361), .A(n11360), .ZN(n11362) );
  XNOR2_X1 U13888 ( .A(n12529), .B(n11016), .ZN(n11372) );
  INV_X1 U13889 ( .A(n15454), .ZN(n12944) );
  AOI22_X1 U13890 ( .A1(n10781), .A2(n13029), .B1(n13027), .B2(n12741), .ZN(
        n11369) );
  XNOR2_X1 U13891 ( .A(n11366), .B(n11016), .ZN(n11367) );
  NAND2_X1 U13892 ( .A1(n11367), .A2(n13032), .ZN(n11368) );
  OAI211_X1 U13893 ( .C1(n11372), .C2(n12944), .A(n11369), .B(n11368), .ZN(
        n15468) );
  NAND2_X1 U13894 ( .A1(n11370), .A2(n15479), .ZN(n15467) );
  OAI22_X1 U13895 ( .A1(n15467), .A2(n12705), .B1(n11027), .B2(n15440), .ZN(
        n11371) );
  OAI21_X1 U13896 ( .B1(n15468), .B2(n11371), .A(n15464), .ZN(n11374) );
  INV_X1 U13897 ( .A(n11372), .ZN(n15470) );
  AND2_X1 U13898 ( .A1(n12528), .A2(n12705), .ZN(n15460) );
  NAND2_X1 U13899 ( .A1(n15470), .A2(n12927), .ZN(n11373) );
  OAI211_X1 U13900 ( .C1(n10510), .C2(n15464), .A(n11374), .B(n11373), .ZN(
        P3_U3232) );
  OAI21_X1 U13901 ( .B1(n11377), .B2(n11376), .A(n11375), .ZN(n15436) );
  OAI211_X1 U13902 ( .C1(n6767), .C2(n12676), .A(n11378), .B(n13032), .ZN(
        n11380) );
  NAND2_X1 U13903 ( .A1(n12737), .A2(n13027), .ZN(n11379) );
  OAI211_X1 U13904 ( .C1(n11622), .C2(n15450), .A(n11380), .B(n11379), .ZN(
        n15435) );
  AOI21_X1 U13905 ( .B1(n15477), .B2(n15436), .A(n15435), .ZN(n11385) );
  AOI22_X1 U13906 ( .A1(n11686), .A2(n11516), .B1(n6791), .B2(
        P3_REG1_REG_6__SCAN_IN), .ZN(n11381) );
  OAI21_X1 U13907 ( .B1(n11385), .B2(n6791), .A(n11381), .ZN(P3_U3465) );
  INV_X1 U13908 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n11382) );
  OAI22_X1 U13909 ( .A1(n15441), .A2(n13144), .B1(n15493), .B2(n11382), .ZN(
        n11383) );
  INV_X1 U13910 ( .A(n11383), .ZN(n11384) );
  OAI21_X1 U13911 ( .B1(n11385), .B2(n15491), .A(n11384), .ZN(P3_U3408) );
  XNOR2_X1 U13912 ( .A(n11386), .B(n12670), .ZN(n15478) );
  INV_X1 U13913 ( .A(n15478), .ZN(n11401) );
  OAI211_X1 U13914 ( .C1(n11389), .C2(n11388), .A(n11387), .B(n13032), .ZN(
        n11392) );
  OAI22_X1 U13915 ( .A1(n15451), .A2(n15452), .B1(n11437), .B2(n15450), .ZN(
        n11390) );
  INV_X1 U13916 ( .A(n11390), .ZN(n11391) );
  NAND2_X1 U13917 ( .A1(n11392), .A2(n11391), .ZN(n15483) );
  INV_X1 U13918 ( .A(n11393), .ZN(n11395) );
  NOR2_X1 U13919 ( .A1(n15486), .A2(n12705), .ZN(n11394) );
  INV_X1 U13920 ( .A(n15442), .ZN(n13008) );
  AOI22_X1 U13921 ( .A1(n13008), .A2(n15480), .B1(n15463), .B2(n11396), .ZN(
        n11397) );
  OAI21_X1 U13922 ( .B1(n11398), .B2(n15464), .A(n11397), .ZN(n11399) );
  AOI21_X1 U13923 ( .B1(n15483), .B2(n15464), .A(n11399), .ZN(n11400) );
  OAI21_X1 U13924 ( .B1(n12088), .B2(n11401), .A(n11400), .ZN(P3_U3229) );
  OAI21_X1 U13925 ( .B1(n11403), .B2(n12673), .A(n11402), .ZN(n11632) );
  OAI211_X1 U13926 ( .C1(n11405), .C2(n11442), .A(n11404), .B(n13032), .ZN(
        n11408) );
  OAI22_X1 U13927 ( .A1(n11444), .A2(n15452), .B1(n11794), .B2(n15450), .ZN(
        n11406) );
  INV_X1 U13928 ( .A(n11406), .ZN(n11407) );
  NAND2_X1 U13929 ( .A1(n11408), .A2(n11407), .ZN(n11629) );
  AOI21_X1 U13930 ( .B1(n15477), .B2(n11632), .A(n11629), .ZN(n11414) );
  INV_X1 U13931 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n11409) );
  OAI22_X1 U13932 ( .A1(n11628), .A2(n13144), .B1(n15493), .B2(n11409), .ZN(
        n11410) );
  INV_X1 U13933 ( .A(n11410), .ZN(n11411) );
  OAI21_X1 U13934 ( .B1(n11414), .B2(n15491), .A(n11411), .ZN(P3_U3411) );
  OAI22_X1 U13935 ( .A1(n13092), .A2(n11628), .B1(n15498), .B2(n9332), .ZN(
        n11412) );
  INV_X1 U13936 ( .A(n11412), .ZN(n11413) );
  OAI21_X1 U13937 ( .B1(n11414), .B2(n6791), .A(n11413), .ZN(P3_U3466) );
  XNOR2_X1 U13938 ( .A(n11746), .B(n13213), .ZN(n11415) );
  NAND2_X1 U13939 ( .A1(n13651), .A2(n13375), .ZN(n11416) );
  NAND2_X1 U13940 ( .A1(n11415), .A2(n11416), .ZN(n11483) );
  INV_X1 U13941 ( .A(n11415), .ZN(n11418) );
  INV_X1 U13942 ( .A(n11416), .ZN(n11417) );
  NAND2_X1 U13943 ( .A1(n11418), .A2(n11417), .ZN(n11419) );
  AND2_X1 U13944 ( .A1(n11483), .A2(n11419), .ZN(n11423) );
  NAND2_X1 U13945 ( .A1(n11421), .A2(n11420), .ZN(n11422) );
  OAI21_X1 U13946 ( .B1(n11423), .B2(n11422), .A(n11484), .ZN(n11424) );
  NAND2_X1 U13947 ( .A1(n11424), .A2(n15193), .ZN(n11429) );
  OAI22_X1 U13948 ( .A1(n11426), .A2(n13303), .B1(n11425), .B2(n13301), .ZN(
        n11561) );
  NAND2_X1 U13949 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3088), .ZN(n15255) );
  OAI21_X1 U13950 ( .B1(n15198), .B2(n11567), .A(n15255), .ZN(n11427) );
  AOI21_X1 U13951 ( .B1(n15190), .B2(n11561), .A(n11427), .ZN(n11428) );
  OAI211_X1 U13952 ( .C1(n11743), .C2(n13331), .A(n11429), .B(n11428), .ZN(
        P2_U3203) );
  INV_X1 U13953 ( .A(n11430), .ZN(n11432) );
  INV_X1 U13954 ( .A(n13415), .ZN(n13419) );
  OAI222_X1 U13955 ( .A1(n13798), .A2(n11433), .B1(n13804), .B2(n11432), .C1(
        P2_U3088), .C2(n13419), .ZN(P2_U3309) );
  INV_X1 U13956 ( .A(n11436), .ZN(n11438) );
  NAND2_X1 U13957 ( .A1(n11438), .A2(n11437), .ZN(n11439) );
  XNOR2_X1 U13958 ( .A(n11516), .B(n12392), .ZN(n11440) );
  XNOR2_X1 U13959 ( .A(n11440), .B(n11444), .ZN(n11520) );
  INV_X1 U13960 ( .A(n11440), .ZN(n11441) );
  XNOR2_X1 U13961 ( .A(n11442), .B(n6818), .ZN(n11572) );
  NAND2_X1 U13962 ( .A1(n11443), .A2(n11572), .ZN(n11575) );
  OAI211_X1 U13963 ( .C1(n11443), .C2(n11572), .A(n11575), .B(n12496), .ZN(
        n11449) );
  OAI22_X1 U13964 ( .A1(n11444), .A2(n12500), .B1(n11794), .B2(n12489), .ZN(
        n11445) );
  AOI211_X1 U13965 ( .C1(n11447), .C2(n12491), .A(n11446), .B(n11445), .ZN(
        n11448) );
  OAI211_X1 U13966 ( .C1(n11627), .C2(n12503), .A(n11449), .B(n11448), .ZN(
        P3_U3153) );
  NAND2_X1 U13967 ( .A1(n11450), .A2(n11453), .ZN(n11451) );
  NAND2_X1 U13968 ( .A1(n11452), .A2(n11451), .ZN(n15363) );
  OR2_X1 U13969 ( .A1(n15363), .A2(n8816), .ZN(n11459) );
  INV_X1 U13970 ( .A(n11453), .ZN(n11454) );
  XNOR2_X1 U13971 ( .A(n11455), .B(n11454), .ZN(n11457) );
  AOI21_X1 U13972 ( .B1(n11457), .B2(n13661), .A(n11456), .ZN(n11458) );
  NAND2_X1 U13973 ( .A1(n11459), .A2(n11458), .ZN(n15369) );
  NAND2_X1 U13974 ( .A1(n15369), .A2(n13643), .ZN(n11468) );
  OAI22_X1 U13975 ( .A1(n13643), .A2(n11461), .B1(n11460), .B2(n13655), .ZN(
        n11466) );
  NAND2_X1 U13976 ( .A1(n15364), .A2(n11462), .ZN(n11463) );
  NAND2_X1 U13977 ( .A1(n11463), .A2(n13604), .ZN(n11464) );
  OR2_X1 U13978 ( .A1(n11564), .A2(n11464), .ZN(n15365) );
  NOR2_X1 U13979 ( .A1(n13612), .A2(n15365), .ZN(n11465) );
  AOI211_X1 U13980 ( .C1(n13641), .C2(n15364), .A(n11466), .B(n11465), .ZN(
        n11467) );
  OAI211_X1 U13981 ( .C1(n15363), .C2(n11588), .A(n11468), .B(n11467), .ZN(
        P2_U3257) );
  NOR2_X1 U13982 ( .A1(n13167), .A2(SI_22_), .ZN(n11469) );
  AOI21_X1 U13983 ( .B1(n11470), .B2(P3_STATE_REG_SCAN_IN), .A(n11469), .ZN(
        n11471) );
  OAI21_X1 U13984 ( .B1(n11472), .B2(n13172), .A(n11471), .ZN(n11473) );
  INV_X1 U13985 ( .A(n11473), .ZN(P3_U3273) );
  INV_X1 U13986 ( .A(n11474), .ZN(n11482) );
  INV_X1 U13987 ( .A(n11475), .ZN(n11477) );
  MUX2_X1 U13988 ( .A(n11477), .B(n11476), .S(n13024), .Z(n11481) );
  AOI22_X1 U13989 ( .A1(n13008), .A2(n11479), .B1(n15463), .B2(n11478), .ZN(
        n11480) );
  OAI211_X1 U13990 ( .C1(n12088), .C2(n11482), .A(n11481), .B(n11480), .ZN(
        P3_U3230) );
  NAND2_X1 U13991 ( .A1(n11484), .A2(n11483), .ZN(n11771) );
  XNOR2_X1 U13992 ( .A(n15370), .B(n13213), .ZN(n11765) );
  NAND2_X1 U13993 ( .A1(n13651), .A2(n13374), .ZN(n11766) );
  XNOR2_X1 U13994 ( .A(n11765), .B(n11766), .ZN(n11770) );
  XNOR2_X1 U13995 ( .A(n11771), .B(n11770), .ZN(n11490) );
  NAND2_X1 U13996 ( .A1(n13336), .A2(n13373), .ZN(n11486) );
  NAND2_X1 U13997 ( .A1(n13337), .A2(n13375), .ZN(n11485) );
  AND2_X1 U13998 ( .A1(n11486), .A2(n11485), .ZN(n11585) );
  NAND2_X1 U13999 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3088), .ZN(n15257)
         );
  NAND2_X1 U14000 ( .A1(n13344), .A2(n11591), .ZN(n11487) );
  OAI211_X1 U14001 ( .C1(n13347), .C2(n11585), .A(n15257), .B(n11487), .ZN(
        n11488) );
  AOI21_X1 U14002 ( .B1(n15370), .B2(n15195), .A(n11488), .ZN(n11489) );
  OAI21_X1 U14003 ( .B1(n11490), .B2(n13349), .A(n11489), .ZN(P2_U3189) );
  NAND2_X1 U14004 ( .A1(n11491), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n11492) );
  NAND2_X1 U14005 ( .A1(n11493), .A2(n11492), .ZN(n15273) );
  INV_X1 U14006 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n14880) );
  MUX2_X1 U14007 ( .A(n14880), .B(P2_REG1_REG_12__SCAN_IN), .S(n15285), .Z(
        n15272) );
  NAND2_X1 U14008 ( .A1(n11494), .A2(n14880), .ZN(n11495) );
  NAND2_X1 U14009 ( .A1(n15275), .A2(n11495), .ZN(n15293) );
  INV_X1 U14010 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n11496) );
  MUX2_X1 U14011 ( .A(n11496), .B(P2_REG1_REG_13__SCAN_IN), .S(n15297), .Z(
        n15294) );
  NAND2_X1 U14012 ( .A1(n15297), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n11497) );
  NAND2_X1 U14013 ( .A1(n15290), .A2(n11497), .ZN(n15309) );
  INV_X1 U14014 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n11498) );
  OR2_X1 U14015 ( .A1(n15317), .A2(n11498), .ZN(n11500) );
  NAND2_X1 U14016 ( .A1(n15317), .A2(n11498), .ZN(n11499) );
  NAND2_X1 U14017 ( .A1(n11500), .A2(n11499), .ZN(n15308) );
  AOI21_X1 U14018 ( .B1(P2_REG1_REG_14__SCAN_IN), .B2(n15317), .A(n15310), 
        .ZN(n11597) );
  XNOR2_X1 U14019 ( .A(n11597), .B(n11596), .ZN(n11502) );
  INV_X1 U14020 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n11501) );
  NOR2_X1 U14021 ( .A1(n11501), .A2(n11502), .ZN(n11598) );
  INV_X1 U14022 ( .A(n15307), .ZN(n15292) );
  AOI211_X1 U14023 ( .C1(n11502), .C2(n11501), .A(n11598), .B(n15292), .ZN(
        n11514) );
  NOR2_X1 U14024 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n11503), .ZN(n11504) );
  AOI21_X1 U14025 ( .B1(n15313), .B2(P2_ADDR_REG_15__SCAN_IN), .A(n11504), 
        .ZN(n11512) );
  NAND2_X1 U14026 ( .A1(n15297), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n11507) );
  AND2_X1 U14027 ( .A1(n11505), .A2(n11758), .ZN(n15277) );
  MUX2_X1 U14028 ( .A(P2_REG2_REG_12__SCAN_IN), .B(n11823), .S(n15285), .Z(
        n15276) );
  OAI21_X1 U14029 ( .B1(n11506), .B2(n15277), .A(n15276), .ZN(n15282) );
  OAI21_X1 U14030 ( .B1(n15285), .B2(P2_REG2_REG_12__SCAN_IN), .A(n15282), 
        .ZN(n15300) );
  MUX2_X1 U14031 ( .A(n11971), .B(P2_REG2_REG_13__SCAN_IN), .S(n15297), .Z(
        n15299) );
  NAND2_X1 U14032 ( .A1(n11507), .A2(n15301), .ZN(n11508) );
  NAND2_X1 U14033 ( .A1(n15317), .A2(n11508), .ZN(n11509) );
  XOR2_X1 U14034 ( .A(n15317), .B(n11508), .Z(n15316) );
  NAND2_X1 U14035 ( .A1(n15316), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n15315) );
  NAND2_X1 U14036 ( .A1(n11509), .A2(n15315), .ZN(n11603) );
  XNOR2_X1 U14037 ( .A(n11596), .B(n11603), .ZN(n11510) );
  NAND2_X1 U14038 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n11510), .ZN(n11605) );
  OAI211_X1 U14039 ( .C1(P2_REG2_REG_15__SCAN_IN), .C2(n11510), .A(n15314), 
        .B(n11605), .ZN(n11511) );
  OAI211_X1 U14040 ( .C1(n15224), .C2(n11596), .A(n11512), .B(n11511), .ZN(
        n11513) );
  OR2_X1 U14041 ( .A1(n11514), .A2(n11513), .ZN(P2_U3229) );
  INV_X1 U14042 ( .A(n15439), .ZN(n11523) );
  NAND2_X1 U14043 ( .A1(n12737), .A2(n12485), .ZN(n11518) );
  AOI21_X1 U14044 ( .B1(n12491), .B2(n11516), .A(n11515), .ZN(n11517) );
  OAI211_X1 U14045 ( .C1(n11622), .C2(n12489), .A(n11518), .B(n11517), .ZN(
        n11522) );
  AOI211_X1 U14046 ( .C1(n11520), .C2(n11519), .A(n12494), .B(n6759), .ZN(
        n11521) );
  AOI211_X1 U14047 ( .C1(n11523), .C2(n12486), .A(n11522), .B(n11521), .ZN(
        n11524) );
  INV_X1 U14048 ( .A(n11524), .ZN(P3_U3179) );
  MUX2_X1 U14049 ( .A(n11525), .B(P3_REG2_REG_0__SCAN_IN), .S(n13024), .Z(
        n11529) );
  OAI22_X1 U14050 ( .A1(n15442), .A2(n11527), .B1(n15440), .B2(n11526), .ZN(
        n11528) );
  OR2_X1 U14051 ( .A1(n11529), .A2(n11528), .ZN(P3_U3233) );
  INV_X1 U14052 ( .A(n11530), .ZN(n11533) );
  OAI222_X1 U14053 ( .A1(n13798), .A2(n11532), .B1(n13804), .B2(n11533), .C1(
        P2_U3088), .C2(n11531), .ZN(P2_U3308) );
  OAI22_X1 U14054 ( .A1(n15442), .A2(n11535), .B1(n11534), .B2(n15440), .ZN(
        n11538) );
  MUX2_X1 U14055 ( .A(P3_REG2_REG_5__SCAN_IN), .B(n11536), .S(n15464), .Z(
        n11537) );
  AOI211_X1 U14056 ( .C1(n13039), .C2(n11539), .A(n11538), .B(n11537), .ZN(
        n11540) );
  INV_X1 U14057 ( .A(n11540), .ZN(P3_U3228) );
  OAI22_X1 U14058 ( .A1(n11557), .A2(n11299), .B1(n11544), .B2(n12284), .ZN(
        n11720) );
  NAND2_X1 U14059 ( .A1(n15141), .A2(n12300), .ZN(n11546) );
  NAND2_X1 U14060 ( .A1(n14225), .A2(n6622), .ZN(n11545) );
  NAND2_X1 U14061 ( .A1(n11546), .A2(n11545), .ZN(n11547) );
  XNOR2_X1 U14062 ( .A(n11547), .B(n12288), .ZN(n11719) );
  XOR2_X1 U14063 ( .A(n11720), .B(n11719), .Z(n11548) );
  OAI211_X1 U14064 ( .C1(n11549), .C2(n11548), .A(n11722), .B(n13912), .ZN(
        n11556) );
  INV_X1 U14065 ( .A(n11550), .ZN(n11554) );
  OAI21_X1 U14066 ( .B1(n13916), .B2(n11552), .A(n11551), .ZN(n11553) );
  AOI21_X1 U14067 ( .B1(n11554), .B2(n13918), .A(n11553), .ZN(n11555) );
  OAI211_X1 U14068 ( .C1(n11557), .C2(n13922), .A(n11556), .B(n11555), .ZN(
        P1_U3213) );
  XNOR2_X1 U14069 ( .A(n11558), .B(n11559), .ZN(n11739) );
  XNOR2_X1 U14070 ( .A(n11560), .B(n11559), .ZN(n11562) );
  AOI21_X1 U14071 ( .B1(n11562), .B2(n13661), .A(n11561), .ZN(n11563) );
  OAI21_X1 U14072 ( .B1(n11739), .B2(n8816), .A(n11563), .ZN(n11740) );
  NAND2_X1 U14073 ( .A1(n11740), .A2(n13643), .ZN(n11571) );
  INV_X1 U14074 ( .A(n11564), .ZN(n11565) );
  NAND2_X1 U14075 ( .A1(n11565), .A2(n11746), .ZN(n11566) );
  AND3_X1 U14076 ( .A1(n11589), .A2(n11566), .A3(n13604), .ZN(n11741) );
  NOR2_X1 U14077 ( .A1(n15330), .A2(n11743), .ZN(n11569) );
  OAI22_X1 U14078 ( .A1(n13643), .A2(n10471), .B1(n11567), .B2(n13655), .ZN(
        n11568) );
  AOI211_X1 U14079 ( .C1(n11741), .C2(n15324), .A(n11569), .B(n11568), .ZN(
        n11570) );
  OAI211_X1 U14080 ( .C1(n11739), .C2(n11588), .A(n11571), .B(n11570), .ZN(
        P2_U3256) );
  INV_X1 U14081 ( .A(n11572), .ZN(n11573) );
  NAND2_X1 U14082 ( .A1(n11573), .A2(n12735), .ZN(n11574) );
  NAND2_X1 U14083 ( .A1(n11575), .A2(n11574), .ZN(n11577) );
  XNOR2_X1 U14084 ( .A(n11685), .B(n6818), .ZN(n11787) );
  XNOR2_X1 U14085 ( .A(n11787), .B(n11794), .ZN(n11576) );
  NAND2_X1 U14086 ( .A1(n11577), .A2(n11576), .ZN(n11790) );
  OAI211_X1 U14087 ( .C1(n11577), .C2(n11576), .A(n11790), .B(n12496), .ZN(
        n11581) );
  OAI22_X1 U14088 ( .A1(n11871), .A2(n12489), .B1(n11622), .B2(n12500), .ZN(
        n11578) );
  AOI211_X1 U14089 ( .C1(n11685), .C2(n12491), .A(n11579), .B(n11578), .ZN(
        n11580) );
  OAI211_X1 U14090 ( .C1(n7578), .C2(n12503), .A(n11581), .B(n11580), .ZN(
        P3_U3161) );
  XNOR2_X1 U14091 ( .A(n11582), .B(n11583), .ZN(n15373) );
  INV_X1 U14092 ( .A(n8816), .ZN(n15361) );
  XNOR2_X1 U14093 ( .A(n11584), .B(n11583), .ZN(n11586) );
  OAI21_X1 U14094 ( .B1(n11586), .B2(n13623), .A(n11585), .ZN(n11587) );
  AOI21_X1 U14095 ( .B1(n15373), .B2(n15361), .A(n11587), .ZN(n15375) );
  INV_X1 U14096 ( .A(n11588), .ZN(n13614) );
  NAND2_X1 U14097 ( .A1(n15370), .A2(n11589), .ZN(n11590) );
  NAND3_X1 U14098 ( .A1(n11759), .A2(n13604), .A3(n11590), .ZN(n15371) );
  AOI22_X1 U14099 ( .A1(n6620), .A2(P2_REG2_REG_10__SCAN_IN), .B1(n11591), 
        .B2(n15326), .ZN(n11593) );
  NAND2_X1 U14100 ( .A1(n13641), .A2(n15370), .ZN(n11592) );
  OAI211_X1 U14101 ( .C1(n15371), .C2(n13612), .A(n11593), .B(n11592), .ZN(
        n11594) );
  AOI21_X1 U14102 ( .B1(n15373), .B2(n13614), .A(n11594), .ZN(n11595) );
  OAI21_X1 U14103 ( .B1(n15375), .B2(n6620), .A(n11595), .ZN(P2_U3255) );
  NOR2_X1 U14104 ( .A1(n11597), .A2(n11596), .ZN(n11599) );
  NOR2_X1 U14105 ( .A1(n11599), .A2(n11598), .ZN(n11602) );
  INV_X1 U14106 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n14864) );
  NOR2_X1 U14107 ( .A1(n11883), .A2(n14864), .ZN(n11600) );
  AOI21_X1 U14108 ( .B1(n11883), .B2(n14864), .A(n11600), .ZN(n11601) );
  NOR2_X1 U14109 ( .A1(n11602), .A2(n11601), .ZN(n11882) );
  AOI211_X1 U14110 ( .C1(n11602), .C2(n11601), .A(n15292), .B(n11882), .ZN(
        n11616) );
  NAND2_X1 U14111 ( .A1(n11604), .A2(n11603), .ZN(n11606) );
  NAND2_X1 U14112 ( .A1(n11606), .A2(n11605), .ZN(n11611) );
  NAND2_X1 U14113 ( .A1(n11883), .A2(n11607), .ZN(n11608) );
  OAI21_X1 U14114 ( .B1(n11883), .B2(n11607), .A(n11608), .ZN(n11610) );
  NAND2_X1 U14115 ( .A1(n11883), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n11609) );
  OAI211_X1 U14116 ( .C1(n11883), .C2(P2_REG2_REG_16__SCAN_IN), .A(n11611), 
        .B(n11609), .ZN(n11879) );
  OAI211_X1 U14117 ( .C1(n11611), .C2(n11610), .A(n11879), .B(n15314), .ZN(
        n11614) );
  NAND2_X1 U14118 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(P2_U3088), .ZN(n14854)
         );
  INV_X1 U14119 ( .A(n14854), .ZN(n11612) );
  AOI21_X1 U14120 ( .B1(n15313), .B2(P2_ADDR_REG_16__SCAN_IN), .A(n11612), 
        .ZN(n11613) );
  OAI211_X1 U14121 ( .C1(n15224), .C2(n11880), .A(n11614), .B(n11613), .ZN(
        n11615) );
  OR2_X1 U14122 ( .A1(n11616), .A2(n11615), .ZN(P2_U3230) );
  OAI21_X1 U14123 ( .B1(n11618), .B2(n12671), .A(n11617), .ZN(n11684) );
  INV_X1 U14124 ( .A(n11684), .ZN(n11626) );
  AOI21_X1 U14125 ( .B1(n12671), .B2(n11620), .A(n11619), .ZN(n11621) );
  OAI222_X1 U14126 ( .A1(n15452), .A2(n11622), .B1(n15450), .B2(n11871), .C1(
        n15457), .C2(n11621), .ZN(n11683) );
  NAND2_X1 U14127 ( .A1(n11683), .A2(n15464), .ZN(n11625) );
  OAI22_X1 U14128 ( .A1(n15442), .A2(n11689), .B1(n7578), .B2(n15440), .ZN(
        n11623) );
  AOI21_X1 U14129 ( .B1(P3_REG2_REG_8__SCAN_IN), .B2(n13024), .A(n11623), .ZN(
        n11624) );
  OAI211_X1 U14130 ( .C1(n12088), .C2(n11626), .A(n11625), .B(n11624), .ZN(
        P3_U3225) );
  OAI22_X1 U14131 ( .A1(n15442), .A2(n11628), .B1(n11627), .B2(n15440), .ZN(
        n11631) );
  MUX2_X1 U14132 ( .A(P3_REG2_REG_7__SCAN_IN), .B(n11629), .S(n15464), .Z(
        n11630) );
  AOI211_X1 U14133 ( .C1(n13039), .C2(n11632), .A(n11631), .B(n11630), .ZN(
        n11633) );
  INV_X1 U14134 ( .A(n11633), .ZN(P3_U3226) );
  XNOR2_X1 U14135 ( .A(n11634), .B(n11636), .ZN(n15171) );
  INV_X1 U14136 ( .A(n15171), .ZN(n11644) );
  AOI211_X1 U14137 ( .C1(n11636), .C2(n11635), .A(n15075), .B(n6758), .ZN(
        n15168) );
  NAND2_X1 U14138 ( .A1(n14223), .A2(n14921), .ZN(n15164) );
  INV_X1 U14139 ( .A(n15164), .ZN(n11637) );
  OAI21_X1 U14140 ( .B1(n15168), .B2(n11637), .A(n14539), .ZN(n11643) );
  OAI22_X1 U14141 ( .A1(n14539), .A2(n11638), .B1(n12063), .B2(n14602), .ZN(
        n11641) );
  XNOR2_X1 U14142 ( .A(n14613), .B(n14029), .ZN(n11639) );
  AOI22_X1 U14143 ( .A1(n11639), .A2(n15086), .B1(n14583), .B2(n14221), .ZN(
        n15165) );
  NOR2_X1 U14144 ( .A1(n15165), .A2(n14557), .ZN(n11640) );
  AOI211_X1 U14145 ( .C1(n15081), .C2(n14029), .A(n11641), .B(n11640), .ZN(
        n11642) );
  OAI211_X1 U14146 ( .C1(n11644), .C2(n15099), .A(n11643), .B(n11642), .ZN(
        P1_U3283) );
  NAND2_X1 U14147 ( .A1(n11645), .A2(n14796), .ZN(n11646) );
  OAI211_X1 U14148 ( .C1(n11647), .C2(n13167), .A(n11646), .B(n12725), .ZN(
        P3_U3272) );
  INV_X1 U14149 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n11896) );
  AOI22_X1 U14150 ( .A1(P3_REG2_REG_12__SCAN_IN), .A2(n11891), .B1(n11901), 
        .B2(n11896), .ZN(n11655) );
  AOI22_X1 U14151 ( .A1(n15416), .A2(n11651), .B1(P3_REG2_REG_10__SCAN_IN), 
        .B2(n11661), .ZN(n15422) );
  NAND2_X1 U14152 ( .A1(n11648), .A2(n11669), .ZN(n11650) );
  NAND2_X1 U14153 ( .A1(n11650), .A2(n11649), .ZN(n15421) );
  NAND2_X1 U14154 ( .A1(n15422), .A2(n15421), .ZN(n15420) );
  OAI21_X1 U14155 ( .B1(n15416), .B2(n11651), .A(n15420), .ZN(n11652) );
  NAND2_X1 U14156 ( .A1(n11652), .A2(n11713), .ZN(n11653) );
  XNOR2_X1 U14157 ( .A(n11652), .B(n11675), .ZN(n11707) );
  NAND2_X1 U14158 ( .A1(P3_REG2_REG_11__SCAN_IN), .A2(n11707), .ZN(n11706) );
  OAI21_X1 U14159 ( .B1(n11655), .B2(n11654), .A(n11895), .ZN(n11681) );
  NOR2_X1 U14160 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11656), .ZN(n12415) );
  AOI21_X1 U14161 ( .B1(n15415), .B2(P3_ADDR_REG_12__SCAN_IN), .A(n12415), 
        .ZN(n11668) );
  MUX2_X1 U14162 ( .A(P3_REG1_REG_10__SCAN_IN), .B(n11657), .S(n11661), .Z(
        n15424) );
  OAI21_X1 U14163 ( .B1(n11660), .B2(n11659), .A(n11658), .ZN(n15425) );
  NAND2_X1 U14164 ( .A1(n15424), .A2(n15425), .ZN(n15423) );
  MUX2_X1 U14165 ( .A(n11663), .B(P3_REG1_REG_12__SCAN_IN), .S(n11901), .Z(
        n11664) );
  NAND2_X1 U14166 ( .A1(n11664), .A2(n11665), .ZN(n11900) );
  OAI21_X1 U14167 ( .B1(n11665), .B2(n11664), .A(n11900), .ZN(n11666) );
  NAND2_X1 U14168 ( .A1(n15426), .A2(n11666), .ZN(n11667) );
  OAI211_X1 U14169 ( .C1(n11925), .C2(n11891), .A(n11668), .B(n11667), .ZN(
        n11680) );
  MUX2_X1 U14170 ( .A(P3_REG2_REG_12__SCAN_IN), .B(P3_REG1_REG_12__SCAN_IN), 
        .S(n13165), .Z(n11892) );
  XNOR2_X1 U14171 ( .A(n11892), .B(n11891), .ZN(n11678) );
  MUX2_X1 U14172 ( .A(P3_REG2_REG_10__SCAN_IN), .B(P3_REG1_REG_10__SCAN_IN), 
        .S(n13165), .Z(n11673) );
  XNOR2_X1 U14173 ( .A(n11673), .B(n15416), .ZN(n15418) );
  INV_X1 U14174 ( .A(n11673), .ZN(n11674) );
  AOI22_X1 U14175 ( .A1(n15419), .A2(n15418), .B1(n15416), .B2(n11674), .ZN(
        n11704) );
  MUX2_X1 U14176 ( .A(P3_REG2_REG_11__SCAN_IN), .B(P3_REG1_REG_11__SCAN_IN), 
        .S(n13165), .Z(n11676) );
  XOR2_X1 U14177 ( .A(n11675), .B(n11676), .Z(n11705) );
  OAI22_X1 U14178 ( .A1(n11704), .A2(n11705), .B1(n11676), .B2(n11713), .ZN(
        n11677) );
  NOR2_X1 U14179 ( .A1(n11677), .A2(n11678), .ZN(n11890) );
  AOI211_X1 U14180 ( .C1(n11678), .C2(n11677), .A(n15406), .B(n11890), .ZN(
        n11679) );
  AOI211_X1 U14181 ( .C1(n15429), .C2(n11681), .A(n11680), .B(n11679), .ZN(
        n11682) );
  INV_X1 U14182 ( .A(n11682), .ZN(P3_U3194) );
  AOI21_X1 U14183 ( .B1(n15477), .B2(n11684), .A(n11683), .ZN(n11692) );
  AOI22_X1 U14184 ( .A1(n11686), .A2(n11685), .B1(n6791), .B2(
        P3_REG1_REG_8__SCAN_IN), .ZN(n11687) );
  OAI21_X1 U14185 ( .B1(n11692), .B2(n6791), .A(n11687), .ZN(P3_U3467) );
  INV_X1 U14186 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n11688) );
  OAI22_X1 U14187 ( .A1(n11689), .A2(n13144), .B1(n15493), .B2(n11688), .ZN(
        n11690) );
  INV_X1 U14188 ( .A(n11690), .ZN(n11691) );
  OAI21_X1 U14189 ( .B1(n11692), .B2(n15491), .A(n11691), .ZN(P3_U3414) );
  XNOR2_X1 U14190 ( .A(n14910), .B(n14221), .ZN(n14180) );
  INV_X1 U14191 ( .A(n14180), .ZN(n11694) );
  XNOR2_X1 U14192 ( .A(n11693), .B(n11694), .ZN(n11805) );
  INV_X1 U14193 ( .A(n11805), .ZN(n11703) );
  XNOR2_X1 U14194 ( .A(n11695), .B(n14180), .ZN(n11696) );
  OAI222_X1 U14195 ( .A1(n14919), .A2(n14898), .B1(n14601), .B2(n14899), .C1(
        n11696), .C2(n15075), .ZN(n11803) );
  NAND2_X1 U14196 ( .A1(n11803), .A2(n14539), .ZN(n11702) );
  AOI211_X1 U14197 ( .C1(n14910), .C2(n11697), .A(n14915), .B(n7085), .ZN(
        n11804) );
  INV_X1 U14198 ( .A(n14910), .ZN(n11698) );
  NOR2_X1 U14199 ( .A1(n11698), .A2(n14570), .ZN(n11700) );
  OAI22_X1 U14200 ( .A1(n14539), .A2(n10180), .B1(n14913), .B2(n14602), .ZN(
        n11699) );
  AOI211_X1 U14201 ( .C1(n11804), .C2(n15090), .A(n11700), .B(n11699), .ZN(
        n11701) );
  OAI211_X1 U14202 ( .C1(n11703), .C2(n15099), .A(n11702), .B(n11701), .ZN(
        P1_U3282) );
  XOR2_X1 U14203 ( .A(n11704), .B(n11705), .Z(n11717) );
  OAI21_X1 U14204 ( .B1(n11707), .B2(P3_REG2_REG_11__SCAN_IN), .A(n11706), 
        .ZN(n11715) );
  NOR2_X1 U14205 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11708), .ZN(n12114) );
  XNOR2_X1 U14206 ( .A(n11709), .B(P3_REG1_REG_11__SCAN_IN), .ZN(n11710) );
  NOR2_X1 U14207 ( .A1(n12841), .A2(n11710), .ZN(n11711) );
  AOI211_X1 U14208 ( .C1(n15415), .C2(P3_ADDR_REG_11__SCAN_IN), .A(n12114), 
        .B(n11711), .ZN(n11712) );
  OAI21_X1 U14209 ( .B1(n11713), .B2(n11925), .A(n11712), .ZN(n11714) );
  AOI21_X1 U14210 ( .B1(n11715), .B2(n15429), .A(n11714), .ZN(n11716) );
  OAI21_X1 U14211 ( .B1(n11717), .B2(n15406), .A(n11716), .ZN(P3_U3193) );
  AOI22_X1 U14212 ( .A1(n14018), .A2(n12300), .B1(n6622), .B2(n14224), .ZN(
        n11718) );
  XNOR2_X1 U14213 ( .A(n11718), .B(n12288), .ZN(n11988) );
  AOI22_X1 U14214 ( .A1(n14018), .A2(n6622), .B1(n12301), .B2(n14224), .ZN(
        n11987) );
  XNOR2_X1 U14215 ( .A(n11988), .B(n11987), .ZN(n11724) );
  NAND2_X1 U14216 ( .A1(n11719), .A2(n11720), .ZN(n11721) );
  AOI21_X1 U14217 ( .B1(n11724), .B2(n11723), .A(n6761), .ZN(n11730) );
  NAND2_X1 U14218 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_U3086), .ZN(n14277) );
  OAI21_X1 U14219 ( .B1(n14897), .B2(n11990), .A(n14277), .ZN(n11725) );
  AOI21_X1 U14220 ( .B1(n13943), .B2(n14225), .A(n11725), .ZN(n11726) );
  OAI21_X1 U14221 ( .B1(n11727), .B2(n14914), .A(n11726), .ZN(n11728) );
  AOI21_X1 U14222 ( .B1(n14018), .B2(n14909), .A(n11728), .ZN(n11729) );
  OAI21_X1 U14223 ( .B1(n11730), .B2(n14904), .A(n11729), .ZN(P1_U3221) );
  XNOR2_X1 U14224 ( .A(n11731), .B(n12565), .ZN(n15488) );
  INV_X1 U14225 ( .A(n12927), .ZN(n12952) );
  OAI211_X1 U14226 ( .C1(n6768), .C2(n12565), .A(n11732), .B(n13032), .ZN(
        n11735) );
  OAI22_X1 U14227 ( .A1(n11794), .A2(n15452), .B1(n12006), .B2(n15450), .ZN(
        n11733) );
  INV_X1 U14228 ( .A(n11733), .ZN(n11734) );
  OAI211_X1 U14229 ( .C1(n12944), .C2(n15488), .A(n11735), .B(n11734), .ZN(
        n15490) );
  NAND2_X1 U14230 ( .A1(n15490), .A2(n15464), .ZN(n11738) );
  OAI22_X1 U14231 ( .A1(n15442), .A2(n15485), .B1(n11798), .B2(n15440), .ZN(
        n11736) );
  AOI21_X1 U14232 ( .B1(P3_REG2_REG_9__SCAN_IN), .B2(n13024), .A(n11736), .ZN(
        n11737) );
  OAI211_X1 U14233 ( .C1(n15488), .C2(n12952), .A(n11738), .B(n11737), .ZN(
        P3_U3224) );
  INV_X1 U14234 ( .A(n11739), .ZN(n11742) );
  AOI211_X1 U14235 ( .C1(n8890), .C2(n11742), .A(n11741), .B(n11740), .ZN(
        n11748) );
  OAI22_X1 U14236 ( .A1(n11743), .A2(n13783), .B1(n15383), .B2(n8499), .ZN(
        n11744) );
  INV_X1 U14237 ( .A(n11744), .ZN(n11745) );
  OAI21_X1 U14238 ( .B1(n11748), .B2(n15382), .A(n11745), .ZN(P2_U3457) );
  AOI22_X1 U14239 ( .A1(n12144), .A2(n11746), .B1(n15389), .B2(
        P2_REG1_REG_9__SCAN_IN), .ZN(n11747) );
  OAI21_X1 U14240 ( .B1(n11748), .B2(n15389), .A(n11747), .ZN(P2_U3508) );
  INV_X1 U14241 ( .A(n11749), .ZN(n11752) );
  INV_X1 U14242 ( .A(n11756), .ZN(n11751) );
  OAI21_X1 U14243 ( .B1(n11752), .B2(n11751), .A(n11750), .ZN(n11755) );
  NAND2_X1 U14244 ( .A1(n13336), .A2(n13372), .ZN(n11754) );
  NAND2_X1 U14245 ( .A1(n13337), .A2(n13374), .ZN(n11753) );
  NAND2_X1 U14246 ( .A1(n11754), .A2(n11753), .ZN(n11782) );
  AOI21_X1 U14247 ( .B1(n11755), .B2(n13661), .A(n11782), .ZN(n15377) );
  XOR2_X1 U14248 ( .A(n11757), .B(n11756), .Z(n15380) );
  NAND2_X1 U14249 ( .A1(n15380), .A2(n15333), .ZN(n11764) );
  OAI22_X1 U14250 ( .A1(n13643), .A2(n11758), .B1(n11779), .B2(n13655), .ZN(
        n11762) );
  INV_X1 U14251 ( .A(n11759), .ZN(n11760) );
  OAI211_X1 U14252 ( .C1(n6889), .C2(n11760), .A(n13604), .B(n11820), .ZN(
        n15376) );
  NOR2_X1 U14253 ( .A1(n15376), .A2(n13612), .ZN(n11761) );
  AOI211_X1 U14254 ( .C1(n13641), .C2(n11783), .A(n11762), .B(n11761), .ZN(
        n11763) );
  OAI211_X1 U14255 ( .C1(n6620), .C2(n15377), .A(n11764), .B(n11763), .ZN(
        P2_U3254) );
  INV_X1 U14256 ( .A(n11765), .ZN(n11768) );
  INV_X1 U14257 ( .A(n11766), .ZN(n11767) );
  NAND2_X1 U14258 ( .A1(n11768), .A2(n11767), .ZN(n11769) );
  XNOR2_X1 U14259 ( .A(n11783), .B(n13213), .ZN(n11772) );
  NAND2_X1 U14260 ( .A1(n13651), .A2(n13373), .ZN(n11773) );
  INV_X1 U14261 ( .A(n11772), .ZN(n11775) );
  INV_X1 U14262 ( .A(n11773), .ZN(n11774) );
  NAND2_X1 U14263 ( .A1(n11775), .A2(n11774), .ZN(n11776) );
  AOI21_X1 U14264 ( .B1(n11778), .B2(n11777), .A(n6762), .ZN(n11786) );
  NOR2_X1 U14265 ( .A1(n15198), .A2(n11779), .ZN(n11780) );
  AOI211_X1 U14266 ( .C1(n15190), .C2(n11782), .A(n11781), .B(n11780), .ZN(
        n11785) );
  NAND2_X1 U14267 ( .A1(n11783), .A2(n15195), .ZN(n11784) );
  OAI211_X1 U14268 ( .C1(n11786), .C2(n13349), .A(n11785), .B(n11784), .ZN(
        P2_U3208) );
  XNOR2_X1 U14269 ( .A(n15485), .B(n12392), .ZN(n11866) );
  XNOR2_X1 U14270 ( .A(n11866), .B(n12734), .ZN(n11793) );
  NAND2_X1 U14271 ( .A1(n11788), .A2(n11787), .ZN(n11789) );
  NAND2_X1 U14272 ( .A1(n11790), .A2(n11789), .ZN(n11792) );
  INV_X1 U14273 ( .A(n6783), .ZN(n11791) );
  AOI21_X1 U14274 ( .B1(n11793), .B2(n11792), .A(n11791), .ZN(n11802) );
  OAI22_X1 U14275 ( .A1(n11794), .A2(n12500), .B1(n12006), .B2(n12489), .ZN(
        n11795) );
  AOI211_X1 U14276 ( .C1(n11797), .C2(n12491), .A(n11796), .B(n11795), .ZN(
        n11801) );
  INV_X1 U14277 ( .A(n11798), .ZN(n11799) );
  NAND2_X1 U14278 ( .A1(n12486), .A2(n11799), .ZN(n11800) );
  OAI211_X1 U14279 ( .C1(n11802), .C2(n12494), .A(n11801), .B(n11800), .ZN(
        P3_U3171) );
  AOI211_X1 U14280 ( .C1(n11805), .C2(n15170), .A(n11804), .B(n11803), .ZN(
        n11809) );
  INV_X1 U14281 ( .A(n14748), .ZN(n14733) );
  NOR2_X1 U14282 ( .A1(n15174), .A2(n7927), .ZN(n11806) );
  AOI21_X1 U14283 ( .B1(n14910), .B2(n14733), .A(n11806), .ZN(n11807) );
  OAI21_X1 U14284 ( .B1(n11809), .B2(n15172), .A(n11807), .ZN(P1_U3492) );
  AOI22_X1 U14285 ( .A1(n14910), .A2(n8887), .B1(n15183), .B2(
        P1_REG1_REG_11__SCAN_IN), .ZN(n11808) );
  OAI21_X1 U14286 ( .B1(n11809), .B2(n15183), .A(n11808), .ZN(P1_U3539) );
  XNOR2_X1 U14287 ( .A(n11810), .B(n11811), .ZN(n14877) );
  NAND2_X1 U14288 ( .A1(n11812), .A2(n11811), .ZN(n11813) );
  NAND3_X1 U14289 ( .A1(n11814), .A2(n13661), .A3(n11813), .ZN(n11818) );
  NAND2_X1 U14290 ( .A1(n13336), .A2(n13371), .ZN(n11816) );
  NAND2_X1 U14291 ( .A1(n13337), .A2(n13373), .ZN(n11815) );
  NAND2_X1 U14292 ( .A1(n11816), .A2(n11815), .ZN(n15191) );
  INV_X1 U14293 ( .A(n15191), .ZN(n11817) );
  NAND2_X1 U14294 ( .A1(n11818), .A2(n11817), .ZN(n11819) );
  AOI21_X1 U14295 ( .B1(n14877), .B2(n15361), .A(n11819), .ZN(n14879) );
  NAND2_X1 U14296 ( .A1(n15194), .A2(n11820), .ZN(n11821) );
  NAND2_X1 U14297 ( .A1(n11821), .A2(n13604), .ZN(n11822) );
  OR2_X1 U14298 ( .A1(n11969), .A2(n11822), .ZN(n14875) );
  OAI22_X1 U14299 ( .A1(n13643), .A2(n11823), .B1(n15197), .B2(n13655), .ZN(
        n11824) );
  AOI21_X1 U14300 ( .B1(n15194), .B2(n13641), .A(n11824), .ZN(n11825) );
  OAI21_X1 U14301 ( .B1(n14875), .B2(n13612), .A(n11825), .ZN(n11826) );
  AOI21_X1 U14302 ( .B1(n14877), .B2(n13614), .A(n11826), .ZN(n11827) );
  OAI21_X1 U14303 ( .B1(n14879), .B2(n6620), .A(n11827), .ZN(P2_U3253) );
  INV_X1 U14304 ( .A(n11828), .ZN(n11831) );
  OAI222_X1 U14305 ( .A1(n13798), .A2(n11830), .B1(n13804), .B2(n11831), .C1(
        P2_U3088), .C2(n11829), .ZN(P2_U3306) );
  INV_X1 U14306 ( .A(n11835), .ZN(n12669) );
  XNOR2_X1 U14307 ( .A(n11833), .B(n12669), .ZN(n11958) );
  INV_X1 U14308 ( .A(n11958), .ZN(n11842) );
  OAI211_X1 U14309 ( .C1(n11836), .C2(n11835), .A(n11834), .B(n13032), .ZN(
        n11838) );
  AOI22_X1 U14310 ( .A1(n12416), .A2(n13029), .B1(n13027), .B2(n12734), .ZN(
        n11837) );
  NAND2_X1 U14311 ( .A1(n11838), .A2(n11837), .ZN(n11957) );
  NAND2_X1 U14312 ( .A1(n11957), .A2(n15464), .ZN(n11841) );
  OAI22_X1 U14313 ( .A1(n15442), .A2(n12574), .B1(n11877), .B2(n15440), .ZN(
        n11839) );
  AOI21_X1 U14314 ( .B1(P3_REG2_REG_10__SCAN_IN), .B2(n13024), .A(n11839), 
        .ZN(n11840) );
  OAI211_X1 U14315 ( .C1(n12088), .C2(n11842), .A(n11841), .B(n11840), .ZN(
        P3_U3223) );
  AOI21_X1 U14316 ( .B1(n14183), .B2(n11843), .A(n6744), .ZN(n14808) );
  AOI22_X1 U14317 ( .A1(n14921), .A2(n14221), .B1(n14922), .B2(n14583), .ZN(
        n11847) );
  XOR2_X1 U14318 ( .A(n14183), .B(n11844), .Z(n11845) );
  NAND2_X1 U14319 ( .A1(n11845), .A2(n14952), .ZN(n11846) );
  OAI211_X1 U14320 ( .C1(n14808), .C2(n15129), .A(n11847), .B(n11846), .ZN(
        n14810) );
  NAND2_X1 U14321 ( .A1(n14810), .A2(n14539), .ZN(n11852) );
  OAI22_X1 U14322 ( .A1(n14539), .A2(n11848), .B1(n13856), .B2(n14602), .ZN(
        n11850) );
  OAI211_X1 U14323 ( .C1(n7084), .C2(n7085), .A(n15086), .B(n11859), .ZN(
        n14809) );
  NOR2_X1 U14324 ( .A1(n14809), .A2(n14557), .ZN(n11849) );
  AOI211_X1 U14325 ( .C1(n15081), .C2(n14040), .A(n11850), .B(n11849), .ZN(
        n11851) );
  OAI211_X1 U14326 ( .C1(n14808), .C2(n15082), .A(n11852), .B(n11851), .ZN(
        P1_U3281) );
  OAI21_X1 U14327 ( .B1(n11855), .B2(n11854), .A(n11853), .ZN(n11980) );
  INV_X1 U14328 ( .A(n11980), .ZN(n11865) );
  XNOR2_X1 U14329 ( .A(n11856), .B(n14185), .ZN(n11857) );
  OAI222_X1 U14330 ( .A1(n14919), .A2(n13904), .B1(n14601), .B2(n14898), .C1(
        n11857), .C2(n15075), .ZN(n11978) );
  NAND2_X1 U14331 ( .A1(n11978), .A2(n14539), .ZN(n11864) );
  INV_X1 U14332 ( .A(n11858), .ZN(n14916) );
  AOI211_X1 U14333 ( .C1(n14043), .C2(n11859), .A(n14915), .B(n11858), .ZN(
        n11979) );
  NOR2_X1 U14334 ( .A1(n14044), .A2(n14570), .ZN(n11862) );
  OAI22_X1 U14335 ( .A1(n14539), .A2(n11860), .B1(n13903), .B2(n14602), .ZN(
        n11861) );
  AOI211_X1 U14336 ( .C1(n11979), .C2(n15090), .A(n11862), .B(n11861), .ZN(
        n11863) );
  OAI211_X1 U14337 ( .C1(n11865), .C2(n15099), .A(n11864), .B(n11863), .ZN(
        P1_U3280) );
  INV_X1 U14338 ( .A(n11866), .ZN(n11867) );
  NAND2_X1 U14339 ( .A1(n11867), .A2(n11871), .ZN(n11868) );
  XNOR2_X1 U14340 ( .A(n11874), .B(n6818), .ZN(n12030) );
  XNOR2_X1 U14341 ( .A(n12030), .B(n12006), .ZN(n11870) );
  OAI211_X1 U14342 ( .C1(n6753), .C2(n11870), .A(n12032), .B(n12496), .ZN(
        n11876) );
  NAND2_X1 U14343 ( .A1(P3_REG3_REG_10__SCAN_IN), .A2(P3_U3151), .ZN(n15432)
         );
  INV_X1 U14344 ( .A(n15432), .ZN(n11873) );
  OAI22_X1 U14345 ( .A1(n11871), .A2(n12500), .B1(n12113), .B2(n12489), .ZN(
        n11872) );
  AOI211_X1 U14346 ( .C1(n11874), .C2(n12491), .A(n11873), .B(n11872), .ZN(
        n11875) );
  OAI211_X1 U14347 ( .C1(n11877), .C2(n12503), .A(n11876), .B(n11875), .ZN(
        P3_U3157) );
  NAND2_X1 U14348 ( .A1(n13407), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n11878) );
  OAI21_X1 U14349 ( .B1(n13407), .B2(P2_REG2_REG_17__SCAN_IN), .A(n11878), 
        .ZN(n13400) );
  OAI21_X1 U14350 ( .B1(n11607), .B2(n11880), .A(n11879), .ZN(n13401) );
  XOR2_X1 U14351 ( .A(n13400), .B(n13401), .Z(n11889) );
  NAND2_X1 U14352 ( .A1(P2_U3088), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n11881)
         );
  OAI21_X1 U14353 ( .B1(n15306), .B2(n14815), .A(n11881), .ZN(n11887) );
  AOI21_X1 U14354 ( .B1(n11883), .B2(P2_REG1_REG_16__SCAN_IN), .A(n11882), 
        .ZN(n11885) );
  XNOR2_X1 U14355 ( .A(n13407), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n11884) );
  NOR2_X1 U14356 ( .A1(n11885), .A2(n11884), .ZN(n13406) );
  AOI211_X1 U14357 ( .C1(n11885), .C2(n11884), .A(n15292), .B(n13406), .ZN(
        n11886) );
  AOI211_X1 U14358 ( .C1(n15318), .C2(n13407), .A(n11887), .B(n11886), .ZN(
        n11888) );
  OAI21_X1 U14359 ( .B1(n11889), .B2(n15298), .A(n11888), .ZN(P2_U3231) );
  MUX2_X1 U14360 ( .A(P3_REG2_REG_13__SCAN_IN), .B(P3_REG1_REG_13__SCAN_IN), 
        .S(n13165), .Z(n11932) );
  XNOR2_X1 U14361 ( .A(n11932), .B(n11899), .ZN(n11893) );
  OAI21_X1 U14362 ( .B1(n11894), .B2(n11893), .A(n11930), .ZN(n11909) );
  NAND2_X1 U14363 ( .A1(P3_REG2_REG_13__SCAN_IN), .A2(n11897), .ZN(n11918) );
  OAI21_X1 U14364 ( .B1(P3_REG2_REG_13__SCAN_IN), .B2(n11897), .A(n11918), 
        .ZN(n11898) );
  NAND2_X1 U14365 ( .A1(n11898), .A2(n15429), .ZN(n11907) );
  AND2_X1 U14366 ( .A1(P3_U3151), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n12043) );
  AOI21_X1 U14367 ( .B1(n15415), .B2(P3_ADDR_REG_13__SCAN_IN), .A(n12043), 
        .ZN(n11906) );
  NAND2_X1 U14368 ( .A1(n15417), .A2(n11899), .ZN(n11905) );
  OAI21_X1 U14369 ( .B1(n11902), .B2(P3_REG1_REG_13__SCAN_IN), .A(n11912), 
        .ZN(n11903) );
  NAND2_X1 U14370 ( .A1(n15426), .A2(n11903), .ZN(n11904) );
  NAND4_X1 U14371 ( .A1(n11907), .A2(n11906), .A3(n11905), .A4(n11904), .ZN(
        n11908) );
  AOI21_X1 U14372 ( .B1(n11909), .B2(n15430), .A(n11908), .ZN(n11910) );
  INV_X1 U14373 ( .A(n11910), .ZN(P3_U3195) );
  NAND2_X1 U14374 ( .A1(n11931), .A2(n11911), .ZN(n11913) );
  NAND2_X1 U14375 ( .A1(n11913), .A2(n11912), .ZN(n11916) );
  OR2_X1 U14376 ( .A1(n12746), .A2(n11914), .ZN(n12743) );
  NAND2_X1 U14377 ( .A1(n12746), .A2(n11914), .ZN(n11915) );
  AND2_X1 U14378 ( .A1(n12743), .A2(n11915), .ZN(n11927) );
  NAND2_X1 U14379 ( .A1(n11927), .A2(n11916), .ZN(n12742) );
  OAI21_X1 U14380 ( .B1(n11916), .B2(n11927), .A(n12742), .ZN(n11937) );
  NAND2_X1 U14381 ( .A1(n11931), .A2(n11917), .ZN(n11919) );
  XNOR2_X1 U14382 ( .A(n12746), .B(P3_REG2_REG_14__SCAN_IN), .ZN(n11926) );
  OAI21_X1 U14383 ( .B1(n11920), .B2(n11926), .A(n12744), .ZN(n11921) );
  NAND2_X1 U14384 ( .A1(n11921), .A2(n15429), .ZN(n11924) );
  NAND2_X1 U14385 ( .A1(P3_U3151), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n12107)
         );
  INV_X1 U14386 ( .A(n12107), .ZN(n11922) );
  AOI21_X1 U14387 ( .B1(n15415), .B2(P3_ADDR_REG_14__SCAN_IN), .A(n11922), 
        .ZN(n11923) );
  OAI211_X1 U14388 ( .C1(n11925), .C2(n12756), .A(n11924), .B(n11923), .ZN(
        n11936) );
  INV_X1 U14389 ( .A(n11926), .ZN(n11929) );
  INV_X1 U14390 ( .A(n11927), .ZN(n11928) );
  MUX2_X1 U14391 ( .A(n11929), .B(n11928), .S(n13165), .Z(n11934) );
  NOR2_X1 U14392 ( .A1(n11933), .A2(n11934), .ZN(n12754) );
  AOI211_X1 U14393 ( .C1(n11934), .C2(n11933), .A(n15406), .B(n12754), .ZN(
        n11935) );
  AOI211_X1 U14394 ( .C1(n15426), .C2(n11937), .A(n11936), .B(n11935), .ZN(
        n11938) );
  INV_X1 U14395 ( .A(n11938), .ZN(P3_U3196) );
  XNOR2_X1 U14396 ( .A(n15194), .B(n13213), .ZN(n11940) );
  NAND2_X1 U14397 ( .A1(n13651), .A2(n13372), .ZN(n11941) );
  NAND2_X1 U14398 ( .A1(n11940), .A2(n11941), .ZN(n15187) );
  NAND2_X1 U14399 ( .A1(n15186), .A2(n15187), .ZN(n11944) );
  INV_X1 U14400 ( .A(n11940), .ZN(n11943) );
  INV_X1 U14401 ( .A(n11941), .ZN(n11942) );
  NAND2_X1 U14402 ( .A1(n11943), .A2(n11942), .ZN(n15188) );
  XNOR2_X1 U14403 ( .A(n11973), .B(n13255), .ZN(n11945) );
  AND2_X1 U14404 ( .A1(n13651), .A2(n13371), .ZN(n11946) );
  NAND2_X1 U14405 ( .A1(n11945), .A2(n11946), .ZN(n13173) );
  INV_X1 U14406 ( .A(n11945), .ZN(n11948) );
  INV_X1 U14407 ( .A(n11946), .ZN(n11947) );
  NAND2_X1 U14408 ( .A1(n11948), .A2(n11947), .ZN(n11949) );
  AND2_X1 U14409 ( .A1(n13173), .A2(n11949), .ZN(n11950) );
  OAI211_X1 U14410 ( .C1(n11951), .C2(n11950), .A(n13174), .B(n15193), .ZN(
        n11956) );
  OAI22_X1 U14411 ( .A1(n11953), .A2(n13301), .B1(n11952), .B2(n13303), .ZN(
        n11964) );
  OAI22_X1 U14412 ( .A1(n15198), .A2(n11970), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n15289), .ZN(n11954) );
  AOI21_X1 U14413 ( .B1(n15190), .B2(n11964), .A(n11954), .ZN(n11955) );
  OAI211_X1 U14414 ( .C1(n14871), .C2(n13331), .A(n11956), .B(n11955), .ZN(
        P2_U3206) );
  INV_X1 U14415 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n11959) );
  AOI21_X1 U14416 ( .B1(n11958), .B2(n15477), .A(n11957), .ZN(n11961) );
  MUX2_X1 U14417 ( .A(n11959), .B(n11961), .S(n15493), .Z(n11960) );
  OAI21_X1 U14418 ( .B1(n13144), .B2(n12574), .A(n11960), .ZN(P3_U3420) );
  MUX2_X1 U14419 ( .A(n11657), .B(n11961), .S(n15498), .Z(n11962) );
  OAI21_X1 U14420 ( .B1(n13092), .B2(n12574), .A(n11962), .ZN(P3_U3469) );
  XNOR2_X1 U14421 ( .A(n11963), .B(n11967), .ZN(n11966) );
  INV_X1 U14422 ( .A(n11964), .ZN(n11965) );
  OAI21_X1 U14423 ( .B1(n11966), .B2(n13623), .A(n11965), .ZN(n14872) );
  INV_X1 U14424 ( .A(n14872), .ZN(n11977) );
  XNOR2_X1 U14425 ( .A(n11968), .B(n11967), .ZN(n14874) );
  OAI211_X1 U14426 ( .C1(n14871), .C2(n11969), .A(n13604), .B(n12020), .ZN(
        n14870) );
  OAI22_X1 U14427 ( .A1(n13643), .A2(n11971), .B1(n11970), .B2(n13655), .ZN(
        n11972) );
  AOI21_X1 U14428 ( .B1(n11973), .B2(n13641), .A(n11972), .ZN(n11974) );
  OAI21_X1 U14429 ( .B1(n14870), .B2(n13612), .A(n11974), .ZN(n11975) );
  AOI21_X1 U14430 ( .B1(n14874), .B2(n15333), .A(n11975), .ZN(n11976) );
  OAI21_X1 U14431 ( .B1(n11977), .B2(n6620), .A(n11976), .ZN(P2_U3252) );
  AOI211_X1 U14432 ( .C1(n15170), .C2(n11980), .A(n11979), .B(n11978), .ZN(
        n11985) );
  AOI22_X1 U14433 ( .A1(n14043), .A2(n8887), .B1(n15183), .B2(
        P1_REG1_REG_13__SCAN_IN), .ZN(n11981) );
  OAI21_X1 U14434 ( .B1(n11985), .B2(n15183), .A(n11981), .ZN(P1_U3541) );
  INV_X1 U14435 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n11982) );
  OAI22_X1 U14436 ( .A1(n14044), .A2(n14748), .B1(n15174), .B2(n11982), .ZN(
        n11983) );
  INV_X1 U14437 ( .A(n11983), .ZN(n11984) );
  OAI21_X1 U14438 ( .B1(n11985), .B2(n15172), .A(n11984), .ZN(P1_U3498) );
  AOI22_X1 U14439 ( .A1(n15156), .A2(n12300), .B1(n6622), .B2(n14223), .ZN(
        n11986) );
  XNOR2_X1 U14440 ( .A(n11986), .B(n12208), .ZN(n12055) );
  NOR2_X1 U14441 ( .A1(n12284), .A2(n11990), .ZN(n11991) );
  AOI21_X1 U14442 ( .B1(n15156), .B2(n6622), .A(n11991), .ZN(n12054) );
  XOR2_X1 U14443 ( .A(n12056), .B(n12055), .Z(n11996) );
  NAND2_X1 U14444 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_U3086), .ZN(n14291) );
  OAI21_X1 U14445 ( .B1(n14897), .B2(n14899), .A(n14291), .ZN(n11992) );
  AOI21_X1 U14446 ( .B1(n13943), .B2(n14224), .A(n11992), .ZN(n11993) );
  OAI21_X1 U14447 ( .B1(n14603), .B2(n14914), .A(n11993), .ZN(n11994) );
  AOI21_X1 U14448 ( .B1(n15156), .B2(n14909), .A(n11994), .ZN(n11995) );
  OAI21_X1 U14449 ( .B1(n11996), .B2(n14904), .A(n11995), .ZN(P1_U3231) );
  NAND2_X1 U14450 ( .A1(n11999), .A2(n14757), .ZN(n11997) );
  OAI211_X1 U14451 ( .C1(n11998), .C2(n14774), .A(n11997), .B(n14209), .ZN(
        P1_U3332) );
  NAND2_X1 U14452 ( .A1(n11999), .A2(n13792), .ZN(n12001) );
  OAI211_X1 U14453 ( .C1(n12002), .C2(n13798), .A(n12001), .B(n12000), .ZN(
        P2_U3304) );
  XNOR2_X1 U14454 ( .A(n12003), .B(n12682), .ZN(n12094) );
  INV_X1 U14455 ( .A(n12094), .ZN(n12010) );
  XOR2_X1 U14456 ( .A(n12682), .B(n12004), .Z(n12005) );
  OAI222_X1 U14457 ( .A1(n15450), .A2(n12081), .B1(n15452), .B2(n12006), .C1(
        n12005), .C2(n15457), .ZN(n12093) );
  NAND2_X1 U14458 ( .A1(n12093), .A2(n15464), .ZN(n12009) );
  OAI22_X1 U14459 ( .A1(n15442), .A2(n12099), .B1(n12115), .B2(n15440), .ZN(
        n12007) );
  AOI21_X1 U14460 ( .B1(P3_REG2_REG_11__SCAN_IN), .B2(n13024), .A(n12007), 
        .ZN(n12008) );
  OAI211_X1 U14461 ( .C1(n12010), .C2(n12088), .A(n12009), .B(n12008), .ZN(
        P3_U3222) );
  INV_X1 U14462 ( .A(n12019), .ZN(n12011) );
  XNOR2_X1 U14463 ( .A(n12012), .B(n12011), .ZN(n12013) );
  NAND2_X1 U14464 ( .A1(n12013), .A2(n13661), .ZN(n12017) );
  NAND2_X1 U14465 ( .A1(n13369), .A2(n13336), .ZN(n12015) );
  NAND2_X1 U14466 ( .A1(n13337), .A2(n13371), .ZN(n12014) );
  NAND2_X1 U14467 ( .A1(n12015), .A2(n12014), .ZN(n14844) );
  INV_X1 U14468 ( .A(n14844), .ZN(n12016) );
  NAND2_X1 U14469 ( .A1(n12017), .A2(n12016), .ZN(n14868) );
  INV_X1 U14470 ( .A(n14868), .ZN(n12027) );
  XOR2_X1 U14471 ( .A(n12019), .B(n12018), .Z(n14869) );
  INV_X1 U14472 ( .A(n14845), .ZN(n14866) );
  INV_X1 U14473 ( .A(n12020), .ZN(n12021) );
  OAI211_X1 U14474 ( .C1(n14866), .C2(n12021), .A(n13604), .B(n12139), .ZN(
        n14865) );
  OAI22_X1 U14475 ( .A1(n13643), .A2(n12022), .B1(n14847), .B2(n13655), .ZN(
        n12023) );
  AOI21_X1 U14476 ( .B1(n14845), .B2(n13641), .A(n12023), .ZN(n12024) );
  OAI21_X1 U14477 ( .B1(n14865), .B2(n13612), .A(n12024), .ZN(n12025) );
  AOI21_X1 U14478 ( .B1(n14869), .B2(n15333), .A(n12025), .ZN(n12026) );
  OAI21_X1 U14479 ( .B1(n6620), .B2(n12027), .A(n12026), .ZN(P2_U3251) );
  XNOR2_X1 U14480 ( .A(n14822), .B(n6818), .ZN(n12029) );
  INV_X1 U14481 ( .A(n12029), .ZN(n12028) );
  NAND2_X1 U14482 ( .A1(n12028), .A2(n12419), .ZN(n12102) );
  NAND2_X1 U14483 ( .A1(n12029), .A2(n12070), .ZN(n12100) );
  NAND2_X1 U14484 ( .A1(n12102), .A2(n12100), .ZN(n12041) );
  NAND2_X1 U14485 ( .A1(n12733), .A2(n12030), .ZN(n12031) );
  XNOR2_X1 U14486 ( .A(n12099), .B(n6818), .ZN(n12034) );
  XNOR2_X1 U14487 ( .A(n12417), .B(n12392), .ZN(n12412) );
  AOI22_X1 U14488 ( .A1(n12113), .A2(n12034), .B1(n12412), .B2(n12081), .ZN(
        n12033) );
  INV_X1 U14489 ( .A(n12412), .ZN(n12038) );
  INV_X1 U14490 ( .A(n12034), .ZN(n12410) );
  NAND2_X1 U14491 ( .A1(n12416), .A2(n12410), .ZN(n12035) );
  NAND2_X1 U14492 ( .A1(n12035), .A2(n12081), .ZN(n12037) );
  INV_X1 U14493 ( .A(n12035), .ZN(n12036) );
  AOI22_X1 U14494 ( .A1(n12038), .A2(n12037), .B1(n12036), .B2(n12732), .ZN(
        n12039) );
  NAND2_X1 U14495 ( .A1(n12040), .A2(n12039), .ZN(n12101) );
  XOR2_X1 U14496 ( .A(n12041), .B(n12101), .Z(n12047) );
  INV_X1 U14497 ( .A(n14822), .ZN(n12085) );
  NOR2_X1 U14498 ( .A1(n12081), .A2(n12500), .ZN(n12042) );
  AOI211_X1 U14499 ( .C1(n12506), .C2(n12731), .A(n12043), .B(n12042), .ZN(
        n12044) );
  OAI21_X1 U14500 ( .B1(n12082), .B2(n12503), .A(n12044), .ZN(n12045) );
  AOI21_X1 U14501 ( .B1(n12085), .B2(n12491), .A(n12045), .ZN(n12046) );
  OAI21_X1 U14502 ( .B1(n12047), .B2(n12494), .A(n12046), .ZN(P3_U3174) );
  INV_X1 U14503 ( .A(n12048), .ZN(n12049) );
  OAI222_X1 U14504 ( .A1(P3_U3151), .A2(n12051), .B1(n13167), .B2(n12050), 
        .C1(n13172), .C2(n12049), .ZN(P3_U3271) );
  INV_X1 U14505 ( .A(n12052), .ZN(n12053) );
  NAND2_X1 U14506 ( .A1(n14029), .A2(n12300), .ZN(n12058) );
  NAND2_X1 U14507 ( .A1(n14222), .A2(n6622), .ZN(n12057) );
  NAND2_X1 U14508 ( .A1(n12058), .A2(n12057), .ZN(n12059) );
  XNOR2_X1 U14509 ( .A(n12059), .B(n12208), .ZN(n12181) );
  NOR2_X1 U14510 ( .A1(n12284), .A2(n14899), .ZN(n12060) );
  AOI21_X1 U14511 ( .B1(n14029), .B2(n6622), .A(n12060), .ZN(n12179) );
  XNOR2_X1 U14512 ( .A(n12181), .B(n12179), .ZN(n12061) );
  OAI211_X1 U14513 ( .C1(n12062), .C2(n12061), .A(n12182), .B(n13912), .ZN(
        n12067) );
  NOR2_X1 U14514 ( .A1(n14914), .A2(n12063), .ZN(n12065) );
  OAI22_X1 U14515 ( .A1(n14897), .A2(n12177), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n7923), .ZN(n12064) );
  AOI211_X1 U14516 ( .C1(n13943), .C2(n14223), .A(n12065), .B(n12064), .ZN(
        n12066) );
  OAI211_X1 U14517 ( .C1(n15167), .C2(n13922), .A(n12067), .B(n12066), .ZN(
        P1_U3217) );
  XNOR2_X1 U14518 ( .A(n12068), .B(n12681), .ZN(n12069) );
  OAI222_X1 U14519 ( .A1(n15450), .A2(n12070), .B1(n15452), .B2(n12113), .C1(
        n12069), .C2(n15457), .ZN(n14828) );
  INV_X1 U14520 ( .A(n14828), .ZN(n12077) );
  OAI21_X1 U14521 ( .B1(n12072), .B2(n12681), .A(n12071), .ZN(n14830) );
  INV_X1 U14522 ( .A(n12073), .ZN(n12418) );
  AOI22_X1 U14523 ( .A1(n13024), .A2(P3_REG2_REG_12__SCAN_IN), .B1(n15463), 
        .B2(n12418), .ZN(n12074) );
  OAI21_X1 U14524 ( .B1(n14827), .B2(n15442), .A(n12074), .ZN(n12075) );
  AOI21_X1 U14525 ( .B1(n14830), .B2(n13039), .A(n12075), .ZN(n12076) );
  OAI21_X1 U14526 ( .B1(n12077), .B2(n13024), .A(n12076), .ZN(P3_U3221) );
  XNOR2_X1 U14527 ( .A(n12078), .B(n12685), .ZN(n14824) );
  INV_X1 U14528 ( .A(n12731), .ZN(n12501) );
  XNOR2_X1 U14529 ( .A(n12079), .B(n12685), .ZN(n12080) );
  OAI222_X1 U14530 ( .A1(n15450), .A2(n12501), .B1(n15452), .B2(n12081), .C1(
        n12080), .C2(n15457), .ZN(n14826) );
  NAND2_X1 U14531 ( .A1(n14826), .A2(n15464), .ZN(n12087) );
  INV_X1 U14532 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n12083) );
  OAI22_X1 U14533 ( .A1(n15464), .A2(n12083), .B1(n12082), .B2(n15440), .ZN(
        n12084) );
  AOI21_X1 U14534 ( .B1(n12085), .B2(n13008), .A(n12084), .ZN(n12086) );
  OAI211_X1 U14535 ( .C1(n12088), .C2(n14824), .A(n12087), .B(n12086), .ZN(
        P3_U3220) );
  INV_X1 U14536 ( .A(n12089), .ZN(n12090) );
  OAI222_X1 U14537 ( .A1(P3_U3151), .A2(n12092), .B1(n13167), .B2(n12091), 
        .C1(n13172), .C2(n12090), .ZN(P3_U3270) );
  INV_X1 U14538 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n12095) );
  AOI21_X1 U14539 ( .B1(n12094), .B2(n15477), .A(n12093), .ZN(n12097) );
  MUX2_X1 U14540 ( .A(n12095), .B(n12097), .S(n15493), .Z(n12096) );
  OAI21_X1 U14541 ( .B1(n13144), .B2(n12099), .A(n12096), .ZN(P3_U3423) );
  MUX2_X1 U14542 ( .A(n11662), .B(n12097), .S(n15498), .Z(n12098) );
  OAI21_X1 U14543 ( .B1(n13092), .B2(n12099), .A(n12098), .ZN(P3_U3470) );
  NAND2_X1 U14544 ( .A1(n12101), .A2(n12100), .ZN(n12103) );
  NAND2_X1 U14545 ( .A1(n12103), .A2(n12102), .ZN(n12105) );
  XNOR2_X1 U14546 ( .A(n12130), .B(n6818), .ZN(n12336) );
  XNOR2_X1 U14547 ( .A(n12336), .B(n12731), .ZN(n12104) );
  NAND2_X1 U14548 ( .A1(n12105), .A2(n12104), .ZN(n12339) );
  OAI211_X1 U14549 ( .C1(n12105), .C2(n12104), .A(n12339), .B(n12496), .ZN(
        n12111) );
  INV_X1 U14550 ( .A(n12106), .ZN(n12128) );
  NAND2_X1 U14551 ( .A1(n12485), .A2(n12419), .ZN(n12108) );
  OAI211_X1 U14552 ( .C1(n12599), .C2(n12489), .A(n12108), .B(n12107), .ZN(
        n12109) );
  AOI21_X1 U14553 ( .B1(n12128), .B2(n12486), .A(n12109), .ZN(n12110) );
  OAI211_X1 U14554 ( .C1(n12509), .C2(n12130), .A(n12111), .B(n12110), .ZN(
        P3_U3155) );
  XNOR2_X1 U14555 ( .A(n12411), .B(n12410), .ZN(n12112) );
  NOR2_X1 U14556 ( .A1(n12112), .A2(n12113), .ZN(n12409) );
  AOI211_X1 U14557 ( .C1(n12113), .C2(n12112), .A(n12494), .B(n12409), .ZN(
        n12123) );
  AOI21_X1 U14558 ( .B1(n12733), .B2(n12485), .A(n12114), .ZN(n12121) );
  INV_X1 U14559 ( .A(n12115), .ZN(n12116) );
  NAND2_X1 U14560 ( .A1(n12486), .A2(n12116), .ZN(n12120) );
  NAND2_X1 U14561 ( .A1(n12491), .A2(n12117), .ZN(n12119) );
  NAND2_X1 U14562 ( .A1(n12732), .A2(n12506), .ZN(n12118) );
  NAND4_X1 U14563 ( .A1(n12121), .A2(n12120), .A3(n12119), .A4(n12118), .ZN(
        n12122) );
  OR2_X1 U14564 ( .A1(n12123), .A2(n12122), .ZN(P3_U3176) );
  INV_X1 U14565 ( .A(n12126), .ZN(n12688) );
  XNOR2_X1 U14566 ( .A(n12124), .B(n12688), .ZN(n12125) );
  AOI222_X1 U14567 ( .A1(n13032), .A2(n12125), .B1(n12419), .B2(n13027), .C1(
        n13028), .C2(n13029), .ZN(n13104) );
  XNOR2_X1 U14568 ( .A(n12127), .B(n12126), .ZN(n13102) );
  AOI22_X1 U14569 ( .A1(n13024), .A2(P3_REG2_REG_14__SCAN_IN), .B1(n15463), 
        .B2(n12128), .ZN(n12129) );
  OAI21_X1 U14570 ( .B1(n12130), .B2(n15442), .A(n12129), .ZN(n12131) );
  AOI21_X1 U14571 ( .B1(n13102), .B2(n13039), .A(n12131), .ZN(n12132) );
  OAI21_X1 U14572 ( .B1(n13104), .B2(n13024), .A(n12132), .ZN(P3_U3219) );
  INV_X1 U14573 ( .A(n12133), .ZN(n12137) );
  OAI222_X1 U14574 ( .A1(n13798), .A2(n6823), .B1(n13804), .B2(n12137), .C1(
        n12136), .C2(P2_U3088), .ZN(P2_U3303) );
  OAI21_X1 U14575 ( .B1(n6743), .B2(n12141), .A(n12138), .ZN(n13637) );
  AOI21_X1 U14576 ( .B1(n13642), .B2(n12139), .A(n13651), .ZN(n12140) );
  AND2_X1 U14577 ( .A1(n12140), .A2(n12162), .ZN(n13645) );
  XNOR2_X1 U14578 ( .A(n12142), .B(n12141), .ZN(n12143) );
  AOI22_X1 U14579 ( .A1(n13368), .A2(n13336), .B1(n13337), .B2(n13370), .ZN(
        n13346) );
  OAI21_X1 U14580 ( .B1(n12143), .B2(n13623), .A(n13346), .ZN(n13644) );
  AOI211_X1 U14581 ( .C1(n15381), .C2(n13637), .A(n13645), .B(n13644), .ZN(
        n12149) );
  AOI22_X1 U14582 ( .A1(n13642), .A2(n12144), .B1(n15389), .B2(
        P2_REG1_REG_15__SCAN_IN), .ZN(n12145) );
  OAI21_X1 U14583 ( .B1(n12149), .B2(n15389), .A(n12145), .ZN(P2_U3514) );
  NOR2_X1 U14584 ( .A1(n15383), .A2(n8583), .ZN(n12146) );
  AOI21_X1 U14585 ( .B1(n13642), .B2(n12147), .A(n12146), .ZN(n12148) );
  OAI21_X1 U14586 ( .B1(n12149), .B2(n15382), .A(n12148), .ZN(P2_U3475) );
  XNOR2_X1 U14587 ( .A(n12150), .B(n12686), .ZN(n12151) );
  AOI222_X1 U14588 ( .A1(n13032), .A2(n12151), .B1(n12731), .B2(n13027), .C1(
        n12730), .C2(n13029), .ZN(n13100) );
  XNOR2_X1 U14589 ( .A(n12152), .B(n12686), .ZN(n13098) );
  NOR2_X1 U14590 ( .A1(n12510), .A2(n15442), .ZN(n12154) );
  INV_X1 U14591 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n12758) );
  OAI22_X1 U14592 ( .A1(n15464), .A2(n12758), .B1(n12502), .B2(n15440), .ZN(
        n12153) );
  AOI211_X1 U14593 ( .C1(n13098), .C2(n13039), .A(n12154), .B(n12153), .ZN(
        n12155) );
  OAI21_X1 U14594 ( .B1(n13100), .B2(n13024), .A(n12155), .ZN(P3_U3218) );
  XOR2_X1 U14595 ( .A(n12158), .B(n12156), .Z(n14863) );
  INV_X1 U14596 ( .A(n14863), .ZN(n12168) );
  OAI211_X1 U14597 ( .C1(n12159), .C2(n12158), .A(n13661), .B(n12157), .ZN(
        n14857) );
  OAI22_X1 U14598 ( .A1(n12161), .A2(n13301), .B1(n12160), .B2(n13303), .ZN(
        n14852) );
  INV_X1 U14599 ( .A(n14852), .ZN(n14858) );
  OAI211_X1 U14600 ( .C1(n13655), .C2(n14856), .A(n14857), .B(n14858), .ZN(
        n12166) );
  INV_X1 U14601 ( .A(n14853), .ZN(n14860) );
  INV_X1 U14602 ( .A(n12162), .ZN(n12163) );
  OAI211_X1 U14603 ( .C1(n14860), .C2(n12163), .A(n13604), .B(n6739), .ZN(
        n14859) );
  NOR2_X1 U14604 ( .A1(n14859), .A2(n13612), .ZN(n12165) );
  OAI22_X1 U14605 ( .A1(n14860), .A2(n15330), .B1(n11607), .B2(n13643), .ZN(
        n12164) );
  AOI211_X1 U14606 ( .C1(n12166), .C2(n13643), .A(n12165), .B(n12164), .ZN(
        n12167) );
  OAI21_X1 U14607 ( .B1(n12168), .B2(n13592), .A(n12167), .ZN(P2_U3249) );
  INV_X1 U14608 ( .A(n12169), .ZN(n12170) );
  OAI222_X1 U14609 ( .A1(n13798), .A2(n12171), .B1(n13804), .B2(n12170), .C1(
        P2_U3088), .C2(n9110), .ZN(P2_U3305) );
  INV_X1 U14610 ( .A(n13793), .ZN(n12172) );
  OAI222_X1 U14611 ( .A1(P1_U3086), .A2(n12173), .B1(n14761), .B2(n12172), 
        .C1(n14774), .C2(n9669), .ZN(P1_U3327) );
  NAND2_X1 U14612 ( .A1(n14910), .A2(n12300), .ZN(n12175) );
  NAND2_X1 U14613 ( .A1(n14221), .A2(n6622), .ZN(n12174) );
  NAND2_X1 U14614 ( .A1(n12175), .A2(n12174), .ZN(n12176) );
  XNOR2_X1 U14615 ( .A(n12176), .B(n12288), .ZN(n12185) );
  NOR2_X1 U14616 ( .A1(n12284), .A2(n12177), .ZN(n12178) );
  AOI21_X1 U14617 ( .B1(n14910), .B2(n6622), .A(n12178), .ZN(n12183) );
  XNOR2_X1 U14618 ( .A(n12185), .B(n12183), .ZN(n14901) );
  INV_X1 U14619 ( .A(n12179), .ZN(n12180) );
  NAND2_X1 U14620 ( .A1(n12181), .A2(n12180), .ZN(n14902) );
  INV_X1 U14621 ( .A(n12183), .ZN(n12184) );
  OR2_X1 U14622 ( .A1(n12185), .A2(n12184), .ZN(n12186) );
  NOR2_X1 U14623 ( .A1(n12284), .A2(n14898), .ZN(n12187) );
  AOI21_X1 U14624 ( .B1(n14040), .B2(n6622), .A(n12187), .ZN(n12192) );
  NAND2_X1 U14625 ( .A1(n14040), .A2(n12300), .ZN(n12189) );
  NAND2_X1 U14626 ( .A1(n14220), .A2(n6622), .ZN(n12188) );
  NAND2_X1 U14627 ( .A1(n12189), .A2(n12188), .ZN(n12190) );
  XNOR2_X1 U14628 ( .A(n12190), .B(n12208), .ZN(n12191) );
  XOR2_X1 U14629 ( .A(n12192), .B(n12191), .Z(n13859) );
  INV_X1 U14630 ( .A(n12191), .ZN(n12193) );
  NOR2_X1 U14631 ( .A1(n12193), .A2(n12192), .ZN(n12194) );
  NOR2_X1 U14632 ( .A1(n12284), .A2(n14887), .ZN(n12195) );
  AOI21_X1 U14633 ( .B1(n14043), .B2(n6622), .A(n12195), .ZN(n12202) );
  OAI22_X1 U14634 ( .A1(n14044), .A2(n12256), .B1(n14887), .B2(n11299), .ZN(
        n12196) );
  XNOR2_X1 U14635 ( .A(n12196), .B(n12208), .ZN(n12201) );
  XOR2_X1 U14636 ( .A(n12202), .B(n12201), .Z(n13901) );
  NAND2_X1 U14637 ( .A1(n14946), .A2(n12300), .ZN(n12198) );
  OR2_X1 U14638 ( .A1(n13904), .A2(n11299), .ZN(n12197) );
  NAND2_X1 U14639 ( .A1(n12198), .A2(n12197), .ZN(n12199) );
  XNOR2_X1 U14640 ( .A(n12199), .B(n12208), .ZN(n12205) );
  NOR2_X1 U14641 ( .A1(n12284), .A2(n13904), .ZN(n12200) );
  AOI21_X1 U14642 ( .B1(n14946), .B2(n6622), .A(n12200), .ZN(n12206) );
  XNOR2_X1 U14643 ( .A(n12205), .B(n12206), .ZN(n14888) );
  INV_X1 U14644 ( .A(n12201), .ZN(n12203) );
  OR2_X1 U14645 ( .A1(n12203), .A2(n12202), .ZN(n14889) );
  INV_X1 U14646 ( .A(n12205), .ZN(n12207) );
  AOI22_X1 U14647 ( .A1(n14590), .A2(n12300), .B1(n6622), .B2(n14567), .ZN(
        n12209) );
  XNOR2_X1 U14648 ( .A(n12209), .B(n12288), .ZN(n12210) );
  AOI22_X1 U14649 ( .A1(n14590), .A2(n6622), .B1(n12301), .B2(n14567), .ZN(
        n13941) );
  NAND2_X1 U14650 ( .A1(n13939), .A2(n13941), .ZN(n12212) );
  NAND2_X1 U14651 ( .A1(n12211), .A2(n12210), .ZN(n13940) );
  NAND2_X1 U14652 ( .A1(n12212), .A2(n13940), .ZN(n13871) );
  NAND2_X1 U14653 ( .A1(n14705), .A2(n12300), .ZN(n12214) );
  NAND2_X1 U14654 ( .A1(n14582), .A2(n6622), .ZN(n12213) );
  NAND2_X1 U14655 ( .A1(n12214), .A2(n12213), .ZN(n12215) );
  XNOR2_X1 U14656 ( .A(n12215), .B(n12288), .ZN(n12216) );
  AOI22_X1 U14657 ( .A1(n14705), .A2(n6622), .B1(n12301), .B2(n14582), .ZN(
        n12217) );
  XNOR2_X1 U14658 ( .A(n12216), .B(n12217), .ZN(n13872) );
  NAND2_X1 U14659 ( .A1(n13871), .A2(n13872), .ZN(n12220) );
  INV_X1 U14660 ( .A(n12216), .ZN(n12218) );
  NAND2_X1 U14661 ( .A1(n12218), .A2(n12217), .ZN(n12219) );
  NAND2_X1 U14662 ( .A1(n12220), .A2(n12219), .ZN(n13878) );
  OAI22_X1 U14663 ( .A1(n14556), .A2(n11299), .B1(n14063), .B2(n12284), .ZN(
        n12225) );
  NAND2_X1 U14664 ( .A1(n14698), .A2(n12300), .ZN(n12222) );
  OR2_X1 U14665 ( .A1(n14063), .A2(n11299), .ZN(n12221) );
  NAND2_X1 U14666 ( .A1(n12222), .A2(n12221), .ZN(n12223) );
  XNOR2_X1 U14667 ( .A(n12223), .B(n12288), .ZN(n12224) );
  XOR2_X1 U14668 ( .A(n12225), .B(n12224), .Z(n13879) );
  NAND2_X1 U14669 ( .A1(n13878), .A2(n13879), .ZN(n12229) );
  INV_X1 U14670 ( .A(n12224), .ZN(n12227) );
  INV_X1 U14671 ( .A(n12225), .ZN(n12226) );
  NAND2_X1 U14672 ( .A1(n12227), .A2(n12226), .ZN(n12228) );
  NAND2_X1 U14673 ( .A1(n12229), .A2(n12228), .ZN(n13923) );
  NAND2_X1 U14674 ( .A1(n14537), .A2(n12300), .ZN(n12231) );
  NAND2_X1 U14675 ( .A1(n6943), .A2(n6622), .ZN(n12230) );
  NAND2_X1 U14676 ( .A1(n12231), .A2(n12230), .ZN(n12232) );
  XNOR2_X1 U14677 ( .A(n12232), .B(n12288), .ZN(n12233) );
  AOI22_X1 U14678 ( .A1(n14537), .A2(n6622), .B1(n12301), .B2(n6943), .ZN(
        n12234) );
  XNOR2_X1 U14679 ( .A(n12233), .B(n12234), .ZN(n13924) );
  INV_X1 U14680 ( .A(n12233), .ZN(n12235) );
  NAND2_X1 U14681 ( .A1(n12235), .A2(n12234), .ZN(n12236) );
  AND2_X1 U14682 ( .A1(n14545), .A2(n12301), .ZN(n12237) );
  AOI21_X1 U14683 ( .B1(n14528), .B2(n6622), .A(n12237), .ZN(n12241) );
  NAND2_X1 U14684 ( .A1(n14528), .A2(n12300), .ZN(n12239) );
  NAND2_X1 U14685 ( .A1(n14545), .A2(n6622), .ZN(n12238) );
  NAND2_X1 U14686 ( .A1(n12239), .A2(n12238), .ZN(n12240) );
  XNOR2_X1 U14687 ( .A(n12240), .B(n12288), .ZN(n12243) );
  XOR2_X1 U14688 ( .A(n12241), .B(n12243), .Z(n13833) );
  INV_X1 U14689 ( .A(n12241), .ZN(n12242) );
  NAND2_X1 U14690 ( .A1(n12243), .A2(n12242), .ZN(n12244) );
  OAI22_X1 U14691 ( .A1(n14674), .A2(n11299), .B1(n14085), .B2(n12284), .ZN(
        n12246) );
  OAI22_X1 U14692 ( .A1(n14674), .A2(n12256), .B1(n14085), .B2(n11299), .ZN(
        n12245) );
  XNOR2_X1 U14693 ( .A(n12245), .B(n12288), .ZN(n12247) );
  XOR2_X1 U14694 ( .A(n12246), .B(n12247), .Z(n13894) );
  NAND2_X1 U14695 ( .A1(n12247), .A2(n12246), .ZN(n12248) );
  AOI22_X1 U14696 ( .A1(n14739), .A2(n12300), .B1(n6622), .B2(n14218), .ZN(
        n12249) );
  XNOR2_X1 U14697 ( .A(n12249), .B(n12288), .ZN(n12252) );
  AOI22_X1 U14698 ( .A1(n14739), .A2(n6622), .B1(n12301), .B2(n14218), .ZN(
        n12251) );
  XNOR2_X1 U14699 ( .A(n12252), .B(n12251), .ZN(n13846) );
  INV_X1 U14700 ( .A(n13846), .ZN(n12250) );
  NAND2_X1 U14701 ( .A1(n12252), .A2(n12251), .ZN(n12253) );
  OAI22_X1 U14702 ( .A1(n14738), .A2(n12256), .B1(n12255), .B2(n11299), .ZN(
        n12257) );
  XNOR2_X1 U14703 ( .A(n12257), .B(n12288), .ZN(n12259) );
  AND2_X1 U14704 ( .A1(n14217), .A2(n12301), .ZN(n12258) );
  AOI21_X1 U14705 ( .B1(n14481), .B2(n6622), .A(n12258), .ZN(n12260) );
  XNOR2_X1 U14706 ( .A(n12259), .B(n12260), .ZN(n13911) );
  INV_X1 U14707 ( .A(n12259), .ZN(n12261) );
  NAND2_X1 U14708 ( .A1(n12261), .A2(n12260), .ZN(n12262) );
  NAND2_X1 U14709 ( .A1(n14732), .A2(n12300), .ZN(n12264) );
  NAND2_X1 U14710 ( .A1(n14216), .A2(n6622), .ZN(n12263) );
  NAND2_X1 U14711 ( .A1(n12264), .A2(n12263), .ZN(n12265) );
  XNOR2_X1 U14712 ( .A(n12265), .B(n12288), .ZN(n12266) );
  AOI22_X1 U14713 ( .A1(n14732), .A2(n6622), .B1(n12301), .B2(n14216), .ZN(
        n12267) );
  XNOR2_X1 U14714 ( .A(n12266), .B(n12267), .ZN(n13817) );
  INV_X1 U14715 ( .A(n12266), .ZN(n12268) );
  NAND2_X1 U14716 ( .A1(n14728), .A2(n12300), .ZN(n12270) );
  NAND2_X1 U14717 ( .A1(n14215), .A2(n6622), .ZN(n12269) );
  NAND2_X1 U14718 ( .A1(n12270), .A2(n12269), .ZN(n12271) );
  XNOR2_X1 U14719 ( .A(n12271), .B(n12288), .ZN(n12272) );
  AOI22_X1 U14720 ( .A1(n14728), .A2(n6622), .B1(n12301), .B2(n14215), .ZN(
        n12273) );
  XNOR2_X1 U14721 ( .A(n12272), .B(n12273), .ZN(n13886) );
  NAND2_X1 U14722 ( .A1(n13885), .A2(n13886), .ZN(n12276) );
  INV_X1 U14723 ( .A(n12272), .ZN(n12274) );
  NAND2_X1 U14724 ( .A1(n12274), .A2(n12273), .ZN(n12275) );
  NAND2_X1 U14725 ( .A1(n14724), .A2(n12300), .ZN(n12278) );
  NAND2_X1 U14726 ( .A1(n14214), .A2(n6622), .ZN(n12277) );
  NAND2_X1 U14727 ( .A1(n12278), .A2(n12277), .ZN(n12279) );
  XNOR2_X1 U14728 ( .A(n12279), .B(n12288), .ZN(n12280) );
  AOI22_X1 U14729 ( .A1(n14724), .A2(n6622), .B1(n12301), .B2(n14214), .ZN(
        n12281) );
  XNOR2_X1 U14730 ( .A(n12280), .B(n12281), .ZN(n13864) );
  INV_X1 U14731 ( .A(n12280), .ZN(n12282) );
  NAND2_X1 U14732 ( .A1(n12282), .A2(n12281), .ZN(n12283) );
  OAI22_X1 U14733 ( .A1(n14639), .A2(n11299), .B1(n12285), .B2(n12284), .ZN(
        n12291) );
  NAND2_X1 U14734 ( .A1(n14419), .A2(n12300), .ZN(n12287) );
  NAND2_X1 U14735 ( .A1(n14213), .A2(n6622), .ZN(n12286) );
  NAND2_X1 U14736 ( .A1(n12287), .A2(n12286), .ZN(n12289) );
  XNOR2_X1 U14737 ( .A(n12289), .B(n12288), .ZN(n12290) );
  XOR2_X1 U14738 ( .A(n12291), .B(n12290), .Z(n13931) );
  INV_X1 U14739 ( .A(n12290), .ZN(n12293) );
  INV_X1 U14740 ( .A(n12291), .ZN(n12292) );
  NAND2_X1 U14741 ( .A1(n14629), .A2(n12300), .ZN(n12295) );
  NAND2_X1 U14742 ( .A1(n14377), .A2(n6622), .ZN(n12294) );
  NAND2_X1 U14743 ( .A1(n12295), .A2(n12294), .ZN(n12296) );
  XNOR2_X1 U14744 ( .A(n12296), .B(n12208), .ZN(n12297) );
  AOI22_X1 U14745 ( .A1(n14629), .A2(n6622), .B1(n12301), .B2(n14377), .ZN(
        n12298) );
  XNOR2_X1 U14746 ( .A(n12297), .B(n12298), .ZN(n13809) );
  INV_X1 U14747 ( .A(n12297), .ZN(n12299) );
  AOI21_X1 U14748 ( .B1(n13808), .B2(n13809), .A(n7570), .ZN(n12306) );
  AOI22_X1 U14749 ( .A1(n14627), .A2(n12300), .B1(n6622), .B2(n14125), .ZN(
        n12304) );
  AOI22_X1 U14750 ( .A1(n14627), .A2(n6622), .B1(n12301), .B2(n14125), .ZN(
        n12302) );
  XNOR2_X1 U14751 ( .A(n12302), .B(n12208), .ZN(n12303) );
  XOR2_X1 U14752 ( .A(n12304), .B(n12303), .Z(n12305) );
  XNOR2_X1 U14753 ( .A(n12306), .B(n12305), .ZN(n12311) );
  NOR2_X1 U14754 ( .A1(n14914), .A2(n14384), .ZN(n12309) );
  AOI22_X1 U14755 ( .A1(n13943), .A2(n14377), .B1(P1_REG3_REG_28__SCAN_IN), 
        .B2(P1_U3086), .ZN(n12307) );
  OAI21_X1 U14756 ( .B1(n14138), .B2(n14897), .A(n12307), .ZN(n12308) );
  AOI211_X1 U14757 ( .C1(n14627), .C2(n14909), .A(n12309), .B(n12308), .ZN(
        n12310) );
  OAI21_X1 U14758 ( .B1(n12311), .B2(n14904), .A(n12310), .ZN(P1_U3220) );
  INV_X1 U14759 ( .A(n12312), .ZN(n12327) );
  INV_X1 U14760 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n12316) );
  OAI222_X1 U14761 ( .A1(n13804), .A2(n14760), .B1(n8368), .B2(P2_U3088), .C1(
        n12316), .C2(n13798), .ZN(P2_U3297) );
  INV_X1 U14762 ( .A(SI_31_), .ZN(n12663) );
  INV_X1 U14763 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n14759) );
  AOI22_X1 U14764 ( .A1(P2_DATAO_REG_30__SCAN_IN), .A2(
        P1_DATAO_REG_30__SCAN_IN), .B1(n12316), .B2(n14759), .ZN(n12658) );
  INV_X1 U14765 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n14753) );
  AOI22_X1 U14766 ( .A1(P1_DATAO_REG_31__SCAN_IN), .A2(n14753), .B1(
        P2_DATAO_REG_31__SCAN_IN), .B2(n12317), .ZN(n12318) );
  XNOR2_X1 U14767 ( .A(n12319), .B(n12318), .ZN(n12664) );
  NAND2_X1 U14768 ( .A1(n12664), .A2(n14796), .ZN(n12324) );
  INV_X1 U14769 ( .A(n12320), .ZN(n12322) );
  OR4_X1 U14770 ( .A1(n12322), .A2(P3_IR_REG_30__SCAN_IN), .A3(n12321), .A4(
        P3_U3151), .ZN(n12323) );
  OAI211_X1 U14771 ( .C1(n12663), .C2(n13167), .A(n12324), .B(n12323), .ZN(
        P3_U3264) );
  OAI222_X1 U14772 ( .A1(n13804), .A2(n12327), .B1(n12326), .B2(P2_U3088), 
        .C1(n12325), .C2(n13798), .ZN(P2_U3307) );
  INV_X1 U14773 ( .A(n12329), .ZN(n12330) );
  NAND2_X1 U14774 ( .A1(n12330), .A2(n15463), .ZN(n12852) );
  NAND2_X1 U14775 ( .A1(n13024), .A2(P3_REG2_REG_29__SCAN_IN), .ZN(n12331) );
  OAI211_X1 U14776 ( .C1(n12332), .C2(n15442), .A(n12852), .B(n12331), .ZN(
        n12333) );
  AOI21_X1 U14777 ( .B1(n12334), .B2(n13039), .A(n12333), .ZN(n12335) );
  OAI21_X1 U14778 ( .B1(n12328), .B2(n13024), .A(n12335), .ZN(P3_U3204) );
  XNOR2_X1 U14779 ( .A(n13111), .B(n12392), .ZN(n12388) );
  XNOR2_X1 U14780 ( .A(n12388), .B(n12891), .ZN(n12390) );
  INV_X1 U14781 ( .A(n12336), .ZN(n12337) );
  NAND2_X1 U14782 ( .A1(n12337), .A2(n12731), .ZN(n12338) );
  NAND2_X1 U14783 ( .A1(n12339), .A2(n12338), .ZN(n12499) );
  XNOR2_X1 U14784 ( .A(n12510), .B(n12392), .ZN(n12340) );
  XNOR2_X1 U14785 ( .A(n12340), .B(n12599), .ZN(n12498) );
  NAND2_X1 U14786 ( .A1(n12340), .A2(n13028), .ZN(n12341) );
  NAND2_X1 U14787 ( .A1(n12497), .A2(n12341), .ZN(n12436) );
  XNOR2_X1 U14788 ( .A(n13093), .B(n12392), .ZN(n12342) );
  XNOR2_X1 U14789 ( .A(n12342), .B(n12730), .ZN(n12435) );
  NAND2_X1 U14790 ( .A1(n12436), .A2(n12435), .ZN(n12434) );
  INV_X1 U14791 ( .A(n12342), .ZN(n12343) );
  NAND2_X1 U14792 ( .A1(n12343), .A2(n12730), .ZN(n12344) );
  NAND2_X1 U14793 ( .A1(n12434), .A2(n12344), .ZN(n12443) );
  XNOR2_X1 U14794 ( .A(n12445), .B(n6818), .ZN(n12345) );
  XNOR2_X1 U14795 ( .A(n12345), .B(n12478), .ZN(n12442) );
  NAND2_X1 U14796 ( .A1(n13030), .A2(n12345), .ZN(n12346) );
  NAND2_X1 U14797 ( .A1(n12441), .A2(n12346), .ZN(n12477) );
  XNOR2_X1 U14798 ( .A(n13009), .B(n6818), .ZN(n12347) );
  XNOR2_X1 U14799 ( .A(n12347), .B(n13017), .ZN(n12476) );
  NAND2_X1 U14800 ( .A1(n12477), .A2(n12476), .ZN(n12475) );
  INV_X1 U14801 ( .A(n13017), .ZN(n12990) );
  NAND2_X1 U14802 ( .A1(n12347), .A2(n12990), .ZN(n12348) );
  NAND2_X1 U14803 ( .A1(n12475), .A2(n12348), .ZN(n12383) );
  XNOR2_X1 U14804 ( .A(n13139), .B(n6818), .ZN(n12349) );
  XNOR2_X1 U14805 ( .A(n12349), .B(n13003), .ZN(n12382) );
  INV_X1 U14806 ( .A(n12349), .ZN(n12350) );
  NAND2_X1 U14807 ( .A1(n12350), .A2(n13003), .ZN(n12351) );
  XNOR2_X1 U14808 ( .A(n12982), .B(n12392), .ZN(n12352) );
  XNOR2_X1 U14809 ( .A(n12352), .B(n12989), .ZN(n12462) );
  INV_X1 U14810 ( .A(n12352), .ZN(n12353) );
  NAND2_X1 U14811 ( .A1(n12353), .A2(n12989), .ZN(n12354) );
  XNOR2_X1 U14812 ( .A(n13134), .B(n12392), .ZN(n12355) );
  XNOR2_X1 U14813 ( .A(n12355), .B(n12954), .ZN(n12403) );
  XNOR2_X1 U14814 ( .A(n12958), .B(n12392), .ZN(n12356) );
  INV_X1 U14815 ( .A(n12356), .ZN(n12357) );
  NOR2_X1 U14816 ( .A1(n12358), .A2(n12357), .ZN(n12359) );
  XNOR2_X1 U14817 ( .A(n13122), .B(n6818), .ZN(n12452) );
  XNOR2_X1 U14818 ( .A(n13126), .B(n6818), .ZN(n12361) );
  OAI22_X1 U14819 ( .A1(n12452), .A2(n12451), .B1(n12955), .B2(n12361), .ZN(
        n12365) );
  OAI21_X1 U14820 ( .B1(n12448), .B2(n12729), .A(n12941), .ZN(n12363) );
  NOR3_X1 U14821 ( .A1(n12448), .A2(n12729), .A3(n12941), .ZN(n12362) );
  AOI21_X1 U14822 ( .B1(n12452), .B2(n12363), .A(n12362), .ZN(n12364) );
  XNOR2_X1 U14823 ( .A(n12908), .B(n12392), .ZN(n12366) );
  XNOR2_X1 U14824 ( .A(n12366), .B(n12728), .ZN(n12428) );
  XNOR2_X1 U14825 ( .A(n12492), .B(n12392), .ZN(n12367) );
  XNOR2_X1 U14826 ( .A(n12367), .B(n12876), .ZN(n12484) );
  INV_X1 U14827 ( .A(n12367), .ZN(n12368) );
  XOR2_X1 U14828 ( .A(n12390), .B(n12391), .Z(n12375) );
  OAI22_X1 U14829 ( .A1(n12876), .A2(n12500), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12369), .ZN(n12371) );
  NOR2_X1 U14830 ( .A1(n12877), .A2(n12489), .ZN(n12370) );
  AOI211_X1 U14831 ( .C1(n12881), .C2(n12486), .A(n12371), .B(n12370), .ZN(
        n12374) );
  NAND2_X1 U14832 ( .A1(n12372), .A2(n12491), .ZN(n12373) );
  OAI211_X1 U14833 ( .C1(n12375), .C2(n12494), .A(n12374), .B(n12373), .ZN(
        P3_U3154) );
  XNOR2_X1 U14834 ( .A(n12450), .B(n12955), .ZN(n12380) );
  AOI22_X1 U14835 ( .A1(n12485), .A2(n12940), .B1(P3_REG3_REG_23__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12377) );
  NAND2_X1 U14836 ( .A1(n12486), .A2(n12945), .ZN(n12376) );
  OAI211_X1 U14837 ( .C1(n12451), .C2(n12489), .A(n12377), .B(n12376), .ZN(
        n12378) );
  AOI21_X1 U14838 ( .B1(n12949), .B2(n12491), .A(n12378), .ZN(n12379) );
  OAI21_X1 U14839 ( .B1(n12380), .B2(n12494), .A(n12379), .ZN(P3_U3156) );
  OAI211_X1 U14840 ( .C1(n12383), .C2(n12382), .A(n12381), .B(n12496), .ZN(
        n12387) );
  NAND2_X1 U14841 ( .A1(P3_U3151), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n12839)
         );
  OAI21_X1 U14842 ( .B1(n13017), .B2(n12500), .A(n12839), .ZN(n12385) );
  NOR2_X1 U14843 ( .A1(n12503), .A2(n12996), .ZN(n12384) );
  AOI211_X1 U14844 ( .C1(n12506), .C2(n12989), .A(n12385), .B(n12384), .ZN(
        n12386) );
  OAI211_X1 U14845 ( .C1(n12509), .C2(n13139), .A(n12387), .B(n12386), .ZN(
        P3_U3159) );
  INV_X1 U14846 ( .A(n12388), .ZN(n12389) );
  XNOR2_X1 U14847 ( .A(n12863), .B(n12392), .ZN(n12393) );
  XNOR2_X1 U14848 ( .A(n12394), .B(n12393), .ZN(n12401) );
  NOR2_X1 U14849 ( .A1(n12859), .A2(n12489), .ZN(n12397) );
  OAI22_X1 U14850 ( .A1(n12891), .A2(n12500), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12395), .ZN(n12396) );
  AOI211_X1 U14851 ( .C1(n12864), .C2(n12486), .A(n12397), .B(n12396), .ZN(
        n12400) );
  NAND2_X1 U14852 ( .A1(n12398), .A2(n12491), .ZN(n12399) );
  OAI211_X1 U14853 ( .C1(n12401), .C2(n12494), .A(n12400), .B(n12399), .ZN(
        P3_U3160) );
  OAI211_X1 U14854 ( .C1(n12404), .C2(n12403), .A(n12402), .B(n12496), .ZN(
        n12408) );
  AOI22_X1 U14855 ( .A1(n12989), .A2(n12485), .B1(P3_REG3_REG_21__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12405) );
  OAI21_X1 U14856 ( .B1(n12967), .B2(n12489), .A(n12405), .ZN(n12406) );
  AOI21_X1 U14857 ( .B1(n12970), .B2(n12486), .A(n12406), .ZN(n12407) );
  OAI211_X1 U14858 ( .C1(n13134), .C2(n12509), .A(n12408), .B(n12407), .ZN(
        P3_U3163) );
  AOI21_X1 U14859 ( .B1(n12411), .B2(n12410), .A(n12409), .ZN(n12414) );
  XNOR2_X1 U14860 ( .A(n12732), .B(n12412), .ZN(n12413) );
  XNOR2_X1 U14861 ( .A(n12414), .B(n12413), .ZN(n12425) );
  AOI21_X1 U14862 ( .B1(n12416), .B2(n12485), .A(n12415), .ZN(n12423) );
  NAND2_X1 U14863 ( .A1(n12491), .A2(n12417), .ZN(n12422) );
  NAND2_X1 U14864 ( .A1(n12486), .A2(n12418), .ZN(n12421) );
  NAND2_X1 U14865 ( .A1(n12506), .A2(n12419), .ZN(n12420) );
  NAND4_X1 U14866 ( .A1(n12423), .A2(n12422), .A3(n12421), .A4(n12420), .ZN(
        n12424) );
  AOI21_X1 U14867 ( .B1(n12425), .B2(n12496), .A(n12424), .ZN(n12426) );
  INV_X1 U14868 ( .A(n12426), .ZN(P3_U3164) );
  XOR2_X1 U14869 ( .A(n12428), .B(n12427), .Z(n12433) );
  AOI22_X1 U14870 ( .A1(n12941), .A2(n12485), .B1(P3_REG3_REG_25__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12430) );
  NAND2_X1 U14871 ( .A1(n12486), .A2(n12909), .ZN(n12429) );
  OAI211_X1 U14872 ( .C1(n12876), .C2(n12489), .A(n12430), .B(n12429), .ZN(
        n12431) );
  AOI21_X1 U14873 ( .B1(n12908), .B2(n12491), .A(n12431), .ZN(n12432) );
  OAI21_X1 U14874 ( .B1(n12433), .B2(n12494), .A(n12432), .ZN(P3_U3165) );
  OAI211_X1 U14875 ( .C1(n12436), .C2(n12435), .A(n12434), .B(n12496), .ZN(
        n12440) );
  NAND2_X1 U14876 ( .A1(P3_U3151), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n12769)
         );
  OAI21_X1 U14877 ( .B1(n12599), .B2(n12500), .A(n12769), .ZN(n12438) );
  NOR2_X1 U14878 ( .A1(n12503), .A2(n13036), .ZN(n12437) );
  AOI211_X1 U14879 ( .C1(n12506), .C2(n13030), .A(n12438), .B(n12437), .ZN(
        n12439) );
  OAI211_X1 U14880 ( .C1(n13035), .C2(n12509), .A(n12440), .B(n12439), .ZN(
        P3_U3166) );
  OAI211_X1 U14881 ( .C1(n12443), .C2(n12442), .A(n12441), .B(n12496), .ZN(
        n12447) );
  AND2_X1 U14882 ( .A1(P3_U3151), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n12797) );
  OAI22_X1 U14883 ( .A1(n13016), .A2(n12500), .B1(n13017), .B2(n12489), .ZN(
        n12444) );
  AOI211_X1 U14884 ( .C1(n12445), .C2(n12491), .A(n12797), .B(n12444), .ZN(
        n12446) );
  OAI211_X1 U14885 ( .C1(n13018), .C2(n12503), .A(n12447), .B(n12446), .ZN(
        P3_U3168) );
  OAI22_X1 U14886 ( .A1(n12450), .A2(n12729), .B1(n12449), .B2(n12448), .ZN(
        n12454) );
  XNOR2_X1 U14887 ( .A(n12452), .B(n12451), .ZN(n12453) );
  XNOR2_X1 U14888 ( .A(n12454), .B(n12453), .ZN(n12460) );
  AOI22_X1 U14889 ( .A1(n12485), .A2(n12729), .B1(P3_REG3_REG_24__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12456) );
  NAND2_X1 U14890 ( .A1(n12486), .A2(n12924), .ZN(n12455) );
  OAI211_X1 U14891 ( .C1(n12920), .C2(n12489), .A(n12456), .B(n12455), .ZN(
        n12457) );
  AOI21_X1 U14892 ( .B1(n12458), .B2(n12491), .A(n12457), .ZN(n12459) );
  OAI21_X1 U14893 ( .B1(n12460), .B2(n12494), .A(n12459), .ZN(P3_U3169) );
  OAI211_X1 U14894 ( .C1(n6784), .C2(n12462), .A(n12461), .B(n12496), .ZN(
        n12468) );
  INV_X1 U14895 ( .A(n12979), .ZN(n12466) );
  AOI22_X1 U14896 ( .A1(n12485), .A2(n13003), .B1(P3_REG3_REG_20__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12464) );
  OAI21_X1 U14897 ( .B1(n12954), .B2(n12489), .A(n12464), .ZN(n12465) );
  AOI21_X1 U14898 ( .B1(n12466), .B2(n12486), .A(n12465), .ZN(n12467) );
  OAI211_X1 U14899 ( .C1(n13078), .C2(n12509), .A(n12468), .B(n12467), .ZN(
        P3_U3173) );
  XNOR2_X1 U14900 ( .A(n12469), .B(n12940), .ZN(n12474) );
  AOI22_X1 U14901 ( .A1(n12977), .A2(n12485), .B1(P3_REG3_REG_22__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12471) );
  NAND2_X1 U14902 ( .A1(n12486), .A2(n12959), .ZN(n12470) );
  OAI211_X1 U14903 ( .C1(n12955), .C2(n12489), .A(n12471), .B(n12470), .ZN(
        n12472) );
  AOI21_X1 U14904 ( .B1(n12958), .B2(n12491), .A(n12472), .ZN(n12473) );
  OAI21_X1 U14905 ( .B1(n12474), .B2(n12494), .A(n12473), .ZN(P3_U3175) );
  OAI211_X1 U14906 ( .C1(n12477), .C2(n12476), .A(n12475), .B(n12496), .ZN(
        n12482) );
  NAND2_X1 U14907 ( .A1(P3_U3151), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n12823)
         );
  OAI21_X1 U14908 ( .B1(n12478), .B2(n12500), .A(n12823), .ZN(n12480) );
  NOR2_X1 U14909 ( .A1(n12503), .A2(n13005), .ZN(n12479) );
  AOI211_X1 U14910 ( .C1(n12506), .C2(n13003), .A(n12480), .B(n12479), .ZN(
        n12481) );
  OAI211_X1 U14911 ( .C1(n13087), .C2(n12509), .A(n12482), .B(n12481), .ZN(
        P3_U3178) );
  XOR2_X1 U14912 ( .A(n12484), .B(n12483), .Z(n12495) );
  AOI22_X1 U14913 ( .A1(n12728), .A2(n12485), .B1(P3_REG3_REG_26__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12488) );
  NAND2_X1 U14914 ( .A1(n12895), .A2(n12486), .ZN(n12487) );
  OAI211_X1 U14915 ( .C1(n12891), .C2(n12489), .A(n12488), .B(n12487), .ZN(
        n12490) );
  AOI21_X1 U14916 ( .B1(n12492), .B2(n12491), .A(n12490), .ZN(n12493) );
  OAI21_X1 U14917 ( .B1(n12495), .B2(n12494), .A(n12493), .ZN(P3_U3180) );
  OAI211_X1 U14918 ( .C1(n12499), .C2(n12498), .A(n12497), .B(n12496), .ZN(
        n12508) );
  NAND2_X1 U14919 ( .A1(P3_U3151), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n12748)
         );
  OAI21_X1 U14920 ( .B1(n12501), .B2(n12500), .A(n12748), .ZN(n12505) );
  NOR2_X1 U14921 ( .A1(n12503), .A2(n12502), .ZN(n12504) );
  AOI211_X1 U14922 ( .C1(n12506), .C2(n12730), .A(n12505), .B(n12504), .ZN(
        n12507) );
  OAI211_X1 U14923 ( .C1(n12510), .C2(n12509), .A(n12508), .B(n12507), .ZN(
        P3_U3181) );
  NAND2_X1 U14924 ( .A1(n12863), .A2(n12872), .ZN(n12700) );
  NAND2_X1 U14925 ( .A1(n6663), .A2(n12641), .ZN(n12888) );
  MUX2_X1 U14926 ( .A(n12512), .B(n12511), .S(n12653), .Z(n12640) );
  INV_X1 U14927 ( .A(n12513), .ZN(n12514) );
  NAND2_X1 U14928 ( .A1(n12517), .A2(n12514), .ZN(n12516) );
  NAND2_X1 U14929 ( .A1(n12516), .A2(n12515), .ZN(n12519) );
  INV_X1 U14930 ( .A(n12517), .ZN(n12518) );
  MUX2_X1 U14931 ( .A(n12519), .B(n12518), .S(n12647), .Z(n12520) );
  INV_X1 U14932 ( .A(n12520), .ZN(n12638) );
  MUX2_X1 U14933 ( .A(n12521), .B(n12522), .S(n12647), .Z(n12633) );
  INV_X1 U14934 ( .A(n12523), .ZN(n12525) );
  OAI21_X1 U14935 ( .B1(n11016), .B2(n12526), .A(n12530), .ZN(n12524) );
  MUX2_X1 U14936 ( .A(n12525), .B(n12524), .S(n12647), .Z(n12540) );
  INV_X1 U14937 ( .A(n12526), .ZN(n12527) );
  OAI22_X1 U14938 ( .A1(n12529), .A2(n12528), .B1(n12722), .B2(n12527), .ZN(
        n12531) );
  NAND2_X1 U14939 ( .A1(n12531), .A2(n12530), .ZN(n12532) );
  NAND2_X1 U14940 ( .A1(n12532), .A2(n15448), .ZN(n12539) );
  NAND2_X1 U14941 ( .A1(n12542), .A2(n12533), .ZN(n12536) );
  NAND2_X1 U14942 ( .A1(n12541), .A2(n12534), .ZN(n12535) );
  MUX2_X1 U14943 ( .A(n12536), .B(n12535), .S(n12647), .Z(n12537) );
  INV_X1 U14944 ( .A(n12537), .ZN(n12538) );
  OAI21_X1 U14945 ( .B1(n12540), .B2(n12539), .A(n12538), .ZN(n12544) );
  MUX2_X1 U14946 ( .A(n12542), .B(n12541), .S(n12653), .Z(n12543) );
  NAND3_X1 U14947 ( .A1(n12544), .A2(n12670), .A3(n12543), .ZN(n12548) );
  MUX2_X1 U14948 ( .A(n12546), .B(n12545), .S(n12647), .Z(n12547) );
  NAND3_X1 U14949 ( .A1(n12548), .A2(n12672), .A3(n12547), .ZN(n12553) );
  NAND2_X1 U14950 ( .A1(n12556), .A2(n12549), .ZN(n12550) );
  NAND2_X1 U14951 ( .A1(n12550), .A2(n12647), .ZN(n12552) );
  INV_X1 U14952 ( .A(n12555), .ZN(n12551) );
  AOI21_X1 U14953 ( .B1(n12553), .B2(n12552), .A(n12551), .ZN(n12560) );
  AOI21_X1 U14954 ( .B1(n12555), .B2(n12554), .A(n12647), .ZN(n12559) );
  INV_X1 U14955 ( .A(n12556), .ZN(n12557) );
  NAND2_X1 U14956 ( .A1(n12557), .A2(n12653), .ZN(n12558) );
  OAI211_X1 U14957 ( .C1(n12560), .C2(n12559), .A(n12673), .B(n12558), .ZN(
        n12564) );
  MUX2_X1 U14958 ( .A(n12562), .B(n12561), .S(n12647), .Z(n12563) );
  NAND3_X1 U14959 ( .A1(n12564), .A2(n12671), .A3(n12563), .ZN(n12569) );
  MUX2_X1 U14960 ( .A(n12567), .B(n12566), .S(n12647), .Z(n12568) );
  NAND3_X1 U14961 ( .A1(n12569), .A2(n7472), .A3(n12568), .ZN(n12573) );
  OR2_X1 U14962 ( .A1(n15485), .A2(n12653), .ZN(n12571) );
  NAND2_X1 U14963 ( .A1(n15485), .A2(n12653), .ZN(n12570) );
  MUX2_X1 U14964 ( .A(n12571), .B(n12570), .S(n12734), .Z(n12572) );
  NAND3_X1 U14965 ( .A1(n12573), .A2(n12669), .A3(n12572), .ZN(n12576) );
  NAND3_X1 U14966 ( .A1(n12733), .A2(n12647), .A3(n12574), .ZN(n12575) );
  NAND2_X1 U14967 ( .A1(n12576), .A2(n12575), .ZN(n12577) );
  NAND2_X1 U14968 ( .A1(n12577), .A2(n12682), .ZN(n12584) );
  NAND2_X1 U14969 ( .A1(n12682), .A2(n7406), .ZN(n12580) );
  NAND3_X1 U14970 ( .A1(n12580), .A2(n12587), .A3(n12579), .ZN(n12581) );
  NAND2_X1 U14971 ( .A1(n12581), .A2(n12653), .ZN(n12583) );
  INV_X1 U14972 ( .A(n12586), .ZN(n12582) );
  AOI21_X1 U14973 ( .B1(n12584), .B2(n12583), .A(n12582), .ZN(n12589) );
  AOI21_X1 U14974 ( .B1(n12586), .B2(n12585), .A(n12653), .ZN(n12588) );
  OAI22_X1 U14975 ( .A1(n12589), .A2(n12588), .B1(n12587), .B2(n12653), .ZN(
        n12590) );
  NAND2_X1 U14976 ( .A1(n12590), .A2(n7481), .ZN(n12594) );
  MUX2_X1 U14977 ( .A(n12592), .B(n12591), .S(n12653), .Z(n12593) );
  NAND3_X1 U14978 ( .A1(n12594), .A2(n12688), .A3(n12593), .ZN(n12598) );
  MUX2_X1 U14979 ( .A(n12596), .B(n12595), .S(n12647), .Z(n12597) );
  NAND3_X1 U14980 ( .A1(n12598), .A2(n12686), .A3(n12597), .ZN(n12602) );
  OAI22_X1 U14981 ( .A1(n13093), .A2(n13016), .B1(n12599), .B2(n13097), .ZN(
        n12600) );
  NAND2_X1 U14982 ( .A1(n12600), .A2(n12653), .ZN(n12601) );
  AOI21_X1 U14983 ( .B1(n12602), .B2(n12601), .A(n7413), .ZN(n12607) );
  AOI21_X1 U14984 ( .B1(n12604), .B2(n12603), .A(n12653), .ZN(n12606) );
  NAND2_X1 U14985 ( .A1(n12730), .A2(n12647), .ZN(n12605) );
  OAI22_X1 U14986 ( .A1(n12607), .A2(n12606), .B1(n13093), .B2(n12605), .ZN(
        n12614) );
  INV_X1 U14987 ( .A(n12608), .ZN(n12613) );
  INV_X1 U14988 ( .A(n12609), .ZN(n12610) );
  AOI21_X1 U14989 ( .B1(n12615), .B2(n12610), .A(n12653), .ZN(n12611) );
  NAND2_X1 U14990 ( .A1(n12612), .A2(n12611), .ZN(n12617) );
  AOI22_X1 U14991 ( .A1(n12614), .A2(n13020), .B1(n12613), .B2(n12617), .ZN(
        n12619) );
  NAND3_X1 U14992 ( .A1(n12621), .A2(n12615), .A3(n12653), .ZN(n12616) );
  NAND2_X1 U14993 ( .A1(n12617), .A2(n12616), .ZN(n12618) );
  OAI21_X1 U14994 ( .B1(n12619), .B2(n9517), .A(n12618), .ZN(n12623) );
  INV_X1 U14995 ( .A(n12983), .ZN(n12976) );
  MUX2_X1 U14996 ( .A(n12621), .B(n12620), .S(n12653), .Z(n12622) );
  NAND3_X1 U14997 ( .A1(n12623), .A2(n12976), .A3(n12622), .ZN(n12627) );
  XNOR2_X1 U14998 ( .A(n13134), .B(n12954), .ZN(n12968) );
  NAND2_X1 U14999 ( .A1(n13078), .A2(n12647), .ZN(n12625) );
  NAND2_X1 U15000 ( .A1(n12982), .A2(n12653), .ZN(n12624) );
  MUX2_X1 U15001 ( .A(n12625), .B(n12624), .S(n12966), .Z(n12626) );
  NAND3_X1 U15002 ( .A1(n12627), .A2(n12968), .A3(n12626), .ZN(n12631) );
  NAND3_X1 U15003 ( .A1(n13134), .A2(n12977), .A3(n12653), .ZN(n12630) );
  NAND3_X1 U15004 ( .A1(n12628), .A2(n12954), .A3(n12647), .ZN(n12629) );
  NAND4_X1 U15005 ( .A1(n12956), .A2(n12631), .A3(n12630), .A4(n12629), .ZN(
        n12632) );
  NAND3_X1 U15006 ( .A1(n12633), .A2(n12937), .A3(n12632), .ZN(n12635) );
  NAND3_X1 U15007 ( .A1(n12949), .A2(n12955), .A3(n12647), .ZN(n12634) );
  NAND2_X1 U15008 ( .A1(n12635), .A2(n12634), .ZN(n12636) );
  NAND2_X1 U15009 ( .A1(n12918), .A2(n12636), .ZN(n12637) );
  NAND3_X1 U15010 ( .A1(n12902), .A2(n12638), .A3(n12637), .ZN(n12639) );
  NAND2_X1 U15011 ( .A1(n12640), .A2(n12639), .ZN(n12643) );
  MUX2_X1 U15012 ( .A(n12641), .B(n6663), .S(n12647), .Z(n12642) );
  OAI21_X1 U15013 ( .B1(n12888), .B2(n12643), .A(n12642), .ZN(n12644) );
  INV_X1 U15014 ( .A(n12644), .ZN(n12645) );
  INV_X1 U15015 ( .A(n12651), .ZN(n12657) );
  NAND3_X1 U15016 ( .A1(n12650), .A2(n12647), .A3(n12646), .ZN(n12649) );
  AND2_X1 U15017 ( .A1(n12649), .A2(n12648), .ZN(n12656) );
  OAI21_X1 U15018 ( .B1(n7030), .B2(n12652), .A(n12651), .ZN(n12654) );
  NAND2_X1 U15019 ( .A1(n12654), .A2(n12653), .ZN(n12655) );
  INV_X1 U15020 ( .A(SI_30_), .ZN(n13155) );
  NAND2_X1 U15021 ( .A1(n14820), .A2(n12666), .ZN(n12696) );
  NAND2_X1 U15022 ( .A1(n12696), .A2(n12660), .ZN(n12709) );
  INV_X1 U15023 ( .A(n12709), .ZN(n12661) );
  NAND2_X1 U15024 ( .A1(n12662), .A2(n12661), .ZN(n12668) );
  INV_X1 U15025 ( .A(n12851), .ZN(n12665) );
  INV_X1 U15026 ( .A(n12666), .ZN(n12727) );
  INV_X1 U15027 ( .A(n12711), .ZN(n12698) );
  AND2_X1 U15028 ( .A1(n12710), .A2(n12698), .ZN(n12667) );
  NAND2_X1 U15029 ( .A1(n12854), .A2(n12851), .ZN(n12708) );
  INV_X1 U15030 ( .A(n12708), .ZN(n12701) );
  NAND3_X1 U15031 ( .A1(n15448), .A2(n12670), .A3(n12669), .ZN(n12675) );
  NAND4_X1 U15032 ( .A1(n12673), .A2(n13020), .A3(n12672), .A4(n12671), .ZN(
        n12674) );
  NOR2_X1 U15033 ( .A1(n12675), .A2(n12674), .ZN(n12683) );
  NOR2_X1 U15034 ( .A1(n12676), .A2(n11016), .ZN(n12679) );
  AND4_X1 U15035 ( .A1(n12679), .A2(n12678), .A3(n12677), .A4(n7472), .ZN(
        n12680) );
  NAND4_X1 U15036 ( .A1(n12683), .A2(n12682), .A3(n12681), .A4(n12680), .ZN(
        n12684) );
  NOR2_X1 U15037 ( .A1(n12685), .A2(n12684), .ZN(n12687) );
  AND4_X1 U15038 ( .A1(n13033), .A2(n12688), .A3(n12687), .A4(n12686), .ZN(
        n12689) );
  AND4_X1 U15039 ( .A1(n12968), .A2(n12995), .A3(n12690), .A4(n12689), .ZN(
        n12691) );
  AND4_X1 U15040 ( .A1(n12937), .A2(n12956), .A3(n12691), .A4(n12976), .ZN(
        n12692) );
  NAND3_X1 U15041 ( .A1(n12902), .A2(n12692), .A3(n12918), .ZN(n12693) );
  NAND3_X1 U15042 ( .A1(n12698), .A2(n12697), .A3(n12696), .ZN(n12699) );
  INV_X1 U15043 ( .A(n12715), .ZN(n12716) );
  NAND2_X1 U15044 ( .A1(n12717), .A2(n12716), .ZN(n12718) );
  NOR3_X1 U15045 ( .A1(n12721), .A2(n12720), .A3(n13162), .ZN(n12724) );
  OAI21_X1 U15046 ( .B1(n12722), .B2(n12725), .A(P3_B_REG_SCAN_IN), .ZN(n12723) );
  OAI22_X1 U15047 ( .A1(n12726), .A2(n12725), .B1(n12724), .B2(n12723), .ZN(
        P3_U3296) );
  MUX2_X1 U15048 ( .A(n12727), .B(P3_DATAO_REG_30__SCAN_IN), .S(n12740), .Z(
        P3_U3521) );
  MUX2_X1 U15049 ( .A(n12904), .B(P3_DATAO_REG_26__SCAN_IN), .S(n12740), .Z(
        P3_U3517) );
  MUX2_X1 U15050 ( .A(n12728), .B(P3_DATAO_REG_25__SCAN_IN), .S(n12740), .Z(
        P3_U3516) );
  MUX2_X1 U15051 ( .A(n12941), .B(P3_DATAO_REG_24__SCAN_IN), .S(n12740), .Z(
        P3_U3515) );
  MUX2_X1 U15052 ( .A(n12729), .B(P3_DATAO_REG_23__SCAN_IN), .S(n12740), .Z(
        P3_U3514) );
  MUX2_X1 U15053 ( .A(n12940), .B(P3_DATAO_REG_22__SCAN_IN), .S(n12740), .Z(
        P3_U3513) );
  MUX2_X1 U15054 ( .A(P3_DATAO_REG_21__SCAN_IN), .B(n12977), .S(P3_U3897), .Z(
        P3_U3512) );
  MUX2_X1 U15055 ( .A(n12989), .B(P3_DATAO_REG_20__SCAN_IN), .S(n12740), .Z(
        P3_U3511) );
  MUX2_X1 U15056 ( .A(n13003), .B(P3_DATAO_REG_19__SCAN_IN), .S(n12740), .Z(
        P3_U3510) );
  MUX2_X1 U15057 ( .A(n12990), .B(P3_DATAO_REG_18__SCAN_IN), .S(n12740), .Z(
        P3_U3509) );
  MUX2_X1 U15058 ( .A(n13030), .B(P3_DATAO_REG_17__SCAN_IN), .S(n12740), .Z(
        P3_U3508) );
  MUX2_X1 U15059 ( .A(n12730), .B(P3_DATAO_REG_16__SCAN_IN), .S(n12740), .Z(
        P3_U3507) );
  MUX2_X1 U15060 ( .A(n13028), .B(P3_DATAO_REG_15__SCAN_IN), .S(n12740), .Z(
        P3_U3506) );
  MUX2_X1 U15061 ( .A(n12731), .B(P3_DATAO_REG_14__SCAN_IN), .S(n12740), .Z(
        P3_U3505) );
  MUX2_X1 U15062 ( .A(n12732), .B(P3_DATAO_REG_12__SCAN_IN), .S(n12740), .Z(
        P3_U3503) );
  MUX2_X1 U15063 ( .A(n12733), .B(P3_DATAO_REG_10__SCAN_IN), .S(n12740), .Z(
        P3_U3501) );
  MUX2_X1 U15064 ( .A(n12734), .B(P3_DATAO_REG_9__SCAN_IN), .S(n12740), .Z(
        P3_U3500) );
  MUX2_X1 U15065 ( .A(n12735), .B(P3_DATAO_REG_7__SCAN_IN), .S(n12740), .Z(
        P3_U3498) );
  MUX2_X1 U15066 ( .A(n12736), .B(P3_DATAO_REG_6__SCAN_IN), .S(n12740), .Z(
        P3_U3497) );
  MUX2_X1 U15067 ( .A(n12737), .B(P3_DATAO_REG_5__SCAN_IN), .S(n12740), .Z(
        P3_U3496) );
  MUX2_X1 U15068 ( .A(n12738), .B(P3_DATAO_REG_4__SCAN_IN), .S(n12740), .Z(
        P3_U3495) );
  MUX2_X1 U15069 ( .A(n12739), .B(P3_DATAO_REG_3__SCAN_IN), .S(n12740), .Z(
        P3_U3494) );
  MUX2_X1 U15070 ( .A(n10781), .B(P3_DATAO_REG_2__SCAN_IN), .S(n12740), .Z(
        P3_U3493) );
  MUX2_X1 U15071 ( .A(n10719), .B(P3_DATAO_REG_1__SCAN_IN), .S(n12740), .Z(
        P3_U3492) );
  MUX2_X1 U15072 ( .A(n12741), .B(P3_DATAO_REG_0__SCAN_IN), .S(n12740), .Z(
        P3_U3491) );
  NAND2_X1 U15073 ( .A1(n12743), .A2(n12742), .ZN(n12772) );
  XNOR2_X1 U15074 ( .A(n12772), .B(n6775), .ZN(n12771) );
  XNOR2_X1 U15075 ( .A(n12771), .B(n12757), .ZN(n12753) );
  INV_X1 U15076 ( .A(P3_REG2_REG_14__SCAN_IN), .ZN(n12745) );
  NAND2_X1 U15077 ( .A1(P3_REG2_REG_15__SCAN_IN), .A2(n12747), .ZN(n12765) );
  OAI21_X1 U15078 ( .B1(n12747), .B2(P3_REG2_REG_15__SCAN_IN), .A(n12765), 
        .ZN(n12751) );
  INV_X1 U15079 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n12749) );
  OAI21_X1 U15080 ( .B1(n15413), .B2(n12749), .A(n12748), .ZN(n12750) );
  AOI21_X1 U15081 ( .B1(n15429), .B2(n12751), .A(n12750), .ZN(n12752) );
  OAI21_X1 U15082 ( .B1(n12753), .B2(n12841), .A(n12752), .ZN(n12762) );
  MUX2_X1 U15083 ( .A(P3_REG2_REG_14__SCAN_IN), .B(P3_REG1_REG_14__SCAN_IN), 
        .S(n13165), .Z(n12755) );
  MUX2_X1 U15084 ( .A(n12758), .B(n12757), .S(n13165), .Z(n12759) );
  AOI211_X1 U15085 ( .C1(n12760), .C2(n12759), .A(n15406), .B(n12782), .ZN(
        n12761) );
  AOI211_X1 U15086 ( .C1(n15417), .C2(n6775), .A(n12762), .B(n12761), .ZN(
        n12763) );
  INV_X1 U15087 ( .A(n12763), .ZN(P3_U3197) );
  INV_X1 U15088 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n12792) );
  AOI22_X1 U15089 ( .A1(P3_REG2_REG_16__SCAN_IN), .A2(n12802), .B1(n12794), 
        .B2(n12792), .ZN(n12768) );
  NAND2_X1 U15090 ( .A1(n12764), .A2(n12784), .ZN(n12766) );
  NAND2_X1 U15091 ( .A1(n12766), .A2(n12765), .ZN(n12767) );
  NAND2_X1 U15092 ( .A1(n12768), .A2(n12767), .ZN(n12791) );
  OAI21_X1 U15093 ( .B1(n12768), .B2(n12767), .A(n12791), .ZN(n12789) );
  NAND2_X1 U15094 ( .A1(n15417), .A2(n12794), .ZN(n12780) );
  INV_X1 U15095 ( .A(n12769), .ZN(n12770) );
  AOI21_X1 U15096 ( .B1(n15415), .B2(P3_ADDR_REG_16__SCAN_IN), .A(n12770), 
        .ZN(n12779) );
  NAND2_X1 U15097 ( .A1(n12771), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n12774) );
  NAND2_X1 U15098 ( .A1(n12772), .A2(n12784), .ZN(n12773) );
  NAND2_X1 U15099 ( .A1(n12774), .A2(n12773), .ZN(n12776) );
  XNOR2_X1 U15100 ( .A(n12794), .B(P3_REG1_REG_16__SCAN_IN), .ZN(n12775) );
  NAND2_X1 U15101 ( .A1(n12775), .A2(n12776), .ZN(n12795) );
  OAI21_X1 U15102 ( .B1(n12776), .B2(n12775), .A(n12795), .ZN(n12777) );
  NAND2_X1 U15103 ( .A1(n15426), .A2(n12777), .ZN(n12778) );
  NAND3_X1 U15104 ( .A1(n12780), .A2(n12779), .A3(n12778), .ZN(n12788) );
  INV_X1 U15105 ( .A(n12781), .ZN(n12783) );
  MUX2_X1 U15106 ( .A(P3_REG2_REG_16__SCAN_IN), .B(P3_REG1_REG_16__SCAN_IN), 
        .S(n13165), .Z(n12803) );
  XNOR2_X1 U15107 ( .A(n12803), .B(n12802), .ZN(n12785) );
  NOR2_X1 U15108 ( .A1(n12786), .A2(n12785), .ZN(n12801) );
  AOI211_X1 U15109 ( .C1(n12786), .C2(n12785), .A(n15406), .B(n12801), .ZN(
        n12787) );
  AOI211_X1 U15110 ( .C1(n15429), .C2(n12789), .A(n12788), .B(n12787), .ZN(
        n12790) );
  INV_X1 U15111 ( .A(n12790), .ZN(P3_U3198) );
  XOR2_X1 U15112 ( .A(P3_REG2_REG_17__SCAN_IN), .B(n12810), .Z(n12809) );
  OR2_X1 U15113 ( .A1(n12794), .A2(n12793), .ZN(n12796) );
  XNOR2_X1 U15114 ( .A(n12816), .B(P3_REG1_REG_17__SCAN_IN), .ZN(n12800) );
  INV_X1 U15115 ( .A(n12797), .ZN(n12799) );
  NAND2_X1 U15116 ( .A1(n15415), .A2(P3_ADDR_REG_17__SCAN_IN), .ZN(n12798) );
  OAI211_X1 U15117 ( .C1(n12841), .C2(n12800), .A(n12799), .B(n12798), .ZN(
        n12807) );
  MUX2_X1 U15118 ( .A(P3_REG2_REG_17__SCAN_IN), .B(P3_REG1_REG_17__SCAN_IN), 
        .S(n13165), .Z(n12812) );
  XNOR2_X1 U15119 ( .A(n12812), .B(n12817), .ZN(n12804) );
  NOR2_X1 U15120 ( .A1(n12805), .A2(n12804), .ZN(n12811) );
  AOI211_X1 U15121 ( .C1(n12805), .C2(n12804), .A(n15406), .B(n12811), .ZN(
        n12806) );
  AOI211_X1 U15122 ( .C1(n15417), .C2(n6866), .A(n12807), .B(n12806), .ZN(
        n12808) );
  OAI21_X1 U15123 ( .B1(n12809), .B2(n15401), .A(n12808), .ZN(P3_U3199) );
  XNOR2_X1 U15124 ( .A(n14799), .B(P3_REG2_REG_18__SCAN_IN), .ZN(n12843) );
  XOR2_X1 U15125 ( .A(n12843), .B(n12844), .Z(n12828) );
  XNOR2_X1 U15126 ( .A(n12829), .B(n14799), .ZN(n12814) );
  MUX2_X1 U15127 ( .A(n13006), .B(n12820), .S(n13165), .Z(n12813) );
  OAI21_X1 U15128 ( .B1(n12814), .B2(n12813), .A(n12830), .ZN(n12815) );
  NAND2_X1 U15129 ( .A1(n12815), .A2(n15430), .ZN(n12827) );
  INV_X1 U15130 ( .A(n14799), .ZN(n12842) );
  NAND2_X1 U15131 ( .A1(n12818), .A2(n12817), .ZN(n12819) );
  XNOR2_X1 U15132 ( .A(n14799), .B(n12820), .ZN(n12835) );
  INV_X1 U15133 ( .A(n12835), .ZN(n12821) );
  XNOR2_X1 U15134 ( .A(n12836), .B(n12821), .ZN(n12824) );
  NAND2_X1 U15135 ( .A1(n15415), .A2(P3_ADDR_REG_18__SCAN_IN), .ZN(n12822) );
  OAI211_X1 U15136 ( .C1(n12841), .C2(n12824), .A(n12823), .B(n12822), .ZN(
        n12825) );
  AOI21_X1 U15137 ( .B1(n12842), .B2(n15417), .A(n12825), .ZN(n12826) );
  OAI211_X1 U15138 ( .C1(n12828), .C2(n15401), .A(n12827), .B(n12826), .ZN(
        P3_U3200) );
  INV_X1 U15139 ( .A(n12829), .ZN(n12831) );
  OAI21_X1 U15140 ( .B1(n12831), .B2(n14799), .A(n12830), .ZN(n12834) );
  XNOR2_X1 U15141 ( .A(n12832), .B(P3_REG2_REG_19__SCAN_IN), .ZN(n12845) );
  XNOR2_X1 U15142 ( .A(n12832), .B(P3_REG1_REG_19__SCAN_IN), .ZN(n12837) );
  MUX2_X1 U15143 ( .A(n12845), .B(n12837), .S(n13165), .Z(n12833) );
  XNOR2_X1 U15144 ( .A(n12834), .B(n12833), .ZN(n12848) );
  AOI22_X1 U15145 ( .A1(n12836), .A2(n12835), .B1(P3_REG1_REG_18__SCAN_IN), 
        .B2(n14799), .ZN(n12838) );
  NAND2_X1 U15146 ( .A1(n15415), .A2(P3_ADDR_REG_19__SCAN_IN), .ZN(n12840) );
  INV_X1 U15147 ( .A(n12849), .ZN(n12850) );
  NAND2_X1 U15148 ( .A1(n12851), .A2(n12850), .ZN(n14817) );
  AOI21_X1 U15149 ( .B1(n12852), .B2(n14817), .A(n13024), .ZN(n12855) );
  AOI21_X1 U15150 ( .B1(n13024), .B2(P3_REG2_REG_31__SCAN_IN), .A(n12855), 
        .ZN(n12853) );
  OAI21_X1 U15151 ( .B1(n12854), .B2(n15442), .A(n12853), .ZN(P3_U3202) );
  AOI21_X1 U15152 ( .B1(n13024), .B2(P3_REG2_REG_30__SCAN_IN), .A(n12855), 
        .ZN(n12856) );
  OAI21_X1 U15153 ( .B1(n12857), .B2(n15442), .A(n12856), .ZN(P3_U3203) );
  AOI21_X1 U15154 ( .B1(n12858), .B2(n7470), .A(n15457), .ZN(n12862) );
  OAI22_X1 U15155 ( .A1(n12859), .A2(n15450), .B1(n12891), .B2(n15452), .ZN(
        n12860) );
  AOI21_X1 U15156 ( .B1(n12862), .B2(n12861), .A(n12860), .ZN(n13041) );
  INV_X1 U15157 ( .A(n13042), .ZN(n12867) );
  AOI22_X1 U15158 ( .A1(n12864), .A2(n15463), .B1(n13024), .B2(
        P3_REG2_REG_28__SCAN_IN), .ZN(n12865) );
  OAI21_X1 U15159 ( .B1(n13107), .B2(n15442), .A(n12865), .ZN(n12866) );
  AOI21_X1 U15160 ( .B1(n12867), .B2(n13039), .A(n12866), .ZN(n12868) );
  OAI21_X1 U15161 ( .B1(n13041), .B2(n13024), .A(n12868), .ZN(P3_U3205) );
  INV_X1 U15162 ( .A(n12869), .ZN(n12870) );
  AOI21_X1 U15163 ( .B1(n12872), .B2(n12871), .A(n12870), .ZN(n12880) );
  AOI21_X1 U15164 ( .B1(n12875), .B2(n12874), .A(n12873), .ZN(n13044) );
  INV_X1 U15165 ( .A(n13044), .ZN(n12884) );
  OAI22_X1 U15166 ( .A1(n12877), .A2(n15450), .B1(n12876), .B2(n15452), .ZN(
        n12878) );
  AOI21_X1 U15167 ( .B1(n12884), .B2(n15454), .A(n12878), .ZN(n12879) );
  OAI21_X1 U15168 ( .B1(n12880), .B2(n15457), .A(n12879), .ZN(n13046) );
  INV_X1 U15169 ( .A(n13046), .ZN(n12886) );
  AOI22_X1 U15170 ( .A1(n12881), .A2(n15463), .B1(n13024), .B2(
        P3_REG2_REG_27__SCAN_IN), .ZN(n12882) );
  OAI21_X1 U15171 ( .B1(n13111), .B2(n15442), .A(n12882), .ZN(n12883) );
  AOI21_X1 U15172 ( .B1(n12884), .B2(n12927), .A(n12883), .ZN(n12885) );
  OAI21_X1 U15173 ( .B1(n12886), .B2(n13024), .A(n12885), .ZN(P3_U3206) );
  XNOR2_X1 U15174 ( .A(n12887), .B(n12888), .ZN(n12894) );
  INV_X1 U15175 ( .A(n12888), .ZN(n12889) );
  XNOR2_X1 U15176 ( .A(n12890), .B(n12889), .ZN(n13050) );
  OAI22_X1 U15177 ( .A1(n12891), .A2(n15450), .B1(n12920), .B2(n15452), .ZN(
        n12892) );
  AOI21_X1 U15178 ( .B1(n13050), .B2(n15454), .A(n12892), .ZN(n12893) );
  OAI21_X1 U15179 ( .B1(n12894), .B2(n15457), .A(n12893), .ZN(n13049) );
  INV_X1 U15180 ( .A(n13049), .ZN(n12899) );
  AOI22_X1 U15181 ( .A1(n12895), .A2(n15463), .B1(n13024), .B2(
        P3_REG2_REG_26__SCAN_IN), .ZN(n12896) );
  OAI21_X1 U15182 ( .B1(n9638), .B2(n15442), .A(n12896), .ZN(n12897) );
  AOI21_X1 U15183 ( .B1(n13050), .B2(n12927), .A(n12897), .ZN(n12898) );
  OAI21_X1 U15184 ( .B1(n12899), .B2(n13024), .A(n12898), .ZN(P3_U3207) );
  XOR2_X1 U15185 ( .A(n12902), .B(n12900), .Z(n12907) );
  OAI211_X1 U15186 ( .C1(n7508), .C2(n7507), .A(n13032), .B(n12903), .ZN(
        n12906) );
  AOI22_X1 U15187 ( .A1(n12904), .A2(n13029), .B1(n13027), .B2(n12941), .ZN(
        n12905) );
  OAI211_X1 U15188 ( .C1(n12944), .C2(n12907), .A(n12906), .B(n12905), .ZN(
        n13053) );
  INV_X1 U15189 ( .A(n13053), .ZN(n12913) );
  INV_X1 U15190 ( .A(n12907), .ZN(n13054) );
  INV_X1 U15191 ( .A(n12908), .ZN(n13118) );
  AOI22_X1 U15192 ( .A1(n13024), .A2(P3_REG2_REG_25__SCAN_IN), .B1(n12909), 
        .B2(n15463), .ZN(n12910) );
  OAI21_X1 U15193 ( .B1(n13118), .B2(n15442), .A(n12910), .ZN(n12911) );
  AOI21_X1 U15194 ( .B1(n13054), .B2(n12927), .A(n12911), .ZN(n12912) );
  OAI21_X1 U15195 ( .B1(n12913), .B2(n13024), .A(n12912), .ZN(P3_U3208) );
  XNOR2_X1 U15196 ( .A(n12915), .B(n12914), .ZN(n12923) );
  INV_X1 U15197 ( .A(n12916), .ZN(n12919) );
  OAI21_X1 U15198 ( .B1(n12919), .B2(n12918), .A(n12917), .ZN(n13058) );
  OAI22_X1 U15199 ( .A1(n12920), .A2(n15450), .B1(n12955), .B2(n15452), .ZN(
        n12921) );
  AOI21_X1 U15200 ( .B1(n13058), .B2(n15454), .A(n12921), .ZN(n12922) );
  OAI21_X1 U15201 ( .B1(n12923), .B2(n15457), .A(n12922), .ZN(n13057) );
  INV_X1 U15202 ( .A(n13057), .ZN(n12929) );
  AOI22_X1 U15203 ( .A1(n13024), .A2(P3_REG2_REG_24__SCAN_IN), .B1(n15463), 
        .B2(n12924), .ZN(n12925) );
  OAI21_X1 U15204 ( .B1(n13122), .B2(n15442), .A(n12925), .ZN(n12926) );
  AOI21_X1 U15205 ( .B1(n13058), .B2(n12927), .A(n12926), .ZN(n12928) );
  OAI21_X1 U15206 ( .B1(n12929), .B2(n13024), .A(n12928), .ZN(P3_U3209) );
  OR2_X1 U15207 ( .A1(n12930), .A2(n12937), .ZN(n12931) );
  NAND2_X1 U15208 ( .A1(n12932), .A2(n12931), .ZN(n13061) );
  OR2_X1 U15209 ( .A1(n12933), .A2(n12934), .ZN(n12936) );
  NAND2_X1 U15210 ( .A1(n12936), .A2(n12935), .ZN(n12938) );
  XNOR2_X1 U15211 ( .A(n12938), .B(n12937), .ZN(n12939) );
  NAND2_X1 U15212 ( .A1(n12939), .A2(n13032), .ZN(n12943) );
  AOI22_X1 U15213 ( .A1(n12941), .A2(n13029), .B1(n13027), .B2(n12940), .ZN(
        n12942) );
  OAI211_X1 U15214 ( .C1(n12944), .C2(n13061), .A(n12943), .B(n12942), .ZN(
        n13062) );
  NAND2_X1 U15215 ( .A1(n13062), .A2(n15464), .ZN(n12951) );
  INV_X1 U15216 ( .A(P3_REG2_REG_23__SCAN_IN), .ZN(n12947) );
  INV_X1 U15217 ( .A(n12945), .ZN(n12946) );
  OAI22_X1 U15218 ( .A1(n15464), .A2(n12947), .B1(n12946), .B2(n15440), .ZN(
        n12948) );
  AOI21_X1 U15219 ( .B1(n12949), .B2(n13008), .A(n12948), .ZN(n12950) );
  OAI211_X1 U15220 ( .C1(n13061), .C2(n12952), .A(n12951), .B(n12950), .ZN(
        P3_U3210) );
  XNOR2_X1 U15221 ( .A(n12933), .B(n12956), .ZN(n12953) );
  OAI222_X1 U15222 ( .A1(n15450), .A2(n12955), .B1(n15452), .B2(n12954), .C1(
        n15457), .C2(n12953), .ZN(n13066) );
  INV_X1 U15223 ( .A(n13066), .ZN(n12963) );
  XOR2_X1 U15224 ( .A(n12957), .B(n12956), .Z(n13067) );
  INV_X1 U15225 ( .A(n12958), .ZN(n13130) );
  AOI22_X1 U15226 ( .A1(n13024), .A2(P3_REG2_REG_22__SCAN_IN), .B1(n15463), 
        .B2(n12959), .ZN(n12960) );
  OAI21_X1 U15227 ( .B1(n13130), .B2(n15442), .A(n12960), .ZN(n12961) );
  AOI21_X1 U15228 ( .B1(n13067), .B2(n13039), .A(n12961), .ZN(n12962) );
  OAI21_X1 U15229 ( .B1(n12963), .B2(n13024), .A(n12962), .ZN(P3_U3211) );
  XOR2_X1 U15230 ( .A(n12968), .B(n12964), .Z(n12965) );
  OAI222_X1 U15231 ( .A1(n15450), .A2(n12967), .B1(n15452), .B2(n12966), .C1(
        n15457), .C2(n12965), .ZN(n13070) );
  INV_X1 U15232 ( .A(n13070), .ZN(n12974) );
  XOR2_X1 U15233 ( .A(n12969), .B(n12968), .Z(n13071) );
  AOI22_X1 U15234 ( .A1(n13024), .A2(P3_REG2_REG_21__SCAN_IN), .B1(n15463), 
        .B2(n12970), .ZN(n12971) );
  OAI21_X1 U15235 ( .B1(n13134), .B2(n15442), .A(n12971), .ZN(n12972) );
  AOI21_X1 U15236 ( .B1(n13071), .B2(n13039), .A(n12972), .ZN(n12973) );
  OAI21_X1 U15237 ( .B1(n12974), .B2(n13024), .A(n12973), .ZN(P3_U3212) );
  XNOR2_X1 U15238 ( .A(n12975), .B(n12976), .ZN(n12978) );
  AOI222_X1 U15239 ( .A1(n13032), .A2(n12978), .B1(n13003), .B2(n13027), .C1(
        n12977), .C2(n13029), .ZN(n13077) );
  INV_X1 U15240 ( .A(P3_REG2_REG_20__SCAN_IN), .ZN(n12980) );
  OAI22_X1 U15241 ( .A1(n15464), .A2(n12980), .B1(n12979), .B2(n15440), .ZN(
        n12981) );
  AOI21_X1 U15242 ( .B1(n12982), .B2(n13008), .A(n12981), .ZN(n12986) );
  NAND2_X1 U15243 ( .A1(n12984), .A2(n12983), .ZN(n13074) );
  NAND3_X1 U15244 ( .A1(n13075), .A2(n13074), .A3(n13039), .ZN(n12985) );
  OAI211_X1 U15245 ( .C1(n13077), .C2(n13024), .A(n12986), .B(n12985), .ZN(
        P3_U3213) );
  INV_X1 U15246 ( .A(n12995), .ZN(n12988) );
  OAI211_X1 U15247 ( .C1(n6745), .C2(n12988), .A(n13032), .B(n12987), .ZN(
        n12992) );
  AOI22_X1 U15248 ( .A1(n13027), .A2(n12990), .B1(n12989), .B2(n13029), .ZN(
        n12991) );
  NAND2_X1 U15249 ( .A1(n12992), .A2(n12991), .ZN(n13079) );
  INV_X1 U15250 ( .A(n13079), .ZN(n13001) );
  NAND2_X1 U15251 ( .A1(n13084), .A2(n12993), .ZN(n12994) );
  XOR2_X1 U15252 ( .A(n12995), .B(n12994), .Z(n13080) );
  NOR2_X1 U15253 ( .A1(n13139), .A2(n15442), .ZN(n12999) );
  INV_X1 U15254 ( .A(P3_REG2_REG_19__SCAN_IN), .ZN(n12997) );
  OAI22_X1 U15255 ( .A1(n15464), .A2(n12997), .B1(n12996), .B2(n15440), .ZN(
        n12998) );
  AOI211_X1 U15256 ( .C1(n13080), .C2(n13039), .A(n12999), .B(n12998), .ZN(
        n13000) );
  OAI21_X1 U15257 ( .B1(n13001), .B2(n13024), .A(n13000), .ZN(P3_U3214) );
  OAI21_X1 U15258 ( .B1(n6651), .B2(n9517), .A(n13002), .ZN(n13004) );
  AOI222_X1 U15259 ( .A1(n13032), .A2(n13004), .B1(n13003), .B2(n13029), .C1(
        n13030), .C2(n13027), .ZN(n13086) );
  OAI22_X1 U15260 ( .A1(n15464), .A2(n13006), .B1(n13005), .B2(n15440), .ZN(
        n13007) );
  AOI21_X1 U15261 ( .B1(n13009), .B2(n13008), .A(n13007), .ZN(n13012) );
  NAND2_X1 U15262 ( .A1(n13010), .A2(n9517), .ZN(n13083) );
  NAND3_X1 U15263 ( .A1(n13084), .A2(n13039), .A3(n13083), .ZN(n13011) );
  OAI211_X1 U15264 ( .C1(n13086), .C2(n13024), .A(n13012), .B(n13011), .ZN(
        P3_U3215) );
  XNOR2_X1 U15265 ( .A(n13014), .B(n13013), .ZN(n13015) );
  OAI222_X1 U15266 ( .A1(n15450), .A2(n13017), .B1(n15452), .B2(n13016), .C1(
        n13015), .C2(n15457), .ZN(n13088) );
  INV_X1 U15267 ( .A(n13088), .ZN(n13025) );
  OAI22_X1 U15268 ( .A1(n15442), .A2(n13145), .B1(n13018), .B2(n15440), .ZN(
        n13019) );
  AOI21_X1 U15269 ( .B1(P3_REG2_REG_17__SCAN_IN), .B2(n13024), .A(n13019), 
        .ZN(n13023) );
  XNOR2_X1 U15270 ( .A(n13021), .B(n13020), .ZN(n13089) );
  NAND2_X1 U15271 ( .A1(n13089), .A2(n13039), .ZN(n13022) );
  OAI211_X1 U15272 ( .C1(n13025), .C2(n13024), .A(n13023), .B(n13022), .ZN(
        P3_U3216) );
  XOR2_X1 U15273 ( .A(n13033), .B(n13026), .Z(n13031) );
  AOI222_X1 U15274 ( .A1(n13032), .A2(n13031), .B1(n13030), .B2(n13029), .C1(
        n13028), .C2(n13027), .ZN(n13096) );
  XNOR2_X1 U15275 ( .A(n13034), .B(n13033), .ZN(n13094) );
  NOR2_X1 U15276 ( .A1(n13035), .A2(n15442), .ZN(n13038) );
  OAI22_X1 U15277 ( .A1(n15464), .A2(n12792), .B1(n13036), .B2(n15440), .ZN(
        n13037) );
  AOI211_X1 U15278 ( .C1(n13094), .C2(n13039), .A(n13038), .B(n13037), .ZN(
        n13040) );
  OAI21_X1 U15279 ( .B1(n13096), .B2(n13024), .A(n13040), .ZN(P3_U3217) );
  INV_X1 U15280 ( .A(n15477), .ZN(n14823) );
  OAI21_X1 U15281 ( .B1(n14823), .B2(n13042), .A(n13041), .ZN(n13105) );
  OAI21_X1 U15282 ( .B1(n13107), .B2(n13092), .A(n13043), .ZN(P3_U3487) );
  INV_X1 U15283 ( .A(n15475), .ZN(n15487) );
  NOR2_X1 U15284 ( .A1(n13044), .A2(n15487), .ZN(n13045) );
  NOR2_X1 U15285 ( .A1(n13046), .A2(n13045), .ZN(n13108) );
  MUX2_X1 U15286 ( .A(n13047), .B(n13108), .S(n15498), .Z(n13048) );
  OAI21_X1 U15287 ( .B1(n13111), .B2(n13092), .A(n13048), .ZN(P3_U3486) );
  AOI21_X1 U15288 ( .B1(n15475), .B2(n13050), .A(n13049), .ZN(n13112) );
  MUX2_X1 U15289 ( .A(n13051), .B(n13112), .S(n15498), .Z(n13052) );
  OAI21_X1 U15290 ( .B1(n9638), .B2(n13092), .A(n13052), .ZN(P3_U3485) );
  INV_X1 U15291 ( .A(P3_REG1_REG_25__SCAN_IN), .ZN(n13055) );
  AOI21_X1 U15292 ( .B1(n15475), .B2(n13054), .A(n13053), .ZN(n13115) );
  MUX2_X1 U15293 ( .A(n13055), .B(n13115), .S(n15498), .Z(n13056) );
  OAI21_X1 U15294 ( .B1(n13118), .B2(n13092), .A(n13056), .ZN(P3_U3484) );
  INV_X1 U15295 ( .A(P3_REG1_REG_24__SCAN_IN), .ZN(n13059) );
  AOI21_X1 U15296 ( .B1(n15475), .B2(n13058), .A(n13057), .ZN(n13119) );
  MUX2_X1 U15297 ( .A(n13059), .B(n13119), .S(n15498), .Z(n13060) );
  OAI21_X1 U15298 ( .B1(n13122), .B2(n13092), .A(n13060), .ZN(P3_U3483) );
  INV_X1 U15299 ( .A(n13061), .ZN(n13063) );
  AOI21_X1 U15300 ( .B1(n15475), .B2(n13063), .A(n13062), .ZN(n13123) );
  MUX2_X1 U15301 ( .A(n13064), .B(n13123), .S(n15498), .Z(n13065) );
  OAI21_X1 U15302 ( .B1(n13126), .B2(n13092), .A(n13065), .ZN(P3_U3482) );
  AOI21_X1 U15303 ( .B1(n15477), .B2(n13067), .A(n13066), .ZN(n13127) );
  MUX2_X1 U15304 ( .A(n13068), .B(n13127), .S(n15498), .Z(n13069) );
  OAI21_X1 U15305 ( .B1(n13130), .B2(n13092), .A(n13069), .ZN(P3_U3481) );
  AOI21_X1 U15306 ( .B1(n13071), .B2(n15477), .A(n13070), .ZN(n13131) );
  MUX2_X1 U15307 ( .A(n13072), .B(n13131), .S(n15498), .Z(n13073) );
  OAI21_X1 U15308 ( .B1(n13134), .B2(n13092), .A(n13073), .ZN(P3_U3480) );
  NAND3_X1 U15309 ( .A1(n13075), .A2(n13074), .A3(n15477), .ZN(n13076) );
  OAI211_X1 U15310 ( .C1(n13078), .C2(n15486), .A(n13077), .B(n13076), .ZN(
        n13135) );
  MUX2_X1 U15311 ( .A(P3_REG1_REG_20__SCAN_IN), .B(n13135), .S(n15498), .Z(
        P3_U3479) );
  AOI21_X1 U15312 ( .B1(n15477), .B2(n13080), .A(n13079), .ZN(n13136) );
  MUX2_X1 U15313 ( .A(n13081), .B(n13136), .S(n15498), .Z(n13082) );
  OAI21_X1 U15314 ( .B1(n13092), .B2(n13139), .A(n13082), .ZN(P3_U3478) );
  NAND3_X1 U15315 ( .A1(n13084), .A2(n15477), .A3(n13083), .ZN(n13085) );
  OAI211_X1 U15316 ( .C1(n13087), .C2(n15486), .A(n13086), .B(n13085), .ZN(
        n13140) );
  MUX2_X1 U15317 ( .A(P3_REG1_REG_18__SCAN_IN), .B(n13140), .S(n15498), .Z(
        P3_U3477) );
  AOI21_X1 U15318 ( .B1(n13089), .B2(n15477), .A(n13088), .ZN(n13141) );
  MUX2_X1 U15319 ( .A(n13090), .B(n13141), .S(n15498), .Z(n13091) );
  OAI21_X1 U15320 ( .B1(n13145), .B2(n13092), .A(n13091), .ZN(P3_U3476) );
  AOI22_X1 U15321 ( .A1(n13094), .A2(n15477), .B1(n15479), .B2(n13093), .ZN(
        n13095) );
  NAND2_X1 U15322 ( .A1(n13096), .A2(n13095), .ZN(n13146) );
  MUX2_X1 U15323 ( .A(P3_REG1_REG_16__SCAN_IN), .B(n13146), .S(n15498), .Z(
        P3_U3475) );
  AOI22_X1 U15324 ( .A1(n13098), .A2(n15477), .B1(n15479), .B2(n13097), .ZN(
        n13099) );
  NAND2_X1 U15325 ( .A1(n13100), .A2(n13099), .ZN(n13147) );
  MUX2_X1 U15326 ( .A(P3_REG1_REG_15__SCAN_IN), .B(n13147), .S(n15498), .Z(
        P3_U3474) );
  AOI22_X1 U15327 ( .A1(n13102), .A2(n15477), .B1(n15479), .B2(n13101), .ZN(
        n13103) );
  NAND2_X1 U15328 ( .A1(n13104), .A2(n13103), .ZN(n13148) );
  MUX2_X1 U15329 ( .A(P3_REG1_REG_14__SCAN_IN), .B(n13148), .S(n15498), .Z(
        P3_U3473) );
  OAI21_X1 U15330 ( .B1(n13107), .B2(n13144), .A(n13106), .ZN(P3_U3455) );
  INV_X1 U15331 ( .A(P3_REG0_REG_27__SCAN_IN), .ZN(n13109) );
  MUX2_X1 U15332 ( .A(n13109), .B(n13108), .S(n15493), .Z(n13110) );
  OAI21_X1 U15333 ( .B1(n13111), .B2(n13144), .A(n13110), .ZN(P3_U3454) );
  INV_X1 U15334 ( .A(P3_REG0_REG_26__SCAN_IN), .ZN(n13113) );
  MUX2_X1 U15335 ( .A(n13113), .B(n13112), .S(n15493), .Z(n13114) );
  OAI21_X1 U15336 ( .B1(n9638), .B2(n13144), .A(n13114), .ZN(P3_U3453) );
  INV_X1 U15337 ( .A(P3_REG0_REG_25__SCAN_IN), .ZN(n13116) );
  MUX2_X1 U15338 ( .A(n13116), .B(n13115), .S(n15493), .Z(n13117) );
  OAI21_X1 U15339 ( .B1(n13118), .B2(n13144), .A(n13117), .ZN(P3_U3452) );
  MUX2_X1 U15340 ( .A(n13120), .B(n13119), .S(n15493), .Z(n13121) );
  OAI21_X1 U15341 ( .B1(n13122), .B2(n13144), .A(n13121), .ZN(P3_U3451) );
  INV_X1 U15342 ( .A(P3_REG0_REG_23__SCAN_IN), .ZN(n13124) );
  MUX2_X1 U15343 ( .A(n13124), .B(n13123), .S(n15493), .Z(n13125) );
  OAI21_X1 U15344 ( .B1(n13126), .B2(n13144), .A(n13125), .ZN(P3_U3450) );
  INV_X1 U15345 ( .A(P3_REG0_REG_22__SCAN_IN), .ZN(n13128) );
  MUX2_X1 U15346 ( .A(n13128), .B(n13127), .S(n15493), .Z(n13129) );
  OAI21_X1 U15347 ( .B1(n13130), .B2(n13144), .A(n13129), .ZN(P3_U3449) );
  INV_X1 U15348 ( .A(P3_REG0_REG_21__SCAN_IN), .ZN(n13132) );
  MUX2_X1 U15349 ( .A(n13132), .B(n13131), .S(n15493), .Z(n13133) );
  OAI21_X1 U15350 ( .B1(n13134), .B2(n13144), .A(n13133), .ZN(P3_U3448) );
  MUX2_X1 U15351 ( .A(P3_REG0_REG_20__SCAN_IN), .B(n13135), .S(n15493), .Z(
        P3_U3447) );
  INV_X1 U15352 ( .A(P3_REG0_REG_19__SCAN_IN), .ZN(n13137) );
  MUX2_X1 U15353 ( .A(n13137), .B(n13136), .S(n15493), .Z(n13138) );
  OAI21_X1 U15354 ( .B1(n13144), .B2(n13139), .A(n13138), .ZN(P3_U3446) );
  MUX2_X1 U15355 ( .A(P3_REG0_REG_18__SCAN_IN), .B(n13140), .S(n15493), .Z(
        P3_U3444) );
  INV_X1 U15356 ( .A(P3_REG0_REG_17__SCAN_IN), .ZN(n13142) );
  MUX2_X1 U15357 ( .A(n13142), .B(n13141), .S(n15493), .Z(n13143) );
  OAI21_X1 U15358 ( .B1(n13145), .B2(n13144), .A(n13143), .ZN(P3_U3441) );
  MUX2_X1 U15359 ( .A(P3_REG0_REG_16__SCAN_IN), .B(n13146), .S(n15493), .Z(
        P3_U3438) );
  MUX2_X1 U15360 ( .A(P3_REG0_REG_15__SCAN_IN), .B(n13147), .S(n15493), .Z(
        P3_U3435) );
  MUX2_X1 U15361 ( .A(P3_REG0_REG_14__SCAN_IN), .B(n13148), .S(n15493), .Z(
        P3_U3432) );
  MUX2_X1 U15362 ( .A(n13150), .B(P3_D_REG_1__SCAN_IN), .S(n13149), .Z(
        P3_U3377) );
  MUX2_X1 U15363 ( .A(P3_D_REG_0__SCAN_IN), .B(n13152), .S(n13151), .Z(
        P3_U3376) );
  INV_X1 U15364 ( .A(n13153), .ZN(n13154) );
  OAI222_X1 U15365 ( .A1(n9199), .A2(P3_U3151), .B1(n13167), .B2(n13155), .C1(
        n13172), .C2(n13154), .ZN(P3_U3265) );
  INV_X1 U15366 ( .A(n13156), .ZN(n13157) );
  OAI222_X1 U15367 ( .A1(n13167), .A2(n13159), .B1(P3_U3151), .B2(n13158), 
        .C1(n13172), .C2(n13157), .ZN(P3_U3266) );
  INV_X1 U15368 ( .A(n13160), .ZN(n13161) );
  OAI222_X1 U15369 ( .A1(n13167), .A2(n13163), .B1(P3_U3151), .B2(n13162), 
        .C1(n13172), .C2(n13161), .ZN(P3_U3267) );
  INV_X1 U15370 ( .A(n13164), .ZN(n13168) );
  OAI222_X1 U15371 ( .A1(n13172), .A2(n13168), .B1(n13167), .B2(n13166), .C1(
        P3_U3151), .C2(n13165), .ZN(P3_U3268) );
  INV_X1 U15372 ( .A(n13169), .ZN(n13171) );
  OAI222_X1 U15373 ( .A1(n6828), .A2(P3_U3151), .B1(n13172), .B2(n13171), .C1(
        n13170), .C2(n13167), .ZN(P3_U3269) );
  INV_X1 U15374 ( .A(n13688), .ZN(n13233) );
  XNOR2_X1 U15375 ( .A(n13557), .B(n13255), .ZN(n13199) );
  NAND2_X1 U15376 ( .A1(n13363), .A2(n13651), .ZN(n13200) );
  XNOR2_X1 U15377 ( .A(n13726), .B(n13255), .ZN(n13196) );
  INV_X1 U15378 ( .A(n13196), .ZN(n13198) );
  NOR2_X1 U15379 ( .A1(n13270), .A2(n13604), .ZN(n13195) );
  INV_X1 U15380 ( .A(n13195), .ZN(n13197) );
  XNOR2_X1 U15381 ( .A(n13731), .B(n13255), .ZN(n13192) );
  INV_X1 U15382 ( .A(n13192), .ZN(n13194) );
  NAND2_X1 U15383 ( .A1(n13365), .A2(n13651), .ZN(n13193) );
  XNOR2_X1 U15384 ( .A(n13630), .B(n13213), .ZN(n13187) );
  NAND2_X1 U15385 ( .A1(n13367), .A2(n13651), .ZN(n13186) );
  XNOR2_X1 U15386 ( .A(n14845), .B(n13213), .ZN(n13177) );
  NAND2_X1 U15387 ( .A1(n13651), .A2(n13370), .ZN(n13176) );
  XNOR2_X1 U15388 ( .A(n13177), .B(n13176), .ZN(n14839) );
  NAND2_X1 U15389 ( .A1(n13177), .A2(n13176), .ZN(n13178) );
  NAND2_X1 U15390 ( .A1(n14842), .A2(n13178), .ZN(n13180) );
  INV_X1 U15391 ( .A(n13180), .ZN(n13182) );
  XOR2_X1 U15392 ( .A(n13255), .B(n13642), .Z(n13179) );
  INV_X1 U15393 ( .A(n13179), .ZN(n13181) );
  NAND2_X1 U15394 ( .A1(n13369), .A2(n13651), .ZN(n13350) );
  XNOR2_X1 U15395 ( .A(n14853), .B(n13255), .ZN(n13183) );
  NAND2_X1 U15396 ( .A1(n13368), .A2(n13651), .ZN(n13184) );
  XNOR2_X1 U15397 ( .A(n13183), .B(n13184), .ZN(n14849) );
  INV_X1 U15398 ( .A(n13183), .ZN(n13185) );
  NAND2_X1 U15399 ( .A1(n13185), .A2(n13184), .ZN(n13287) );
  XNOR2_X1 U15400 ( .A(n13187), .B(n13186), .ZN(n13288) );
  XNOR2_X1 U15401 ( .A(n13609), .B(n13213), .ZN(n13189) );
  NAND2_X1 U15402 ( .A1(n13366), .A2(n13651), .ZN(n13188) );
  NOR2_X1 U15403 ( .A1(n13189), .A2(n13188), .ZN(n13190) );
  AOI21_X1 U15404 ( .B1(n13189), .B2(n13188), .A(n13190), .ZN(n13325) );
  INV_X1 U15405 ( .A(n13190), .ZN(n13191) );
  XOR2_X1 U15406 ( .A(n13193), .B(n13192), .Z(n13247) );
  XNOR2_X1 U15407 ( .A(n13196), .B(n13195), .ZN(n13311) );
  XNOR2_X1 U15408 ( .A(n13199), .B(n13200), .ZN(n13268) );
  NOR2_X1 U15409 ( .A1(n13271), .A2(n13604), .ZN(n13318) );
  INV_X1 U15410 ( .A(n13318), .ZN(n13201) );
  INV_X1 U15411 ( .A(n13203), .ZN(n13204) );
  NAND2_X1 U15412 ( .A1(n13204), .A2(n6664), .ZN(n13235) );
  XNOR2_X1 U15413 ( .A(n13524), .B(n13255), .ZN(n13237) );
  AND2_X1 U15414 ( .A1(n13361), .A2(n13651), .ZN(n13236) );
  NAND2_X1 U15415 ( .A1(n13234), .A2(n13206), .ZN(n13208) );
  NAND2_X1 U15416 ( .A1(n13208), .A2(n13207), .ZN(n13297) );
  XNOR2_X1 U15417 ( .A(n13703), .B(n13213), .ZN(n13210) );
  NAND2_X1 U15418 ( .A1(n13651), .A2(n13360), .ZN(n13209) );
  NOR2_X1 U15419 ( .A1(n13210), .A2(n13209), .ZN(n13211) );
  AOI21_X1 U15420 ( .B1(n13210), .B2(n13209), .A(n13211), .ZN(n13300) );
  NAND2_X1 U15421 ( .A1(n13297), .A2(n13300), .ZN(n13298) );
  INV_X1 U15422 ( .A(n13211), .ZN(n13212) );
  NAND2_X1 U15423 ( .A1(n13298), .A2(n13212), .ZN(n13276) );
  XNOR2_X1 U15424 ( .A(n13698), .B(n13213), .ZN(n13215) );
  NAND2_X1 U15425 ( .A1(n13651), .A2(n13359), .ZN(n13214) );
  NOR2_X1 U15426 ( .A1(n13215), .A2(n13214), .ZN(n13216) );
  AOI21_X1 U15427 ( .B1(n13215), .B2(n13214), .A(n13216), .ZN(n13279) );
  NAND2_X1 U15428 ( .A1(n13276), .A2(n13279), .ZN(n13277) );
  INV_X1 U15429 ( .A(n13216), .ZN(n13217) );
  NAND2_X1 U15430 ( .A1(n13277), .A2(n13217), .ZN(n13332) );
  INV_X1 U15431 ( .A(n13332), .ZN(n13219) );
  NAND2_X1 U15432 ( .A1(n13651), .A2(n13358), .ZN(n13220) );
  XNOR2_X1 U15433 ( .A(n6882), .B(n13255), .ZN(n13222) );
  XOR2_X1 U15434 ( .A(n13220), .B(n13222), .Z(n13335) );
  INV_X1 U15435 ( .A(n13335), .ZN(n13218) );
  INV_X1 U15436 ( .A(n13220), .ZN(n13221) );
  XNOR2_X1 U15437 ( .A(n13688), .B(n13255), .ZN(n13225) );
  AND2_X1 U15438 ( .A1(n13651), .A2(n13357), .ZN(n13224) );
  NAND2_X1 U15439 ( .A1(n13225), .A2(n13224), .ZN(n13252) );
  OAI21_X1 U15440 ( .B1(n13225), .B2(n13224), .A(n13252), .ZN(n13226) );
  NAND2_X1 U15441 ( .A1(n13228), .A2(n13227), .ZN(n13232) );
  OAI22_X1 U15442 ( .A1(n13280), .A2(n13303), .B1(n13254), .B2(n13301), .ZN(
        n13464) );
  OAI22_X1 U15443 ( .A1(n15198), .A2(n13469), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13229), .ZN(n13230) );
  AOI21_X1 U15444 ( .B1(n15190), .B2(n13464), .A(n13230), .ZN(n13231) );
  OAI211_X1 U15445 ( .C1(n13233), .C2(n13331), .A(n13232), .B(n13231), .ZN(
        P2_U3186) );
  NAND2_X1 U15446 ( .A1(n13234), .A2(n13235), .ZN(n13239) );
  XNOR2_X1 U15447 ( .A(n13237), .B(n13236), .ZN(n13238) );
  XNOR2_X1 U15448 ( .A(n13239), .B(n13238), .ZN(n13244) );
  AND2_X1 U15449 ( .A1(n13336), .A2(n13360), .ZN(n13240) );
  AOI21_X1 U15450 ( .B1(n13362), .B2(n13337), .A(n13240), .ZN(n13709) );
  AOI22_X1 U15451 ( .A1(n13344), .A2(n13523), .B1(P2_REG3_REG_23__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13241) );
  OAI21_X1 U15452 ( .B1(n13709), .B2(n13347), .A(n13241), .ZN(n13242) );
  AOI21_X1 U15453 ( .B1(n13524), .B2(n15195), .A(n13242), .ZN(n13243) );
  OAI21_X1 U15454 ( .B1(n13244), .B2(n13349), .A(n13243), .ZN(P2_U3188) );
  AOI21_X1 U15455 ( .B1(n13247), .B2(n13246), .A(n13245), .ZN(n13251) );
  OAI22_X1 U15456 ( .A1(n13270), .A2(n13301), .B1(n13292), .B2(n13303), .ZN(
        n13579) );
  NAND2_X1 U15457 ( .A1(n15190), .A2(n13579), .ZN(n13248) );
  NAND2_X1 U15458 ( .A1(P2_U3088), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n13432)
         );
  OAI211_X1 U15459 ( .C1(n15198), .C2(n13584), .A(n13248), .B(n13432), .ZN(
        n13249) );
  AOI21_X1 U15460 ( .B1(n13731), .B2(n15195), .A(n13249), .ZN(n13250) );
  OAI21_X1 U15461 ( .B1(n13251), .B2(n13349), .A(n13250), .ZN(P2_U3191) );
  NAND2_X1 U15462 ( .A1(n13253), .A2(n13252), .ZN(n13259) );
  NOR2_X1 U15463 ( .A1(n13254), .A2(n13604), .ZN(n13256) );
  XOR2_X1 U15464 ( .A(n13256), .B(n13255), .Z(n13257) );
  XNOR2_X1 U15465 ( .A(n13455), .B(n13257), .ZN(n13258) );
  XNOR2_X1 U15466 ( .A(n13259), .B(n13258), .ZN(n13266) );
  NAND2_X1 U15467 ( .A1(n13336), .A2(n13356), .ZN(n13261) );
  NAND2_X1 U15468 ( .A1(n13337), .A2(n13357), .ZN(n13260) );
  NAND2_X1 U15469 ( .A1(n13261), .A2(n13260), .ZN(n13458) );
  OAI22_X1 U15470 ( .A1(n15198), .A2(n13449), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13262), .ZN(n13264) );
  NOR2_X1 U15471 ( .A1(n13762), .A2(n13331), .ZN(n13263) );
  AOI211_X1 U15472 ( .C1(n15190), .C2(n13458), .A(n13264), .B(n13263), .ZN(
        n13265) );
  OAI21_X1 U15473 ( .B1(n13266), .B2(n13349), .A(n13265), .ZN(P2_U3192) );
  OAI211_X1 U15474 ( .C1(n13269), .C2(n13268), .A(n13267), .B(n15193), .ZN(
        n13275) );
  OAI22_X1 U15475 ( .A1(n13271), .A2(n13301), .B1(n13270), .B2(n13303), .ZN(
        n13550) );
  OAI22_X1 U15476 ( .A1(n15198), .A2(n13558), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13272), .ZN(n13273) );
  AOI21_X1 U15477 ( .B1(n13550), .B2(n15190), .A(n13273), .ZN(n13274) );
  OAI211_X1 U15478 ( .C1(n7270), .C2(n13331), .A(n13275), .B(n13274), .ZN(
        P2_U3195) );
  INV_X1 U15479 ( .A(n13698), .ZN(n13498) );
  OAI211_X1 U15480 ( .C1(n13276), .C2(n13279), .A(n13278), .B(n15193), .ZN(
        n13286) );
  OAI22_X1 U15481 ( .A1(n13281), .A2(n13303), .B1(n13280), .B2(n13301), .ZN(
        n13493) );
  INV_X1 U15482 ( .A(n13496), .ZN(n13283) );
  OAI22_X1 U15483 ( .A1(n15198), .A2(n13283), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13282), .ZN(n13284) );
  AOI21_X1 U15484 ( .B1(n15190), .B2(n13493), .A(n13284), .ZN(n13285) );
  OAI211_X1 U15485 ( .C1(n13498), .C2(n13331), .A(n13286), .B(n13285), .ZN(
        P2_U3197) );
  AND3_X1 U15486 ( .A1(n14848), .A2(n13288), .A3(n13287), .ZN(n13289) );
  OAI21_X1 U15487 ( .B1(n13290), .B2(n13289), .A(n15193), .ZN(n13296) );
  OAI22_X1 U15488 ( .A1(n13292), .A2(n13301), .B1(n13291), .B2(n13303), .ZN(
        n13621) );
  OAI22_X1 U15489 ( .A1(n15198), .A2(n13626), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13293), .ZN(n13294) );
  AOI21_X1 U15490 ( .B1(n15190), .B2(n13621), .A(n13294), .ZN(n13295) );
  OAI211_X1 U15491 ( .C1(n7272), .C2(n13331), .A(n13296), .B(n13295), .ZN(
        P2_U3200) );
  OAI211_X1 U15492 ( .C1(n13297), .C2(n13300), .A(n13299), .B(n15193), .ZN(
        n13308) );
  OAI22_X1 U15493 ( .A1(n13304), .A2(n13303), .B1(n13302), .B2(n13301), .ZN(
        n13505) );
  INV_X1 U15494 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n13305) );
  OAI22_X1 U15495 ( .A1(n15198), .A2(n13512), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13305), .ZN(n13306) );
  AOI21_X1 U15496 ( .B1(n13505), .B2(n15190), .A(n13306), .ZN(n13307) );
  OAI211_X1 U15497 ( .C1(n6884), .C2(n13331), .A(n13308), .B(n13307), .ZN(
        P2_U3201) );
  AOI21_X1 U15498 ( .B1(n13311), .B2(n13310), .A(n13309), .ZN(n13315) );
  AOI22_X1 U15499 ( .A1(n13363), .A2(n13336), .B1(n13337), .B2(n13365), .ZN(
        n13566) );
  AOI22_X1 U15500 ( .A1(n13344), .A2(n13570), .B1(P2_REG3_REG_20__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13312) );
  OAI21_X1 U15501 ( .B1(n13347), .B2(n13566), .A(n13312), .ZN(n13313) );
  AOI21_X1 U15502 ( .B1(n13726), .B2(n15195), .A(n13313), .ZN(n13314) );
  OAI21_X1 U15503 ( .B1(n13315), .B2(n13349), .A(n13314), .ZN(P2_U3205) );
  INV_X1 U15504 ( .A(n13234), .ZN(n13316) );
  AOI21_X1 U15505 ( .B1(n13318), .B2(n13317), .A(n13316), .ZN(n13323) );
  AOI22_X1 U15506 ( .A1(n13361), .A2(n13336), .B1(n13337), .B2(n13363), .ZN(
        n13535) );
  INV_X1 U15507 ( .A(n13319), .ZN(n13538) );
  AOI22_X1 U15508 ( .A1(n13344), .A2(n13538), .B1(P2_REG3_REG_22__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13320) );
  OAI21_X1 U15509 ( .B1(n13535), .B2(n13347), .A(n13320), .ZN(n13321) );
  AOI21_X1 U15510 ( .B1(n13716), .B2(n15195), .A(n13321), .ZN(n13322) );
  OAI21_X1 U15511 ( .B1(n13323), .B2(n13349), .A(n13322), .ZN(P2_U3207) );
  INV_X1 U15512 ( .A(n13609), .ZN(n13739) );
  OAI211_X1 U15513 ( .C1(n13326), .C2(n13325), .A(n6830), .B(n15193), .ZN(
        n13330) );
  AND2_X1 U15514 ( .A1(P2_U3088), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n13410) );
  AND2_X1 U15515 ( .A1(n13367), .A2(n13337), .ZN(n13327) );
  AOI21_X1 U15516 ( .B1(n13365), .B2(n13336), .A(n13327), .ZN(n13601) );
  NOR2_X1 U15517 ( .A1(n13347), .A2(n13601), .ZN(n13328) );
  AOI211_X1 U15518 ( .C1(n13344), .C2(n13608), .A(n13410), .B(n13328), .ZN(
        n13329) );
  OAI211_X1 U15519 ( .C1(n13739), .C2(n13331), .A(n13330), .B(n13329), .ZN(
        P2_U3210) );
  INV_X1 U15520 ( .A(n13333), .ZN(n13334) );
  AOI21_X1 U15521 ( .B1(n13335), .B2(n13332), .A(n13334), .ZN(n13342) );
  AOI22_X1 U15522 ( .A1(n13337), .A2(n13359), .B1(n13336), .B2(n13357), .ZN(
        n13487) );
  INV_X1 U15523 ( .A(n13338), .ZN(n13482) );
  AOI22_X1 U15524 ( .A1(n13344), .A2(n13482), .B1(P2_REG3_REG_26__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13339) );
  OAI21_X1 U15525 ( .B1(n13347), .B2(n13487), .A(n13339), .ZN(n13340) );
  AOI21_X1 U15526 ( .B1(n13694), .B2(n15195), .A(n13340), .ZN(n13341) );
  OAI21_X1 U15527 ( .B1(n13342), .B2(n13349), .A(n13341), .ZN(P2_U3212) );
  INV_X1 U15528 ( .A(n13639), .ZN(n13343) );
  AOI22_X1 U15529 ( .A1(n13344), .A2(n13343), .B1(P2_REG3_REG_15__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13345) );
  OAI21_X1 U15530 ( .B1(n13347), .B2(n13346), .A(n13345), .ZN(n13353) );
  AOI211_X1 U15531 ( .C1(n13351), .C2(n13350), .A(n13349), .B(n13348), .ZN(
        n13352) );
  AOI211_X1 U15532 ( .C1(n13642), .C2(n15195), .A(n13353), .B(n13352), .ZN(
        n13354) );
  INV_X1 U15533 ( .A(n13354), .ZN(P2_U3213) );
  MUX2_X1 U15534 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n13436), .S(n6623), .Z(
        P2_U3562) );
  MUX2_X1 U15535 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n13355), .S(n6623), .Z(
        P2_U3561) );
  MUX2_X1 U15536 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n13356), .S(n6623), .Z(
        P2_U3560) );
  MUX2_X1 U15537 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n13357), .S(n6623), .Z(
        P2_U3558) );
  MUX2_X1 U15538 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n13358), .S(n6623), .Z(
        P2_U3557) );
  MUX2_X1 U15539 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n13359), .S(n6623), .Z(
        P2_U3556) );
  MUX2_X1 U15540 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n13360), .S(n6623), .Z(
        P2_U3555) );
  MUX2_X1 U15541 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(n13361), .S(n6623), .Z(
        P2_U3554) );
  MUX2_X1 U15542 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n13362), .S(n6623), .Z(
        P2_U3553) );
  MUX2_X1 U15543 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n13363), .S(n6623), .Z(
        P2_U3552) );
  MUX2_X1 U15544 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n13364), .S(n6623), .Z(
        P2_U3551) );
  MUX2_X1 U15545 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n13365), .S(n6623), .Z(
        P2_U3550) );
  MUX2_X1 U15546 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n13366), .S(n6623), .Z(
        P2_U3549) );
  MUX2_X1 U15547 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n13367), .S(n6623), .Z(
        P2_U3548) );
  MUX2_X1 U15548 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n13368), .S(n6623), .Z(
        P2_U3547) );
  MUX2_X1 U15549 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n13369), .S(n6623), .Z(
        P2_U3546) );
  MUX2_X1 U15550 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n13370), .S(n6623), .Z(
        P2_U3545) );
  MUX2_X1 U15551 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n13371), .S(n6623), .Z(
        P2_U3544) );
  MUX2_X1 U15552 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n13372), .S(n6623), .Z(
        P2_U3543) );
  MUX2_X1 U15553 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n13373), .S(n6623), .Z(
        P2_U3542) );
  MUX2_X1 U15554 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n13374), .S(n6623), .Z(
        P2_U3541) );
  MUX2_X1 U15555 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n13375), .S(n6623), .Z(
        P2_U3540) );
  MUX2_X1 U15556 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n13376), .S(n6623), .Z(
        P2_U3539) );
  MUX2_X1 U15557 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n13377), .S(n6623), .Z(
        P2_U3538) );
  MUX2_X1 U15558 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n13378), .S(n6623), .Z(
        P2_U3537) );
  MUX2_X1 U15559 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(n13379), .S(n6623), .Z(
        P2_U3536) );
  MUX2_X1 U15560 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n13380), .S(n6623), .Z(
        P2_U3535) );
  MUX2_X1 U15561 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(n13381), .S(n6623), .Z(
        P2_U3534) );
  MUX2_X1 U15562 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(n13382), .S(n6623), .Z(
        P2_U3533) );
  MUX2_X1 U15563 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n13383), .S(n6623), .Z(
        P2_U3532) );
  MUX2_X1 U15564 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n13384), .S(n6623), .Z(
        P2_U3531) );
  INV_X1 U15565 ( .A(n13385), .ZN(n13390) );
  NOR3_X1 U15566 ( .A1(n13388), .A2(n13387), .A3(n13386), .ZN(n13389) );
  NOR3_X1 U15567 ( .A1(n15298), .A2(n13390), .A3(n13389), .ZN(n13391) );
  AOI21_X1 U15568 ( .B1(n15318), .B2(n13392), .A(n13391), .ZN(n13399) );
  NOR2_X1 U15569 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8468), .ZN(n13393) );
  AOI21_X1 U15570 ( .B1(n15313), .B2(P2_ADDR_REG_7__SCAN_IN), .A(n13393), .ZN(
        n13398) );
  OAI211_X1 U15571 ( .C1(n13396), .C2(n13395), .A(n15307), .B(n13394), .ZN(
        n13397) );
  NAND3_X1 U15572 ( .A1(n13399), .A2(n13398), .A3(n13397), .ZN(P2_U3221) );
  INV_X1 U15573 ( .A(n13400), .ZN(n13402) );
  NAND2_X1 U15574 ( .A1(n13402), .A2(n13401), .ZN(n13403) );
  OAI21_X1 U15575 ( .B1(n13404), .B2(n8622), .A(n13403), .ZN(n13414) );
  XNOR2_X1 U15576 ( .A(n13415), .B(n13414), .ZN(n13405) );
  NOR2_X1 U15577 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n13405), .ZN(n13416) );
  AOI21_X1 U15578 ( .B1(n13405), .B2(P2_REG2_REG_18__SCAN_IN), .A(n13416), 
        .ZN(n13413) );
  AOI21_X1 U15579 ( .B1(n13407), .B2(P2_REG1_REG_17__SCAN_IN), .A(n13406), 
        .ZN(n13420) );
  XNOR2_X1 U15580 ( .A(n13419), .B(n13420), .ZN(n13408) );
  NOR2_X1 U15581 ( .A1(n13742), .A2(n13408), .ZN(n13421) );
  AOI211_X1 U15582 ( .C1(n13408), .C2(n13742), .A(n13421), .B(n15292), .ZN(
        n13409) );
  AOI211_X1 U15583 ( .C1(n13415), .C2(n15318), .A(n13410), .B(n13409), .ZN(
        n13412) );
  NAND2_X1 U15584 ( .A1(n15313), .A2(P2_ADDR_REG_18__SCAN_IN), .ZN(n13411) );
  OAI211_X1 U15585 ( .C1(n13413), .C2(n15298), .A(n13412), .B(n13411), .ZN(
        P2_U3232) );
  NOR2_X1 U15586 ( .A1(n13415), .A2(n13414), .ZN(n13417) );
  NOR2_X1 U15587 ( .A1(n13417), .A2(n13416), .ZN(n13418) );
  XOR2_X1 U15588 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n13418), .Z(n13424) );
  NOR2_X1 U15589 ( .A1(n13420), .A2(n13419), .ZN(n13422) );
  NOR2_X1 U15590 ( .A1(n13422), .A2(n13421), .ZN(n13423) );
  XNOR2_X1 U15591 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n13423), .ZN(n13427) );
  AOI22_X1 U15592 ( .A1(n13424), .A2(n15314), .B1(n15307), .B2(n13427), .ZN(
        n13431) );
  INV_X1 U15593 ( .A(n13424), .ZN(n13425) );
  AOI21_X1 U15594 ( .B1(n15314), .B2(n13425), .A(n15318), .ZN(n13426) );
  OAI21_X1 U15595 ( .B1(n13427), .B2(n15292), .A(n13426), .ZN(n13428) );
  INV_X1 U15596 ( .A(n13428), .ZN(n13430) );
  MUX2_X1 U15597 ( .A(n13431), .B(n13430), .S(n13429), .Z(n13433) );
  OAI211_X1 U15598 ( .C1(n13434), .C2(n15306), .A(n13433), .B(n13432), .ZN(
        P2_U3233) );
  NAND2_X1 U15599 ( .A1(n13757), .A2(n13441), .ZN(n13440) );
  XNOR2_X1 U15600 ( .A(n9128), .B(n13440), .ZN(n13435) );
  NAND2_X1 U15601 ( .A1(n13668), .A2(n15324), .ZN(n13439) );
  AND2_X1 U15602 ( .A1(n13437), .A2(n13436), .ZN(n13667) );
  INV_X1 U15603 ( .A(n13667), .ZN(n13671) );
  NOR2_X1 U15604 ( .A1(n6620), .A2(n13671), .ZN(n13443) );
  AOI21_X1 U15605 ( .B1(n6620), .B2(P2_REG2_REG_31__SCAN_IN), .A(n13443), .ZN(
        n13438) );
  OAI211_X1 U15606 ( .C1(n13753), .C2(n15330), .A(n13439), .B(n13438), .ZN(
        P2_U3234) );
  OAI211_X1 U15607 ( .C1(n13757), .C2(n13441), .A(n13604), .B(n13440), .ZN(
        n13672) );
  NOR2_X1 U15608 ( .A1(n13643), .A2(n13442), .ZN(n13444) );
  AOI211_X1 U15609 ( .C1(n13445), .C2(n13641), .A(n13444), .B(n13443), .ZN(
        n13446) );
  OAI21_X1 U15610 ( .B1(n13672), .B2(n13612), .A(n13446), .ZN(P2_U3235) );
  OAI22_X1 U15611 ( .A1(n13643), .A2(n13450), .B1(n13449), .B2(n13655), .ZN(
        n13454) );
  AOI21_X1 U15612 ( .B1(n13455), .B2(n6883), .A(n13651), .ZN(n13451) );
  NAND2_X1 U15613 ( .A1(n13452), .A2(n13451), .ZN(n13680) );
  NOR2_X1 U15614 ( .A1(n13680), .A2(n13612), .ZN(n13453) );
  AOI211_X1 U15615 ( .C1(n13641), .C2(n13455), .A(n13454), .B(n13453), .ZN(
        n13462) );
  AOI21_X1 U15616 ( .B1(n13457), .B2(n13456), .A(n13623), .ZN(n13460) );
  OR2_X1 U15617 ( .A1(n13681), .A2(n6620), .ZN(n13461) );
  OAI211_X1 U15618 ( .C1(n13682), .C2(n13592), .A(n13462), .B(n13461), .ZN(
        P2_U3237) );
  XNOR2_X1 U15619 ( .A(n13463), .B(n13474), .ZN(n13465) );
  AOI21_X1 U15620 ( .B1(n13465), .B2(n13661), .A(n13464), .ZN(n13690) );
  NAND2_X1 U15621 ( .A1(n13688), .A2(n13480), .ZN(n13466) );
  NAND2_X1 U15622 ( .A1(n13466), .A2(n13604), .ZN(n13467) );
  NOR2_X1 U15623 ( .A1(n13468), .A2(n13467), .ZN(n13687) );
  NAND2_X1 U15624 ( .A1(n13688), .A2(n13641), .ZN(n13472) );
  NOR2_X1 U15625 ( .A1(n13655), .A2(n13469), .ZN(n13470) );
  AOI21_X1 U15626 ( .B1(n6620), .B2(P2_REG2_REG_27__SCAN_IN), .A(n13470), .ZN(
        n13471) );
  NAND2_X1 U15627 ( .A1(n13472), .A2(n13471), .ZN(n13473) );
  AOI21_X1 U15628 ( .B1(n13687), .B2(n15324), .A(n13473), .ZN(n13477) );
  NAND2_X1 U15629 ( .A1(n13475), .A2(n13474), .ZN(n13685) );
  NAND3_X1 U15630 ( .A1(n13686), .A2(n13685), .A3(n15333), .ZN(n13476) );
  OAI211_X1 U15631 ( .C1(n13690), .C2(n6620), .A(n13477), .B(n13476), .ZN(
        P2_U3238) );
  XOR2_X1 U15632 ( .A(n13478), .B(n13486), .Z(n13696) );
  INV_X1 U15633 ( .A(n13480), .ZN(n13481) );
  AOI211_X1 U15634 ( .C1(n13694), .C2(n13495), .A(n13651), .B(n13481), .ZN(
        n13693) );
  AOI22_X1 U15635 ( .A1(n6620), .A2(P2_REG2_REG_26__SCAN_IN), .B1(n13482), 
        .B2(n15326), .ZN(n13483) );
  OAI21_X1 U15636 ( .B1(n8876), .B2(n15330), .A(n13483), .ZN(n13484) );
  AOI21_X1 U15637 ( .B1(n13693), .B2(n15324), .A(n13484), .ZN(n13490) );
  XOR2_X1 U15638 ( .A(n13486), .B(n13485), .Z(n13488) );
  OAI21_X1 U15639 ( .B1(n13488), .B2(n13623), .A(n13487), .ZN(n13692) );
  NAND2_X1 U15640 ( .A1(n13692), .A2(n13643), .ZN(n13489) );
  OAI211_X1 U15641 ( .C1(n13696), .C2(n13592), .A(n13490), .B(n13489), .ZN(
        P2_U3239) );
  XNOR2_X1 U15642 ( .A(n13492), .B(n13491), .ZN(n13494) );
  AOI21_X1 U15643 ( .B1(n13494), .B2(n13661), .A(n13493), .ZN(n13699) );
  AOI211_X1 U15644 ( .C1(n13698), .C2(n13514), .A(n13651), .B(n13479), .ZN(
        n13697) );
  AOI22_X1 U15645 ( .A1(n6620), .A2(P2_REG2_REG_25__SCAN_IN), .B1(n13496), 
        .B2(n15326), .ZN(n13497) );
  OAI21_X1 U15646 ( .B1(n13498), .B2(n15330), .A(n13497), .ZN(n13502) );
  XNOR2_X1 U15647 ( .A(n13499), .B(n13500), .ZN(n13701) );
  NOR2_X1 U15648 ( .A1(n13701), .A2(n13592), .ZN(n13501) );
  AOI211_X1 U15649 ( .C1(n13697), .C2(n15324), .A(n13502), .B(n13501), .ZN(
        n13503) );
  OAI21_X1 U15650 ( .B1(n6620), .B2(n13699), .A(n13503), .ZN(P2_U3240) );
  XNOR2_X1 U15651 ( .A(n13507), .B(n13504), .ZN(n13506) );
  AOI21_X1 U15652 ( .B1(n13506), .B2(n13661), .A(n13505), .ZN(n13705) );
  NAND2_X1 U15653 ( .A1(n13508), .A2(n13507), .ZN(n13509) );
  NAND2_X1 U15654 ( .A1(n13510), .A2(n13509), .ZN(n13706) );
  NAND2_X1 U15655 ( .A1(n6620), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n13511) );
  OAI21_X1 U15656 ( .B1(n13655), .B2(n13512), .A(n13511), .ZN(n13513) );
  AOI21_X1 U15657 ( .B1(n13703), .B2(n13641), .A(n13513), .ZN(n13517) );
  AOI21_X1 U15658 ( .B1(n13703), .B2(n13522), .A(n13651), .ZN(n13515) );
  AND2_X1 U15659 ( .A1(n13515), .A2(n13514), .ZN(n13702) );
  NAND2_X1 U15660 ( .A1(n13702), .A2(n15324), .ZN(n13516) );
  OAI211_X1 U15661 ( .C1(n13706), .C2(n13592), .A(n13517), .B(n13516), .ZN(
        n13518) );
  INV_X1 U15662 ( .A(n13518), .ZN(n13519) );
  OAI21_X1 U15663 ( .B1(n6620), .B2(n13705), .A(n13519), .ZN(P2_U3241) );
  INV_X1 U15664 ( .A(n13527), .ZN(n13520) );
  XNOR2_X1 U15665 ( .A(n13521), .B(n13520), .ZN(n13707) );
  OAI211_X1 U15666 ( .C1(n6734), .C2(n13770), .A(n13604), .B(n13522), .ZN(
        n13708) );
  AOI22_X1 U15667 ( .A1(n6620), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n13523), 
        .B2(n15326), .ZN(n13526) );
  NAND2_X1 U15668 ( .A1(n13524), .A2(n13641), .ZN(n13525) );
  OAI211_X1 U15669 ( .C1(n13708), .C2(n13612), .A(n13526), .B(n13525), .ZN(
        n13531) );
  XNOR2_X1 U15670 ( .A(n13528), .B(n13527), .ZN(n13529) );
  NAND2_X1 U15671 ( .A1(n13529), .A2(n13661), .ZN(n13710) );
  AOI21_X1 U15672 ( .B1(n13710), .B2(n13709), .A(n6620), .ZN(n13530) );
  AOI211_X1 U15673 ( .C1(n15333), .C2(n13707), .A(n13531), .B(n13530), .ZN(
        n13532) );
  INV_X1 U15674 ( .A(n13532), .ZN(P2_U3242) );
  XNOR2_X1 U15675 ( .A(n13534), .B(n13533), .ZN(n13537) );
  INV_X1 U15676 ( .A(n13535), .ZN(n13536) );
  AOI21_X1 U15677 ( .B1(n13537), .B2(n13661), .A(n13536), .ZN(n13717) );
  AOI211_X1 U15678 ( .C1(n13716), .C2(n13555), .A(n13651), .B(n6734), .ZN(
        n13715) );
  INV_X1 U15679 ( .A(n13716), .ZN(n13540) );
  AOI22_X1 U15680 ( .A1(n6620), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n13538), 
        .B2(n15326), .ZN(n13539) );
  OAI21_X1 U15681 ( .B1(n13540), .B2(n15330), .A(n13539), .ZN(n13546) );
  NAND2_X1 U15682 ( .A1(n13542), .A2(n13541), .ZN(n13543) );
  NAND2_X1 U15683 ( .A1(n13544), .A2(n13543), .ZN(n13719) );
  NOR2_X1 U15684 ( .A1(n13719), .A2(n13592), .ZN(n13545) );
  AOI211_X1 U15685 ( .C1(n13715), .C2(n15324), .A(n13546), .B(n13545), .ZN(
        n13547) );
  OAI21_X1 U15686 ( .B1(n6620), .B2(n13717), .A(n13547), .ZN(P2_U3243) );
  XNOR2_X1 U15687 ( .A(n13549), .B(n13548), .ZN(n13552) );
  INV_X1 U15688 ( .A(n13550), .ZN(n13551) );
  OAI21_X1 U15689 ( .B1(n13552), .B2(n13623), .A(n13551), .ZN(n13720) );
  INV_X1 U15690 ( .A(n13720), .ZN(n13564) );
  XNOR2_X1 U15691 ( .A(n13554), .B(n13553), .ZN(n13722) );
  INV_X1 U15692 ( .A(n13555), .ZN(n13556) );
  AOI211_X1 U15693 ( .C1(n13557), .C2(n13569), .A(n13651), .B(n13556), .ZN(
        n13721) );
  NAND2_X1 U15694 ( .A1(n13721), .A2(n15324), .ZN(n13561) );
  INV_X1 U15695 ( .A(n13558), .ZN(n13559) );
  AOI22_X1 U15696 ( .A1(n6620), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n13559), 
        .B2(n15326), .ZN(n13560) );
  OAI211_X1 U15697 ( .C1(n7270), .C2(n15330), .A(n13561), .B(n13560), .ZN(
        n13562) );
  AOI21_X1 U15698 ( .B1(n15333), .B2(n13722), .A(n13562), .ZN(n13563) );
  OAI21_X1 U15699 ( .B1(n6620), .B2(n13564), .A(n13563), .ZN(P2_U3244) );
  XNOR2_X1 U15700 ( .A(n13565), .B(n13573), .ZN(n13568) );
  INV_X1 U15701 ( .A(n13566), .ZN(n13567) );
  AOI21_X1 U15702 ( .B1(n13568), .B2(n13661), .A(n13567), .ZN(n13727) );
  AOI211_X1 U15703 ( .C1(n13726), .C2(n13589), .A(n13651), .B(n7271), .ZN(
        n13725) );
  AOI22_X1 U15704 ( .A1(n6620), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n13570), 
        .B2(n15326), .ZN(n13571) );
  OAI21_X1 U15705 ( .B1(n13572), .B2(n15330), .A(n13571), .ZN(n13576) );
  XOR2_X1 U15706 ( .A(n13574), .B(n13573), .Z(n13729) );
  NOR2_X1 U15707 ( .A1(n13729), .A2(n13592), .ZN(n13575) );
  AOI211_X1 U15708 ( .C1(n13725), .C2(n15324), .A(n13576), .B(n13575), .ZN(
        n13577) );
  OAI21_X1 U15709 ( .B1(n6620), .B2(n13727), .A(n13577), .ZN(P2_U3245) );
  XOR2_X1 U15710 ( .A(n13578), .B(n13581), .Z(n13580) );
  AOI21_X1 U15711 ( .B1(n13580), .B2(n13661), .A(n13579), .ZN(n13733) );
  XNOR2_X1 U15712 ( .A(n13582), .B(n13581), .ZN(n13735) );
  NAND2_X1 U15713 ( .A1(n6620), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n13583) );
  OAI21_X1 U15714 ( .B1(n13655), .B2(n13584), .A(n13583), .ZN(n13585) );
  AOI21_X1 U15715 ( .B1(n13731), .B2(n13641), .A(n13585), .ZN(n13591) );
  OR2_X1 U15716 ( .A1(n13606), .A2(n13586), .ZN(n13587) );
  AND3_X1 U15717 ( .A1(n13589), .A2(n13604), .A3(n13587), .ZN(n13730) );
  NAND2_X1 U15718 ( .A1(n13730), .A2(n15324), .ZN(n13590) );
  OAI211_X1 U15719 ( .C1(n13735), .C2(n13592), .A(n13591), .B(n13590), .ZN(
        n13593) );
  INV_X1 U15720 ( .A(n13593), .ZN(n13594) );
  OAI21_X1 U15721 ( .B1(n6620), .B2(n13733), .A(n13594), .ZN(P2_U3246) );
  XNOR2_X1 U15722 ( .A(n13596), .B(n13595), .ZN(n13603) );
  NAND2_X1 U15723 ( .A1(n13598), .A2(n13597), .ZN(n13599) );
  NAND2_X1 U15724 ( .A1(n13600), .A2(n13599), .ZN(n13736) );
  NAND2_X1 U15725 ( .A1(n13736), .A2(n15361), .ZN(n13602) );
  OAI211_X1 U15726 ( .C1(n13623), .C2(n13603), .A(n13602), .B(n13601), .ZN(
        n13741) );
  INV_X1 U15727 ( .A(n13741), .ZN(n13616) );
  NAND2_X1 U15728 ( .A1(n13609), .A2(n13632), .ZN(n13605) );
  NAND2_X1 U15729 ( .A1(n13605), .A2(n13604), .ZN(n13607) );
  OR2_X1 U15730 ( .A1(n13607), .A2(n13606), .ZN(n13737) );
  AOI22_X1 U15731 ( .A1(n6620), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n13608), 
        .B2(n15326), .ZN(n13611) );
  NAND2_X1 U15732 ( .A1(n13609), .A2(n13641), .ZN(n13610) );
  OAI211_X1 U15733 ( .C1(n13737), .C2(n13612), .A(n13611), .B(n13610), .ZN(
        n13613) );
  AOI21_X1 U15734 ( .B1(n13736), .B2(n13614), .A(n13613), .ZN(n13615) );
  OAI21_X1 U15735 ( .B1(n13616), .B2(n6620), .A(n13615), .ZN(P2_U3247) );
  INV_X1 U15736 ( .A(n13617), .ZN(n13618) );
  AOI21_X1 U15737 ( .B1(n13620), .B2(n13619), .A(n13618), .ZN(n13624) );
  INV_X1 U15738 ( .A(n13621), .ZN(n13622) );
  OAI21_X1 U15739 ( .B1(n13624), .B2(n13623), .A(n13622), .ZN(n13744) );
  NAND2_X1 U15740 ( .A1(n13744), .A2(n13643), .ZN(n13636) );
  NAND2_X1 U15741 ( .A1(n6620), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n13625) );
  OAI21_X1 U15742 ( .B1(n13655), .B2(n13626), .A(n13625), .ZN(n13627) );
  AOI21_X1 U15743 ( .B1(n13630), .B2(n13641), .A(n13627), .ZN(n13635) );
  XNOR2_X1 U15744 ( .A(n13629), .B(n13628), .ZN(n13746) );
  NAND2_X1 U15745 ( .A1(n13746), .A2(n15333), .ZN(n13634) );
  AOI21_X1 U15746 ( .B1(n13630), .B2(n6739), .A(n13651), .ZN(n13631) );
  AND2_X1 U15747 ( .A1(n13632), .A2(n13631), .ZN(n13745) );
  NAND2_X1 U15748 ( .A1(n13745), .A2(n15324), .ZN(n13633) );
  NAND4_X1 U15749 ( .A1(n13636), .A2(n13635), .A3(n13634), .A4(n13633), .ZN(
        P2_U3248) );
  NAND2_X1 U15750 ( .A1(n13637), .A2(n15333), .ZN(n13649) );
  NAND2_X1 U15751 ( .A1(n6620), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n13638) );
  OAI21_X1 U15752 ( .B1(n13655), .B2(n13639), .A(n13638), .ZN(n13640) );
  AOI21_X1 U15753 ( .B1(n13642), .B2(n13641), .A(n13640), .ZN(n13648) );
  NAND2_X1 U15754 ( .A1(n13644), .A2(n13643), .ZN(n13647) );
  NAND2_X1 U15755 ( .A1(n13645), .A2(n15324), .ZN(n13646) );
  NAND4_X1 U15756 ( .A1(n13649), .A2(n13648), .A3(n13647), .A4(n13646), .ZN(
        P2_U3250) );
  AOI211_X1 U15757 ( .C1(n15354), .C2(n13652), .A(n13651), .B(n13650), .ZN(
        n15353) );
  OAI21_X1 U15758 ( .B1(n13654), .B2(n6621), .A(n13653), .ZN(n15360) );
  AOI22_X1 U15759 ( .A1(n15324), .A2(n15353), .B1(n15333), .B2(n15360), .ZN(
        n13666) );
  INV_X1 U15760 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n13656) );
  OAI22_X1 U15761 ( .A1(n15330), .A2(n10651), .B1(n13656), .B2(n13655), .ZN(
        n13657) );
  INV_X1 U15762 ( .A(n13657), .ZN(n13665) );
  XNOR2_X1 U15763 ( .A(n13659), .B(n13658), .ZN(n13662) );
  AOI21_X1 U15764 ( .B1(n13662), .B2(n13661), .A(n13660), .ZN(n15352) );
  MUX2_X1 U15765 ( .A(n15352), .B(n13663), .S(n6620), .Z(n13664) );
  NAND3_X1 U15766 ( .A1(n13666), .A2(n13665), .A3(n13664), .ZN(P2_U3263) );
  INV_X1 U15767 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n13669) );
  NOR2_X1 U15768 ( .A1(n13668), .A2(n13667), .ZN(n13750) );
  MUX2_X1 U15769 ( .A(n13669), .B(n13750), .S(n15392), .Z(n13670) );
  OAI21_X1 U15770 ( .B1(n13753), .B2(n13749), .A(n13670), .ZN(P2_U3530) );
  INV_X1 U15771 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n13673) );
  AND2_X1 U15772 ( .A1(n13672), .A2(n13671), .ZN(n13754) );
  MUX2_X1 U15773 ( .A(n13673), .B(n13754), .S(n15392), .Z(n13674) );
  OAI21_X1 U15774 ( .B1(n13757), .B2(n13749), .A(n13674), .ZN(P2_U3529) );
  AOI21_X1 U15775 ( .B1(n15355), .B2(n13676), .A(n13675), .ZN(n13677) );
  OAI211_X1 U15776 ( .C1(n13734), .C2(n13679), .A(n13678), .B(n13677), .ZN(
        n13758) );
  MUX2_X1 U15777 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n13758), .S(n15392), .Z(
        P2_U3528) );
  OAI211_X1 U15778 ( .C1(n13682), .C2(n13734), .A(n13681), .B(n13680), .ZN(
        n13759) );
  MUX2_X1 U15779 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n13759), .S(n15392), .Z(
        n13683) );
  INV_X1 U15780 ( .A(n13683), .ZN(n13684) );
  NAND3_X1 U15781 ( .A1(n13686), .A2(n15381), .A3(n13685), .ZN(n13691) );
  AOI21_X1 U15782 ( .B1(n15355), .B2(n13688), .A(n13687), .ZN(n13689) );
  NAND3_X1 U15783 ( .A1(n13691), .A2(n13690), .A3(n13689), .ZN(n13763) );
  MUX2_X1 U15784 ( .A(n13763), .B(P2_REG1_REG_27__SCAN_IN), .S(n15389), .Z(
        P2_U3526) );
  AOI211_X1 U15785 ( .C1(n15355), .C2(n6882), .A(n13693), .B(n13692), .ZN(
        n13695) );
  OAI21_X1 U15786 ( .B1(n13734), .B2(n13696), .A(n13695), .ZN(n13764) );
  MUX2_X1 U15787 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n13764), .S(n15392), .Z(
        P2_U3525) );
  AOI21_X1 U15788 ( .B1(n15355), .B2(n13698), .A(n13697), .ZN(n13700) );
  OAI211_X1 U15789 ( .C1(n13734), .C2(n13701), .A(n13700), .B(n13699), .ZN(
        n13765) );
  MUX2_X1 U15790 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n13765), .S(n15392), .Z(
        P2_U3524) );
  AOI21_X1 U15791 ( .B1(n15355), .B2(n13703), .A(n13702), .ZN(n13704) );
  OAI211_X1 U15792 ( .C1(n13706), .C2(n13734), .A(n13705), .B(n13704), .ZN(
        n13766) );
  MUX2_X1 U15793 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n13766), .S(n15392), .Z(
        P2_U3523) );
  NAND2_X1 U15794 ( .A1(n13707), .A2(n15381), .ZN(n13712) );
  AND3_X1 U15795 ( .A1(n13710), .A2(n13709), .A3(n13708), .ZN(n13711) );
  NAND2_X1 U15796 ( .A1(n13712), .A2(n13711), .ZN(n13767) );
  MUX2_X1 U15797 ( .A(n13767), .B(P2_REG1_REG_23__SCAN_IN), .S(n15389), .Z(
        n13713) );
  INV_X1 U15798 ( .A(n13713), .ZN(n13714) );
  OAI21_X1 U15799 ( .B1(n13770), .B2(n13749), .A(n13714), .ZN(P2_U3522) );
  AOI21_X1 U15800 ( .B1(n15355), .B2(n13716), .A(n13715), .ZN(n13718) );
  OAI211_X1 U15801 ( .C1(n13734), .C2(n13719), .A(n13718), .B(n13717), .ZN(
        n13771) );
  MUX2_X1 U15802 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n13771), .S(n15392), .Z(
        P2_U3521) );
  AOI211_X1 U15803 ( .C1(n15381), .C2(n13722), .A(n13721), .B(n13720), .ZN(
        n13772) );
  MUX2_X1 U15804 ( .A(n13723), .B(n13772), .S(n15392), .Z(n13724) );
  OAI21_X1 U15805 ( .B1(n7270), .B2(n13749), .A(n13724), .ZN(P2_U3520) );
  AOI21_X1 U15806 ( .B1(n15355), .B2(n13726), .A(n13725), .ZN(n13728) );
  OAI211_X1 U15807 ( .C1(n13734), .C2(n13729), .A(n13728), .B(n13727), .ZN(
        n13775) );
  MUX2_X1 U15808 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n13775), .S(n15392), .Z(
        P2_U3519) );
  AOI21_X1 U15809 ( .B1(n15355), .B2(n13731), .A(n13730), .ZN(n13732) );
  OAI211_X1 U15810 ( .C1(n13735), .C2(n13734), .A(n13733), .B(n13732), .ZN(
        n13776) );
  MUX2_X1 U15811 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n13776), .S(n15392), .Z(
        P2_U3518) );
  INV_X1 U15812 ( .A(n15355), .ZN(n15378) );
  NAND2_X1 U15813 ( .A1(n13736), .A2(n8890), .ZN(n13738) );
  OAI211_X1 U15814 ( .C1(n13739), .C2(n15378), .A(n13738), .B(n13737), .ZN(
        n13740) );
  NOR2_X1 U15815 ( .A1(n13741), .A2(n13740), .ZN(n13777) );
  MUX2_X1 U15816 ( .A(n13742), .B(n13777), .S(n15392), .Z(n13743) );
  INV_X1 U15817 ( .A(n13743), .ZN(P2_U3517) );
  INV_X1 U15818 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n13747) );
  AOI211_X1 U15819 ( .C1(n15381), .C2(n13746), .A(n13745), .B(n13744), .ZN(
        n13780) );
  MUX2_X1 U15820 ( .A(n13747), .B(n13780), .S(n15392), .Z(n13748) );
  OAI21_X1 U15821 ( .B1(n7272), .B2(n13749), .A(n13748), .ZN(P2_U3516) );
  INV_X1 U15822 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n13751) );
  MUX2_X1 U15823 ( .A(n13751), .B(n13750), .S(n15383), .Z(n13752) );
  OAI21_X1 U15824 ( .B1(n13753), .B2(n13783), .A(n13752), .ZN(P2_U3498) );
  MUX2_X1 U15825 ( .A(n13755), .B(n13754), .S(n15383), .Z(n13756) );
  OAI21_X1 U15826 ( .B1(n13757), .B2(n13783), .A(n13756), .ZN(P2_U3497) );
  MUX2_X1 U15827 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n13758), .S(n15383), .Z(
        P2_U3496) );
  MUX2_X1 U15828 ( .A(n13759), .B(P2_REG0_REG_28__SCAN_IN), .S(n15382), .Z(
        n13760) );
  INV_X1 U15829 ( .A(n13760), .ZN(n13761) );
  OAI21_X1 U15830 ( .B1(n13762), .B2(n13783), .A(n13761), .ZN(P2_U3495) );
  MUX2_X1 U15831 ( .A(n13763), .B(P2_REG0_REG_27__SCAN_IN), .S(n15382), .Z(
        P2_U3494) );
  MUX2_X1 U15832 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n13764), .S(n15383), .Z(
        P2_U3493) );
  MUX2_X1 U15833 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n13765), .S(n15383), .Z(
        P2_U3492) );
  MUX2_X1 U15834 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n13766), .S(n15383), .Z(
        P2_U3491) );
  MUX2_X1 U15835 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n13767), .S(n15383), .Z(
        n13768) );
  INV_X1 U15836 ( .A(n13768), .ZN(n13769) );
  OAI21_X1 U15837 ( .B1(n13770), .B2(n13783), .A(n13769), .ZN(P2_U3490) );
  MUX2_X1 U15838 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n13771), .S(n15383), .Z(
        P2_U3489) );
  INV_X1 U15839 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n13773) );
  MUX2_X1 U15840 ( .A(n13773), .B(n13772), .S(n15383), .Z(n13774) );
  OAI21_X1 U15841 ( .B1(n7270), .B2(n13783), .A(n13774), .ZN(P2_U3488) );
  MUX2_X1 U15842 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n13775), .S(n15383), .Z(
        P2_U3487) );
  MUX2_X1 U15843 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n13776), .S(n15383), .Z(
        P2_U3486) );
  INV_X1 U15844 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n13778) );
  MUX2_X1 U15845 ( .A(n13778), .B(n13777), .S(n15383), .Z(n13779) );
  INV_X1 U15846 ( .A(n13779), .ZN(P2_U3484) );
  INV_X1 U15847 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n13781) );
  MUX2_X1 U15848 ( .A(n13781), .B(n13780), .S(n15383), .Z(n13782) );
  OAI21_X1 U15849 ( .B1(n7272), .B2(n13783), .A(n13782), .ZN(P2_U3481) );
  INV_X1 U15850 ( .A(n13784), .ZN(n13788) );
  NOR4_X1 U15851 ( .A1(n8365), .A2(P2_IR_REG_30__SCAN_IN), .A3(P2_U3088), .A4(
        n8803), .ZN(n13785) );
  AOI21_X1 U15852 ( .B1(n13786), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n13785), 
        .ZN(n13787) );
  OAI21_X1 U15853 ( .B1(n13788), .B2(n13804), .A(n13787), .ZN(P2_U3296) );
  INV_X1 U15854 ( .A(n13789), .ZN(n14763) );
  OAI222_X1 U15855 ( .A1(n13804), .A2(n14763), .B1(n13791), .B2(P2_U3088), 
        .C1(n13790), .C2(n13798), .ZN(P2_U3298) );
  NAND2_X1 U15856 ( .A1(n13793), .A2(n13792), .ZN(n13795) );
  OAI211_X1 U15857 ( .C1(n8218), .C2(n13798), .A(n13795), .B(n13794), .ZN(
        P2_U3299) );
  INV_X1 U15858 ( .A(n13796), .ZN(n14766) );
  OAI222_X1 U15859 ( .A1(n13798), .A2(n13797), .B1(n13804), .B2(n14766), .C1(
        P2_U3088), .C2(n8868), .ZN(P2_U3300) );
  INV_X1 U15860 ( .A(n13799), .ZN(n14769) );
  OAI222_X1 U15861 ( .A1(n13804), .A2(n14769), .B1(P2_U3088), .B2(n13801), 
        .C1(n13800), .C2(n13798), .ZN(P2_U3301) );
  INV_X1 U15862 ( .A(n13802), .ZN(n14772) );
  OAI222_X1 U15863 ( .A1(n13798), .A2(n13805), .B1(n13804), .B2(n14772), .C1(
        n13803), .C2(P2_U3088), .ZN(P2_U3302) );
  INV_X1 U15864 ( .A(n13806), .ZN(n13807) );
  MUX2_X1 U15865 ( .A(n13807), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3327) );
  XOR2_X1 U15866 ( .A(n13809), .B(n13808), .Z(n13815) );
  NAND2_X1 U15867 ( .A1(n14213), .A2(n14921), .ZN(n13811) );
  NAND2_X1 U15868 ( .A1(n14125), .A2(n14583), .ZN(n13810) );
  NAND2_X1 U15869 ( .A1(n13811), .A2(n13810), .ZN(n14396) );
  AOI22_X1 U15870 ( .A1(n13934), .A2(n14396), .B1(P1_REG3_REG_27__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13812) );
  OAI21_X1 U15871 ( .B1(n14400), .B2(n14914), .A(n13812), .ZN(n13813) );
  AOI21_X1 U15872 ( .B1(n14629), .B2(n14909), .A(n13813), .ZN(n13814) );
  OAI21_X1 U15873 ( .B1(n13815), .B2(n14904), .A(n13814), .ZN(P1_U3214) );
  XOR2_X1 U15874 ( .A(n13817), .B(n13816), .Z(n13823) );
  NAND2_X1 U15875 ( .A1(n14217), .A2(n14921), .ZN(n13819) );
  NAND2_X1 U15876 ( .A1(n14215), .A2(n14583), .ZN(n13818) );
  NAND2_X1 U15877 ( .A1(n13819), .A2(n13818), .ZN(n14460) );
  AOI22_X1 U15878 ( .A1(n14460), .A2(n13934), .B1(P1_REG3_REG_23__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13820) );
  OAI21_X1 U15879 ( .B1(n14467), .B2(n14914), .A(n13820), .ZN(n13821) );
  AOI21_X1 U15880 ( .B1(n14732), .B2(n14909), .A(n13821), .ZN(n13822) );
  OAI21_X1 U15881 ( .B1(n13823), .B2(n14904), .A(n13822), .ZN(P1_U3216) );
  OAI211_X1 U15882 ( .C1(n13826), .C2(n13825), .A(n13824), .B(n13912), .ZN(
        n13832) );
  AOI22_X1 U15883 ( .A1(n13943), .A2(n14230), .B1(n14909), .B2(n13984), .ZN(
        n13831) );
  AOI22_X1 U15884 ( .A1(n13827), .A2(n6624), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        P1_U3086), .ZN(n13830) );
  INV_X1 U15885 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n13828) );
  NAND2_X1 U15886 ( .A1(n13918), .A2(n13828), .ZN(n13829) );
  NAND4_X1 U15887 ( .A1(n13832), .A2(n13831), .A3(n13830), .A4(n13829), .ZN(
        P1_U3218) );
  AOI21_X1 U15888 ( .B1(n13834), .B2(n13833), .A(n14904), .ZN(n13836) );
  NAND2_X1 U15889 ( .A1(n13836), .A2(n13835), .ZN(n13842) );
  OR2_X1 U15890 ( .A1(n14085), .A2(n14919), .ZN(n13838) );
  NAND2_X1 U15891 ( .A1(n6943), .A2(n14921), .ZN(n13837) );
  NAND2_X1 U15892 ( .A1(n13838), .A2(n13837), .ZN(n14680) );
  NOR2_X1 U15893 ( .A1(n13839), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14338) );
  NOR2_X1 U15894 ( .A1(n14914), .A2(n14529), .ZN(n13840) );
  AOI211_X1 U15895 ( .C1(n14680), .C2(n13934), .A(n14338), .B(n13840), .ZN(
        n13841) );
  OAI211_X1 U15896 ( .C1(n6915), .C2(n13922), .A(n13842), .B(n13841), .ZN(
        P1_U3219) );
  INV_X1 U15897 ( .A(n13843), .ZN(n13844) );
  AOI21_X1 U15898 ( .B1(n13846), .B2(n13845), .A(n13844), .ZN(n13852) );
  NOR2_X1 U15899 ( .A1(n14914), .A2(n14501), .ZN(n13850) );
  NOR2_X1 U15900 ( .A1(n14085), .A2(n14601), .ZN(n13847) );
  AOI21_X1 U15901 ( .B1(n14217), .B2(n14583), .A(n13847), .ZN(n14497) );
  INV_X1 U15902 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n13848) );
  OAI22_X1 U15903 ( .A1(n14497), .A2(n13916), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13848), .ZN(n13849) );
  AOI211_X1 U15904 ( .C1(n14739), .C2(n14909), .A(n13850), .B(n13849), .ZN(
        n13851) );
  OAI21_X1 U15905 ( .B1(n13852), .B2(n14904), .A(n13851), .ZN(P1_U3223) );
  OAI21_X1 U15906 ( .B1(n14897), .B2(n14887), .A(n13853), .ZN(n13854) );
  AOI21_X1 U15907 ( .B1(n13943), .B2(n14221), .A(n13854), .ZN(n13855) );
  OAI21_X1 U15908 ( .B1(n13856), .B2(n14914), .A(n13855), .ZN(n13861) );
  AOI211_X1 U15909 ( .C1(n13859), .C2(n13858), .A(n14904), .B(n6827), .ZN(
        n13860) );
  AOI211_X1 U15910 ( .C1(n14040), .C2(n14909), .A(n13861), .B(n13860), .ZN(
        n13862) );
  INV_X1 U15911 ( .A(n13862), .ZN(P1_U3224) );
  XOR2_X1 U15912 ( .A(n13864), .B(n13863), .Z(n13870) );
  NAND2_X1 U15913 ( .A1(n14215), .A2(n14921), .ZN(n13866) );
  NAND2_X1 U15914 ( .A1(n14213), .A2(n14583), .ZN(n13865) );
  NAND2_X1 U15915 ( .A1(n13866), .A2(n13865), .ZN(n14426) );
  AOI22_X1 U15916 ( .A1(n13934), .A2(n14426), .B1(P1_REG3_REG_25__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13867) );
  OAI21_X1 U15917 ( .B1(n14433), .B2(n14914), .A(n13867), .ZN(n13868) );
  AOI21_X1 U15918 ( .B1(n14724), .B2(n14909), .A(n13868), .ZN(n13869) );
  OAI21_X1 U15919 ( .B1(n13870), .B2(n14904), .A(n13869), .ZN(P1_U3225) );
  XOR2_X1 U15920 ( .A(n13871), .B(n13872), .Z(n13877) );
  NOR2_X1 U15921 ( .A1(n14914), .A2(n14572), .ZN(n13875) );
  NAND2_X1 U15922 ( .A1(n13943), .A2(n14567), .ZN(n13873) );
  NAND2_X1 U15923 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n15039)
         );
  OAI211_X1 U15924 ( .C1(n14063), .C2(n14897), .A(n13873), .B(n15039), .ZN(
        n13874) );
  AOI211_X1 U15925 ( .C1(n14705), .C2(n14909), .A(n13875), .B(n13874), .ZN(
        n13876) );
  OAI21_X1 U15926 ( .B1(n13877), .B2(n14904), .A(n13876), .ZN(P1_U3226) );
  XOR2_X1 U15927 ( .A(n13878), .B(n13879), .Z(n13884) );
  NAND2_X1 U15928 ( .A1(n13943), .A2(n14582), .ZN(n13880) );
  NAND2_X1 U15929 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n15053)
         );
  OAI211_X1 U15930 ( .C1(n14551), .C2(n14897), .A(n13880), .B(n15053), .ZN(
        n13882) );
  NOR2_X1 U15931 ( .A1(n14556), .A2(n13922), .ZN(n13881) );
  AOI211_X1 U15932 ( .C1(n13918), .C2(n14552), .A(n13882), .B(n13881), .ZN(
        n13883) );
  OAI21_X1 U15933 ( .B1(n13884), .B2(n14904), .A(n13883), .ZN(P1_U3228) );
  XOR2_X1 U15934 ( .A(n13886), .B(n13885), .Z(n13892) );
  NAND2_X1 U15935 ( .A1(n14216), .A2(n14921), .ZN(n13888) );
  NAND2_X1 U15936 ( .A1(n14214), .A2(n14583), .ZN(n13887) );
  NAND2_X1 U15937 ( .A1(n13888), .A2(n13887), .ZN(n14444) );
  AOI22_X1 U15938 ( .A1(n14444), .A2(n13934), .B1(P1_REG3_REG_24__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13889) );
  OAI21_X1 U15939 ( .B1(n14452), .B2(n14914), .A(n13889), .ZN(n13890) );
  AOI21_X1 U15940 ( .B1(n14728), .B2(n14909), .A(n13890), .ZN(n13891) );
  OAI21_X1 U15941 ( .B1(n13892), .B2(n14904), .A(n13891), .ZN(P1_U3229) );
  OAI211_X1 U15942 ( .C1(n13895), .C2(n13894), .A(n13893), .B(n13912), .ZN(
        n13899) );
  AOI22_X1 U15943 ( .A1(n14218), .A2(n14583), .B1(n14921), .B2(n14545), .ZN(
        n14672) );
  OAI22_X1 U15944 ( .A1(n14672), .A2(n13916), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13896), .ZN(n13897) );
  AOI21_X1 U15945 ( .B1(n14513), .B2(n13918), .A(n13897), .ZN(n13898) );
  OAI211_X1 U15946 ( .C1(n14674), .C2(n13922), .A(n13899), .B(n13898), .ZN(
        P1_U3233) );
  AOI21_X1 U15947 ( .B1(n13900), .B2(n13901), .A(n14904), .ZN(n13902) );
  NAND2_X1 U15948 ( .A1(n13902), .A2(n14890), .ZN(n13908) );
  NOR2_X1 U15949 ( .A1(n14914), .A2(n13903), .ZN(n13906) );
  NAND2_X1 U15950 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3086), .ZN(n14994)
         );
  OAI21_X1 U15951 ( .B1(n14897), .B2(n13904), .A(n14994), .ZN(n13905) );
  AOI211_X1 U15952 ( .C1(n13943), .C2(n14220), .A(n13906), .B(n13905), .ZN(
        n13907) );
  OAI211_X1 U15953 ( .C1(n14044), .C2(n13922), .A(n13908), .B(n13907), .ZN(
        P1_U3234) );
  OAI21_X1 U15954 ( .B1(n13911), .B2(n13910), .A(n13909), .ZN(n13913) );
  NAND2_X1 U15955 ( .A1(n13913), .A2(n13912), .ZN(n13921) );
  INV_X1 U15956 ( .A(n14479), .ZN(n13919) );
  AND2_X1 U15957 ( .A1(n14218), .A2(n14921), .ZN(n13914) );
  AOI21_X1 U15958 ( .B1(n14216), .B2(n14583), .A(n13914), .ZN(n14663) );
  INV_X1 U15959 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n13915) );
  OAI22_X1 U15960 ( .A1(n14663), .A2(n13916), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13915), .ZN(n13917) );
  AOI21_X1 U15961 ( .B1(n13919), .B2(n13918), .A(n13917), .ZN(n13920) );
  OAI211_X1 U15962 ( .C1(n13922), .C2(n14738), .A(n13921), .B(n13920), .ZN(
        P1_U3235) );
  XOR2_X1 U15963 ( .A(n13923), .B(n13924), .Z(n13929) );
  NOR2_X1 U15964 ( .A1(n14914), .A2(n14538), .ZN(n13927) );
  NAND2_X1 U15965 ( .A1(n13943), .A2(n14566), .ZN(n13925) );
  NAND2_X1 U15966 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n15068)
         );
  OAI211_X1 U15967 ( .C1(n14062), .C2(n14897), .A(n13925), .B(n15068), .ZN(
        n13926) );
  AOI211_X1 U15968 ( .C1(n14537), .C2(n14909), .A(n13927), .B(n13926), .ZN(
        n13928) );
  OAI21_X1 U15969 ( .B1(n13929), .B2(n14904), .A(n13928), .ZN(P1_U3238) );
  XOR2_X1 U15970 ( .A(n13931), .B(n13930), .Z(n13938) );
  NAND2_X1 U15971 ( .A1(n14214), .A2(n14921), .ZN(n13933) );
  NAND2_X1 U15972 ( .A1(n14377), .A2(n14583), .ZN(n13932) );
  NAND2_X1 U15973 ( .A1(n13933), .A2(n13932), .ZN(n14415) );
  AOI22_X1 U15974 ( .A1(n13934), .A2(n14415), .B1(P1_REG3_REG_26__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13935) );
  OAI21_X1 U15975 ( .B1(n14416), .B2(n14914), .A(n13935), .ZN(n13936) );
  AOI21_X1 U15976 ( .B1(n14419), .B2(n14909), .A(n13936), .ZN(n13937) );
  OAI21_X1 U15977 ( .B1(n13938), .B2(n14904), .A(n13937), .ZN(P1_U3240) );
  NAND2_X1 U15978 ( .A1(n13939), .A2(n13940), .ZN(n13942) );
  XNOR2_X1 U15979 ( .A(n13942), .B(n13941), .ZN(n13948) );
  NOR2_X1 U15980 ( .A1(n14914), .A2(n14585), .ZN(n13946) );
  NAND2_X1 U15981 ( .A1(n13943), .A2(n14584), .ZN(n13944) );
  NAND2_X1 U15982 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n15021)
         );
  OAI211_X1 U15983 ( .C1(n14550), .C2(n14897), .A(n13944), .B(n15021), .ZN(
        n13945) );
  AOI211_X1 U15984 ( .C1(n14590), .C2(n14909), .A(n13946), .B(n13945), .ZN(
        n13947) );
  OAI21_X1 U15985 ( .B1(n13948), .B2(n14904), .A(n13947), .ZN(P1_U3241) );
  INV_X1 U15986 ( .A(n13959), .ZN(n14156) );
  OAI21_X1 U15987 ( .B1(n14156), .B2(n14776), .A(n13949), .ZN(n13950) );
  AND2_X1 U15988 ( .A1(n13951), .A2(n13950), .ZN(n14160) );
  INV_X1 U15989 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n13952) );
  OR2_X1 U15990 ( .A1(n13953), .A2(n13952), .ZN(n13958) );
  INV_X1 U15991 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n14344) );
  OR2_X1 U15992 ( .A1(n13954), .A2(n14344), .ZN(n13957) );
  OR2_X1 U15993 ( .A1(n6617), .A2(n13955), .ZN(n13956) );
  AND3_X1 U15994 ( .A1(n13958), .A2(n13957), .A3(n13956), .ZN(n14347) );
  INV_X1 U15995 ( .A(n14347), .ZN(n14211) );
  NAND2_X1 U15996 ( .A1(n13960), .A2(n14155), .ZN(n14131) );
  NAND2_X1 U15997 ( .A1(n14131), .A2(n13959), .ZN(n14134) );
  NAND2_X1 U15998 ( .A1(n13960), .A2(n14156), .ZN(n13961) );
  NAND2_X1 U15999 ( .A1(n13784), .A2(n7767), .ZN(n13963) );
  OR2_X1 U16000 ( .A1(n8083), .A2(n14753), .ZN(n13962) );
  MUX2_X1 U16001 ( .A(n14211), .B(n14136), .S(n14711), .Z(n13964) );
  OR2_X1 U16002 ( .A1(n14091), .A2(n14347), .ZN(n14132) );
  NAND2_X1 U16003 ( .A1(n13964), .A2(n14132), .ZN(n14163) );
  MUX2_X1 U16004 ( .A(n13966), .B(n13965), .S(n13973), .Z(n13972) );
  NAND2_X1 U16005 ( .A1(n15098), .A2(n10390), .ZN(n13968) );
  NAND2_X1 U16006 ( .A1(n13968), .A2(n13967), .ZN(n13971) );
  NAND2_X1 U16007 ( .A1(n14091), .A2(n13976), .ZN(n13974) );
  AND2_X1 U16008 ( .A1(n13975), .A2(n13974), .ZN(n13979) );
  MUX2_X1 U16009 ( .A(n13976), .B(n15111), .S(n14091), .Z(n13977) );
  OAI21_X1 U16010 ( .B1(n13980), .B2(n13979), .A(n13977), .ZN(n13982) );
  NAND3_X1 U16011 ( .A1(n13980), .A2(n13979), .A3(n13978), .ZN(n13981) );
  NAND3_X1 U16012 ( .A1(n13982), .A2(n13981), .A3(n14170), .ZN(n13989) );
  NAND2_X1 U16013 ( .A1(n14136), .A2(n13983), .ZN(n13987) );
  NAND2_X1 U16014 ( .A1(n14091), .A2(n13984), .ZN(n13986) );
  MUX2_X1 U16015 ( .A(n13987), .B(n13986), .S(n13985), .Z(n13988) );
  NAND2_X1 U16016 ( .A1(n13989), .A2(n13988), .ZN(n13993) );
  MUX2_X1 U16017 ( .A(n6624), .B(n13990), .S(n14091), .Z(n13994) );
  NAND2_X1 U16018 ( .A1(n13993), .A2(n13994), .ZN(n13992) );
  MUX2_X1 U16019 ( .A(n13990), .B(n6624), .S(n14091), .Z(n13991) );
  NAND2_X1 U16020 ( .A1(n13992), .A2(n13991), .ZN(n13998) );
  INV_X1 U16021 ( .A(n13993), .ZN(n13996) );
  INV_X1 U16022 ( .A(n13994), .ZN(n13995) );
  NAND2_X1 U16023 ( .A1(n13996), .A2(n13995), .ZN(n13997) );
  NAND2_X1 U16024 ( .A1(n13998), .A2(n13997), .ZN(n14002) );
  MUX2_X1 U16025 ( .A(n13999), .B(n14227), .S(n14091), .Z(n14003) );
  NAND2_X1 U16026 ( .A1(n14002), .A2(n14003), .ZN(n14001) );
  MUX2_X1 U16027 ( .A(n13999), .B(n14227), .S(n14136), .Z(n14000) );
  NAND2_X1 U16028 ( .A1(n14001), .A2(n14000), .ZN(n14007) );
  INV_X1 U16029 ( .A(n14002), .ZN(n14005) );
  INV_X1 U16030 ( .A(n14003), .ZN(n14004) );
  MUX2_X1 U16031 ( .A(n14226), .B(n15083), .S(n14091), .Z(n14009) );
  MUX2_X1 U16032 ( .A(n15083), .B(n14226), .S(n14091), .Z(n14008) );
  MUX2_X1 U16033 ( .A(n14225), .B(n15141), .S(n14136), .Z(n14013) );
  NAND2_X1 U16034 ( .A1(n14012), .A2(n14013), .ZN(n14011) );
  MUX2_X1 U16035 ( .A(n14225), .B(n15141), .S(n14091), .Z(n14010) );
  NAND2_X1 U16036 ( .A1(n14011), .A2(n14010), .ZN(n14017) );
  INV_X1 U16037 ( .A(n14012), .ZN(n14015) );
  INV_X1 U16038 ( .A(n14013), .ZN(n14014) );
  NAND2_X1 U16039 ( .A1(n14015), .A2(n14014), .ZN(n14016) );
  MUX2_X1 U16040 ( .A(n14224), .B(n14018), .S(n14091), .Z(n14020) );
  MUX2_X1 U16041 ( .A(n14224), .B(n14018), .S(n14136), .Z(n14019) );
  MUX2_X1 U16042 ( .A(n14223), .B(n15156), .S(n14136), .Z(n14024) );
  NAND2_X1 U16043 ( .A1(n14023), .A2(n14024), .ZN(n14022) );
  MUX2_X1 U16044 ( .A(n14223), .B(n15156), .S(n14091), .Z(n14021) );
  NAND2_X1 U16045 ( .A1(n14022), .A2(n14021), .ZN(n14028) );
  INV_X1 U16046 ( .A(n14023), .ZN(n14026) );
  INV_X1 U16047 ( .A(n14024), .ZN(n14025) );
  NAND2_X1 U16048 ( .A1(n14026), .A2(n14025), .ZN(n14027) );
  MUX2_X1 U16049 ( .A(n14222), .B(n14029), .S(n14091), .Z(n14031) );
  MUX2_X1 U16050 ( .A(n14222), .B(n14029), .S(n14136), .Z(n14030) );
  MUX2_X1 U16051 ( .A(n14221), .B(n14910), .S(n14136), .Z(n14035) );
  NAND2_X1 U16052 ( .A1(n14034), .A2(n14035), .ZN(n14033) );
  MUX2_X1 U16053 ( .A(n14221), .B(n14910), .S(n14091), .Z(n14032) );
  NAND2_X1 U16054 ( .A1(n14033), .A2(n14032), .ZN(n14039) );
  INV_X1 U16055 ( .A(n14034), .ZN(n14037) );
  INV_X1 U16056 ( .A(n14035), .ZN(n14036) );
  NAND2_X1 U16057 ( .A1(n14037), .A2(n14036), .ZN(n14038) );
  MUX2_X1 U16058 ( .A(n14220), .B(n14040), .S(n14091), .Z(n14042) );
  MUX2_X1 U16059 ( .A(n14220), .B(n14040), .S(n14136), .Z(n14041) );
  MUX2_X1 U16060 ( .A(n14922), .B(n14043), .S(n14136), .Z(n14046) );
  MUX2_X1 U16061 ( .A(n14887), .B(n14044), .S(n14091), .Z(n14045) );
  OAI21_X1 U16062 ( .B1(n14047), .B2(n14046), .A(n14045), .ZN(n14049) );
  NAND2_X1 U16063 ( .A1(n14047), .A2(n14046), .ZN(n14048) );
  NAND2_X1 U16064 ( .A1(n14049), .A2(n14048), .ZN(n14050) );
  NAND2_X1 U16065 ( .A1(n14057), .A2(n14051), .ZN(n14052) );
  NAND2_X1 U16066 ( .A1(n14052), .A2(n14091), .ZN(n14054) );
  AOI21_X1 U16067 ( .B1(n14056), .B2(n14055), .A(n14091), .ZN(n14058) );
  OR3_X1 U16068 ( .A1(n14698), .A2(n14063), .A3(n14136), .ZN(n14060) );
  NAND3_X1 U16069 ( .A1(n14698), .A2(n14063), .A3(n14136), .ZN(n14059) );
  AND2_X1 U16070 ( .A1(n14060), .A2(n14059), .ZN(n14075) );
  MUX2_X1 U16071 ( .A(n14582), .B(n14705), .S(n14136), .Z(n14073) );
  NAND2_X1 U16072 ( .A1(n14705), .A2(n14091), .ZN(n14065) );
  NAND2_X1 U16073 ( .A1(n14136), .A2(n14582), .ZN(n14072) );
  NAND3_X1 U16074 ( .A1(n14073), .A2(n14065), .A3(n14072), .ZN(n14061) );
  OR2_X1 U16075 ( .A1(n14528), .A2(n14062), .ZN(n14081) );
  AOI21_X1 U16076 ( .B1(n14081), .B2(n14067), .A(n14091), .ZN(n14070) );
  NAND2_X1 U16077 ( .A1(n14698), .A2(n14063), .ZN(n14064) );
  OAI21_X1 U16078 ( .B1(n14073), .B2(n14065), .A(n14064), .ZN(n14066) );
  NAND3_X1 U16079 ( .A1(n14067), .A2(n14075), .A3(n14066), .ZN(n14068) );
  NAND2_X1 U16080 ( .A1(n14068), .A2(n14082), .ZN(n14069) );
  NOR2_X1 U16081 ( .A1(n14070), .A2(n14069), .ZN(n14080) );
  OAI21_X1 U16082 ( .B1(n14073), .B2(n14072), .A(n14071), .ZN(n14074) );
  NAND2_X1 U16083 ( .A1(n14075), .A2(n14074), .ZN(n14076) );
  NAND2_X1 U16084 ( .A1(n14076), .A2(n14078), .ZN(n14077) );
  OAI21_X1 U16085 ( .B1(n14091), .B2(n14078), .A(n14077), .ZN(n14079) );
  MUX2_X1 U16086 ( .A(n14082), .B(n14081), .S(n14091), .Z(n14083) );
  NAND2_X1 U16087 ( .A1(n14084), .A2(n14083), .ZN(n14088) );
  MUX2_X1 U16088 ( .A(n14085), .B(n14674), .S(n14091), .Z(n14087) );
  INV_X1 U16089 ( .A(n14085), .ZN(n14219) );
  MUX2_X1 U16090 ( .A(n14219), .B(n14518), .S(n14136), .Z(n14086) );
  OAI21_X1 U16091 ( .B1(n14088), .B2(n14087), .A(n14086), .ZN(n14090) );
  NAND2_X1 U16092 ( .A1(n14088), .A2(n14087), .ZN(n14089) );
  NAND2_X1 U16093 ( .A1(n14090), .A2(n14089), .ZN(n14093) );
  MUX2_X1 U16094 ( .A(n14218), .B(n14739), .S(n14136), .Z(n14094) );
  MUX2_X1 U16095 ( .A(n14218), .B(n14739), .S(n14091), .Z(n14092) );
  INV_X1 U16096 ( .A(n14094), .ZN(n14095) );
  MUX2_X1 U16097 ( .A(n14217), .B(n14481), .S(n14091), .Z(n14098) );
  MUX2_X1 U16098 ( .A(n14217), .B(n14481), .S(n14136), .Z(n14096) );
  MUX2_X1 U16099 ( .A(n14216), .B(n14732), .S(n14136), .Z(n14100) );
  MUX2_X1 U16100 ( .A(n14216), .B(n14732), .S(n14091), .Z(n14099) );
  MUX2_X1 U16101 ( .A(n14215), .B(n14728), .S(n14091), .Z(n14104) );
  MUX2_X1 U16102 ( .A(n14215), .B(n14728), .S(n14136), .Z(n14101) );
  NAND2_X1 U16103 ( .A1(n14102), .A2(n14101), .ZN(n14108) );
  INV_X1 U16104 ( .A(n14103), .ZN(n14106) );
  INV_X1 U16105 ( .A(n14104), .ZN(n14105) );
  NAND2_X1 U16106 ( .A1(n14106), .A2(n14105), .ZN(n14107) );
  NAND2_X1 U16107 ( .A1(n14108), .A2(n14107), .ZN(n14110) );
  MUX2_X1 U16108 ( .A(n14214), .B(n14724), .S(n14136), .Z(n14111) );
  MUX2_X1 U16109 ( .A(n14214), .B(n14724), .S(n14091), .Z(n14109) );
  INV_X1 U16110 ( .A(n14111), .ZN(n14112) );
  MUX2_X1 U16111 ( .A(n14213), .B(n14419), .S(n14091), .Z(n14115) );
  MUX2_X1 U16112 ( .A(n14213), .B(n14419), .S(n14136), .Z(n14113) );
  INV_X1 U16113 ( .A(n14115), .ZN(n14116) );
  MUX2_X1 U16114 ( .A(n14377), .B(n14629), .S(n14136), .Z(n14120) );
  NAND2_X1 U16115 ( .A1(n14119), .A2(n14120), .ZN(n14118) );
  MUX2_X1 U16116 ( .A(n14377), .B(n14629), .S(n14091), .Z(n14117) );
  NAND2_X1 U16117 ( .A1(n14118), .A2(n14117), .ZN(n14124) );
  INV_X1 U16118 ( .A(n14120), .ZN(n14121) );
  MUX2_X1 U16119 ( .A(n14125), .B(n14627), .S(n14091), .Z(n14140) );
  MUX2_X1 U16120 ( .A(n14125), .B(n14627), .S(n14136), .Z(n14126) );
  OR2_X1 U16121 ( .A1(n8083), .A2(n14759), .ZN(n14128) );
  INV_X1 U16122 ( .A(n14212), .ZN(n14130) );
  AOI21_X1 U16123 ( .B1(n14132), .B2(n14131), .A(n14130), .ZN(n14133) );
  NAND2_X1 U16124 ( .A1(n14347), .A2(n14134), .ZN(n14135) );
  AND2_X1 U16125 ( .A1(n14135), .A2(n14212), .ZN(n14137) );
  MUX2_X1 U16126 ( .A(n14137), .B(n14715), .S(n14136), .Z(n14147) );
  MUX2_X1 U16127 ( .A(n14138), .B(n14365), .S(n14091), .Z(n14144) );
  INV_X1 U16128 ( .A(n14138), .ZN(n14376) );
  MUX2_X1 U16129 ( .A(n14376), .B(n14139), .S(n14136), .Z(n14143) );
  AOI22_X1 U16130 ( .A1(n14149), .A2(n14147), .B1(n14144), .B2(n14143), .ZN(
        n14142) );
  INV_X1 U16131 ( .A(n14143), .ZN(n14146) );
  INV_X1 U16132 ( .A(n14144), .ZN(n14145) );
  NAND2_X1 U16133 ( .A1(n14146), .A2(n14145), .ZN(n14148) );
  NAND2_X1 U16134 ( .A1(n14149), .A2(n14148), .ZN(n14153) );
  INV_X1 U16135 ( .A(n14147), .ZN(n14152) );
  INV_X1 U16136 ( .A(n14148), .ZN(n14151) );
  INV_X1 U16137 ( .A(n14149), .ZN(n14150) );
  NAND3_X1 U16138 ( .A1(n14159), .A2(n14160), .A3(n14163), .ZN(n14157) );
  NAND2_X1 U16139 ( .A1(n14156), .A2(n14155), .ZN(n14200) );
  OAI211_X1 U16140 ( .C1(n14160), .C2(n14163), .A(n14157), .B(n14200), .ZN(
        n14158) );
  INV_X1 U16141 ( .A(n14158), .ZN(n14205) );
  XNOR2_X1 U16142 ( .A(n14711), .B(n14347), .ZN(n14198) );
  INV_X1 U16143 ( .A(n14198), .ZN(n14162) );
  INV_X1 U16144 ( .A(n14160), .ZN(n14161) );
  NOR2_X1 U16145 ( .A1(n14162), .A2(n14161), .ZN(n14164) );
  NOR2_X1 U16146 ( .A1(n14166), .A2(n14165), .ZN(n14204) );
  XOR2_X1 U16147 ( .A(n14212), .B(n14715), .Z(n14197) );
  INV_X1 U16148 ( .A(n14543), .ZN(n14189) );
  AND2_X1 U16149 ( .A1(n14168), .A2(n15098), .ZN(n14171) );
  NAND4_X1 U16150 ( .A1(n14172), .A2(n14171), .A3(n14170), .A4(n14169), .ZN(
        n14173) );
  NOR2_X1 U16151 ( .A1(n14174), .A2(n14173), .ZN(n14177) );
  NAND4_X1 U16152 ( .A1(n14178), .A2(n14177), .A3(n14176), .A4(n14175), .ZN(
        n14179) );
  NOR2_X1 U16153 ( .A1(n14607), .A2(n14179), .ZN(n14182) );
  NAND4_X1 U16154 ( .A1(n14183), .A2(n14182), .A3(n14181), .A4(n14180), .ZN(
        n14184) );
  NOR2_X1 U16155 ( .A1(n14931), .A2(n14184), .ZN(n14186) );
  NAND4_X1 U16156 ( .A1(n14187), .A2(n14592), .A3(n14186), .A4(n14185), .ZN(
        n14188) );
  NOR4_X1 U16157 ( .A1(n14523), .A2(n14560), .A3(n14189), .A4(n14188), .ZN(
        n14190) );
  NAND4_X1 U16158 ( .A1(n14191), .A2(n14512), .A3(n14190), .A4(n14496), .ZN(
        n14192) );
  NOR4_X1 U16159 ( .A1(n14430), .A2(n14441), .A3(n14463), .A4(n14192), .ZN(
        n14194) );
  NAND4_X1 U16160 ( .A1(n14372), .A2(n14194), .A3(n14411), .A4(n14193), .ZN(
        n14195) );
  NOR4_X1 U16161 ( .A1(n14198), .A2(n14197), .A3(n14196), .A4(n14195), .ZN(
        n14199) );
  XNOR2_X1 U16162 ( .A(n14199), .B(n14917), .ZN(n14202) );
  INV_X1 U16163 ( .A(n14200), .ZN(n14201) );
  NOR3_X1 U16164 ( .A1(n14206), .A2(n6625), .A3(n14601), .ZN(n14208) );
  OAI21_X1 U16165 ( .B1(n14209), .B2(n14776), .A(P1_B_REG_SCAN_IN), .ZN(n14207) );
  OAI22_X1 U16166 ( .A1(n14210), .A2(n14209), .B1(n14208), .B2(n14207), .ZN(
        P1_U3242) );
  MUX2_X1 U16167 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n14211), .S(n14232), .Z(
        P1_U3591) );
  MUX2_X1 U16168 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n14212), .S(P1_U4016), .Z(
        P1_U3590) );
  MUX2_X1 U16169 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n14376), .S(P1_U4016), .Z(
        P1_U3589) );
  MUX2_X1 U16170 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n14377), .S(P1_U4016), .Z(
        P1_U3587) );
  MUX2_X1 U16171 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n14213), .S(P1_U4016), .Z(
        P1_U3586) );
  MUX2_X1 U16172 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n14214), .S(P1_U4016), .Z(
        P1_U3585) );
  MUX2_X1 U16173 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n14215), .S(P1_U4016), .Z(
        P1_U3584) );
  MUX2_X1 U16174 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n14216), .S(P1_U4016), .Z(
        P1_U3583) );
  MUX2_X1 U16175 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n14217), .S(P1_U4016), .Z(
        P1_U3582) );
  MUX2_X1 U16176 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n14218), .S(P1_U4016), .Z(
        P1_U3581) );
  MUX2_X1 U16177 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n14219), .S(P1_U4016), .Z(
        P1_U3580) );
  MUX2_X1 U16178 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n14545), .S(P1_U4016), .Z(
        P1_U3579) );
  MUX2_X1 U16179 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n6943), .S(P1_U4016), .Z(
        P1_U3578) );
  MUX2_X1 U16180 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n14566), .S(P1_U4016), .Z(
        P1_U3577) );
  MUX2_X1 U16181 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n14582), .S(P1_U4016), .Z(
        P1_U3576) );
  MUX2_X1 U16182 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n14567), .S(P1_U4016), .Z(
        P1_U3575) );
  MUX2_X1 U16183 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n14584), .S(P1_U4016), .Z(
        P1_U3574) );
  MUX2_X1 U16184 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n14922), .S(P1_U4016), .Z(
        P1_U3573) );
  MUX2_X1 U16185 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n14220), .S(P1_U4016), .Z(
        P1_U3572) );
  MUX2_X1 U16186 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n14221), .S(P1_U4016), .Z(
        P1_U3571) );
  MUX2_X1 U16187 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n14222), .S(P1_U4016), .Z(
        P1_U3570) );
  MUX2_X1 U16188 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n14223), .S(P1_U4016), .Z(
        P1_U3569) );
  MUX2_X1 U16189 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n14224), .S(P1_U4016), .Z(
        P1_U3568) );
  MUX2_X1 U16190 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n14225), .S(P1_U4016), .Z(
        P1_U3567) );
  MUX2_X1 U16191 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n14226), .S(P1_U4016), .Z(
        P1_U3566) );
  MUX2_X1 U16192 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n14227), .S(P1_U4016), .Z(
        P1_U3565) );
  MUX2_X1 U16193 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n6624), .S(n14232), .Z(
        P1_U3564) );
  MUX2_X1 U16194 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n14229), .S(n14232), .Z(
        P1_U3563) );
  MUX2_X1 U16195 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n14230), .S(n14232), .Z(
        P1_U3562) );
  MUX2_X1 U16196 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n14231), .S(n14232), .Z(
        P1_U3561) );
  MUX2_X1 U16197 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n14233), .S(n14232), .Z(
        P1_U3560) );
  OAI211_X1 U16198 ( .C1(n14236), .C2(n14235), .A(n15012), .B(n14234), .ZN(
        n14244) );
  OAI211_X1 U16199 ( .C1(n14239), .C2(n14238), .A(n15015), .B(n14237), .ZN(
        n14243) );
  AOI22_X1 U16200 ( .A1(n14981), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n14242) );
  NAND2_X1 U16201 ( .A1(n15067), .A2(n14240), .ZN(n14241) );
  NAND4_X1 U16202 ( .A1(n14244), .A2(n14243), .A3(n14242), .A4(n14241), .ZN(
        P1_U3244) );
  AOI211_X1 U16203 ( .C1(n14247), .C2(n14246), .A(n14245), .B(n15056), .ZN(
        n14248) );
  INV_X1 U16204 ( .A(n14248), .ZN(n14258) );
  NAND2_X1 U16205 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_U3086), .ZN(n14249) );
  OAI21_X1 U16206 ( .B1(n15070), .B2(n14250), .A(n14249), .ZN(n14251) );
  AOI21_X1 U16207 ( .B1(n14252), .B2(n15067), .A(n14251), .ZN(n14257) );
  OAI211_X1 U16208 ( .C1(n14255), .C2(n14254), .A(n15012), .B(n14253), .ZN(
        n14256) );
  NAND3_X1 U16209 ( .A1(n14258), .A2(n14257), .A3(n14256), .ZN(P1_U3246) );
  OAI21_X1 U16210 ( .B1(n14261), .B2(n14260), .A(n14259), .ZN(n14262) );
  NAND2_X1 U16211 ( .A1(n14262), .A2(n15015), .ZN(n14272) );
  OAI21_X1 U16212 ( .B1(n15070), .B2(n14264), .A(n14263), .ZN(n14265) );
  AOI21_X1 U16213 ( .B1(n14266), .B2(n15067), .A(n14265), .ZN(n14271) );
  OAI211_X1 U16214 ( .C1(n14269), .C2(n14268), .A(n15012), .B(n14267), .ZN(
        n14270) );
  NAND3_X1 U16215 ( .A1(n14272), .A2(n14271), .A3(n14270), .ZN(P1_U3248) );
  OAI21_X1 U16216 ( .B1(n14275), .B2(n14274), .A(n14273), .ZN(n14276) );
  NAND2_X1 U16217 ( .A1(n14276), .A2(n15015), .ZN(n14286) );
  INV_X1 U16218 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n14278) );
  OAI21_X1 U16219 ( .B1(n15070), .B2(n14278), .A(n14277), .ZN(n14279) );
  AOI21_X1 U16220 ( .B1(n14280), .B2(n15067), .A(n14279), .ZN(n14285) );
  OAI211_X1 U16221 ( .C1(n14283), .C2(n14282), .A(n14281), .B(n15012), .ZN(
        n14284) );
  NAND3_X1 U16222 ( .A1(n14286), .A2(n14285), .A3(n14284), .ZN(P1_U3251) );
  OAI21_X1 U16223 ( .B1(n14289), .B2(n14288), .A(n14287), .ZN(n14290) );
  NAND2_X1 U16224 ( .A1(n14290), .A2(n15015), .ZN(n14300) );
  OAI21_X1 U16225 ( .B1(n15070), .B2(n14292), .A(n14291), .ZN(n14293) );
  AOI21_X1 U16226 ( .B1(n14294), .B2(n15067), .A(n14293), .ZN(n14299) );
  OAI211_X1 U16227 ( .C1(n14297), .C2(n14296), .A(n14295), .B(n15012), .ZN(
        n14298) );
  NAND3_X1 U16228 ( .A1(n14300), .A2(n14299), .A3(n14298), .ZN(P1_U3252) );
  XNOR2_X1 U16229 ( .A(n15052), .B(P1_REG2_REG_17__SCAN_IN), .ZN(n15048) );
  NAND2_X1 U16230 ( .A1(n14316), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n14301) );
  OAI21_X1 U16231 ( .B1(n14316), .B2(P1_REG2_REG_16__SCAN_IN), .A(n14301), 
        .ZN(n15029) );
  NAND2_X1 U16232 ( .A1(n15000), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n14307) );
  MUX2_X1 U16233 ( .A(P1_REG2_REG_13__SCAN_IN), .B(n11860), .S(n14993), .Z(
        n14302) );
  INV_X1 U16234 ( .A(n14302), .ZN(n14986) );
  OAI21_X1 U16235 ( .B1(n14319), .B2(P1_REG2_REG_12__SCAN_IN), .A(n14303), 
        .ZN(n14987) );
  NOR2_X1 U16236 ( .A1(n14986), .A2(n14987), .ZN(n14985) );
  AOI21_X1 U16237 ( .B1(n14993), .B2(P1_REG2_REG_13__SCAN_IN), .A(n14985), 
        .ZN(n15004) );
  INV_X1 U16238 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n14304) );
  MUX2_X1 U16239 ( .A(P1_REG2_REG_14__SCAN_IN), .B(n14304), .S(n15000), .Z(
        n14305) );
  INV_X1 U16240 ( .A(n14305), .ZN(n15003) );
  NOR2_X1 U16241 ( .A1(n15004), .A2(n15003), .ZN(n15002) );
  INV_X1 U16242 ( .A(n15002), .ZN(n14306) );
  NAND2_X1 U16243 ( .A1(n14307), .A2(n14306), .ZN(n14308) );
  INV_X1 U16244 ( .A(n14322), .ZN(n15019) );
  XNOR2_X1 U16245 ( .A(n14308), .B(n15019), .ZN(n15011) );
  NAND2_X1 U16246 ( .A1(n15011), .A2(n8008), .ZN(n14311) );
  INV_X1 U16247 ( .A(n14308), .ZN(n14309) );
  NAND2_X1 U16248 ( .A1(n14309), .A2(n15019), .ZN(n14310) );
  NAND2_X1 U16249 ( .A1(n14311), .A2(n14310), .ZN(n15030) );
  NOR2_X1 U16250 ( .A1(n15029), .A2(n15030), .ZN(n15031) );
  AOI21_X1 U16251 ( .B1(n14316), .B2(P1_REG2_REG_16__SCAN_IN), .A(n15031), 
        .ZN(n15049) );
  NOR2_X1 U16252 ( .A1(n15048), .A2(n15049), .ZN(n15047) );
  AOI21_X1 U16253 ( .B1(n15052), .B2(P1_REG2_REG_17__SCAN_IN), .A(n15047), 
        .ZN(n14312) );
  NOR2_X1 U16254 ( .A1(n14312), .A2(n14329), .ZN(n14313) );
  XNOR2_X1 U16255 ( .A(n14312), .B(n14329), .ZN(n15063) );
  NOR2_X1 U16256 ( .A1(n15062), .A2(n15063), .ZN(n15061) );
  XNOR2_X1 U16257 ( .A(P1_REG2_REG_19__SCAN_IN), .B(n14314), .ZN(n14336) );
  INV_X1 U16258 ( .A(n14336), .ZN(n14334) );
  INV_X1 U16259 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n15058) );
  INV_X1 U16260 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n14315) );
  XNOR2_X1 U16261 ( .A(n15052), .B(n14315), .ZN(n15043) );
  NAND2_X1 U16262 ( .A1(n14316), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n14327) );
  XNOR2_X1 U16263 ( .A(n14316), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n15024) );
  OR2_X1 U16264 ( .A1(n15000), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n14321) );
  MUX2_X1 U16265 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n14317), .S(n15000), .Z(
        n14999) );
  OAI21_X1 U16266 ( .B1(n14319), .B2(P1_REG1_REG_12__SCAN_IN), .A(n14318), 
        .ZN(n14990) );
  MUX2_X1 U16267 ( .A(n14320), .B(P1_REG1_REG_13__SCAN_IN), .S(n14993), .Z(
        n14989) );
  NOR2_X1 U16268 ( .A1(n14990), .A2(n14989), .ZN(n14988) );
  NAND2_X1 U16269 ( .A1(n14999), .A2(n14998), .ZN(n14997) );
  NAND2_X1 U16270 ( .A1(n14321), .A2(n14997), .ZN(n14323) );
  XNOR2_X1 U16271 ( .A(n14323), .B(n14322), .ZN(n15014) );
  NAND2_X1 U16272 ( .A1(n15014), .A2(n8007), .ZN(n14325) );
  NAND2_X1 U16273 ( .A1(n14323), .A2(n15019), .ZN(n14324) );
  NAND2_X1 U16274 ( .A1(n14325), .A2(n14324), .ZN(n15025) );
  NOR2_X1 U16275 ( .A1(n15024), .A2(n15025), .ZN(n15026) );
  INV_X1 U16276 ( .A(n15026), .ZN(n14326) );
  NAND2_X1 U16277 ( .A1(n14327), .A2(n14326), .ZN(n15042) );
  AND2_X1 U16278 ( .A1(n15052), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n14328) );
  XNOR2_X1 U16279 ( .A(n14330), .B(n14329), .ZN(n15059) );
  NOR2_X1 U16280 ( .A1(n15058), .A2(n15059), .ZN(n15057) );
  NOR2_X1 U16281 ( .A1(n14330), .A2(n14329), .ZN(n14331) );
  NOR2_X1 U16282 ( .A1(n15057), .A2(n14331), .ZN(n14332) );
  XNOR2_X1 U16283 ( .A(n14332), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n14335) );
  OAI21_X1 U16284 ( .B1(n14335), .B2(n15056), .A(n15037), .ZN(n14333) );
  AOI22_X1 U16285 ( .A1(n14336), .A2(n15012), .B1(n14335), .B2(n15015), .ZN(
        n14337) );
  INV_X1 U16286 ( .A(n14338), .ZN(n14339) );
  OAI211_X1 U16287 ( .C1(n14341), .C2(n15070), .A(n14340), .B(n14339), .ZN(
        P1_U3262) );
  XNOR2_X1 U16288 ( .A(n14342), .B(n14711), .ZN(n14343) );
  NAND2_X1 U16289 ( .A1(n14343), .A2(n15086), .ZN(n14618) );
  NOR2_X1 U16290 ( .A1(n14539), .A2(n14344), .ZN(n14348) );
  INV_X1 U16291 ( .A(n14345), .ZN(n14346) );
  OR2_X1 U16292 ( .A1(n14347), .A2(n14346), .ZN(n14621) );
  NOR2_X1 U16293 ( .A1(n15105), .A2(n14621), .ZN(n14354) );
  AOI211_X1 U16294 ( .C1(n14711), .C2(n15081), .A(n14348), .B(n14354), .ZN(
        n14349) );
  OAI21_X1 U16295 ( .B1(n14618), .B2(n14557), .A(n14349), .ZN(P1_U3263) );
  NAND2_X1 U16296 ( .A1(n14350), .A2(n14715), .ZN(n14351) );
  NAND3_X1 U16297 ( .A1(n14352), .A2(n15086), .A3(n14351), .ZN(n14622) );
  NOR2_X1 U16298 ( .A1(n14539), .A2(n14353), .ZN(n14355) );
  AOI211_X1 U16299 ( .C1(n14715), .C2(n15081), .A(n14355), .B(n14354), .ZN(
        n14356) );
  OAI21_X1 U16300 ( .B1(n14622), .B2(n14557), .A(n14356), .ZN(P1_U3264) );
  INV_X1 U16301 ( .A(n14357), .ZN(n14371) );
  AND2_X1 U16302 ( .A1(n14539), .A2(n14952), .ZN(n14561) );
  OAI22_X1 U16303 ( .A1(n14360), .A2(n14359), .B1(n14358), .B2(n14602), .ZN(
        n14363) );
  NOR2_X1 U16304 ( .A1(n15105), .A2(n14361), .ZN(n14362) );
  AOI211_X1 U16305 ( .C1(n15105), .C2(P1_REG2_REG_29__SCAN_IN), .A(n14363), 
        .B(n14362), .ZN(n14364) );
  OAI21_X1 U16306 ( .B1(n14365), .B2(n14570), .A(n14364), .ZN(n14368) );
  NOR2_X1 U16307 ( .A1(n14366), .A2(n14557), .ZN(n14367) );
  AOI211_X1 U16308 ( .C1(n14369), .C2(n14561), .A(n14368), .B(n14367), .ZN(
        n14370) );
  OAI21_X1 U16309 ( .B1(n14371), .B2(n15099), .A(n14370), .ZN(P1_U3356) );
  INV_X1 U16310 ( .A(n14372), .ZN(n14381) );
  NAND3_X1 U16311 ( .A1(n7567), .A2(n14381), .A3(n14373), .ZN(n14374) );
  NAND2_X1 U16312 ( .A1(n14376), .A2(n14583), .ZN(n14379) );
  INV_X1 U16313 ( .A(n14628), .ZN(n14389) );
  AND2_X1 U16314 ( .A1(n14627), .A2(n14403), .ZN(n14382) );
  OR3_X1 U16315 ( .A1(n14383), .A2(n14382), .A3(n14915), .ZN(n14625) );
  OAI22_X1 U16316 ( .A1(n14539), .A2(n14385), .B1(n14384), .B2(n14602), .ZN(
        n14386) );
  AOI21_X1 U16317 ( .B1(n14627), .B2(n15081), .A(n14386), .ZN(n14387) );
  OAI21_X1 U16318 ( .B1(n14625), .B2(n14557), .A(n14387), .ZN(n14388) );
  AOI21_X1 U16319 ( .B1(n14389), .B2(n14609), .A(n14388), .ZN(n14390) );
  OAI21_X1 U16320 ( .B1(n6724), .B2(n15105), .A(n14390), .ZN(P1_U3265) );
  OR2_X1 U16321 ( .A1(n14391), .A2(n14394), .ZN(n14392) );
  INV_X1 U16322 ( .A(n14630), .ZN(n14408) );
  NAND2_X1 U16323 ( .A1(n14630), .A2(n15162), .ZN(n14399) );
  AOI21_X1 U16324 ( .B1(n14397), .B2(n14952), .A(n14396), .ZN(n14398) );
  NAND2_X1 U16325 ( .A1(n14399), .A2(n14398), .ZN(n14634) );
  NAND2_X1 U16326 ( .A1(n14634), .A2(n14539), .ZN(n14407) );
  OAI22_X1 U16327 ( .A1(n14539), .A2(n14401), .B1(n14400), .B2(n14602), .ZN(
        n14405) );
  NAND2_X1 U16328 ( .A1(n14413), .A2(n14629), .ZN(n14402) );
  NAND3_X1 U16329 ( .A1(n14403), .A2(n15086), .A3(n14402), .ZN(n14631) );
  NOR2_X1 U16330 ( .A1(n14631), .A2(n14557), .ZN(n14404) );
  AOI211_X1 U16331 ( .C1(n15081), .C2(n14629), .A(n14405), .B(n14404), .ZN(
        n14406) );
  OAI211_X1 U16332 ( .C1(n14408), .C2(n15082), .A(n14407), .B(n14406), .ZN(
        P1_U3266) );
  XNOR2_X1 U16333 ( .A(n14410), .B(n14409), .ZN(n14643) );
  XNOR2_X1 U16334 ( .A(n14412), .B(n14411), .ZN(n14641) );
  OAI211_X1 U16335 ( .C1(n14639), .C2(n6639), .A(n15086), .B(n14413), .ZN(
        n14638) );
  NOR2_X1 U16336 ( .A1(n14539), .A2(n14414), .ZN(n14418) );
  INV_X1 U16337 ( .A(n14415), .ZN(n14637) );
  OAI22_X1 U16338 ( .A1(n15105), .A2(n14637), .B1(n14416), .B2(n14602), .ZN(
        n14417) );
  AOI211_X1 U16339 ( .C1(n14419), .C2(n15081), .A(n14418), .B(n14417), .ZN(
        n14420) );
  OAI21_X1 U16340 ( .B1(n14638), .B2(n14557), .A(n14420), .ZN(n14421) );
  AOI21_X1 U16341 ( .B1(n14641), .B2(n14609), .A(n14421), .ZN(n14422) );
  OAI21_X1 U16342 ( .B1(n14643), .B2(n15100), .A(n14422), .ZN(P1_U3267) );
  NAND2_X1 U16343 ( .A1(n14423), .A2(n14430), .ZN(n14424) );
  NAND2_X1 U16344 ( .A1(n14425), .A2(n14424), .ZN(n14427) );
  OAI21_X1 U16345 ( .B1(n14428), .B2(n14430), .A(n14429), .ZN(n14646) );
  INV_X1 U16346 ( .A(n14646), .ZN(n14438) );
  NAND2_X1 U16347 ( .A1(n14724), .A2(n14450), .ZN(n14431) );
  NAND2_X1 U16348 ( .A1(n14431), .A2(n15086), .ZN(n14432) );
  OR2_X1 U16349 ( .A1(n6639), .A2(n14432), .ZN(n14644) );
  OAI22_X1 U16350 ( .A1(n14539), .A2(n14434), .B1(n14433), .B2(n14602), .ZN(
        n14435) );
  AOI21_X1 U16351 ( .B1(n14724), .B2(n15081), .A(n14435), .ZN(n14436) );
  OAI21_X1 U16352 ( .B1(n14644), .B2(n14557), .A(n14436), .ZN(n14437) );
  AOI21_X1 U16353 ( .B1(n14438), .B2(n14609), .A(n14437), .ZN(n14439) );
  OAI21_X1 U16354 ( .B1(n15105), .B2(n14645), .A(n14439), .ZN(P1_U3268) );
  NAND2_X1 U16355 ( .A1(n14441), .A2(n14440), .ZN(n14442) );
  NAND3_X1 U16356 ( .A1(n14443), .A2(n14952), .A3(n14442), .ZN(n14446) );
  INV_X1 U16357 ( .A(n14444), .ZN(n14445) );
  AND2_X1 U16358 ( .A1(n14446), .A2(n14445), .ZN(n14651) );
  NAND2_X1 U16359 ( .A1(n14448), .A2(n14447), .ZN(n14449) );
  NAND2_X1 U16360 ( .A1(n6705), .A2(n14449), .ZN(n14649) );
  AOI21_X1 U16361 ( .B1(n14728), .B2(n14465), .A(n14915), .ZN(n14451) );
  NAND2_X1 U16362 ( .A1(n14451), .A2(n14450), .ZN(n14650) );
  OAI22_X1 U16363 ( .A1(n14539), .A2(n14453), .B1(n14452), .B2(n14602), .ZN(
        n14454) );
  AOI21_X1 U16364 ( .B1(n14728), .B2(n15081), .A(n14454), .ZN(n14455) );
  OAI21_X1 U16365 ( .B1(n14650), .B2(n14557), .A(n14455), .ZN(n14456) );
  AOI21_X1 U16366 ( .B1(n14649), .B2(n14609), .A(n14456), .ZN(n14457) );
  OAI21_X1 U16367 ( .B1(n15105), .B2(n14651), .A(n14457), .ZN(P1_U3269) );
  XNOR2_X1 U16368 ( .A(n14459), .B(n14458), .ZN(n14461) );
  AOI21_X1 U16369 ( .B1(n14461), .B2(n14952), .A(n14460), .ZN(n14656) );
  OAI21_X1 U16370 ( .B1(n14464), .B2(n14463), .A(n14462), .ZN(n14657) );
  INV_X1 U16371 ( .A(n14657), .ZN(n14472) );
  AOI21_X1 U16372 ( .B1(n14476), .B2(n14732), .A(n14915), .ZN(n14466) );
  NAND2_X1 U16373 ( .A1(n14466), .A2(n14465), .ZN(n14655) );
  INV_X1 U16374 ( .A(n14467), .ZN(n14468) );
  AOI22_X1 U16375 ( .A1(n14468), .A2(n15102), .B1(P1_REG2_REG_23__SCAN_IN), 
        .B2(n15105), .ZN(n14470) );
  NAND2_X1 U16376 ( .A1(n14732), .A2(n15081), .ZN(n14469) );
  OAI211_X1 U16377 ( .C1(n14655), .C2(n14557), .A(n14470), .B(n14469), .ZN(
        n14471) );
  AOI21_X1 U16378 ( .B1(n14472), .B2(n14609), .A(n14471), .ZN(n14473) );
  OAI21_X1 U16379 ( .B1(n15105), .B2(n14656), .A(n14473), .ZN(P1_U3270) );
  OAI21_X1 U16380 ( .B1(n14475), .B2(n14484), .A(n14474), .ZN(n14660) );
  AOI21_X1 U16381 ( .B1(n6735), .B2(n14481), .A(n14915), .ZN(n14477) );
  NAND2_X1 U16382 ( .A1(n14477), .A2(n14476), .ZN(n14661) );
  OAI22_X1 U16383 ( .A1(n14479), .A2(n14602), .B1(n14478), .B2(n14539), .ZN(
        n14480) );
  AOI21_X1 U16384 ( .B1(n14481), .B2(n15081), .A(n14480), .ZN(n14482) );
  OAI21_X1 U16385 ( .B1(n14661), .B2(n14557), .A(n14482), .ZN(n14490) );
  NAND2_X1 U16386 ( .A1(n14494), .A2(n14483), .ZN(n14485) );
  NAND2_X1 U16387 ( .A1(n14485), .A2(n14484), .ZN(n14487) );
  NAND2_X1 U16388 ( .A1(n14487), .A2(n14486), .ZN(n14488) );
  NAND2_X1 U16389 ( .A1(n14488), .A2(n14952), .ZN(n14662) );
  AOI21_X1 U16390 ( .B1(n14662), .B2(n14663), .A(n15105), .ZN(n14489) );
  AOI211_X1 U16391 ( .C1(n14609), .C2(n14660), .A(n14490), .B(n14489), .ZN(
        n14491) );
  INV_X1 U16392 ( .A(n14491), .ZN(P1_U3271) );
  INV_X1 U16393 ( .A(n14496), .ZN(n14492) );
  XNOR2_X1 U16394 ( .A(n14493), .B(n14492), .ZN(n14669) );
  OAI211_X1 U16395 ( .C1(n14496), .C2(n14495), .A(n14494), .B(n14952), .ZN(
        n14498) );
  AND2_X1 U16396 ( .A1(n14498), .A2(n14497), .ZN(n14668) );
  INV_X1 U16397 ( .A(n14668), .ZN(n14505) );
  AOI21_X1 U16398 ( .B1(n6738), .B2(n14739), .A(n14915), .ZN(n14499) );
  NAND2_X1 U16399 ( .A1(n14499), .A2(n6735), .ZN(n14667) );
  INV_X1 U16400 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n14500) );
  OAI22_X1 U16401 ( .A1(n14501), .A2(n14602), .B1(n14539), .B2(n14500), .ZN(
        n14502) );
  AOI21_X1 U16402 ( .B1(n14739), .B2(n15081), .A(n14502), .ZN(n14503) );
  OAI21_X1 U16403 ( .B1(n14667), .B2(n14557), .A(n14503), .ZN(n14504) );
  AOI21_X1 U16404 ( .B1(n14505), .B2(n14539), .A(n14504), .ZN(n14506) );
  OAI21_X1 U16405 ( .B1(n14669), .B2(n15099), .A(n14506), .ZN(P1_U3272) );
  OAI21_X1 U16406 ( .B1(n14512), .B2(n14508), .A(n14507), .ZN(n14678) );
  INV_X1 U16407 ( .A(n14509), .ZN(n14510) );
  AOI21_X1 U16408 ( .B1(n14512), .B2(n14511), .A(n14510), .ZN(n14676) );
  OAI211_X1 U16409 ( .C1(n14674), .C2(n14527), .A(n15086), .B(n6738), .ZN(
        n14673) );
  INV_X1 U16410 ( .A(n14672), .ZN(n14514) );
  AOI22_X1 U16411 ( .A1(n14514), .A2(n14539), .B1(n14513), .B2(n15102), .ZN(
        n14515) );
  OAI21_X1 U16412 ( .B1(n14516), .B2(n14539), .A(n14515), .ZN(n14517) );
  AOI21_X1 U16413 ( .B1(n14518), .B2(n15081), .A(n14517), .ZN(n14519) );
  OAI21_X1 U16414 ( .B1(n14673), .B2(n14557), .A(n14519), .ZN(n14520) );
  AOI21_X1 U16415 ( .B1(n14676), .B2(n14609), .A(n14520), .ZN(n14521) );
  OAI21_X1 U16416 ( .B1(n15100), .B2(n14678), .A(n14521), .ZN(P1_U3273) );
  XNOR2_X1 U16417 ( .A(n14522), .B(n14523), .ZN(n14679) );
  NAND2_X1 U16418 ( .A1(n14524), .A2(n14523), .ZN(n14525) );
  AOI21_X1 U16419 ( .B1(n14526), .B2(n14525), .A(n15075), .ZN(n14682) );
  OAI21_X1 U16420 ( .B1(n14682), .B2(n14680), .A(n14539), .ZN(n14534) );
  AOI211_X1 U16421 ( .C1(n14528), .C2(n14536), .A(n14915), .B(n14527), .ZN(
        n14681) );
  NOR2_X1 U16422 ( .A1(n6915), .A2(n14570), .ZN(n14532) );
  OAI22_X1 U16423 ( .A1(n14539), .A2(n14530), .B1(n14529), .B2(n14602), .ZN(
        n14531) );
  AOI211_X1 U16424 ( .C1(n14681), .C2(n15090), .A(n14532), .B(n14531), .ZN(
        n14533) );
  OAI211_X1 U16425 ( .C1(n14679), .C2(n15099), .A(n14534), .B(n14533), .ZN(
        P1_U3274) );
  XNOR2_X1 U16426 ( .A(n14535), .B(n14543), .ZN(n14693) );
  AOI211_X1 U16427 ( .C1(n14537), .C2(n14555), .A(n14915), .B(n6910), .ZN(
        n14690) );
  INV_X1 U16428 ( .A(n14537), .ZN(n14688) );
  NOR2_X1 U16429 ( .A1(n14688), .A2(n14570), .ZN(n14541) );
  OAI22_X1 U16430 ( .A1(n14539), .A2(n15062), .B1(n14538), .B2(n14602), .ZN(
        n14540) );
  AOI211_X1 U16431 ( .C1(n14690), .C2(n15090), .A(n14541), .B(n14540), .ZN(
        n14548) );
  OAI211_X1 U16432 ( .C1(n14544), .C2(n14543), .A(n14952), .B(n14542), .ZN(
        n14691) );
  AOI22_X1 U16433 ( .A1(n14545), .A2(n14583), .B1(n14566), .B2(n14921), .ZN(
        n14687) );
  AOI21_X1 U16434 ( .B1(n14691), .B2(n14687), .A(n15105), .ZN(n14546) );
  INV_X1 U16435 ( .A(n14546), .ZN(n14547) );
  OAI211_X1 U16436 ( .C1(n14693), .C2(n15099), .A(n14548), .B(n14547), .ZN(
        P1_U3275) );
  XNOR2_X1 U16437 ( .A(n14549), .B(n14560), .ZN(n14696) );
  INV_X1 U16438 ( .A(n14696), .ZN(n14564) );
  OAI22_X1 U16439 ( .A1(n14551), .A2(n14919), .B1(n14550), .B2(n14601), .ZN(
        n14697) );
  AOI21_X1 U16440 ( .B1(n14552), .B2(n15102), .A(n14697), .ZN(n14554) );
  NAND2_X1 U16441 ( .A1(n15105), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n14553) );
  OAI21_X1 U16442 ( .B1(n14554), .B2(n15105), .A(n14553), .ZN(n14559) );
  OAI211_X1 U16443 ( .C1(n14556), .C2(n14569), .A(n15086), .B(n14555), .ZN(
        n14699) );
  NOR2_X1 U16444 ( .A1(n14699), .A2(n14557), .ZN(n14558) );
  AOI211_X1 U16445 ( .C1(n15081), .C2(n14698), .A(n14559), .B(n14558), .ZN(
        n14563) );
  NAND2_X1 U16446 ( .A1(n6747), .A2(n14560), .ZN(n14695) );
  NAND3_X1 U16447 ( .A1(n14695), .A2(n14561), .A3(n14694), .ZN(n14562) );
  OAI211_X1 U16448 ( .C1(n14564), .C2(n15099), .A(n14563), .B(n14562), .ZN(
        P1_U3276) );
  XNOR2_X1 U16449 ( .A(n14565), .B(n14577), .ZN(n14568) );
  AOI222_X1 U16450 ( .A1(n14952), .A2(n14568), .B1(n14567), .B2(n14921), .C1(
        n14566), .C2(n14583), .ZN(n14707) );
  AOI211_X1 U16451 ( .C1(n14705), .C2(n14587), .A(n14915), .B(n14569), .ZN(
        n14704) );
  INV_X1 U16452 ( .A(n14705), .ZN(n14571) );
  NOR2_X1 U16453 ( .A1(n14571), .A2(n14570), .ZN(n14575) );
  INV_X1 U16454 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n14573) );
  OAI22_X1 U16455 ( .A1(n14539), .A2(n14573), .B1(n14572), .B2(n14602), .ZN(
        n14574) );
  AOI211_X1 U16456 ( .C1(n14704), .C2(n15090), .A(n14575), .B(n14574), .ZN(
        n14580) );
  OAI21_X1 U16457 ( .B1(n14578), .B2(n14577), .A(n14576), .ZN(n14703) );
  NAND2_X1 U16458 ( .A1(n14703), .A2(n14609), .ZN(n14579) );
  OAI211_X1 U16459 ( .C1(n14707), .C2(n15105), .A(n14580), .B(n14579), .ZN(
        P1_U3277) );
  OAI21_X1 U16460 ( .B1(n6742), .B2(n7104), .A(n14581), .ZN(n14943) );
  INV_X1 U16461 ( .A(n14943), .ZN(n14595) );
  AOI22_X1 U16462 ( .A1(n14584), .A2(n14921), .B1(n14583), .B2(n14582), .ZN(
        n14936) );
  OAI21_X1 U16463 ( .B1(n14585), .B2(n14602), .A(n14936), .ZN(n14586) );
  MUX2_X1 U16464 ( .A(P1_REG2_REG_15__SCAN_IN), .B(n14586), .S(n14539), .Z(
        n14589) );
  INV_X1 U16465 ( .A(n14590), .ZN(n14938) );
  OAI211_X1 U16466 ( .C1(n14938), .C2(n6736), .A(n14587), .B(n15086), .ZN(
        n14937) );
  NOR2_X1 U16467 ( .A1(n14937), .A2(n14557), .ZN(n14588) );
  AOI211_X1 U16468 ( .C1(n15081), .C2(n14590), .A(n14589), .B(n14588), .ZN(
        n14594) );
  INV_X1 U16469 ( .A(n14591), .ZN(n14939) );
  NOR2_X1 U16470 ( .A1(n6646), .A2(n14592), .ZN(n14940) );
  OR3_X1 U16471 ( .A1(n14939), .A2(n14940), .A3(n15100), .ZN(n14593) );
  OAI211_X1 U16472 ( .C1(n14595), .C2(n15099), .A(n14594), .B(n14593), .ZN(
        P1_U3278) );
  INV_X1 U16473 ( .A(n14596), .ZN(n14597) );
  AOI21_X1 U16474 ( .B1(n14607), .B2(n14598), .A(n14597), .ZN(n14599) );
  OAI222_X1 U16475 ( .A1(n14919), .A2(n14899), .B1(n14601), .B2(n14600), .C1(
        n15075), .C2(n14599), .ZN(n15153) );
  NAND2_X1 U16476 ( .A1(n15153), .A2(n14539), .ZN(n14617) );
  OAI22_X1 U16477 ( .A1(n14539), .A2(n14604), .B1(n14603), .B2(n14602), .ZN(
        n14606) );
  AOI21_X1 U16478 ( .B1(n15156), .B2(n15081), .A(n14606), .ZN(n14616) );
  XOR2_X1 U16479 ( .A(n14608), .B(n14607), .Z(n15158) );
  INV_X1 U16480 ( .A(n15158), .ZN(n15161) );
  NAND2_X1 U16481 ( .A1(n15161), .A2(n14609), .ZN(n14615) );
  NAND2_X1 U16482 ( .A1(n15156), .A2(n14610), .ZN(n14611) );
  NAND2_X1 U16483 ( .A1(n14611), .A2(n15086), .ZN(n14612) );
  NOR2_X1 U16484 ( .A1(n14613), .A2(n14612), .ZN(n15154) );
  NAND2_X1 U16485 ( .A1(n15154), .A2(n15090), .ZN(n14614) );
  NAND4_X1 U16486 ( .A1(n14617), .A2(n14616), .A3(n14615), .A4(n14614), .ZN(
        P1_U3284) );
  NAND2_X1 U16487 ( .A1(n14618), .A2(n14621), .ZN(n14709) );
  MUX2_X1 U16488 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n14709), .S(n15185), .Z(
        n14619) );
  AOI21_X1 U16489 ( .B1(n8887), .B2(n14711), .A(n14619), .ZN(n14620) );
  INV_X1 U16490 ( .A(n14620), .ZN(P1_U3559) );
  NAND2_X1 U16491 ( .A1(n14622), .A2(n14621), .ZN(n14713) );
  MUX2_X1 U16492 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n14713), .S(n15185), .Z(
        n14623) );
  AOI21_X1 U16493 ( .B1(n8887), .B2(n14715), .A(n14623), .ZN(n14624) );
  INV_X1 U16494 ( .A(n14624), .ZN(P1_U3558) );
  INV_X1 U16495 ( .A(n14625), .ZN(n14626) );
  MUX2_X1 U16496 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n14717), .S(n15185), .Z(
        P1_U3556) );
  INV_X1 U16497 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n14635) );
  NAND2_X1 U16498 ( .A1(n14630), .A2(n15137), .ZN(n14632) );
  NAND2_X1 U16499 ( .A1(n14632), .A2(n14631), .ZN(n14633) );
  MUX2_X1 U16500 ( .A(n14635), .B(n14718), .S(n15185), .Z(n14636) );
  INV_X1 U16501 ( .A(n15155), .ZN(n15166) );
  OAI211_X1 U16502 ( .C1(n14639), .C2(n15166), .A(n14638), .B(n14637), .ZN(
        n14640) );
  AOI21_X1 U16503 ( .B1(n14641), .B2(n15170), .A(n14640), .ZN(n14642) );
  OAI21_X1 U16504 ( .B1(n15075), .B2(n14643), .A(n14642), .ZN(n14721) );
  MUX2_X1 U16505 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n14721), .S(n15185), .Z(
        P1_U3554) );
  MUX2_X1 U16506 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n14722), .S(n15185), .Z(
        n14647) );
  AOI21_X1 U16507 ( .B1(n8887), .B2(n14724), .A(n14647), .ZN(n14648) );
  INV_X1 U16508 ( .A(n14648), .ZN(P1_U3553) );
  NAND2_X1 U16509 ( .A1(n14649), .A2(n15170), .ZN(n14652) );
  NAND3_X1 U16510 ( .A1(n14652), .A2(n14651), .A3(n14650), .ZN(n14726) );
  MUX2_X1 U16511 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n14726), .S(n15185), .Z(
        n14653) );
  AOI21_X1 U16512 ( .B1(n8887), .B2(n14728), .A(n14653), .ZN(n14654) );
  INV_X1 U16513 ( .A(n14654), .ZN(P1_U3552) );
  OAI211_X1 U16514 ( .C1(n14657), .C2(n14949), .A(n14656), .B(n14655), .ZN(
        n14730) );
  MUX2_X1 U16515 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n14730), .S(n15185), .Z(
        n14658) );
  AOI21_X1 U16516 ( .B1(n8887), .B2(n14732), .A(n14658), .ZN(n14659) );
  INV_X1 U16517 ( .A(n14659), .ZN(P1_U3551) );
  NAND2_X1 U16518 ( .A1(n14660), .A2(n15170), .ZN(n14664) );
  NAND4_X1 U16519 ( .A1(n14664), .A2(n14663), .A3(n14662), .A4(n14661), .ZN(
        n14735) );
  MUX2_X1 U16520 ( .A(n14735), .B(P1_REG1_REG_22__SCAN_IN), .S(n15183), .Z(
        n14665) );
  INV_X1 U16521 ( .A(n14665), .ZN(n14666) );
  OAI21_X1 U16522 ( .B1(n14686), .B2(n14738), .A(n14666), .ZN(P1_U3550) );
  OAI211_X1 U16523 ( .C1(n14949), .C2(n14669), .A(n14668), .B(n14667), .ZN(
        n14740) );
  MUX2_X1 U16524 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n14740), .S(n15185), .Z(
        n14670) );
  AOI21_X1 U16525 ( .B1(n8887), .B2(n14739), .A(n14670), .ZN(n14671) );
  INV_X1 U16526 ( .A(n14671), .ZN(P1_U3549) );
  OAI211_X1 U16527 ( .C1(n14674), .C2(n15166), .A(n14673), .B(n14672), .ZN(
        n14675) );
  AOI21_X1 U16528 ( .B1(n14676), .B2(n15170), .A(n14675), .ZN(n14677) );
  OAI21_X1 U16529 ( .B1(n15075), .B2(n14678), .A(n14677), .ZN(n14744) );
  MUX2_X1 U16530 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n14744), .S(n15185), .Z(
        P1_U3548) );
  INV_X1 U16531 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n14684) );
  NOR2_X1 U16532 ( .A1(n14679), .A2(n14949), .ZN(n14683) );
  NOR4_X1 U16533 ( .A1(n14683), .A2(n14682), .A3(n14681), .A4(n14680), .ZN(
        n14745) );
  MUX2_X1 U16534 ( .A(n14684), .B(n14745), .S(n15185), .Z(n14685) );
  OAI21_X1 U16535 ( .B1(n6915), .B2(n14686), .A(n14685), .ZN(P1_U3547) );
  OAI21_X1 U16536 ( .B1(n14688), .B2(n15166), .A(n14687), .ZN(n14689) );
  NOR2_X1 U16537 ( .A1(n14690), .A2(n14689), .ZN(n14692) );
  OAI211_X1 U16538 ( .C1(n14949), .C2(n14693), .A(n14692), .B(n14691), .ZN(
        n14749) );
  MUX2_X1 U16539 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n14749), .S(n15185), .Z(
        P1_U3546) );
  NAND3_X1 U16540 ( .A1(n14695), .A2(n14952), .A3(n14694), .ZN(n14702) );
  NAND2_X1 U16541 ( .A1(n14696), .A2(n15170), .ZN(n14701) );
  AOI21_X1 U16542 ( .B1(n14698), .B2(n15155), .A(n14697), .ZN(n14700) );
  NAND4_X1 U16543 ( .A1(n14702), .A2(n14701), .A3(n14700), .A4(n14699), .ZN(
        n14750) );
  MUX2_X1 U16544 ( .A(n14750), .B(P1_REG1_REG_17__SCAN_IN), .S(n15183), .Z(
        P1_U3545) );
  INV_X1 U16545 ( .A(n14703), .ZN(n14708) );
  AOI21_X1 U16546 ( .B1(n14705), .B2(n15155), .A(n14704), .ZN(n14706) );
  OAI211_X1 U16547 ( .C1(n14949), .C2(n14708), .A(n14707), .B(n14706), .ZN(
        n14751) );
  MUX2_X1 U16548 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n14751), .S(n15185), .Z(
        P1_U3544) );
  MUX2_X1 U16549 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n14709), .S(n15174), .Z(
        n14710) );
  AOI21_X1 U16550 ( .B1(n14733), .B2(n14711), .A(n14710), .ZN(n14712) );
  INV_X1 U16551 ( .A(n14712), .ZN(P1_U3527) );
  MUX2_X1 U16552 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n14713), .S(n15174), .Z(
        n14714) );
  AOI21_X1 U16553 ( .B1(n14733), .B2(n14715), .A(n14714), .ZN(n14716) );
  INV_X1 U16554 ( .A(n14716), .ZN(P1_U3526) );
  MUX2_X1 U16555 ( .A(n14719), .B(n14718), .S(n15174), .Z(n14720) );
  MUX2_X1 U16556 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n14721), .S(n15174), .Z(
        P1_U3522) );
  MUX2_X1 U16557 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n14722), .S(n15174), .Z(
        n14723) );
  AOI21_X1 U16558 ( .B1(n14733), .B2(n14724), .A(n14723), .ZN(n14725) );
  INV_X1 U16559 ( .A(n14725), .ZN(P1_U3521) );
  MUX2_X1 U16560 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n14726), .S(n15174), .Z(
        n14727) );
  AOI21_X1 U16561 ( .B1(n14733), .B2(n14728), .A(n14727), .ZN(n14729) );
  INV_X1 U16562 ( .A(n14729), .ZN(P1_U3520) );
  MUX2_X1 U16563 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n14730), .S(n15174), .Z(
        n14731) );
  AOI21_X1 U16564 ( .B1(n14733), .B2(n14732), .A(n14731), .ZN(n14734) );
  INV_X1 U16565 ( .A(n14734), .ZN(P1_U3519) );
  MUX2_X1 U16566 ( .A(n14735), .B(P1_REG0_REG_22__SCAN_IN), .S(n15172), .Z(
        n14736) );
  INV_X1 U16567 ( .A(n14736), .ZN(n14737) );
  OAI21_X1 U16568 ( .B1(n14748), .B2(n14738), .A(n14737), .ZN(P1_U3518) );
  INV_X1 U16569 ( .A(n14740), .ZN(n14742) );
  MUX2_X1 U16570 ( .A(n14742), .B(n14741), .S(n15172), .Z(n14743) );
  OAI21_X1 U16571 ( .B1(n6912), .B2(n14748), .A(n14743), .ZN(P1_U3517) );
  MUX2_X1 U16572 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n14744), .S(n15174), .Z(
        P1_U3516) );
  MUX2_X1 U16573 ( .A(n14746), .B(n14745), .S(n15174), .Z(n14747) );
  OAI21_X1 U16574 ( .B1(n6915), .B2(n14748), .A(n14747), .ZN(P1_U3515) );
  MUX2_X1 U16575 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n14749), .S(n15174), .Z(
        P1_U3513) );
  MUX2_X1 U16576 ( .A(n14750), .B(P1_REG0_REG_17__SCAN_IN), .S(n15172), .Z(
        P1_U3510) );
  MUX2_X1 U16577 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n14751), .S(n15174), .Z(
        P1_U3507) );
  NAND3_X1 U16578 ( .A1(n14752), .A2(P1_IR_REG_31__SCAN_IN), .A3(
        P1_STATE_REG_SCAN_IN), .ZN(n14754) );
  OAI22_X1 U16579 ( .A1(n14755), .A2(n14754), .B1(n14753), .B2(n14774), .ZN(
        n14756) );
  AOI21_X1 U16580 ( .B1(n13784), .B2(n14757), .A(n14756), .ZN(n14758) );
  INV_X1 U16581 ( .A(n14758), .ZN(P1_U3324) );
  OAI222_X1 U16582 ( .A1(n7705), .A2(P1_U3086), .B1(n14761), .B2(n14760), .C1(
        n14759), .C2(n14774), .ZN(P1_U3325) );
  OAI222_X1 U16583 ( .A1(P1_U3086), .A2(n14770), .B1(n14761), .B2(n14769), 
        .C1(n14768), .C2(n14774), .ZN(P1_U3329) );
  INV_X1 U16584 ( .A(n8325), .ZN(n14771) );
  MUX2_X1 U16585 ( .A(n14776), .B(n14775), .S(P1_U3086), .Z(P1_U3333) );
  INV_X1 U16586 ( .A(n14777), .ZN(n14778) );
  MUX2_X1 U16587 ( .A(n14778), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  OAI21_X1 U16588 ( .B1(n14781), .B2(n14780), .A(n14779), .ZN(n14782) );
  XNOR2_X1 U16589 ( .A(n14782), .B(P2_ADDR_REG_18__SCAN_IN), .ZN(SUB_1596_U62)
         );
  AOI21_X1 U16590 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n14783) );
  OAI21_X1 U16591 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(n14783), 
        .ZN(U28) );
  AOI21_X1 U16592 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(
        P3_RD_REG_SCAN_IN), .ZN(n14784) );
  OAI21_X1 U16593 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(n14784), 
        .ZN(U29) );
  OAI21_X1 U16594 ( .B1(n14787), .B2(n14786), .A(n14785), .ZN(n14788) );
  XNOR2_X1 U16595 ( .A(n14788), .B(P2_ADDR_REG_2__SCAN_IN), .ZN(SUB_1596_U61)
         );
  AOI21_X1 U16596 ( .B1(n14791), .B2(n14790), .A(n14789), .ZN(SUB_1596_U57) );
  OAI21_X1 U16597 ( .B1(n14794), .B2(n14793), .A(n14792), .ZN(SUB_1596_U55) );
  AOI22_X1 U16598 ( .A1(n14797), .A2(n14796), .B1(SI_18_), .B2(n14795), .ZN(
        n14798) );
  OAI21_X1 U16599 ( .B1(P3_U3151), .B2(n14799), .A(n14798), .ZN(P3_U3277) );
  OAI21_X1 U16600 ( .B1(n14802), .B2(n14801), .A(n14800), .ZN(n14803) );
  XNOR2_X1 U16601 ( .A(n14803), .B(P2_ADDR_REG_9__SCAN_IN), .ZN(SUB_1596_U54)
         );
  OAI222_X1 U16602 ( .A1(n15271), .A2(n14807), .B1(n15271), .B2(n14806), .C1(
        n14805), .C2(n14804), .ZN(SUB_1596_U70) );
  INV_X1 U16603 ( .A(n14808), .ZN(n14812) );
  OAI21_X1 U16604 ( .B1(n7084), .B2(n15166), .A(n14809), .ZN(n14811) );
  AOI211_X1 U16605 ( .C1(n15137), .C2(n14812), .A(n14811), .B(n14810), .ZN(
        n14813) );
  AOI22_X1 U16606 ( .A1(n15174), .A2(n14813), .B1(n7948), .B2(n15172), .ZN(
        P1_U3495) );
  AOI22_X1 U16607 ( .A1(n15185), .A2(n14813), .B1(n11270), .B2(n15183), .ZN(
        P1_U3540) );
  OAI21_X1 U16608 ( .B1(n14816), .B2(n14815), .A(n14814), .ZN(SUB_1596_U63) );
  INV_X1 U16609 ( .A(n14817), .ZN(n14819) );
  AOI21_X1 U16610 ( .B1(n14818), .B2(n15479), .A(n14819), .ZN(n14832) );
  AOI22_X1 U16611 ( .A1(n15498), .A2(n14832), .B1(n11248), .B2(n6791), .ZN(
        P3_U3490) );
  AOI21_X1 U16612 ( .B1(n14820), .B2(n15479), .A(n14819), .ZN(n14834) );
  AOI22_X1 U16613 ( .A1(n15498), .A2(n14834), .B1(n14821), .B2(n6791), .ZN(
        P3_U3489) );
  OAI22_X1 U16614 ( .A1(n14824), .A2(n14823), .B1(n15486), .B2(n14822), .ZN(
        n14825) );
  NOR2_X1 U16615 ( .A1(n14826), .A2(n14825), .ZN(n14836) );
  AOI22_X1 U16616 ( .A1(n15498), .A2(n14836), .B1(n9422), .B2(n6791), .ZN(
        P3_U3472) );
  NOR2_X1 U16617 ( .A1(n14827), .A2(n15486), .ZN(n14829) );
  AOI211_X1 U16618 ( .C1(n15477), .C2(n14830), .A(n14829), .B(n14828), .ZN(
        n14838) );
  AOI22_X1 U16619 ( .A1(n15498), .A2(n14838), .B1(n11663), .B2(n6791), .ZN(
        P3_U3471) );
  INV_X1 U16620 ( .A(P3_REG0_REG_31__SCAN_IN), .ZN(n14831) );
  AOI22_X1 U16621 ( .A1(n15493), .A2(n14832), .B1(n14831), .B2(n15491), .ZN(
        P3_U3458) );
  INV_X1 U16622 ( .A(P3_REG0_REG_30__SCAN_IN), .ZN(n14833) );
  AOI22_X1 U16623 ( .A1(n15493), .A2(n14834), .B1(n14833), .B2(n15491), .ZN(
        P3_U3457) );
  INV_X1 U16624 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n14835) );
  AOI22_X1 U16625 ( .A1(n15493), .A2(n14836), .B1(n14835), .B2(n15491), .ZN(
        P3_U3429) );
  AOI22_X1 U16626 ( .A1(n15493), .A2(n14838), .B1(n14837), .B2(n15491), .ZN(
        P3_U3426) );
  NAND2_X1 U16627 ( .A1(n14840), .A2(n14839), .ZN(n14841) );
  NAND2_X1 U16628 ( .A1(n14842), .A2(n14841), .ZN(n14843) );
  AOI222_X1 U16629 ( .A1(n15195), .A2(n14845), .B1(n14844), .B2(n15190), .C1(
        n14843), .C2(n15193), .ZN(n14846) );
  NAND2_X1 U16630 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3088), .ZN(n15321)
         );
  OAI211_X1 U16631 ( .C1(n15198), .C2(n14847), .A(n14846), .B(n15321), .ZN(
        P2_U3187) );
  OAI21_X1 U16632 ( .B1(n14850), .B2(n14849), .A(n14848), .ZN(n14851) );
  AOI222_X1 U16633 ( .A1(n15195), .A2(n14853), .B1(n14852), .B2(n15190), .C1(
        n14851), .C2(n15193), .ZN(n14855) );
  OAI211_X1 U16634 ( .C1(n15198), .C2(n14856), .A(n14855), .B(n14854), .ZN(
        P2_U3198) );
  INV_X1 U16635 ( .A(n14857), .ZN(n14862) );
  OAI211_X1 U16636 ( .C1(n14860), .C2(n15378), .A(n14859), .B(n14858), .ZN(
        n14861) );
  AOI211_X1 U16637 ( .C1(n14863), .C2(n15381), .A(n14862), .B(n14861), .ZN(
        n14882) );
  AOI22_X1 U16638 ( .A1(n15392), .A2(n14882), .B1(n14864), .B2(n15389), .ZN(
        P2_U3515) );
  OAI21_X1 U16639 ( .B1(n14866), .B2(n15378), .A(n14865), .ZN(n14867) );
  AOI211_X1 U16640 ( .C1(n14869), .C2(n15381), .A(n14868), .B(n14867), .ZN(
        n14883) );
  AOI22_X1 U16641 ( .A1(n15392), .A2(n14883), .B1(n11498), .B2(n15389), .ZN(
        P2_U3513) );
  OAI21_X1 U16642 ( .B1(n14871), .B2(n15378), .A(n14870), .ZN(n14873) );
  AOI211_X1 U16643 ( .C1(n15381), .C2(n14874), .A(n14873), .B(n14872), .ZN(
        n14885) );
  AOI22_X1 U16644 ( .A1(n15392), .A2(n14885), .B1(n11496), .B2(n15389), .ZN(
        P2_U3512) );
  OAI21_X1 U16645 ( .B1(n6888), .B2(n15378), .A(n14875), .ZN(n14876) );
  AOI21_X1 U16646 ( .B1(n14877), .B2(n8890), .A(n14876), .ZN(n14878) );
  AND2_X1 U16647 ( .A1(n14879), .A2(n14878), .ZN(n14886) );
  AOI22_X1 U16648 ( .A1(n15392), .A2(n14886), .B1(n14880), .B2(n15389), .ZN(
        P2_U3511) );
  INV_X1 U16649 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n14881) );
  AOI22_X1 U16650 ( .A1(n15383), .A2(n14882), .B1(n14881), .B2(n15382), .ZN(
        P2_U3478) );
  AOI22_X1 U16651 ( .A1(n15383), .A2(n14883), .B1(n8568), .B2(n15382), .ZN(
        P2_U3472) );
  INV_X1 U16652 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n14884) );
  AOI22_X1 U16653 ( .A1(n15383), .A2(n14885), .B1(n14884), .B2(n15382), .ZN(
        P2_U3469) );
  AOI22_X1 U16654 ( .A1(n15383), .A2(n14886), .B1(n8542), .B2(n15382), .ZN(
        P2_U3466) );
  OAI22_X1 U16655 ( .A1(n14900), .A2(n14887), .B1(n14920), .B2(n14897), .ZN(
        n14895) );
  AOI21_X1 U16656 ( .B1(n14890), .B2(n14889), .A(n14888), .ZN(n14891) );
  INV_X1 U16657 ( .A(n14891), .ZN(n14893) );
  AOI21_X1 U16658 ( .B1(n14893), .B2(n14892), .A(n14904), .ZN(n14894) );
  AOI211_X1 U16659 ( .C1(n14946), .C2(n14909), .A(n14895), .B(n14894), .ZN(
        n14896) );
  NAND2_X1 U16660 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n15008)
         );
  OAI211_X1 U16661 ( .C1(n14914), .C2(n14918), .A(n14896), .B(n15008), .ZN(
        P1_U3215) );
  OAI22_X1 U16662 ( .A1(n14900), .A2(n14899), .B1(n14898), .B2(n14897), .ZN(
        n14908) );
  AOI21_X1 U16663 ( .B1(n12182), .B2(n14902), .A(n14901), .ZN(n14903) );
  INV_X1 U16664 ( .A(n14903), .ZN(n14906) );
  AOI21_X1 U16665 ( .B1(n14906), .B2(n14905), .A(n14904), .ZN(n14907) );
  AOI211_X1 U16666 ( .C1(n14910), .C2(n14909), .A(n14908), .B(n14907), .ZN(
        n14912) );
  OAI211_X1 U16667 ( .C1(n14914), .C2(n14913), .A(n14912), .B(n14911), .ZN(
        P1_U3236) );
  AOI211_X1 U16668 ( .C1(n14946), .C2(n14916), .A(n14915), .B(n6736), .ZN(
        n14944) );
  NAND2_X1 U16669 ( .A1(n14944), .A2(n14917), .ZN(n14927) );
  INV_X1 U16670 ( .A(n14918), .ZN(n14925) );
  OR2_X1 U16671 ( .A1(n14920), .A2(n14919), .ZN(n14924) );
  NAND2_X1 U16672 ( .A1(n14922), .A2(n14921), .ZN(n14923) );
  NAND2_X1 U16673 ( .A1(n14924), .A2(n14923), .ZN(n14945) );
  AOI21_X1 U16674 ( .B1(n14925), .B2(n15102), .A(n14945), .ZN(n14926) );
  OAI211_X1 U16675 ( .C1(n8300), .C2(n14928), .A(n14927), .B(n14926), .ZN(
        n14934) );
  OAI21_X1 U16676 ( .B1(n6652), .B2(n14931), .A(n14929), .ZN(n14948) );
  XNOR2_X1 U16677 ( .A(n14931), .B(n14930), .ZN(n14951) );
  INV_X1 U16678 ( .A(n14951), .ZN(n14932) );
  OAI22_X1 U16679 ( .A1(n14948), .A2(n15099), .B1(n14932), .B2(n15100), .ZN(
        n14933) );
  AOI221_X1 U16680 ( .B1(P1_REG2_REG_14__SCAN_IN), .B2(n15105), .C1(n14934), 
        .C2(n14539), .A(n14933), .ZN(n14935) );
  INV_X1 U16681 ( .A(n14935), .ZN(P1_U3279) );
  OAI211_X1 U16682 ( .C1(n14938), .C2(n15166), .A(n14937), .B(n14936), .ZN(
        n14942) );
  NOR3_X1 U16683 ( .A1(n14940), .A2(n14939), .A3(n15075), .ZN(n14941) );
  AOI211_X1 U16684 ( .C1(n15170), .C2(n14943), .A(n14942), .B(n14941), .ZN(
        n14953) );
  AOI22_X1 U16685 ( .A1(n15185), .A2(n14953), .B1(n8007), .B2(n15183), .ZN(
        P1_U3543) );
  AOI211_X1 U16686 ( .C1(n14946), .C2(n15155), .A(n14945), .B(n14944), .ZN(
        n14947) );
  OAI21_X1 U16687 ( .B1(n14949), .B2(n14948), .A(n14947), .ZN(n14950) );
  AOI21_X1 U16688 ( .B1(n14952), .B2(n14951), .A(n14950), .ZN(n14954) );
  AOI22_X1 U16689 ( .A1(n15185), .A2(n14954), .B1(n14317), .B2(n15183), .ZN(
        P1_U3542) );
  AOI22_X1 U16690 ( .A1(n15174), .A2(n14953), .B1(n8009), .B2(n15172), .ZN(
        P1_U3504) );
  AOI22_X1 U16691 ( .A1(n15174), .A2(n14954), .B1(n7985), .B2(n15172), .ZN(
        P1_U3501) );
  OAI21_X1 U16692 ( .B1(n14957), .B2(n14956), .A(n14955), .ZN(n14958) );
  XNOR2_X1 U16693 ( .A(n14958), .B(P2_ADDR_REG_11__SCAN_IN), .ZN(SUB_1596_U69)
         );
  OAI21_X1 U16694 ( .B1(n14960), .B2(n15288), .A(n14959), .ZN(SUB_1596_U68) );
  OAI21_X1 U16695 ( .B1(n14963), .B2(n14962), .A(n14961), .ZN(n14964) );
  XNOR2_X1 U16696 ( .A(n14964), .B(P2_ADDR_REG_13__SCAN_IN), .ZN(SUB_1596_U67)
         );
  OAI21_X1 U16697 ( .B1(n14967), .B2(n14966), .A(n14965), .ZN(n14968) );
  XNOR2_X1 U16698 ( .A(n14968), .B(P2_ADDR_REG_14__SCAN_IN), .ZN(SUB_1596_U66)
         );
  OAI21_X1 U16699 ( .B1(n14971), .B2(n14970), .A(n14969), .ZN(n14972) );
  XNOR2_X1 U16700 ( .A(n14972), .B(P2_ADDR_REG_15__SCAN_IN), .ZN(SUB_1596_U65)
         );
  AOI21_X1 U16701 ( .B1(n14975), .B2(n14974), .A(n14973), .ZN(n14976) );
  XOR2_X1 U16702 ( .A(P2_ADDR_REG_16__SCAN_IN), .B(n14976), .Z(SUB_1596_U64)
         );
  OAI21_X1 U16703 ( .B1(n14978), .B2(P1_REG1_REG_0__SCAN_IN), .A(n14977), .ZN(
        n14980) );
  XNOR2_X1 U16704 ( .A(n14980), .B(n14979), .ZN(n14984) );
  AOI22_X1 U16705 ( .A1(n14981), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n14982) );
  OAI21_X1 U16706 ( .B1(n14984), .B2(n14983), .A(n14982), .ZN(P1_U3243) );
  AOI211_X1 U16707 ( .C1(n14987), .C2(n14986), .A(n14985), .B(n15060), .ZN(
        n14992) );
  AOI211_X1 U16708 ( .C1(n14990), .C2(n14989), .A(n14988), .B(n15056), .ZN(
        n14991) );
  AOI211_X1 U16709 ( .C1(n15067), .C2(n14993), .A(n14992), .B(n14991), .ZN(
        n14995) );
  OAI211_X1 U16710 ( .C1(n14996), .C2(n15070), .A(n14995), .B(n14994), .ZN(
        P1_U3256) );
  OAI21_X1 U16711 ( .B1(n14999), .B2(n14998), .A(n14997), .ZN(n15007) );
  INV_X1 U16712 ( .A(n15000), .ZN(n15001) );
  NOR2_X1 U16713 ( .A1(n15037), .A2(n15001), .ZN(n15006) );
  AOI211_X1 U16714 ( .C1(n15004), .C2(n15003), .A(n15002), .B(n15060), .ZN(
        n15005) );
  AOI211_X1 U16715 ( .C1(n15015), .C2(n15007), .A(n15006), .B(n15005), .ZN(
        n15009) );
  OAI211_X1 U16716 ( .C1(n15010), .C2(n15070), .A(n15009), .B(n15008), .ZN(
        P1_U3257) );
  XNOR2_X1 U16717 ( .A(n15011), .B(n8008), .ZN(n15013) );
  NAND2_X1 U16718 ( .A1(n15013), .A2(n15012), .ZN(n15018) );
  XNOR2_X1 U16719 ( .A(n15014), .B(n8007), .ZN(n15016) );
  NAND2_X1 U16720 ( .A1(n15016), .A2(n15015), .ZN(n15017) );
  OAI211_X1 U16721 ( .C1(n15037), .C2(n15019), .A(n15018), .B(n15017), .ZN(
        n15020) );
  INV_X1 U16722 ( .A(n15020), .ZN(n15022) );
  OAI211_X1 U16723 ( .C1(n15023), .C2(n15070), .A(n15022), .B(n15021), .ZN(
        P1_U3258) );
  NAND2_X1 U16724 ( .A1(n15025), .A2(n15024), .ZN(n15028) );
  NOR2_X1 U16725 ( .A1(n15056), .A2(n15026), .ZN(n15027) );
  NAND2_X1 U16726 ( .A1(n15028), .A2(n15027), .ZN(n15035) );
  NAND2_X1 U16727 ( .A1(n15030), .A2(n15029), .ZN(n15033) );
  NOR2_X1 U16728 ( .A1(n15060), .A2(n15031), .ZN(n15032) );
  NAND2_X1 U16729 ( .A1(n15033), .A2(n15032), .ZN(n15034) );
  OAI211_X1 U16730 ( .C1(n15037), .C2(n15036), .A(n15035), .B(n15034), .ZN(
        n15038) );
  INV_X1 U16731 ( .A(n15038), .ZN(n15040) );
  OAI211_X1 U16732 ( .C1(n15041), .C2(n15070), .A(n15040), .B(n15039), .ZN(
        P1_U3259) );
  INV_X1 U16733 ( .A(n15042), .ZN(n15046) );
  INV_X1 U16734 ( .A(n15043), .ZN(n15045) );
  AOI211_X1 U16735 ( .C1(n15046), .C2(n15045), .A(n15044), .B(n15056), .ZN(
        n15051) );
  AOI211_X1 U16736 ( .C1(n15049), .C2(n15048), .A(n15047), .B(n15060), .ZN(
        n15050) );
  AOI211_X1 U16737 ( .C1(n15067), .C2(n15052), .A(n15051), .B(n15050), .ZN(
        n15054) );
  OAI211_X1 U16738 ( .C1(n15055), .C2(n15070), .A(n15054), .B(n15053), .ZN(
        P1_U3260) );
  INV_X1 U16739 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n15071) );
  AOI211_X1 U16740 ( .C1(n15059), .C2(n15058), .A(n15057), .B(n15056), .ZN(
        n15065) );
  AOI211_X1 U16741 ( .C1(n15063), .C2(n15062), .A(n15061), .B(n15060), .ZN(
        n15064) );
  AOI211_X1 U16742 ( .C1(n15067), .C2(n15066), .A(n15065), .B(n15064), .ZN(
        n15069) );
  OAI211_X1 U16743 ( .C1(n15071), .C2(n15070), .A(n15069), .B(n15068), .ZN(
        P1_U3261) );
  XNOR2_X1 U16744 ( .A(n15072), .B(n15073), .ZN(n15136) );
  XNOR2_X1 U16745 ( .A(n15074), .B(n15073), .ZN(n15076) );
  NOR2_X1 U16746 ( .A1(n15076), .A2(n15075), .ZN(n15077) );
  AOI211_X1 U16747 ( .C1(n15162), .C2(n15136), .A(n15078), .B(n15077), .ZN(
        n15133) );
  INV_X1 U16748 ( .A(n15079), .ZN(n15080) );
  AOI222_X1 U16749 ( .A1(n15083), .A2(n15081), .B1(P1_REG2_REG_6__SCAN_IN), 
        .B2(n15105), .C1(n15102), .C2(n15080), .ZN(n15093) );
  INV_X1 U16750 ( .A(n15082), .ZN(n15091) );
  INV_X1 U16751 ( .A(n15083), .ZN(n15132) );
  INV_X1 U16752 ( .A(n15084), .ZN(n15088) );
  INV_X1 U16753 ( .A(n15085), .ZN(n15087) );
  OAI211_X1 U16754 ( .C1(n15132), .C2(n15088), .A(n15087), .B(n15086), .ZN(
        n15131) );
  INV_X1 U16755 ( .A(n15131), .ZN(n15089) );
  AOI22_X1 U16756 ( .A1(n15136), .A2(n15091), .B1(n15090), .B2(n15089), .ZN(
        n15092) );
  OAI211_X1 U16757 ( .C1(n15105), .C2(n15133), .A(n15093), .B(n15092), .ZN(
        P1_U3287) );
  INV_X1 U16758 ( .A(n15094), .ZN(n15096) );
  AOI21_X1 U16759 ( .B1(n15097), .B2(n15096), .A(n15095), .ZN(n15104) );
  AOI21_X1 U16760 ( .B1(n15100), .B2(n15099), .A(n15098), .ZN(n15101) );
  AOI21_X1 U16761 ( .B1(n15102), .B2(P1_REG3_REG_0__SCAN_IN), .A(n15101), .ZN(
        n15103) );
  OAI221_X1 U16762 ( .B1(n15105), .B2(n15104), .C1(n14539), .C2(n7731), .A(
        n15103), .ZN(P1_U3293) );
  AND2_X1 U16763 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n15109), .ZN(P1_U3294) );
  AND2_X1 U16764 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n15109), .ZN(P1_U3295) );
  INV_X1 U16765 ( .A(n15109), .ZN(n15108) );
  NOR2_X1 U16766 ( .A1(n15108), .A2(n15106), .ZN(P1_U3296) );
  AND2_X1 U16767 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n15109), .ZN(P1_U3297) );
  AND2_X1 U16768 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n15109), .ZN(P1_U3298) );
  AND2_X1 U16769 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n15109), .ZN(P1_U3299) );
  AND2_X1 U16770 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n15109), .ZN(P1_U3300) );
  AND2_X1 U16771 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n15109), .ZN(P1_U3301) );
  AND2_X1 U16772 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n15109), .ZN(P1_U3302) );
  AND2_X1 U16773 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n15109), .ZN(P1_U3303) );
  AND2_X1 U16774 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n15109), .ZN(P1_U3304) );
  AND2_X1 U16775 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n15109), .ZN(P1_U3305) );
  AND2_X1 U16776 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n15109), .ZN(P1_U3306) );
  AND2_X1 U16777 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n15109), .ZN(P1_U3307) );
  AND2_X1 U16778 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n15109), .ZN(P1_U3308) );
  AND2_X1 U16779 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n15109), .ZN(P1_U3309) );
  AND2_X1 U16780 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n15109), .ZN(P1_U3310) );
  AND2_X1 U16781 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n15109), .ZN(P1_U3311) );
  AND2_X1 U16782 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n15109), .ZN(P1_U3312) );
  AND2_X1 U16783 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n15109), .ZN(P1_U3313) );
  AND2_X1 U16784 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n15109), .ZN(P1_U3314) );
  AND2_X1 U16785 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n15109), .ZN(P1_U3315) );
  AND2_X1 U16786 ( .A1(n15109), .A2(P1_D_REG_9__SCAN_IN), .ZN(P1_U3316) );
  NOR2_X1 U16787 ( .A1(n15108), .A2(n15107), .ZN(P1_U3317) );
  AND2_X1 U16788 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n15109), .ZN(P1_U3318) );
  AND2_X1 U16789 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n15109), .ZN(P1_U3319) );
  AND2_X1 U16790 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n15109), .ZN(P1_U3320) );
  AND2_X1 U16791 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n15109), .ZN(P1_U3321) );
  AND2_X1 U16792 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n15109), .ZN(P1_U3322) );
  AND2_X1 U16793 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n15109), .ZN(P1_U3323) );
  OAI21_X1 U16794 ( .B1(n15111), .B2(n15166), .A(n15110), .ZN(n15112) );
  AOI21_X1 U16795 ( .B1(n15113), .B2(n15137), .A(n15112), .ZN(n15114) );
  AND2_X1 U16796 ( .A1(n15115), .A2(n15114), .ZN(n15176) );
  AOI22_X1 U16797 ( .A1(n15174), .A2(n15176), .B1(n7741), .B2(n15172), .ZN(
        P1_U3465) );
  OAI21_X1 U16798 ( .B1(n15117), .B2(n15166), .A(n15116), .ZN(n15119) );
  AOI211_X1 U16799 ( .C1(n15120), .C2(n15170), .A(n15119), .B(n15118), .ZN(
        n15177) );
  INV_X1 U16800 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n15121) );
  AOI22_X1 U16801 ( .A1(n15174), .A2(n15177), .B1(n15121), .B2(n15172), .ZN(
        P1_U3471) );
  INV_X1 U16802 ( .A(n15126), .ZN(n15128) );
  OAI21_X1 U16803 ( .B1(n15123), .B2(n15166), .A(n15122), .ZN(n15125) );
  AOI211_X1 U16804 ( .C1(n15137), .C2(n15126), .A(n15125), .B(n15124), .ZN(
        n15127) );
  OAI21_X1 U16805 ( .B1(n15129), .B2(n15128), .A(n15127), .ZN(n15130) );
  INV_X1 U16806 ( .A(n15130), .ZN(n15178) );
  AOI22_X1 U16807 ( .A1(n15174), .A2(n15178), .B1(n7814), .B2(n15172), .ZN(
        P1_U3474) );
  OAI21_X1 U16808 ( .B1(n15132), .B2(n15166), .A(n15131), .ZN(n15135) );
  INV_X1 U16809 ( .A(n15133), .ZN(n15134) );
  AOI211_X1 U16810 ( .C1(n15137), .C2(n15136), .A(n15135), .B(n15134), .ZN(
        n15179) );
  INV_X1 U16811 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n15138) );
  AOI22_X1 U16812 ( .A1(n15174), .A2(n15179), .B1(n15138), .B2(n15172), .ZN(
        P1_U3477) );
  INV_X1 U16813 ( .A(n15143), .ZN(n15145) );
  AOI211_X1 U16814 ( .C1(n15141), .C2(n15155), .A(n15140), .B(n15139), .ZN(
        n15142) );
  OAI21_X1 U16815 ( .B1(n15159), .B2(n15143), .A(n15142), .ZN(n15144) );
  AOI21_X1 U16816 ( .B1(n15162), .B2(n15145), .A(n15144), .ZN(n15180) );
  INV_X1 U16817 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n15146) );
  AOI22_X1 U16818 ( .A1(n15174), .A2(n15180), .B1(n15146), .B2(n15172), .ZN(
        P1_U3480) );
  OAI211_X1 U16819 ( .C1(n6920), .C2(n15166), .A(n15148), .B(n15147), .ZN(
        n15150) );
  AOI211_X1 U16820 ( .C1(n15151), .C2(n15170), .A(n15150), .B(n15149), .ZN(
        n15181) );
  INV_X1 U16821 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n15152) );
  AOI22_X1 U16822 ( .A1(n15174), .A2(n15181), .B1(n15152), .B2(n15172), .ZN(
        P1_U3483) );
  AOI211_X1 U16823 ( .C1(n15156), .C2(n15155), .A(n15154), .B(n15153), .ZN(
        n15157) );
  OAI21_X1 U16824 ( .B1(n15159), .B2(n15158), .A(n15157), .ZN(n15160) );
  AOI21_X1 U16825 ( .B1(n15162), .B2(n15161), .A(n15160), .ZN(n15182) );
  INV_X1 U16826 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n15163) );
  AOI22_X1 U16827 ( .A1(n15174), .A2(n15182), .B1(n15163), .B2(n15172), .ZN(
        P1_U3486) );
  OAI211_X1 U16828 ( .C1(n15167), .C2(n15166), .A(n15165), .B(n15164), .ZN(
        n15169) );
  AOI211_X1 U16829 ( .C1(n15171), .C2(n15170), .A(n15169), .B(n15168), .ZN(
        n15184) );
  INV_X1 U16830 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n15173) );
  AOI22_X1 U16831 ( .A1(n15174), .A2(n15184), .B1(n15173), .B2(n15172), .ZN(
        P1_U3489) );
  AOI22_X1 U16832 ( .A1(n15185), .A2(n15176), .B1(n15175), .B2(n15183), .ZN(
        P1_U3530) );
  AOI22_X1 U16833 ( .A1(n15185), .A2(n15177), .B1(n9916), .B2(n15183), .ZN(
        P1_U3532) );
  AOI22_X1 U16834 ( .A1(n15185), .A2(n15178), .B1(n9918), .B2(n15183), .ZN(
        P1_U3533) );
  AOI22_X1 U16835 ( .A1(n15185), .A2(n15179), .B1(n9913), .B2(n15183), .ZN(
        P1_U3534) );
  AOI22_X1 U16836 ( .A1(n15185), .A2(n15180), .B1(n10377), .B2(n15183), .ZN(
        P1_U3535) );
  AOI22_X1 U16837 ( .A1(n15185), .A2(n15181), .B1(n10991), .B2(n15183), .ZN(
        P1_U3536) );
  AOI22_X1 U16838 ( .A1(n15185), .A2(n15182), .B1(n10992), .B2(n15183), .ZN(
        P1_U3537) );
  AOI22_X1 U16839 ( .A1(n15185), .A2(n15184), .B1(n10987), .B2(n15183), .ZN(
        P1_U3538) );
  NOR2_X1 U16840 ( .A1(n15313), .A2(n6623), .ZN(P2_U3087) );
  NAND2_X1 U16841 ( .A1(n15188), .A2(n15187), .ZN(n15189) );
  XNOR2_X1 U16842 ( .A(n15186), .B(n15189), .ZN(n15192) );
  AOI222_X1 U16843 ( .A1(n15195), .A2(n15194), .B1(n15193), .B2(n15192), .C1(
        n15191), .C2(n15190), .ZN(n15196) );
  NAND2_X1 U16844 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3088), .ZN(n15286)
         );
  OAI211_X1 U16845 ( .C1(n15198), .C2(n15197), .A(n15196), .B(n15286), .ZN(
        P2_U3196) );
  AOI22_X1 U16846 ( .A1(P2_REG2_REG_0__SCAN_IN), .A2(n15314), .B1(n15307), 
        .B2(P2_REG1_REG_0__SCAN_IN), .ZN(n15202) );
  OAI22_X1 U16847 ( .A1(P2_REG1_REG_0__SCAN_IN), .A2(n15292), .B1(n15298), 
        .B2(P2_REG2_REG_0__SCAN_IN), .ZN(n15199) );
  NOR2_X1 U16848 ( .A1(n15318), .A2(n15199), .ZN(n15201) );
  AOI22_X1 U16849 ( .A1(n15313), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3088), .ZN(n15200) );
  OAI221_X1 U16850 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(n15202), .C1(n8396), .C2(
        n15201), .A(n15200), .ZN(P2_U3214) );
  INV_X1 U16851 ( .A(n15203), .ZN(n15205) );
  NAND2_X1 U16852 ( .A1(n15205), .A2(n15204), .ZN(n15206) );
  NAND3_X1 U16853 ( .A1(n15307), .A2(n15207), .A3(n15206), .ZN(n15210) );
  NAND2_X1 U16854 ( .A1(n15318), .A2(n15208), .ZN(n15209) );
  OAI211_X1 U16855 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n15211), .A(n15210), .B(
        n15209), .ZN(n15212) );
  INV_X1 U16856 ( .A(n15212), .ZN(n15217) );
  AND2_X1 U16857 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n15215) );
  OAI211_X1 U16858 ( .C1(n15215), .C2(n15214), .A(n15314), .B(n15213), .ZN(
        n15216) );
  OAI211_X1 U16859 ( .C1(n15306), .C2(n15218), .A(n15217), .B(n15216), .ZN(
        P2_U3215) );
  AOI22_X1 U16860 ( .A1(n15313), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3088), .ZN(n15231) );
  OAI211_X1 U16861 ( .C1(n15221), .C2(n15220), .A(n15307), .B(n15219), .ZN(
        n15222) );
  OAI21_X1 U16862 ( .B1(n15224), .B2(n15223), .A(n15222), .ZN(n15225) );
  INV_X1 U16863 ( .A(n15225), .ZN(n15230) );
  OAI211_X1 U16864 ( .C1(n15228), .C2(n15227), .A(n15314), .B(n15226), .ZN(
        n15229) );
  NAND3_X1 U16865 ( .A1(n15231), .A2(n15230), .A3(n15229), .ZN(P2_U3216) );
  INV_X1 U16866 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n15514) );
  OAI211_X1 U16867 ( .C1(n15234), .C2(n15233), .A(n15307), .B(n15232), .ZN(
        n15239) );
  NAND3_X1 U16868 ( .A1(n15236), .A2(n15235), .A3(n8867), .ZN(n15237) );
  AND3_X1 U16869 ( .A1(n15239), .A2(n15238), .A3(n15237), .ZN(n15244) );
  OAI211_X1 U16870 ( .C1(n15242), .C2(n15241), .A(n15314), .B(n15240), .ZN(
        n15243) );
  OAI211_X1 U16871 ( .C1(n15306), .C2(n15514), .A(n15244), .B(n15243), .ZN(
        P2_U3217) );
  OAI21_X1 U16872 ( .B1(n15247), .B2(n15246), .A(n15245), .ZN(n15254) );
  NAND2_X1 U16873 ( .A1(n15249), .A2(n15248), .ZN(n15250) );
  NAND2_X1 U16874 ( .A1(n15251), .A2(n15250), .ZN(n15252) );
  AOI222_X1 U16875 ( .A1(n15254), .A2(n15314), .B1(n15253), .B2(n15318), .C1(
        n15252), .C2(n15307), .ZN(n15256) );
  OAI211_X1 U16876 ( .C1(n7052), .C2(n15306), .A(n15256), .B(n15255), .ZN(
        P2_U3223) );
  INV_X1 U16877 ( .A(n15257), .ZN(n15263) );
  INV_X1 U16878 ( .A(n15258), .ZN(n15259) );
  AOI211_X1 U16879 ( .C1(n15261), .C2(n15260), .A(n15292), .B(n15259), .ZN(
        n15262) );
  AOI211_X1 U16880 ( .C1(n15318), .C2(n15264), .A(n15263), .B(n15262), .ZN(
        n15270) );
  AOI211_X1 U16881 ( .C1(n15267), .C2(n15266), .A(n15298), .B(n15265), .ZN(
        n15268) );
  INV_X1 U16882 ( .A(n15268), .ZN(n15269) );
  OAI211_X1 U16883 ( .C1(n15306), .C2(n15271), .A(n15270), .B(n15269), .ZN(
        P2_U3224) );
  NAND2_X1 U16884 ( .A1(n15273), .A2(n15272), .ZN(n15274) );
  AOI21_X1 U16885 ( .B1(n15275), .B2(n15274), .A(n15292), .ZN(n15284) );
  INV_X1 U16886 ( .A(n15276), .ZN(n15279) );
  INV_X1 U16887 ( .A(n15277), .ZN(n15278) );
  NAND3_X1 U16888 ( .A1(n15280), .A2(n15279), .A3(n15278), .ZN(n15281) );
  AOI21_X1 U16889 ( .B1(n15282), .B2(n15281), .A(n15298), .ZN(n15283) );
  AOI211_X1 U16890 ( .C1(n15318), .C2(n15285), .A(n15284), .B(n15283), .ZN(
        n15287) );
  OAI211_X1 U16891 ( .C1(n15288), .C2(n15306), .A(n15287), .B(n15286), .ZN(
        P2_U3226) );
  NOR2_X1 U16892 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n15289), .ZN(n15296) );
  INV_X1 U16893 ( .A(n15290), .ZN(n15291) );
  AOI211_X1 U16894 ( .C1(n15294), .C2(n15293), .A(n15292), .B(n15291), .ZN(
        n15295) );
  AOI211_X1 U16895 ( .C1(n15318), .C2(n15297), .A(n15296), .B(n15295), .ZN(
        n15304) );
  AOI21_X1 U16896 ( .B1(n15300), .B2(n15299), .A(n15298), .ZN(n15302) );
  NAND2_X1 U16897 ( .A1(n15302), .A2(n15301), .ZN(n15303) );
  OAI211_X1 U16898 ( .C1(n15306), .C2(n15305), .A(n15304), .B(n15303), .ZN(
        P2_U3227) );
  OAI21_X1 U16899 ( .B1(n15309), .B2(n15308), .A(n15307), .ZN(n15311) );
  NOR2_X1 U16900 ( .A1(n15311), .A2(n15310), .ZN(n15312) );
  AOI21_X1 U16901 ( .B1(n15313), .B2(P2_ADDR_REG_14__SCAN_IN), .A(n15312), 
        .ZN(n15322) );
  OAI211_X1 U16902 ( .C1(n15316), .C2(P2_REG2_REG_14__SCAN_IN), .A(n15315), 
        .B(n15314), .ZN(n15320) );
  NAND2_X1 U16903 ( .A1(n15318), .A2(n15317), .ZN(n15319) );
  NAND4_X1 U16904 ( .A1(n15322), .A2(n15321), .A3(n15320), .A4(n15319), .ZN(
        P2_U3228) );
  INV_X1 U16905 ( .A(n15323), .ZN(n15331) );
  NAND2_X1 U16906 ( .A1(n15325), .A2(n15324), .ZN(n15329) );
  AOI22_X1 U16907 ( .A1(n6620), .A2(P2_REG2_REG_7__SCAN_IN), .B1(n15327), .B2(
        n15326), .ZN(n15328) );
  OAI211_X1 U16908 ( .C1(n15331), .C2(n15330), .A(n15329), .B(n15328), .ZN(
        n15332) );
  AOI21_X1 U16909 ( .B1(n15334), .B2(n15333), .A(n15332), .ZN(n15335) );
  OAI21_X1 U16910 ( .B1(n6620), .B2(n15336), .A(n15335), .ZN(P2_U3258) );
  AND2_X1 U16911 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n15343), .ZN(P2_U3266) );
  AND2_X1 U16912 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n15343), .ZN(P2_U3267) );
  AND2_X1 U16913 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n15343), .ZN(P2_U3268) );
  NOR2_X1 U16914 ( .A1(n15342), .A2(n15338), .ZN(P2_U3269) );
  AND2_X1 U16915 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n15343), .ZN(P2_U3270) );
  AND2_X1 U16916 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n15343), .ZN(P2_U3271) );
  NOR2_X1 U16917 ( .A1(n15342), .A2(n15339), .ZN(P2_U3272) );
  AND2_X1 U16918 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n15343), .ZN(P2_U3273) );
  NOR2_X1 U16919 ( .A1(n15342), .A2(n15340), .ZN(P2_U3274) );
  AND2_X1 U16920 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n15343), .ZN(P2_U3275) );
  AND2_X1 U16921 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n15343), .ZN(P2_U3276) );
  AND2_X1 U16922 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n15343), .ZN(P2_U3277) );
  AND2_X1 U16923 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n15343), .ZN(P2_U3278) );
  AND2_X1 U16924 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n15343), .ZN(P2_U3279) );
  AND2_X1 U16925 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n15343), .ZN(P2_U3280) );
  AND2_X1 U16926 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n15343), .ZN(P2_U3281) );
  AND2_X1 U16927 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n15343), .ZN(P2_U3282) );
  NOR2_X1 U16928 ( .A1(n15342), .A2(n15341), .ZN(P2_U3283) );
  AND2_X1 U16929 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n15343), .ZN(P2_U3284) );
  AND2_X1 U16930 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n15343), .ZN(P2_U3285) );
  AND2_X1 U16931 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n15343), .ZN(P2_U3286) );
  AND2_X1 U16932 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n15343), .ZN(P2_U3287) );
  AND2_X1 U16933 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n15343), .ZN(P2_U3288) );
  AND2_X1 U16934 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n15343), .ZN(P2_U3289) );
  AND2_X1 U16935 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n15343), .ZN(P2_U3290) );
  AND2_X1 U16936 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n15343), .ZN(P2_U3291) );
  AND2_X1 U16937 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n15343), .ZN(P2_U3292) );
  AND2_X1 U16938 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n15343), .ZN(P2_U3293) );
  AND2_X1 U16939 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n15343), .ZN(P2_U3294) );
  AND2_X1 U16940 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n15343), .ZN(P2_U3295) );
  AOI22_X1 U16941 ( .A1(n15349), .A2(n15345), .B1(n15344), .B2(n15346), .ZN(
        P2_U3416) );
  AOI22_X1 U16942 ( .A1(n15349), .A2(n15348), .B1(n15347), .B2(n15346), .ZN(
        P2_U3417) );
  INV_X1 U16943 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n15350) );
  AOI22_X1 U16944 ( .A1(n15383), .A2(n15351), .B1(n15350), .B2(n15382), .ZN(
        P2_U3430) );
  INV_X1 U16945 ( .A(n15352), .ZN(n15359) );
  INV_X1 U16946 ( .A(n15360), .ZN(n15357) );
  AOI21_X1 U16947 ( .B1(n15355), .B2(n15354), .A(n15353), .ZN(n15356) );
  OAI21_X1 U16948 ( .B1(n15357), .B2(n15362), .A(n15356), .ZN(n15358) );
  AOI211_X1 U16949 ( .C1(n15361), .C2(n15360), .A(n15359), .B(n15358), .ZN(
        n15385) );
  AOI22_X1 U16950 ( .A1(n15383), .A2(n15385), .B1(n8398), .B2(n15382), .ZN(
        P2_U3436) );
  NOR2_X1 U16951 ( .A1(n15363), .A2(n15362), .ZN(n15368) );
  INV_X1 U16952 ( .A(n15364), .ZN(n15366) );
  OAI21_X1 U16953 ( .B1(n15366), .B2(n15378), .A(n15365), .ZN(n15367) );
  NOR3_X1 U16954 ( .A1(n15369), .A2(n15368), .A3(n15367), .ZN(n15387) );
  AOI22_X1 U16955 ( .A1(n15383), .A2(n15387), .B1(n8487), .B2(n15382), .ZN(
        P2_U3454) );
  OAI21_X1 U16956 ( .B1(n7268), .B2(n15378), .A(n15371), .ZN(n15372) );
  AOI21_X1 U16957 ( .B1(n15373), .B2(n8890), .A(n15372), .ZN(n15374) );
  AND2_X1 U16958 ( .A1(n15375), .A2(n15374), .ZN(n15388) );
  AOI22_X1 U16959 ( .A1(n15383), .A2(n15388), .B1(n8513), .B2(n15382), .ZN(
        P2_U3460) );
  OAI211_X1 U16960 ( .C1(n6889), .C2(n15378), .A(n15377), .B(n15376), .ZN(
        n15379) );
  AOI21_X1 U16961 ( .B1(n15381), .B2(n15380), .A(n15379), .ZN(n15391) );
  AOI22_X1 U16962 ( .A1(n15383), .A2(n15391), .B1(n8525), .B2(n15382), .ZN(
        P2_U3463) );
  AOI22_X1 U16963 ( .A1(n15392), .A2(n15385), .B1(n15384), .B2(n15389), .ZN(
        P2_U3501) );
  AOI22_X1 U16964 ( .A1(n15392), .A2(n15387), .B1(n15386), .B2(n15389), .ZN(
        P2_U3507) );
  AOI22_X1 U16965 ( .A1(n15392), .A2(n15388), .B1(n10482), .B2(n15389), .ZN(
        P2_U3509) );
  AOI22_X1 U16966 ( .A1(n15392), .A2(n15391), .B1(n15390), .B2(n15389), .ZN(
        P2_U3510) );
  NOR2_X1 U16967 ( .A1(P3_U3897), .A2(n15415), .ZN(P3_U3150) );
  AOI21_X1 U16968 ( .B1(n15395), .B2(n15394), .A(n15393), .ZN(n15402) );
  OAI21_X1 U16969 ( .B1(n15398), .B2(n15397), .A(n15396), .ZN(n15399) );
  NAND2_X1 U16970 ( .A1(n15426), .A2(n15399), .ZN(n15400) );
  OAI21_X1 U16971 ( .B1(n15402), .B2(n15401), .A(n15400), .ZN(n15409) );
  AOI21_X1 U16972 ( .B1(n15405), .B2(n15404), .A(n15403), .ZN(n15407) );
  NOR2_X1 U16973 ( .A1(n15407), .A2(n15406), .ZN(n15408) );
  AOI211_X1 U16974 ( .C1(n15417), .C2(n15410), .A(n15409), .B(n15408), .ZN(
        n15412) );
  OAI211_X1 U16975 ( .C1(n15414), .C2(n15413), .A(n15412), .B(n15411), .ZN(
        P3_U3186) );
  AOI22_X1 U16976 ( .A1(n15417), .A2(n15416), .B1(n15415), .B2(
        P3_ADDR_REG_10__SCAN_IN), .ZN(n15434) );
  XNOR2_X1 U16977 ( .A(n15419), .B(n15418), .ZN(n15431) );
  OAI21_X1 U16978 ( .B1(n15422), .B2(n15421), .A(n15420), .ZN(n15428) );
  OAI21_X1 U16979 ( .B1(n15425), .B2(n15424), .A(n15423), .ZN(n15427) );
  AOI222_X1 U16980 ( .A1(n15431), .A2(n15430), .B1(n15429), .B2(n15428), .C1(
        n15427), .C2(n15426), .ZN(n15433) );
  NAND3_X1 U16981 ( .A1(n15434), .A2(n15433), .A3(n15432), .ZN(P3_U3192) );
  AOI21_X1 U16982 ( .B1(n15437), .B2(n15436), .A(n15435), .ZN(n15438) );
  OAI222_X1 U16983 ( .A1(n15442), .A2(n15441), .B1(n15440), .B2(n15439), .C1(
        n13024), .C2(n15438), .ZN(n15443) );
  INV_X1 U16984 ( .A(n15443), .ZN(n15444) );
  OAI21_X1 U16985 ( .B1(n15464), .B2(n15445), .A(n15444), .ZN(P3_U3227) );
  XNOR2_X1 U16986 ( .A(n15446), .B(n15448), .ZN(n15456) );
  OAI21_X1 U16987 ( .B1(n15449), .B2(n15448), .A(n15447), .ZN(n15474) );
  OAI22_X1 U16988 ( .A1(n10678), .A2(n15452), .B1(n15451), .B2(n15450), .ZN(
        n15453) );
  AOI21_X1 U16989 ( .B1(n15474), .B2(n15454), .A(n15453), .ZN(n15455) );
  OAI21_X1 U16990 ( .B1(n15457), .B2(n15456), .A(n15455), .ZN(n15472) );
  NOR2_X1 U16991 ( .A1(n15458), .A2(n15486), .ZN(n15473) );
  AOI22_X1 U16992 ( .A1(n15474), .A2(n15460), .B1(n15473), .B2(n15459), .ZN(
        n15461) );
  INV_X1 U16993 ( .A(n15461), .ZN(n15462) );
  AOI211_X1 U16994 ( .C1(n15463), .C2(P3_REG3_REG_2__SCAN_IN), .A(n15472), .B(
        n15462), .ZN(n15465) );
  AOI22_X1 U16995 ( .A1(n13024), .A2(n10532), .B1(n15465), .B2(n15464), .ZN(
        P3_U3231) );
  INV_X1 U16996 ( .A(n15467), .ZN(n15469) );
  AOI211_X1 U16997 ( .C1(n15475), .C2(n15470), .A(n15469), .B(n15468), .ZN(
        n15494) );
  INV_X1 U16998 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n15471) );
  AOI22_X1 U16999 ( .A1(n15493), .A2(n15494), .B1(n15471), .B2(n15491), .ZN(
        P3_U3393) );
  AOI211_X1 U17000 ( .C1(n15475), .C2(n15474), .A(n15473), .B(n15472), .ZN(
        n15495) );
  INV_X1 U17001 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n15476) );
  AOI22_X1 U17002 ( .A1(n15493), .A2(n15495), .B1(n15476), .B2(n15491), .ZN(
        P3_U3396) );
  AND2_X1 U17003 ( .A1(n15478), .A2(n15477), .ZN(n15482) );
  AND2_X1 U17004 ( .A1(n15480), .A2(n15479), .ZN(n15481) );
  NOR3_X1 U17005 ( .A1(n15483), .A2(n15482), .A3(n15481), .ZN(n15496) );
  INV_X1 U17006 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n15484) );
  AOI22_X1 U17007 ( .A1(n15493), .A2(n15496), .B1(n15484), .B2(n15491), .ZN(
        P3_U3402) );
  OAI22_X1 U17008 ( .A1(n15488), .A2(n15487), .B1(n15486), .B2(n15485), .ZN(
        n15489) );
  NOR2_X1 U17009 ( .A1(n15490), .A2(n15489), .ZN(n15497) );
  INV_X1 U17010 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n15492) );
  AOI22_X1 U17011 ( .A1(n15493), .A2(n15497), .B1(n15492), .B2(n15491), .ZN(
        P3_U3417) );
  AOI22_X1 U17012 ( .A1(n15498), .A2(n15494), .B1(n10509), .B2(n6791), .ZN(
        P3_U3460) );
  AOI22_X1 U17013 ( .A1(n15498), .A2(n15495), .B1(n10516), .B2(n6791), .ZN(
        P3_U3461) );
  AOI22_X1 U17014 ( .A1(n15498), .A2(n15496), .B1(n10800), .B2(n6791), .ZN(
        P3_U3463) );
  AOI22_X1 U17015 ( .A1(n15498), .A2(n15497), .B1(n9198), .B2(n6791), .ZN(
        P3_U3468) );
  AOI21_X1 U17016 ( .B1(n15501), .B2(n15500), .A(n15499), .ZN(SUB_1596_U53) );
  AOI21_X1 U17017 ( .B1(n15504), .B2(n15503), .A(n15502), .ZN(SUB_1596_U59) );
  OAI21_X1 U17018 ( .B1(n15507), .B2(n15506), .A(n15505), .ZN(SUB_1596_U58) );
  AOI21_X1 U17019 ( .B1(n15510), .B2(n15509), .A(n15508), .ZN(SUB_1596_U56) );
  AOI21_X1 U17020 ( .B1(n15513), .B2(n15512), .A(n15511), .ZN(n15515) );
  XNOR2_X1 U17021 ( .A(n15515), .B(n15514), .ZN(SUB_1596_U60) );
  AOI21_X1 U17022 ( .B1(n15518), .B2(n15517), .A(n15516), .ZN(SUB_1596_U5) );
  INV_X1 U7375 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n8803) );
  OR2_X1 U9498 ( .A1(n9584), .A2(n7195), .ZN(n7192) );
  CLKBUF_X2 U7368 ( .A(n12208), .Z(n12288) );
  CLKBUF_X1 U7381 ( .A(n12360), .Z(n6818) );
  CLKBUF_X1 U7616 ( .A(n9250), .Z(n10506) );
  CLKBUF_X1 U8354 ( .A(n13857), .Z(n6827) );
  XNOR2_X1 U8749 ( .A(n12659), .B(n7189), .ZN(n13153) );
  CLKBUF_X1 U8815 ( .A(n13324), .Z(n6830) );
  CLKBUF_X3 U9303 ( .A(n8415), .Z(n9090) );
  INV_X2 U9497 ( .A(n15105), .ZN(n14539) );
endmodule

