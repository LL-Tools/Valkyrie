

module b20_C_2inp_gates_syn ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, ADD_1068_U4, 
        ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58, ADD_1068_U59, 
        ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63, ADD_1068_U47, 
        ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51, ADD_1068_U52, 
        ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46, U126, U123, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439, P1_U3440, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462, P1_U3465, P1_U3468, 
        P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, 
        P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3509, 
        P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, 
        P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, 
        P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, 
        P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, 
        P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, 
        P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, 
        P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3554, P1_U3555, 
        P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, 
        P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, 
        P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, 
        P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, 
        P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U3973, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376, P2_U3377, P2_U3263, 
        P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, 
        P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, 
        P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, 
        P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, 
        P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399, P2_U3402, P2_U3405, 
        P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420, P2_U3423, P2_U3426, 
        P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441, P2_U3444, P2_U3446, 
        P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451, P2_U3452, P2_U3453, 
        P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458, P2_U3459, P2_U3460, 
        P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465, P2_U3466, P2_U3467, 
        P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472, P2_U3473, P2_U3474, 
        P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479, P2_U3480, P2_U3481, 
        P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486, P2_U3487, P2_U3488, 
        P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, 
        P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, 
        P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, 
        P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3491, P2_U3492, 
        P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, 
        P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, 
        P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, 
        P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, 
        P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180, P2_U3179, P2_U3178, 
        P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, P2_U3171, 
        P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, P2_U3164, 
        P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, P2_U3157, 
        P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151, P2_U3150, P2_U3893, 
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, 
        keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, 
        keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, 
        keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, 
        keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, 
        keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, 
        keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, 
        keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, 
        keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, 
        keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, 
        keyinput60, keyinput61, keyinput62, keyinput63 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278,
         n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288,
         n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298,
         n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308,
         n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318,
         n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328,
         n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338,
         n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348,
         n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358,
         n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368,
         n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378,
         n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388,
         n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398,
         n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408,
         n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418,
         n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428,
         n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438,
         n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448,
         n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458,
         n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468,
         n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478,
         n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488,
         n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498,
         n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508,
         n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518,
         n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528,
         n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538,
         n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548,
         n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558,
         n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568,
         n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578,
         n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588,
         n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598,
         n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608,
         n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618,
         n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628,
         n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638,
         n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648,
         n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658,
         n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668,
         n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678,
         n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688,
         n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698,
         n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708,
         n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718,
         n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728,
         n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738,
         n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748,
         n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758,
         n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768,
         n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778,
         n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788,
         n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798,
         n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808,
         n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818,
         n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828,
         n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838,
         n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848,
         n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858,
         n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868,
         n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878,
         n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888,
         n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898,
         n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908,
         n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918,
         n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928,
         n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938,
         n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948,
         n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958,
         n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968,
         n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978,
         n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988,
         n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998,
         n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008,
         n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018,
         n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028,
         n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038,
         n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048,
         n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058,
         n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068,
         n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078,
         n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088,
         n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098,
         n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108,
         n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118,
         n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128,
         n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138,
         n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148,
         n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158,
         n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168,
         n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178,
         n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188,
         n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198,
         n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208,
         n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218,
         n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228,
         n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238,
         n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248,
         n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258,
         n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268,
         n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278,
         n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288,
         n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298,
         n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308,
         n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318,
         n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328,
         n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338,
         n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348,
         n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358,
         n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368,
         n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378,
         n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388,
         n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398,
         n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408,
         n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418,
         n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428,
         n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438,
         n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448,
         n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458,
         n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468,
         n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478,
         n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488,
         n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498,
         n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508,
         n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518,
         n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528,
         n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538,
         n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548,
         n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558,
         n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568,
         n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578,
         n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588,
         n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598,
         n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608,
         n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618,
         n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628,
         n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638,
         n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648,
         n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658,
         n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668,
         n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678,
         n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688,
         n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698,
         n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708,
         n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718,
         n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728,
         n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738,
         n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748,
         n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758,
         n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768,
         n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778,
         n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788,
         n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798,
         n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808,
         n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818,
         n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828,
         n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838,
         n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848,
         n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858,
         n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868,
         n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878,
         n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888,
         n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898,
         n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908,
         n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918,
         n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928,
         n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938,
         n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948,
         n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958,
         n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968,
         n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978,
         n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988,
         n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998,
         n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008,
         n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018,
         n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028,
         n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038,
         n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048,
         n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058,
         n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068,
         n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078,
         n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088,
         n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098,
         n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108,
         n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118,
         n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128,
         n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138,
         n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148,
         n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158,
         n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168,
         n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178,
         n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188,
         n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198,
         n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208,
         n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218,
         n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228,
         n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238,
         n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248,
         n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258,
         n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268,
         n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278,
         n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288,
         n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298,
         n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308,
         n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318,
         n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328,
         n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338,
         n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348,
         n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358,
         n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368,
         n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378,
         n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388,
         n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398,
         n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408,
         n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418,
         n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428,
         n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438,
         n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448,
         n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458,
         n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468,
         n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478,
         n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488,
         n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498,
         n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508,
         n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518,
         n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528,
         n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538,
         n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548,
         n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558,
         n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568,
         n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578,
         n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588,
         n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598,
         n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608,
         n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618,
         n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628,
         n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638,
         n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648,
         n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658,
         n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668,
         n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678,
         n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688,
         n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698,
         n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708,
         n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718,
         n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728,
         n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738,
         n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748,
         n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758,
         n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768,
         n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778,
         n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788,
         n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798,
         n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808,
         n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818,
         n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828,
         n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838,
         n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848,
         n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858,
         n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868,
         n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878,
         n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888,
         n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898,
         n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908,
         n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918,
         n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928,
         n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938,
         n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948,
         n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958,
         n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968,
         n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978,
         n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988,
         n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998,
         n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008,
         n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018,
         n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028,
         n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038,
         n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048,
         n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058,
         n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068,
         n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078,
         n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088,
         n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098,
         n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108,
         n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118,
         n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128,
         n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138,
         n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148,
         n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158,
         n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168,
         n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178,
         n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188,
         n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198,
         n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208,
         n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218,
         n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228,
         n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238,
         n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248,
         n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258,
         n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268,
         n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278,
         n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288,
         n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298,
         n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308,
         n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318,
         n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328,
         n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338,
         n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348,
         n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358,
         n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368,
         n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378,
         n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388,
         n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398,
         n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408,
         n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418,
         n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428,
         n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438,
         n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448,
         n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458,
         n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468,
         n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478,
         n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488,
         n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498,
         n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508,
         n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518,
         n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528,
         n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538,
         n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548,
         n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558,
         n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568,
         n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578,
         n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588,
         n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598,
         n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608,
         n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618,
         n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628,
         n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638,
         n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648,
         n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658,
         n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668,
         n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678,
         n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688,
         n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698,
         n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708,
         n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718,
         n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728,
         n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738,
         n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748,
         n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758,
         n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768,
         n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778,
         n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788,
         n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798,
         n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808,
         n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818,
         n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828,
         n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838,
         n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848,
         n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858,
         n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868,
         n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878,
         n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888,
         n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898,
         n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908,
         n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918,
         n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928,
         n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938,
         n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948,
         n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958,
         n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968,
         n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978,
         n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988,
         n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998,
         n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008,
         n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018,
         n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028,
         n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038,
         n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048,
         n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058,
         n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068,
         n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078,
         n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088,
         n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098,
         n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108,
         n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118,
         n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128,
         n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138,
         n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148,
         n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158,
         n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168,
         n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178,
         n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188,
         n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198,
         n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208,
         n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218,
         n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228,
         n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238,
         n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248,
         n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258,
         n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268,
         n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278,
         n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288,
         n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298,
         n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308,
         n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318,
         n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328,
         n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338,
         n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348,
         n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358,
         n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368,
         n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378,
         n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388,
         n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398,
         n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408,
         n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418,
         n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428,
         n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438,
         n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448,
         n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458,
         n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468,
         n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478,
         n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488,
         n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498,
         n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508,
         n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518,
         n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528,
         n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538,
         n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548,
         n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558,
         n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568,
         n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578,
         n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588,
         n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598,
         n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608,
         n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618,
         n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628,
         n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638,
         n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648,
         n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658,
         n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668,
         n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678,
         n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688,
         n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698,
         n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708,
         n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718,
         n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728,
         n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738,
         n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748,
         n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758,
         n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768,
         n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778,
         n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788,
         n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798,
         n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808,
         n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818,
         n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828,
         n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838,
         n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848,
         n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858,
         n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868,
         n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878,
         n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888,
         n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898,
         n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908,
         n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918,
         n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928,
         n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938,
         n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948,
         n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958,
         n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968,
         n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978,
         n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988,
         n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998,
         n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008,
         n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018,
         n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028,
         n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038,
         n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048,
         n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058,
         n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068,
         n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078,
         n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088,
         n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098,
         n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108,
         n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118,
         n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128,
         n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138,
         n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9149,
         n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159,
         n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169,
         n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179,
         n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189,
         n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199,
         n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209,
         n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219,
         n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229,
         n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239,
         n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249,
         n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259,
         n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9269, n9270,
         n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280,
         n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290,
         n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300,
         n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310,
         n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320,
         n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330,
         n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340,
         n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350,
         n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360,
         n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370,
         n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380,
         n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390,
         n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400,
         n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410,
         n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420,
         n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430,
         n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440,
         n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450,
         n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460,
         n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470,
         n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480,
         n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490,
         n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500,
         n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510,
         n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520,
         n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530,
         n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540,
         n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550,
         n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560,
         n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570,
         n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580,
         n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590,
         n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600,
         n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610,
         n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620,
         n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630,
         n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640,
         n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650,
         n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660,
         n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670,
         n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680,
         n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690,
         n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700,
         n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710,
         n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720,
         n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730,
         n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740,
         n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750,
         n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760,
         n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770,
         n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780,
         n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790,
         n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800,
         n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810,
         n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820,
         n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830,
         n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840,
         n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850,
         n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860,
         n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870,
         n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9881,
         n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891,
         n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901,
         n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911,
         n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921,
         n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931,
         n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941,
         n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951,
         n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961,
         n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971,
         n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981,
         n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991,
         n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245;

  AOI22_X1 U4775 ( .A1(n7519), .A2(n7520), .B1(P2_REG1_REG_12__SCAN_IN), .B2(
        n7521), .ZN(n5129) );
  XNOR2_X1 U4776 ( .A(n4808), .B(n5065), .ZN(n7047) );
  BUF_X2 U4777 ( .A(n6423), .Z(n4391) );
  INV_X1 U4778 ( .A(n9334), .ZN(n6398) );
  INV_X2 U4779 ( .A(n8504), .ZN(n8440) );
  AND2_X1 U4780 ( .A1(n6978), .A2(n5943), .ZN(n7111) );
  INV_X1 U4781 ( .A(n7103), .ZN(n7226) );
  CLKBUF_X1 U4782 ( .A(n6323), .Z(n6486) );
  BUF_X1 U4783 ( .A(n5938), .Z(n9337) );
  NOR2_X1 U4784 ( .A1(n5084), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n5087) );
  AND3_X1 U4785 ( .A1(n5977), .A2(n5975), .A3(n4349), .ZN(n7344) );
  NAND2_X1 U4786 ( .A1(n5043), .A2(n5076), .ZN(n7068) );
  NAND2_X1 U4787 ( .A1(n5875), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n6145) );
  AND2_X1 U4788 ( .A1(n5855), .A2(n5854), .ZN(n8022) );
  XNOR2_X1 U4790 ( .A(n5895), .B(P1_IR_REG_19__SCAN_IN), .ZN(n5897) );
  AND3_X1 U4791 ( .A1(n5824), .A2(n6032), .A3(n5823), .ZN(n5825) );
  INV_X1 U4792 ( .A(n9003), .ZN(n4269) );
  AND3_X2 U4793 ( .A1(n4738), .A2(n4739), .A3(n4737), .ZN(n4939) );
  XNOR2_X1 U4794 ( .A(n5495), .B(n5128), .ZN(n7474) );
  MUX2_X2 U4795 ( .A(n9175), .B(P2_REG1_REG_25__SCAN_IN), .S(n4269), .Z(n8943)
         );
  OAI21_X1 U4796 ( .B1(n7876), .B2(n8049), .A(n7875), .ZN(n7883) );
  AOI21_X1 U4797 ( .B1(n4435), .B2(n7874), .A(n4434), .ZN(n7876) );
  AOI21_X1 U4798 ( .B1(n8401), .B2(n8400), .A(n8399), .ZN(n8405) );
  NAND2_X1 U4799 ( .A1(n5938), .A2(n6000), .ZN(n5931) );
  OR2_X1 U4800 ( .A1(n6477), .A2(n8022), .ZN(n5904) );
  NAND2_X2 U4801 ( .A1(n5905), .A2(n5904), .ZN(n6000) );
  NAND2_X1 U4802 ( .A1(n4411), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n6236) );
  NAND2_X1 U4803 ( .A1(n10122), .A2(n7504), .ZN(n7807) );
  CLKBUF_X3 U4804 ( .A(n9285), .Z(n4271) );
  NAND2_X1 U4805 ( .A1(n8605), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n8640) );
  AND2_X1 U4806 ( .A1(n5740), .A2(n5739), .ZN(n6686) );
  AND2_X1 U4807 ( .A1(n8425), .A2(n8420), .ZN(n8705) );
  INV_X1 U4808 ( .A(n8435), .ZN(n5587) );
  AND2_X1 U4809 ( .A1(n7178), .A2(n8313), .ZN(n8481) );
  INV_X1 U4810 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n5023) );
  OR2_X1 U4811 ( .A1(n5032), .A2(P2_IR_REG_16__SCAN_IN), .ZN(n5103) );
  OR2_X1 U4814 ( .A1(n6030), .A2(n5228), .ZN(n5910) );
  OR2_X1 U4815 ( .A1(n6414), .A2(n6413), .ZN(n6440) );
  NOR2_X1 U4816 ( .A1(n6462), .A2(n7683), .ZN(n5869) );
  NOR2_X1 U4817 ( .A1(n9796), .A2(n9631), .ZN(n7953) );
  INV_X1 U4818 ( .A(n10017), .ZN(n9766) );
  OR2_X1 U4819 ( .A1(n9795), .A2(n4447), .ZN(n4297) );
  INV_X1 U4820 ( .A(n7493), .ZN(n10092) );
  BUF_X1 U4821 ( .A(n5360), .Z(n5794) );
  AND4_X1 U4822 ( .A1(n5433), .A2(n5432), .A3(n5431), .A4(n5430), .ZN(n8906)
         );
  INV_X1 U4823 ( .A(n8169), .ZN(n6663) );
  NAND2_X1 U4824 ( .A1(n6319), .A2(n6318), .ZN(n9829) );
  CLKBUF_X3 U4825 ( .A(n5991), .Z(n7881) );
  AND4_X1 U4826 ( .A1(n6067), .A2(n6066), .A3(n6065), .A4(n6064), .ZN(n9975)
         );
  INV_X1 U4827 ( .A(n10039), .ZN(n10027) );
  NAND2_X1 U4828 ( .A1(n6059), .A2(n6058), .ZN(n7429) );
  INV_X1 U4829 ( .A(n5794), .ZN(n6710) );
  INV_X1 U4830 ( .A(n6621), .ZN(n8537) );
  CLKBUF_X3 U4831 ( .A(n9285), .Z(n4270) );
  INV_X2 U4832 ( .A(n4984), .ZN(n10070) );
  BUF_X1 U4833 ( .A(n5349), .Z(n8456) );
  OR2_X1 U4835 ( .A1(n10000), .A2(n10001), .ZN(n10002) );
  INV_X2 U4836 ( .A(n5369), .ZN(n5429) );
  INV_X4 U4837 ( .A(n6150), .ZN(n6423) );
  AND2_X2 U4838 ( .A1(n9555), .A2(n9556), .ZN(n9553) );
  NOR2_X2 U4839 ( .A1(n5100), .A2(n4436), .ZN(n8573) );
  NAND2_X2 U4840 ( .A1(n9638), .A2(n4735), .ZN(n4734) );
  NAND2_X2 U4841 ( .A1(n9640), .A2(n9639), .ZN(n9638) );
  OAI222_X1 U4842 ( .A1(n7680), .A2(n7540), .B1(P1_U3086), .B2(n6477), .C1(
        n9897), .C2(n7539), .ZN(P1_U3334) );
  INV_X2 U4843 ( .A(n8022), .ZN(n6480) );
  NAND2_X1 U4844 ( .A1(n5438), .A2(n5271), .ZN(n5453) );
  INV_X2 U4845 ( .A(n5371), .ZN(n5379) );
  NAND2_X2 U4847 ( .A1(n5027), .A2(n5208), .ZN(n9285) );
  NAND2_X2 U4848 ( .A1(n5869), .A2(n7709), .ZN(n6738) );
  XNOR2_X2 U4849 ( .A(n5868), .B(P1_IR_REG_25__SCAN_IN), .ZN(n7709) );
  BUF_X2 U4850 ( .A(n9552), .Z(n4422) );
  NAND2_X1 U4852 ( .A1(n7226), .A2(n6963), .ZN(n8298) );
  NAND2_X2 U4853 ( .A1(n9881), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5883) );
  NAND2_X2 U4854 ( .A1(n5215), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5211) );
  NAND2_X2 U4855 ( .A1(n8721), .A2(n8473), .ZN(n8716) );
  AOI21_X2 U4856 ( .B1(P1_REG1_REG_6__SCAN_IN), .B2(n6925), .A(n6919), .ZN(
        n6935) );
  BUF_X4 U4857 ( .A(n8456), .Z(n4272) );
  NAND2_X2 U4858 ( .A1(n5909), .A2(n5936), .ZN(n5969) );
  XNOR2_X2 U4859 ( .A(n5949), .B(P1_IR_REG_2__SCAN_IN), .ZN(n9522) );
  XNOR2_X2 U4860 ( .A(n5886), .B(P1_IR_REG_29__SCAN_IN), .ZN(n9888) );
  OAI21_X1 U4861 ( .B1(n7883), .B2(n8004), .A(n4863), .ZN(n4862) );
  OAI21_X1 U4862 ( .B1(n6735), .B2(n4269), .A(n4512), .ZN(n6727) );
  OAI21_X1 U4863 ( .B1(n8423), .B2(n4907), .A(n4906), .ZN(n4905) );
  XNOR2_X1 U4864 ( .A(n5749), .B(n5747), .ZN(n8271) );
  NOR2_X1 U4865 ( .A1(n7953), .A2(n7952), .ZN(n9604) );
  NAND2_X1 U4866 ( .A1(n8565), .A2(n4437), .ZN(n8539) );
  NAND2_X1 U4867 ( .A1(n6633), .A2(n6632), .ZN(n8824) );
  NAND2_X1 U4868 ( .A1(n5713), .A2(n5712), .ZN(n5733) );
  NAND2_X1 U4869 ( .A1(n5486), .A2(n5485), .ZN(n8164) );
  NOR2_X1 U4870 ( .A1(n6752), .A2(n4678), .ZN(n9905) );
  NOR2_X1 U4871 ( .A1(n7127), .A2(n8481), .ZN(n4626) );
  AND2_X1 U4872 ( .A1(n8334), .A2(n8902), .ZN(n8479) );
  OR2_X1 U4873 ( .A1(n6625), .A2(n8898), .ZN(n8860) );
  NAND2_X2 U4874 ( .A1(n9499), .A2(n7360), .ZN(n7788) );
  NAND2_X1 U4875 ( .A1(n7344), .A2(n7493), .ZN(n10007) );
  NOR2_X1 U4876 ( .A1(n8535), .A2(n7257), .ZN(n7192) );
  NAND2_X1 U4877 ( .A1(n6807), .A2(n6555), .ZN(n6095) );
  INV_X1 U4878 ( .A(n10018), .ZN(n10096) );
  INV_X2 U4879 ( .A(n5457), .ZN(n5442) );
  AND4_X1 U4880 ( .A1(n5997), .A2(n5996), .A3(n4305), .A4(n5995), .ZN(n7356)
         );
  NOR2_X1 U4881 ( .A1(n7346), .A2(n7642), .ZN(n7637) );
  BUF_X2 U4882 ( .A(n6000), .Z(n6426) );
  INV_X1 U4883 ( .A(n8222), .ZN(n8891) );
  INV_X1 U4884 ( .A(n8889), .ZN(n8345) );
  AND4_X1 U4885 ( .A1(n5451), .A2(n5450), .A3(n5449), .A4(n5448), .ZN(n8222)
         );
  NAND4_X1 U4886 ( .A1(n5468), .A2(n5467), .A3(n5466), .A4(n5465), .ZN(n8916)
         );
  NAND2_X1 U4887 ( .A1(n6914), .A2(n7019), .ZN(n7099) );
  INV_X1 U4888 ( .A(n8538), .ZN(n6880) );
  AND4_X2 U4889 ( .A1(n5353), .A2(n5352), .A3(n5351), .A4(n5350), .ZN(n6963)
         );
  NAND4_X1 U4890 ( .A1(n5348), .A2(n5347), .A3(n5346), .A4(n5345), .ZN(n8538)
         );
  INV_X2 U4891 ( .A(n7877), .ZN(n7882) );
  CLKBUF_X2 U4893 ( .A(n5387), .Z(n8435) );
  MUX2_X1 U4894 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5834), .S(
        P1_IR_REG_27__SCAN_IN), .Z(n5839) );
  AND3_X1 U4895 ( .A1(n4989), .A2(n4988), .A3(n4987), .ZN(n4992) );
  NOR2_X1 U4896 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n5829) );
  NOR2_X1 U4897 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_16__SCAN_IN), .ZN(
        n5827) );
  NOR2_X1 U4898 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_IR_REG_20__SCAN_IN), .ZN(
        n5828) );
  INV_X2 U4899 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n5884) );
  XOR2_X1 U4900 ( .A(n9604), .B(n9602), .Z(n9798) );
  NAND2_X1 U4901 ( .A1(n5751), .A2(n4310), .ZN(n8145) );
  AND2_X1 U4902 ( .A1(n7884), .A2(n4864), .ZN(n4863) );
  NAND2_X1 U4903 ( .A1(n8271), .A2(n8178), .ZN(n5751) );
  AND2_X1 U4904 ( .A1(n4606), .A2(n8614), .ZN(n5102) );
  NAND2_X1 U4905 ( .A1(n4834), .A2(n4284), .ZN(n9602) );
  AOI21_X1 U4906 ( .B1(n5705), .B2(n5704), .A(n4535), .ZN(n4532) );
  OAI21_X1 U4907 ( .B1(n8205), .B2(n4531), .A(n4530), .ZN(n5749) );
  NOR2_X1 U4908 ( .A1(n4604), .A2(n4367), .ZN(n4603) );
  NOR2_X1 U4909 ( .A1(n8427), .A2(n8414), .ZN(n8684) );
  NAND2_X1 U4910 ( .A1(n6547), .A2(n6546), .ZN(n8004) );
  NAND2_X1 U4911 ( .A1(n9368), .A2(n4300), .ZN(n4702) );
  NAND2_X1 U4912 ( .A1(n8732), .A2(n8733), .ZN(n6681) );
  AND2_X1 U4913 ( .A1(n5761), .A2(n5760), .ZN(n6689) );
  OR2_X1 U4914 ( .A1(n5089), .A2(n8544), .ZN(n4437) );
  XNOR2_X1 U4915 ( .A(n5759), .B(n5758), .ZN(n9282) );
  AND2_X1 U4916 ( .A1(n6447), .A2(n6446), .ZN(n9631) );
  AND2_X1 U4917 ( .A1(n7853), .A2(n9705), .ZN(n8040) );
  NAND2_X1 U4918 ( .A1(n6397), .A2(n6396), .ZN(n9804) );
  NOR2_X1 U4919 ( .A1(n4445), .A2(n8636), .ZN(n4444) );
  XNOR2_X1 U4920 ( .A(n5752), .B(n6515), .ZN(n7727) );
  NOR2_X1 U4921 ( .A1(n9824), .A2(n8062), .ZN(n7889) );
  XNOR2_X1 U4922 ( .A(n5733), .B(n5732), .ZN(n7708) );
  MUX2_X1 U4923 ( .A(n8631), .B(n8630), .S(n8629), .Z(n8636) );
  NAND2_X1 U4924 ( .A1(n6029), .A2(n7313), .ZN(n7323) );
  NOR2_X1 U4925 ( .A1(n9903), .A2(n4365), .ZN(n6595) );
  XNOR2_X1 U4926 ( .A(n5627), .B(n5626), .ZN(n7517) );
  NAND2_X1 U4927 ( .A1(n5612), .A2(n5611), .ZN(n9207) );
  NOR2_X1 U4928 ( .A1(n9905), .A2(n9904), .ZN(n9903) );
  NAND2_X2 U4929 ( .A1(n4377), .A2(n5308), .ZN(n9213) );
  OAI21_X1 U4930 ( .B1(n7203), .B2(n4614), .A(n4612), .ZN(n5082) );
  NAND2_X1 U4931 ( .A1(n4497), .A2(n6296), .ZN(n9834) );
  OAI21_X1 U4932 ( .B1(n5647), .B2(n5639), .A(n5640), .ZN(n5625) );
  AND2_X1 U4933 ( .A1(n5589), .A2(n5588), .ZN(n9220) );
  NAND2_X1 U4934 ( .A1(n7288), .A2(n8450), .ZN(n4377) );
  NOR3_X1 U4935 ( .A1(n4930), .A2(n4931), .A3(n4929), .ZN(n4928) );
  OAI21_X1 U4936 ( .B1(n5669), .B2(n5668), .A(n5667), .ZN(n5700) );
  NAND2_X1 U4937 ( .A1(n4883), .A2(n4889), .ZN(n5647) );
  XNOR2_X1 U4938 ( .A(n5608), .B(n5607), .ZN(n7288) );
  NAND2_X1 U4939 ( .A1(n4880), .A2(n4884), .ZN(n5669) );
  OAI21_X1 U4940 ( .B1(n5585), .B2(n5302), .A(n5301), .ZN(n5608) );
  NAND2_X1 U4941 ( .A1(n5574), .A2(n5573), .ZN(n9223) );
  AND2_X1 U4942 ( .A1(n4754), .A2(n4753), .ZN(n7230) );
  NAND2_X1 U4943 ( .A1(n5298), .A2(n4881), .ZN(n4880) );
  NAND2_X1 U4944 ( .A1(n5298), .A2(n5297), .ZN(n5585) );
  AND2_X1 U4945 ( .A1(n7928), .A2(n7924), .ZN(n7969) );
  OAI21_X1 U4946 ( .B1(n4790), .B2(n7271), .A(n4783), .ZN(n5127) );
  OAI211_X1 U4947 ( .C1(n7077), .C2(n4794), .A(n4380), .B(
        P2_REG1_REG_9__SCAN_IN), .ZN(n4790) );
  NAND2_X1 U4948 ( .A1(n7077), .A2(n4792), .ZN(n4380) );
  INV_X1 U4949 ( .A(n10140), .ZN(n9311) );
  AND2_X1 U4950 ( .A1(n5503), .A2(n5502), .ZN(n8169) );
  OR2_X2 U4951 ( .A1(n7079), .A2(n7080), .ZN(n7077) );
  NAND2_X1 U4952 ( .A1(n6125), .A2(n6124), .ZN(n9445) );
  AND2_X1 U4953 ( .A1(n5497), .A2(n5496), .ZN(n8340) );
  AND2_X1 U4954 ( .A1(n7161), .A2(n4291), .ZN(n4755) );
  AND2_X1 U4955 ( .A1(n7788), .A2(n7914), .ZN(n7798) );
  OR2_X1 U4956 ( .A1(n5741), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n5764) );
  NAND2_X1 U4957 ( .A1(n4557), .A2(n4556), .ZN(n5512) );
  OAI21_X1 U4958 ( .B1(n7370), .B2(n7348), .A(n7371), .ZN(n10044) );
  AND2_X1 U4959 ( .A1(n8316), .A2(n8313), .ZN(n6622) );
  OR2_X1 U4960 ( .A1(n10122), .A2(n7504), .ZN(n7502) );
  NAND2_X2 U4961 ( .A1(n6095), .A2(n6094), .ZN(n10122) );
  INV_X1 U4962 ( .A(n7592), .ZN(n10104) );
  NOR2_X1 U4963 ( .A1(n4793), .A2(n4286), .ZN(n4792) );
  INV_X1 U4964 ( .A(n8302), .ZN(n8486) );
  NAND2_X1 U4965 ( .A1(n6010), .A2(n6011), .ZN(n7592) );
  INV_X1 U4966 ( .A(n5363), .ZN(n5457) );
  AND4_X1 U4967 ( .A1(n6105), .A2(n6104), .A3(n6103), .A4(n6102), .ZN(n7504)
         );
  AND4_X1 U4968 ( .A1(n6085), .A2(n6084), .A3(n6083), .A4(n6082), .ZN(n9974)
         );
  AND4_X1 U4969 ( .A1(n6017), .A2(n6018), .A3(n6016), .A4(n6019), .ZN(n7359)
         );
  AND4_X1 U4970 ( .A1(n6046), .A2(n6045), .A3(n6044), .A4(n6043), .ZN(n7586)
         );
  NAND2_X1 U4971 ( .A1(n5972), .A2(n5971), .ZN(n7493) );
  NAND4_X2 U4972 ( .A1(n5957), .A2(n5956), .A3(n5955), .A4(n5954), .ZN(n7352)
         );
  AND3_X2 U4973 ( .A1(n5344), .A2(n5343), .A3(n5342), .ZN(n10164) );
  AND4_X1 U4974 ( .A1(n5375), .A2(n5374), .A3(n5373), .A4(n5372), .ZN(n6914)
         );
  XNOR2_X1 U4975 ( .A(n5067), .B(n9109), .ZN(n5454) );
  AOI21_X1 U4976 ( .B1(n4886), .B2(n4889), .A(n4885), .ZN(n4884) );
  AOI21_X1 U4977 ( .B1(n4501), .B2(n4499), .A(n4559), .ZN(n4498) );
  NAND2_X1 U4978 ( .A1(n5866), .A2(n5865), .ZN(n7683) );
  INV_X2 U4979 ( .A(n5358), .ZN(n8450) );
  NAND2_X1 U4980 ( .A1(n5360), .A2(n6778), .ZN(n5358) );
  NAND2_X1 U4981 ( .A1(n4389), .A2(n4386), .ZN(n6462) );
  NAND2_X2 U4982 ( .A1(n8525), .A2(n8295), .ZN(n8504) );
  INV_X1 U4983 ( .A(n6099), .ZN(n5875) );
  INV_X1 U4984 ( .A(n5645), .ZN(n4885) );
  NAND2_X1 U4985 ( .A1(n5216), .A2(n9269), .ZN(n9277) );
  XNOR2_X1 U4986 ( .A(n5021), .B(n5020), .ZN(n5190) );
  NAND2_X1 U4987 ( .A1(n5214), .A2(n5213), .ZN(n5216) );
  OAI21_X1 U4988 ( .B1(n5609), .B2(n5249), .A(n5248), .ZN(n5263) );
  NAND2_X2 U4989 ( .A1(n6779), .A2(P1_U3086), .ZN(n9897) );
  OR2_X1 U4990 ( .A1(n5042), .A2(P2_IR_REG_3__SCAN_IN), .ZN(n5076) );
  INV_X1 U4991 ( .A(n4385), .ZN(n4704) );
  OR2_X1 U4992 ( .A1(n5079), .A2(P2_IR_REG_11__SCAN_IN), .ZN(n5084) );
  NAND2_X1 U4993 ( .A1(n5826), .A2(n5825), .ZN(n5844) );
  NAND2_X1 U4994 ( .A1(n4980), .A2(n4995), .ZN(n4624) );
  NAND2_X1 U4995 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n5209), .ZN(n5213) );
  NAND4_X1 U4996 ( .A1(n5846), .A2(n5828), .A3(n5827), .A4(n5829), .ZN(n4893)
         );
  NOR2_X1 U4997 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .ZN(
        n4739) );
  INV_X4 U4998 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  NOR2_X1 U4999 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n4738) );
  INV_X1 U5000 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5900) );
  NOR2_X1 U5001 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_6__SCAN_IN), .ZN(
        n5824) );
  INV_X1 U5002 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5310) );
  NOR2_X1 U5003 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n4990) );
  NOR2_X1 U5004 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), .ZN(
        n4991) );
  INV_X1 U5005 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n5008) );
  INV_X1 U5006 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5009) );
  INV_X1 U5007 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5863) );
  INV_X1 U5008 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n5210) );
  NOR2_X1 U5009 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_5__SCAN_IN), .ZN(
        n4742) );
  NOR2_X1 U5010 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_9__SCAN_IN), .ZN(
        n4740) );
  INV_X1 U5011 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5867) );
  NOR2_X1 U5012 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .ZN(
        n4741) );
  INV_X1 U5013 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n5226) );
  NOR2_X1 U5014 ( .A1(n7063), .A2(n7064), .ZN(n7062) );
  AOI21_X1 U5015 ( .B1(n8808), .B2(n8369), .A(n8367), .ZN(n8799) );
  OAI21_X1 U5016 ( .B1(n9337), .B2(n5927), .A(n5937), .ZN(n5939) );
  NAND2_X1 U5017 ( .A1(n10001), .A2(n7586), .ZN(n7794) );
  NAND2_X1 U5018 ( .A1(n4734), .A2(n4299), .ZN(n9603) );
  NAND2_X1 U5019 ( .A1(n5938), .A2(n6000), .ZN(n4273) );
  AOI21_X4 U5020 ( .B1(n7428), .B2(n7424), .A(n7425), .ZN(n9401) );
  INV_X2 U5021 ( .A(n6963), .ZN(n4967) );
  NOR2_X2 U5022 ( .A1(n6932), .A2(n6931), .ZN(n6930) );
  AND2_X2 U5023 ( .A1(n9744), .A2(n9731), .ZN(n9729) );
  AND2_X1 U5024 ( .A1(n6480), .A2(n5897), .ZN(n7949) );
  OAI21_X2 U5025 ( .B1(n7323), .B2(n6052), .A(n6055), .ZN(n7428) );
  XNOR2_X1 U5026 ( .A(n5111), .B(n5110), .ZN(n5312) );
  OAI211_X2 U5028 ( .C1(n5764), .C2(n4515), .A(n5746), .B(n4514), .ZN(n8699)
         );
  OAI21_X2 U5029 ( .B1(n8706), .B2(n4960), .A(n4957), .ZN(n8653) );
  AOI21_X2 U5030 ( .B1(n8716), .B2(n8428), .A(n8472), .ZN(n8706) );
  NAND2_X1 U5031 ( .A1(n7978), .A2(n7867), .ZN(n7898) );
  NAND2_X1 U5032 ( .A1(n5529), .A2(SI_14_), .ZN(n4879) );
  OR2_X1 U5033 ( .A1(n9834), .A2(n9717), .ZN(n7956) );
  OR2_X1 U5034 ( .A1(n5994), .A2(n5913), .ZN(n5917) );
  OR2_X1 U5035 ( .A1(n5992), .A2(n9502), .ZN(n5918) );
  NAND2_X1 U5036 ( .A1(n6041), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5915) );
  AND4_X1 U5037 ( .A1(n5540), .A2(n5539), .A3(n5538), .A4(n5537), .ZN(n6667)
         );
  NAND2_X1 U5038 ( .A1(n6854), .A2(n6855), .ZN(n6853) );
  AND2_X1 U5039 ( .A1(n7940), .A2(n7943), .ZN(n8077) );
  OR2_X1 U5040 ( .A1(n8015), .A2(n9891), .ZN(n10048) );
  AND2_X1 U5041 ( .A1(n6500), .A2(n9891), .ZN(n10010) );
  NAND2_X1 U5042 ( .A1(n4919), .A2(n4918), .ZN(n8300) );
  NAND2_X1 U5043 ( .A1(n8296), .A2(n8295), .ZN(n4919) );
  NAND2_X1 U5044 ( .A1(n8297), .A2(n7518), .ZN(n4918) );
  AND2_X1 U5045 ( .A1(n8881), .A2(n8328), .ZN(n8330) );
  INV_X1 U5046 ( .A(n6682), .ZN(n4656) );
  AOI21_X1 U5047 ( .B1(n4891), .B2(n5302), .A(n4890), .ZN(n4889) );
  INV_X1 U5048 ( .A(n5606), .ZN(n4890) );
  INV_X1 U5049 ( .A(n4879), .ZN(n4878) );
  AOI21_X1 U5050 ( .B1(n4748), .B2(n4749), .A(n4746), .ZN(n4745) );
  INV_X1 U5051 ( .A(n8098), .ZN(n4746) );
  AND2_X1 U5052 ( .A1(n8411), .A2(n8417), .ZN(n4904) );
  INV_X1 U5053 ( .A(n4613), .ZN(n4612) );
  OAI21_X1 U5054 ( .B1(n7280), .B2(n4614), .A(n5078), .ZN(n4613) );
  NAND2_X1 U5055 ( .A1(n5083), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n4609) );
  NOR2_X1 U5056 ( .A1(n5460), .A2(n7271), .ZN(n4788) );
  AND2_X1 U5057 ( .A1(n9165), .A2(n8274), .ZN(n8413) );
  OR2_X1 U5058 ( .A1(n9165), .A2(n8274), .ZN(n8430) );
  OR2_X1 U5059 ( .A1(n4986), .A2(n6691), .ZN(n8669) );
  NAND2_X1 U5060 ( .A1(n9171), .A2(n8178), .ZN(n8417) );
  AND2_X1 U5061 ( .A1(n6686), .A2(n8699), .ZN(n8427) );
  INV_X1 U5062 ( .A(n6679), .ZN(n4638) );
  NOR2_X1 U5063 ( .A1(n6671), .A2(n4645), .ZN(n4644) );
  INV_X1 U5064 ( .A(n6668), .ZN(n4645) );
  OR2_X1 U5065 ( .A1(n9223), .A2(n8778), .ZN(n8375) );
  OR2_X1 U5066 ( .A1(n9229), .A2(n8286), .ZN(n8371) );
  AND2_X1 U5067 ( .A1(n7873), .A2(n7877), .ZN(n4434) );
  NOR2_X1 U5068 ( .A1(n9629), .A2(n4736), .ZN(n4735) );
  INV_X1 U5069 ( .A(n8045), .ZN(n4736) );
  AND2_X1 U5070 ( .A1(n9796), .A2(n9631), .ZN(n7952) );
  OR2_X1 U5071 ( .A1(n9809), .A2(n9673), .ZN(n8044) );
  NOR2_X1 U5072 ( .A1(n9311), .A2(n9407), .ZN(n4896) );
  NOR2_X1 U5073 ( .A1(n9660), .A2(n4899), .ZN(n9595) );
  INV_X1 U5074 ( .A(n4901), .ZN(n4900) );
  INV_X1 U5075 ( .A(n9657), .ZN(n9630) );
  NAND2_X1 U5076 ( .A1(n6513), .A2(n6511), .ZN(n5752) );
  AND2_X1 U5077 ( .A1(n6510), .A2(n5738), .ZN(n6515) );
  NAND2_X1 U5078 ( .A1(n4704), .A2(n4703), .ZN(n6201) );
  AND2_X1 U5079 ( .A1(n4293), .A2(n5845), .ZN(n4703) );
  NAND2_X1 U5080 ( .A1(n4875), .A2(n4879), .ZN(n5557) );
  OAI21_X1 U5081 ( .B1(n5494), .B2(n4549), .A(n4331), .ZN(n4875) );
  NAND2_X1 U5082 ( .A1(n4555), .A2(n4550), .ZN(n4549) );
  XNOR2_X1 U5083 ( .A(n5275), .B(SI_9_), .ZN(n5458) );
  OR2_X1 U5084 ( .A1(n6138), .A2(P1_IR_REG_10__SCAN_IN), .ZN(n6163) );
  NOR2_X1 U5085 ( .A1(n5324), .A2(n5256), .ZN(n5255) );
  INV_X1 U5086 ( .A(n5603), .ZN(n4762) );
  NOR2_X1 U5087 ( .A1(n5484), .A2(n4770), .ZN(n4769) );
  NOR2_X1 U5088 ( .A1(n5443), .A2(n4771), .ZN(n4770) );
  AOI21_X1 U5089 ( .B1(n4533), .B2(n4535), .A(n4321), .ZN(n4530) );
  INV_X1 U5090 ( .A(n4533), .ZN(n4531) );
  INV_X1 U5091 ( .A(n6644), .ZN(n4515) );
  NAND2_X1 U5092 ( .A1(n6853), .A2(n5118), .ZN(n5120) );
  OR2_X1 U5093 ( .A1(n5797), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n8088) );
  NAND2_X1 U5094 ( .A1(n5722), .A2(n5721), .ZN(n5741) );
  INV_X1 U5095 ( .A(n5723), .ZN(n5722) );
  NAND2_X1 U5096 ( .A1(n8791), .A2(n8789), .ZN(n6669) );
  NAND2_X1 U5097 ( .A1(n6802), .A2(n5808), .ZN(n6715) );
  NAND2_X1 U5098 ( .A1(n6643), .A2(n6642), .ZN(n6726) );
  XNOR2_X1 U5099 ( .A(n9159), .B(n8470), .ZN(n8655) );
  NAND2_X1 U5100 ( .A1(n8673), .A2(n8917), .ZN(n8675) );
  OR2_X1 U5101 ( .A1(n9178), .A2(n8711), .ZN(n8425) );
  INV_X1 U5102 ( .A(n4663), .ZN(n4662) );
  OAI21_X1 U5103 ( .B1(n4665), .B2(n4664), .A(n8365), .ZN(n4663) );
  INV_X1 U5104 ( .A(n4668), .ZN(n4667) );
  OAI21_X1 U5105 ( .B1(n8477), .B2(n8476), .A(n4322), .ZN(n4668) );
  OR2_X1 U5106 ( .A1(n9248), .A2(n8847), .ZN(n6632) );
  NAND2_X1 U5107 ( .A1(n8836), .A2(n6631), .ZN(n6633) );
  NAND2_X1 U5108 ( .A1(n7542), .A2(n7518), .ZN(n7396) );
  INV_X1 U5109 ( .A(n6161), .ZN(n5907) );
  AND2_X1 U5110 ( .A1(n4695), .A2(n6395), .ZN(n4691) );
  INV_X1 U5111 ( .A(n6221), .ZN(n5876) );
  INV_X1 U5112 ( .A(n6563), .ZN(n7878) );
  NAND2_X1 U5113 ( .A1(n9885), .A2(n5887), .ZN(n5994) );
  NAND2_X1 U5114 ( .A1(n9885), .A2(n9888), .ZN(n5992) );
  NAND2_X1 U5115 ( .A1(n9587), .A2(n9586), .ZN(n9588) );
  AOI21_X1 U5116 ( .B1(n4829), .B2(n4830), .A(n4827), .ZN(n4826) );
  NAND2_X1 U5117 ( .A1(n9683), .A2(n8041), .ZN(n9671) );
  AND2_X1 U5118 ( .A1(n8040), .A2(n4716), .ZN(n4721) );
  NAND2_X1 U5119 ( .A1(n7997), .A2(n9727), .ZN(n4716) );
  NAND2_X1 U5120 ( .A1(n4337), .A2(n4822), .ZN(n4815) );
  NAND2_X1 U5121 ( .A1(n9724), .A2(n9740), .ZN(n4822) );
  INV_X1 U5122 ( .A(n8061), .ZN(n4817) );
  NAND2_X1 U5123 ( .A1(n9834), .A2(n9754), .ZN(n4823) );
  NAND2_X1 U5124 ( .A1(n7834), .A2(n9772), .ZN(n4824) );
  OAI22_X2 U5125 ( .A1(n9760), .A2(n8059), .B1(n9755), .B2(n9843), .ZN(n9743)
         );
  NAND2_X1 U5126 ( .A1(n10053), .A2(n10078), .ZN(n10136) );
  AND2_X1 U5127 ( .A1(n6738), .A2(n6737), .ZN(n6818) );
  XNOR2_X1 U5128 ( .A(n6007), .B(P1_IR_REG_4__SCAN_IN), .ZN(n9552) );
  INV_X1 U5129 ( .A(n8724), .ZN(n8747) );
  NAND2_X1 U5130 ( .A1(n8053), .A2(n8052), .ZN(n8054) );
  OAI21_X1 U5131 ( .B1(n8311), .B2(n8310), .A(n8309), .ZN(n8319) );
  AND2_X1 U5132 ( .A1(n4920), .A2(n4913), .ZN(n8311) );
  NAND2_X1 U5133 ( .A1(n8303), .A2(n8304), .ZN(n4920) );
  AOI21_X1 U5134 ( .B1(n4398), .B2(n4302), .A(n8504), .ZN(n8338) );
  OR2_X1 U5135 ( .A1(n8387), .A2(n4424), .ZN(n4376) );
  NAND2_X1 U5136 ( .A1(n4426), .A2(n4425), .ZN(n4424) );
  NAND2_X1 U5137 ( .A1(n7865), .A2(n7864), .ZN(n7870) );
  AND2_X1 U5138 ( .A1(n6510), .A2(n6509), .ZN(n6514) );
  AOI21_X1 U5139 ( .B1(n8408), .B2(n8409), .A(n4332), .ZN(n4460) );
  NOR2_X1 U5140 ( .A1(n8744), .A2(n4450), .ZN(n4449) );
  NOR2_X1 U5141 ( .A1(n8733), .A2(n4452), .ZN(n4451) );
  INV_X1 U5142 ( .A(n8755), .ZN(n4453) );
  INV_X1 U5143 ( .A(n6652), .ZN(n4627) );
  NOR2_X1 U5144 ( .A1(n4633), .A2(n7192), .ZN(n4632) );
  NOR2_X1 U5145 ( .A1(n6688), .A2(n4652), .ZN(n4651) );
  INV_X1 U5146 ( .A(n6684), .ZN(n4652) );
  OR2_X1 U5147 ( .A1(n8668), .A2(n6687), .ZN(n6688) );
  AND2_X1 U5148 ( .A1(n7181), .A2(n7136), .ZN(n4633) );
  OR2_X1 U5149 ( .A1(n7136), .A2(n7181), .ZN(n4635) );
  NOR2_X1 U5150 ( .A1(n4893), .A2(n5831), .ZN(n5832) );
  NAND2_X1 U5151 ( .A1(n5733), .A2(n5732), .ZN(n6513) );
  NOR2_X2 U5152 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), .ZN(
        n5846) );
  NOR2_X1 U5153 ( .A1(n5607), .A2(n4892), .ZN(n4891) );
  INV_X1 U5154 ( .A(n5301), .ZN(n4892) );
  NAND2_X1 U5155 ( .A1(n5304), .A2(n5303), .ZN(n5606) );
  INV_X1 U5156 ( .A(n5570), .ZN(n4483) );
  OAI21_X1 U5157 ( .B1(n4276), .B2(n4878), .A(n5285), .ZN(n4877) );
  INV_X1 U5158 ( .A(n5291), .ZN(n4874) );
  NAND2_X1 U5159 ( .A1(n5294), .A2(n5293), .ZN(n5297) );
  NAND2_X1 U5160 ( .A1(n5609), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n5248) );
  INV_X1 U5161 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4488) );
  INV_X1 U5162 ( .A(P2_RD_REG_SCAN_IN), .ZN(n5224) );
  AOI211_X1 U5163 ( .C1(n5526), .C2(n5525), .A(n8235), .B(n8238), .ZN(n5527)
         );
  NAND2_X1 U5164 ( .A1(n5597), .A2(n4548), .ZN(n4547) );
  INV_X1 U5165 ( .A(n8195), .ZN(n4548) );
  INV_X1 U5166 ( .A(n7139), .ZN(n4752) );
  AOI21_X1 U5167 ( .B1(n4788), .B2(n4786), .A(n4359), .ZN(n4785) );
  INV_X1 U5168 ( .A(n4798), .ZN(n4786) );
  INV_X1 U5169 ( .A(n5096), .ZN(n4598) );
  NAND2_X1 U5170 ( .A1(n4590), .A2(n4591), .ZN(n4589) );
  OR2_X1 U5171 ( .A1(n6726), .A2(n8531), .ZN(n8500) );
  AND2_X1 U5172 ( .A1(n9191), .A2(n8712), .ZN(n8403) );
  NOR2_X1 U5173 ( .A1(n4281), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n5614) );
  NOR2_X1 U5174 ( .A1(n5565), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n4516) );
  INV_X1 U5175 ( .A(n5504), .ZN(n5203) );
  INV_X1 U5176 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n4520) );
  INV_X1 U5177 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n5200) );
  INV_X1 U5178 ( .A(n5427), .ZN(n5201) );
  INV_X1 U5179 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n4521) );
  INV_X1 U5180 ( .A(n8430), .ZN(n4958) );
  INV_X1 U5181 ( .A(n4965), .ZN(n4959) );
  AND2_X1 U5182 ( .A1(n8945), .A2(n8725), .ZN(n8472) );
  NOR2_X1 U5183 ( .A1(n6683), .A2(n4659), .ZN(n4658) );
  INV_X1 U5184 ( .A(n6680), .ZN(n4659) );
  OR2_X1 U5185 ( .A1(n9191), .A2(n8712), .ZN(n8473) );
  OR2_X1 U5186 ( .A1(n8954), .A2(n8253), .ZN(n8400) );
  OR2_X1 U5187 ( .A1(n9207), .A2(n8769), .ZN(n8398) );
  NOR2_X1 U5188 ( .A1(n4949), .A2(n4948), .ZN(n4947) );
  INV_X1 U5189 ( .A(n8474), .ZN(n4953) );
  INV_X1 U5190 ( .A(n8503), .ZN(n6702) );
  NOR2_X1 U5191 ( .A1(n4323), .A2(P2_IR_REG_25__SCAN_IN), .ZN(n4971) );
  INV_X1 U5192 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n5019) );
  NOR2_X1 U5193 ( .A1(n5309), .A2(P2_IR_REG_20__SCAN_IN), .ZN(n5014) );
  OR2_X1 U5194 ( .A1(n5056), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n5059) );
  INV_X1 U5195 ( .A(n6259), .ZN(n4701) );
  INV_X1 U5196 ( .A(n7698), .ZN(n4684) );
  OR2_X1 U5197 ( .A1(n8085), .A2(n9591), .ZN(n7940) );
  INV_X1 U5198 ( .A(n9642), .ZN(n8074) );
  OR2_X1 U5199 ( .A1(n9804), .A2(n9630), .ZN(n8045) );
  NOR2_X1 U5200 ( .A1(n9848), .A2(n9852), .ZN(n4894) );
  NAND2_X1 U5201 ( .A1(n9852), .A2(n9491), .ZN(n4860) );
  NOR2_X1 U5202 ( .A1(n9852), .A2(n9491), .ZN(n7714) );
  INV_X1 U5203 ( .A(n7686), .ZN(n4858) );
  AND2_X1 U5204 ( .A1(n4338), .A2(n4841), .ZN(n4839) );
  NOR2_X1 U5205 ( .A1(n7456), .A2(n7457), .ZN(n4837) );
  NAND2_X1 U5206 ( .A1(n9445), .A2(n7457), .ZN(n7825) );
  NAND2_X1 U5207 ( .A1(n7584), .A2(n7912), .ZN(n7407) );
  AND2_X1 U5208 ( .A1(n7910), .A2(n7906), .ZN(n4975) );
  OAI21_X1 U5209 ( .B1(n4985), .B2(n4712), .A(n10007), .ZN(n4711) );
  AND2_X1 U5210 ( .A1(n10044), .A2(n7905), .ZN(n4710) );
  NAND2_X1 U5211 ( .A1(n9500), .A2(n10096), .ZN(n7910) );
  OR2_X1 U5212 ( .A1(n7353), .A2(n7352), .ZN(n7491) );
  AND2_X1 U5213 ( .A1(n6572), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6737) );
  INV_X1 U5215 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n4390) );
  INV_X1 U5216 ( .A(n5860), .ZN(n4388) );
  NAND2_X1 U5217 ( .A1(n5676), .A2(n5675), .ZN(n5711) );
  NAND2_X1 U5218 ( .A1(n5700), .A2(n5699), .ZN(n5676) );
  AND2_X1 U5219 ( .A1(n5712), .A2(n5680), .ZN(n5710) );
  NAND2_X1 U5220 ( .A1(n5649), .A2(n5648), .ZN(n5667) );
  INV_X1 U5221 ( .A(n5279), .ZN(n4502) );
  INV_X1 U5222 ( .A(n4870), .ZN(n4499) );
  NAND2_X1 U5223 ( .A1(n5277), .A2(SI_10_), .ZN(n5279) );
  AND2_X1 U5224 ( .A1(n5278), .A2(n5276), .ZN(n4870) );
  INV_X1 U5225 ( .A(n5470), .ZN(n5278) );
  OAI21_X1 U5226 ( .B1(n6779), .B2(n4463), .A(n4462), .ZN(n5269) );
  NAND2_X1 U5227 ( .A1(n6779), .A2(P2_DATAO_REG_7__SCAN_IN), .ZN(n4462) );
  NAND2_X1 U5228 ( .A1(n4421), .A2(n4420), .ZN(n6031) );
  INV_X1 U5229 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n4420) );
  INV_X1 U5230 ( .A(n5987), .ZN(n4421) );
  OAI21_X1 U5231 ( .B1(n5609), .B2(P1_DATAO_REG_4__SCAN_IN), .A(n5242), .ZN(
        n5259) );
  INV_X1 U5232 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n5936) );
  NAND2_X1 U5233 ( .A1(n4765), .A2(n4764), .ZN(n4763) );
  INV_X1 U5234 ( .A(n5604), .ZN(n4764) );
  INV_X1 U5235 ( .A(n5709), .ZN(n4535) );
  NOR2_X1 U5236 ( .A1(n4758), .A2(n8229), .ZN(n4757) );
  AND2_X1 U5237 ( .A1(n4773), .A2(n4767), .ZN(n4766) );
  NOR2_X1 U5238 ( .A1(n4298), .A2(n4774), .ZN(n4773) );
  NAND2_X1 U5239 ( .A1(n4769), .A2(n4771), .ZN(n4767) );
  NAND2_X1 U5240 ( .A1(n4747), .A2(n4745), .ZN(n5544) );
  AND2_X1 U5241 ( .A1(n5036), .A2(n4810), .ZN(n4620) );
  OAI21_X1 U5242 ( .B1(n4270), .B2(n4468), .A(n4467), .ZN(n5135) );
  NAND2_X1 U5243 ( .A1(n9285), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n4467) );
  NAND2_X1 U5244 ( .A1(n5122), .A2(n5121), .ZN(n7030) );
  NAND2_X1 U5245 ( .A1(n7065), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5122) );
  NAND2_X1 U5246 ( .A1(n4615), .A2(n6890), .ZN(n6894) );
  NAND2_X1 U5247 ( .A1(n6887), .A2(n4809), .ZN(n4808) );
  OR2_X1 U5248 ( .A1(n6804), .A2(n9137), .ZN(n4809) );
  AND2_X1 U5249 ( .A1(n4972), .A2(n7280), .ZN(n7204) );
  OAI21_X1 U5250 ( .B1(n7208), .B2(n7207), .A(n7206), .ZN(n7275) );
  NAND2_X1 U5251 ( .A1(n5072), .A2(n4796), .ZN(n7280) );
  OR2_X1 U5252 ( .A1(n5454), .A2(n5126), .ZN(n4798) );
  NAND2_X1 U5253 ( .A1(n5081), .A2(n5495), .ZN(n5083) );
  NAND2_X1 U5254 ( .A1(n5089), .A2(n8544), .ZN(n8565) );
  AND2_X1 U5255 ( .A1(n5099), .A2(n5553), .ZN(n4436) );
  NAND2_X1 U5256 ( .A1(n8573), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n8599) );
  NAND2_X1 U5257 ( .A1(n5182), .A2(n5183), .ZN(n8628) );
  NAND2_X1 U5258 ( .A1(n8627), .A2(n5586), .ZN(n8624) );
  INV_X1 U5259 ( .A(n8403), .ZN(n8715) );
  NAND2_X1 U5260 ( .A1(n5614), .A2(n4522), .ZN(n5693) );
  AND2_X1 U5261 ( .A1(n4524), .A2(n4523), .ZN(n4522) );
  INV_X1 U5262 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n4523) );
  NOR2_X1 U5263 ( .A1(n6634), .A2(n8368), .ZN(n4956) );
  AOI21_X1 U5264 ( .B1(n8377), .B2(n8381), .A(n4945), .ZN(n4955) );
  INV_X1 U5265 ( .A(n8375), .ZN(n4945) );
  NAND2_X1 U5266 ( .A1(n5203), .A2(n9113), .ZN(n5519) );
  OR2_X1 U5267 ( .A1(n5487), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5504) );
  OR2_X1 U5268 ( .A1(n5477), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5487) );
  OR2_X1 U5269 ( .A1(n5441), .A2(n5440), .ZN(n7445) );
  OR2_X1 U5270 ( .A1(n5419), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5427) );
  NAND2_X1 U5271 ( .A1(n4937), .A2(n6969), .ZN(n8293) );
  NAND2_X1 U5272 ( .A1(n8656), .A2(n8917), .ZN(n8658) );
  AND2_X1 U5273 ( .A1(n8429), .A2(n8430), .ZN(n8671) );
  OR2_X1 U5274 ( .A1(n8667), .A2(n8668), .ZN(n8670) );
  INV_X1 U5275 ( .A(n8671), .ZN(n8665) );
  NOR2_X1 U5276 ( .A1(n8427), .A2(n4966), .ZN(n4965) );
  INV_X1 U5277 ( .A(n8425), .ZN(n4966) );
  AOI21_X1 U5278 ( .B1(n8420), .B2(n8417), .A(n8427), .ZN(n4964) );
  NAND2_X1 U5279 ( .A1(n8686), .A2(n8917), .ZN(n8689) );
  INV_X1 U5280 ( .A(n8417), .ZN(n8414) );
  OR2_X1 U5281 ( .A1(n8667), .A2(n8705), .ZN(n8696) );
  AOI21_X1 U5282 ( .B1(n4640), .B2(n4643), .A(n4638), .ZN(n4637) );
  INV_X1 U5283 ( .A(n6670), .ZN(n4643) );
  NAND2_X1 U5284 ( .A1(n8402), .A2(n8404), .ZN(n8733) );
  AND3_X1 U5285 ( .A1(n5594), .A2(n5593), .A3(n5592), .ZN(n8768) );
  INV_X1 U5286 ( .A(n8917), .ZN(n8848) );
  OR2_X1 U5287 ( .A1(n6708), .A2(n8504), .ZN(n8905) );
  OAI21_X1 U5288 ( .B1(n4955), .B2(n4953), .A(n8384), .ZN(n4949) );
  NOR2_X1 U5289 ( .A1(n4953), .A2(n4954), .ZN(n4951) );
  INV_X1 U5290 ( .A(n4956), .ZN(n4954) );
  AOI21_X1 U5292 ( .B1(n4667), .B2(n8477), .A(n4329), .ZN(n4665) );
  AND2_X1 U5293 ( .A1(n8365), .A2(n8364), .ZN(n8809) );
  NAND2_X1 U5294 ( .A1(n6666), .A2(n6665), .ZN(n8828) );
  NAND2_X1 U5295 ( .A1(n8169), .A2(n8355), .ZN(n6665) );
  NAND2_X1 U5296 ( .A1(n4969), .A2(n4968), .ZN(n8843) );
  AND2_X1 U5297 ( .A1(n6708), .A2(n8440), .ZN(n8917) );
  INV_X1 U5298 ( .A(n8905), .ZN(n8890) );
  OR3_X1 U5299 ( .A1(n4274), .A2(n8525), .A3(n6702), .ZN(n7397) );
  INV_X1 U5300 ( .A(n8887), .ZN(n8911) );
  NOR2_X1 U5301 ( .A1(P2_IR_REG_24__SCAN_IN), .A2(P2_IR_REG_25__SCAN_IN), .ZN(
        n4933) );
  AND2_X1 U5302 ( .A1(n4939), .A2(n4980), .ZN(n4446) );
  INV_X1 U5303 ( .A(n5079), .ZN(n4934) );
  NAND2_X1 U5304 ( .A1(n5038), .A2(n5037), .ZN(n5042) );
  NAND2_X1 U5305 ( .A1(n6198), .A2(n6197), .ZN(n9368) );
  BUF_X1 U5306 ( .A(n6150), .Z(n6389) );
  NAND2_X1 U5307 ( .A1(n4413), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n6401) );
  OR2_X1 U5308 ( .A1(n7769), .A2(n7756), .ZN(n4699) );
  NAND2_X1 U5309 ( .A1(n4698), .A2(n4696), .ZN(n4695) );
  INV_X1 U5310 ( .A(n6394), .ZN(n4696) );
  INV_X1 U5311 ( .A(n6169), .ZN(n4411) );
  NOR2_X1 U5312 ( .A1(n4684), .A2(n4681), .ZN(n4680) );
  INV_X1 U5313 ( .A(n6152), .ZN(n4681) );
  OR2_X1 U5314 ( .A1(n4684), .A2(n6160), .ZN(n4683) );
  CLKBUF_X1 U5315 ( .A(n9307), .Z(n9308) );
  XNOR2_X1 U5316 ( .A(n4459), .B(n9335), .ZN(n5944) );
  OR2_X1 U5317 ( .A1(n9337), .A2(n5961), .ZN(n5963) );
  XNOR2_X1 U5318 ( .A(n5960), .B(n9335), .ZN(n5966) );
  AND2_X1 U5319 ( .A1(n7946), .A2(n8010), .ZN(n8018) );
  AND4_X1 U5320 ( .A1(n6244), .A2(n6243), .A3(n6242), .A4(n6241), .ZN(n9425)
         );
  OR2_X1 U5321 ( .A1(n6924), .A2(n6923), .ZN(n4574) );
  NOR2_X1 U5322 ( .A1(n6945), .A2(n4676), .ZN(n9567) );
  AND2_X1 U5323 ( .A1(n6948), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n4676) );
  AND2_X1 U5324 ( .A1(n6745), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n4675) );
  OR2_X1 U5325 ( .A1(n6756), .A2(n6757), .ZN(n4571) );
  AND2_X1 U5326 ( .A1(n4571), .A2(n4570), .ZN(n9902) );
  NAND2_X1 U5327 ( .A1(n6758), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n4570) );
  OR2_X1 U5328 ( .A1(n9902), .A2(n9901), .ZN(n4569) );
  INV_X1 U5329 ( .A(n4565), .ZN(n4564) );
  AOI21_X1 U5330 ( .B1(n4563), .B2(n4565), .A(n4562), .ZN(n4561) );
  NOR2_X1 U5331 ( .A1(n9660), .A2(n4901), .ZN(n9624) );
  NAND2_X1 U5332 ( .A1(n6412), .A2(n6411), .ZN(n9800) );
  INV_X1 U5333 ( .A(n4730), .ZN(n4729) );
  OAI21_X1 U5334 ( .B1(n4732), .B2(n9668), .A(n8044), .ZN(n4730) );
  NAND2_X1 U5335 ( .A1(n4855), .A2(n4847), .ZN(n4846) );
  INV_X1 U5336 ( .A(n4851), .ZN(n4847) );
  OR2_X1 U5337 ( .A1(n4849), .A2(n8069), .ZN(n4845) );
  INV_X1 U5338 ( .A(n4850), .ZN(n4849) );
  OAI21_X1 U5339 ( .B1(n4851), .B2(n4853), .A(n8070), .ZN(n4850) );
  AND2_X1 U5340 ( .A1(n8045), .A2(n7954), .ZN(n9639) );
  NAND2_X1 U5341 ( .A1(n9655), .A2(n8042), .ZN(n4732) );
  NOR2_X1 U5342 ( .A1(n9669), .A2(n8043), .ZN(n9656) );
  OAI22_X1 U5343 ( .A1(n8068), .A2(n4852), .B1(n9679), .B2(n8067), .ZN(n4851)
         );
  NAND2_X1 U5344 ( .A1(n8066), .A2(n8065), .ZN(n4852) );
  NOR2_X1 U5345 ( .A1(n8068), .A2(n4854), .ZN(n4853) );
  INV_X1 U5346 ( .A(n8065), .ZN(n4854) );
  NOR2_X1 U5347 ( .A1(n9671), .A2(n9670), .ZN(n9669) );
  NOR2_X1 U5348 ( .A1(n8039), .A2(n4719), .ZN(n4718) );
  INV_X1 U5349 ( .A(n9684), .ZN(n4719) );
  OR2_X1 U5350 ( .A1(n8063), .A2(n8062), .ZN(n4977) );
  NOR2_X1 U5351 ( .A1(n4815), .A2(n4311), .ZN(n4813) );
  NAND2_X1 U5352 ( .A1(n4819), .A2(n4823), .ZN(n4818) );
  INV_X1 U5353 ( .A(n4821), .ZN(n4819) );
  AOI21_X1 U5354 ( .B1(n4824), .B2(n8060), .A(n4327), .ZN(n4821) );
  INV_X1 U5355 ( .A(n6299), .ZN(n5878) );
  NAND2_X1 U5356 ( .A1(n7956), .A2(n7997), .ZN(n9727) );
  AND2_X1 U5358 ( .A1(n7842), .A2(n7991), .ZN(n8057) );
  OR2_X1 U5359 ( .A1(n7685), .A2(n9425), .ZN(n4979) );
  AND4_X1 U5360 ( .A1(n6225), .A2(n6224), .A3(n6223), .A4(n6222), .ZN(n9291)
         );
  NAND2_X1 U5361 ( .A1(n7461), .A2(n7459), .ZN(n4840) );
  NAND2_X1 U5362 ( .A1(n10140), .A2(n7506), .ZN(n4841) );
  AND2_X1 U5363 ( .A1(n7822), .A2(n7825), .ZN(n7968) );
  AND2_X1 U5364 ( .A1(n9984), .A2(n4896), .ZN(n7562) );
  AND2_X1 U5365 ( .A1(n4835), .A2(n4292), .ZN(n7554) );
  INV_X1 U5366 ( .A(n10010), .ZN(n10050) );
  OR2_X1 U5367 ( .A1(n10062), .A2(n8022), .ZN(n10039) );
  NAND2_X1 U5368 ( .A1(n7346), .A2(n10058), .ZN(n10035) );
  INV_X1 U5369 ( .A(n10048), .ZN(n10009) );
  INV_X1 U5370 ( .A(n9579), .ZN(n7946) );
  NAND2_X1 U5371 ( .A1(n6437), .A2(n6436), .ZN(n9796) );
  NAND2_X1 U5372 ( .A1(n6282), .A2(n6281), .ZN(n7834) );
  XNOR2_X1 U5373 ( .A(n6554), .B(n6553), .ZN(n9267) );
  OAI21_X1 U5374 ( .B1(n6550), .B2(n6549), .A(n6548), .ZN(n6554) );
  XNOR2_X1 U5375 ( .A(n6550), .B(n6549), .ZN(n9272) );
  XNOR2_X1 U5376 ( .A(n6530), .B(n6529), .ZN(n9275) );
  XNOR2_X1 U5377 ( .A(n5711), .B(n5710), .ZN(n7669) );
  NAND2_X1 U5378 ( .A1(n4704), .A2(n4293), .ZN(n6199) );
  NAND3_X1 U5379 ( .A1(n4537), .A2(n4536), .A3(n4538), .ZN(n7157) );
  NAND2_X1 U5380 ( .A1(n4540), .A2(n4539), .ZN(n4538) );
  OR2_X1 U5381 ( .A1(n5557), .A2(n4544), .ZN(n4537) );
  XNOR2_X1 U5382 ( .A(n5515), .B(n4283), .ZN(n6180) );
  AND2_X1 U5383 ( .A1(n6140), .A2(n6163), .ZN(n6770) );
  AND2_X1 U5384 ( .A1(n5267), .A2(n5413), .ZN(n5268) );
  OR2_X1 U5385 ( .A1(n6056), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n6118) );
  AOI21_X1 U5386 ( .B1(n5385), .B2(n5326), .A(n5325), .ZN(n5328) );
  INV_X1 U5387 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n5909) );
  OAI21_X1 U5388 ( .B1(n8164), .B2(n4749), .A(n4748), .ZN(n8097) );
  AND2_X1 U5389 ( .A1(n5690), .A2(n5689), .ZN(n8702) );
  INV_X1 U5390 ( .A(n8734), .ZN(n8712) );
  AND2_X1 U5391 ( .A1(n5729), .A2(n5728), .ZN(n8711) );
  AND2_X1 U5392 ( .A1(n5653), .A2(n5652), .ZN(n8259) );
  AND3_X1 U5393 ( .A1(n5579), .A2(n5578), .A3(n5577), .ZN(n8778) );
  AND2_X1 U5394 ( .A1(n5770), .A2(n5769), .ZN(n8274) );
  NAND2_X1 U5395 ( .A1(n5791), .A2(n10165), .ZN(n8276) );
  AND3_X1 U5396 ( .A1(n5569), .A2(n5568), .A3(n5567), .ZN(n8286) );
  NAND2_X1 U5397 ( .A1(n5803), .A2(n5802), .ZN(n8673) );
  INV_X1 U5398 ( .A(n8274), .ZN(n8686) );
  OR2_X1 U5399 ( .A1(n5742), .A2(n4515), .ZN(n4514) );
  INV_X1 U5400 ( .A(n8711), .ZN(n8687) );
  INV_X1 U5401 ( .A(n8702), .ZN(n8725) );
  NAND2_X1 U5402 ( .A1(n5660), .A2(n5659), .ZN(n8724) );
  NAND2_X1 U5403 ( .A1(n5223), .A2(n5222), .ZN(n8757) );
  INV_X1 U5404 ( .A(n8286), .ZN(n8811) );
  INV_X1 U5405 ( .A(n6667), .ZN(n8830) );
  INV_X1 U5406 ( .A(P2_U3893), .ZN(n8623) );
  OR2_X1 U5407 ( .A1(P2_U3150), .A2(n5194), .ZN(n8634) );
  AOI21_X1 U5408 ( .B1(n7047), .B2(P2_REG1_REG_7__SCAN_IN), .A(n4807), .ZN(
        n7079) );
  AND2_X1 U5409 ( .A1(n4808), .A2(n6791), .ZN(n4807) );
  OR2_X1 U5410 ( .A1(n4798), .A2(n4796), .ZN(n4795) );
  NAND2_X1 U5411 ( .A1(n7077), .A2(n4286), .ZN(n4791) );
  AOI21_X1 U5412 ( .B1(n4583), .B2(n4579), .A(n4578), .ZN(n5198) );
  NAND2_X1 U5413 ( .A1(n4584), .A2(n4368), .ZN(n4583) );
  NAND2_X1 U5414 ( .A1(n8622), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n4781) );
  AOI21_X1 U5415 ( .B1(n4780), .B2(n4779), .A(n4369), .ZN(n4778) );
  INV_X1 U5416 ( .A(n9153), .ZN(n8928) );
  NAND2_X1 U5417 ( .A1(n9157), .A2(n9003), .ZN(n8931) );
  OR2_X1 U5418 ( .A1(n4269), .A2(n7396), .ZN(n8996) );
  NAND2_X1 U5419 ( .A1(n4671), .A2(n4471), .ZN(n6735) );
  AND2_X1 U5420 ( .A1(n4670), .A2(n4673), .ZN(n4471) );
  NAND2_X1 U5421 ( .A1(n4672), .A2(n8999), .ZN(n4671) );
  INV_X1 U5422 ( .A(n6726), .ZN(n8089) );
  NAND2_X1 U5423 ( .A1(n6640), .A2(n6639), .ZN(n9159) );
  INV_X1 U5424 ( .A(n8361), .ZN(n9241) );
  NAND2_X1 U5425 ( .A1(n7288), .A2(n6555), .ZN(n4497) );
  NAND2_X1 U5426 ( .A1(n4394), .A2(n4393), .ZN(n4392) );
  NAND2_X1 U5427 ( .A1(n6076), .A2(n6555), .ZN(n6079) );
  AND3_X1 U5428 ( .A1(n6269), .A2(n6268), .A3(n6267), .ZN(n9453) );
  AND2_X1 U5429 ( .A1(n6440), .A2(n6415), .ZN(n9632) );
  AOI21_X1 U5430 ( .B1(n4410), .B2(n8004), .A(n4408), .ZN(n7885) );
  NAND2_X1 U5431 ( .A1(n4862), .A2(n7984), .ZN(n4861) );
  NAND2_X1 U5432 ( .A1(n6407), .A2(n6406), .ZN(n9657) );
  INV_X1 U5433 ( .A(n9709), .ZN(n9489) );
  INV_X1 U5434 ( .A(n9291), .ZN(n9491) );
  AND2_X1 U5435 ( .A1(n4422), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n4560) );
  AND2_X1 U5436 ( .A1(n4574), .A2(n4573), .ZN(n6932) );
  NAND2_X1 U5437 ( .A1(n6925), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n4573) );
  AND2_X1 U5438 ( .A1(n6936), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n4677) );
  NOR2_X1 U5439 ( .A1(n6947), .A2(n6946), .ZN(n6945) );
  NOR2_X1 U5440 ( .A1(n6765), .A2(n6766), .ZN(n6764) );
  NOR2_X1 U5441 ( .A1(n6753), .A2(n6754), .ZN(n6752) );
  OR2_X1 U5442 ( .A1(n9961), .A2(n9960), .ZN(n9963) );
  AND2_X1 U5443 ( .A1(n6832), .A2(n6827), .ZN(n9964) );
  NAND2_X1 U5444 ( .A1(n4567), .A2(n4565), .ZN(n9956) );
  NAND2_X1 U5445 ( .A1(n4567), .A2(n6583), .ZN(n9954) );
  NAND2_X1 U5446 ( .A1(n6607), .A2(n6606), .ZN(n9970) );
  NAND2_X1 U5447 ( .A1(n9594), .A2(n9593), .ZN(n9790) );
  AND2_X1 U5448 ( .A1(n9592), .A2(n4982), .ZN(n9593) );
  NAND2_X1 U5449 ( .A1(n4825), .A2(n4829), .ZN(n9584) );
  OR2_X1 U5450 ( .A1(n9622), .A2(n4830), .ZN(n4825) );
  OAI21_X1 U5451 ( .B1(n9611), .B2(n9610), .A(n9609), .ZN(n9794) );
  NOR2_X1 U5452 ( .A1(n9605), .A2(n9604), .ZN(n9610) );
  NOR2_X1 U5453 ( .A1(n9799), .A2(n4406), .ZN(n9633) );
  NOR2_X1 U5454 ( .A1(n4407), .A2(n10068), .ZN(n4406) );
  INV_X1 U5455 ( .A(n9632), .ZN(n4407) );
  OAI21_X1 U5456 ( .B1(n7945), .B2(n10139), .A(n7777), .ZN(n6614) );
  NAND2_X1 U5457 ( .A1(n4727), .A2(n9787), .ZN(n9863) );
  AOI21_X1 U5458 ( .B1(n9783), .B2(n10136), .A(n4334), .ZN(n4727) );
  NAND2_X1 U5459 ( .A1(n8085), .A2(n9858), .ZN(n9785) );
  INV_X1 U5460 ( .A(n8293), .ZN(n8294) );
  NAND2_X1 U5461 ( .A1(n8301), .A2(n8440), .ZN(n4915) );
  AOI21_X1 U5462 ( .B1(n4917), .B2(n4916), .A(n4914), .ZN(n4913) );
  NOR2_X1 U5463 ( .A1(n8301), .A2(n8440), .ZN(n4916) );
  NAND2_X1 U5464 ( .A1(n8486), .A2(n4915), .ZN(n4914) );
  NAND2_X1 U5465 ( .A1(n8300), .A2(n8299), .ZN(n4917) );
  OR2_X1 U5466 ( .A1(n7796), .A2(n7795), .ZN(n7800) );
  OAI21_X1 U5467 ( .B1(n8319), .B2(n4328), .A(n4909), .ZN(n4911) );
  AOI21_X1 U5468 ( .B1(n4944), .B2(n8317), .A(n4910), .ZN(n4909) );
  INV_X1 U5469 ( .A(n8330), .ZN(n8332) );
  NAND2_X1 U5470 ( .A1(n4482), .A2(n4481), .ZN(n7836) );
  NAND2_X1 U5471 ( .A1(n7829), .A2(n7877), .ZN(n4481) );
  NOR2_X1 U5472 ( .A1(n8351), .A2(n8352), .ZN(n4401) );
  NOR2_X1 U5473 ( .A1(n8809), .A2(n8366), .ZN(n4932) );
  NAND2_X1 U5474 ( .A1(n4926), .A2(n4318), .ZN(n4925) );
  NAND2_X1 U5475 ( .A1(n8823), .A2(n8359), .ZN(n4926) );
  NAND2_X1 U5476 ( .A1(n8389), .A2(n8440), .ZN(n4425) );
  AND2_X1 U5477 ( .A1(n7849), .A2(n7956), .ZN(n4443) );
  NOR2_X1 U5478 ( .A1(n4717), .A2(n4478), .ZN(n4477) );
  NAND2_X1 U5479 ( .A1(n7996), .A2(n7882), .ZN(n4478) );
  NAND2_X1 U5480 ( .A1(n4376), .A2(n4304), .ZN(n8395) );
  INV_X1 U5481 ( .A(n4376), .ZN(n8394) );
  INV_X1 U5482 ( .A(n8800), .ZN(n4452) );
  INV_X1 U5483 ( .A(n7888), .ZN(n4473) );
  INV_X1 U5484 ( .A(n5637), .ZN(n5643) );
  INV_X1 U5485 ( .A(n5551), .ZN(n5556) );
  INV_X1 U5486 ( .A(n7281), .ZN(n4614) );
  AND2_X1 U5487 ( .A1(n5613), .A2(n5630), .ZN(n4526) );
  INV_X1 U5488 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n4987) );
  NOR2_X2 U5489 ( .A1(P2_IR_REG_14__SCAN_IN), .A2(P2_IR_REG_13__SCAN_IN), .ZN(
        n5028) );
  NAND2_X1 U5490 ( .A1(n6478), .A2(n7985), .ZN(n5902) );
  OAI21_X1 U5491 ( .B1(n4866), .B2(n7898), .A(n4865), .ZN(n4435) );
  NAND2_X1 U5492 ( .A1(n7898), .A2(n7882), .ZN(n4865) );
  NOR2_X1 U5493 ( .A1(n7953), .A2(n4296), .ZN(n4867) );
  INV_X1 U5494 ( .A(n7905), .ZN(n4712) );
  NAND2_X1 U5495 ( .A1(n10011), .A2(n10092), .ZN(n7906) );
  OR2_X1 U5496 ( .A1(n5991), .A2(n5914), .ZN(n5916) );
  NOR2_X1 U5497 ( .A1(n4887), .A2(n4882), .ZN(n4881) );
  INV_X1 U5498 ( .A(n5297), .ZN(n4882) );
  NAND2_X1 U5499 ( .A1(n4889), .A2(n4888), .ZN(n4887) );
  INV_X1 U5500 ( .A(n5646), .ZN(n4888) );
  NOR2_X1 U5501 ( .A1(n4891), .A2(n5646), .ZN(n4886) );
  NAND2_X1 U5502 ( .A1(n5556), .A2(n5287), .ZN(n4545) );
  INV_X1 U5503 ( .A(n4545), .ZN(n4543) );
  INV_X1 U5504 ( .A(n4553), .ZN(n4552) );
  OAI21_X1 U5505 ( .B1(n4294), .B2(n4554), .A(n4276), .ZN(n4553) );
  INV_X1 U5506 ( .A(n5493), .ZN(n4550) );
  INV_X1 U5507 ( .A(n5445), .ZN(n4771) );
  INV_X1 U5508 ( .A(n5483), .ZN(n4774) );
  INV_X1 U5509 ( .A(n4547), .ZN(n5598) );
  AND2_X1 U5510 ( .A1(n4534), .A2(n8175), .ZN(n4533) );
  NAND2_X1 U5511 ( .A1(n5709), .A2(n5703), .ZN(n4534) );
  INV_X1 U5512 ( .A(n8428), .ZN(n4907) );
  NOR2_X1 U5513 ( .A1(n8426), .A2(n8427), .ZN(n4906) );
  AND2_X1 U5514 ( .A1(n8497), .A2(n4449), .ZN(n8498) );
  NAND2_X1 U5515 ( .A1(n5055), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n4617) );
  INV_X1 U5516 ( .A(n4795), .ZN(n4793) );
  AND2_X1 U5517 ( .A1(n5100), .A2(n4607), .ZN(n4604) );
  NAND2_X1 U5518 ( .A1(n8638), .A2(n5108), .ZN(n4591) );
  AND2_X1 U5519 ( .A1(n4526), .A2(n4525), .ZN(n4524) );
  INV_X1 U5520 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n4525) );
  NOR2_X1 U5521 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(P2_REG3_REG_12__SCAN_IN), 
        .ZN(n4519) );
  AOI21_X1 U5522 ( .B1(n4632), .B2(n4629), .A(n4295), .ZN(n4628) );
  OR2_X1 U5523 ( .A1(n4630), .A2(n4627), .ZN(n4354) );
  INV_X1 U5524 ( .A(n4635), .ZN(n4629) );
  NAND2_X1 U5525 ( .A1(n6621), .A2(n7171), .ZN(n6652) );
  XNOR2_X1 U5526 ( .A(n8538), .B(n10164), .ZN(n8302) );
  NAND2_X1 U5527 ( .A1(n4651), .A2(n4655), .ZN(n4649) );
  NAND2_X1 U5528 ( .A1(n4653), .A2(n6684), .ZN(n8667) );
  NAND2_X1 U5529 ( .A1(n4657), .A2(n4654), .ZN(n4653) );
  AND2_X1 U5530 ( .A1(n9185), .A2(n8702), .ZN(n8471) );
  AND2_X1 U5531 ( .A1(n6673), .A2(n4641), .ZN(n4640) );
  NAND2_X1 U5532 ( .A1(n4642), .A2(n6670), .ZN(n4641) );
  INV_X1 U5533 ( .A(n4644), .ZN(n4642) );
  INV_X1 U5534 ( .A(n6672), .ZN(n8386) );
  AND2_X1 U5535 ( .A1(n8364), .A2(n4667), .ZN(n4661) );
  OR2_X1 U5536 ( .A1(n4295), .A2(n7192), .ZN(n8478) );
  NAND2_X1 U5537 ( .A1(n4634), .A2(n4631), .ZN(n7193) );
  INV_X1 U5538 ( .A(n4633), .ZN(n4631) );
  NAND2_X1 U5539 ( .A1(n7176), .A2(n4635), .ZN(n4634) );
  INV_X1 U5540 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n4737) );
  AND2_X1 U5541 ( .A1(n6738), .A2(n6996), .ZN(n5905) );
  AND2_X1 U5542 ( .A1(n6391), .A2(n6390), .ZN(n6392) );
  INV_X1 U5543 ( .A(n10049), .ZN(n4427) );
  OR2_X1 U5544 ( .A1(n8015), .A2(n6478), .ZN(n6566) );
  AOI21_X1 U5545 ( .B1(n7999), .B2(n7899), .A(n7898), .ZN(n8000) );
  NAND2_X1 U5546 ( .A1(n6041), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n5974) );
  AND2_X1 U5547 ( .A1(n4569), .A2(n4568), .ZN(n6580) );
  NAND2_X1 U5548 ( .A1(n9908), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n4568) );
  INV_X1 U5549 ( .A(n9940), .ZN(n4563) );
  INV_X1 U5550 ( .A(n6584), .ZN(n4562) );
  NAND2_X1 U5551 ( .A1(n9599), .A2(n9488), .ZN(n8048) );
  NAND2_X1 U5552 ( .A1(n9626), .A2(n9650), .ZN(n4901) );
  NAND2_X1 U5553 ( .A1(n4844), .A2(n8071), .ZN(n4843) );
  NAND2_X1 U5554 ( .A1(n4845), .A2(n4846), .ZN(n4844) );
  INV_X1 U5555 ( .A(n4732), .ZN(n4731) );
  NOR2_X1 U5556 ( .A1(n6359), .A2(n6358), .ZN(n4413) );
  OR2_X1 U5557 ( .A1(n9814), .A2(n8067), .ZN(n7858) );
  NOR2_X1 U5558 ( .A1(n9824), .A2(n9829), .ZN(n4897) );
  INV_X1 U5559 ( .A(n4486), .ZN(n4723) );
  OAI21_X1 U5560 ( .B1(n9727), .B2(n7996), .A(n7997), .ZN(n4486) );
  OR2_X1 U5561 ( .A1(n9843), .A2(n9453), .ZN(n7994) );
  NOR2_X1 U5562 ( .A1(n7970), .A2(n4715), .ZN(n4713) );
  INV_X1 U5563 ( .A(n6062), .ZN(n5874) );
  NAND2_X1 U5564 ( .A1(n5873), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n6062) );
  INV_X1 U5565 ( .A(n6039), .ZN(n5873) );
  NAND2_X1 U5566 ( .A1(n7372), .A2(n4985), .ZN(n7908) );
  NOR2_X1 U5567 ( .A1(n7903), .A2(n10058), .ZN(n7641) );
  NAND2_X1 U5568 ( .A1(n9628), .A2(n9629), .ZN(n4511) );
  NAND2_X1 U5569 ( .A1(n9638), .A2(n8045), .ZN(n9628) );
  NAND3_X1 U5570 ( .A1(n9679), .A2(n9729), .A3(n4277), .ZN(n9674) );
  INV_X1 U5571 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5836) );
  AND2_X1 U5572 ( .A1(n6518), .A2(n4363), .ZN(n6525) );
  OR2_X1 U5573 ( .A1(n6516), .A2(n6515), .ZN(n6517) );
  AND2_X1 U5574 ( .A1(n6511), .A2(n5718), .ZN(n5732) );
  NAND2_X1 U5575 ( .A1(n5667), .A2(n5651), .ZN(n5668) );
  NAND2_X1 U5576 ( .A1(n5585), .A2(n4891), .ZN(n4883) );
  NAND2_X1 U5577 ( .A1(n5606), .A2(n5306), .ZN(n5607) );
  INV_X1 U5578 ( .A(n5584), .ZN(n5302) );
  XNOR2_X1 U5579 ( .A(n5299), .B(SI_18_), .ZN(n5584) );
  AOI21_X1 U5580 ( .B1(n4876), .B2(n4878), .A(n4874), .ZN(n4873) );
  INV_X1 U5581 ( .A(n4877), .ZN(n4876) );
  NAND2_X1 U5582 ( .A1(n5297), .A2(n5296), .ZN(n5570) );
  INV_X1 U5583 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n4705) );
  NAND2_X1 U5584 ( .A1(n5559), .A2(n4287), .ZN(n4544) );
  NOR2_X1 U5585 ( .A1(n5559), .A2(n4543), .ZN(n4542) );
  OAI21_X1 U5586 ( .B1(n5559), .B2(n4287), .A(n4545), .ZN(n4539) );
  NAND2_X1 U5587 ( .A1(n4541), .A2(n4543), .ZN(n4540) );
  INV_X1 U5588 ( .A(n5559), .ZN(n4541) );
  NAND2_X1 U5589 ( .A1(n5281), .A2(SI_12_), .ZN(n5511) );
  NAND2_X1 U5590 ( .A1(n5473), .A2(n5279), .ZN(n5494) );
  NAND2_X1 U5591 ( .A1(n5251), .A2(n5250), .ZN(n5327) );
  OAI211_X1 U5592 ( .C1(n4494), .C2(P1_DATAO_REG_2__SCAN_IN), .A(n4491), .B(
        n4490), .ZN(n5231) );
  NAND2_X1 U5593 ( .A1(n4492), .A2(n4496), .ZN(n4491) );
  AOI21_X1 U5594 ( .B1(n5527), .B2(n4307), .A(n4279), .ZN(n4748) );
  INV_X1 U5595 ( .A(n5527), .ZN(n4749) );
  OR2_X1 U5596 ( .A1(n7137), .A2(n7139), .ZN(n4756) );
  NAND2_X1 U5597 ( .A1(n4529), .A2(n4324), .ZN(n4758) );
  NAND2_X1 U5598 ( .A1(n5604), .A2(n4761), .ZN(n4529) );
  XNOR2_X1 U5599 ( .A(n5442), .B(n10164), .ZN(n5378) );
  NAND2_X1 U5600 ( .A1(n4547), .A2(n4546), .ZN(n8261) );
  AOI21_X1 U5601 ( .B1(n5597), .B2(n8183), .A(n5599), .ZN(n4546) );
  NAND2_X1 U5602 ( .A1(n4751), .A2(n7231), .ZN(n4753) );
  AOI21_X1 U5603 ( .B1(n4750), .B2(n4278), .A(n7232), .ZN(n4754) );
  INV_X1 U5604 ( .A(n4755), .ZN(n4751) );
  AND2_X1 U5605 ( .A1(n8462), .A2(n8461), .ZN(n8648) );
  AND2_X1 U5606 ( .A1(n8462), .A2(n6650), .ZN(n8531) );
  NAND2_X1 U5607 ( .A1(n4455), .A2(n4454), .ZN(n6855) );
  NAND2_X1 U5608 ( .A1(n6851), .A2(n5113), .ZN(n4454) );
  OR2_X1 U5609 ( .A1(n6851), .A2(n5113), .ZN(n4455) );
  OAI21_X1 U5610 ( .B1(n7067), .B2(n4595), .A(n4592), .ZN(n7036) );
  INV_X1 U5611 ( .A(n7033), .ZN(n4595) );
  AND2_X1 U5612 ( .A1(n7032), .A2(n4593), .ZN(n4592) );
  NAND2_X1 U5613 ( .A1(n7067), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n7066) );
  NOR3_X1 U5614 ( .A1(n7062), .A2(n7025), .A3(n7024), .ZN(n7023) );
  NOR2_X1 U5615 ( .A1(n7028), .A2(n4316), .ZN(n5124) );
  NAND2_X1 U5616 ( .A1(n4616), .A2(n6891), .ZN(n6986) );
  INV_X1 U5617 ( .A(n4617), .ZN(n4616) );
  AOI21_X1 U5618 ( .B1(n7275), .B2(n7274), .A(n7273), .ZN(n7480) );
  OAI21_X1 U5619 ( .B1(n7480), .B2(n7479), .A(n7478), .ZN(n7524) );
  INV_X1 U5620 ( .A(n4609), .ZN(n4608) );
  INV_X1 U5621 ( .A(n4784), .ZN(n4783) );
  INV_X1 U5622 ( .A(n4788), .ZN(n4787) );
  OAI21_X1 U5623 ( .B1(n8547), .B2(n8546), .A(n8545), .ZN(n8560) );
  NAND2_X1 U5624 ( .A1(n4799), .A2(n8544), .ZN(n4806) );
  INV_X1 U5625 ( .A(n8566), .ZN(n4601) );
  AOI21_X1 U5626 ( .B1(n8560), .B2(n8559), .A(n8558), .ZN(n8579) );
  OAI211_X1 U5627 ( .C1(n8540), .C2(n4802), .A(n4805), .B(n4800), .ZN(n4804)
         );
  NAND2_X1 U5628 ( .A1(n8557), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n4805) );
  NAND2_X1 U5629 ( .A1(n8555), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n4802) );
  NAND2_X1 U5630 ( .A1(n4801), .A2(n8555), .ZN(n4800) );
  OAI21_X1 U5631 ( .B1(n8579), .B2(n8578), .A(n8577), .ZN(n8592) );
  OAI21_X1 U5632 ( .B1(n8608), .B2(n8607), .A(n8606), .ZN(n8610) );
  INV_X1 U5633 ( .A(n4589), .ZN(n4582) );
  NAND2_X1 U5634 ( .A1(n4588), .A2(n5186), .ZN(n4587) );
  INV_X1 U5635 ( .A(n4591), .ZN(n4588) );
  INV_X1 U5636 ( .A(n4282), .ZN(n4584) );
  AND2_X1 U5637 ( .A1(n8622), .A2(n8614), .ZN(n4779) );
  AND2_X1 U5638 ( .A1(n8500), .A2(n8466), .ZN(n6699) );
  NAND2_X1 U5639 ( .A1(n5763), .A2(n5762), .ZN(n5797) );
  INV_X1 U5640 ( .A(n5764), .ZN(n5763) );
  NAND2_X1 U5641 ( .A1(n5684), .A2(n5683), .ZN(n5723) );
  INV_X1 U5642 ( .A(n5693), .ZN(n5684) );
  NAND2_X1 U5643 ( .A1(n5614), .A2(n4524), .ZN(n5691) );
  NAND2_X1 U5644 ( .A1(n4516), .A2(n5206), .ZN(n5590) );
  INV_X1 U5645 ( .A(n4516), .ZN(n5575) );
  NAND2_X1 U5646 ( .A1(n5205), .A2(n5204), .ZN(n5565) );
  INV_X1 U5647 ( .A(n5545), .ZN(n5205) );
  NAND2_X1 U5648 ( .A1(n5203), .A2(n4517), .ZN(n5545) );
  AND2_X1 U5649 ( .A1(n4519), .A2(n4518), .ZN(n4517) );
  INV_X1 U5650 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n4518) );
  NAND2_X1 U5651 ( .A1(n5203), .A2(n4519), .ZN(n5535) );
  AND2_X1 U5652 ( .A1(n8327), .A2(n8902), .ZN(n8879) );
  INV_X1 U5653 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5202) );
  NAND2_X1 U5654 ( .A1(n5201), .A2(n4290), .ZN(n5463) );
  CLKBUF_X1 U5655 ( .A(n7384), .Z(n7385) );
  NAND2_X1 U5656 ( .A1(n5201), .A2(n5200), .ZN(n5446) );
  INV_X1 U5657 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5199) );
  NAND2_X1 U5658 ( .A1(n7142), .A2(n4521), .ZN(n5401) );
  NAND2_X1 U5659 ( .A1(n4625), .A2(n6652), .ZN(n7176) );
  INV_X1 U5660 ( .A(n4626), .ZN(n4625) );
  OR2_X1 U5661 ( .A1(n7011), .A2(n7010), .ZN(n7017) );
  AND2_X1 U5662 ( .A1(n7007), .A2(n5772), .ZN(n6713) );
  INV_X1 U5663 ( .A(n4962), .ZN(n4960) );
  AOI21_X1 U5664 ( .B1(n4962), .B2(n4959), .A(n4958), .ZN(n4957) );
  NOR2_X1 U5665 ( .A1(n4964), .A2(n8413), .ZN(n4962) );
  NOR2_X1 U5666 ( .A1(n8472), .A2(n8471), .ZN(n8717) );
  NAND2_X1 U5667 ( .A1(n6672), .A2(n8400), .ZN(n8744) );
  OR2_X1 U5668 ( .A1(n4947), .A2(n6636), .ZN(n4946) );
  INV_X1 U5669 ( .A(n4274), .ZN(n6701) );
  NAND2_X1 U5670 ( .A1(n6669), .A2(n4644), .ZN(n4639) );
  AND2_X1 U5671 ( .A1(n5621), .A2(n5620), .ZN(n8769) );
  AND2_X1 U5672 ( .A1(n8371), .A2(n8374), .ZN(n8800) );
  NAND2_X1 U5673 ( .A1(n8843), .A2(n8356), .ZN(n8836) );
  OR2_X1 U5674 ( .A1(n6720), .A2(n8463), .ZN(n7012) );
  OR3_X1 U5675 ( .A1(n4274), .A2(n7542), .A3(n8510), .ZN(n6728) );
  INV_X1 U5676 ( .A(n6866), .ZN(n5359) );
  NAND2_X1 U5677 ( .A1(n5794), .A2(n9287), .ZN(n4935) );
  AND2_X1 U5678 ( .A1(n4971), .A2(n5020), .ZN(n4970) );
  AND2_X1 U5679 ( .A1(n4998), .A2(n4997), .ZN(n5316) );
  AND2_X1 U5680 ( .A1(n5097), .A2(n5095), .ZN(n5532) );
  OR2_X1 U5681 ( .A1(n5063), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n5070) );
  XNOR2_X1 U5682 ( .A(n5057), .B(P2_IR_REG_6__SCAN_IN), .ZN(n6804) );
  INV_X1 U5683 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5048) );
  NAND2_X1 U5684 ( .A1(n5034), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4458) );
  AND2_X1 U5685 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n4811) );
  NAND2_X1 U5686 ( .A1(n4938), .A2(n5023), .ZN(n4618) );
  INV_X1 U5687 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n6234) );
  INV_X1 U5688 ( .A(n5931), .ZN(n9334) );
  INV_X1 U5689 ( .A(n4423), .ZN(n6421) );
  AND2_X1 U5690 ( .A1(n6272), .A2(n6271), .ZN(n9383) );
  AND2_X1 U5691 ( .A1(n6376), .A2(n6375), .ZN(n7760) );
  NAND2_X1 U5692 ( .A1(n7753), .A2(n4693), .ZN(n4692) );
  XNOR2_X1 U5693 ( .A(n5459), .B(n5458), .ZN(n6076) );
  NAND2_X1 U5694 ( .A1(n4412), .A2(n4314), .ZN(n6169) );
  INV_X1 U5695 ( .A(n6145), .ZN(n4412) );
  NAND2_X1 U5696 ( .A1(n4466), .A2(n4465), .ZN(n6237) );
  NOR2_X1 U5697 ( .A1(n6235), .A2(n6234), .ZN(n4465) );
  INV_X1 U5698 ( .A(n6236), .ZN(n4466) );
  NAND2_X1 U5699 ( .A1(n4464), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n6221) );
  INV_X1 U5700 ( .A(n6237), .ZN(n4464) );
  OR2_X1 U5701 ( .A1(n6494), .A2(n6492), .ZN(n6502) );
  NAND2_X1 U5702 ( .A1(n7945), .A2(n7882), .ZN(n4409) );
  INV_X1 U5703 ( .A(n7883), .ZN(n4410) );
  AND3_X1 U5704 ( .A1(n6209), .A2(n6208), .A3(n6207), .ZN(n9476) );
  NAND2_X1 U5705 ( .A1(n6323), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5996) );
  OAI21_X1 U5706 ( .B1(n4422), .B2(n5993), .A(n4428), .ZN(n9547) );
  NAND2_X1 U5707 ( .A1(n9552), .A2(n5993), .ZN(n4428) );
  AND2_X1 U5708 ( .A1(n9548), .A2(n9547), .ZN(n9550) );
  NOR2_X1 U5709 ( .A1(n6768), .A2(n6769), .ZN(n6767) );
  AND2_X1 U5710 ( .A1(n6745), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n4572) );
  XNOR2_X1 U5711 ( .A(n7107), .B(n6580), .ZN(n9914) );
  NOR2_X1 U5712 ( .A1(n4418), .A2(n7721), .ZN(n4448) );
  NAND2_X1 U5713 ( .A1(n4418), .A2(n4417), .ZN(n4416) );
  INV_X1 U5714 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n4417) );
  AND2_X1 U5715 ( .A1(n4566), .A2(n6583), .ZN(n4565) );
  INV_X1 U5716 ( .A(n9953), .ZN(n4566) );
  NAND2_X1 U5717 ( .A1(n9939), .A2(n9940), .ZN(n4567) );
  NAND2_X1 U5718 ( .A1(n9595), .A2(n9784), .ZN(n8082) );
  NOR2_X1 U5719 ( .A1(n8082), .A2(n8004), .ZN(n6611) );
  INV_X1 U5720 ( .A(n8077), .ZN(n8049) );
  NAND2_X1 U5721 ( .A1(n9488), .A2(n10010), .ZN(n8053) );
  NAND2_X1 U5722 ( .A1(n4832), .A2(n4289), .ZN(n4829) );
  NAND2_X1 U5723 ( .A1(n4833), .A2(n4284), .ZN(n4832) );
  INV_X1 U5724 ( .A(n9604), .ZN(n4833) );
  NAND2_X1 U5725 ( .A1(n4289), .A2(n4831), .ZN(n4830) );
  INV_X1 U5726 ( .A(n8075), .ZN(n4831) );
  INV_X1 U5727 ( .A(n8046), .ZN(n4733) );
  NOR2_X1 U5728 ( .A1(n9660), .A2(n9804), .ZN(n9645) );
  XNOR2_X1 U5729 ( .A(n9800), .B(n8074), .ZN(n9629) );
  INV_X1 U5730 ( .A(n4413), .ZN(n6380) );
  AND2_X1 U5731 ( .A1(n6387), .A2(n6386), .ZN(n9673) );
  NAND2_X1 U5732 ( .A1(n9729), .A2(n9724), .ZN(n9718) );
  NAND2_X1 U5733 ( .A1(n9729), .A2(n4897), .ZN(n9699) );
  OR2_X1 U5734 ( .A1(n6321), .A2(n6320), .ZN(n6341) );
  OAI21_X1 U5735 ( .B1(n4404), .B2(n9727), .A(n4723), .ZN(n9715) );
  INV_X1 U5736 ( .A(n9834), .ZN(n9731) );
  NOR2_X2 U5737 ( .A1(n4895), .A2(n7834), .ZN(n9744) );
  AND2_X1 U5738 ( .A1(n7994), .A2(n7957), .ZN(n9769) );
  NAND2_X1 U5739 ( .A1(n7691), .A2(n4894), .ZN(n9761) );
  NAND2_X1 U5740 ( .A1(n4335), .A2(n4860), .ZN(n4857) );
  NAND2_X1 U5741 ( .A1(n7691), .A2(n9486), .ZN(n7719) );
  NAND2_X1 U5742 ( .A1(n9430), .A2(n7700), .ZN(n7924) );
  NAND2_X1 U5743 ( .A1(n7461), .A2(n9494), .ZN(n7827) );
  NAND2_X1 U5744 ( .A1(n9984), .A2(n4317), .ZN(n7617) );
  AND2_X1 U5745 ( .A1(n7464), .A2(n7822), .ZN(n7465) );
  OR2_X1 U5746 ( .A1(n7463), .A2(n7823), .ZN(n7464) );
  CLKBUF_X1 U5747 ( .A(n7624), .Z(n7623) );
  AOI21_X1 U5748 ( .B1(n7965), .B2(n4839), .A(n4837), .ZN(n4836) );
  AND2_X1 U5749 ( .A1(n7827), .A2(n7923), .ZN(n4983) );
  NAND2_X1 U5750 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n6014) );
  NAND2_X1 U5751 ( .A1(n5872), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n6039) );
  INV_X1 U5752 ( .A(n6014), .ZN(n5872) );
  NAND2_X1 U5753 ( .A1(n7583), .A2(n7373), .ZN(n7584) );
  CLKBUF_X1 U5754 ( .A(n7488), .Z(n10021) );
  AND2_X1 U5755 ( .A1(n10086), .A2(n7641), .ZN(n10038) );
  INV_X1 U5756 ( .A(n7949), .ZN(n7000) );
  NAND2_X1 U5757 ( .A1(n4509), .A2(n4507), .ZN(n9799) );
  INV_X1 U5758 ( .A(n4508), .ZN(n4507) );
  NAND2_X1 U5759 ( .A1(n4510), .A2(n10013), .ZN(n4509) );
  OAI22_X1 U5760 ( .A1(n9631), .A2(n10048), .B1(n10050), .B2(n9630), .ZN(n4508) );
  AND2_X1 U5761 ( .A1(n9800), .A2(n9858), .ZN(n4505) );
  NAND2_X1 U5762 ( .A1(n4872), .A2(n6378), .ZN(n9809) );
  NAND2_X1 U5763 ( .A1(n7669), .A2(n6555), .ZN(n4872) );
  INV_X1 U5764 ( .A(n9445), .ZN(n7456) );
  AND2_X1 U5765 ( .A1(n6459), .A2(n7728), .ZN(n6817) );
  XNOR2_X1 U5766 ( .A(n6525), .B(n6524), .ZN(n9278) );
  NAND2_X1 U5767 ( .A1(n5753), .A2(n6510), .ZN(n5759) );
  NOR2_X1 U5768 ( .A1(n4388), .A2(n4387), .ZN(n4386) );
  OR2_X1 U5769 ( .A1(n5859), .A2(n4390), .ZN(n4389) );
  NOR2_X1 U5770 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n4387) );
  NAND2_X1 U5771 ( .A1(n5861), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5864) );
  NAND2_X1 U5772 ( .A1(n5864), .A2(n5863), .ZN(n5866) );
  OAI21_X2 U5773 ( .B1(n6201), .B2(P1_IR_REG_17__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5894) );
  INV_X1 U5774 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n6216) );
  INV_X1 U5775 ( .A(n4501), .ZN(n4500) );
  NOR2_X1 U5776 ( .A1(n5493), .A2(n4502), .ZN(n4501) );
  OAI21_X1 U5777 ( .B1(n5277), .B2(SI_10_), .A(n5279), .ZN(n5470) );
  NAND2_X1 U5778 ( .A1(n4871), .A2(n4870), .ZN(n5473) );
  CLKBUF_X1 U5779 ( .A(n6076), .Z(n6815) );
  NAND2_X1 U5780 ( .A1(n6031), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6007) );
  NAND2_X1 U5781 ( .A1(n5257), .A2(SI_3_), .ZN(n5392) );
  NAND2_X1 U5782 ( .A1(n5259), .A2(n5243), .ZN(n5395) );
  INV_X1 U5783 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5970) );
  NAND2_X1 U5784 ( .A1(n5969), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5949) );
  NAND2_X1 U5786 ( .A1(n4775), .A2(n5443), .ZN(n7449) );
  INV_X1 U5787 ( .A(n7451), .ZN(n4775) );
  NAND2_X1 U5788 ( .A1(n5751), .A2(n5750), .ZN(n4528) );
  AND4_X1 U5789 ( .A1(n5492), .A2(n5491), .A3(n5490), .A4(n5489), .ZN(n8846)
         );
  NAND2_X1 U5790 ( .A1(n4763), .A2(n5603), .ZN(n8123) );
  NAND2_X1 U5791 ( .A1(n4763), .A2(n4761), .ZN(n8124) );
  INV_X1 U5792 ( .A(n8699), .ZN(n8178) );
  INV_X1 U5793 ( .A(n4532), .ZN(n8174) );
  NAND2_X1 U5794 ( .A1(n4756), .A2(n4755), .ZN(n7233) );
  AND2_X1 U5795 ( .A1(n5636), .A2(n5635), .ZN(n8253) );
  NAND2_X1 U5796 ( .A1(n4759), .A2(n4760), .ZN(n8228) );
  INV_X1 U5797 ( .A(n4758), .ZN(n4760) );
  AND4_X1 U5798 ( .A1(n5509), .A2(n5508), .A3(n5507), .A4(n5506), .ZN(n8355)
         );
  OR2_X1 U5799 ( .A1(n8113), .A2(n8345), .ZN(n5485) );
  OAI21_X1 U5800 ( .B1(n7451), .B2(n4768), .A(n4766), .ZN(n5486) );
  INV_X1 U5801 ( .A(n4769), .ZN(n4768) );
  INV_X1 U5802 ( .A(n8283), .ZN(n8266) );
  XNOR2_X1 U5803 ( .A(n5013), .B(P2_IR_REG_22__SCAN_IN), .ZN(n8525) );
  NAND2_X1 U5804 ( .A1(n5698), .A2(n5697), .ZN(n8734) );
  INV_X1 U5805 ( .A(n8253), .ZN(n8758) );
  INV_X1 U5806 ( .A(n8355), .ZN(n8829) );
  OAI22_X1 U5807 ( .A1(n6850), .A2(n6849), .B1(n5138), .B2(n5137), .ZN(n7063)
         );
  XNOR2_X1 U5808 ( .A(n5120), .B(n5119), .ZN(n7065) );
  XNOR2_X1 U5809 ( .A(n5124), .B(n5052), .ZN(n6985) );
  AND2_X1 U5810 ( .A1(n4621), .A2(n7088), .ZN(n7054) );
  NAND2_X1 U5811 ( .A1(n7203), .A2(n7280), .ZN(n4611) );
  AND2_X1 U5812 ( .A1(n4790), .A2(n4797), .ZN(n7270) );
  NAND2_X1 U5813 ( .A1(n4789), .A2(n4796), .ZN(n4797) );
  XNOR2_X1 U5814 ( .A(n4804), .B(n8576), .ZN(n8572) );
  NAND2_X1 U5815 ( .A1(n8599), .A2(n8597), .ZN(n4602) );
  OR2_X1 U5816 ( .A1(n8637), .A2(n8635), .ZN(n4445) );
  NAND2_X1 U5817 ( .A1(n4780), .A2(n8614), .ZN(n4782) );
  AOI21_X1 U5818 ( .B1(n8640), .B2(n8639), .A(n8638), .ZN(n8643) );
  INV_X1 U5819 ( .A(n6711), .ZN(n4673) );
  NAND2_X1 U5820 ( .A1(n5764), .A2(n5742), .ZN(n8693) );
  NAND2_X1 U5821 ( .A1(n6669), .A2(n6668), .ZN(n8776) );
  NAND2_X1 U5822 ( .A1(n4952), .A2(n4955), .ZN(n8780) );
  NAND2_X1 U5823 ( .A1(n4470), .A2(n4956), .ZN(n4952) );
  NAND2_X1 U5824 ( .A1(n8993), .A2(n5790), .ZN(n10165) );
  INV_X1 U5825 ( .A(n8784), .ZN(n8921) );
  INV_X1 U5826 ( .A(n10165), .ZN(n8920) );
  NAND2_X2 U5827 ( .A1(n7017), .A2(n10165), .ZN(n10171) );
  INV_X1 U5828 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n4513) );
  AND2_X1 U5829 ( .A1(n5682), .A2(n5681), .ZN(n8945) );
  INV_X1 U5830 ( .A(n8996), .ZN(n8979) );
  INV_X1 U5831 ( .A(n8507), .ZN(n9152) );
  NAND2_X1 U5832 ( .A1(n8437), .A2(n8436), .ZN(n9153) );
  AOI21_X1 U5833 ( .B1(n8660), .B2(n8887), .A(n8659), .ZN(n9157) );
  NAND2_X1 U5834 ( .A1(n8658), .A2(n8657), .ZN(n8659) );
  NAND2_X1 U5835 ( .A1(n8675), .A2(n8674), .ZN(n8676) );
  NAND2_X1 U5836 ( .A1(n8699), .A2(n8890), .ZN(n8674) );
  NAND2_X1 U5837 ( .A1(n4963), .A2(n4961), .ZN(n8666) );
  INV_X1 U5838 ( .A(n4964), .ZN(n4961) );
  NAND2_X1 U5839 ( .A1(n8706), .A2(n4965), .ZN(n4963) );
  INV_X1 U5840 ( .A(n6686), .ZN(n9171) );
  NAND2_X1 U5841 ( .A1(n8689), .A2(n8688), .ZN(n8690) );
  NAND2_X1 U5842 ( .A1(n8687), .A2(n8890), .ZN(n8688) );
  AOI21_X1 U5843 ( .B1(n8706), .B2(n8425), .A(n8410), .ZN(n8682) );
  INV_X1 U5844 ( .A(n8945), .ZN(n9185) );
  NAND2_X1 U5845 ( .A1(n5702), .A2(n5701), .ZN(n9191) );
  NAND2_X1 U5846 ( .A1(n6681), .A2(n6680), .ZN(n8722) );
  INV_X1 U5847 ( .A(n8259), .ZN(n9197) );
  AOI21_X1 U5848 ( .B1(n4951), .B2(n4470), .A(n4949), .ZN(n8765) );
  AOI21_X1 U5849 ( .B1(n4470), .B2(n8374), .A(n8377), .ZN(n8790) );
  NAND2_X1 U5850 ( .A1(n5562), .A2(n5561), .ZN(n9229) );
  NAND2_X1 U5851 ( .A1(n5555), .A2(n5554), .ZN(n9235) );
  NAND2_X1 U5852 ( .A1(n4666), .A2(n4665), .ZN(n8810) );
  NAND2_X1 U5853 ( .A1(n8828), .A2(n4667), .ZN(n4666) );
  AOI21_X1 U5854 ( .B1(n8828), .B2(n8476), .A(n8477), .ZN(n8817) );
  NAND2_X1 U5855 ( .A1(n5518), .A2(n5517), .ZN(n9248) );
  INV_X1 U5856 ( .A(n8340), .ZN(n8349) );
  INV_X1 U5857 ( .A(n9264), .ZN(n9247) );
  OR2_X1 U5858 ( .A1(n10188), .A2(n7396), .ZN(n9264) );
  NAND2_X1 U5859 ( .A1(n6796), .A2(n4744), .ZN(n6809) );
  BUF_X1 U5860 ( .A(n5215), .Z(n9269) );
  INV_X1 U5861 ( .A(n5316), .ZN(n7731) );
  NAND2_X1 U5862 ( .A1(n4776), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5002) );
  INV_X1 U5863 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n7613) );
  INV_X1 U5864 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7543) );
  INV_X1 U5865 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n9007) );
  XNOR2_X1 U5866 ( .A(n5311), .B(n5310), .ZN(n8503) );
  INV_X1 U5867 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n9118) );
  INV_X1 U5868 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n7145) );
  INV_X1 U5869 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n7158) );
  INV_X1 U5870 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n9108) );
  NAND2_X2 U5871 ( .A1(n5039), .A2(n5042), .ZN(n6851) );
  NAND2_X1 U5872 ( .A1(n4457), .A2(n4456), .ZN(n5039) );
  NAND2_X1 U5873 ( .A1(n5037), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4456) );
  NAND2_X1 U5874 ( .A1(n4458), .A2(P2_IR_REG_2__SCAN_IN), .ZN(n4457) );
  AND2_X1 U5875 ( .A1(n5893), .A2(n5892), .ZN(n9709) );
  NAND2_X1 U5876 ( .A1(n9308), .A2(n6152), .ZN(n4685) );
  AOI21_X1 U5877 ( .B1(n4691), .B2(n4694), .A(n9360), .ZN(n4689) );
  INV_X1 U5878 ( .A(n4691), .ZN(n4690) );
  NAND2_X1 U5879 ( .A1(n6204), .A2(n6203), .ZN(n9848) );
  NAND2_X1 U5880 ( .A1(n4702), .A2(n6259), .ZN(n9386) );
  NAND2_X1 U5881 ( .A1(n4692), .A2(n4695), .ZN(n7761) );
  NOR2_X1 U5882 ( .A1(n9393), .A2(n4687), .ZN(n4686) );
  INV_X1 U5883 ( .A(n5985), .ZN(n4687) );
  AND2_X1 U5884 ( .A1(n6305), .A2(n6304), .ZN(n9717) );
  AND2_X1 U5885 ( .A1(n4683), .A2(n6179), .ZN(n4682) );
  NAND2_X1 U5886 ( .A1(n5944), .A2(n5946), .ZN(n5947) );
  INV_X1 U5887 ( .A(n5945), .ZN(n5946) );
  INV_X1 U5888 ( .A(n9474), .ZN(n9458) );
  INV_X1 U5889 ( .A(n9451), .ZN(n9477) );
  INV_X1 U5890 ( .A(n9479), .ZN(n9468) );
  NOR2_X1 U5891 ( .A1(n6502), .A2(n6493), .ZN(n9474) );
  AND2_X1 U5892 ( .A1(n7251), .A2(n7250), .ZN(n9591) );
  NAND2_X1 U5893 ( .A1(n6420), .A2(n6419), .ZN(n9642) );
  INV_X1 U5894 ( .A(n9673), .ZN(n9641) );
  INV_X1 U5895 ( .A(n7504), .ZN(n9498) );
  NAND2_X1 U5896 ( .A1(n6041), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5957) );
  OR2_X1 U5897 ( .A1(n5992), .A2(n10043), .ZN(n5956) );
  OR2_X1 U5898 ( .A1(n5994), .A2(n5952), .ZN(n5955) );
  INV_X1 U5899 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n5229) );
  NAND2_X1 U5900 ( .A1(n6041), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5924) );
  OR2_X1 U5901 ( .A1(n5992), .A2(n10067), .ZN(n5926) );
  OR2_X1 U5902 ( .A1(n5994), .A2(n5921), .ZN(n5925) );
  OR2_X1 U5903 ( .A1(n6738), .A2(n6979), .ZN(n9501) );
  OAI21_X1 U5904 ( .B1(n9522), .B2(n5952), .A(n4414), .ZN(n9528) );
  NAND2_X1 U5905 ( .A1(n9522), .A2(n5952), .ZN(n4414) );
  OAI21_X1 U5906 ( .B1(n9522), .B2(n10148), .A(n4419), .ZN(n9525) );
  NAND2_X1 U5907 ( .A1(n9522), .A2(n10148), .ZN(n4419) );
  OAI21_X1 U5908 ( .B1(n9552), .B2(n10151), .A(n4395), .ZN(n9556) );
  NAND2_X1 U5909 ( .A1(n9552), .A2(n10151), .ZN(n4395) );
  NOR2_X1 U5910 ( .A1(n9553), .A2(n4674), .ZN(n6904) );
  AND2_X1 U5911 ( .A1(n4422), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n4674) );
  NOR2_X1 U5912 ( .A1(n6904), .A2(n6903), .ZN(n6902) );
  AND2_X1 U5913 ( .A1(n6908), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n4575) );
  INV_X1 U5914 ( .A(n4574), .ZN(n6922) );
  NOR2_X1 U5915 ( .A1(n6944), .A2(n6943), .ZN(n6942) );
  NOR2_X1 U5916 ( .A1(n6764), .A2(n4358), .ZN(n6741) );
  NOR2_X1 U5917 ( .A1(n6741), .A2(n6740), .ZN(n6739) );
  INV_X1 U5918 ( .A(n4571), .ZN(n6755) );
  AND2_X1 U5919 ( .A1(n6758), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n4678) );
  INV_X1 U5920 ( .A(n4569), .ZN(n9900) );
  INV_X1 U5921 ( .A(n9964), .ZN(n9915) );
  NAND2_X1 U5922 ( .A1(n6558), .A2(n6557), .ZN(n9579) );
  NAND2_X1 U5923 ( .A1(n6438), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n8081) );
  INV_X1 U5924 ( .A(n6440), .ZN(n6438) );
  NAND2_X1 U5925 ( .A1(n6532), .A2(n6531), .ZN(n8085) );
  OAI21_X1 U5926 ( .B1(n9682), .B2(n4846), .A(n4845), .ZN(n9637) );
  INV_X1 U5927 ( .A(n9809), .ZN(n9664) );
  OR2_X1 U5928 ( .A1(n9669), .A2(n4732), .ZN(n9654) );
  INV_X1 U5929 ( .A(n4848), .ZN(n9653) );
  AOI21_X1 U5930 ( .B1(n9682), .B2(n4853), .A(n4851), .ZN(n4848) );
  AND2_X1 U5931 ( .A1(n4720), .A2(n4724), .ZN(n9685) );
  AND2_X1 U5932 ( .A1(n4814), .A2(n4812), .ZN(n9698) );
  INV_X1 U5933 ( .A(n4815), .ZN(n4812) );
  NAND2_X1 U5934 ( .A1(n4816), .A2(n4818), .ZN(n9713) );
  NAND2_X1 U5935 ( .A1(n9743), .A2(n4355), .ZN(n4816) );
  AND2_X1 U5936 ( .A1(n4404), .A2(n7996), .ZN(n9737) );
  NAND2_X1 U5937 ( .A1(n4820), .A2(n4824), .ZN(n9728) );
  OR2_X1 U5938 ( .A1(n9743), .A2(n8060), .ZN(n4820) );
  CLKBUF_X1 U5939 ( .A(n7993), .Z(n7717) );
  NAND2_X1 U5940 ( .A1(n7684), .A2(n4979), .ZN(n4859) );
  OAI21_X1 U5941 ( .B1(n7554), .B2(n7965), .A(n4841), .ZN(n7458) );
  AND2_X1 U5942 ( .A1(n9984), .A2(n10131), .ZN(n7560) );
  NAND2_X1 U5943 ( .A1(n5990), .A2(n5989), .ZN(n10018) );
  AND2_X1 U5944 ( .A1(n10070), .A2(n10041), .ZN(n10017) );
  CLKBUF_X1 U5945 ( .A(n7370), .Z(n4405) );
  NAND2_X1 U5946 ( .A1(n6477), .A2(n7985), .ZN(n10062) );
  AND2_X1 U5947 ( .A1(n6818), .A2(n6602), .ZN(n6482) );
  NOR2_X1 U5948 ( .A1(n9789), .A2(n4978), .ZN(n9792) );
  NOR2_X1 U5949 ( .A1(n9794), .A2(n4297), .ZN(n9797) );
  AND2_X1 U5950 ( .A1(n9796), .A2(n9858), .ZN(n4447) );
  NAND2_X1 U5951 ( .A1(n4506), .A2(n4503), .ZN(n9866) );
  INV_X1 U5952 ( .A(n9799), .ZN(n4506) );
  INV_X1 U5953 ( .A(n4504), .ZN(n4503) );
  OAI21_X1 U5954 ( .B1(n9801), .B2(n9861), .A(n4320), .ZN(n4504) );
  INV_X1 U5955 ( .A(n10076), .ZN(n10074) );
  NAND2_X1 U5956 ( .A1(n5866), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5868) );
  XNOR2_X1 U5957 ( .A(n5700), .B(n5699), .ZN(n7610) );
  INV_X1 U5958 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7289) );
  INV_X1 U5959 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n9104) );
  INV_X1 U5960 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n9072) );
  AND2_X1 U5961 ( .A1(n6166), .A2(n6181), .ZN(n7305) );
  AND2_X1 U5962 ( .A1(n6093), .A2(n6092), .ZN(n6948) );
  INV_X1 U5963 ( .A(n5435), .ZN(n5437) );
  CLKBUF_X1 U5964 ( .A(n5434), .Z(n5435) );
  XNOR2_X1 U5965 ( .A(n6057), .B(P1_IR_REG_7__SCAN_IN), .ZN(n6936) );
  XNOR2_X1 U5966 ( .A(n6034), .B(P1_IR_REG_6__SCAN_IN), .ZN(n6925) );
  CLKBUF_X1 U5967 ( .A(n9522), .Z(n4431) );
  NAND2_X1 U5968 ( .A1(n5909), .A2(n5884), .ZN(n4429) );
  OAI211_X1 U5969 ( .C1(n7077), .C2(n4796), .A(n4795), .B(n4791), .ZN(n7202)
         );
  OAI211_X1 U5970 ( .C1(n5132), .C2(n8645), .A(n4415), .B(n4379), .ZN(P2_U3201) );
  OR2_X1 U5971 ( .A1(n5197), .A2(n8626), .ZN(n4379) );
  AND2_X1 U5972 ( .A1(n5198), .A2(n5196), .ZN(n4415) );
  NAND2_X1 U5973 ( .A1(n4269), .A2(n4513), .ZN(n4512) );
  AOI211_X1 U5974 ( .C1(n8034), .C2(n8033), .A(n8032), .B(n8031), .ZN(n8035)
         );
  AND3_X1 U5975 ( .A1(n9967), .A2(n9966), .A3(n9965), .ZN(n9969) );
  AOI21_X1 U5976 ( .B1(n6609), .B2(n6294), .A(n6608), .ZN(n4378) );
  NAND2_X1 U5977 ( .A1(n10160), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n4725) );
  NAND2_X1 U5978 ( .A1(n9863), .A2(n10162), .ZN(n4726) );
  NAND2_X1 U5979 ( .A1(n6617), .A2(n6616), .ZN(P1_U3520) );
  NAND2_X1 U5980 ( .A1(n4382), .A2(n4381), .ZN(P1_U3519) );
  NAND2_X1 U5981 ( .A1(n10144), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n4381) );
  NAND2_X1 U5982 ( .A1(n9863), .A2(n10145), .ZN(n4382) );
  INV_X1 U5983 ( .A(n8312), .ZN(n4944) );
  AND2_X1 U5984 ( .A1(n4599), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n4275) );
  INV_X1 U5985 ( .A(n8823), .ZN(n4930) );
  OR2_X1 U5986 ( .A1(n5529), .A2(SI_14_), .ZN(n4276) );
  INV_X1 U5987 ( .A(n7834), .ZN(n9747) );
  AND2_X1 U5988 ( .A1(n4897), .A2(n9695), .ZN(n4277) );
  INV_X1 U5989 ( .A(n7759), .ZN(n4698) );
  INV_X1 U5990 ( .A(n8320), .ZN(n4910) );
  INV_X1 U5991 ( .A(n8004), .ZN(n7945) );
  INV_X1 U5992 ( .A(n6455), .ZN(n4394) );
  AND4_X1 U5993 ( .A1(n6189), .A2(n6188), .A3(n6187), .A4(n6186), .ZN(n7700)
         );
  AND2_X1 U5994 ( .A1(n4752), .A2(n7231), .ZN(n4278) );
  AND2_X1 U5995 ( .A1(n5528), .A2(n8847), .ZN(n4279) );
  INV_X1 U5996 ( .A(n4694), .ZN(n4693) );
  NAND2_X1 U5997 ( .A1(n4698), .A2(n4309), .ZN(n4694) );
  NAND2_X1 U5998 ( .A1(n4811), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n4810) );
  NAND2_X1 U5999 ( .A1(n5284), .A2(n5283), .ZN(n5513) );
  AND2_X1 U6000 ( .A1(n4647), .A2(n6778), .ZN(n4280) );
  NAND2_X1 U6001 ( .A1(n4608), .A2(n7529), .ZN(n7475) );
  INV_X1 U6002 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n9105) );
  OR2_X1 U6003 ( .A1(n6294), .A2(n7886), .ZN(n7877) );
  INV_X2 U6004 ( .A(n10188), .ZN(n10185) );
  INV_X1 U6005 ( .A(n8598), .ZN(n4607) );
  INV_X2 U6006 ( .A(n5991), .ZN(n6060) );
  INV_X1 U6007 ( .A(n5457), .ZN(n8132) );
  AND2_X1 U6008 ( .A1(n5534), .A2(n5533), .ZN(n8361) );
  INV_X1 U6009 ( .A(n5460), .ZN(n4796) );
  NAND2_X1 U6010 ( .A1(n4639), .A2(n6670), .ZN(n8741) );
  OR2_X1 U6011 ( .A1(n5590), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n4281) );
  AND2_X1 U6012 ( .A1(n8639), .A2(n5108), .ZN(n4282) );
  XNOR2_X1 U6013 ( .A(n5016), .B(P2_IR_REG_21__SCAN_IN), .ZN(n8295) );
  NAND2_X1 U6014 ( .A1(n5514), .A2(n5513), .ZN(n4283) );
  INV_X1 U6015 ( .A(n8875), .ZN(n9260) );
  INV_X1 U6016 ( .A(n7136), .ZN(n8536) );
  AND4_X1 U6017 ( .A1(n5405), .A2(n5404), .A3(n5403), .A4(n5402), .ZN(n7136)
         );
  OR2_X1 U6018 ( .A1(n9626), .A2(n8074), .ZN(n4284) );
  INV_X1 U6019 ( .A(n5349), .ZN(n5368) );
  NAND2_X1 U6020 ( .A1(n5614), .A2(n5613), .ZN(n4285) );
  AND2_X1 U6021 ( .A1(n4798), .A2(n4796), .ZN(n4286) );
  XNOR2_X1 U6022 ( .A(n5280), .B(SI_11_), .ZN(n5493) );
  OR2_X1 U6023 ( .A1(n5556), .A2(n5287), .ZN(n4287) );
  INV_X1 U6024 ( .A(n8477), .ZN(n4669) );
  AND2_X1 U6025 ( .A1(n7456), .A2(n4896), .ZN(n4288) );
  NAND2_X1 U6026 ( .A1(n9619), .A2(n9631), .ZN(n4289) );
  AND2_X1 U6027 ( .A1(n5200), .A2(n4520), .ZN(n4290) );
  NOR2_X1 U6028 ( .A1(n4385), .A2(P1_IR_REG_14__SCAN_IN), .ZN(n6215) );
  NOR2_X1 U6029 ( .A1(n7946), .A2(n8010), .ZN(n8016) );
  NAND2_X1 U6030 ( .A1(n5391), .A2(n8537), .ZN(n4291) );
  OR2_X1 U6031 ( .A1(n9407), .A2(n9497), .ZN(n4292) );
  AND2_X1 U6032 ( .A1(n6216), .A2(n4705), .ZN(n4293) );
  INV_X1 U6033 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n5035) );
  OAI21_X1 U6034 ( .B1(n9682), .B2(n8066), .A(n8065), .ZN(n9667) );
  NAND2_X1 U6035 ( .A1(n4859), .A2(n7686), .ZN(n7715) );
  AND2_X1 U6036 ( .A1(n4556), .A2(n5513), .ZN(n4294) );
  INV_X1 U6037 ( .A(n7997), .ZN(n4717) );
  AND2_X1 U6038 ( .A1(n8535), .A2(n7257), .ZN(n4295) );
  AND2_X1 U6039 ( .A1(n7888), .A2(n7882), .ZN(n4296) );
  INV_X1 U6040 ( .A(n8476), .ZN(n4929) );
  AND3_X1 U6041 ( .A1(n8112), .A2(n8222), .A3(n8110), .ZN(n4298) );
  AND2_X1 U6042 ( .A1(n9604), .A2(n4733), .ZN(n4299) );
  NAND2_X1 U6043 ( .A1(n6168), .A2(n6167), .ZN(n7705) );
  INV_X1 U6044 ( .A(n7705), .ZN(n7461) );
  INV_X1 U6045 ( .A(n9772), .ZN(n9739) );
  NAND2_X1 U6046 ( .A1(n6233), .A2(n6232), .ZN(n9857) );
  AND2_X1 U6047 ( .A1(n6255), .A2(n6248), .ZN(n4300) );
  AND3_X1 U6048 ( .A1(n8135), .A2(n8140), .A3(n8216), .ZN(n4301) );
  AOI21_X1 U6049 ( .B1(n8055), .B2(n10013), .A(n8054), .ZN(n9787) );
  NOR2_X1 U6050 ( .A1(n8490), .A2(n8336), .ZN(n4302) );
  NOR2_X1 U6051 ( .A1(n8046), .A2(n7869), .ZN(n4303) );
  AND2_X1 U6052 ( .A1(n8390), .A2(n8474), .ZN(n4304) );
  OR2_X1 U6053 ( .A1(n6442), .A2(n10014), .ZN(n4305) );
  INV_X1 U6054 ( .A(n9767), .ZN(n9843) );
  AND2_X1 U6055 ( .A1(n6263), .A2(n6262), .ZN(n9767) );
  NAND2_X1 U6056 ( .A1(n6491), .A2(n6490), .ZN(n9488) );
  AND2_X1 U6057 ( .A1(n4894), .A2(n9767), .ZN(n4306) );
  OR2_X1 U6058 ( .A1(n9213), .A2(n8779), .ZN(n8391) );
  INV_X1 U6059 ( .A(n9695), .ZN(n9819) );
  AND2_X1 U6060 ( .A1(n5843), .A2(n5842), .ZN(n9695) );
  AND2_X1 U6061 ( .A1(n6142), .A2(n6141), .ZN(n10140) );
  NAND2_X1 U6062 ( .A1(n8163), .A2(n8236), .ZN(n4307) );
  OR2_X1 U6063 ( .A1(n5034), .A2(n5134), .ZN(n4308) );
  AND2_X1 U6064 ( .A1(n7757), .A2(n4699), .ZN(n4309) );
  AND2_X1 U6065 ( .A1(n5750), .A2(n5789), .ZN(n4310) );
  NAND2_X1 U6066 ( .A1(n9729), .A2(n4277), .ZN(n4898) );
  INV_X1 U6067 ( .A(n8359), .ZN(n4931) );
  AND2_X1 U6068 ( .A1(n6219), .A2(n6218), .ZN(n9486) );
  INV_X1 U6069 ( .A(n9486), .ZN(n9852) );
  NAND2_X1 U6070 ( .A1(n9814), .A2(n8067), .ZN(n8042) );
  AND2_X1 U6071 ( .A1(n8063), .A2(n8062), .ZN(n4311) );
  AND4_X1 U6072 ( .A1(n8383), .A2(n8382), .A3(n8390), .A4(n8474), .ZN(n4312)
         );
  NAND2_X1 U6073 ( .A1(n8048), .A2(n7978), .ZN(n9586) );
  INV_X1 U6074 ( .A(n9586), .ZN(n4827) );
  AND2_X1 U6075 ( .A1(n7969), .A2(n7827), .ZN(n4313) );
  AND2_X1 U6076 ( .A1(P1_REG3_REG_10__SCAN_IN), .A2(P1_REG3_REG_11__SCAN_IN), 
        .ZN(n4314) );
  AND2_X1 U6077 ( .A1(n4692), .A2(n4691), .ZN(n4315) );
  AND2_X1 U6078 ( .A1(n7037), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n4316) );
  AND2_X1 U6079 ( .A1(n6522), .A2(n6521), .ZN(n9599) );
  INV_X1 U6080 ( .A(n9599), .ZN(n9788) );
  AND2_X1 U6081 ( .A1(n4288), .A2(n7461), .ZN(n4317) );
  OR2_X1 U6082 ( .A1(n4930), .A2(n4669), .ZN(n4318) );
  OR2_X1 U6083 ( .A1(n4554), .A2(n4558), .ZN(n4319) );
  NOR2_X1 U6084 ( .A1(n4973), .A2(n4505), .ZN(n4320) );
  NOR2_X1 U6085 ( .A1(n5731), .A2(n8687), .ZN(n4321) );
  INV_X1 U6086 ( .A(n4655), .ZN(n4654) );
  OR2_X1 U6087 ( .A1(n6685), .A2(n4656), .ZN(n4655) );
  OR2_X1 U6088 ( .A1(n8361), .A2(n6667), .ZN(n4322) );
  NAND2_X1 U6089 ( .A1(n5019), .A2(n5018), .ZN(n4323) );
  INV_X1 U6090 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n4995) );
  OR2_X1 U6091 ( .A1(n5605), .A2(n8779), .ZN(n4324) );
  AND2_X1 U6092 ( .A1(n6697), .A2(n8673), .ZN(n4325) );
  NOR2_X1 U6093 ( .A1(n7418), .A2(n9976), .ZN(n4326) );
  AND2_X1 U6094 ( .A1(n9731), .A2(n9717), .ZN(n4327) );
  AND2_X1 U6095 ( .A1(n9220), .A2(n8793), .ZN(n8475) );
  OR2_X1 U6096 ( .A1(n8314), .A2(n4912), .ZN(n4328) );
  INV_X1 U6097 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n5037) );
  NOR2_X1 U6098 ( .A1(n9241), .A2(n8830), .ZN(n4329) );
  INV_X1 U6099 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n5000) );
  AND2_X1 U6100 ( .A1(n4932), .A2(n4927), .ZN(n4330) );
  AND2_X1 U6101 ( .A1(n4552), .A2(n4319), .ZN(n4331) );
  AND2_X1 U6102 ( .A1(n8407), .A2(n8440), .ZN(n4332) );
  AND2_X1 U6103 ( .A1(n6435), .A2(n6434), .ZN(n6456) );
  INV_X1 U6104 ( .A(n6456), .ZN(n4393) );
  AND2_X1 U6105 ( .A1(n4823), .A2(n8061), .ZN(n4333) );
  NAND2_X1 U6106 ( .A1(n9786), .A2(n9785), .ZN(n4334) );
  INV_X1 U6107 ( .A(n4559), .ZN(n4558) );
  NOR2_X1 U6108 ( .A1(n5280), .A2(SI_11_), .ZN(n4559) );
  INV_X1 U6109 ( .A(n5871), .ZN(n6150) );
  NAND2_X1 U6110 ( .A1(n6357), .A2(n6356), .ZN(n9814) );
  INV_X1 U6111 ( .A(n4555), .ZN(n4554) );
  NAND2_X1 U6112 ( .A1(n4336), .A2(n5513), .ZN(n4555) );
  OR2_X1 U6113 ( .A1(n7714), .A2(n4858), .ZN(n4335) );
  NAND2_X1 U6114 ( .A1(n5511), .A2(n5514), .ZN(n4336) );
  INV_X1 U6115 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n4938) );
  OR2_X1 U6116 ( .A1(n4818), .A2(n4817), .ZN(n4337) );
  OR2_X1 U6117 ( .A1(n9445), .A2(n9495), .ZN(n4338) );
  AND2_X1 U6118 ( .A1(n5392), .A2(n5384), .ZN(n4339) );
  AND2_X1 U6119 ( .A1(n5034), .A2(n4618), .ZN(n4340) );
  AND2_X1 U6120 ( .A1(n7923), .A2(n7825), .ZN(n4341) );
  NOR2_X1 U6121 ( .A1(n8122), .A2(n4762), .ZN(n4761) );
  AND2_X1 U6122 ( .A1(n8565), .A2(n5096), .ZN(n4342) );
  AND2_X1 U6123 ( .A1(n7822), .A2(n7823), .ZN(n4343) );
  NOR2_X1 U6124 ( .A1(n8046), .A2(n7866), .ZN(n4344) );
  AND2_X1 U6125 ( .A1(n7837), .A2(n7924), .ZN(n4345) );
  INV_X1 U6126 ( .A(n8069), .ZN(n4855) );
  INV_X1 U6127 ( .A(n8364), .ZN(n4664) );
  AND2_X1 U6128 ( .A1(n7955), .A2(n7994), .ZN(n4346) );
  AND2_X1 U6129 ( .A1(n4333), .A2(n4824), .ZN(n4347) );
  OR2_X1 U6130 ( .A1(n9857), .A2(n9425), .ZN(n7929) );
  AND2_X1 U6131 ( .A1(n4860), .A2(n4979), .ZN(n4348) );
  AND2_X1 U6132 ( .A1(n5976), .A2(n5974), .ZN(n4349) );
  AND2_X1 U6133 ( .A1(n4839), .A2(n4292), .ZN(n4350) );
  AND2_X1 U6134 ( .A1(n4290), .A2(n5202), .ZN(n4351) );
  AND2_X1 U6135 ( .A1(n4602), .A2(n4607), .ZN(n4352) );
  AND2_X1 U6136 ( .A1(n7840), .A2(n7929), .ZN(n4353) );
  OR2_X1 U6137 ( .A1(n9430), .A2(n7700), .ZN(n7928) );
  NAND2_X1 U6138 ( .A1(n7908), .A2(n7905), .ZN(n7487) );
  NAND2_X1 U6139 ( .A1(n9984), .A2(n4288), .ZN(n7412) );
  INV_X1 U6140 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n4463) );
  INV_X1 U6141 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n4496) );
  INV_X1 U6142 ( .A(n10068), .ZN(n10015) );
  NAND2_X1 U6143 ( .A1(n10027), .A2(n6482), .ZN(n10068) );
  AOI21_X1 U6144 ( .B1(n9972), .B2(n7419), .A(n4326), .ZN(n7509) );
  AOI21_X1 U6145 ( .B1(n7598), .B2(n8493), .A(n6662), .ZN(n8844) );
  INV_X1 U6146 ( .A(n4743), .ZN(n5772) );
  NAND2_X1 U6147 ( .A1(n4685), .A2(n6160), .ZN(n7697) );
  NAND2_X1 U6148 ( .A1(n4969), .A2(n6629), .ZN(n8840) );
  NAND2_X1 U6149 ( .A1(n7691), .A2(n4306), .ZN(n4895) );
  AND2_X1 U6150 ( .A1(n4824), .A2(n4823), .ZN(n4355) );
  AND2_X1 U6151 ( .A1(n4600), .A2(n4596), .ZN(n4356) );
  AND2_X1 U6152 ( .A1(n4611), .A2(n7281), .ZN(n4357) );
  AND2_X1 U6153 ( .A1(n6770), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n4358) );
  INV_X1 U6154 ( .A(n4772), .ZN(n8109) );
  NAND2_X1 U6155 ( .A1(n7449), .A2(n5445), .ZN(n4772) );
  INV_X1 U6156 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n9113) );
  NOR2_X1 U6157 ( .A1(n5474), .A2(n9024), .ZN(n4359) );
  OAI21_X1 U6158 ( .B1(n4744), .B2(P2_D_REG_0__SCAN_IN), .A(n6800), .ZN(n4743)
         );
  OR2_X1 U6159 ( .A1(n9664), .A2(n9485), .ZN(n4360) );
  AND2_X1 U6160 ( .A1(n6770), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n4361) );
  AND2_X1 U6161 ( .A1(n5083), .A2(n7529), .ZN(n4362) );
  AND2_X1 U6162 ( .A1(n6517), .A2(n6519), .ZN(n4363) );
  NOR2_X1 U6163 ( .A1(n5190), .A2(P2_U3151), .ZN(n4364) );
  INV_X1 U6164 ( .A(n10162), .ZN(n10160) );
  INV_X1 U6165 ( .A(n5186), .ZN(n4590) );
  NAND2_X1 U6166 ( .A1(n6036), .A2(n6035), .ZN(n10001) );
  INV_X1 U6167 ( .A(n10001), .ZN(n7360) );
  AND2_X1 U6168 ( .A1(n9908), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n4365) );
  INV_X1 U6169 ( .A(n6914), .ZN(n4937) );
  INV_X1 U6170 ( .A(n10013), .ZN(n10047) );
  NAND2_X1 U6171 ( .A1(n7986), .A2(n7001), .ZN(n10013) );
  XOR2_X1 U6172 ( .A(n4274), .B(n8960), .Z(n4366) );
  NAND2_X2 U6173 ( .A1(n6184), .A2(n6183), .ZN(n9430) );
  NAND2_X1 U6174 ( .A1(n4688), .A2(n5985), .ZN(n9392) );
  AND2_X1 U6175 ( .A1(n8589), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n4367) );
  OR2_X1 U6176 ( .A1(n4589), .A2(n4586), .ZN(n4368) );
  AND2_X1 U6177 ( .A1(n8629), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n4369) );
  OR2_X1 U6178 ( .A1(n10185), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n4370) );
  AND2_X1 U6179 ( .A1(n8589), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n4371) );
  AND2_X1 U6180 ( .A1(n5055), .A2(n6891), .ZN(n4372) );
  AND2_X1 U6181 ( .A1(n4756), .A2(n4291), .ZN(n4373) );
  OR2_X1 U6182 ( .A1(n8614), .A2(n5180), .ZN(n4374) );
  INV_X1 U6183 ( .A(n6777), .ZN(n4647) );
  INV_X1 U6184 ( .A(n4744), .ZN(n6795) );
  NAND2_X1 U6185 ( .A1(n5315), .A2(n5316), .ZN(n4744) );
  INV_X1 U6186 ( .A(n7159), .ZN(n4418) );
  INV_X1 U6187 ( .A(n7985), .ZN(n7886) );
  XNOR2_X1 U6188 ( .A(n5901), .B(n5900), .ZN(n7985) );
  INV_X1 U6189 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n7142) );
  INV_X1 U6190 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n4495) );
  INV_X1 U6191 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n4594) );
  INV_X1 U6192 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n4468) );
  INV_X1 U6193 ( .A(n8641), .ZN(n4586) );
  NAND2_X1 U6194 ( .A1(n8641), .A2(n4582), .ZN(n4581) );
  NOR2_X2 U6195 ( .A1(n5131), .A2(n4270), .ZN(n8641) );
  NAND2_X1 U6196 ( .A1(n4551), .A2(n4555), .ZN(n5531) );
  INV_X1 U6197 ( .A(n5499), .ZN(n4557) );
  AOI21_X1 U6198 ( .B1(n4902), .B2(n8449), .A(n8448), .ZN(n8520) );
  AND2_X1 U6199 ( .A1(n8422), .A2(n8421), .ZN(n4908) );
  OAI211_X2 U6200 ( .C1(n5908), .C2(n5909), .A(n5969), .B(n4429), .ZN(n6780)
         );
  NAND3_X1 U6201 ( .A1(n4375), .A2(n6601), .A3(n9948), .ZN(n4430) );
  NAND2_X1 U6202 ( .A1(n6603), .A2(n9957), .ZN(n4375) );
  NOR2_X2 U6203 ( .A1(n9931), .A2(n9930), .ZN(n9929) );
  NOR2_X1 U6204 ( .A1(n9550), .A2(n4560), .ZN(n6907) );
  OAI21_X1 U6205 ( .B1(n7305), .B2(P1_REG2_REG_12__SCAN_IN), .A(n7298), .ZN(
        n6756) );
  NOR2_X1 U6206 ( .A1(n6742), .A2(n4572), .ZN(n7299) );
  NOR2_X1 U6207 ( .A1(n6905), .A2(n4575), .ZN(n6924) );
  NAND2_X1 U6208 ( .A1(n4378), .A2(n6610), .ZN(P1_U3262) );
  INV_X1 U6209 ( .A(n8388), .ZN(n4426) );
  OAI21_X1 U6210 ( .B1(n8423), .B2(n8412), .A(n4904), .ZN(n4903) );
  NAND2_X1 U6211 ( .A1(n4810), .A2(n4340), .ZN(n6866) );
  AOI21_X1 U6212 ( .B1(n8586), .B2(n8587), .A(n4371), .ZN(n5130) );
  NAND2_X1 U6213 ( .A1(n4384), .A2(n4383), .ZN(n7363) );
  NAND2_X1 U6214 ( .A1(n7581), .A2(n7357), .ZN(n4383) );
  AND2_X1 U6215 ( .A1(n7361), .A2(n9999), .ZN(n4384) );
  INV_X2 U6216 ( .A(n7344), .ZN(n10011) );
  NAND2_X2 U6217 ( .A1(n8073), .A2(n8072), .ZN(n9622) );
  NAND2_X1 U6218 ( .A1(n4838), .A2(n4836), .ZN(n7614) );
  NAND2_X1 U6219 ( .A1(n4835), .A2(n4350), .ZN(n4838) );
  OAI21_X1 U6220 ( .B1(n7614), .B2(n4983), .A(n4840), .ZN(n7616) );
  AOI21_X1 U6221 ( .B1(n9682), .B2(n4845), .A(n4843), .ZN(n4842) );
  NAND3_X1 U6222 ( .A1(n7490), .A2(n10019), .A3(n7491), .ZN(n7354) );
  NAND2_X1 U6223 ( .A1(n7146), .A2(n7147), .ZN(n4688) );
  AOI21_X1 U6224 ( .B1(n6317), .B2(n6316), .A(n9324), .ZN(n9416) );
  OAI21_X2 U6225 ( .B1(n7407), .B2(n7919), .A(n7918), .ZN(n7462) );
  OAI21_X1 U6226 ( .B1(n7753), .B2(n4690), .A(n4689), .ZN(n4697) );
  NOR2_X2 U6227 ( .A1(n9460), .A2(n4392), .ZN(n9352) );
  NAND2_X2 U6228 ( .A1(n5896), .A2(n7949), .ZN(n7420) );
  NAND2_X1 U6229 ( .A1(n9748), .A2(n7995), .ZN(n9751) );
  NAND2_X1 U6230 ( .A1(n4679), .A2(n4682), .ZN(n9422) );
  NOR2_X2 U6231 ( .A1(n9463), .A2(n6432), .ZN(n9460) );
  AND4_X2 U6232 ( .A1(n5915), .A2(n5917), .A3(n5916), .A4(n5918), .ZN(n10049)
         );
  NAND2_X1 U6233 ( .A1(n6337), .A2(n6336), .ZN(n9353) );
  OAI21_X2 U6234 ( .B1(n9353), .B2(n9354), .A(n6355), .ZN(n7753) );
  NOR2_X1 U6235 ( .A1(n5844), .A2(n4893), .ZN(n5898) );
  NAND2_X1 U6236 ( .A1(n4427), .A2(n5871), .ZN(n4981) );
  NAND2_X1 U6237 ( .A1(n4688), .A2(n4686), .ZN(n9394) );
  BUF_X2 U6238 ( .A(n5844), .Z(n4385) );
  NAND2_X1 U6239 ( .A1(n6025), .A2(n6026), .ZN(n7312) );
  NAND2_X1 U6240 ( .A1(n9394), .A2(n6005), .ZN(n6025) );
  NOR2_X1 U6241 ( .A1(n6273), .A2(n4701), .ZN(n4700) );
  XNOR2_X1 U6242 ( .A(n5944), .B(n5945), .ZN(n7112) );
  AOI21_X2 U6243 ( .B1(n9300), .B2(n9299), .A(n9298), .ZN(n9302) );
  NAND2_X1 U6244 ( .A1(n5942), .A2(n5935), .ZN(n6976) );
  NAND3_X1 U6245 ( .A1(n7767), .A2(n7766), .A3(n4360), .ZN(P1_U3229) );
  NAND2_X1 U6246 ( .A1(n7755), .A2(n7754), .ZN(n7770) );
  NAND2_X1 U6247 ( .A1(n6975), .A2(n6976), .ZN(n6978) );
  NAND2_X1 U6248 ( .A1(n4657), .A2(n6682), .ZN(n8709) );
  OAI21_X1 U6249 ( .B1(n4626), .B2(n4354), .A(n4628), .ZN(n6653) );
  OAI21_X1 U6250 ( .B1(n7290), .B2(n7390), .A(n6654), .ZN(n7384) );
  NAND2_X1 U6251 ( .A1(n5116), .A2(n6866), .ZN(n5115) );
  NOR2_X1 U6252 ( .A1(n6886), .A2(n6885), .ZN(n7050) );
  OAI21_X1 U6253 ( .B1(n8604), .B2(n8967), .A(n4782), .ZN(n8621) );
  OAI21_X1 U6254 ( .B1(n4600), .B2(n4598), .A(n4597), .ZN(n5099) );
  NAND2_X1 U6255 ( .A1(n7036), .A2(n5047), .ZN(n5054) );
  NAND2_X1 U6256 ( .A1(n4622), .A2(n5065), .ZN(n4621) );
  NAND2_X1 U6257 ( .A1(n4396), .A2(n8431), .ZN(n4902) );
  NAND3_X1 U6258 ( .A1(n4905), .A2(n4903), .A3(n4908), .ZN(n4396) );
  OAI211_X1 U6259 ( .C1(n8520), .C2(n8519), .A(n4397), .B(n8518), .ZN(n8521)
         );
  NAND3_X1 U6260 ( .A1(n8520), .A2(n8517), .A3(n8516), .ZN(n4397) );
  INV_X1 U6261 ( .A(n8337), .ZN(n4398) );
  NAND2_X1 U6262 ( .A1(n4399), .A2(n8358), .ZN(n8360) );
  NAND2_X1 U6263 ( .A1(n4400), .A2(n6630), .ZN(n4399) );
  NAND2_X1 U6264 ( .A1(n4402), .A2(n4401), .ZN(n4400) );
  NAND2_X1 U6265 ( .A1(n8353), .A2(n8354), .ZN(n4402) );
  NAND2_X1 U6266 ( .A1(n8397), .A2(n4403), .ZN(n8401) );
  NAND2_X1 U6267 ( .A1(n8396), .A2(n4312), .ZN(n4403) );
  NAND2_X1 U6268 ( .A1(n8380), .A2(n8379), .ZN(n8396) );
  NAND2_X2 U6269 ( .A1(n7688), .A2(n7972), .ZN(n7716) );
  NAND2_X1 U6270 ( .A1(n9585), .A2(n4827), .ZN(n9589) );
  NAND2_X2 U6271 ( .A1(n7624), .A2(n4313), .ZN(n7655) );
  NAND2_X1 U6272 ( .A1(n5907), .A2(n6777), .ZN(n5912) );
  NAND2_X2 U6273 ( .A1(n7793), .A2(n7913), .ZN(n7583) );
  NAND2_X1 U6274 ( .A1(n4728), .A2(n4729), .ZN(n9640) );
  NAND2_X1 U6275 ( .A1(n4722), .A2(n4721), .ZN(n4720) );
  NAND2_X1 U6276 ( .A1(n5878), .A2(n5877), .ZN(n6321) );
  NAND2_X1 U6277 ( .A1(n5876), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n6265) );
  NAND2_X1 U6278 ( .A1(n5874), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n6097) );
  OR2_X1 U6279 ( .A1(n7808), .A2(n7803), .ZN(n7402) );
  NAND2_X1 U6280 ( .A1(n4720), .A2(n4718), .ZN(n9683) );
  INV_X1 U6281 ( .A(n6341), .ZN(n5879) );
  NAND2_X1 U6282 ( .A1(n5235), .A2(SI_1_), .ZN(n5335) );
  NAND3_X1 U6283 ( .A1(n9579), .A2(n4409), .A3(n9487), .ZN(n4408) );
  NAND2_X1 U6284 ( .A1(n7655), .A2(n4713), .ZN(n4714) );
  NAND2_X1 U6285 ( .A1(n9751), .A2(n4723), .ZN(n4722) );
  NAND2_X1 U6286 ( .A1(n9671), .A2(n4731), .ZN(n4728) );
  NAND2_X1 U6287 ( .A1(n4734), .A2(n4511), .ZN(n4510) );
  NAND2_X1 U6288 ( .A1(n5434), .A2(n5270), .ZN(n5438) );
  NAND2_X1 U6289 ( .A1(n6399), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n6414) );
  NOR2_X1 U6290 ( .A1(n9913), .A2(n9914), .ZN(n9912) );
  NOR2_X2 U6291 ( .A1(n9929), .A2(n4448), .ZN(n9939) );
  NAND4_X1 U6292 ( .A1(n4446), .A2(n4933), .A3(n4994), .A4(n5074), .ZN(n5026)
         );
  OAI21_X1 U6293 ( .B1(n7050), .B2(n7049), .A(n7048), .ZN(n7083) );
  INV_X2 U6294 ( .A(n6477), .ZN(n5896) );
  NAND2_X1 U6295 ( .A1(n4484), .A2(n4483), .ZN(n5298) );
  NAND2_X1 U6296 ( .A1(n4651), .A2(n4658), .ZN(n4650) );
  OAI21_X1 U6297 ( .B1(n5609), .B2(n5245), .A(n5244), .ZN(n5257) );
  INV_X1 U6298 ( .A(n5182), .ZN(n5185) );
  NAND2_X1 U6299 ( .A1(n8610), .A2(n4374), .ZN(n5182) );
  NOR2_X1 U6300 ( .A1(n6696), .A2(n6695), .ZN(n8654) );
  NAND2_X1 U6301 ( .A1(n9537), .A2(n9538), .ZN(n9536) );
  NAND2_X1 U6302 ( .A1(n9925), .A2(n4416), .ZN(n9942) );
  NAND2_X1 U6303 ( .A1(n9942), .A2(n9943), .ZN(n6598) );
  NOR2_X1 U6304 ( .A1(n6739), .A2(n4675), .ZN(n7303) );
  NOR2_X1 U6305 ( .A1(n6933), .A2(n4677), .ZN(n6947) );
  AOI21_X1 U6306 ( .B1(n6908), .B2(P1_REG1_REG_5__SCAN_IN), .A(n6902), .ZN(
        n6921) );
  NAND2_X1 U6307 ( .A1(n5987), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4576) );
  OAI22_X1 U6308 ( .A1(n6604), .A2(n9915), .B1(n6603), .B2(n9928), .ZN(n6609)
         );
  XNOR2_X1 U6309 ( .A(n6600), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n6604) );
  NAND2_X1 U6310 ( .A1(n9927), .A2(n9926), .ZN(n9925) );
  NOR2_X1 U6311 ( .A1(n9916), .A2(n6596), .ZN(n9927) );
  XNOR2_X1 U6312 ( .A(n6595), .B(n7107), .ZN(n9918) );
  NAND2_X1 U6313 ( .A1(n7303), .A2(n7304), .ZN(n7302) );
  NAND2_X1 U6314 ( .A1(n9567), .A2(n9566), .ZN(n9565) );
  NAND2_X1 U6315 ( .A1(n4528), .A2(n5788), .ZN(n4527) );
  NAND2_X1 U6316 ( .A1(n4759), .A2(n4757), .ZN(n8226) );
  OAI21_X1 U6317 ( .B1(n5927), .B2(n6150), .A(n5932), .ZN(n5933) );
  NAND2_X1 U6318 ( .A1(n5919), .A2(n4981), .ZN(n4459) );
  NAND2_X1 U6319 ( .A1(n5857), .A2(n5856), .ZN(n5861) );
  NAND2_X1 U6320 ( .A1(n5898), .A2(n5900), .ZN(n6475) );
  INV_X1 U6321 ( .A(n6475), .ZN(n5857) );
  NAND2_X1 U6322 ( .A1(n6540), .A2(n6539), .ZN(n6550) );
  XNOR2_X1 U6323 ( .A(n6585), .B(P1_REG2_REG_19__SCAN_IN), .ZN(n6603) );
  NAND2_X1 U6324 ( .A1(n4577), .A2(n5970), .ZN(n5987) );
  NAND2_X1 U6325 ( .A1(n9528), .A2(n9527), .ZN(n9526) );
  NAND2_X1 U6326 ( .A1(n4430), .A2(n6602), .ZN(n6610) );
  NAND2_X1 U6327 ( .A1(n7299), .A2(n7300), .ZN(n7298) );
  NAND2_X1 U6328 ( .A1(n9539), .A2(n6578), .ZN(n9548) );
  NOR2_X1 U6329 ( .A1(n6744), .A2(n6743), .ZN(n6742) );
  NAND2_X1 U6330 ( .A1(n7852), .A2(n4432), .ZN(n4479) );
  NAND3_X1 U6331 ( .A1(n4476), .A2(n4442), .A3(n7851), .ZN(n4432) );
  NAND2_X1 U6332 ( .A1(n4433), .A2(n4346), .ZN(n7835) );
  NAND2_X1 U6333 ( .A1(n7833), .A2(n7957), .ZN(n4433) );
  XNOR2_X2 U6334 ( .A(n5852), .B(n5851), .ZN(n6477) );
  INV_X2 U6335 ( .A(n7356), .ZN(n9500) );
  INV_X1 U6336 ( .A(n4928), .ZN(n4927) );
  NAND2_X1 U6337 ( .A1(n4610), .A2(n7530), .ZN(n7533) );
  INV_X1 U6338 ( .A(n5082), .ZN(n5081) );
  OAI211_X1 U6339 ( .C1(n8646), .C2(n8645), .A(n8644), .B(n4444), .ZN(P2_U3200) );
  NAND2_X1 U6340 ( .A1(n5240), .A2(n4469), .ZN(n5385) );
  NAND3_X1 U6341 ( .A1(n4475), .A2(n5268), .A3(n4438), .ZN(n5434) );
  NAND2_X1 U6342 ( .A1(n5325), .A2(n5262), .ZN(n4438) );
  NAND2_X1 U6343 ( .A1(n5625), .A2(n5624), .ZN(n5627) );
  INV_X1 U6344 ( .A(n4632), .ZN(n4630) );
  NAND2_X1 U6345 ( .A1(n4660), .A2(n4662), .ZN(n8801) );
  NAND2_X1 U6346 ( .A1(n5258), .A2(n5395), .ZN(n5261) );
  NOR2_X1 U6347 ( .A1(n7885), .A2(n4861), .ZN(n7989) );
  NAND2_X1 U6348 ( .A1(n4439), .A2(n4353), .ZN(n7845) );
  NAND2_X1 U6349 ( .A1(n4480), .A2(n4345), .ZN(n4439) );
  NAND2_X1 U6350 ( .A1(n4440), .A2(n7827), .ZN(n7828) );
  NAND2_X1 U6351 ( .A1(n7826), .A2(n4341), .ZN(n4440) );
  CLKBUF_X2 U6352 ( .A(n10049), .Z(n4441) );
  OAI21_X1 U6353 ( .B1(n7850), .B2(n7934), .A(n4443), .ZN(n4442) );
  NAND4_X2 U6354 ( .A1(n5926), .A2(n5925), .A3(n5924), .A4(n5923), .ZN(n7346)
         );
  AOI21_X2 U6355 ( .B1(n5026), .B2(n5025), .A(n5024), .ZN(n5027) );
  AOI21_X2 U6356 ( .B1(n7993), .B2(n8057), .A(n7992), .ZN(n9770) );
  NAND2_X1 U6357 ( .A1(n9541), .A2(n9540), .ZN(n9539) );
  NAND4_X1 U6358 ( .A1(n8767), .A2(n4453), .A3(n8781), .A4(n4451), .ZN(n4450)
         );
  NOR2_X1 U6359 ( .A1(n6767), .A2(n4361), .ZN(n6744) );
  AOI21_X1 U6360 ( .B1(n6948), .B2(P1_REG2_REG_8__SCAN_IN), .A(n6942), .ZN(
        n9562) );
  OAI21_X1 U6361 ( .B1(n8572), .B2(n8973), .A(n4803), .ZN(n8586) );
  NAND2_X1 U6362 ( .A1(n6888), .A2(n6889), .ZN(n6887) );
  NAND2_X1 U6363 ( .A1(n7824), .A2(n4343), .ZN(n7826) );
  OAI21_X1 U6364 ( .B1(n7832), .B2(n7900), .A(n7930), .ZN(n7833) );
  NAND2_X1 U6365 ( .A1(n7836), .A2(n7928), .ZN(n4480) );
  INV_X1 U6366 ( .A(n10044), .ZN(n7372) );
  NAND2_X1 U6367 ( .A1(n4485), .A2(n4873), .ZN(n5571) );
  NOR3_X1 U6368 ( .A1(n8386), .A2(n8440), .A3(n8389), .ZN(n8387) );
  AND2_X1 U6369 ( .A1(n4461), .A2(n4460), .ZN(n8423) );
  NAND2_X1 U6370 ( .A1(n8406), .A2(n8504), .ZN(n4461) );
  NAND2_X1 U6371 ( .A1(n7467), .A2(n4983), .ZN(n7624) );
  NAND2_X1 U6372 ( .A1(n9770), .A2(n9769), .ZN(n9748) );
  NAND2_X1 U6373 ( .A1(n5879), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n6343) );
  INV_X1 U6374 ( .A(n6401), .ZN(n6399) );
  NAND2_X1 U6375 ( .A1(n4828), .A2(n4826), .ZN(n9583) );
  NAND2_X1 U6376 ( .A1(n4726), .A2(n4725), .ZN(P1_U3551) );
  NOR2_X2 U6377 ( .A1(n5079), .A2(n4624), .ZN(n4623) );
  NAND2_X2 U6378 ( .A1(n4939), .A2(n5073), .ZN(n5079) );
  NAND2_X1 U6379 ( .A1(n5531), .A2(n4876), .ZN(n4485) );
  INV_X1 U6380 ( .A(n5571), .ZN(n4484) );
  NAND2_X1 U6381 ( .A1(n4557), .A2(n4294), .ZN(n4551) );
  NOR2_X1 U6382 ( .A1(n5234), .A2(n5233), .ZN(n5240) );
  NAND3_X1 U6383 ( .A1(n5354), .A2(n5336), .A3(n5339), .ZN(n4469) );
  NAND2_X1 U6384 ( .A1(n4950), .A2(n4946), .ZN(n8753) );
  INV_X1 U6385 ( .A(n8091), .ZN(n4672) );
  NAND2_X1 U6386 ( .A1(n7835), .A2(n4477), .ZN(n4476) );
  OAI21_X2 U6387 ( .B1(n4710), .B2(n4711), .A(n4975), .ZN(n7793) );
  NAND2_X1 U6388 ( .A1(n4868), .A2(n4867), .ZN(n4866) );
  NAND2_X1 U6389 ( .A1(n7868), .A2(n8045), .ZN(n4869) );
  AOI21_X1 U6390 ( .B1(n4474), .B2(n4303), .A(n4472), .ZN(n7872) );
  NAND2_X1 U6391 ( .A1(n4473), .A2(n7877), .ZN(n4472) );
  NAND2_X1 U6392 ( .A1(n7870), .A2(n8045), .ZN(n4474) );
  NAND2_X1 U6393 ( .A1(n7910), .A2(n7913), .ZN(n10024) );
  NAND2_X1 U6394 ( .A1(n7509), .A2(n7510), .ZN(n4835) );
  NAND2_X1 U6395 ( .A1(n5255), .A2(n5385), .ZN(n4475) );
  INV_X2 U6396 ( .A(n5307), .ZN(n5252) );
  NAND2_X1 U6397 ( .A1(n4489), .A2(n4488), .ZN(n4487) );
  NAND2_X1 U6398 ( .A1(n4869), .A2(n4344), .ZN(n4868) );
  INV_X1 U6399 ( .A(n7870), .ZN(n7868) );
  NAND2_X1 U6400 ( .A1(n7828), .A2(n7882), .ZN(n4482) );
  AND4_X2 U6401 ( .A1(n4709), .A2(n4708), .A3(n4707), .A4(n4706), .ZN(n5826)
         );
  NAND2_X1 U6402 ( .A1(n4479), .A2(n7855), .ZN(n7856) );
  NAND2_X4 U6403 ( .A1(n4493), .A2(n4494), .ZN(n5307) );
  NAND2_X2 U6404 ( .A1(n5225), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n4494) );
  NAND2_X2 U6405 ( .A1(n4487), .A2(n5226), .ZN(n4493) );
  INV_X2 U6406 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n4489) );
  NAND3_X1 U6407 ( .A1(n4493), .A2(n4494), .A3(n4495), .ZN(n4490) );
  INV_X1 U6408 ( .A(n4493), .ZN(n4492) );
  OAI21_X2 U6409 ( .B1(n4871), .B2(n4500), .A(n4498), .ZN(n5499) );
  NAND2_X1 U6410 ( .A1(n5201), .A2(n4351), .ZN(n5477) );
  NAND3_X1 U6411 ( .A1(n7142), .A2(n4521), .A3(n5199), .ZN(n5419) );
  NAND2_X1 U6412 ( .A1(n5614), .A2(n4526), .ZN(n5654) );
  NAND3_X1 U6413 ( .A1(n8145), .A2(n4527), .A3(n8216), .ZN(n5822) );
  NAND2_X1 U6414 ( .A1(n5557), .A2(n4542), .ZN(n4536) );
  INV_X1 U6415 ( .A(n5498), .ZN(n4556) );
  OAI21_X1 U6416 ( .B1(n9939), .B2(n4564), .A(n4561), .ZN(n6585) );
  XNOR2_X2 U6417 ( .A(n4576), .B(P1_IR_REG_3__SCAN_IN), .ZN(n9535) );
  INV_X1 U6418 ( .A(n5969), .ZN(n4577) );
  OAI22_X1 U6419 ( .A1(n8640), .A2(n4581), .B1(n4587), .B2(n4586), .ZN(n4578)
         );
  NAND2_X1 U6420 ( .A1(n4282), .A2(n4580), .ZN(n4579) );
  NAND2_X1 U6421 ( .A1(n8640), .A2(n4585), .ZN(n4580) );
  NOR2_X1 U6422 ( .A1(n4586), .A2(n4590), .ZN(n4585) );
  NAND2_X1 U6423 ( .A1(n7033), .A2(n4594), .ZN(n4593) );
  NAND2_X1 U6424 ( .A1(n8539), .A2(n8565), .ZN(n4596) );
  NAND2_X1 U6425 ( .A1(n8539), .A2(n4342), .ZN(n4597) );
  INV_X1 U6426 ( .A(n8539), .ZN(n4599) );
  AOI21_X1 U6427 ( .B1(n8565), .B2(n8837), .A(n4601), .ZN(n4600) );
  OAI21_X2 U6428 ( .B1(n8599), .B2(n8598), .A(n4603), .ZN(n4606) );
  NOR2_X2 U6429 ( .A1(n5102), .A2(n4605), .ZN(n8605) );
  NOR2_X1 U6430 ( .A1(n4606), .A2(n8614), .ZN(n4605) );
  NAND2_X1 U6431 ( .A1(n4609), .A2(n7529), .ZN(n4610) );
  NAND2_X1 U6432 ( .A1(n4617), .A2(n6891), .ZN(n4615) );
  AND2_X1 U6433 ( .A1(n4308), .A2(n4619), .ZN(n6870) );
  NAND3_X1 U6434 ( .A1(n4308), .A2(P2_REG2_REG_1__SCAN_IN), .A3(n4619), .ZN(
        n6869) );
  NAND2_X1 U6435 ( .A1(n4620), .A2(n4340), .ZN(n4619) );
  NAND2_X1 U6436 ( .A1(n5066), .A2(n6791), .ZN(n7088) );
  NAND3_X1 U6437 ( .A1(n4621), .A2(P2_REG2_REG_7__SCAN_IN), .A3(n7088), .ZN(
        n7053) );
  INV_X1 U6438 ( .A(n5066), .ZN(n4622) );
  AND2_X2 U6439 ( .A1(n4623), .A2(n4994), .ZN(n4999) );
  AND4_X2 U6440 ( .A1(n5310), .A2(n4993), .A3(n5008), .A4(n5009), .ZN(n4980)
         );
  AND3_X2 U6441 ( .A1(n4742), .A2(n4740), .A3(n4741), .ZN(n5073) );
  NAND2_X1 U6442 ( .A1(n6669), .A2(n4640), .ZN(n4636) );
  NAND2_X1 U6443 ( .A1(n4636), .A2(n4637), .ZN(n8732) );
  NAND3_X2 U6444 ( .A1(n5362), .A2(n5361), .A3(n4646), .ZN(n7103) );
  NAND2_X1 U6445 ( .A1(n4280), .A2(n5360), .ZN(n4646) );
  INV_X1 U6446 ( .A(n6681), .ZN(n4648) );
  OAI21_X1 U6447 ( .B1(n4650), .B2(n4648), .A(n4649), .ZN(n6696) );
  NAND2_X1 U6448 ( .A1(n6681), .A2(n4658), .ZN(n4657) );
  NAND2_X1 U6449 ( .A1(n8828), .A2(n4661), .ZN(n4660) );
  NAND2_X1 U6450 ( .A1(n6712), .A2(n8887), .ZN(n4670) );
  AND2_X1 U6451 ( .A1(n4670), .A2(n4673), .ZN(n8094) );
  OAI21_X1 U6452 ( .B1(n6735), .B2(n10188), .A(n4370), .ZN(n6736) );
  NAND2_X1 U6453 ( .A1(n9307), .A2(n4680), .ZN(n4679) );
  INV_X1 U6454 ( .A(n4697), .ZN(n9463) );
  NAND2_X1 U6455 ( .A1(n4702), .A2(n4700), .ZN(n6277) );
  NOR2_X2 U6456 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n4706) );
  NOR2_X2 U6457 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n4707) );
  NOR2_X2 U6458 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .ZN(
        n4708) );
  NOR2_X1 U6459 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n4709) );
  INV_X2 U6460 ( .A(n6574), .ZN(n6295) );
  NAND2_X2 U6461 ( .A1(n6484), .A2(n6827), .ZN(n6574) );
  NAND3_X1 U6462 ( .A1(n6828), .A2(n6827), .A3(n9505), .ZN(n5911) );
  NAND2_X2 U6463 ( .A1(n5839), .A2(n5838), .ZN(n6827) );
  XNOR2_X2 U6464 ( .A(n5841), .B(n5840), .ZN(n6484) );
  AND2_X2 U6465 ( .A1(n4714), .A2(n7929), .ZN(n7688) );
  NAND2_X1 U6466 ( .A1(n7655), .A2(n7924), .ZN(n7656) );
  INV_X1 U6467 ( .A(n4714), .ZN(n7687) );
  INV_X1 U6468 ( .A(n7924), .ZN(n4715) );
  INV_X1 U6469 ( .A(n8039), .ZN(n4724) );
  INV_X1 U6470 ( .A(n4734), .ZN(n9627) );
  NOR2_X1 U6471 ( .A1(n9627), .A2(n8046), .ZN(n9605) );
  NAND2_X1 U6472 ( .A1(n8164), .A2(n4748), .ZN(n4747) );
  INV_X1 U6473 ( .A(n7137), .ZN(n4750) );
  INV_X1 U6474 ( .A(n4756), .ZN(n7138) );
  INV_X1 U6475 ( .A(n8260), .ZN(n4765) );
  NAND2_X1 U6476 ( .A1(n8260), .A2(n4761), .ZN(n4759) );
  NAND2_X1 U6477 ( .A1(n8145), .A2(n4301), .ZN(n8144) );
  NAND3_X1 U6478 ( .A1(n4934), .A2(n4994), .A3(n4980), .ZN(n4776) );
  XNOR2_X1 U6479 ( .A(n5130), .B(n5572), .ZN(n8604) );
  XNOR2_X1 U6480 ( .A(n4777), .B(n4366), .ZN(n5132) );
  OAI21_X1 U6481 ( .B1(n8604), .B2(n4781), .A(n4778), .ZN(n4777) );
  INV_X1 U6482 ( .A(n5130), .ZN(n4780) );
  NAND2_X1 U6483 ( .A1(n7077), .A2(n4798), .ZN(n4789) );
  OAI21_X1 U6484 ( .B1(n7077), .B2(n4787), .A(n4785), .ZN(n4784) );
  NAND2_X1 U6485 ( .A1(n4795), .A2(n4796), .ZN(n4794) );
  INV_X1 U6486 ( .A(n4806), .ZN(n4801) );
  INV_X1 U6487 ( .A(n5129), .ZN(n4799) );
  OAI21_X1 U6488 ( .B1(n8540), .B2(n9021), .A(n4806), .ZN(n8554) );
  NAND2_X1 U6489 ( .A1(n4804), .A2(n8576), .ZN(n4803) );
  AND2_X1 U6490 ( .A1(n7030), .A2(n7031), .ZN(n7028) );
  AND2_X2 U6491 ( .A1(n7914), .A2(n7912), .ZN(n7373) );
  NAND2_X1 U6492 ( .A1(n7359), .A2(n7592), .ZN(n7912) );
  NAND2_X1 U6493 ( .A1(n7358), .A2(n10104), .ZN(n7914) );
  INV_X2 U6494 ( .A(n7359), .ZN(n7358) );
  NAND2_X1 U6495 ( .A1(n9743), .A2(n4347), .ZN(n4814) );
  NAND2_X1 U6496 ( .A1(n4814), .A2(n4813), .ZN(n8064) );
  NAND2_X1 U6497 ( .A1(n9622), .A2(n4829), .ZN(n4828) );
  OR2_X1 U6498 ( .A1(n9622), .A2(n8075), .ZN(n4834) );
  INV_X1 U6499 ( .A(n4842), .ZN(n8073) );
  NAND2_X1 U6500 ( .A1(n7684), .A2(n4348), .ZN(n4856) );
  NAND2_X1 U6501 ( .A1(n4856), .A2(n4857), .ZN(n8058) );
  NAND2_X1 U6502 ( .A1(n8004), .A2(n7877), .ZN(n4864) );
  NAND2_X1 U6503 ( .A1(n4871), .A2(n5276), .ZN(n5471) );
  NAND2_X2 U6504 ( .A1(n5459), .A2(n5458), .ZN(n4871) );
  INV_X2 U6505 ( .A(n7903), .ZN(n7370) );
  NAND3_X2 U6506 ( .A1(n5912), .A2(n5911), .A3(n5910), .ZN(n7903) );
  INV_X1 U6507 ( .A(n4895), .ZN(n9764) );
  INV_X1 U6508 ( .A(n4898), .ZN(n9690) );
  OR3_X1 U6509 ( .A1(n9660), .A2(n9796), .A3(n4901), .ZN(n9612) );
  NAND3_X1 U6510 ( .A1(n4900), .A2(n9619), .A3(n9599), .ZN(n4899) );
  AOI21_X1 U6511 ( .B1(n4911), .B2(n8315), .A(n8321), .ZN(n8326) );
  INV_X1 U6512 ( .A(n8313), .ZN(n4912) );
  NAND2_X1 U6513 ( .A1(n4923), .A2(n4921), .ZN(n8378) );
  INV_X1 U6514 ( .A(n4922), .ZN(n4921) );
  OAI21_X1 U6515 ( .B1(n8373), .B2(n4330), .A(n8792), .ZN(n4922) );
  NAND3_X1 U6516 ( .A1(n8360), .A2(n4925), .A3(n4924), .ZN(n4923) );
  INV_X1 U6517 ( .A(n8373), .ZN(n4924) );
  INV_X1 U6518 ( .A(n6969), .ZN(n7019) );
  NAND2_X1 U6519 ( .A1(n4936), .A2(n4935), .ZN(n6969) );
  OR2_X1 U6520 ( .A1(n5794), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n4936) );
  OAI21_X1 U6521 ( .B1(n7125), .B2(n4941), .A(n4940), .ZN(n7194) );
  AOI21_X1 U6522 ( .B1(n6622), .B2(n8307), .A(n4944), .ZN(n4940) );
  INV_X1 U6523 ( .A(n6622), .ZN(n4941) );
  OAI211_X1 U6524 ( .C1(n4944), .C2(n6622), .A(n4942), .B(n8317), .ZN(n6623)
         );
  NAND2_X1 U6525 ( .A1(n7125), .A2(n4943), .ZN(n4942) );
  AND2_X1 U6526 ( .A1(n8306), .A2(n8312), .ZN(n4943) );
  INV_X1 U6527 ( .A(n8391), .ZN(n4948) );
  NAND3_X1 U6528 ( .A1(n8390), .A2(n4951), .A3(n8799), .ZN(n4950) );
  AOI21_X2 U6529 ( .B1(n8653), .B2(n6641), .A(n4325), .ZN(n8465) );
  INV_X1 U6530 ( .A(n8484), .ZN(n6620) );
  NAND2_X2 U6531 ( .A1(n8299), .A2(n8298), .ZN(n8484) );
  NAND2_X2 U6532 ( .A1(n4967), .A2(n7103), .ZN(n8299) );
  AND2_X1 U6533 ( .A1(n6630), .A2(n6629), .ZN(n4968) );
  NAND2_X1 U6534 ( .A1(n7595), .A2(n7597), .ZN(n4969) );
  AND2_X2 U6535 ( .A1(n4999), .A2(n4970), .ZN(n5212) );
  NAND2_X1 U6536 ( .A1(n4999), .A2(n4971), .ZN(n5208) );
  AND2_X1 U6537 ( .A1(n5364), .A2(n4967), .ZN(n5365) );
  CLKBUF_X1 U6538 ( .A(n6201), .Z(n6260) );
  INV_X1 U6539 ( .A(n6025), .ZN(n6028) );
  OAI211_X1 U6540 ( .C1(n8702), .C2(n8905), .A(n8701), .B(n8700), .ZN(n9175)
         );
  NAND2_X1 U6541 ( .A1(n5896), .A2(n7886), .ZN(n8015) );
  AOI21_X1 U6542 ( .B1(n8691), .B2(n8887), .A(n8690), .ZN(n9169) );
  XNOR2_X1 U6543 ( .A(n8685), .B(n8684), .ZN(n8691) );
  NAND2_X1 U6544 ( .A1(n6876), .A2(n6878), .ZN(n6877) );
  AOI21_X1 U6545 ( .B1(n8677), .B2(n8887), .A(n8676), .ZN(n9163) );
  XNOR2_X1 U6546 ( .A(n8672), .B(n8671), .ZN(n8677) );
  INV_X4 U6547 ( .A(n6000), .ZN(n9335) );
  OR2_X1 U6548 ( .A1(n5991), .A2(n5953), .ZN(n5954) );
  INV_X1 U6549 ( .A(n9790), .ZN(n9791) );
  NOR2_X2 U6550 ( .A1(n5904), .A2(n5870), .ZN(n5871) );
  CLKBUF_X1 U6551 ( .A(n9748), .Z(n9768) );
  INV_X1 U6552 ( .A(n7969), .ZN(n7615) );
  NAND2_X1 U6553 ( .A1(n9781), .A2(n10145), .ZN(n6571) );
  NAND2_X1 U6554 ( .A1(n9582), .A2(n6565), .ZN(n9781) );
  NAND2_X1 U6555 ( .A1(n9782), .A2(n10145), .ZN(n6617) );
  NAND2_X1 U6556 ( .A1(n5711), .A2(n5710), .ZN(n5713) );
  NAND2_X1 U6557 ( .A1(n7780), .A2(n6615), .ZN(n9782) );
  NAND2_X1 U6558 ( .A1(n5385), .A2(n4339), .ZN(n5393) );
  OR2_X1 U6559 ( .A1(n5385), .A2(n4339), .ZN(n5386) );
  INV_X2 U6560 ( .A(n4441), .ZN(n7348) );
  OAI21_X1 U6561 ( .B1(n6479), .B2(n9352), .A(n9474), .ZN(n6508) );
  NAND2_X1 U6562 ( .A1(n5512), .A2(n5511), .ZN(n5515) );
  NAND2_X1 U6563 ( .A1(n5512), .A2(n5500), .ZN(n6842) );
  INV_X1 U6564 ( .A(n9800), .ZN(n9626) );
  INV_X1 U6565 ( .A(n9460), .ZN(n9465) );
  OAI21_X1 U6566 ( .B1(n9460), .B2(n6456), .A(n6455), .ZN(n6454) );
  OAI21_X1 U6567 ( .B1(n5212), .B2(n5023), .A(P2_IR_REG_29__SCAN_IN), .ZN(
        n5214) );
  NAND2_X1 U6568 ( .A1(n9603), .A2(n10013), .ZN(n9611) );
  INV_X1 U6569 ( .A(n9814), .ZN(n9679) );
  INV_X1 U6570 ( .A(n9273), .ZN(n5218) );
  OAI21_X1 U6571 ( .B1(n9584), .B2(n9586), .A(n9583), .ZN(n9793) );
  OR2_X1 U6572 ( .A1(n6786), .A2(n6161), .ZN(n6011) );
  OR2_X1 U6573 ( .A1(n5986), .A2(n6161), .ZN(n5990) );
  OR2_X1 U6574 ( .A1(n6782), .A2(n6161), .ZN(n5971) );
  NAND2_X2 U6576 ( .A1(n6339), .A2(n6338), .ZN(n9824) );
  CLKBUF_X1 U6577 ( .A(n7386), .Z(n8859) );
  INV_X1 U6578 ( .A(n7887), .ZN(n8038) );
  INV_X1 U6579 ( .A(n9888), .ZN(n5887) );
  OR2_X1 U6580 ( .A1(n5072), .A2(n4796), .ZN(n4972) );
  NOR3_X1 U6581 ( .A1(n9624), .A2(n9623), .A3(n10039), .ZN(n4973) );
  AND2_X2 U6582 ( .A1(n6995), .A2(n6569), .ZN(n10145) );
  AND2_X2 U6583 ( .A1(n6725), .A2(n7011), .ZN(n9003) );
  INV_X1 U6584 ( .A(n9425), .ZN(n9492) );
  OR2_X1 U6585 ( .A1(n8089), .A2(n9264), .ZN(n4974) );
  OR2_X1 U6586 ( .A1(n8089), .A2(n8996), .ZN(n4976) );
  AND2_X1 U6587 ( .A1(n9788), .A2(n9858), .ZN(n4978) );
  OR2_X1 U6588 ( .A1(n9591), .A2(n10048), .ZN(n4982) );
  OR2_X1 U6589 ( .A1(n10062), .A2(n6478), .ZN(n10139) );
  INV_X1 U6590 ( .A(n5239), .ZN(n5354) );
  OAI211_X1 U6591 ( .C1(n5609), .C2(P1_DATAO_REG_0__SCAN_IN), .A(SI_0_), .B(
        n5238), .ZN(n5239) );
  INV_X1 U6592 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n5245) );
  INV_X1 U6593 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n5249) );
  INV_X1 U6594 ( .A(n9581), .ZN(n10031) );
  INV_X1 U6595 ( .A(n8841), .ZN(n6630) );
  INV_X1 U6596 ( .A(n6294), .ZN(n6602) );
  AND2_X2 U6597 ( .A1(n7379), .A2(n10068), .ZN(n4984) );
  OR2_X1 U6598 ( .A1(n7352), .A2(n10086), .ZN(n4985) );
  INV_X1 U6599 ( .A(n8085), .ZN(n9784) );
  INV_X1 U6600 ( .A(n9824), .ZN(n8063) );
  AND2_X1 U6601 ( .A1(n6686), .A2(n8178), .ZN(n4986) );
  INV_X1 U6602 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n4993) );
  NOR2_X1 U6603 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n5823) );
  AND2_X1 U6604 ( .A1(n8743), .A2(n8744), .ZN(n6673) );
  INV_X1 U6605 ( .A(n9686), .ZN(n8062) );
  NAND2_X1 U6606 ( .A1(n5053), .A2(n5052), .ZN(n5055) );
  NAND2_X1 U6607 ( .A1(n7637), .A2(n7960), .ZN(n7371) );
  INV_X1 U6608 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n5273) );
  NAND2_X1 U6609 ( .A1(n5609), .A2(n5241), .ZN(n5242) );
  OR2_X1 U6610 ( .A1(n5425), .A2(n7390), .ZN(n5426) );
  AND2_X1 U6611 ( .A1(n6694), .A2(n6693), .ZN(n6695) );
  AND2_X1 U6612 ( .A1(n5771), .A2(n6797), .ZN(n7007) );
  NAND2_X1 U6613 ( .A1(n8875), .A2(n8889), .ZN(n6660) );
  INV_X1 U6614 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5018) );
  INV_X1 U6615 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n6096) );
  AND2_X1 U6616 ( .A1(n9752), .A2(n7994), .ZN(n7995) );
  INV_X1 U6617 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5840) );
  INV_X1 U6618 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n5856) );
  INV_X1 U6619 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n5845) );
  NAND2_X1 U6620 ( .A1(n7261), .A2(n5426), .ZN(n7451) );
  NAND2_X1 U6621 ( .A1(n5360), .A2(n6779), .ZN(n5387) );
  OR2_X1 U6622 ( .A1(n6722), .A2(n4743), .ZN(n6724) );
  NAND2_X1 U6623 ( .A1(n8686), .A2(n8890), .ZN(n8657) );
  NAND3_X2 U6624 ( .A1(n7420), .A2(n5902), .A3(n6738), .ZN(n5938) );
  INV_X1 U6625 ( .A(n9462), .ZN(n6430) );
  INV_X1 U6626 ( .A(n5939), .ZN(n5940) );
  INV_X1 U6627 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n6235) );
  INV_X1 U6628 ( .A(n9488), .ZN(n9607) );
  NAND2_X1 U6629 ( .A1(n6525), .A2(n6524), .ZN(n6536) );
  NAND2_X1 U6630 ( .A1(n5300), .A2(SI_18_), .ZN(n5301) );
  AND2_X1 U6631 ( .A1(n5804), .A2(n6732), .ZN(n8283) );
  NAND2_X1 U6632 ( .A1(n8250), .A2(n5666), .ZN(n8205) );
  INV_X1 U6633 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5020) );
  INV_X1 U6634 ( .A(n8757), .ZN(n8779) );
  INV_X1 U6635 ( .A(n8673), .ZN(n8470) );
  INV_X1 U6636 ( .A(n7396), .ZN(n8998) );
  NAND2_X1 U6637 ( .A1(n6431), .A2(n6430), .ZN(n6432) );
  NAND2_X1 U6638 ( .A1(n6028), .A2(n6027), .ZN(n7313) );
  OR2_X1 U6639 ( .A1(n6502), .A2(n6501), .ZN(n9454) );
  OR2_X1 U6640 ( .A1(n9615), .A2(n6442), .ZN(n6447) );
  INV_X1 U6641 ( .A(n6442), .ZN(n7243) );
  NOR2_X1 U6642 ( .A1(n6581), .A2(n9912), .ZN(n9931) );
  INV_X1 U6643 ( .A(n9796), .ZN(n9619) );
  INV_X1 U6644 ( .A(n9804), .ZN(n9650) );
  AND2_X1 U6645 ( .A1(n7823), .A2(n7820), .ZN(n7965) );
  OAI21_X1 U6646 ( .B1(n7946), .B2(n10139), .A(n7777), .ZN(n6564) );
  INV_X1 U6647 ( .A(n10139), .ZN(n9858) );
  INV_X1 U6648 ( .A(n7709), .ZN(n6457) );
  AND2_X1 U6649 ( .A1(n5675), .A2(n5674), .ZN(n5699) );
  OAI21_X1 U6650 ( .B1(n5281), .B2(SI_12_), .A(n5511), .ZN(n5498) );
  XNOR2_X1 U6651 ( .A(n5272), .B(SI_8_), .ZN(n5452) );
  OAI21_X1 U6652 ( .B1(n6689), .B2(n8291), .A(n5819), .ZN(n5820) );
  INV_X1 U6653 ( .A(n8285), .ZN(n8264) );
  OR2_X1 U6654 ( .A1(n8182), .A2(n8280), .ZN(n8281) );
  INV_X1 U6655 ( .A(n8634), .ZN(n8611) );
  NAND2_X1 U6656 ( .A1(n6703), .A2(n8469), .ZN(n8887) );
  NAND2_X1 U6657 ( .A1(n4269), .A2(n8929), .ZN(n8930) );
  NOR2_X1 U6658 ( .A1(n8648), .A2(n8647), .ZN(n9150) );
  AND2_X1 U6659 ( .A1(n8715), .A2(n8473), .ZN(n8723) );
  AND2_X1 U6660 ( .A1(n8894), .A2(n7397), .ZN(n7596) );
  INV_X1 U6661 ( .A(n7596), .ZN(n8999) );
  INV_X1 U6662 ( .A(n7397), .ZN(n8993) );
  AND2_X1 U6663 ( .A1(n6499), .A2(n8021), .ZN(n9479) );
  INV_X1 U6664 ( .A(n9485), .ZN(n9444) );
  INV_X1 U6665 ( .A(n9454), .ZN(n9482) );
  OAI21_X1 U6666 ( .B1(n7989), .B2(n7985), .A(n5896), .ZN(n7887) );
  OR2_X1 U6667 ( .A1(n9646), .A2(n6442), .ZN(n6407) );
  INV_X1 U6668 ( .A(n9928), .ZN(n9957) );
  AND2_X1 U6669 ( .A1(n6605), .A2(n6606), .ZN(n6832) );
  INV_X1 U6670 ( .A(n9948), .ZN(n9959) );
  OAI21_X1 U6671 ( .B1(n9970), .B2(n5226), .A(n9328), .ZN(n6608) );
  AND2_X1 U6672 ( .A1(n8044), .A2(n7894), .ZN(n9655) );
  AND2_X1 U6673 ( .A1(n7955), .A2(n7996), .ZN(n9752) );
  AND2_X1 U6674 ( .A1(n10070), .A2(n7421), .ZN(n10032) );
  INV_X1 U6675 ( .A(n6564), .ZN(n6565) );
  AOI21_X1 U6676 ( .B1(n6817), .B2(n6463), .A(n6821), .ZN(n7365) );
  INV_X1 U6677 ( .A(n10136), .ZN(n9861) );
  NOR2_X1 U6678 ( .A1(n6568), .A2(n7366), .ZN(n6995) );
  INV_X1 U6679 ( .A(n8216), .ZN(n8279) );
  INV_X1 U6680 ( .A(n8276), .ZN(n8291) );
  INV_X1 U6681 ( .A(n8768), .ZN(n8793) );
  INV_X1 U6682 ( .A(n7445), .ZN(n7553) );
  NAND2_X1 U6683 ( .A1(n10171), .A2(n7124), .ZN(n8855) );
  INV_X1 U6684 ( .A(n10171), .ZN(n10174) );
  NAND2_X1 U6685 ( .A1(n8931), .A2(n8930), .ZN(n8933) );
  NAND2_X1 U6686 ( .A1(n9003), .A2(n8999), .ZN(n8985) );
  XOR2_X1 U6688 ( .A(n8655), .B(n8653), .Z(n9162) );
  OR2_X1 U6689 ( .A1(n10188), .A2(n7596), .ZN(n9255) );
  AND2_X1 U6690 ( .A1(n6734), .A2(n6733), .ZN(n10188) );
  AND2_X1 U6691 ( .A1(n5809), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6802) );
  INV_X1 U6692 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n8096) );
  INV_X1 U6693 ( .A(n6506), .ZN(n6507) );
  AND2_X1 U6694 ( .A1(n6483), .A2(n10068), .ZN(n9485) );
  INV_X1 U6695 ( .A(n9631), .ZN(n9590) );
  INV_X1 U6696 ( .A(n9717), .ZN(n9754) );
  INV_X1 U6697 ( .A(n9974), .ZN(n9497) );
  INV_X1 U6698 ( .A(n10032), .ZN(n9780) );
  AND2_X2 U6699 ( .A1(n6995), .A2(n7365), .ZN(n10162) );
  OAI211_X1 U6700 ( .C1(n9793), .C2(n9861), .A(n9792), .B(n9791), .ZN(n9864)
         );
  INV_X1 U6701 ( .A(n10145), .ZN(n10144) );
  AND2_X1 U6702 ( .A1(n6819), .A2(n6818), .ZN(n10076) );
  NAND2_X1 U6703 ( .A1(n5332), .A2(n5412), .ZN(n6786) );
  AND2_X1 U6704 ( .A1(n5011), .A2(n6802), .ZN(P2_U3893) );
  INV_X1 U6705 ( .A(n9501), .ZN(P1_U3973) );
  NAND2_X1 U6706 ( .A1(n6571), .A2(n6570), .ZN(P1_U3521) );
  INV_X1 U6707 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n4989) );
  INV_X1 U6708 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n4988) );
  NAND4_X1 U6709 ( .A1(n4992), .A2(n4991), .A3(n4990), .A4(n5028), .ZN(n5007)
         );
  INV_X1 U6710 ( .A(n5007), .ZN(n4994) );
  NAND2_X1 U6711 ( .A1(n5026), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4996) );
  OR2_X1 U6712 ( .A1(n4996), .A2(n5019), .ZN(n4998) );
  NAND2_X1 U6713 ( .A1(n4996), .A2(n5019), .ZN(n4997) );
  INV_X1 U6714 ( .A(n4999), .ZN(n5003) );
  NAND2_X1 U6715 ( .A1(n5003), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5001) );
  XNOR2_X1 U6716 ( .A(n5001), .B(n5000), .ZN(n7712) );
  INV_X1 U6717 ( .A(n7712), .ZN(n5006) );
  MUX2_X1 U6718 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5002), .S(
        P2_IR_REG_24__SCAN_IN), .Z(n5004) );
  NAND2_X1 U6719 ( .A1(n5004), .A2(n5003), .ZN(n5313) );
  INV_X1 U6720 ( .A(n5313), .ZN(n5005) );
  NAND3_X1 U6721 ( .A1(n5316), .A2(n5006), .A3(n5005), .ZN(n5808) );
  INV_X1 U6722 ( .A(n5808), .ZN(n5011) );
  OR2_X1 U6723 ( .A1(n5079), .A2(n5007), .ZN(n5309) );
  NAND2_X1 U6724 ( .A1(n5014), .A2(n5008), .ZN(n5012) );
  OAI21_X1 U6725 ( .B1(n5012), .B2(P2_IR_REG_22__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5010) );
  XNOR2_X1 U6726 ( .A(n5010), .B(n5009), .ZN(n5809) );
  INV_X1 U6727 ( .A(n5809), .ZN(n7611) );
  OR2_X1 U6728 ( .A1(n5808), .A2(n7611), .ZN(n5189) );
  NAND2_X1 U6729 ( .A1(n5012), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5013) );
  INV_X1 U6730 ( .A(n5014), .ZN(n5015) );
  NAND2_X1 U6731 ( .A1(n5015), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5016) );
  NAND2_X1 U6732 ( .A1(n8440), .A2(n5809), .ZN(n5017) );
  NAND2_X1 U6733 ( .A1(n5189), .A2(n5017), .ZN(n5192) );
  NAND2_X1 U6734 ( .A1(n5208), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5021) );
  AND2_X1 U6735 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), .ZN(
        n5025) );
  NAND2_X1 U6736 ( .A1(P2_IR_REG_26__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), 
        .ZN(n5022) );
  AOI22_X1 U6737 ( .A1(P2_IR_REG_27__SCAN_IN), .A2(n5023), .B1(n5022), .B2(
        P2_IR_REG_31__SCAN_IN), .ZN(n5024) );
  NAND2_X2 U6738 ( .A1(n5190), .A2(n9285), .ZN(n5360) );
  OAI21_X1 U6739 ( .B1(n5192), .B2(n6710), .A(P2_STATE_REG_SCAN_IN), .ZN(
        P2_U3150) );
  INV_X1 U6740 ( .A(n5028), .ZN(n5029) );
  NOR2_X1 U6741 ( .A1(n5029), .A2(P2_IR_REG_15__SCAN_IN), .ZN(n5030) );
  NAND2_X1 U6742 ( .A1(n5087), .A2(n5030), .ZN(n5032) );
  NAND2_X1 U6743 ( .A1(n5032), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5031) );
  MUX2_X1 U6744 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5031), .S(
        P2_IR_REG_16__SCAN_IN), .Z(n5033) );
  AND2_X1 U6745 ( .A1(n5033), .A2(n5103), .ZN(n5560) );
  INV_X1 U6746 ( .A(n5560), .ZN(n8589) );
  NAND2_X1 U6747 ( .A1(n5035), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5036) );
  INV_X1 U6748 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n5134) );
  NAND2_X1 U6749 ( .A1(n6869), .A2(n4308), .ZN(n6857) );
  INV_X1 U6750 ( .A(n5034), .ZN(n5038) );
  INV_X1 U6751 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n10173) );
  XNOR2_X1 U6752 ( .A(n6851), .B(n10173), .ZN(n6858) );
  NAND2_X1 U6753 ( .A1(n6857), .A2(n6858), .ZN(n6856) );
  NAND2_X1 U6754 ( .A1(n6851), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n5040) );
  NAND2_X1 U6755 ( .A1(n6856), .A2(n5040), .ZN(n5044) );
  NAND2_X1 U6756 ( .A1(n5042), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5041) );
  MUX2_X1 U6757 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5041), .S(
        P2_IR_REG_3__SCAN_IN), .Z(n5043) );
  NAND2_X1 U6758 ( .A1(n5044), .A2(n7068), .ZN(n7033) );
  OR2_X1 U6759 ( .A1(n5044), .A2(n7068), .ZN(n5045) );
  AND2_X1 U6760 ( .A1(n7033), .A2(n5045), .ZN(n7067) );
  NAND2_X1 U6761 ( .A1(n5076), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5046) );
  XNOR2_X2 U6762 ( .A(n5046), .B(n5048), .ZN(n7037) );
  INV_X1 U6763 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n7217) );
  XNOR2_X1 U6764 ( .A(n7037), .B(n7217), .ZN(n7032) );
  NAND2_X1 U6765 ( .A1(n7037), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5047) );
  INV_X1 U6766 ( .A(n5054), .ZN(n5053) );
  INV_X1 U6767 ( .A(n5076), .ZN(n5049) );
  NAND2_X1 U6768 ( .A1(n5049), .A2(n5048), .ZN(n5056) );
  NAND2_X1 U6769 ( .A1(n5056), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5051) );
  INV_X1 U6770 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5050) );
  XNOR2_X1 U6771 ( .A(n5051), .B(n5050), .ZN(n6785) );
  INV_X1 U6772 ( .A(n6785), .ZN(n5052) );
  NAND2_X1 U6773 ( .A1(n5054), .A2(n6785), .ZN(n6891) );
  NAND2_X1 U6774 ( .A1(n5059), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5057) );
  XNOR2_X1 U6775 ( .A(n6804), .B(P2_REG2_REG_6__SCAN_IN), .ZN(n6890) );
  INV_X1 U6776 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n7338) );
  OR2_X1 U6777 ( .A1(n6804), .A2(n7338), .ZN(n5058) );
  NAND2_X1 U6778 ( .A1(n6894), .A2(n5058), .ZN(n5066) );
  INV_X1 U6779 ( .A(n5059), .ZN(n5061) );
  INV_X1 U6780 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5060) );
  NAND2_X1 U6781 ( .A1(n5061), .A2(n5060), .ZN(n5063) );
  NAND2_X1 U6782 ( .A1(n5063), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5062) );
  MUX2_X1 U6783 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5062), .S(
        P2_IR_REG_7__SCAN_IN), .Z(n5064) );
  NAND2_X1 U6784 ( .A1(n5064), .A2(n5070), .ZN(n6791) );
  INV_X1 U6785 ( .A(n6791), .ZN(n5065) );
  NAND2_X1 U6786 ( .A1(n7053), .A2(n7088), .ZN(n5068) );
  NAND2_X1 U6787 ( .A1(n5070), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5067) );
  XNOR2_X1 U6788 ( .A(n5454), .B(P2_REG2_REG_8__SCAN_IN), .ZN(n7087) );
  NAND2_X1 U6789 ( .A1(n5068), .A2(n7087), .ZN(n7091) );
  INV_X1 U6790 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n8918) );
  OR2_X1 U6791 ( .A1(n5454), .A2(n8918), .ZN(n5069) );
  NAND2_X1 U6792 ( .A1(n7091), .A2(n5069), .ZN(n5072) );
  OAI21_X1 U6793 ( .B1(n5070), .B2(n9109), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n5071) );
  XNOR2_X1 U6794 ( .A(n5071), .B(P2_IR_REG_9__SCAN_IN), .ZN(n5460) );
  NAND2_X2 U6795 ( .A1(n7204), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n7203) );
  BUF_X1 U6796 ( .A(n5073), .Z(n5074) );
  INV_X1 U6797 ( .A(n5074), .ZN(n5075) );
  OAI21_X1 U6798 ( .B1(n5076), .B2(n5075), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n5077) );
  XNOR2_X1 U6799 ( .A(n5077), .B(P2_IR_REG_10__SCAN_IN), .ZN(n5474) );
  XNOR2_X1 U6800 ( .A(n5474), .B(P2_REG2_REG_10__SCAN_IN), .ZN(n7281) );
  INV_X1 U6801 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n8873) );
  OR2_X1 U6802 ( .A1(n5474), .A2(n8873), .ZN(n5078) );
  NAND2_X1 U6803 ( .A1(n5079), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5080) );
  XNOR2_X1 U6804 ( .A(n5080), .B(P2_IR_REG_11__SCAN_IN), .ZN(n5495) );
  INV_X1 U6805 ( .A(n5495), .ZN(n7477) );
  NAND2_X1 U6806 ( .A1(n5082), .A2(n7477), .ZN(n7529) );
  NAND2_X1 U6807 ( .A1(n5084), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5085) );
  XNOR2_X1 U6808 ( .A(n5085), .B(P2_IR_REG_12__SCAN_IN), .ZN(n5501) );
  XNOR2_X1 U6809 ( .A(n5501), .B(P2_REG2_REG_12__SCAN_IN), .ZN(n7530) );
  INV_X1 U6810 ( .A(n5501), .ZN(n7521) );
  NAND2_X1 U6811 ( .A1(n7521), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n5086) );
  NAND2_X1 U6812 ( .A1(n7533), .A2(n5086), .ZN(n5089) );
  INV_X1 U6813 ( .A(n5087), .ZN(n5088) );
  NAND2_X1 U6814 ( .A1(n5088), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5091) );
  XNOR2_X1 U6815 ( .A(n5091), .B(P2_IR_REG_13__SCAN_IN), .ZN(n5516) );
  INV_X1 U6816 ( .A(n5516), .ZN(n8544) );
  INV_X1 U6817 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n8837) );
  INV_X1 U6818 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5090) );
  NAND2_X1 U6819 ( .A1(n5091), .A2(n5090), .ZN(n5092) );
  NAND2_X1 U6820 ( .A1(n5092), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5094) );
  INV_X1 U6821 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5093) );
  NAND2_X1 U6822 ( .A1(n5094), .A2(n5093), .ZN(n5097) );
  OR2_X1 U6823 ( .A1(n5094), .A2(n5093), .ZN(n5095) );
  XNOR2_X1 U6824 ( .A(n5532), .B(P2_REG2_REG_14__SCAN_IN), .ZN(n8566) );
  INV_X1 U6825 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n8825) );
  OR2_X1 U6826 ( .A1(n5532), .A2(n8825), .ZN(n5096) );
  NAND2_X1 U6827 ( .A1(n5097), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5098) );
  XNOR2_X1 U6828 ( .A(n5098), .B(P2_IR_REG_15__SCAN_IN), .ZN(n5553) );
  NOR2_X1 U6829 ( .A1(n5099), .A2(n5553), .ZN(n5100) );
  INV_X1 U6830 ( .A(n5100), .ZN(n8597) );
  INV_X1 U6831 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8804) );
  XNOR2_X1 U6832 ( .A(n5560), .B(n8804), .ZN(n8598) );
  NAND2_X1 U6833 ( .A1(n5103), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5101) );
  XNOR2_X1 U6834 ( .A(n5101), .B(P2_IR_REG_17__SCAN_IN), .ZN(n5572) );
  INV_X1 U6835 ( .A(n5102), .ZN(n8639) );
  OAI21_X2 U6836 ( .B1(n5103), .B2(P2_IR_REG_17__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5105) );
  INV_X1 U6837 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5104) );
  NAND2_X1 U6838 ( .A1(n5105), .A2(n5104), .ZN(n5109) );
  OR2_X1 U6839 ( .A1(n5105), .A2(n5104), .ZN(n5106) );
  AND2_X1 U6840 ( .A1(n5109), .A2(n5106), .ZN(n5586) );
  INV_X1 U6841 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n5181) );
  OR2_X1 U6842 ( .A1(n5586), .A2(n5181), .ZN(n5108) );
  NAND2_X1 U6843 ( .A1(n5586), .A2(n5181), .ZN(n5107) );
  NAND2_X1 U6844 ( .A1(n5108), .A2(n5107), .ZN(n8638) );
  NAND2_X1 U6845 ( .A1(n5109), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5111) );
  INV_X1 U6846 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5110) );
  XNOR2_X1 U6847 ( .A(n4274), .B(P2_REG2_REG_19__SCAN_IN), .ZN(n5186) );
  INV_X1 U6848 ( .A(n5192), .ZN(n5112) );
  NAND2_X1 U6849 ( .A1(n5112), .A2(n4364), .ZN(n5131) );
  INV_X1 U6850 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n5126) );
  INV_X1 U6851 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n9137) );
  INV_X1 U6852 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n5113) );
  INV_X1 U6853 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n5133) );
  OR2_X1 U6854 ( .A1(n5034), .A2(n5133), .ZN(n5116) );
  NAND3_X1 U6855 ( .A1(n5034), .A2(P2_REG1_REG_0__SCAN_IN), .A3(n5035), .ZN(
        n5114) );
  NAND2_X1 U6856 ( .A1(n5115), .A2(n5114), .ZN(n6868) );
  NAND2_X1 U6857 ( .A1(n6868), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5117) );
  NAND2_X1 U6858 ( .A1(n5117), .A2(n5116), .ZN(n6854) );
  NAND2_X1 U6859 ( .A1(n6851), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5118) );
  INV_X1 U6860 ( .A(n7068), .ZN(n5119) );
  NAND2_X1 U6861 ( .A1(n5120), .A2(n7068), .ZN(n5121) );
  INV_X1 U6862 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n5123) );
  MUX2_X1 U6863 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n5123), .S(n7037), .Z(n7031)
         );
  INV_X1 U6864 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n5125) );
  OAI22_X1 U6865 ( .A1(n6985), .A2(n5125), .B1(n5052), .B2(n5124), .ZN(n6888)
         );
  MUX2_X1 U6866 ( .A(n9137), .B(P2_REG1_REG_6__SCAN_IN), .S(n6804), .Z(n6889)
         );
  MUX2_X1 U6867 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n5126), .S(n5454), .Z(n7080)
         );
  XOR2_X1 U6868 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n5474), .Z(n7271) );
  INV_X1 U6869 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n9024) );
  INV_X1 U6870 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n7602) );
  INV_X1 U6871 ( .A(n5127), .ZN(n5128) );
  OAI22_X1 U6872 ( .A1(n7474), .A2(n7602), .B1(n5495), .B2(n5128), .ZN(n7519)
         );
  XNOR2_X1 U6873 ( .A(n5501), .B(P2_REG1_REG_12__SCAN_IN), .ZN(n7520) );
  XNOR2_X1 U6874 ( .A(n5129), .B(n5516), .ZN(n8540) );
  INV_X1 U6875 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n9021) );
  XNOR2_X1 U6876 ( .A(n5532), .B(P2_REG1_REG_14__SCAN_IN), .ZN(n8555) );
  INV_X1 U6877 ( .A(n5532), .ZN(n8557) );
  INV_X1 U6878 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n8973) );
  XNOR2_X1 U6879 ( .A(n5560), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n8587) );
  INV_X1 U6880 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n8967) );
  XNOR2_X1 U6881 ( .A(n5586), .B(P2_REG1_REG_18__SCAN_IN), .ZN(n8622) );
  INV_X1 U6882 ( .A(n5586), .ZN(n8629) );
  INV_X1 U6883 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n8960) );
  INV_X1 U6884 ( .A(n5131), .ZN(n6845) );
  NAND2_X1 U6885 ( .A1(n6845), .A2(n4270), .ZN(n8645) );
  MUX2_X1 U6886 ( .A(P2_REG2_REG_17__SCAN_IN), .B(P2_REG1_REG_17__SCAN_IN), 
        .S(n4271), .Z(n5180) );
  INV_X1 U6887 ( .A(n5572), .ZN(n8614) );
  MUX2_X1 U6888 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n4270), .Z(n5140) );
  XNOR2_X1 U6889 ( .A(n5135), .B(n5359), .ZN(n6865) );
  MUX2_X1 U6890 ( .A(n5134), .B(n5133), .S(n4271), .Z(n6843) );
  NAND2_X1 U6891 ( .A1(n6843), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n6864) );
  AOI22_X1 U6892 ( .A1(n6865), .A2(n6864), .B1(n5135), .B2(n6866), .ZN(n6850)
         );
  MUX2_X1 U6893 ( .A(P2_REG2_REG_2__SCAN_IN), .B(P2_REG1_REG_2__SCAN_IN), .S(
        n4270), .Z(n5136) );
  XNOR2_X1 U6894 ( .A(n5136), .B(n6851), .ZN(n6849) );
  INV_X1 U6895 ( .A(n6851), .ZN(n5138) );
  INV_X1 U6896 ( .A(n5136), .ZN(n5137) );
  MUX2_X1 U6897 ( .A(P2_REG2_REG_3__SCAN_IN), .B(P2_REG1_REG_3__SCAN_IN), .S(
        n4270), .Z(n5139) );
  XNOR2_X1 U6898 ( .A(n5139), .B(n7068), .ZN(n7064) );
  NOR2_X1 U6899 ( .A1(n5139), .A2(n7068), .ZN(n7025) );
  XNOR2_X1 U6900 ( .A(n5140), .B(n7037), .ZN(n7024) );
  AOI21_X1 U6901 ( .B1(n5140), .B2(n7037), .A(n7023), .ZN(n6984) );
  MUX2_X1 U6902 ( .A(P2_REG2_REG_5__SCAN_IN), .B(P2_REG1_REG_5__SCAN_IN), .S(
        n4271), .Z(n5141) );
  XNOR2_X1 U6903 ( .A(n5141), .B(n6785), .ZN(n6983) );
  INV_X1 U6904 ( .A(n5141), .ZN(n5142) );
  OAI22_X1 U6905 ( .A1(n6984), .A2(n6983), .B1(n5052), .B2(n5142), .ZN(n6886)
         );
  MUX2_X1 U6906 ( .A(n7338), .B(n9137), .S(n4270), .Z(n5143) );
  NAND2_X1 U6907 ( .A1(n5143), .A2(n6804), .ZN(n5144) );
  OAI21_X1 U6908 ( .B1(n5143), .B2(n6804), .A(n5144), .ZN(n6885) );
  INV_X1 U6909 ( .A(n5144), .ZN(n7049) );
  INV_X1 U6910 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n9074) );
  INV_X1 U6911 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n7046) );
  MUX2_X1 U6912 ( .A(n9074), .B(n7046), .S(n4271), .Z(n5145) );
  NAND2_X1 U6913 ( .A1(n5145), .A2(n5065), .ZN(n7082) );
  INV_X1 U6914 ( .A(n5145), .ZN(n5146) );
  NAND2_X1 U6915 ( .A1(n5146), .A2(n6791), .ZN(n5147) );
  AND2_X1 U6916 ( .A1(n7082), .A2(n5147), .ZN(n7048) );
  MUX2_X1 U6917 ( .A(n8918), .B(n5126), .S(n4271), .Z(n5148) );
  NAND2_X1 U6918 ( .A1(n5148), .A2(n5454), .ZN(n5151) );
  INV_X1 U6919 ( .A(n5148), .ZN(n5149) );
  INV_X1 U6920 ( .A(n5454), .ZN(n7086) );
  NAND2_X1 U6921 ( .A1(n5149), .A2(n7086), .ZN(n5150) );
  NAND2_X1 U6922 ( .A1(n5151), .A2(n5150), .ZN(n7081) );
  AOI21_X1 U6923 ( .B1(n7083), .B2(n7082), .A(n7081), .ZN(n7208) );
  INV_X1 U6924 ( .A(n5151), .ZN(n7207) );
  INV_X1 U6925 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n8896) );
  INV_X1 U6926 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n8994) );
  MUX2_X1 U6927 ( .A(n8896), .B(n8994), .S(n4271), .Z(n5152) );
  NAND2_X1 U6928 ( .A1(n5152), .A2(n5460), .ZN(n7274) );
  INV_X1 U6929 ( .A(n5152), .ZN(n5153) );
  NAND2_X1 U6930 ( .A1(n5153), .A2(n4796), .ZN(n5154) );
  AND2_X1 U6931 ( .A1(n7274), .A2(n5154), .ZN(n7206) );
  MUX2_X1 U6932 ( .A(n8873), .B(n9024), .S(n4271), .Z(n5155) );
  NAND2_X1 U6933 ( .A1(n5155), .A2(n5474), .ZN(n5158) );
  INV_X1 U6934 ( .A(n5155), .ZN(n5156) );
  INV_X1 U6935 ( .A(n5474), .ZN(n7272) );
  NAND2_X1 U6936 ( .A1(n5156), .A2(n7272), .ZN(n5157) );
  NAND2_X1 U6937 ( .A1(n5158), .A2(n5157), .ZN(n7273) );
  INV_X1 U6938 ( .A(n5158), .ZN(n7479) );
  INV_X1 U6939 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n9110) );
  MUX2_X1 U6940 ( .A(n9110), .B(n7602), .S(n4270), .Z(n5159) );
  NAND2_X1 U6941 ( .A1(n5159), .A2(n5495), .ZN(n7523) );
  INV_X1 U6942 ( .A(n5159), .ZN(n5160) );
  NAND2_X1 U6943 ( .A1(n5160), .A2(n7477), .ZN(n5161) );
  AND2_X1 U6944 ( .A1(n7523), .A2(n5161), .ZN(n7478) );
  INV_X1 U6945 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n8851) );
  INV_X1 U6946 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n8983) );
  MUX2_X1 U6947 ( .A(n8851), .B(n8983), .S(n4271), .Z(n5162) );
  NAND2_X1 U6948 ( .A1(n5162), .A2(n5501), .ZN(n5165) );
  INV_X1 U6949 ( .A(n5162), .ZN(n5163) );
  NAND2_X1 U6950 ( .A1(n5163), .A2(n7521), .ZN(n5164) );
  NAND2_X1 U6951 ( .A1(n5165), .A2(n5164), .ZN(n7522) );
  AOI21_X1 U6952 ( .B1(n7524), .B2(n7523), .A(n7522), .ZN(n8547) );
  INV_X1 U6953 ( .A(n5165), .ZN(n8546) );
  MUX2_X1 U6954 ( .A(n8837), .B(n9021), .S(n4270), .Z(n5166) );
  NAND2_X1 U6955 ( .A1(n5166), .A2(n5516), .ZN(n8559) );
  INV_X1 U6956 ( .A(n5166), .ZN(n5167) );
  NAND2_X1 U6957 ( .A1(n5167), .A2(n8544), .ZN(n5168) );
  AND2_X1 U6958 ( .A1(n8559), .A2(n5168), .ZN(n8545) );
  INV_X1 U6959 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n8976) );
  MUX2_X1 U6960 ( .A(n8825), .B(n8976), .S(n4270), .Z(n5169) );
  NAND2_X1 U6961 ( .A1(n5169), .A2(n5532), .ZN(n5172) );
  INV_X1 U6962 ( .A(n5169), .ZN(n5170) );
  NAND2_X1 U6963 ( .A1(n5170), .A2(n8557), .ZN(n5171) );
  NAND2_X1 U6964 ( .A1(n5172), .A2(n5171), .ZN(n8558) );
  INV_X1 U6965 ( .A(n5172), .ZN(n8578) );
  INV_X1 U6966 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n8813) );
  MUX2_X1 U6967 ( .A(n8813), .B(n8973), .S(n4271), .Z(n5173) );
  NAND2_X1 U6968 ( .A1(n5173), .A2(n5553), .ZN(n8591) );
  INV_X1 U6969 ( .A(n5553), .ZN(n8576) );
  INV_X1 U6970 ( .A(n5173), .ZN(n5174) );
  NAND2_X1 U6971 ( .A1(n8576), .A2(n5174), .ZN(n5175) );
  AND2_X1 U6972 ( .A1(n8591), .A2(n5175), .ZN(n8577) );
  INV_X1 U6973 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8970) );
  MUX2_X1 U6974 ( .A(n8804), .B(n8970), .S(n4270), .Z(n5176) );
  NAND2_X1 U6975 ( .A1(n5176), .A2(n5560), .ZN(n5179) );
  INV_X1 U6976 ( .A(n5176), .ZN(n5177) );
  NAND2_X1 U6977 ( .A1(n5177), .A2(n8589), .ZN(n5178) );
  NAND2_X1 U6978 ( .A1(n5179), .A2(n5178), .ZN(n8590) );
  AOI21_X1 U6979 ( .B1(n8592), .B2(n8591), .A(n8590), .ZN(n8608) );
  INV_X1 U6980 ( .A(n5179), .ZN(n8607) );
  XNOR2_X1 U6981 ( .A(n5180), .B(n5572), .ZN(n8606) );
  INV_X1 U6982 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8965) );
  MUX2_X1 U6983 ( .A(n5181), .B(n8965), .S(n4271), .Z(n5183) );
  INV_X1 U6984 ( .A(n5183), .ZN(n5184) );
  NAND2_X1 U6985 ( .A1(n5185), .A2(n5184), .ZN(n8627) );
  NAND2_X1 U6986 ( .A1(n8628), .A2(n8624), .ZN(n5188) );
  INV_X1 U6987 ( .A(n4271), .ZN(n5792) );
  MUX2_X1 U6988 ( .A(n4366), .B(n5186), .S(n5792), .Z(n5187) );
  XNOR2_X1 U6989 ( .A(n5188), .B(n5187), .ZN(n5197) );
  NAND2_X1 U6990 ( .A1(P2_U3893), .A2(n5190), .ZN(n8626) );
  INV_X1 U6991 ( .A(n5189), .ZN(n5194) );
  INV_X1 U6992 ( .A(n5190), .ZN(n8522) );
  OR2_X1 U6993 ( .A1(n4271), .A2(P2_U3151), .ZN(n5191) );
  NOR3_X1 U6994 ( .A1(n5192), .A2(n8522), .A3(n5191), .ZN(n5193) );
  AOI21_X2 U6995 ( .B1(n4364), .B2(n5194), .A(n5193), .ZN(n8615) );
  NAND2_X1 U6996 ( .A1(P2_U3151), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8127) );
  OAI21_X1 U6997 ( .B1(n8615), .B2(n4274), .A(n8127), .ZN(n5195) );
  AOI21_X1 U6998 ( .B1(P2_ADDR_REG_19__SCAN_IN), .B2(n8611), .A(n5195), .ZN(
        n5196) );
  INV_X1 U6999 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n5204) );
  INV_X1 U7000 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n5206) );
  INV_X1 U7001 ( .A(n5614), .ZN(n5615) );
  NAND2_X1 U7002 ( .A1(n4281), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n5207) );
  NAND2_X1 U7003 ( .A1(n5615), .A2(n5207), .ZN(n8773) );
  INV_X1 U7004 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5209) );
  NAND2_X1 U7005 ( .A1(n5212), .A2(n5209), .ZN(n5215) );
  XNOR2_X2 U7006 ( .A(n5211), .B(n5210), .ZN(n9273) );
  INV_X1 U7007 ( .A(n9277), .ZN(n5217) );
  AND2_X2 U7008 ( .A1(n5218), .A2(n5217), .ZN(n5370) );
  BUF_X4 U7009 ( .A(n5370), .Z(n6644) );
  NAND2_X1 U7010 ( .A1(n8773), .A2(n6644), .ZN(n5223) );
  AND2_X2 U7011 ( .A1(n5217), .A2(n9273), .ZN(n5349) );
  AND2_X2 U7012 ( .A1(n5218), .A2(n9277), .ZN(n5371) );
  INV_X4 U7013 ( .A(n5379), .ZN(n8457) );
  NAND2_X1 U7014 ( .A1(n8457), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n5220) );
  AND2_X2 U7015 ( .A1(n9273), .A2(n9277), .ZN(n5369) );
  NAND2_X1 U7016 ( .A1(n5369), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n5219) );
  OAI211_X1 U7017 ( .C1(n5368), .C2(n8960), .A(n5220), .B(n5219), .ZN(n5221)
         );
  INV_X1 U7018 ( .A(n5221), .ZN(n5222) );
  NAND2_X1 U7019 ( .A1(n5224), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n5225) );
  INV_X1 U7020 ( .A(SI_2_), .ZN(n5227) );
  NAND2_X1 U7021 ( .A1(n5231), .A2(n5227), .ZN(n5339) );
  INV_X1 U7022 ( .A(n5339), .ZN(n5230) );
  INV_X1 U7023 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n5228) );
  OAI22_X2 U7024 ( .A1(n5252), .A2(n5229), .B1(n5228), .B2(n5307), .ZN(n5235)
         );
  NOR2_X1 U7025 ( .A1(n5230), .A2(n5335), .ZN(n5234) );
  INV_X1 U7026 ( .A(n5231), .ZN(n5232) );
  NAND2_X1 U7027 ( .A1(n5232), .A2(SI_2_), .ZN(n5338) );
  INV_X1 U7028 ( .A(n5338), .ZN(n5233) );
  INV_X1 U7029 ( .A(n5235), .ZN(n5237) );
  INV_X1 U7030 ( .A(SI_1_), .ZN(n5236) );
  NAND2_X1 U7031 ( .A1(n5237), .A2(n5236), .ZN(n5336) );
  INV_X4 U7032 ( .A(n5307), .ZN(n5609) );
  INV_X1 U7033 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5366) );
  INV_X1 U7034 ( .A(SI_0_), .ZN(n5928) );
  INV_X1 U7035 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5929) );
  NAND2_X1 U7036 ( .A1(n5252), .A2(n5929), .ZN(n5238) );
  INV_X1 U7037 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6790) );
  INV_X1 U7038 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n5241) );
  INV_X1 U7039 ( .A(SI_4_), .ZN(n5243) );
  NAND2_X1 U7040 ( .A1(n5609), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n5244) );
  INV_X1 U7041 ( .A(n5257), .ZN(n5247) );
  INV_X1 U7042 ( .A(SI_3_), .ZN(n5246) );
  NAND2_X1 U7043 ( .A1(n5247), .A2(n5246), .ZN(n5384) );
  NAND2_X1 U7044 ( .A1(n5395), .A2(n5384), .ZN(n5324) );
  INV_X1 U7045 ( .A(n5263), .ZN(n5251) );
  INV_X1 U7046 ( .A(SI_5_), .ZN(n5250) );
  INV_X1 U7047 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6806) );
  INV_X1 U7048 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n5253) );
  MUX2_X1 U7049 ( .A(n6806), .B(n5253), .S(n5252), .Z(n5265) );
  INV_X1 U7050 ( .A(SI_6_), .ZN(n5254) );
  NAND2_X2 U7051 ( .A1(n5265), .A2(n5254), .ZN(n5414) );
  NAND2_X1 U7052 ( .A1(n5327), .A2(n5414), .ZN(n5256) );
  INV_X1 U7053 ( .A(n5256), .ZN(n5262) );
  INV_X1 U7054 ( .A(n5392), .ZN(n5258) );
  INV_X1 U7055 ( .A(n5259), .ZN(n5260) );
  NAND2_X1 U7056 ( .A1(n5260), .A2(SI_4_), .ZN(n5394) );
  NAND2_X1 U7057 ( .A1(n5261), .A2(n5394), .ZN(n5325) );
  NAND2_X1 U7058 ( .A1(n5263), .A2(SI_5_), .ZN(n5411) );
  INV_X1 U7059 ( .A(n5411), .ZN(n5264) );
  NAND2_X1 U7060 ( .A1(n5264), .A2(n5414), .ZN(n5267) );
  INV_X1 U7061 ( .A(n5265), .ZN(n5266) );
  NAND2_X1 U7062 ( .A1(n5266), .A2(SI_6_), .ZN(n5413) );
  INV_X8 U7063 ( .A(n5307), .ZN(n6779) );
  NAND2_X1 U7064 ( .A1(n5269), .A2(SI_7_), .ZN(n5271) );
  OAI21_X1 U7065 ( .B1(n5269), .B2(SI_7_), .A(n5271), .ZN(n5436) );
  INV_X1 U7066 ( .A(n5436), .ZN(n5270) );
  MUX2_X1 U7067 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .S(n6779), .Z(n5272) );
  OAI22_X2 U7068 ( .A1(n5453), .A2(n5452), .B1(SI_8_), .B2(n5272), .ZN(n5459)
         );
  MUX2_X1 U7069 ( .A(n9108), .B(n5273), .S(n6779), .Z(n5275) );
  INV_X1 U7070 ( .A(SI_9_), .ZN(n5274) );
  NAND2_X1 U7071 ( .A1(n5275), .A2(n5274), .ZN(n5276) );
  MUX2_X1 U7072 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .S(n6779), .Z(n5277) );
  MUX2_X1 U7073 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .S(n6779), .Z(n5280) );
  MUX2_X1 U7074 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .S(n6779), .Z(n5281) );
  MUX2_X1 U7075 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n6779), .Z(n5282) );
  NAND2_X1 U7076 ( .A1(n5282), .A2(SI_13_), .ZN(n5514) );
  INV_X1 U7077 ( .A(n5282), .ZN(n5284) );
  INV_X1 U7078 ( .A(SI_13_), .ZN(n5283) );
  MUX2_X1 U7079 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n6779), .Z(n5529) );
  MUX2_X1 U7080 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .S(n6779), .Z(n5551) );
  INV_X1 U7081 ( .A(SI_15_), .ZN(n5287) );
  MUX2_X1 U7082 ( .A(n7158), .B(n9072), .S(n6779), .Z(n5558) );
  INV_X1 U7083 ( .A(SI_16_), .ZN(n5286) );
  AOI22_X1 U7084 ( .A1(n5556), .A2(n5287), .B1(n5558), .B2(n5286), .ZN(n5285)
         );
  OAI21_X1 U7085 ( .B1(n5556), .B2(n5287), .A(n5286), .ZN(n5290) );
  INV_X1 U7086 ( .A(n5558), .ZN(n5289) );
  AND2_X1 U7087 ( .A1(SI_16_), .A2(SI_15_), .ZN(n5288) );
  AOI22_X1 U7088 ( .A1(n5290), .A2(n5289), .B1(n5551), .B2(n5288), .ZN(n5291)
         );
  INV_X1 U7089 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n5292) );
  MUX2_X1 U7090 ( .A(n7145), .B(n5292), .S(n6779), .Z(n5294) );
  INV_X1 U7091 ( .A(SI_17_), .ZN(n5293) );
  INV_X1 U7092 ( .A(n5294), .ZN(n5295) );
  NAND2_X1 U7093 ( .A1(n5295), .A2(SI_17_), .ZN(n5296) );
  MUX2_X1 U7094 ( .A(n9118), .B(n9104), .S(n6779), .Z(n5299) );
  INV_X1 U7095 ( .A(n5299), .ZN(n5300) );
  MUX2_X1 U7096 ( .A(n8096), .B(n7289), .S(n6779), .Z(n5304) );
  INV_X1 U7097 ( .A(SI_19_), .ZN(n5303) );
  INV_X1 U7098 ( .A(n5304), .ZN(n5305) );
  NAND2_X1 U7099 ( .A1(n5305), .A2(SI_19_), .ZN(n5306) );
  AOI22_X1 U7100 ( .A1(n5587), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n6701), .B2(
        n6710), .ZN(n5308) );
  NAND2_X1 U7101 ( .A1(n5309), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5311) );
  NAND2_X1 U7102 ( .A1(n5312), .A2(n8503), .ZN(n6618) );
  XNOR2_X1 U7103 ( .A(n5313), .B(P2_B_REG_SCAN_IN), .ZN(n5314) );
  NAND2_X1 U7104 ( .A1(n5314), .A2(n7712), .ZN(n5315) );
  INV_X1 U7105 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n6803) );
  NAND2_X1 U7106 ( .A1(n7731), .A2(n5313), .ZN(n6800) );
  INV_X1 U7107 ( .A(n8295), .ZN(n7518) );
  NAND2_X1 U7108 ( .A1(n7518), .A2(n6702), .ZN(n8510) );
  INV_X1 U7109 ( .A(n8510), .ZN(n5317) );
  NAND2_X1 U7110 ( .A1(n5772), .A2(n5317), .ZN(n5318) );
  NAND2_X1 U7111 ( .A1(n8295), .A2(n8503), .ZN(n8463) );
  NAND3_X1 U7112 ( .A1(n6618), .A2(n5318), .A3(n8463), .ZN(n5363) );
  XNOR2_X1 U7113 ( .A(n9213), .B(n8132), .ZN(n5605) );
  NAND2_X1 U7114 ( .A1(n5349), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n5323) );
  NAND2_X1 U7115 ( .A1(n5401), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5319) );
  NAND2_X1 U7116 ( .A1(n5419), .A2(n5319), .ZN(n7256) );
  NAND2_X1 U7117 ( .A1(n6644), .A2(n7256), .ZN(n5322) );
  NAND2_X1 U7118 ( .A1(n8457), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n5321) );
  NAND2_X1 U7119 ( .A1(n5369), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5320) );
  NAND4_X1 U7120 ( .A1(n5323), .A2(n5322), .A3(n5321), .A4(n5320), .ZN(n8535)
         );
  INV_X1 U7121 ( .A(n8535), .ZN(n7292) );
  INV_X1 U7122 ( .A(n5324), .ZN(n5326) );
  NAND2_X1 U7123 ( .A1(n5411), .A2(n5327), .ZN(n5329) );
  NAND2_X1 U7124 ( .A1(n5328), .A2(n5329), .ZN(n5332) );
  INV_X1 U7125 ( .A(n5328), .ZN(n5331) );
  INV_X1 U7126 ( .A(n5329), .ZN(n5330) );
  NAND2_X1 U7127 ( .A1(n5331), .A2(n5330), .ZN(n5412) );
  OR2_X1 U7128 ( .A1(n5358), .A2(n6786), .ZN(n5334) );
  OR2_X1 U7129 ( .A1(n8435), .A2(n5249), .ZN(n5333) );
  OAI211_X1 U7130 ( .C1(n5794), .C2(n6785), .A(n5334), .B(n5333), .ZN(n7257)
         );
  INV_X1 U7131 ( .A(n7257), .ZN(n7199) );
  XNOR2_X1 U7132 ( .A(n7199), .B(n8132), .ZN(n5409) );
  INV_X1 U7133 ( .A(n5409), .ZN(n5410) );
  NAND2_X1 U7134 ( .A1(n5336), .A2(n5335), .ZN(n5355) );
  INV_X1 U7135 ( .A(n5355), .ZN(n5337) );
  NAND2_X1 U7136 ( .A1(n5337), .A2(n5354), .ZN(n5357) );
  NAND2_X1 U7137 ( .A1(n5357), .A2(n5335), .ZN(n5341) );
  AND2_X1 U7138 ( .A1(n5339), .A2(n5338), .ZN(n5340) );
  XNOR2_X1 U7139 ( .A(n5341), .B(n5340), .ZN(n6789) );
  OR2_X1 U7140 ( .A1(n5358), .A2(n6789), .ZN(n5344) );
  OR2_X1 U7141 ( .A1(n8435), .A2(n4496), .ZN(n5343) );
  OR2_X1 U7142 ( .A1(n5794), .A2(n6851), .ZN(n5342) );
  NAND2_X1 U7143 ( .A1(n5349), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5348) );
  NAND2_X1 U7144 ( .A1(n5370), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n5347) );
  NAND2_X1 U7145 ( .A1(n5371), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n5346) );
  NAND2_X1 U7146 ( .A1(n5369), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5345) );
  NAND2_X1 U7147 ( .A1(n5349), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5353) );
  NAND2_X1 U7148 ( .A1(n5369), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n5352) );
  NAND2_X1 U7149 ( .A1(n5370), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n5351) );
  NAND2_X1 U7150 ( .A1(n5371), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n5350) );
  NAND2_X1 U7151 ( .A1(n5355), .A2(n5239), .ZN(n5356) );
  AND2_X1 U7152 ( .A1(n5357), .A2(n5356), .ZN(n6777) );
  OR2_X1 U7153 ( .A1(n5387), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n5362) );
  OR2_X1 U7154 ( .A1(n5360), .A2(n5359), .ZN(n5361) );
  XNOR2_X1 U7155 ( .A(n7103), .B(n5363), .ZN(n5364) );
  NOR2_X1 U7156 ( .A1(n4967), .A2(n5364), .ZN(n5376) );
  NOR2_X1 U7157 ( .A1(n5376), .A2(n5365), .ZN(n6876) );
  NAND2_X1 U7158 ( .A1(n6778), .A2(SI_0_), .ZN(n5367) );
  XNOR2_X1 U7159 ( .A(n5367), .B(n5366), .ZN(n9287) );
  NAND2_X1 U7160 ( .A1(n5349), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5375) );
  NAND2_X1 U7161 ( .A1(n5369), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5374) );
  NAND2_X1 U7162 ( .A1(n5370), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n5373) );
  NAND2_X1 U7163 ( .A1(n5371), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5372) );
  OAI21_X1 U7164 ( .B1(n7019), .B2(n5442), .A(n7099), .ZN(n6878) );
  INV_X1 U7165 ( .A(n5376), .ZN(n5377) );
  NAND2_X1 U7166 ( .A1(n6877), .A2(n5377), .ZN(n6959) );
  XNOR2_X1 U7167 ( .A(n5378), .B(n6880), .ZN(n6961) );
  NAND2_X1 U7168 ( .A1(n6959), .A2(n6961), .ZN(n6960) );
  OAI21_X1 U7169 ( .B1(n5378), .B2(n8538), .A(n6960), .ZN(n7137) );
  NAND2_X1 U7170 ( .A1(n8456), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5383) );
  NAND2_X1 U7171 ( .A1(n6644), .A2(n7142), .ZN(n5382) );
  NAND2_X1 U7172 ( .A1(n8457), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n5381) );
  NAND2_X1 U7173 ( .A1(n5369), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5380) );
  AND4_X2 U7174 ( .A1(n5383), .A2(n5382), .A3(n5381), .A4(n5380), .ZN(n6621)
         );
  NAND2_X1 U7175 ( .A1(n5386), .A2(n5393), .ZN(n6782) );
  OR2_X1 U7176 ( .A1(n5358), .A2(n6782), .ZN(n5389) );
  OR2_X1 U7178 ( .A1(n8452), .A2(n5245), .ZN(n5388) );
  OAI211_X1 U7179 ( .C1(n5794), .C2(n7068), .A(n5389), .B(n5388), .ZN(n7132)
         );
  XNOR2_X1 U7180 ( .A(n5442), .B(n7132), .ZN(n5390) );
  XNOR2_X1 U7181 ( .A(n6621), .B(n5390), .ZN(n7139) );
  INV_X1 U7182 ( .A(n5390), .ZN(n5391) );
  NAND2_X1 U7183 ( .A1(n5393), .A2(n5392), .ZN(n5397) );
  AND2_X1 U7184 ( .A1(n5395), .A2(n5394), .ZN(n5396) );
  XNOR2_X1 U7185 ( .A(n5397), .B(n5396), .ZN(n5986) );
  OR2_X1 U7186 ( .A1(n5986), .A2(n5358), .ZN(n5399) );
  OR2_X1 U7187 ( .A1(n8452), .A2(n6790), .ZN(n5398) );
  OAI211_X1 U7188 ( .C1(n5794), .C2(n7037), .A(n5399), .B(n5398), .ZN(n7219)
         );
  XNOR2_X1 U7189 ( .A(n5442), .B(n7219), .ZN(n5406) );
  INV_X1 U7190 ( .A(n5406), .ZN(n5407) );
  NAND2_X1 U7191 ( .A1(n5349), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5405) );
  NAND2_X1 U7192 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n5400) );
  NAND2_X1 U7193 ( .A1(n5401), .A2(n5400), .ZN(n7218) );
  NAND2_X1 U7194 ( .A1(n6644), .A2(n7218), .ZN(n5404) );
  NAND2_X1 U7195 ( .A1(n5369), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n5403) );
  NAND2_X1 U7196 ( .A1(n8457), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5402) );
  AND2_X1 U7197 ( .A1(n7136), .A2(n5406), .ZN(n5408) );
  AOI21_X1 U7198 ( .B1(n5407), .B2(n8536), .A(n5408), .ZN(n7161) );
  INV_X1 U7199 ( .A(n5408), .ZN(n7231) );
  XNOR2_X1 U7200 ( .A(n5409), .B(n8535), .ZN(n7232) );
  AOI21_X1 U7201 ( .B1(n7292), .B2(n5410), .A(n7230), .ZN(n7263) );
  AOI22_X1 U7202 ( .A1(n5587), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n6804), .B2(
        n6710), .ZN(n5418) );
  NAND2_X1 U7203 ( .A1(n5412), .A2(n5411), .ZN(n5416) );
  NAND2_X1 U7204 ( .A1(n5414), .A2(n5413), .ZN(n5415) );
  XNOR2_X2 U7205 ( .A(n5416), .B(n5415), .ZN(n6793) );
  NAND2_X1 U7206 ( .A1(n6793), .A2(n8450), .ZN(n5417) );
  NAND2_X1 U7207 ( .A1(n5418), .A2(n5417), .ZN(n7340) );
  XNOR2_X1 U7208 ( .A(n7340), .B(n8132), .ZN(n5425) );
  NAND2_X1 U7209 ( .A1(n4272), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5424) );
  NAND2_X1 U7210 ( .A1(n5419), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5420) );
  NAND2_X1 U7211 ( .A1(n5427), .A2(n5420), .ZN(n7339) );
  NAND2_X1 U7212 ( .A1(n6644), .A2(n7339), .ZN(n5423) );
  NAND2_X1 U7213 ( .A1(n8457), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n5422) );
  NAND2_X1 U7214 ( .A1(n8455), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5421) );
  NAND4_X1 U7215 ( .A1(n5424), .A2(n5423), .A3(n5422), .A4(n5421), .ZN(n8534)
         );
  XNOR2_X1 U7216 ( .A(n5425), .B(n8534), .ZN(n7262) );
  NAND2_X1 U7217 ( .A1(n7263), .A2(n7262), .ZN(n7261) );
  INV_X1 U7218 ( .A(n8534), .ZN(n7390) );
  NAND2_X1 U7219 ( .A1(n4272), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n5433) );
  NAND2_X1 U7220 ( .A1(n5427), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5428) );
  NAND2_X1 U7221 ( .A1(n5446), .A2(n5428), .ZN(n7550) );
  NAND2_X1 U7222 ( .A1(n6644), .A2(n7550), .ZN(n5432) );
  NAND2_X1 U7223 ( .A1(n8457), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n5431) );
  INV_X2 U7224 ( .A(n5429), .ZN(n8455) );
  NAND2_X1 U7225 ( .A1(n8455), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5430) );
  NAND2_X1 U7226 ( .A1(n5437), .A2(n5436), .ZN(n5439) );
  NAND2_X1 U7227 ( .A1(n5439), .A2(n5438), .ZN(n6792) );
  NOR2_X1 U7228 ( .A1(n6792), .A2(n5358), .ZN(n5441) );
  OAI22_X1 U7229 ( .A1(n8452), .A2(n4463), .B1(n6791), .B2(n5794), .ZN(n5440)
         );
  XNOR2_X1 U7230 ( .A(n5442), .B(n7445), .ZN(n5444) );
  XNOR2_X1 U7231 ( .A(n8906), .B(n5444), .ZN(n7450) );
  INV_X1 U7232 ( .A(n7450), .ZN(n5443) );
  NAND2_X1 U7233 ( .A1(n8906), .A2(n5444), .ZN(n5445) );
  NAND2_X1 U7234 ( .A1(n4272), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5451) );
  NAND2_X1 U7235 ( .A1(n5446), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5447) );
  NAND2_X1 U7236 ( .A1(n5463), .A2(n5447), .ZN(n8919) );
  NAND2_X1 U7237 ( .A1(n6644), .A2(n8919), .ZN(n5450) );
  NAND2_X1 U7238 ( .A1(n8457), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n5449) );
  NAND2_X1 U7239 ( .A1(n8455), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n5448) );
  XNOR2_X1 U7240 ( .A(n5453), .B(n5452), .ZN(n6807) );
  NAND2_X1 U7241 ( .A1(n6807), .A2(n8450), .ZN(n5456) );
  AOI22_X1 U7242 ( .A1(n5587), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n5454), .B2(
        n6710), .ZN(n5455) );
  NAND2_X1 U7243 ( .A1(n5456), .A2(n5455), .ZN(n8997) );
  XNOR2_X1 U7244 ( .A(n8997), .B(n8132), .ZN(n8110) );
  NAND2_X1 U7245 ( .A1(n6815), .A2(n8450), .ZN(n5462) );
  AOI22_X1 U7246 ( .A1(n5587), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n5460), .B2(
        n6710), .ZN(n5461) );
  NAND2_X1 U7247 ( .A1(n5462), .A2(n5461), .ZN(n8898) );
  XNOR2_X1 U7248 ( .A(n8898), .B(n8132), .ZN(n8111) );
  INV_X1 U7249 ( .A(n8111), .ZN(n5469) );
  NAND2_X1 U7250 ( .A1(n4272), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n5468) );
  NAND2_X1 U7251 ( .A1(n5463), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n5464) );
  NAND2_X1 U7252 ( .A1(n5477), .A2(n5464), .ZN(n8897) );
  NAND2_X1 U7253 ( .A1(n6644), .A2(n8897), .ZN(n5467) );
  NAND2_X1 U7254 ( .A1(n8457), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n5466) );
  NAND2_X1 U7255 ( .A1(n8455), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5465) );
  NAND2_X1 U7256 ( .A1(n5469), .A2(n8916), .ZN(n8112) );
  OAI21_X1 U7257 ( .B1(n8222), .B2(n8110), .A(n8112), .ZN(n5484) );
  NAND2_X1 U7258 ( .A1(n5471), .A2(n5470), .ZN(n5472) );
  NAND2_X1 U7259 ( .A1(n5473), .A2(n5472), .ZN(n6825) );
  OR2_X1 U7260 ( .A1(n6825), .A2(n5358), .ZN(n5476) );
  AOI22_X1 U7261 ( .A1(n5587), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n5474), .B2(
        n6710), .ZN(n5475) );
  NAND2_X2 U7262 ( .A1(n5476), .A2(n5475), .ZN(n8875) );
  XNOR2_X1 U7263 ( .A(n8875), .B(n8132), .ZN(n8113) );
  NAND2_X1 U7264 ( .A1(n4272), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n5482) );
  NAND2_X1 U7265 ( .A1(n5477), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5478) );
  NAND2_X1 U7266 ( .A1(n5487), .A2(n5478), .ZN(n8874) );
  NAND2_X1 U7267 ( .A1(n6644), .A2(n8874), .ZN(n5481) );
  NAND2_X1 U7268 ( .A1(n8457), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n5480) );
  NAND2_X1 U7269 ( .A1(n8455), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5479) );
  NAND4_X1 U7270 ( .A1(n5482), .A2(n5481), .A3(n5480), .A4(n5479), .ZN(n8889)
         );
  INV_X1 U7271 ( .A(n8916), .ZN(n6625) );
  AOI22_X1 U7272 ( .A1(n8113), .A2(n8345), .B1(n6625), .B2(n8111), .ZN(n5483)
         );
  NAND2_X1 U7273 ( .A1(n4272), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n5492) );
  NAND2_X1 U7274 ( .A1(n8457), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n5491) );
  NAND2_X1 U7275 ( .A1(n5487), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5488) );
  NAND2_X1 U7276 ( .A1(n5504), .A2(n5488), .ZN(n7634) );
  NAND2_X1 U7277 ( .A1(n6644), .A2(n7634), .ZN(n5490) );
  NAND2_X1 U7278 ( .A1(n8455), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5489) );
  XNOR2_X1 U7279 ( .A(n5494), .B(n5493), .ZN(n6835) );
  NAND2_X1 U7280 ( .A1(n6835), .A2(n8450), .ZN(n5497) );
  AOI22_X1 U7281 ( .A1(n5587), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n5495), .B2(
        n6710), .ZN(n5496) );
  NOR2_X1 U7282 ( .A1(n8340), .A2(n8846), .ZN(n6662) );
  AOI21_X2 U7283 ( .B1(n8846), .B2(n8340), .A(n6662), .ZN(n8493) );
  XNOR2_X1 U7284 ( .A(n8493), .B(n5457), .ZN(n8163) );
  NAND2_X1 U7285 ( .A1(n5499), .A2(n5498), .ZN(n5500) );
  OR2_X1 U7286 ( .A1(n6842), .A2(n5358), .ZN(n5503) );
  AOI22_X1 U7287 ( .A1(n5587), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n5501), .B2(
        n6710), .ZN(n5502) );
  XNOR2_X1 U7288 ( .A(n8169), .B(n5457), .ZN(n5510) );
  NAND2_X1 U7289 ( .A1(n8457), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n5509) );
  NAND2_X1 U7290 ( .A1(n4272), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n5508) );
  NAND2_X1 U7291 ( .A1(n5504), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5505) );
  NAND2_X1 U7292 ( .A1(n5519), .A2(n5505), .ZN(n8849) );
  NAND2_X1 U7293 ( .A1(n6644), .A2(n8849), .ZN(n5507) );
  NAND2_X1 U7294 ( .A1(n8455), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5506) );
  NAND2_X1 U7295 ( .A1(n5510), .A2(n8355), .ZN(n8236) );
  INV_X1 U7296 ( .A(n8236), .ZN(n8165) );
  NOR2_X1 U7297 ( .A1(n8165), .A2(n8846), .ZN(n5526) );
  INV_X1 U7298 ( .A(n8163), .ZN(n5525) );
  NOR2_X1 U7299 ( .A1(n5510), .A2(n8355), .ZN(n8235) );
  NAND2_X1 U7300 ( .A1(n6180), .A2(n8450), .ZN(n5518) );
  AOI22_X1 U7301 ( .A1(n5587), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n5516), .B2(
        n6710), .ZN(n5517) );
  XNOR2_X1 U7302 ( .A(n9248), .B(n8132), .ZN(n5528) );
  NAND2_X1 U7303 ( .A1(n4272), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n5524) );
  NAND2_X1 U7304 ( .A1(n5519), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n5520) );
  NAND2_X1 U7305 ( .A1(n5535), .A2(n5520), .ZN(n8832) );
  NAND2_X1 U7306 ( .A1(n6644), .A2(n8832), .ZN(n5523) );
  NAND2_X1 U7307 ( .A1(n8455), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5522) );
  NAND2_X1 U7308 ( .A1(n8457), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n5521) );
  NAND4_X1 U7309 ( .A1(n5524), .A2(n5523), .A3(n5522), .A4(n5521), .ZN(n8819)
         );
  INV_X1 U7310 ( .A(n8819), .ZN(n8847) );
  XNOR2_X1 U7311 ( .A(n5528), .B(n8847), .ZN(n8238) );
  XNOR2_X1 U7312 ( .A(n5529), .B(SI_14_), .ZN(n5530) );
  XNOR2_X1 U7313 ( .A(n5531), .B(n5530), .ZN(n6957) );
  NAND2_X1 U7314 ( .A1(n6957), .A2(n8450), .ZN(n5534) );
  AOI22_X1 U7315 ( .A1(n5587), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n5532), .B2(
        n6710), .ZN(n5533) );
  XNOR2_X1 U7316 ( .A(n8361), .B(n5442), .ZN(n5541) );
  NAND2_X1 U7317 ( .A1(n4272), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n5540) );
  NAND2_X1 U7318 ( .A1(n5535), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5536) );
  NAND2_X1 U7319 ( .A1(n5545), .A2(n5536), .ZN(n8821) );
  NAND2_X1 U7320 ( .A1(n6644), .A2(n8821), .ZN(n5539) );
  NAND2_X1 U7321 ( .A1(n8457), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n5538) );
  NAND2_X1 U7322 ( .A1(n8455), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5537) );
  XNOR2_X1 U7323 ( .A(n5541), .B(n6667), .ZN(n8098) );
  INV_X1 U7324 ( .A(n5541), .ZN(n5542) );
  NAND2_X1 U7325 ( .A1(n5542), .A2(n6667), .ZN(n5543) );
  NAND2_X1 U7326 ( .A1(n5544), .A2(n5543), .ZN(n8182) );
  NAND2_X1 U7327 ( .A1(n4272), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n5550) );
  NAND2_X1 U7328 ( .A1(n5545), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5546) );
  NAND2_X1 U7329 ( .A1(n5565), .A2(n5546), .ZN(n8814) );
  NAND2_X1 U7330 ( .A1(n6644), .A2(n8814), .ZN(n5549) );
  NAND2_X1 U7331 ( .A1(n8457), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n5548) );
  NAND2_X1 U7332 ( .A1(n8455), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n5547) );
  NAND4_X1 U7333 ( .A1(n5550), .A2(n5549), .A3(n5548), .A4(n5547), .ZN(n8818)
         );
  XNOR2_X1 U7334 ( .A(n5551), .B(SI_15_), .ZN(n5552) );
  XNOR2_X1 U7335 ( .A(n5557), .B(n5552), .ZN(n7106) );
  NAND2_X1 U7336 ( .A1(n7106), .A2(n8450), .ZN(n5555) );
  AOI22_X1 U7337 ( .A1(n5587), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n5553), .B2(
        n6710), .ZN(n5554) );
  XNOR2_X1 U7338 ( .A(n9235), .B(n8132), .ZN(n5595) );
  XOR2_X1 U7339 ( .A(n8818), .B(n5595), .Z(n8280) );
  XNOR2_X1 U7340 ( .A(n5558), .B(SI_16_), .ZN(n5559) );
  NAND2_X1 U7341 ( .A1(n7157), .A2(n8450), .ZN(n5562) );
  AOI22_X1 U7342 ( .A1(n5587), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n5560), .B2(
        n6710), .ZN(n5561) );
  XNOR2_X1 U7343 ( .A(n9229), .B(n5457), .ZN(n8184) );
  NAND2_X1 U7344 ( .A1(n4272), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n5564) );
  NAND2_X1 U7345 ( .A1(n8457), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n5563) );
  AND2_X1 U7346 ( .A1(n5564), .A2(n5563), .ZN(n5569) );
  NAND2_X1 U7347 ( .A1(n5565), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5566) );
  NAND2_X1 U7348 ( .A1(n5575), .A2(n5566), .ZN(n8805) );
  NAND2_X1 U7349 ( .A1(n8805), .A2(n6644), .ZN(n5568) );
  NAND2_X1 U7350 ( .A1(n8455), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n5567) );
  NAND2_X1 U7351 ( .A1(n8184), .A2(n8811), .ZN(n8196) );
  XNOR2_X1 U7352 ( .A(n5571), .B(n5570), .ZN(n7122) );
  NAND2_X1 U7353 ( .A1(n7122), .A2(n8450), .ZN(n5574) );
  AOI22_X1 U7354 ( .A1(n5587), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n5572), .B2(
        n6710), .ZN(n5573) );
  XNOR2_X1 U7355 ( .A(n9223), .B(n8132), .ZN(n5581) );
  INV_X1 U7356 ( .A(n5581), .ZN(n5580) );
  NAND2_X1 U7357 ( .A1(n5575), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n5576) );
  NAND2_X1 U7358 ( .A1(n5590), .A2(n5576), .ZN(n8796) );
  NAND2_X1 U7359 ( .A1(n8796), .A2(n6644), .ZN(n5579) );
  AOI22_X1 U7360 ( .A1(P2_REG1_REG_17__SCAN_IN), .A2(n4272), .B1(n8457), .B2(
        P2_REG2_REG_17__SCAN_IN), .ZN(n5578) );
  NAND2_X1 U7361 ( .A1(n5369), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n5577) );
  INV_X1 U7362 ( .A(n8778), .ZN(n8802) );
  NAND2_X1 U7363 ( .A1(n5580), .A2(n8802), .ZN(n8193) );
  AND2_X1 U7364 ( .A1(n8196), .A2(n8193), .ZN(n5597) );
  OR2_X1 U7365 ( .A1(n8184), .A2(n8811), .ZN(n8195) );
  OR2_X1 U7366 ( .A1(n8280), .A2(n5598), .ZN(n5582) );
  NAND2_X1 U7367 ( .A1(n5581), .A2(n8778), .ZN(n8192) );
  INV_X1 U7368 ( .A(n8192), .ZN(n5599) );
  OR2_X1 U7369 ( .A1(n5582), .A2(n5599), .ZN(n5583) );
  NOR2_X1 U7370 ( .A1(n8182), .A2(n5583), .ZN(n8260) );
  XNOR2_X1 U7371 ( .A(n5585), .B(n5584), .ZN(n7191) );
  NAND2_X1 U7372 ( .A1(n7191), .A2(n8450), .ZN(n5589) );
  AOI22_X1 U7373 ( .A1(n5587), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n5586), .B2(
        n6710), .ZN(n5588) );
  XNOR2_X1 U7374 ( .A(n9220), .B(n5442), .ZN(n5601) );
  NAND2_X1 U7375 ( .A1(n5590), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5591) );
  NAND2_X1 U7376 ( .A1(n4281), .A2(n5591), .ZN(n8782) );
  NAND2_X1 U7377 ( .A1(n8782), .A2(n6644), .ZN(n5594) );
  AOI22_X1 U7378 ( .A1(P2_REG1_REG_18__SCAN_IN), .A2(n4272), .B1(n8457), .B2(
        P2_REG2_REG_18__SCAN_IN), .ZN(n5593) );
  NAND2_X1 U7379 ( .A1(n8455), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n5592) );
  XNOR2_X1 U7380 ( .A(n5601), .B(n8793), .ZN(n8263) );
  INV_X1 U7381 ( .A(n8263), .ZN(n5600) );
  INV_X1 U7382 ( .A(n5595), .ZN(n5596) );
  NAND2_X1 U7383 ( .A1(n5596), .A2(n8818), .ZN(n8183) );
  NAND2_X1 U7384 ( .A1(n5600), .A2(n8261), .ZN(n5604) );
  INV_X1 U7385 ( .A(n5601), .ZN(n5602) );
  NAND2_X1 U7386 ( .A1(n5602), .A2(n8768), .ZN(n5603) );
  XNOR2_X1 U7387 ( .A(n5605), .B(n8779), .ZN(n8122) );
  INV_X1 U7388 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7335) );
  INV_X1 U7389 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7401) );
  MUX2_X1 U7390 ( .A(n7335), .B(n7401), .S(n6779), .Z(n5640) );
  XNOR2_X1 U7391 ( .A(n5640), .B(SI_20_), .ZN(n5610) );
  XNOR2_X1 U7392 ( .A(n5647), .B(n5610), .ZN(n7334) );
  NAND2_X1 U7393 ( .A1(n7334), .A2(n8450), .ZN(n5612) );
  OR2_X1 U7394 ( .A1(n8435), .A2(n7335), .ZN(n5611) );
  XNOR2_X1 U7395 ( .A(n9207), .B(n8132), .ZN(n5622) );
  INV_X1 U7396 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n5613) );
  NAND2_X1 U7397 ( .A1(n5615), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n5616) );
  NAND2_X1 U7398 ( .A1(n4285), .A2(n5616), .ZN(n8761) );
  NAND2_X1 U7399 ( .A1(n8761), .A2(n6644), .ZN(n5621) );
  INV_X1 U7400 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n9206) );
  NAND2_X1 U7401 ( .A1(n4272), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n5618) );
  NAND2_X1 U7402 ( .A1(n8457), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n5617) );
  OAI211_X1 U7403 ( .C1(n9206), .C2(n5429), .A(n5618), .B(n5617), .ZN(n5619)
         );
  INV_X1 U7404 ( .A(n5619), .ZN(n5620) );
  XNOR2_X1 U7405 ( .A(n5622), .B(n8769), .ZN(n8229) );
  NAND2_X1 U7406 ( .A1(n5622), .A2(n8769), .ZN(n5623) );
  NAND2_X1 U7407 ( .A1(n8226), .A2(n5623), .ZN(n8156) );
  INV_X1 U7408 ( .A(SI_20_), .ZN(n5639) );
  NAND2_X1 U7409 ( .A1(n5647), .A2(n5639), .ZN(n5624) );
  INV_X1 U7410 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7540) );
  MUX2_X1 U7411 ( .A(n9007), .B(n7540), .S(n6779), .Z(n5637) );
  XNOR2_X1 U7412 ( .A(n5637), .B(SI_21_), .ZN(n5626) );
  NAND2_X1 U7413 ( .A1(n7517), .A2(n8450), .ZN(n5629) );
  OR2_X1 U7414 ( .A1(n8452), .A2(n9007), .ZN(n5628) );
  NAND2_X2 U7415 ( .A1(n5629), .A2(n5628), .ZN(n8954) );
  INV_X1 U7416 ( .A(n8954), .ZN(n6678) );
  XNOR2_X1 U7417 ( .A(n6678), .B(n5442), .ZN(n5661) );
  INV_X1 U7418 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n5630) );
  NAND2_X1 U7419 ( .A1(n4285), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n5631) );
  NAND2_X1 U7420 ( .A1(n5654), .A2(n5631), .ZN(n8748) );
  NAND2_X1 U7421 ( .A1(n8748), .A2(n6644), .ZN(n5636) );
  INV_X1 U7422 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n9062) );
  NAND2_X1 U7423 ( .A1(n4272), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n5633) );
  NAND2_X1 U7424 ( .A1(n8455), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n5632) );
  OAI211_X1 U7425 ( .C1(n5379), .C2(n9062), .A(n5633), .B(n5632), .ZN(n5634)
         );
  INV_X1 U7426 ( .A(n5634), .ZN(n5635) );
  XNOR2_X1 U7427 ( .A(n5661), .B(n8253), .ZN(n8157) );
  NAND2_X1 U7428 ( .A1(n8156), .A2(n8157), .ZN(n8247) );
  INV_X1 U7429 ( .A(n5640), .ZN(n5642) );
  OAI22_X1 U7430 ( .A1(n5642), .A2(SI_20_), .B1(n5643), .B2(SI_21_), .ZN(n5646) );
  INV_X1 U7431 ( .A(SI_21_), .ZN(n5638) );
  OAI21_X1 U7432 ( .B1(n5640), .B2(n5639), .A(n5638), .ZN(n5644) );
  AND2_X1 U7433 ( .A1(SI_21_), .A2(SI_20_), .ZN(n5641) );
  AOI22_X1 U7434 ( .A1(n5644), .A2(n5643), .B1(n5642), .B2(n5641), .ZN(n5645)
         );
  INV_X1 U7435 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7545) );
  MUX2_X1 U7436 ( .A(n7543), .B(n7545), .S(n6779), .Z(n5649) );
  INV_X1 U7437 ( .A(SI_22_), .ZN(n5648) );
  INV_X1 U7438 ( .A(n5649), .ZN(n5650) );
  NAND2_X1 U7439 ( .A1(n5650), .A2(SI_22_), .ZN(n5651) );
  XNOR2_X1 U7440 ( .A(n5669), .B(n5668), .ZN(n7541) );
  NAND2_X1 U7441 ( .A1(n7541), .A2(n8450), .ZN(n5653) );
  OR2_X1 U7442 ( .A1(n8435), .A2(n7543), .ZN(n5652) );
  XNOR2_X1 U7443 ( .A(n8259), .B(n5442), .ZN(n5665) );
  NAND2_X1 U7444 ( .A1(n5654), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n5655) );
  NAND2_X1 U7445 ( .A1(n5691), .A2(n5655), .ZN(n8252) );
  NAND2_X1 U7446 ( .A1(n8252), .A2(n6644), .ZN(n5660) );
  INV_X1 U7447 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n9094) );
  NAND2_X1 U7448 ( .A1(n8457), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n5657) );
  NAND2_X1 U7449 ( .A1(n5369), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n5656) );
  OAI211_X1 U7450 ( .C1(n5368), .C2(n9094), .A(n5657), .B(n5656), .ZN(n5658)
         );
  INV_X1 U7451 ( .A(n5658), .ZN(n5659) );
  XNOR2_X1 U7452 ( .A(n5665), .B(n8724), .ZN(n8248) );
  INV_X1 U7453 ( .A(n8248), .ZN(n5663) );
  INV_X1 U7454 ( .A(n5661), .ZN(n5662) );
  NAND2_X1 U7455 ( .A1(n5662), .A2(n8253), .ZN(n8246) );
  AND2_X1 U7456 ( .A1(n5663), .A2(n8246), .ZN(n5664) );
  NAND2_X1 U7457 ( .A1(n8247), .A2(n5664), .ZN(n8250) );
  NAND2_X1 U7458 ( .A1(n5665), .A2(n8724), .ZN(n5666) );
  INV_X1 U7459 ( .A(n8205), .ZN(n5705) );
  INV_X1 U7460 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n5670) );
  MUX2_X1 U7461 ( .A(n7613), .B(n5670), .S(n6779), .Z(n5672) );
  INV_X1 U7462 ( .A(SI_23_), .ZN(n5671) );
  NAND2_X1 U7463 ( .A1(n5672), .A2(n5671), .ZN(n5675) );
  INV_X1 U7464 ( .A(n5672), .ZN(n5673) );
  NAND2_X1 U7465 ( .A1(n5673), .A2(SI_23_), .ZN(n5674) );
  INV_X1 U7466 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7670) );
  INV_X1 U7467 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7681) );
  MUX2_X1 U7468 ( .A(n7670), .B(n7681), .S(n6779), .Z(n5678) );
  INV_X1 U7469 ( .A(SI_24_), .ZN(n5677) );
  NAND2_X1 U7470 ( .A1(n5678), .A2(n5677), .ZN(n5712) );
  INV_X1 U7471 ( .A(n5678), .ZN(n5679) );
  NAND2_X1 U7472 ( .A1(n5679), .A2(SI_24_), .ZN(n5680) );
  NAND2_X1 U7473 ( .A1(n7669), .A2(n8450), .ZN(n5682) );
  OR2_X1 U7474 ( .A1(n8435), .A2(n7670), .ZN(n5681) );
  XNOR2_X1 U7475 ( .A(n9185), .B(n5442), .ZN(n8208) );
  INV_X1 U7476 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n5683) );
  NAND2_X1 U7477 ( .A1(n5693), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n5685) );
  NAND2_X1 U7478 ( .A1(n5723), .A2(n5685), .ZN(n8714) );
  NAND2_X1 U7479 ( .A1(n8714), .A2(n6644), .ZN(n5690) );
  INV_X1 U7480 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n9184) );
  NAND2_X1 U7481 ( .A1(n5349), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n5687) );
  NAND2_X1 U7482 ( .A1(n8457), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n5686) );
  OAI211_X1 U7483 ( .C1(n9184), .C2(n5429), .A(n5687), .B(n5686), .ZN(n5688)
         );
  INV_X1 U7484 ( .A(n5688), .ZN(n5689) );
  NAND2_X1 U7485 ( .A1(n5691), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5692) );
  NAND2_X1 U7486 ( .A1(n5693), .A2(n5692), .ZN(n8728) );
  NAND2_X1 U7487 ( .A1(n8728), .A2(n6644), .ZN(n5698) );
  INV_X1 U7488 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n9190) );
  NAND2_X1 U7489 ( .A1(n5349), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n5695) );
  NAND2_X1 U7490 ( .A1(n8457), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n5694) );
  OAI211_X1 U7491 ( .C1(n9190), .C2(n5429), .A(n5695), .B(n5694), .ZN(n5696)
         );
  INV_X1 U7492 ( .A(n5696), .ZN(n5697) );
  NAND2_X1 U7493 ( .A1(n7610), .A2(n8450), .ZN(n5702) );
  OR2_X1 U7494 ( .A1(n8435), .A2(n7613), .ZN(n5701) );
  XNOR2_X1 U7495 ( .A(n9191), .B(n5442), .ZN(n5706) );
  OAI22_X1 U7496 ( .A1(n8208), .A2(n8702), .B1(n8712), .B2(n5706), .ZN(n5703)
         );
  INV_X1 U7497 ( .A(n5703), .ZN(n5704) );
  INV_X1 U7498 ( .A(n5706), .ZN(n8206) );
  OAI21_X1 U7499 ( .B1(n8206), .B2(n8734), .A(n8725), .ZN(n5708) );
  NOR2_X1 U7500 ( .A1(n8725), .A2(n8734), .ZN(n5707) );
  AOI22_X1 U7501 ( .A1(n8208), .A2(n5708), .B1(n5707), .B2(n5706), .ZN(n5709)
         );
  INV_X1 U7502 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7711) );
  INV_X1 U7503 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n5714) );
  MUX2_X1 U7504 ( .A(n7711), .B(n5714), .S(n6779), .Z(n5716) );
  INV_X1 U7505 ( .A(SI_25_), .ZN(n5715) );
  NAND2_X1 U7506 ( .A1(n5716), .A2(n5715), .ZN(n6511) );
  INV_X1 U7507 ( .A(n5716), .ZN(n5717) );
  NAND2_X1 U7508 ( .A1(n5717), .A2(SI_25_), .ZN(n5718) );
  NAND2_X1 U7509 ( .A1(n7708), .A2(n8450), .ZN(n5720) );
  OR2_X1 U7510 ( .A1(n8452), .A2(n7711), .ZN(n5719) );
  NAND2_X2 U7511 ( .A1(n5720), .A2(n5719), .ZN(n9178) );
  XNOR2_X1 U7512 ( .A(n9178), .B(n8132), .ZN(n5730) );
  INV_X1 U7513 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n5721) );
  NAND2_X1 U7514 ( .A1(n5723), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n5724) );
  NAND2_X1 U7515 ( .A1(n5741), .A2(n5724), .ZN(n8704) );
  NAND2_X1 U7516 ( .A1(n8704), .A2(n6644), .ZN(n5729) );
  INV_X1 U7517 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n9177) );
  NAND2_X1 U7518 ( .A1(n4272), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n5726) );
  NAND2_X1 U7519 ( .A1(n8457), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n5725) );
  OAI211_X1 U7520 ( .C1(n9177), .C2(n5429), .A(n5726), .B(n5725), .ZN(n5727)
         );
  INV_X1 U7521 ( .A(n5727), .ZN(n5728) );
  XNOR2_X1 U7522 ( .A(n5730), .B(n8687), .ZN(n8175) );
  INV_X1 U7523 ( .A(n5730), .ZN(n5731) );
  INV_X1 U7524 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n7730) );
  INV_X1 U7525 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n5734) );
  MUX2_X1 U7526 ( .A(n7730), .B(n5734), .S(n6779), .Z(n5736) );
  INV_X1 U7527 ( .A(SI_26_), .ZN(n5735) );
  NAND2_X1 U7528 ( .A1(n5736), .A2(n5735), .ZN(n6510) );
  INV_X1 U7529 ( .A(n5736), .ZN(n5737) );
  NAND2_X1 U7530 ( .A1(n5737), .A2(SI_26_), .ZN(n5738) );
  NAND2_X1 U7531 ( .A1(n7727), .A2(n8450), .ZN(n5740) );
  OR2_X1 U7532 ( .A1(n8452), .A2(n7730), .ZN(n5739) );
  XNOR2_X1 U7533 ( .A(n6686), .B(n5442), .ZN(n5747) );
  NAND2_X1 U7534 ( .A1(n5741), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n5742) );
  INV_X1 U7535 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n9170) );
  NAND2_X1 U7536 ( .A1(n5349), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n5744) );
  NAND2_X1 U7537 ( .A1(n8457), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n5743) );
  OAI211_X1 U7538 ( .C1(n9170), .C2(n5429), .A(n5744), .B(n5743), .ZN(n5745)
         );
  INV_X1 U7539 ( .A(n5745), .ZN(n5746) );
  INV_X1 U7540 ( .A(n5747), .ZN(n5748) );
  NAND2_X1 U7541 ( .A1(n5749), .A2(n5748), .ZN(n5750) );
  NAND2_X1 U7542 ( .A1(n5752), .A2(n6515), .ZN(n5753) );
  INV_X1 U7543 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n9284) );
  INV_X1 U7544 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n5754) );
  MUX2_X1 U7545 ( .A(n9284), .B(n5754), .S(n6779), .Z(n5756) );
  INV_X1 U7546 ( .A(SI_27_), .ZN(n5755) );
  NAND2_X1 U7547 ( .A1(n5756), .A2(n5755), .ZN(n6509) );
  INV_X1 U7548 ( .A(n5756), .ZN(n5757) );
  NAND2_X1 U7549 ( .A1(n5757), .A2(SI_27_), .ZN(n6519) );
  AND2_X1 U7550 ( .A1(n6509), .A2(n6519), .ZN(n5758) );
  NAND2_X1 U7551 ( .A1(n9282), .A2(n8450), .ZN(n5761) );
  OR2_X1 U7552 ( .A1(n8452), .A2(n9284), .ZN(n5760) );
  XNOR2_X1 U7553 ( .A(n6689), .B(n5442), .ZN(n8138) );
  INV_X1 U7554 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n5762) );
  NAND2_X1 U7555 ( .A1(n5764), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n5765) );
  NAND2_X1 U7556 ( .A1(n5797), .A2(n5765), .ZN(n8679) );
  NAND2_X1 U7557 ( .A1(n8679), .A2(n6644), .ZN(n5770) );
  INV_X1 U7558 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n9164) );
  NAND2_X1 U7559 ( .A1(n5349), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n5767) );
  NAND2_X1 U7560 ( .A1(n8457), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n5766) );
  OAI211_X1 U7561 ( .C1(n9164), .C2(n5429), .A(n5767), .B(n5766), .ZN(n5768)
         );
  INV_X1 U7562 ( .A(n5768), .ZN(n5769) );
  NAND2_X1 U7563 ( .A1(n8138), .A2(n8686), .ZN(n8135) );
  OAI21_X1 U7564 ( .B1(n8138), .B2(n8686), .A(n8135), .ZN(n5788) );
  INV_X1 U7565 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n6799) );
  NAND2_X1 U7566 ( .A1(n6795), .A2(n6799), .ZN(n5771) );
  NAND2_X1 U7567 ( .A1(n7731), .A2(n7712), .ZN(n6797) );
  NOR2_X1 U7568 ( .A1(P2_D_REG_27__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .ZN(
        n9107) );
  NOR4_X1 U7569 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_2__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n5775) );
  NOR4_X1 U7570 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_12__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n5774) );
  NOR4_X1 U7571 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_22__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n5773) );
  NAND4_X1 U7572 ( .A1(n9107), .A2(n5775), .A3(n5774), .A4(n5773), .ZN(n5781)
         );
  NOR4_X1 U7573 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_21__SCAN_IN), .ZN(n5779) );
  NOR4_X1 U7574 ( .A1(P2_D_REG_23__SCAN_IN), .A2(P2_D_REG_9__SCAN_IN), .A3(
        P2_D_REG_15__SCAN_IN), .A4(P2_D_REG_17__SCAN_IN), .ZN(n5778) );
  NOR4_X1 U7575 ( .A1(P2_D_REG_19__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_6__SCAN_IN), .A4(P2_D_REG_5__SCAN_IN), .ZN(n5777) );
  NOR4_X1 U7576 ( .A1(P2_D_REG_8__SCAN_IN), .A2(P2_D_REG_20__SCAN_IN), .A3(
        P2_D_REG_11__SCAN_IN), .A4(P2_D_REG_10__SCAN_IN), .ZN(n5776) );
  NAND4_X1 U7577 ( .A1(n5779), .A2(n5778), .A3(n5777), .A4(n5776), .ZN(n5780)
         );
  OAI21_X1 U7578 ( .B1(n5781), .B2(n5780), .A(n6795), .ZN(n6716) );
  NAND2_X1 U7579 ( .A1(n6713), .A2(n6716), .ZN(n5807) );
  NOR2_X1 U7580 ( .A1(n5807), .A2(n6715), .ZN(n6730) );
  INV_X1 U7581 ( .A(n8525), .ZN(n7542) );
  AND2_X1 U7582 ( .A1(n8504), .A2(n7396), .ZN(n5782) );
  NAND2_X1 U7583 ( .A1(n6728), .A2(n5782), .ZN(n5806) );
  INV_X1 U7584 ( .A(n5806), .ZN(n5783) );
  NAND2_X1 U7585 ( .A1(n6730), .A2(n5783), .ZN(n5787) );
  INV_X1 U7586 ( .A(n7007), .ZN(n5784) );
  NAND3_X1 U7587 ( .A1(n5784), .A2(n4743), .A3(n6716), .ZN(n5814) );
  NOR2_X1 U7588 ( .A1(n5814), .A2(n6715), .ZN(n6732) );
  INV_X1 U7589 ( .A(n6728), .ZN(n5785) );
  NAND2_X1 U7590 ( .A1(n6732), .A2(n5785), .ZN(n5786) );
  NAND2_X1 U7591 ( .A1(n5787), .A2(n5786), .ZN(n8216) );
  INV_X1 U7592 ( .A(n5788), .ZN(n5789) );
  NAND2_X1 U7593 ( .A1(n6730), .A2(n8998), .ZN(n5791) );
  NOR2_X1 U7594 ( .A1(n6715), .A2(n8295), .ZN(n5790) );
  NAND2_X1 U7595 ( .A1(n4274), .A2(n8525), .ZN(n6720) );
  NAND2_X1 U7596 ( .A1(n8522), .A2(n5792), .ZN(n5793) );
  NAND2_X1 U7597 ( .A1(n5794), .A2(n5793), .ZN(n6708) );
  INV_X1 U7598 ( .A(n6708), .ZN(n5795) );
  NOR2_X1 U7599 ( .A1(n7012), .A2(n5795), .ZN(n5796) );
  NAND2_X1 U7600 ( .A1(n5796), .A2(n6732), .ZN(n8285) );
  NAND2_X1 U7601 ( .A1(n5797), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n5798) );
  NAND2_X1 U7602 ( .A1(n8088), .A2(n5798), .ZN(n8662) );
  NAND2_X1 U7603 ( .A1(n8662), .A2(n6644), .ZN(n5803) );
  INV_X1 U7604 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n9158) );
  NAND2_X1 U7605 ( .A1(n5349), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n5800) );
  NAND2_X1 U7606 ( .A1(n8457), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n5799) );
  OAI211_X1 U7607 ( .C1(n9158), .C2(n5429), .A(n5800), .B(n5799), .ZN(n5801)
         );
  INV_X1 U7608 ( .A(n5801), .ZN(n5802) );
  NOR2_X1 U7609 ( .A1(n7012), .A2(n6708), .ZN(n5804) );
  INV_X1 U7610 ( .A(n5814), .ZN(n5812) );
  NAND2_X1 U7611 ( .A1(n6701), .A2(n8503), .ZN(n5805) );
  NAND2_X1 U7612 ( .A1(n5805), .A2(n8998), .ZN(n10163) );
  NAND2_X1 U7613 ( .A1(n5806), .A2(n10163), .ZN(n6731) );
  NAND2_X1 U7614 ( .A1(n6731), .A2(n5807), .ZN(n5811) );
  NAND2_X1 U7615 ( .A1(n6618), .A2(n8440), .ZN(n6718) );
  AND3_X1 U7616 ( .A1(n6718), .A2(n5809), .A3(n5808), .ZN(n5810) );
  OAI211_X1 U7617 ( .C1(n5812), .C2(n6728), .A(n5811), .B(n5810), .ZN(n5813)
         );
  NAND2_X1 U7618 ( .A1(n5813), .A2(P2_STATE_REG_SCAN_IN), .ZN(n5816) );
  NOR2_X1 U7619 ( .A1(n7012), .A2(n6715), .ZN(n8523) );
  NAND2_X1 U7620 ( .A1(n8523), .A2(n5814), .ZN(n5815) );
  NAND2_X2 U7621 ( .A1(n5816), .A2(n5815), .ZN(n8288) );
  AOI22_X1 U7622 ( .A1(n8679), .A2(n8288), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3151), .ZN(n5817) );
  OAI21_X1 U7623 ( .B1(n8178), .B2(n8266), .A(n5817), .ZN(n5818) );
  AOI21_X1 U7624 ( .B1(n8264), .B2(n8673), .A(n5818), .ZN(n5819) );
  INV_X1 U7625 ( .A(n5820), .ZN(n5821) );
  NAND2_X1 U7626 ( .A1(n5822), .A2(n5821), .ZN(P2_U3154) );
  INV_X2 U7627 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  NOR2_X2 U7628 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_4__SCAN_IN), .ZN(
        n6032) );
  INV_X1 U7629 ( .A(n5844), .ZN(n5833) );
  NOR2_X1 U7630 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), .ZN(
        n5830) );
  NAND4_X1 U7631 ( .A1(n5830), .A2(n5900), .A3(n5863), .A4(n5867), .ZN(n5831)
         );
  NAND2_X1 U7632 ( .A1(n5833), .A2(n5832), .ZN(n5835) );
  NAND2_X1 U7633 ( .A1(n5860), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5834) );
  INV_X1 U7634 ( .A(n5835), .ZN(n5837) );
  NAND2_X1 U7635 ( .A1(n5837), .A2(n5836), .ZN(n5881) );
  BUF_X1 U7636 ( .A(n5881), .Z(n5838) );
  NAND2_X2 U7637 ( .A1(n5838), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5841) );
  NAND2_X2 U7638 ( .A1(n6574), .A2(n6779), .ZN(n6161) );
  BUF_X4 U7639 ( .A(n5907), .Z(n6555) );
  NAND2_X1 U7640 ( .A1(n7541), .A2(n6555), .ZN(n5843) );
  NAND2_X2 U7641 ( .A1(n6574), .A2(n6778), .ZN(n6030) );
  INV_X2 U7642 ( .A(n6030), .ZN(n5988) );
  NAND2_X1 U7643 ( .A1(n5988), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n5842) );
  INV_X1 U7644 ( .A(n5846), .ZN(n5847) );
  NAND2_X1 U7645 ( .A1(n5847), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5848) );
  NAND2_X1 U7646 ( .A1(n5894), .A2(n5848), .ZN(n5853) );
  INV_X1 U7647 ( .A(n5853), .ZN(n5850) );
  INV_X1 U7648 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5849) );
  NAND2_X1 U7649 ( .A1(n5850), .A2(n5849), .ZN(n5855) );
  INV_X1 U7650 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5851) );
  NAND2_X1 U7651 ( .A1(n5853), .A2(P1_IR_REG_20__SCAN_IN), .ZN(n5854) );
  NAND2_X1 U7652 ( .A1(n5863), .A2(n5867), .ZN(n5858) );
  OAI21_X1 U7653 ( .B1(n5861), .B2(n5858), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n5859) );
  INV_X1 U7654 ( .A(n5864), .ZN(n5862) );
  NAND2_X1 U7655 ( .A1(n5862), .A2(P1_IR_REG_24__SCAN_IN), .ZN(n5865) );
  INV_X1 U7656 ( .A(n6738), .ZN(n5870) );
  OR2_X2 U7657 ( .A1(n6097), .A2(n6096), .ZN(n6099) );
  INV_X1 U7658 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n6264) );
  OR2_X2 U7659 ( .A1(n6265), .A2(n6264), .ZN(n6299) );
  AND2_X1 U7660 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(P1_REG3_REG_19__SCAN_IN), 
        .ZN(n5877) );
  INV_X1 U7661 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n6320) );
  INV_X1 U7662 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n9038) );
  OR2_X2 U7663 ( .A1(n6343), .A2(n9038), .ZN(n6359) );
  NAND2_X1 U7664 ( .A1(n6343), .A2(n9038), .ZN(n5880) );
  NAND2_X1 U7665 ( .A1(n6359), .A2(n5880), .ZN(n9691) );
  NOR2_X2 U7666 ( .A1(n5881), .A2(P1_IR_REG_28__SCAN_IN), .ZN(n5885) );
  INV_X1 U7667 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n5882) );
  NAND2_X1 U7668 ( .A1(n5885), .A2(n5882), .ZN(n9881) );
  XNOR2_X2 U7669 ( .A(n5883), .B(P1_IR_REG_30__SCAN_IN), .ZN(n9885) );
  OR2_X2 U7670 ( .A1(n5885), .A2(n5884), .ZN(n5886) );
  OR2_X1 U7671 ( .A1(n9691), .A2(n6442), .ZN(n5893) );
  INV_X1 U7672 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n9115) );
  BUF_X4 U7673 ( .A(n5994), .Z(n6563) );
  NAND2_X1 U7674 ( .A1(n7878), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n5890) );
  INV_X1 U7675 ( .A(n9885), .ZN(n5888) );
  AND2_X2 U7676 ( .A1(n5888), .A2(n9888), .ZN(n6041) );
  NAND2_X1 U7678 ( .A1(n6486), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n5889) );
  OAI211_X1 U7679 ( .C1(n7881), .C2(n9115), .A(n5890), .B(n5889), .ZN(n5891)
         );
  INV_X1 U7680 ( .A(n5891), .ZN(n5892) );
  INV_X1 U7681 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n6278) );
  NAND2_X1 U7682 ( .A1(n5894), .A2(n6278), .ZN(n6280) );
  NAND2_X1 U7683 ( .A1(n6280), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5895) );
  INV_X2 U7684 ( .A(n5897), .ZN(n6294) );
  AND2_X2 U7685 ( .A1(n6294), .A2(n6480), .ZN(n6478) );
  INV_X1 U7686 ( .A(n5898), .ZN(n5899) );
  NAND2_X1 U7687 ( .A1(n5899), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5901) );
  NOR2_X1 U7688 ( .A1(n9709), .A2(n4423), .ZN(n5903) );
  AOI21_X1 U7689 ( .B1(n9819), .B2(n6423), .A(n5903), .ZN(n7769) );
  NAND2_X1 U7690 ( .A1(n6294), .A2(n7886), .ZN(n6996) );
  OAI22_X1 U7691 ( .A1(n9695), .A2(n9334), .B1(n9709), .B2(n6389), .ZN(n5906)
         );
  XNOR2_X1 U7692 ( .A(n5906), .B(n9335), .ZN(n7756) );
  NAND2_X1 U7693 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5908) );
  INV_X1 U7694 ( .A(n6780), .ZN(n9505) );
  NAND2_X1 U7695 ( .A1(n4273), .A2(n7903), .ZN(n5919) );
  INV_X1 U7696 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n9502) );
  INV_X1 U7697 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n5913) );
  INV_X1 U7698 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n5914) );
  NAND2_X1 U7699 ( .A1(n5871), .A2(n7903), .ZN(n5920) );
  OAI21_X1 U7700 ( .B1(n9337), .B2(n10049), .A(n5920), .ZN(n5945) );
  INV_X1 U7701 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n10067) );
  INV_X1 U7702 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n5921) );
  INV_X1 U7703 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n5922) );
  OR2_X1 U7704 ( .A1(n5991), .A2(n5922), .ZN(n5923) );
  INV_X1 U7705 ( .A(n7346), .ZN(n5927) );
  NOR2_X1 U7706 ( .A1(n6778), .A2(n5928), .ZN(n5930) );
  XNOR2_X1 U7707 ( .A(n5930), .B(n5929), .ZN(n9899) );
  MUX2_X1 U7708 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9899), .S(n6574), .Z(n10058)
         );
  NAND2_X1 U7709 ( .A1(n4273), .A2(n10058), .ZN(n5932) );
  INV_X1 U7710 ( .A(n5933), .ZN(n5942) );
  INV_X1 U7711 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n5934) );
  OR2_X1 U7712 ( .A1(n6738), .A2(n5934), .ZN(n5935) );
  NAND2_X1 U7713 ( .A1(n5871), .A2(n10058), .ZN(n5941) );
  OR2_X1 U7714 ( .A1(n6738), .A2(n5936), .ZN(n5937) );
  NAND2_X1 U7715 ( .A1(n5941), .A2(n5940), .ZN(n6975) );
  NAND2_X1 U7716 ( .A1(n5942), .A2(n9335), .ZN(n5943) );
  NAND2_X1 U7717 ( .A1(n7112), .A2(n7111), .ZN(n5948) );
  NAND2_X1 U7718 ( .A1(n5948), .A2(n5947), .ZN(n7117) );
  OR2_X1 U7719 ( .A1(n6789), .A2(n6161), .ZN(n5951) );
  AOI22_X1 U7720 ( .A1(n5988), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(n6295), .B2(
        n4431), .ZN(n5950) );
  AND2_X2 U7721 ( .A1(n5951), .A2(n5950), .ZN(n10086) );
  INV_X1 U7722 ( .A(n10086), .ZN(n7353) );
  NAND2_X1 U7723 ( .A1(n5931), .A2(n7353), .ZN(n5959) );
  INV_X1 U7724 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n10043) );
  INV_X1 U7725 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n5952) );
  INV_X1 U7726 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n5953) );
  NAND2_X1 U7727 ( .A1(n6423), .A2(n7352), .ZN(n5958) );
  NAND2_X1 U7728 ( .A1(n5959), .A2(n5958), .ZN(n5960) );
  INV_X1 U7729 ( .A(n7352), .ZN(n5961) );
  NAND2_X1 U7730 ( .A1(n6423), .A2(n7353), .ZN(n5962) );
  NAND2_X1 U7731 ( .A1(n5963), .A2(n5962), .ZN(n5964) );
  XNOR2_X1 U7732 ( .A(n5966), .B(n5964), .ZN(n7116) );
  NAND2_X1 U7733 ( .A1(n7117), .A2(n7116), .ZN(n5968) );
  INV_X1 U7734 ( .A(n5964), .ZN(n5965) );
  NAND2_X1 U7735 ( .A1(n5966), .A2(n5965), .ZN(n5967) );
  NAND2_X1 U7736 ( .A1(n5968), .A2(n5967), .ZN(n7146) );
  AOI22_X1 U7737 ( .A1(n5988), .A2(P2_DATAO_REG_3__SCAN_IN), .B1(n6295), .B2(
        n9535), .ZN(n5972) );
  NAND2_X1 U7738 ( .A1(n5931), .A2(n7493), .ZN(n5979) );
  OR2_X1 U7739 ( .A1(n6442), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n5977) );
  INV_X1 U7740 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n5973) );
  OR2_X1 U7741 ( .A1(n5991), .A2(n5973), .ZN(n5976) );
  INV_X1 U7742 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n7496) );
  OR2_X1 U7743 ( .A1(n6563), .A2(n7496), .ZN(n5975) );
  NAND2_X1 U7744 ( .A1(n6423), .A2(n10011), .ZN(n5978) );
  NAND2_X1 U7745 ( .A1(n5979), .A2(n5978), .ZN(n5980) );
  XNOR2_X1 U7746 ( .A(n5980), .B(n9335), .ZN(n5984) );
  NAND2_X1 U7747 ( .A1(n6423), .A2(n7493), .ZN(n5981) );
  OAI21_X1 U7748 ( .B1(n9337), .B2(n7344), .A(n5981), .ZN(n5982) );
  XNOR2_X1 U7749 ( .A(n5984), .B(n5982), .ZN(n7147) );
  INV_X1 U7750 ( .A(n5982), .ZN(n5983) );
  NAND2_X1 U7751 ( .A1(n5984), .A2(n5983), .ZN(n5985) );
  AOI22_X1 U7752 ( .A1(n5988), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n6295), .B2(
        n4422), .ZN(n5989) );
  NAND2_X1 U7753 ( .A1(n5931), .A2(n10018), .ZN(n5999) );
  NAND2_X1 U7754 ( .A1(n6060), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5997) );
  OAI21_X1 U7755 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(n6014), .ZN(n10014) );
  INV_X1 U7756 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n5993) );
  OR2_X1 U7757 ( .A1(n6563), .A2(n5993), .ZN(n5995) );
  NAND2_X1 U7758 ( .A1(n9500), .A2(n6423), .ZN(n5998) );
  NAND2_X1 U7759 ( .A1(n5999), .A2(n5998), .ZN(n6001) );
  XNOR2_X1 U7760 ( .A(n6001), .B(n6426), .ZN(n6004) );
  NAND2_X1 U7761 ( .A1(n6423), .A2(n10018), .ZN(n6002) );
  OAI21_X1 U7762 ( .B1(n4423), .B2(n7356), .A(n6002), .ZN(n6003) );
  XNOR2_X1 U7763 ( .A(n6004), .B(n6003), .ZN(n9393) );
  NAND2_X1 U7764 ( .A1(n6004), .A2(n6003), .ZN(n6005) );
  INV_X1 U7765 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n6006) );
  NAND2_X1 U7766 ( .A1(n6007), .A2(n6006), .ZN(n6008) );
  NAND2_X1 U7767 ( .A1(n6008), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6009) );
  XNOR2_X2 U7768 ( .A(n6009), .B(P1_IR_REG_5__SCAN_IN), .ZN(n6908) );
  AOI22_X1 U7769 ( .A1(n5988), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n6295), .B2(
        n6908), .ZN(n6010) );
  NAND2_X1 U7770 ( .A1(n6398), .A2(n7592), .ZN(n6021) );
  NAND2_X1 U7771 ( .A1(n6323), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6019) );
  INV_X1 U7772 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n6012) );
  OR2_X1 U7773 ( .A1(n7881), .A2(n6012), .ZN(n6018) );
  INV_X1 U7774 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n6013) );
  NAND2_X1 U7775 ( .A1(n6014), .A2(n6013), .ZN(n6015) );
  NAND2_X1 U7776 ( .A1(n6039), .A2(n6015), .ZN(n7590) );
  OR2_X1 U7777 ( .A1(n6442), .A2(n7590), .ZN(n6017) );
  INV_X1 U7778 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n7589) );
  OR2_X1 U7779 ( .A1(n6563), .A2(n7589), .ZN(n6016) );
  NAND2_X1 U7780 ( .A1(n7358), .A2(n6423), .ZN(n6020) );
  NAND2_X1 U7781 ( .A1(n6021), .A2(n6020), .ZN(n6022) );
  XNOR2_X1 U7782 ( .A(n6022), .B(n6426), .ZN(n6026) );
  NAND2_X1 U7783 ( .A1(n7358), .A2(n6421), .ZN(n6024) );
  NAND2_X1 U7784 ( .A1(n7592), .A2(n4391), .ZN(n6023) );
  AND2_X1 U7785 ( .A1(n6024), .A2(n6023), .ZN(n7314) );
  NAND2_X1 U7786 ( .A1(n7312), .A2(n7314), .ZN(n6029) );
  INV_X1 U7787 ( .A(n6026), .ZN(n6027) );
  NAND2_X1 U7788 ( .A1(n6793), .A2(n6555), .ZN(n6036) );
  INV_X2 U7789 ( .A(n6030), .ZN(n6556) );
  INV_X1 U7790 ( .A(n6031), .ZN(n6033) );
  NAND2_X1 U7791 ( .A1(n6033), .A2(n6032), .ZN(n6056) );
  NAND2_X1 U7792 ( .A1(n6056), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6034) );
  AOI22_X1 U7793 ( .A1(n6556), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n6295), .B2(
        n6925), .ZN(n6035) );
  NAND2_X1 U7794 ( .A1(n6398), .A2(n10001), .ZN(n6048) );
  INV_X1 U7795 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n6037) );
  OR2_X1 U7796 ( .A1(n6563), .A2(n6037), .ZN(n6046) );
  INV_X1 U7797 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n6038) );
  NAND2_X1 U7798 ( .A1(n6039), .A2(n6038), .ZN(n6040) );
  NAND2_X1 U7799 ( .A1(n6062), .A2(n6040), .ZN(n9994) );
  OR2_X1 U7800 ( .A1(n6442), .A2(n9994), .ZN(n6045) );
  INV_X1 U7801 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n6042) );
  OR2_X1 U7802 ( .A1(n7247), .A2(n6042), .ZN(n6044) );
  NAND2_X1 U7803 ( .A1(n6060), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n6043) );
  NAND2_X1 U7805 ( .A1(n9499), .A2(n4391), .ZN(n6047) );
  NAND2_X1 U7806 ( .A1(n6048), .A2(n6047), .ZN(n6049) );
  XNOR2_X1 U7807 ( .A(n6049), .B(n9335), .ZN(n7325) );
  NAND2_X1 U7808 ( .A1(n9499), .A2(n6421), .ZN(n6051) );
  NAND2_X1 U7809 ( .A1(n10001), .A2(n4391), .ZN(n6050) );
  AND2_X1 U7810 ( .A1(n6051), .A2(n6050), .ZN(n7324) );
  AND2_X1 U7811 ( .A1(n7325), .A2(n7324), .ZN(n6052) );
  INV_X1 U7812 ( .A(n7325), .ZN(n6054) );
  INV_X1 U7813 ( .A(n7324), .ZN(n6053) );
  NAND2_X1 U7814 ( .A1(n6054), .A2(n6053), .ZN(n6055) );
  OR2_X1 U7815 ( .A1(n6792), .A2(n6161), .ZN(n6059) );
  NAND2_X1 U7816 ( .A1(n6118), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6057) );
  AOI22_X1 U7817 ( .A1(n6556), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n6295), .B2(
        n6936), .ZN(n6058) );
  NAND2_X1 U7818 ( .A1(n6398), .A2(n7429), .ZN(n6069) );
  NAND2_X1 U7819 ( .A1(n6060), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n6067) );
  INV_X1 U7820 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n6591) );
  OR2_X1 U7821 ( .A1(n7247), .A2(n6591), .ZN(n6066) );
  INV_X1 U7822 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n6061) );
  NAND2_X1 U7823 ( .A1(n6062), .A2(n6061), .ZN(n6063) );
  NAND2_X1 U7824 ( .A1(n6097), .A2(n6063), .ZN(n7433) );
  OR2_X1 U7825 ( .A1(n6442), .A2(n7433), .ZN(n6065) );
  INV_X1 U7826 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n6579) );
  OR2_X1 U7827 ( .A1(n6563), .A2(n6579), .ZN(n6064) );
  INV_X1 U7828 ( .A(n9975), .ZN(n9992) );
  NAND2_X1 U7829 ( .A1(n9992), .A2(n4391), .ZN(n6068) );
  NAND2_X1 U7830 ( .A1(n6069), .A2(n6068), .ZN(n6070) );
  XNOR2_X1 U7831 ( .A(n6070), .B(n6426), .ZN(n6075) );
  INV_X1 U7832 ( .A(n6075), .ZN(n6073) );
  NAND2_X1 U7833 ( .A1(n4391), .A2(n7429), .ZN(n6071) );
  OAI21_X1 U7834 ( .B1(n4423), .B2(n9975), .A(n6071), .ZN(n6074) );
  INV_X1 U7835 ( .A(n6074), .ZN(n6072) );
  NAND2_X1 U7836 ( .A1(n6073), .A2(n6072), .ZN(n7424) );
  AND2_X1 U7837 ( .A1(n6075), .A2(n6074), .ZN(n7425) );
  OAI21_X1 U7838 ( .B1(n6118), .B2(P1_IR_REG_7__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6091) );
  INV_X1 U7839 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n6119) );
  NAND2_X1 U7840 ( .A1(n6091), .A2(n6119), .ZN(n6093) );
  NAND2_X1 U7841 ( .A1(n6093), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6077) );
  XNOR2_X1 U7842 ( .A(n6077), .B(P1_IR_REG_9__SCAN_IN), .ZN(n9572) );
  AOI22_X1 U7843 ( .A1(n9572), .A2(n6295), .B1(n6556), .B2(
        P2_DATAO_REG_9__SCAN_IN), .ZN(n6078) );
  NAND2_X2 U7844 ( .A1(n6079), .A2(n6078), .ZN(n9407) );
  NAND2_X1 U7845 ( .A1(n9407), .A2(n6398), .ZN(n6087) );
  NAND2_X1 U7846 ( .A1(n6060), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n6085) );
  INV_X1 U7847 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n6592) );
  OR2_X1 U7848 ( .A1(n7247), .A2(n6592), .ZN(n6084) );
  INV_X1 U7849 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n7511) );
  OR2_X1 U7850 ( .A1(n6563), .A2(n7511), .ZN(n6083) );
  INV_X1 U7851 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n6080) );
  NAND2_X1 U7852 ( .A1(n6099), .A2(n6080), .ZN(n6081) );
  NAND2_X1 U7853 ( .A1(n6145), .A2(n6081), .ZN(n9408) );
  OR2_X1 U7854 ( .A1(n6442), .A2(n9408), .ZN(n6082) );
  NAND2_X1 U7855 ( .A1(n9497), .A2(n4391), .ZN(n6086) );
  NAND2_X1 U7856 ( .A1(n6087), .A2(n6086), .ZN(n6088) );
  XNOR2_X1 U7857 ( .A(n6088), .B(n6426), .ZN(n6112) );
  NAND2_X1 U7858 ( .A1(n9407), .A2(n4391), .ZN(n6090) );
  NAND2_X1 U7859 ( .A1(n9497), .A2(n6421), .ZN(n6089) );
  NAND2_X1 U7860 ( .A1(n6090), .A2(n6089), .ZN(n9403) );
  OR2_X1 U7861 ( .A1(n6091), .A2(n6119), .ZN(n6092) );
  AOI22_X1 U7862 ( .A1(n6556), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n6295), .B2(
        n6948), .ZN(n6094) );
  NAND2_X1 U7863 ( .A1(n10122), .A2(n4391), .ZN(n6107) );
  NAND2_X1 U7864 ( .A1(n6323), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6105) );
  NAND2_X1 U7865 ( .A1(n6097), .A2(n6096), .ZN(n6098) );
  NAND2_X1 U7866 ( .A1(n6099), .A2(n6098), .ZN(n9982) );
  OR2_X1 U7867 ( .A1(n6442), .A2(n9982), .ZN(n6104) );
  INV_X1 U7868 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n6100) );
  OR2_X1 U7869 ( .A1(n6563), .A2(n6100), .ZN(n6103) );
  INV_X1 U7870 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n6101) );
  OR2_X1 U7871 ( .A1(n7881), .A2(n6101), .ZN(n6102) );
  NAND2_X1 U7872 ( .A1(n9498), .A2(n6421), .ZN(n6106) );
  NAND2_X1 U7873 ( .A1(n6107), .A2(n6106), .ZN(n7672) );
  NAND2_X1 U7874 ( .A1(n10122), .A2(n6398), .ZN(n6109) );
  NAND2_X1 U7875 ( .A1(n9498), .A2(n4391), .ZN(n6108) );
  NAND2_X1 U7876 ( .A1(n6109), .A2(n6108), .ZN(n6110) );
  XNOR2_X1 U7877 ( .A(n6110), .B(n6426), .ZN(n6113) );
  AOI22_X1 U7878 ( .A1(n6112), .A2(n9403), .B1(n7672), .B2(n6113), .ZN(n6111)
         );
  NAND2_X1 U7879 ( .A1(n9401), .A2(n6111), .ZN(n6117) );
  INV_X1 U7880 ( .A(n6112), .ZN(n9404) );
  OAI21_X1 U7881 ( .B1(n6113), .B2(n7672), .A(n9403), .ZN(n6115) );
  NOR2_X1 U7882 ( .A1(n9403), .A2(n7672), .ZN(n6114) );
  INV_X1 U7883 ( .A(n6113), .ZN(n9402) );
  AOI22_X1 U7884 ( .A1(n9404), .A2(n6115), .B1(n6114), .B2(n9402), .ZN(n6116)
         );
  NAND2_X1 U7885 ( .A1(n6117), .A2(n6116), .ZN(n9307) );
  NAND2_X1 U7886 ( .A1(n6835), .A2(n6555), .ZN(n6125) );
  INV_X1 U7887 ( .A(n6118), .ZN(n6122) );
  INV_X1 U7888 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n6120) );
  INV_X1 U7889 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n9022) );
  AND3_X1 U7890 ( .A1(n6120), .A2(n9022), .A3(n6119), .ZN(n6121) );
  NAND2_X1 U7891 ( .A1(n6122), .A2(n6121), .ZN(n6138) );
  NAND2_X1 U7892 ( .A1(n6163), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6123) );
  XNOR2_X1 U7893 ( .A(n6123), .B(P1_IR_REG_11__SCAN_IN), .ZN(n6745) );
  AOI22_X1 U7894 ( .A1(n6556), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n6745), .B2(
        n6295), .ZN(n6124) );
  NAND2_X1 U7895 ( .A1(n9445), .A2(n6398), .ZN(n6134) );
  NAND2_X1 U7896 ( .A1(n6323), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n6132) );
  INV_X1 U7897 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n7411) );
  OR2_X1 U7898 ( .A1(n6563), .A2(n7411), .ZN(n6131) );
  INV_X1 U7899 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n6144) );
  INV_X1 U7900 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n6126) );
  OAI21_X1 U7901 ( .B1(n6145), .B2(n6144), .A(n6126), .ZN(n6127) );
  NAND2_X1 U7902 ( .A1(n6127), .A2(n6169), .ZN(n9442) );
  OR2_X1 U7903 ( .A1(n6442), .A2(n9442), .ZN(n6130) );
  INV_X1 U7904 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n6128) );
  OR2_X1 U7905 ( .A1(n7881), .A2(n6128), .ZN(n6129) );
  NAND4_X1 U7906 ( .A1(n6132), .A2(n6131), .A3(n6130), .A4(n6129), .ZN(n9495)
         );
  NAND2_X1 U7907 ( .A1(n4391), .A2(n9495), .ZN(n6133) );
  NAND2_X1 U7908 ( .A1(n6134), .A2(n6133), .ZN(n6135) );
  XNOR2_X1 U7909 ( .A(n6135), .B(n6426), .ZN(n9436) );
  NAND2_X1 U7910 ( .A1(n9445), .A2(n4391), .ZN(n6137) );
  NAND2_X1 U7911 ( .A1(n6421), .A2(n9495), .ZN(n6136) );
  NAND2_X1 U7912 ( .A1(n6137), .A2(n6136), .ZN(n6156) );
  OR2_X1 U7913 ( .A1(n6825), .A2(n6161), .ZN(n6142) );
  NAND2_X1 U7914 ( .A1(n6138), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6139) );
  MUX2_X1 U7915 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6139), .S(
        P1_IR_REG_10__SCAN_IN), .Z(n6140) );
  AOI22_X1 U7916 ( .A1(n6556), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n6770), .B2(
        n6295), .ZN(n6141) );
  NAND2_X1 U7917 ( .A1(n6486), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n6149) );
  INV_X1 U7918 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n6143) );
  OR2_X1 U7919 ( .A1(n7881), .A2(n6143), .ZN(n6148) );
  XNOR2_X1 U7920 ( .A(n6145), .B(n6144), .ZN(n9312) );
  OR2_X1 U7921 ( .A1(n6442), .A2(n9312), .ZN(n6147) );
  INV_X1 U7922 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n7563) );
  OR2_X1 U7923 ( .A1(n6563), .A2(n7563), .ZN(n6146) );
  NAND4_X1 U7924 ( .A1(n6149), .A2(n6148), .A3(n6147), .A4(n6146), .ZN(n9496)
         );
  INV_X1 U7925 ( .A(n9496), .ZN(n7506) );
  OAI22_X1 U7926 ( .A1(n10140), .A2(n6389), .B1(n7506), .B2(n4423), .ZN(n9309)
         );
  OAI22_X1 U7927 ( .A1(n10140), .A2(n9334), .B1(n7506), .B2(n6389), .ZN(n6151)
         );
  XNOR2_X1 U7928 ( .A(n6151), .B(n6426), .ZN(n6153) );
  AOI22_X1 U7929 ( .A1(n9436), .A2(n6156), .B1(n9309), .B2(n6153), .ZN(n6152)
         );
  INV_X1 U7930 ( .A(n9436), .ZN(n6159) );
  INV_X1 U7931 ( .A(n6153), .ZN(n9434) );
  INV_X1 U7932 ( .A(n9309), .ZN(n6154) );
  NAND2_X1 U7933 ( .A1(n9434), .A2(n6154), .ZN(n6155) );
  NAND2_X1 U7934 ( .A1(n6155), .A2(n6156), .ZN(n6158) );
  INV_X1 U7935 ( .A(n6155), .ZN(n6157) );
  INV_X1 U7936 ( .A(n6156), .ZN(n9435) );
  AOI22_X1 U7937 ( .A1(n6159), .A2(n6158), .B1(n6157), .B2(n9435), .ZN(n6160)
         );
  INV_X1 U7938 ( .A(n6842), .ZN(n6162) );
  NAND2_X1 U7939 ( .A1(n6162), .A2(n6555), .ZN(n6168) );
  OAI21_X1 U7940 ( .B1(n6163), .B2(P1_IR_REG_11__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6165) );
  INV_X1 U7941 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n6164) );
  OR2_X1 U7942 ( .A1(n6165), .A2(n6164), .ZN(n6166) );
  NAND2_X1 U7943 ( .A1(n6165), .A2(n6164), .ZN(n6181) );
  AOI22_X1 U7944 ( .A1(n7305), .A2(n6295), .B1(n6556), .B2(
        P2_DATAO_REG_12__SCAN_IN), .ZN(n6167) );
  NAND2_X1 U7945 ( .A1(n6060), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n6174) );
  INV_X1 U7946 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n6594) );
  OR2_X1 U7947 ( .A1(n7247), .A2(n6594), .ZN(n6173) );
  INV_X1 U7948 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n9032) );
  NAND2_X1 U7949 ( .A1(n6169), .A2(n9032), .ZN(n6170) );
  NAND2_X1 U7950 ( .A1(n6236), .A2(n6170), .ZN(n7703) );
  OR2_X1 U7951 ( .A1(n6442), .A2(n7703), .ZN(n6172) );
  INV_X1 U7952 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n7570) );
  OR2_X1 U7953 ( .A1(n6563), .A2(n7570), .ZN(n6171) );
  NAND4_X1 U7954 ( .A1(n6174), .A2(n6173), .A3(n6172), .A4(n6171), .ZN(n9494)
         );
  INV_X1 U7955 ( .A(n9494), .ZN(n7459) );
  OAI22_X1 U7956 ( .A1(n7461), .A2(n9334), .B1(n7459), .B2(n6389), .ZN(n6175)
         );
  XNOR2_X1 U7957 ( .A(n6175), .B(n9335), .ZN(n6178) );
  OAI22_X1 U7958 ( .A1(n7461), .A2(n6389), .B1(n7459), .B2(n4423), .ZN(n6176)
         );
  XNOR2_X1 U7959 ( .A(n6178), .B(n6176), .ZN(n7698) );
  INV_X1 U7960 ( .A(n6176), .ZN(n6177) );
  NAND2_X1 U7961 ( .A1(n6178), .A2(n6177), .ZN(n6179) );
  NAND2_X1 U7962 ( .A1(n6180), .A2(n6555), .ZN(n6184) );
  NAND2_X1 U7963 ( .A1(n6181), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6182) );
  XNOR2_X1 U7964 ( .A(n6182), .B(P1_IR_REG_13__SCAN_IN), .ZN(n6758) );
  AOI22_X1 U7965 ( .A1(n6758), .A2(n6295), .B1(n6556), .B2(
        P2_DATAO_REG_13__SCAN_IN), .ZN(n6183) );
  NAND2_X1 U7966 ( .A1(n9430), .A2(n6398), .ZN(n6191) );
  NAND2_X1 U7967 ( .A1(n6486), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n6189) );
  INV_X1 U7968 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n7620) );
  OR2_X1 U7969 ( .A1(n6563), .A2(n7620), .ZN(n6188) );
  XNOR2_X1 U7970 ( .A(n6236), .B(n6235), .ZN(n9428) );
  OR2_X1 U7971 ( .A1(n6442), .A2(n9428), .ZN(n6187) );
  INV_X1 U7972 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n6185) );
  OR2_X1 U7973 ( .A1(n7881), .A2(n6185), .ZN(n6186) );
  INV_X1 U7974 ( .A(n7700), .ZN(n9493) );
  NAND2_X1 U7975 ( .A1(n9493), .A2(n4391), .ZN(n6190) );
  NAND2_X1 U7976 ( .A1(n6191), .A2(n6190), .ZN(n6192) );
  XNOR2_X1 U7977 ( .A(n6192), .B(n6426), .ZN(n6194) );
  NOR2_X1 U7978 ( .A1(n4423), .A2(n7700), .ZN(n6193) );
  AOI21_X1 U7979 ( .B1(n9430), .B2(n6423), .A(n6193), .ZN(n6195) );
  XNOR2_X1 U7980 ( .A(n6194), .B(n6195), .ZN(n9423) );
  NAND2_X1 U7981 ( .A1(n9422), .A2(n9423), .ZN(n6198) );
  INV_X1 U7982 ( .A(n6194), .ZN(n6196) );
  NAND2_X1 U7983 ( .A1(n6196), .A2(n6195), .ZN(n6197) );
  NAND2_X1 U7984 ( .A1(n7157), .A2(n6555), .ZN(n6204) );
  NAND2_X1 U7985 ( .A1(n6199), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6200) );
  MUX2_X1 U7986 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6200), .S(
        P1_IR_REG_16__SCAN_IN), .Z(n6202) );
  AND2_X1 U7987 ( .A1(n6202), .A2(n6260), .ZN(n7159) );
  AOI22_X1 U7988 ( .A1(n6556), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n6295), .B2(
        n7159), .ZN(n6203) );
  NAND2_X1 U7989 ( .A1(n9848), .A2(n6398), .ZN(n6211) );
  AOI22_X1 U7990 ( .A1(n6060), .A2(P1_REG0_REG_16__SCAN_IN), .B1(n6486), .B2(
        P1_REG1_REG_16__SCAN_IN), .ZN(n6209) );
  INV_X1 U7991 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n6205) );
  NAND2_X1 U7992 ( .A1(n6221), .A2(n6205), .ZN(n6206) );
  NAND2_X1 U7993 ( .A1(n6265), .A2(n6206), .ZN(n9379) );
  OR2_X1 U7994 ( .A1(n9379), .A2(n6442), .ZN(n6208) );
  INV_X1 U7995 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n7721) );
  OR2_X1 U7996 ( .A1(n6563), .A2(n7721), .ZN(n6207) );
  INV_X1 U7997 ( .A(n9476), .ZN(n9771) );
  NAND2_X1 U7998 ( .A1(n9771), .A2(n4391), .ZN(n6210) );
  NAND2_X1 U7999 ( .A1(n6211), .A2(n6210), .ZN(n6212) );
  XNOR2_X1 U8000 ( .A(n6212), .B(n6426), .ZN(n9374) );
  NAND2_X1 U8001 ( .A1(n9848), .A2(n4391), .ZN(n6214) );
  NAND2_X1 U8002 ( .A1(n9771), .A2(n6421), .ZN(n6213) );
  NAND2_X1 U8003 ( .A1(n6214), .A2(n6213), .ZN(n9373) );
  NAND2_X1 U8004 ( .A1(n7106), .A2(n6555), .ZN(n6219) );
  OR2_X1 U8005 ( .A1(n6215), .A2(n5884), .ZN(n6217) );
  XNOR2_X1 U8006 ( .A(n6217), .B(n6216), .ZN(n7107) );
  INV_X1 U8007 ( .A(n7107), .ZN(n9921) );
  AOI22_X1 U8008 ( .A1(n6556), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n6295), .B2(
        n9921), .ZN(n6218) );
  OR2_X1 U8009 ( .A1(n9486), .A2(n6389), .ZN(n6227) );
  INV_X1 U8010 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n9128) );
  NAND2_X1 U8011 ( .A1(n6237), .A2(n9128), .ZN(n6220) );
  NAND2_X1 U8012 ( .A1(n6221), .A2(n6220), .ZN(n9478) );
  OR2_X1 U8013 ( .A1(n9478), .A2(n6442), .ZN(n6225) );
  NAND2_X1 U8014 ( .A1(n6060), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n6224) );
  INV_X1 U8015 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n9917) );
  OR2_X1 U8016 ( .A1(n7247), .A2(n9917), .ZN(n6223) );
  NAND2_X1 U8017 ( .A1(n7878), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n6222) );
  NAND2_X1 U8018 ( .A1(n9491), .A2(n6421), .ZN(n6226) );
  NAND2_X1 U8019 ( .A1(n6227), .A2(n6226), .ZN(n6249) );
  OAI22_X1 U8020 ( .A1(n9486), .A2(n9334), .B1(n9291), .B2(n6389), .ZN(n6228)
         );
  XNOR2_X1 U8021 ( .A(n6228), .B(n6426), .ZN(n9371) );
  AOI22_X1 U8022 ( .A1(n9374), .A2(n9373), .B1(n6249), .B2(n9371), .ZN(n6255)
         );
  NAND2_X1 U8023 ( .A1(n6957), .A2(n6555), .ZN(n6233) );
  NAND2_X1 U8024 ( .A1(n4385), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6229) );
  MUX2_X1 U8025 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6229), .S(
        P1_IR_REG_14__SCAN_IN), .Z(n6230) );
  INV_X1 U8026 ( .A(n6230), .ZN(n6231) );
  NOR2_X1 U8027 ( .A1(n6231), .A2(n6215), .ZN(n9908) );
  AOI22_X1 U8028 ( .A1(n6556), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n6295), .B2(
        n9908), .ZN(n6232) );
  NAND2_X1 U8029 ( .A1(n6486), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n6244) );
  OAI21_X1 U8030 ( .B1(n6236), .B2(n6235), .A(n6234), .ZN(n6238) );
  NAND2_X1 U8031 ( .A1(n6238), .A2(n6237), .ZN(n9294) );
  OR2_X1 U8032 ( .A1(n9294), .A2(n6442), .ZN(n6243) );
  INV_X1 U8033 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n6239) );
  OR2_X1 U8034 ( .A1(n6563), .A2(n6239), .ZN(n6242) );
  INV_X1 U8035 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n6240) );
  OR2_X1 U8036 ( .A1(n7881), .A2(n6240), .ZN(n6241) );
  OAI22_X1 U8037 ( .A1(n7685), .A2(n9334), .B1(n9425), .B2(n6389), .ZN(n6245)
         );
  XNOR2_X1 U8038 ( .A(n6245), .B(n6426), .ZN(n9366) );
  OR2_X1 U8039 ( .A1(n7685), .A2(n6389), .ZN(n6247) );
  NAND2_X1 U8040 ( .A1(n9492), .A2(n6421), .ZN(n6246) );
  NAND2_X1 U8041 ( .A1(n6247), .A2(n6246), .ZN(n9289) );
  NAND2_X1 U8042 ( .A1(n9366), .A2(n9289), .ZN(n6248) );
  INV_X1 U8043 ( .A(n9374), .ZN(n6254) );
  INV_X1 U8044 ( .A(n9371), .ZN(n9370) );
  INV_X1 U8045 ( .A(n6249), .ZN(n9473) );
  NAND2_X1 U8046 ( .A1(n9370), .A2(n9473), .ZN(n6250) );
  NAND2_X1 U8047 ( .A1(n6250), .A2(n9373), .ZN(n6253) );
  INV_X1 U8048 ( .A(n6250), .ZN(n6252) );
  INV_X1 U8049 ( .A(n9373), .ZN(n6251) );
  AOI22_X1 U8050 ( .A1(n6254), .A2(n6253), .B1(n6252), .B2(n6251), .ZN(n6258)
         );
  INV_X1 U8051 ( .A(n6255), .ZN(n6256) );
  OR3_X1 U8052 ( .A1(n6256), .A2(n9289), .A3(n9366), .ZN(n6257) );
  AND2_X1 U8053 ( .A1(n6258), .A2(n6257), .ZN(n6259) );
  NAND2_X1 U8054 ( .A1(n7122), .A2(n6555), .ZN(n6263) );
  NAND2_X1 U8055 ( .A1(n6260), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6261) );
  XNOR2_X1 U8056 ( .A(n6261), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9938) );
  AOI22_X1 U8057 ( .A1(n6556), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n6295), .B2(
        n9938), .ZN(n6262) );
  NAND2_X1 U8058 ( .A1(n6265), .A2(n6264), .ZN(n6266) );
  AND2_X1 U8059 ( .A1(n6299), .A2(n6266), .ZN(n9775) );
  NAND2_X1 U8060 ( .A1(n9775), .A2(n7243), .ZN(n6269) );
  AOI22_X1 U8061 ( .A1(n6060), .A2(P1_REG0_REG_17__SCAN_IN), .B1(n6486), .B2(
        P1_REG1_REG_17__SCAN_IN), .ZN(n6268) );
  INV_X1 U8062 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n9765) );
  OR2_X1 U8063 ( .A1(n6563), .A2(n9765), .ZN(n6267) );
  OAI22_X1 U8064 ( .A1(n9767), .A2(n9334), .B1(n9453), .B2(n6389), .ZN(n6270)
         );
  XNOR2_X1 U8065 ( .A(n6270), .B(n9335), .ZN(n9384) );
  OR2_X1 U8066 ( .A1(n9767), .A2(n6389), .ZN(n6272) );
  OR2_X1 U8067 ( .A1(n9453), .A2(n4423), .ZN(n6271) );
  AND2_X1 U8068 ( .A1(n9384), .A2(n9383), .ZN(n6273) );
  INV_X1 U8069 ( .A(n9384), .ZN(n6275) );
  INV_X1 U8070 ( .A(n9383), .ZN(n6274) );
  NAND2_X1 U8071 ( .A1(n6275), .A2(n6274), .ZN(n6276) );
  NAND2_X1 U8072 ( .A1(n6277), .A2(n6276), .ZN(n9318) );
  NAND2_X1 U8073 ( .A1(n7191), .A2(n6555), .ZN(n6282) );
  OR2_X1 U8074 ( .A1(n5894), .A2(n6278), .ZN(n6279) );
  AND2_X1 U8075 ( .A1(n6280), .A2(n6279), .ZN(n9958) );
  AOI22_X1 U8076 ( .A1(n6556), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n9958), .B2(
        n6295), .ZN(n6281) );
  NAND2_X1 U8077 ( .A1(n7834), .A2(n6398), .ZN(n6289) );
  XNOR2_X1 U8078 ( .A(n6299), .B(P1_REG3_REG_18__SCAN_IN), .ZN(n9745) );
  NAND2_X1 U8079 ( .A1(n9745), .A2(n7243), .ZN(n6287) );
  INV_X1 U8080 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n9129) );
  NAND2_X1 U8081 ( .A1(n6323), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n6284) );
  NAND2_X1 U8082 ( .A1(n7878), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n6283) );
  OAI211_X1 U8083 ( .C1(n9129), .C2(n7881), .A(n6284), .B(n6283), .ZN(n6285)
         );
  INV_X1 U8084 ( .A(n6285), .ZN(n6286) );
  NAND2_X1 U8085 ( .A1(n6287), .A2(n6286), .ZN(n9772) );
  NAND2_X1 U8086 ( .A1(n9772), .A2(n4391), .ZN(n6288) );
  NAND2_X1 U8087 ( .A1(n6289), .A2(n6288), .ZN(n6290) );
  XNOR2_X1 U8088 ( .A(n6290), .B(n9335), .ZN(n9319) );
  NAND2_X1 U8089 ( .A1(n7834), .A2(n4391), .ZN(n6292) );
  NAND2_X1 U8090 ( .A1(n9772), .A2(n6421), .ZN(n6291) );
  AND2_X1 U8091 ( .A1(n6292), .A2(n6291), .ZN(n6309) );
  NAND2_X1 U8092 ( .A1(n9319), .A2(n6309), .ZN(n6293) );
  NAND2_X1 U8093 ( .A1(n9318), .A2(n6293), .ZN(n6317) );
  AOI22_X1 U8094 ( .A1(n6602), .A2(n6295), .B1(n6556), .B2(
        P2_DATAO_REG_19__SCAN_IN), .ZN(n6296) );
  INV_X1 U8095 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n6298) );
  INV_X1 U8096 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n6297) );
  OAI21_X1 U8097 ( .B1(n6299), .B2(n6298), .A(n6297), .ZN(n6300) );
  NAND2_X1 U8098 ( .A1(n6321), .A2(n6300), .ZN(n9732) );
  OR2_X1 U8099 ( .A1(n9732), .A2(n6442), .ZN(n6305) );
  INV_X1 U8100 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n9733) );
  NAND2_X1 U8101 ( .A1(n6060), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n6302) );
  NAND2_X1 U8102 ( .A1(n6486), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n6301) );
  OAI211_X1 U8103 ( .C1(n9733), .C2(n6563), .A(n6302), .B(n6301), .ZN(n6303)
         );
  INV_X1 U8104 ( .A(n6303), .ZN(n6304) );
  OAI22_X1 U8105 ( .A1(n9731), .A2(n9334), .B1(n9717), .B2(n6389), .ZN(n6306)
         );
  XNOR2_X1 U8106 ( .A(n6306), .B(n6426), .ZN(n6312) );
  OR2_X1 U8107 ( .A1(n9731), .A2(n6389), .ZN(n6308) );
  NAND2_X1 U8108 ( .A1(n9754), .A2(n6421), .ZN(n6307) );
  NAND2_X1 U8109 ( .A1(n6308), .A2(n6307), .ZN(n6313) );
  NAND2_X1 U8110 ( .A1(n6312), .A2(n6313), .ZN(n9323) );
  INV_X1 U8111 ( .A(n9319), .ZN(n6310) );
  INV_X1 U8112 ( .A(n6309), .ZN(n9450) );
  NAND2_X1 U8113 ( .A1(n6310), .A2(n9450), .ZN(n6311) );
  AND2_X1 U8114 ( .A1(n9323), .A2(n6311), .ZN(n6316) );
  INV_X1 U8115 ( .A(n6312), .ZN(n6315) );
  INV_X1 U8116 ( .A(n6313), .ZN(n6314) );
  AND2_X1 U8117 ( .A1(n6315), .A2(n6314), .ZN(n9324) );
  NAND2_X1 U8118 ( .A1(n7334), .A2(n6555), .ZN(n6319) );
  NAND2_X1 U8119 ( .A1(n5988), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n6318) );
  NAND2_X1 U8120 ( .A1(n9829), .A2(n6398), .ZN(n6330) );
  NAND2_X1 U8121 ( .A1(n6321), .A2(n6320), .ZN(n6322) );
  AND2_X1 U8122 ( .A1(n6341), .A2(n6322), .ZN(n9721) );
  NAND2_X1 U8123 ( .A1(n9721), .A2(n7243), .ZN(n6328) );
  INV_X1 U8124 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n9095) );
  NAND2_X1 U8125 ( .A1(n7878), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n6325) );
  NAND2_X1 U8126 ( .A1(n6486), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n6324) );
  OAI211_X1 U8127 ( .C1(n7881), .C2(n9095), .A(n6325), .B(n6324), .ZN(n6326)
         );
  INV_X1 U8128 ( .A(n6326), .ZN(n6327) );
  NAND2_X1 U8129 ( .A1(n6328), .A2(n6327), .ZN(n9490) );
  NAND2_X1 U8130 ( .A1(n9490), .A2(n4391), .ZN(n6329) );
  NAND2_X1 U8131 ( .A1(n6330), .A2(n6329), .ZN(n6331) );
  XNOR2_X1 U8132 ( .A(n6331), .B(n9335), .ZN(n9414) );
  AND2_X1 U8133 ( .A1(n9490), .A2(n6421), .ZN(n6332) );
  AOI21_X1 U8134 ( .B1(n9829), .B2(n4391), .A(n6332), .ZN(n6334) );
  NAND2_X1 U8135 ( .A1(n9414), .A2(n6334), .ZN(n6333) );
  NAND2_X1 U8136 ( .A1(n9416), .A2(n6333), .ZN(n6337) );
  INV_X1 U8137 ( .A(n9414), .ZN(n6335) );
  INV_X1 U8138 ( .A(n6334), .ZN(n9413) );
  NAND2_X1 U8139 ( .A1(n6335), .A2(n9413), .ZN(n6336) );
  NAND2_X1 U8140 ( .A1(n7517), .A2(n6555), .ZN(n6339) );
  NAND2_X1 U8141 ( .A1(n5988), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n6338) );
  NAND2_X1 U8142 ( .A1(n9824), .A2(n5931), .ZN(n6350) );
  INV_X1 U8143 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n6340) );
  NAND2_X1 U8144 ( .A1(n6341), .A2(n6340), .ZN(n6342) );
  NAND2_X1 U8145 ( .A1(n6343), .A2(n6342), .ZN(n9701) );
  OR2_X1 U8146 ( .A1(n9701), .A2(n6442), .ZN(n6348) );
  INV_X1 U8147 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n9702) );
  NAND2_X1 U8148 ( .A1(n6060), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n6345) );
  INV_X1 U8149 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n9097) );
  OR2_X1 U8150 ( .A1(n7247), .A2(n9097), .ZN(n6344) );
  OAI211_X1 U8151 ( .C1(n9702), .C2(n6563), .A(n6345), .B(n6344), .ZN(n6346)
         );
  INV_X1 U8152 ( .A(n6346), .ZN(n6347) );
  NAND2_X1 U8153 ( .A1(n6348), .A2(n6347), .ZN(n9686) );
  NAND2_X1 U8154 ( .A1(n9686), .A2(n4391), .ZN(n6349) );
  NAND2_X1 U8155 ( .A1(n6350), .A2(n6349), .ZN(n6351) );
  XNOR2_X1 U8156 ( .A(n6351), .B(n9335), .ZN(n6354) );
  AND2_X1 U8157 ( .A1(n9686), .A2(n6421), .ZN(n6352) );
  AOI21_X1 U8158 ( .B1(n9824), .B2(n6423), .A(n6352), .ZN(n6353) );
  XNOR2_X1 U8159 ( .A(n6354), .B(n6353), .ZN(n9354) );
  NAND2_X1 U8160 ( .A1(n6354), .A2(n6353), .ZN(n6355) );
  NAND2_X1 U8161 ( .A1(n7610), .A2(n6555), .ZN(n6357) );
  NAND2_X1 U8162 ( .A1(n5988), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n6356) );
  NAND2_X1 U8163 ( .A1(n9814), .A2(n6398), .ZN(n6368) );
  INV_X1 U8164 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n6358) );
  NAND2_X1 U8165 ( .A1(n6359), .A2(n6358), .ZN(n6360) );
  AND2_X1 U8166 ( .A1(n6380), .A2(n6360), .ZN(n9676) );
  NAND2_X1 U8167 ( .A1(n9676), .A2(n7243), .ZN(n6366) );
  INV_X1 U8168 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n6363) );
  NAND2_X1 U8169 ( .A1(n6060), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n6362) );
  NAND2_X1 U8170 ( .A1(n6486), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n6361) );
  OAI211_X1 U8171 ( .C1(n6363), .C2(n6563), .A(n6362), .B(n6361), .ZN(n6364)
         );
  INV_X1 U8172 ( .A(n6364), .ZN(n6365) );
  NAND2_X1 U8173 ( .A1(n6366), .A2(n6365), .ZN(n9687) );
  NAND2_X1 U8174 ( .A1(n9687), .A2(n4391), .ZN(n6367) );
  NAND2_X1 U8175 ( .A1(n6368), .A2(n6367), .ZN(n6369) );
  XNOR2_X1 U8176 ( .A(n6369), .B(n6426), .ZN(n6373) );
  NAND2_X1 U8177 ( .A1(n9814), .A2(n4391), .ZN(n6371) );
  NAND2_X1 U8178 ( .A1(n9687), .A2(n6421), .ZN(n6370) );
  NAND2_X1 U8179 ( .A1(n6371), .A2(n6370), .ZN(n6374) );
  NAND2_X1 U8180 ( .A1(n6373), .A2(n6374), .ZN(n7757) );
  INV_X1 U8181 ( .A(n7756), .ZN(n7754) );
  INV_X1 U8182 ( .A(n7769), .ZN(n6372) );
  NOR2_X1 U8183 ( .A1(n7754), .A2(n6372), .ZN(n6377) );
  INV_X1 U8184 ( .A(n6373), .ZN(n6376) );
  INV_X1 U8185 ( .A(n6374), .ZN(n6375) );
  AOI21_X1 U8186 ( .B1(n6377), .B2(n7757), .A(n7760), .ZN(n6394) );
  NAND2_X1 U8187 ( .A1(n5988), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n6378) );
  INV_X1 U8188 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n6379) );
  NAND2_X1 U8189 ( .A1(n6380), .A2(n6379), .ZN(n6381) );
  NAND2_X1 U8190 ( .A1(n6401), .A2(n6381), .ZN(n7763) );
  OR2_X1 U8191 ( .A1(n7763), .A2(n6442), .ZN(n6387) );
  INV_X1 U8192 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n6384) );
  NAND2_X1 U8193 ( .A1(n6060), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n6383) );
  NAND2_X1 U8194 ( .A1(n6486), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n6382) );
  OAI211_X1 U8195 ( .C1(n6384), .C2(n6563), .A(n6383), .B(n6382), .ZN(n6385)
         );
  INV_X1 U8196 ( .A(n6385), .ZN(n6386) );
  OAI22_X1 U8197 ( .A1(n9664), .A2(n9334), .B1(n9673), .B2(n6389), .ZN(n6388)
         );
  XNOR2_X1 U8198 ( .A(n6388), .B(n9335), .ZN(n6393) );
  OR2_X1 U8199 ( .A1(n9664), .A2(n6389), .ZN(n6391) );
  NAND2_X1 U8200 ( .A1(n9641), .A2(n6421), .ZN(n6390) );
  NAND2_X1 U8201 ( .A1(n6393), .A2(n6392), .ZN(n6395) );
  OAI21_X1 U8202 ( .B1(n6393), .B2(n6392), .A(n6395), .ZN(n7759) );
  NAND2_X1 U8203 ( .A1(n7708), .A2(n6555), .ZN(n6397) );
  NAND2_X1 U8204 ( .A1(n5988), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n6396) );
  NAND2_X1 U8205 ( .A1(n9804), .A2(n5931), .ZN(n6409) );
  INV_X1 U8206 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n6400) );
  NAND2_X1 U8207 ( .A1(n6401), .A2(n6400), .ZN(n6402) );
  NAND2_X1 U8208 ( .A1(n6414), .A2(n6402), .ZN(n9646) );
  INV_X1 U8209 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n9071) );
  NAND2_X1 U8210 ( .A1(n6486), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n6404) );
  NAND2_X1 U8211 ( .A1(n7878), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n6403) );
  OAI211_X1 U8212 ( .C1(n7881), .C2(n9071), .A(n6404), .B(n6403), .ZN(n6405)
         );
  INV_X1 U8213 ( .A(n6405), .ZN(n6406) );
  NAND2_X1 U8214 ( .A1(n9657), .A2(n4391), .ZN(n6408) );
  NAND2_X1 U8215 ( .A1(n6409), .A2(n6408), .ZN(n6410) );
  XNOR2_X1 U8216 ( .A(n6410), .B(n6426), .ZN(n6429) );
  OAI22_X1 U8217 ( .A1(n9650), .A2(n6389), .B1(n9630), .B2(n4423), .ZN(n6428)
         );
  XNOR2_X1 U8218 ( .A(n6429), .B(n6428), .ZN(n9360) );
  NAND2_X1 U8219 ( .A1(n7727), .A2(n6555), .ZN(n6412) );
  NAND2_X1 U8220 ( .A1(n5988), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n6411) );
  INV_X1 U8221 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n6413) );
  NAND2_X1 U8222 ( .A1(n6414), .A2(n6413), .ZN(n6415) );
  NAND2_X1 U8223 ( .A1(n9632), .A2(n7243), .ZN(n6420) );
  INV_X1 U8224 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n9625) );
  NAND2_X1 U8225 ( .A1(n6486), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n6417) );
  NAND2_X1 U8226 ( .A1(n6060), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n6416) );
  OAI211_X1 U8227 ( .C1(n9625), .C2(n6563), .A(n6417), .B(n6416), .ZN(n6418)
         );
  INV_X1 U8228 ( .A(n6418), .ZN(n6419) );
  AND2_X1 U8229 ( .A1(n9642), .A2(n6421), .ZN(n6422) );
  AOI21_X1 U8230 ( .B1(n9800), .B2(n4391), .A(n6422), .ZN(n6433) );
  NAND2_X1 U8231 ( .A1(n9800), .A2(n5931), .ZN(n6425) );
  NAND2_X1 U8232 ( .A1(n9642), .A2(n4391), .ZN(n6424) );
  NAND2_X1 U8233 ( .A1(n6425), .A2(n6424), .ZN(n6427) );
  XNOR2_X1 U8234 ( .A(n6427), .B(n6426), .ZN(n6435) );
  XOR2_X1 U8235 ( .A(n6433), .B(n6435), .Z(n9461) );
  INV_X1 U8236 ( .A(n9461), .ZN(n6431) );
  NOR2_X1 U8237 ( .A1(n6429), .A2(n6428), .ZN(n9462) );
  INV_X1 U8238 ( .A(n6433), .ZN(n6434) );
  NAND2_X1 U8239 ( .A1(n9282), .A2(n6555), .ZN(n6437) );
  NAND2_X1 U8240 ( .A1(n6556), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n6436) );
  NAND2_X1 U8241 ( .A1(n9796), .A2(n5931), .ZN(n6449) );
  INV_X1 U8242 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n6439) );
  NAND2_X1 U8243 ( .A1(n6440), .A2(n6439), .ZN(n6441) );
  NAND2_X1 U8244 ( .A1(n8081), .A2(n6441), .ZN(n9615) );
  INV_X1 U8245 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n9114) );
  NAND2_X1 U8246 ( .A1(n6060), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n6444) );
  NAND2_X1 U8247 ( .A1(n7878), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n6443) );
  OAI211_X1 U8248 ( .C1(n7247), .C2(n9114), .A(n6444), .B(n6443), .ZN(n6445)
         );
  INV_X1 U8249 ( .A(n6445), .ZN(n6446) );
  NAND2_X1 U8250 ( .A1(n9590), .A2(n4391), .ZN(n6448) );
  NAND2_X1 U8251 ( .A1(n6449), .A2(n6448), .ZN(n6450) );
  XNOR2_X1 U8252 ( .A(n6450), .B(n9335), .ZN(n6453) );
  NOR2_X1 U8253 ( .A1(n9631), .A2(n4423), .ZN(n6451) );
  AOI21_X1 U8254 ( .B1(n9796), .B2(n6423), .A(n6451), .ZN(n6452) );
  NAND2_X1 U8255 ( .A1(n6453), .A2(n6452), .ZN(n9345) );
  OAI21_X1 U8256 ( .B1(n6453), .B2(n6452), .A(n9345), .ZN(n6455) );
  INV_X1 U8257 ( .A(n6454), .ZN(n6479) );
  NAND2_X1 U8258 ( .A1(n6457), .A2(P1_B_REG_SCAN_IN), .ZN(n6458) );
  MUX2_X1 U8259 ( .A(P1_B_REG_SCAN_IN), .B(n6458), .S(n7683), .Z(n6459) );
  INV_X1 U8260 ( .A(n6462), .ZN(n7728) );
  INV_X1 U8261 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n6460) );
  NAND2_X1 U8262 ( .A1(n6817), .A2(n6460), .ZN(n6461) );
  NAND2_X1 U8263 ( .A1(n6457), .A2(n6462), .ZN(n9879) );
  NAND2_X1 U8264 ( .A1(n6461), .A2(n9879), .ZN(n7364) );
  INV_X1 U8265 ( .A(n7364), .ZN(n6474) );
  INV_X1 U8266 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n6463) );
  AND2_X1 U8267 ( .A1(n6462), .A2(n7683), .ZN(n6821) );
  NOR4_X1 U8268 ( .A1(P1_D_REG_4__SCAN_IN), .A2(P1_D_REG_5__SCAN_IN), .A3(
        P1_D_REG_6__SCAN_IN), .A4(P1_D_REG_7__SCAN_IN), .ZN(n6472) );
  NOR4_X1 U8269 ( .A1(P1_D_REG_8__SCAN_IN), .A2(P1_D_REG_9__SCAN_IN), .A3(
        P1_D_REG_10__SCAN_IN), .A4(P1_D_REG_11__SCAN_IN), .ZN(n6471) );
  OR4_X1 U8270 ( .A1(P1_D_REG_28__SCAN_IN), .A2(P1_D_REG_2__SCAN_IN), .A3(
        P1_D_REG_13__SCAN_IN), .A4(P1_D_REG_3__SCAN_IN), .ZN(n6469) );
  NOR4_X1 U8271 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_18__SCAN_IN), .A3(
        P1_D_REG_19__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n6467) );
  NOR4_X1 U8272 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_12__SCAN_IN), .A3(
        P1_D_REG_14__SCAN_IN), .A4(P1_D_REG_16__SCAN_IN), .ZN(n6466) );
  NOR4_X1 U8273 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_27__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n6465) );
  NOR4_X1 U8274 ( .A1(P1_D_REG_21__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_23__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n6464) );
  NAND4_X1 U8275 ( .A1(n6467), .A2(n6466), .A3(n6465), .A4(n6464), .ZN(n6468)
         );
  NOR4_X1 U8276 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        n6469), .A4(n6468), .ZN(n6470) );
  NAND3_X1 U8277 ( .A1(n6472), .A2(n6471), .A3(n6470), .ZN(n6473) );
  NAND2_X1 U8278 ( .A1(n6817), .A2(n6473), .ZN(n6567) );
  NAND3_X1 U8279 ( .A1(n6474), .A2(n7365), .A3(n6567), .ZN(n6494) );
  NAND2_X1 U8280 ( .A1(n6475), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6476) );
  XNOR2_X1 U8281 ( .A(n6476), .B(n5856), .ZN(n6572) );
  INV_X1 U8282 ( .A(n6818), .ZN(n6492) );
  NAND2_X1 U8283 ( .A1(n10139), .A2(n8015), .ZN(n6493) );
  INV_X1 U8284 ( .A(n6502), .ZN(n6481) );
  NOR2_X1 U8285 ( .A1(n10062), .A2(n6480), .ZN(n10041) );
  NAND2_X1 U8286 ( .A1(n6481), .A2(n10041), .ZN(n6483) );
  INV_X1 U8287 ( .A(n6828), .ZN(n9891) );
  NAND2_X1 U8288 ( .A1(n10009), .A2(n6478), .ZN(n6485) );
  NOR2_X2 U8289 ( .A1(n6502), .A2(n6485), .ZN(n9451) );
  XNOR2_X1 U8290 ( .A(n8081), .B(P1_REG3_REG_28__SCAN_IN), .ZN(n9596) );
  NAND2_X1 U8291 ( .A1(n9596), .A2(n7243), .ZN(n6491) );
  INV_X1 U8292 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n9092) );
  NAND2_X1 U8293 ( .A1(n6486), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n6488) );
  NAND2_X1 U8294 ( .A1(n7878), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n6487) );
  OAI211_X1 U8295 ( .C1(n7881), .C2(n9092), .A(n6488), .B(n6487), .ZN(n6489)
         );
  INV_X1 U8296 ( .A(n6489), .ZN(n6490) );
  INV_X1 U8297 ( .A(n6478), .ZN(n6997) );
  OR2_X1 U8298 ( .A1(n8015), .A2(n6997), .ZN(n10063) );
  NOR2_X1 U8299 ( .A1(n10063), .A2(n6492), .ZN(n8027) );
  OR2_X1 U8300 ( .A1(n8027), .A2(n10041), .ZN(n6496) );
  INV_X1 U8301 ( .A(n6493), .ZN(n6495) );
  OAI21_X1 U8302 ( .B1(n6496), .B2(n6495), .A(n6494), .ZN(n6498) );
  AND2_X1 U8303 ( .A1(n6566), .A2(n6738), .ZN(n6497) );
  NAND2_X1 U8304 ( .A1(n6498), .A2(n6497), .ZN(n6980) );
  NAND2_X1 U8305 ( .A1(n6980), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6499) );
  OR2_X1 U8306 ( .A1(n6572), .A2(P1_U3086), .ZN(n8021) );
  INV_X1 U8307 ( .A(n8015), .ZN(n6500) );
  NAND2_X1 U8308 ( .A1(n10010), .A2(n6478), .ZN(n6501) );
  AOI22_X1 U8309 ( .A1(n9642), .A2(n9482), .B1(P1_REG3_REG_27__SCAN_IN), .B2(
        P1_U3086), .ZN(n6503) );
  OAI21_X1 U8310 ( .B1(n9479), .B2(n9615), .A(n6503), .ZN(n6504) );
  AOI21_X1 U8311 ( .B1(n9451), .B2(n9488), .A(n6504), .ZN(n6505) );
  OAI21_X1 U8312 ( .B1(n9619), .B2(n9485), .A(n6505), .ZN(n6506) );
  NAND2_X1 U8313 ( .A1(n6508), .A2(n6507), .ZN(P1_U3214) );
  AND2_X1 U8314 ( .A1(n6511), .A2(n6514), .ZN(n6512) );
  NAND2_X1 U8315 ( .A1(n6513), .A2(n6512), .ZN(n6518) );
  INV_X1 U8316 ( .A(n6514), .ZN(n6516) );
  INV_X1 U8317 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n6638) );
  INV_X1 U8318 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n6520) );
  MUX2_X1 U8319 ( .A(n6638), .B(n6520), .S(n6779), .Z(n6527) );
  XNOR2_X1 U8320 ( .A(n6527), .B(SI_28_), .ZN(n6524) );
  NAND2_X1 U8321 ( .A1(n9278), .A2(n6555), .ZN(n6522) );
  NAND2_X1 U8322 ( .A1(n6556), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n6521) );
  NAND2_X1 U8323 ( .A1(n10038), .A2(n10092), .ZN(n10025) );
  NOR2_X2 U8324 ( .A1(n10025), .A2(n10018), .ZN(n10026) );
  NAND2_X1 U8325 ( .A1(n10026), .A2(n10104), .ZN(n10000) );
  NOR2_X4 U8327 ( .A1(n9985), .A2(n10122), .ZN(n9984) );
  INV_X1 U8328 ( .A(n9407), .ZN(n10131) );
  NOR2_X2 U8329 ( .A1(n7617), .A2(n9430), .ZN(n7651) );
  AND2_X2 U8330 ( .A1(n7651), .A2(n7685), .ZN(n7691) );
  INV_X1 U8331 ( .A(n9829), .ZN(n9724) );
  NOR2_X2 U8332 ( .A1(n9674), .A2(n9809), .ZN(n6523) );
  INV_X1 U8333 ( .A(n6523), .ZN(n9660) );
  INV_X1 U8334 ( .A(SI_28_), .ZN(n6526) );
  NAND2_X1 U8335 ( .A1(n6527), .A2(n6526), .ZN(n6535) );
  NAND2_X1 U8336 ( .A1(n6536), .A2(n6535), .ZN(n6530) );
  INV_X1 U8337 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n9276) );
  INV_X1 U8338 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n6528) );
  MUX2_X1 U8339 ( .A(n9276), .B(n6528), .S(n6779), .Z(n6537) );
  XNOR2_X1 U8340 ( .A(n6537), .B(SI_29_), .ZN(n6529) );
  NAND2_X1 U8341 ( .A1(n9275), .A2(n6555), .ZN(n6532) );
  NAND2_X1 U8342 ( .A1(n6556), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n6531) );
  INV_X1 U8343 ( .A(SI_29_), .ZN(n6533) );
  NAND2_X1 U8344 ( .A1(n6537), .A2(n6533), .ZN(n6534) );
  NAND3_X1 U8345 ( .A1(n6536), .A2(n6535), .A3(n6534), .ZN(n6540) );
  INV_X1 U8346 ( .A(n6537), .ZN(n6538) );
  NAND2_X1 U8347 ( .A1(n6538), .A2(SI_29_), .ZN(n6539) );
  INV_X1 U8348 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n6541) );
  INV_X1 U8349 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n9274) );
  MUX2_X1 U8350 ( .A(n6541), .B(n9274), .S(n6778), .Z(n6543) );
  INV_X1 U8351 ( .A(SI_30_), .ZN(n6542) );
  NAND2_X1 U8352 ( .A1(n6543), .A2(n6542), .ZN(n6548) );
  INV_X1 U8353 ( .A(n6543), .ZN(n6544) );
  NAND2_X1 U8354 ( .A1(n6544), .A2(SI_30_), .ZN(n6545) );
  NAND2_X1 U8355 ( .A1(n6548), .A2(n6545), .ZN(n6549) );
  NAND2_X1 U8356 ( .A1(n9272), .A2(n6555), .ZN(n6547) );
  NAND2_X1 U8357 ( .A1(n6556), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n6546) );
  INV_X1 U8358 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n6551) );
  INV_X1 U8359 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n8451) );
  MUX2_X1 U8360 ( .A(n6551), .B(n8451), .S(n6778), .Z(n6552) );
  XNOR2_X1 U8361 ( .A(n6552), .B(SI_31_), .ZN(n6553) );
  NAND2_X1 U8362 ( .A1(n9267), .A2(n6555), .ZN(n6558) );
  NAND2_X1 U8363 ( .A1(n6556), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n6557) );
  XNOR2_X1 U8364 ( .A(n9579), .B(n6611), .ZN(n6559) );
  NAND2_X1 U8365 ( .A1(n6559), .A2(n10027), .ZN(n9582) );
  INV_X1 U8366 ( .A(n6827), .ZN(n9895) );
  AOI21_X1 U8367 ( .B1(n9895), .B2(P1_B_REG_SCAN_IN), .A(n10048), .ZN(n8051)
         );
  INV_X1 U8368 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n9576) );
  NAND2_X1 U8369 ( .A1(n6486), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n6562) );
  INV_X1 U8370 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n6560) );
  OR2_X1 U8371 ( .A1(n7881), .A2(n6560), .ZN(n6561) );
  OAI211_X1 U8372 ( .C1(n6563), .C2(n9576), .A(n6562), .B(n6561), .ZN(n8010)
         );
  NAND2_X1 U8373 ( .A1(n8051), .A2(n8010), .ZN(n7777) );
  OAI21_X1 U8374 ( .B1(n10039), .B2(n6294), .A(n7364), .ZN(n6568) );
  NAND3_X1 U8375 ( .A1(n6567), .A2(n6566), .A3(n6818), .ZN(n7366) );
  INV_X1 U8376 ( .A(n7365), .ZN(n6569) );
  NAND2_X1 U8377 ( .A1(n10144), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n6570) );
  INV_X1 U8378 ( .A(n6572), .ZN(n6573) );
  OR2_X1 U8379 ( .A1(n8015), .A2(n6573), .ZN(n6575) );
  AND2_X1 U8380 ( .A1(n6575), .A2(n6574), .ZN(n6605) );
  INV_X1 U8381 ( .A(n8021), .ZN(n8014) );
  OR2_X1 U8382 ( .A1(n6818), .A2(n8014), .ZN(n6606) );
  NOR2_X1 U8383 ( .A1(n6828), .A2(n6827), .ZN(n8026) );
  NAND2_X1 U8384 ( .A1(n6832), .A2(n8026), .ZN(n9928) );
  XNOR2_X1 U8385 ( .A(n9938), .B(n9765), .ZN(n9940) );
  XNOR2_X1 U8386 ( .A(n6780), .B(P1_REG2_REG_1__SCAN_IN), .ZN(n9507) );
  AND2_X1 U8387 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n9514) );
  NAND2_X1 U8388 ( .A1(n9507), .A2(n9514), .ZN(n9506) );
  NAND2_X1 U8389 ( .A1(n9505), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6576) );
  NAND2_X1 U8390 ( .A1(n9506), .A2(n6576), .ZN(n9527) );
  NAND2_X1 U8391 ( .A1(n4431), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6577) );
  NAND2_X1 U8392 ( .A1(n9526), .A2(n6577), .ZN(n9540) );
  XNOR2_X1 U8393 ( .A(n9535), .B(n7496), .ZN(n9541) );
  NAND2_X1 U8394 ( .A1(n9535), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6578) );
  MUX2_X1 U8395 ( .A(n7589), .B(P1_REG2_REG_5__SCAN_IN), .S(n6908), .Z(n6906)
         );
  NOR2_X1 U8396 ( .A1(n6907), .A2(n6906), .ZN(n6905) );
  XNOR2_X1 U8397 ( .A(n6925), .B(P1_REG2_REG_6__SCAN_IN), .ZN(n6923) );
  MUX2_X1 U8398 ( .A(n6579), .B(P1_REG2_REG_7__SCAN_IN), .S(n6936), .Z(n6931)
         );
  AOI21_X1 U8399 ( .B1(P1_REG2_REG_7__SCAN_IN), .B2(n6936), .A(n6930), .ZN(
        n6944) );
  XNOR2_X1 U8400 ( .A(n6948), .B(P1_REG2_REG_8__SCAN_IN), .ZN(n6943) );
  XNOR2_X1 U8401 ( .A(n9572), .B(n7511), .ZN(n9563) );
  NAND2_X1 U8402 ( .A1(n9562), .A2(n9563), .ZN(n9561) );
  OAI21_X1 U8403 ( .B1(n9572), .B2(P1_REG2_REG_9__SCAN_IN), .A(n9561), .ZN(
        n6768) );
  XNOR2_X1 U8404 ( .A(n6770), .B(P1_REG2_REG_10__SCAN_IN), .ZN(n6769) );
  XNOR2_X1 U8405 ( .A(n6745), .B(P1_REG2_REG_11__SCAN_IN), .ZN(n6743) );
  XNOR2_X1 U8406 ( .A(n7305), .B(n7570), .ZN(n7300) );
  XNOR2_X1 U8407 ( .A(n6758), .B(P1_REG2_REG_13__SCAN_IN), .ZN(n6757) );
  XNOR2_X1 U8408 ( .A(n9908), .B(P1_REG2_REG_14__SCAN_IN), .ZN(n9901) );
  NOR2_X1 U8409 ( .A1(n6580), .A2(n7107), .ZN(n6581) );
  INV_X1 U8410 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n9913) );
  NAND2_X1 U8411 ( .A1(n7159), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n6582) );
  OAI21_X1 U8412 ( .B1(n7159), .B2(P1_REG2_REG_16__SCAN_IN), .A(n6582), .ZN(
        n9930) );
  OR2_X1 U8413 ( .A1(n9938), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n6583) );
  NAND2_X1 U8414 ( .A1(n9958), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n6584) );
  OAI21_X1 U8415 ( .B1(n9958), .B2(P1_REG2_REG_18__SCAN_IN), .A(n6584), .ZN(
        n9953) );
  NAND2_X1 U8416 ( .A1(n9958), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n6599) );
  OAI21_X1 U8417 ( .B1(n9958), .B2(P1_REG1_REG_18__SCAN_IN), .A(n6599), .ZN(
        n9960) );
  INV_X1 U8418 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n6586) );
  XNOR2_X1 U8419 ( .A(n9938), .B(n6586), .ZN(n9943) );
  XOR2_X1 U8420 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n7159), .Z(n9926) );
  INV_X1 U8421 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n10148) );
  XNOR2_X1 U8422 ( .A(n6780), .B(P1_REG1_REG_1__SCAN_IN), .ZN(n9510) );
  AND2_X1 U8423 ( .A1(P1_REG1_REG_0__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n9509) );
  NAND2_X1 U8424 ( .A1(n9510), .A2(n9509), .ZN(n9508) );
  NAND2_X1 U8425 ( .A1(n9505), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6587) );
  NAND2_X1 U8426 ( .A1(n9508), .A2(n6587), .ZN(n9524) );
  NAND2_X1 U8427 ( .A1(n9525), .A2(n9524), .ZN(n9523) );
  NAND2_X1 U8428 ( .A1(n4431), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6588) );
  NAND2_X1 U8429 ( .A1(n9523), .A2(n6588), .ZN(n9537) );
  INV_X1 U8430 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6589) );
  XNOR2_X1 U8431 ( .A(n9535), .B(n6589), .ZN(n9538) );
  NAND2_X1 U8432 ( .A1(n9535), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6590) );
  NAND2_X1 U8433 ( .A1(n9536), .A2(n6590), .ZN(n9555) );
  INV_X1 U8434 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n10151) );
  XNOR2_X1 U8435 ( .A(n6908), .B(P1_REG1_REG_5__SCAN_IN), .ZN(n6903) );
  XNOR2_X1 U8436 ( .A(n6925), .B(P1_REG1_REG_6__SCAN_IN), .ZN(n6920) );
  NOR2_X1 U8437 ( .A1(n6921), .A2(n6920), .ZN(n6919) );
  MUX2_X1 U8438 ( .A(n6591), .B(P1_REG1_REG_7__SCAN_IN), .S(n6936), .Z(n6934)
         );
  NOR2_X1 U8439 ( .A1(n6935), .A2(n6934), .ZN(n6933) );
  XNOR2_X1 U8440 ( .A(n6948), .B(P1_REG1_REG_8__SCAN_IN), .ZN(n6946) );
  MUX2_X1 U8441 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n6592), .S(n9572), .Z(n9566)
         );
  OAI21_X1 U8442 ( .B1(n9572), .B2(P1_REG1_REG_9__SCAN_IN), .A(n9565), .ZN(
        n6765) );
  INV_X1 U8443 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n6593) );
  MUX2_X1 U8444 ( .A(n6593), .B(P1_REG1_REG_10__SCAN_IN), .S(n6770), .Z(n6766)
         );
  XNOR2_X1 U8445 ( .A(n6745), .B(P1_REG1_REG_11__SCAN_IN), .ZN(n6740) );
  XNOR2_X1 U8446 ( .A(n7305), .B(n6594), .ZN(n7304) );
  OAI21_X1 U8447 ( .B1(n7305), .B2(P1_REG1_REG_12__SCAN_IN), .A(n7302), .ZN(
        n6753) );
  XNOR2_X1 U8448 ( .A(n6758), .B(P1_REG1_REG_13__SCAN_IN), .ZN(n6754) );
  XNOR2_X1 U8449 ( .A(n9908), .B(P1_REG1_REG_14__SCAN_IN), .ZN(n9904) );
  NOR2_X1 U8450 ( .A1(n6595), .A2(n7107), .ZN(n6596) );
  NOR2_X1 U8451 ( .A1(n9917), .A2(n9918), .ZN(n9916) );
  OR2_X1 U8452 ( .A1(n9938), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n6597) );
  NAND2_X1 U8453 ( .A1(n6598), .A2(n6597), .ZN(n9961) );
  NAND2_X1 U8454 ( .A1(n9963), .A2(n6599), .ZN(n6600) );
  NAND2_X1 U8455 ( .A1(n9964), .A2(n6604), .ZN(n6601) );
  NAND2_X1 U8456 ( .A1(n6832), .A2(n6828), .ZN(n9948) );
  INV_X1 U8457 ( .A(n6605), .ZN(n6607) );
  NAND2_X1 U8458 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9328) );
  INV_X1 U8459 ( .A(n8082), .ZN(n6613) );
  INV_X1 U8460 ( .A(n6611), .ZN(n6612) );
  OAI211_X1 U8461 ( .C1(n6613), .C2(n7945), .A(n6612), .B(n10027), .ZN(n7780)
         );
  INV_X1 U8462 ( .A(n6614), .ZN(n6615) );
  NAND2_X1 U8463 ( .A1(n10144), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n6616) );
  NAND2_X1 U8464 ( .A1(n6720), .A2(n6618), .ZN(n6619) );
  NAND3_X1 U8465 ( .A1(n7012), .A2(n7396), .A3(n6619), .ZN(n8894) );
  INV_X1 U8466 ( .A(n7099), .ZN(n8297) );
  NAND2_X1 U8467 ( .A1(n6620), .A2(n8297), .ZN(n7097) );
  NAND2_X1 U8468 ( .A1(n7097), .A2(n8298), .ZN(n7184) );
  NAND2_X1 U8469 ( .A1(n7184), .A2(n8486), .ZN(n7125) );
  NAND2_X1 U8470 ( .A1(n6621), .A2(n7132), .ZN(n7178) );
  INV_X1 U8471 ( .A(n10164), .ZN(n6965) );
  NAND2_X1 U8472 ( .A1(n6880), .A2(n6965), .ZN(n7126) );
  AND2_X1 U8473 ( .A1(n7178), .A2(n7126), .ZN(n8306) );
  INV_X1 U8474 ( .A(n7219), .ZN(n7181) );
  NAND2_X1 U8475 ( .A1(n8536), .A2(n7181), .ZN(n8316) );
  INV_X1 U8476 ( .A(n7132), .ZN(n7171) );
  NAND2_X1 U8477 ( .A1(n8537), .A2(n7171), .ZN(n8313) );
  NAND2_X1 U8478 ( .A1(n7136), .A2(n7219), .ZN(n8312) );
  NAND2_X1 U8479 ( .A1(n8535), .A2(n7199), .ZN(n8317) );
  NAND2_X1 U8480 ( .A1(n7292), .A2(n7257), .ZN(n8320) );
  NAND2_X1 U8481 ( .A1(n6623), .A2(n8320), .ZN(n7294) );
  INV_X1 U8482 ( .A(n7340), .ZN(n7295) );
  NOR2_X1 U8483 ( .A1(n8534), .A2(n7295), .ZN(n8321) );
  NAND2_X1 U8484 ( .A1(n8534), .A2(n7295), .ZN(n8315) );
  OAI21_X1 U8485 ( .B1(n7294), .B2(n8321), .A(n8315), .ZN(n7386) );
  NAND2_X1 U8486 ( .A1(n9260), .A2(n8889), .ZN(n8491) );
  AND2_X1 U8487 ( .A1(n8491), .A2(n8860), .ZN(n8331) );
  INV_X1 U8488 ( .A(n8997), .ZN(n8151) );
  NAND2_X1 U8489 ( .A1(n8891), .A2(n8151), .ZN(n8327) );
  INV_X1 U8490 ( .A(n8906), .ZN(n8533) );
  NAND2_X1 U8491 ( .A1(n8533), .A2(n7553), .ZN(n8902) );
  NAND2_X1 U8492 ( .A1(n8331), .A2(n8879), .ZN(n6628) );
  NAND2_X1 U8493 ( .A1(n8906), .A2(n7445), .ZN(n8334) );
  INV_X1 U8494 ( .A(n8334), .ZN(n6624) );
  NAND2_X1 U8495 ( .A1(n8222), .A2(n8997), .ZN(n8333) );
  INV_X1 U8496 ( .A(n8333), .ZN(n8878) );
  AOI21_X1 U8497 ( .B1(n6624), .B2(n8327), .A(n8878), .ZN(n6626) );
  NAND2_X1 U8498 ( .A1(n8898), .A2(n6625), .ZN(n8335) );
  AND2_X2 U8499 ( .A1(n8860), .A2(n8335), .ZN(n8881) );
  NAND2_X1 U8500 ( .A1(n6626), .A2(n8881), .ZN(n8856) );
  AND2_X1 U8501 ( .A1(n8875), .A2(n8345), .ZN(n8490) );
  AOI21_X1 U8502 ( .B1(n8331), .B2(n8856), .A(n8490), .ZN(n6627) );
  OAI21_X2 U8503 ( .B1(n6628), .B2(n7386), .A(n6627), .ZN(n7595) );
  INV_X1 U8504 ( .A(n8493), .ZN(n7597) );
  NAND2_X1 U8505 ( .A1(n8349), .A2(n8846), .ZN(n6629) );
  XNOR2_X1 U8506 ( .A(n6663), .B(n8355), .ZN(n8841) );
  NAND2_X1 U8507 ( .A1(n8169), .A2(n8829), .ZN(n8356) );
  INV_X1 U8508 ( .A(n9248), .ZN(n8241) );
  NAND2_X1 U8509 ( .A1(n9248), .A2(n8847), .ZN(n6631) );
  XNOR2_X1 U8510 ( .A(n9241), .B(n8830), .ZN(n8823) );
  NOR2_X1 U8511 ( .A1(n9241), .A2(n6667), .ZN(n8362) );
  AOI21_X2 U8512 ( .B1(n8824), .B2(n8823), .A(n8362), .ZN(n8808) );
  INV_X1 U8513 ( .A(n9235), .ZN(n8292) );
  NAND2_X1 U8514 ( .A1(n8292), .A2(n8818), .ZN(n8369) );
  NOR2_X1 U8515 ( .A1(n8292), .A2(n8818), .ZN(n8367) );
  NAND2_X1 U8516 ( .A1(n9229), .A2(n8286), .ZN(n8374) );
  INV_X1 U8517 ( .A(n8371), .ZN(n8377) );
  NAND2_X1 U8518 ( .A1(n9223), .A2(n8778), .ZN(n8381) );
  INV_X1 U8519 ( .A(n8381), .ZN(n6634) );
  INV_X1 U8520 ( .A(n9220), .ZN(n6635) );
  NAND2_X1 U8521 ( .A1(n6635), .A2(n8768), .ZN(n8474) );
  NAND2_X1 U8522 ( .A1(n9213), .A2(n8779), .ZN(n8390) );
  INV_X1 U8523 ( .A(n8390), .ZN(n6636) );
  INV_X1 U8524 ( .A(n8398), .ZN(n8392) );
  NAND2_X1 U8525 ( .A1(n9207), .A2(n8769), .ZN(n8383) );
  OAI21_X2 U8526 ( .B1(n8753), .B2(n8392), .A(n8383), .ZN(n8740) );
  NAND2_X1 U8527 ( .A1(n8954), .A2(n8253), .ZN(n6672) );
  OAI21_X1 U8528 ( .B1(n8740), .B2(n8386), .A(n8400), .ZN(n8731) );
  NAND2_X1 U8529 ( .A1(n9197), .A2(n8747), .ZN(n8404) );
  NAND2_X1 U8530 ( .A1(n8259), .A2(n8724), .ZN(n8402) );
  INV_X1 U8531 ( .A(n8402), .ZN(n6637) );
  AOI21_X2 U8532 ( .B1(n8731), .B2(n8404), .A(n6637), .ZN(n8721) );
  NOR2_X1 U8533 ( .A1(n8471), .A2(n8403), .ZN(n8428) );
  NAND2_X1 U8534 ( .A1(n9178), .A2(n8711), .ZN(n8420) );
  INV_X1 U8535 ( .A(n8420), .ZN(n8410) );
  INV_X2 U8536 ( .A(n6689), .ZN(n9165) );
  NAND2_X1 U8537 ( .A1(n9278), .A2(n8450), .ZN(n6640) );
  OR2_X1 U8538 ( .A1(n8435), .A2(n6638), .ZN(n6639) );
  NAND2_X1 U8539 ( .A1(n9159), .A2(n8470), .ZN(n6641) );
  INV_X1 U8540 ( .A(n9159), .ZN(n6697) );
  NAND2_X1 U8541 ( .A1(n9275), .A2(n8450), .ZN(n6643) );
  OR2_X1 U8542 ( .A1(n8452), .A2(n9276), .ZN(n6642) );
  INV_X1 U8543 ( .A(n8088), .ZN(n6645) );
  NAND2_X1 U8544 ( .A1(n6645), .A2(n6644), .ZN(n8462) );
  INV_X1 U8545 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n6648) );
  NAND2_X1 U8546 ( .A1(n5349), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n6647) );
  NAND2_X1 U8547 ( .A1(n8457), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n6646) );
  OAI211_X1 U8548 ( .C1(n5429), .C2(n6648), .A(n6647), .B(n6646), .ZN(n6649)
         );
  INV_X1 U8549 ( .A(n6649), .ZN(n6650) );
  NAND2_X1 U8550 ( .A1(n6726), .A2(n8531), .ZN(n8466) );
  INV_X1 U8551 ( .A(n6699), .ZN(n6651) );
  XNOR2_X1 U8552 ( .A(n8465), .B(n6651), .ZN(n8091) );
  NOR2_X1 U8553 ( .A1(n6914), .A2(n6969), .ZN(n7100) );
  OAI22_X1 U8554 ( .A1(n6620), .A2(n7100), .B1(n7226), .B2(n4967), .ZN(n7185)
         );
  AOI22_X1 U8555 ( .A1(n7185), .A2(n8302), .B1(n6880), .B2(n10164), .ZN(n7127)
         );
  INV_X1 U8556 ( .A(n6653), .ZN(n7290) );
  OAI21_X1 U8557 ( .B1(n6653), .B2(n8534), .A(n7340), .ZN(n6654) );
  NAND2_X1 U8558 ( .A1(n8333), .A2(n8327), .ZN(n8908) );
  NAND2_X1 U8559 ( .A1(n8906), .A2(n7553), .ZN(n8909) );
  NAND3_X1 U8560 ( .A1(n8479), .A2(n8908), .A3(n8909), .ZN(n6656) );
  AND2_X1 U8561 ( .A1(n8891), .A2(n8997), .ZN(n8884) );
  AOI21_X1 U8562 ( .B1(n8916), .B2(n8898), .A(n8884), .ZN(n6655) );
  AND2_X1 U8563 ( .A1(n6656), .A2(n6655), .ZN(n6658) );
  INV_X1 U8564 ( .A(n6658), .ZN(n8862) );
  NAND2_X1 U8565 ( .A1(n8908), .A2(n8909), .ZN(n8883) );
  NOR2_X1 U8566 ( .A1(n8898), .A2(n8916), .ZN(n8864) );
  NOR2_X1 U8567 ( .A1(n8875), .A2(n8889), .ZN(n6657) );
  AOI211_X1 U8568 ( .C1(n6658), .C2(n8883), .A(n8864), .B(n6657), .ZN(n6659)
         );
  OAI21_X1 U8569 ( .B1(n7384), .B2(n8862), .A(n6659), .ZN(n6661) );
  NAND2_X1 U8570 ( .A1(n6661), .A2(n6660), .ZN(n7598) );
  NAND2_X1 U8571 ( .A1(n6663), .A2(n8829), .ZN(n6664) );
  NAND2_X1 U8572 ( .A1(n8844), .A2(n6664), .ZN(n6666) );
  NAND2_X1 U8573 ( .A1(n9248), .A2(n8819), .ZN(n8476) );
  NOR2_X1 U8574 ( .A1(n9248), .A2(n8819), .ZN(n8477) );
  NAND2_X1 U8575 ( .A1(n9235), .A2(n8818), .ZN(n8364) );
  OR2_X1 U8576 ( .A1(n9235), .A2(n8818), .ZN(n8365) );
  INV_X1 U8577 ( .A(n9229), .ZN(n8187) );
  OAI22_X1 U8578 ( .A1(n8801), .A2(n8800), .B1(n8286), .B2(n8187), .ZN(n8791)
         );
  NAND2_X1 U8579 ( .A1(n8375), .A2(n8381), .ZN(n8789) );
  NAND2_X1 U8580 ( .A1(n9223), .A2(n8802), .ZN(n6668) );
  NOR2_X1 U8581 ( .A1(n9220), .A2(n8768), .ZN(n6671) );
  NAND2_X1 U8582 ( .A1(n9220), .A2(n8768), .ZN(n6670) );
  NAND2_X1 U8583 ( .A1(n8398), .A2(n8383), .ZN(n8755) );
  NAND2_X1 U8584 ( .A1(n9213), .A2(n8757), .ZN(n6674) );
  AND2_X1 U8585 ( .A1(n8755), .A2(n6674), .ZN(n8743) );
  NAND2_X1 U8586 ( .A1(n8391), .A2(n8390), .ZN(n8764) );
  INV_X1 U8587 ( .A(n6674), .ZN(n8754) );
  NOR2_X1 U8588 ( .A1(n8764), .A2(n8754), .ZN(n6675) );
  NAND2_X1 U8589 ( .A1(n8755), .A2(n6675), .ZN(n6677) );
  INV_X1 U8590 ( .A(n8769), .ZN(n8532) );
  OR2_X1 U8591 ( .A1(n9207), .A2(n8532), .ZN(n6676) );
  NAND2_X1 U8592 ( .A1(n6677), .A2(n6676), .ZN(n8742) );
  AOI22_X1 U8593 ( .A1(n8744), .A2(n8742), .B1(n8253), .B2(n6678), .ZN(n6679)
         );
  NAND2_X1 U8594 ( .A1(n8259), .A2(n8747), .ZN(n6680) );
  NOR2_X1 U8595 ( .A1(n9191), .A2(n8734), .ZN(n6683) );
  NAND2_X1 U8596 ( .A1(n9191), .A2(n8734), .ZN(n6682) );
  NOR2_X1 U8597 ( .A1(n8945), .A2(n8702), .ZN(n6685) );
  NAND2_X1 U8598 ( .A1(n8945), .A2(n8702), .ZN(n6684) );
  OR2_X1 U8599 ( .A1(n8705), .A2(n4986), .ZN(n8668) );
  NAND2_X1 U8600 ( .A1(n6689), .A2(n8274), .ZN(n6694) );
  INV_X1 U8601 ( .A(n6694), .ZN(n6687) );
  OR2_X1 U8602 ( .A1(n6689), .A2(n8274), .ZN(n6692) );
  NAND2_X1 U8603 ( .A1(n9178), .A2(n8687), .ZN(n8683) );
  NAND2_X1 U8604 ( .A1(n9171), .A2(n8699), .ZN(n6690) );
  AND2_X1 U8605 ( .A1(n8683), .A2(n6690), .ZN(n6691) );
  NAND2_X1 U8606 ( .A1(n6692), .A2(n8669), .ZN(n6693) );
  NOR2_X1 U8607 ( .A1(n9159), .A2(n8673), .ZN(n6698) );
  OAI22_X1 U8608 ( .A1(n8654), .A2(n6698), .B1(n6697), .B2(n8470), .ZN(n6700)
         );
  XNOR2_X1 U8609 ( .A(n6700), .B(n6699), .ZN(n6712) );
  NAND2_X1 U8610 ( .A1(n6701), .A2(n8525), .ZN(n6703) );
  NAND2_X1 U8611 ( .A1(n8295), .A2(n6702), .ZN(n8469) );
  INV_X1 U8612 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n9156) );
  NAND2_X1 U8613 ( .A1(n4272), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n6705) );
  NAND2_X1 U8614 ( .A1(n8457), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n6704) );
  OAI211_X1 U8615 ( .C1(n9156), .C2(n5429), .A(n6705), .B(n6704), .ZN(n6706)
         );
  INV_X1 U8616 ( .A(n6706), .ZN(n6707) );
  AND2_X1 U8617 ( .A1(n8462), .A2(n6707), .ZN(n8438) );
  INV_X1 U8618 ( .A(P2_B_REG_SCAN_IN), .ZN(n6709) );
  OAI21_X1 U8619 ( .B1(n6710), .B2(n6709), .A(n8917), .ZN(n8647) );
  OAI22_X1 U8620 ( .A1(n8470), .A2(n8905), .B1(n8438), .B2(n8647), .ZN(n6711)
         );
  INV_X1 U8621 ( .A(n6713), .ZN(n6714) );
  OAI21_X1 U8622 ( .B1(n8295), .B2(n7397), .A(n6714), .ZN(n6719) );
  INV_X1 U8623 ( .A(n6715), .ZN(n6796) );
  AND2_X1 U8624 ( .A1(n6796), .A2(n6716), .ZN(n6717) );
  NAND2_X1 U8625 ( .A1(n6718), .A2(n6717), .ZN(n7009) );
  NOR2_X1 U8626 ( .A1(n6719), .A2(n7009), .ZN(n6725) );
  OR2_X1 U8627 ( .A1(n6720), .A2(n8503), .ZN(n6721) );
  NAND2_X1 U8628 ( .A1(n6721), .A2(n8504), .ZN(n6722) );
  NAND2_X1 U8629 ( .A1(n6722), .A2(n7007), .ZN(n6723) );
  NAND2_X1 U8630 ( .A1(n6724), .A2(n6723), .ZN(n7011) );
  NAND2_X1 U8631 ( .A1(n6727), .A2(n4976), .ZN(P2_U3488) );
  NAND2_X1 U8632 ( .A1(n7012), .A2(n6728), .ZN(n6729) );
  NAND2_X1 U8633 ( .A1(n6730), .A2(n6729), .ZN(n6734) );
  NAND2_X1 U8634 ( .A1(n6732), .A2(n6731), .ZN(n6733) );
  NAND2_X1 U8635 ( .A1(n6736), .A2(n4974), .ZN(P2_U3456) );
  INV_X1 U8636 ( .A(n6737), .ZN(n6979) );
  AOI211_X1 U8637 ( .C1(n6741), .C2(n6740), .A(n9915), .B(n6739), .ZN(n6751)
         );
  AOI211_X1 U8638 ( .C1(n6744), .C2(n6743), .A(n9928), .B(n6742), .ZN(n6750)
         );
  INV_X1 U8639 ( .A(n6745), .ZN(n6836) );
  NOR2_X1 U8640 ( .A1(n9948), .A2(n6836), .ZN(n6749) );
  INV_X1 U8641 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n6747) );
  AND2_X1 U8642 ( .A1(P1_U3086), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n9439) );
  INV_X1 U8643 ( .A(n9439), .ZN(n6746) );
  OAI21_X1 U8644 ( .B1(n9970), .B2(n6747), .A(n6746), .ZN(n6748) );
  OR4_X1 U8645 ( .A1(n6751), .A2(n6750), .A3(n6749), .A4(n6748), .ZN(P1_U3254)
         );
  AOI211_X1 U8646 ( .C1(n6754), .C2(n6753), .A(n9915), .B(n6752), .ZN(n6763)
         );
  AOI211_X1 U8647 ( .C1(n6757), .C2(n6756), .A(n9928), .B(n6755), .ZN(n6762)
         );
  INV_X1 U8648 ( .A(n6758), .ZN(n6954) );
  NOR2_X1 U8649 ( .A1(n9948), .A2(n6954), .ZN(n6761) );
  INV_X1 U8650 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n6759) );
  NAND2_X1 U8651 ( .A1(P1_U3086), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n9424) );
  OAI21_X1 U8652 ( .B1(n9970), .B2(n6759), .A(n9424), .ZN(n6760) );
  OR4_X1 U8653 ( .A1(n6763), .A2(n6762), .A3(n6761), .A4(n6760), .ZN(P1_U3256)
         );
  AOI211_X1 U8654 ( .C1(n6766), .C2(n6765), .A(n9915), .B(n6764), .ZN(n6776)
         );
  AOI211_X1 U8655 ( .C1(n6769), .C2(n6768), .A(n9928), .B(n6767), .ZN(n6775)
         );
  INV_X1 U8656 ( .A(n6770), .ZN(n6824) );
  NOR2_X1 U8657 ( .A1(n9948), .A2(n6824), .ZN(n6774) );
  INV_X1 U8658 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n6772) );
  AND2_X1 U8659 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n9314) );
  INV_X1 U8660 ( .A(n9314), .ZN(n6771) );
  OAI21_X1 U8661 ( .B1(n9970), .B2(n6772), .A(n6771), .ZN(n6773) );
  OR4_X1 U8662 ( .A1(n6776), .A2(n6775), .A3(n6774), .A4(n6773), .ZN(P1_U3253)
         );
  NAND2_X1 U8663 ( .A1(n6778), .A2(P2_U3151), .ZN(n9286) );
  NOR2_X1 U8664 ( .A1(n6778), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9279) );
  INV_X2 U8665 ( .A(n9279), .ZN(n9283) );
  OAI222_X1 U8666 ( .A1(n9286), .A2(n4647), .B1(n9283), .B2(n5229), .C1(n6866), 
        .C2(P2_U3151), .ZN(P2_U3294) );
  OAI222_X1 U8667 ( .A1(n9286), .A2(n6782), .B1(P2_U3151), .B2(n7068), .C1(
        n5245), .C2(n9283), .ZN(P2_U3292) );
  NOR2_X2 U8668 ( .A1(n6779), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9894) );
  INV_X1 U8669 ( .A(n9894), .ZN(n7680) );
  OAI222_X1 U8670 ( .A1(n9897), .A2(n4647), .B1(n7680), .B2(n5228), .C1(
        P1_U3086), .C2(n6780), .ZN(P1_U3354) );
  AOI22_X1 U8671 ( .A1(n9894), .A2(P2_DATAO_REG_3__SCAN_IN), .B1(n9535), .B2(
        P1_STATE_REG_SCAN_IN), .ZN(n6781) );
  OAI21_X1 U8672 ( .B1(n6782), .B2(n9897), .A(n6781), .ZN(P1_U3352) );
  AOI22_X1 U8673 ( .A1(n9894), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(n4431), .B2(
        P1_STATE_REG_SCAN_IN), .ZN(n6783) );
  OAI21_X1 U8674 ( .B1(n6789), .B2(n9897), .A(n6783), .ZN(P1_U3353) );
  AOI22_X1 U8675 ( .A1(n6908), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n9894), .ZN(n6784) );
  OAI21_X1 U8676 ( .B1(n6786), .B2(n9897), .A(n6784), .ZN(P1_U3350) );
  OAI222_X1 U8677 ( .A1(n9286), .A2(n6786), .B1(P2_U3151), .B2(n6785), .C1(
        n5249), .C2(n9283), .ZN(P2_U3290) );
  AOI22_X1 U8678 ( .A1(n4422), .A2(P1_STATE_REG_SCAN_IN), .B1(n9894), .B2(
        P2_DATAO_REG_4__SCAN_IN), .ZN(n6787) );
  OAI21_X1 U8679 ( .B1(n5986), .B2(n9897), .A(n6787), .ZN(P1_U3351) );
  AOI22_X1 U8680 ( .A1(n6936), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n9894), .ZN(n6788) );
  OAI21_X1 U8681 ( .B1(n6792), .B2(n9897), .A(n6788), .ZN(P1_U3348) );
  INV_X1 U8682 ( .A(n9286), .ZN(n7609) );
  INV_X1 U8683 ( .A(n7609), .ZN(n9281) );
  OAI222_X1 U8684 ( .A1(n9283), .A2(n4496), .B1(n9281), .B2(n6789), .C1(n6851), 
        .C2(P2_U3151), .ZN(P2_U3293) );
  OAI222_X1 U8685 ( .A1(n9283), .A2(n6790), .B1(n9281), .B2(n5986), .C1(n7037), 
        .C2(P2_U3151), .ZN(P2_U3291) );
  OAI222_X1 U8686 ( .A1(n9286), .A2(n6792), .B1(P2_U3151), .B2(n6791), .C1(
        n4463), .C2(n9283), .ZN(P2_U3288) );
  INV_X1 U8687 ( .A(n6793), .ZN(n6805) );
  AOI22_X1 U8688 ( .A1(n6925), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n9894), .ZN(n6794) );
  OAI21_X1 U8689 ( .B1(n6805), .B2(n9897), .A(n6794), .ZN(P1_U3349) );
  INV_X1 U8690 ( .A(n6797), .ZN(n6798) );
  AOI22_X1 U8691 ( .A1(n6809), .A2(n6799), .B1(n6802), .B2(n6798), .ZN(
        P2_U3377) );
  INV_X1 U8692 ( .A(n6800), .ZN(n6801) );
  AOI22_X1 U8693 ( .A1(n6809), .A2(n6803), .B1(n6802), .B2(n6801), .ZN(
        P2_U3376) );
  INV_X1 U8694 ( .A(n6804), .ZN(n6896) );
  OAI222_X1 U8695 ( .A1(n9283), .A2(n6806), .B1(n9281), .B2(n6805), .C1(n6896), 
        .C2(P2_U3151), .ZN(P2_U3289) );
  AND2_X1 U8696 ( .A1(n6809), .A2(P2_D_REG_23__SCAN_IN), .ZN(P2_U3242) );
  AND2_X1 U8697 ( .A1(n6809), .A2(P2_D_REG_12__SCAN_IN), .ZN(P2_U3253) );
  AND2_X1 U8698 ( .A1(n6809), .A2(P2_D_REG_24__SCAN_IN), .ZN(P2_U3241) );
  AND2_X1 U8699 ( .A1(n6809), .A2(P2_D_REG_15__SCAN_IN), .ZN(P2_U3250) );
  AND2_X1 U8700 ( .A1(n6809), .A2(P2_D_REG_30__SCAN_IN), .ZN(P2_U3235) );
  AND2_X1 U8701 ( .A1(n6809), .A2(P2_D_REG_29__SCAN_IN), .ZN(P2_U3236) );
  AND2_X1 U8702 ( .A1(n6809), .A2(P2_D_REG_7__SCAN_IN), .ZN(P2_U3258) );
  AND2_X1 U8703 ( .A1(n6809), .A2(P2_D_REG_6__SCAN_IN), .ZN(P2_U3259) );
  AND2_X1 U8704 ( .A1(n6809), .A2(P2_D_REG_26__SCAN_IN), .ZN(P2_U3239) );
  AND2_X1 U8705 ( .A1(n6809), .A2(P2_D_REG_4__SCAN_IN), .ZN(P2_U3261) );
  AND2_X1 U8706 ( .A1(n6809), .A2(P2_D_REG_2__SCAN_IN), .ZN(P2_U3263) );
  AND2_X1 U8707 ( .A1(n6809), .A2(P2_D_REG_14__SCAN_IN), .ZN(P2_U3251) );
  AND2_X1 U8708 ( .A1(n6809), .A2(P2_D_REG_13__SCAN_IN), .ZN(P2_U3252) );
  AND2_X1 U8709 ( .A1(n6809), .A2(P2_D_REG_21__SCAN_IN), .ZN(P2_U3244) );
  AND2_X1 U8710 ( .A1(n6809), .A2(P2_D_REG_10__SCAN_IN), .ZN(P2_U3255) );
  AND2_X1 U8711 ( .A1(n6809), .A2(P2_D_REG_22__SCAN_IN), .ZN(P2_U3243) );
  AND2_X1 U8712 ( .A1(n6809), .A2(P2_D_REG_9__SCAN_IN), .ZN(P2_U3256) );
  AND2_X1 U8713 ( .A1(n6809), .A2(P2_D_REG_8__SCAN_IN), .ZN(P2_U3257) );
  AND2_X1 U8714 ( .A1(n6809), .A2(P2_D_REG_20__SCAN_IN), .ZN(P2_U3245) );
  AND2_X1 U8715 ( .A1(n6809), .A2(P2_D_REG_31__SCAN_IN), .ZN(P2_U3234) );
  AND2_X1 U8716 ( .A1(n6809), .A2(P2_D_REG_5__SCAN_IN), .ZN(P2_U3260) );
  AND2_X1 U8717 ( .A1(n6809), .A2(P2_D_REG_19__SCAN_IN), .ZN(P2_U3246) );
  AND2_X1 U8718 ( .A1(n6809), .A2(P2_D_REG_18__SCAN_IN), .ZN(P2_U3247) );
  AND2_X1 U8719 ( .A1(n6809), .A2(P2_D_REG_17__SCAN_IN), .ZN(P2_U3248) );
  AND2_X1 U8720 ( .A1(n6809), .A2(P2_D_REG_16__SCAN_IN), .ZN(P2_U3249) );
  AND2_X1 U8721 ( .A1(n6809), .A2(P2_D_REG_11__SCAN_IN), .ZN(P2_U3254) );
  INV_X1 U8722 ( .A(n6807), .ZN(n6811) );
  AOI22_X1 U8723 ( .A1(n6948), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n9894), .ZN(n6808) );
  OAI21_X1 U8724 ( .B1(n6811), .B2(n9897), .A(n6808), .ZN(P1_U3347) );
  INV_X1 U8725 ( .A(n6809), .ZN(n6810) );
  INV_X1 U8726 ( .A(P2_D_REG_28__SCAN_IN), .ZN(n9061) );
  NOR2_X1 U8727 ( .A1(n6810), .A2(n9061), .ZN(P2_U3237) );
  INV_X1 U8728 ( .A(P2_D_REG_27__SCAN_IN), .ZN(n9025) );
  NOR2_X1 U8729 ( .A1(n6810), .A2(n9025), .ZN(P2_U3238) );
  INV_X1 U8730 ( .A(P2_D_REG_25__SCAN_IN), .ZN(n9033) );
  NOR2_X1 U8731 ( .A1(n6810), .A2(n9033), .ZN(P2_U3240) );
  INV_X1 U8732 ( .A(P2_D_REG_3__SCAN_IN), .ZN(n9008) );
  NOR2_X1 U8733 ( .A1(n6810), .A2(n9008), .ZN(P2_U3262) );
  INV_X1 U8734 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6812) );
  OAI222_X1 U8735 ( .A1(n9283), .A2(n6812), .B1(n9281), .B2(n6811), .C1(n7086), 
        .C2(P2_U3151), .ZN(P2_U3287) );
  NAND2_X1 U8736 ( .A1(n7348), .A2(P1_U3973), .ZN(n6813) );
  OAI21_X1 U8737 ( .B1(P1_U3973), .B2(n5229), .A(n6813), .ZN(P1_U3555) );
  NAND2_X1 U8738 ( .A1(n8010), .A2(P1_U3973), .ZN(n6814) );
  OAI21_X1 U8739 ( .B1(P1_U3973), .B2(n8451), .A(n6814), .ZN(P1_U3585) );
  INV_X1 U8740 ( .A(n6815), .ZN(n6822) );
  AOI22_X1 U8741 ( .A1(n9572), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n9894), .ZN(n6816) );
  OAI21_X1 U8742 ( .B1(n6822), .B2(n9897), .A(n6816), .ZN(P1_U3346) );
  INV_X1 U8743 ( .A(n6817), .ZN(n6819) );
  NAND2_X1 U8744 ( .A1(n10074), .A2(P1_D_REG_0__SCAN_IN), .ZN(n6820) );
  OAI21_X1 U8745 ( .B1(n10074), .B2(n6821), .A(n6820), .ZN(P1_U3439) );
  OAI222_X1 U8746 ( .A1(n9286), .A2(n6822), .B1(P2_U3151), .B2(n4796), .C1(
        n9108), .C2(n9283), .ZN(P2_U3286) );
  INV_X1 U8747 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6823) );
  OAI222_X1 U8748 ( .A1(n9286), .A2(n6825), .B1(P2_U3151), .B2(n7272), .C1(
        n6823), .C2(n9283), .ZN(P2_U3285) );
  INV_X1 U8749 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n6826) );
  OAI222_X1 U8750 ( .A1(n7680), .A2(n6826), .B1(n9897), .B2(n6825), .C1(n6824), 
        .C2(P1_U3086), .ZN(P1_U3345) );
  INV_X1 U8751 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n6834) );
  NOR2_X1 U8752 ( .A1(n6827), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n6829) );
  NOR2_X1 U8753 ( .A1(n6829), .A2(n6828), .ZN(n9516) );
  OAI21_X1 U8754 ( .B1(n9895), .B2(P1_REG1_REG_0__SCAN_IN), .A(n9516), .ZN(
        n6830) );
  XNOR2_X1 U8755 ( .A(n6830), .B(P1_IR_REG_0__SCAN_IN), .ZN(n6831) );
  AOI22_X1 U8756 ( .A1(n6832), .A2(n6831), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        P1_U3086), .ZN(n6833) );
  OAI21_X1 U8757 ( .B1(n9970), .B2(n6834), .A(n6833), .ZN(P1_U3243) );
  INV_X1 U8758 ( .A(n9970), .ZN(n9546) );
  NOR2_X1 U8759 ( .A1(n9546), .A2(P1_U3973), .ZN(P1_U3085) );
  INV_X1 U8760 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6837) );
  INV_X1 U8761 ( .A(n6835), .ZN(n6838) );
  OAI222_X1 U8762 ( .A1(n7680), .A2(n6837), .B1(n9897), .B2(n6838), .C1(
        P1_U3086), .C2(n6836), .ZN(P1_U3344) );
  INV_X1 U8763 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6839) );
  OAI222_X1 U8764 ( .A1(n9283), .A2(n6839), .B1(n9281), .B2(n6838), .C1(n7477), 
        .C2(P2_U3151), .ZN(P2_U3284) );
  AOI22_X1 U8765 ( .A1(n7305), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n9894), .ZN(n6840) );
  OAI21_X1 U8766 ( .B1(n6842), .B2(n9897), .A(n6840), .ZN(P1_U3343) );
  INV_X1 U8767 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6841) );
  OAI222_X1 U8768 ( .A1(n9286), .A2(n6842), .B1(P2_U3151), .B2(n7521), .C1(
        n6841), .C2(n9283), .ZN(P2_U3283) );
  INV_X1 U8769 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n6848) );
  INV_X1 U8770 ( .A(n8615), .ZN(n8631) );
  AOI22_X1 U8771 ( .A1(n8631), .A2(P2_IR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3151), .ZN(n6847) );
  INV_X1 U8772 ( .A(n8626), .ZN(n7084) );
  OAI21_X1 U8773 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(n6843), .A(n6864), .ZN(n6844) );
  OAI21_X1 U8774 ( .B1(n6845), .B2(n7084), .A(n6844), .ZN(n6846) );
  OAI211_X1 U8775 ( .C1(n6848), .C2(n8634), .A(n6847), .B(n6846), .ZN(P2_U3182) );
  XNOR2_X1 U8776 ( .A(n6850), .B(n6849), .ZN(n6863) );
  INV_X1 U8777 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n10166) );
  OAI22_X1 U8778 ( .A1(n8615), .A2(n6851), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10166), .ZN(n6852) );
  AOI21_X1 U8779 ( .B1(n8611), .B2(P2_ADDR_REG_2__SCAN_IN), .A(n6852), .ZN(
        n6862) );
  INV_X1 U8780 ( .A(n8645), .ZN(n8541) );
  OAI21_X1 U8781 ( .B1(n6855), .B2(n6854), .A(n6853), .ZN(n6860) );
  OAI21_X1 U8782 ( .B1(n6858), .B2(n6857), .A(n6856), .ZN(n6859) );
  AOI22_X1 U8783 ( .A1(n8541), .A2(n6860), .B1(n8641), .B2(n6859), .ZN(n6861)
         );
  OAI211_X1 U8784 ( .C1(n8626), .C2(n6863), .A(n6862), .B(n6861), .ZN(P2_U3184) );
  XNOR2_X1 U8785 ( .A(n6865), .B(n6864), .ZN(n6875) );
  INV_X1 U8786 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n6884) );
  OAI22_X1 U8787 ( .A1(n8615), .A2(n6866), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6884), .ZN(n6867) );
  AOI21_X1 U8788 ( .B1(n8611), .B2(P2_ADDR_REG_1__SCAN_IN), .A(n6867), .ZN(
        n6874) );
  XNOR2_X1 U8789 ( .A(n6868), .B(P2_REG1_REG_1__SCAN_IN), .ZN(n6872) );
  OAI21_X1 U8790 ( .B1(P2_REG2_REG_1__SCAN_IN), .B2(n6870), .A(n6869), .ZN(
        n6871) );
  AOI22_X1 U8791 ( .A1(n8541), .A2(n6872), .B1(n8641), .B2(n6871), .ZN(n6873)
         );
  OAI211_X1 U8792 ( .C1(n8626), .C2(n6875), .A(n6874), .B(n6873), .ZN(P2_U3183) );
  NOR2_X1 U8793 ( .A1(n8288), .A2(P2_U3151), .ZN(n6968) );
  OAI21_X1 U8794 ( .B1(n6876), .B2(n6878), .A(n6877), .ZN(n6879) );
  NAND2_X1 U8795 ( .A1(n6879), .A2(n8216), .ZN(n6883) );
  OAI22_X1 U8796 ( .A1(n8266), .A2(n6914), .B1(n6880), .B2(n8285), .ZN(n6881)
         );
  AOI21_X1 U8797 ( .B1(n7226), .B2(n8276), .A(n6881), .ZN(n6882) );
  OAI211_X1 U8798 ( .C1(n6968), .C2(n6884), .A(n6883), .B(n6882), .ZN(P2_U3162) );
  AOI21_X1 U8799 ( .B1(n6886), .B2(n6885), .A(n7050), .ZN(n6901) );
  OAI21_X1 U8800 ( .B1(n6889), .B2(n6888), .A(n6887), .ZN(n6899) );
  INV_X1 U8801 ( .A(n6890), .ZN(n6892) );
  NAND3_X1 U8802 ( .A1(n6986), .A2(n6892), .A3(n6891), .ZN(n6893) );
  AOI21_X1 U8803 ( .B1(n6894), .B2(n6893), .A(n4586), .ZN(n6898) );
  NAND2_X1 U8804 ( .A1(P2_U3151), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n7265) );
  NAND2_X1 U8805 ( .A1(n8611), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n6895) );
  OAI211_X1 U8806 ( .C1(n8615), .C2(n6896), .A(n7265), .B(n6895), .ZN(n6897)
         );
  AOI211_X1 U8807 ( .C1(n6899), .C2(n8541), .A(n6898), .B(n6897), .ZN(n6900)
         );
  OAI21_X1 U8808 ( .B1(n6901), .B2(n8626), .A(n6900), .ZN(P2_U3188) );
  AOI211_X1 U8809 ( .C1(n6904), .C2(n6903), .A(n6902), .B(n9915), .ZN(n6913)
         );
  AOI211_X1 U8810 ( .C1(n6907), .C2(n6906), .A(n6905), .B(n9928), .ZN(n6912)
         );
  INV_X1 U8811 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n6910) );
  NAND2_X1 U8812 ( .A1(n9959), .A2(n6908), .ZN(n6909) );
  NAND2_X1 U8813 ( .A1(P1_U3086), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n7316) );
  OAI211_X1 U8814 ( .C1(n6910), .C2(n9970), .A(n6909), .B(n7316), .ZN(n6911)
         );
  OR3_X1 U8815 ( .A1(n6913), .A2(n6912), .A3(n6911), .ZN(P1_U3248) );
  AND2_X1 U8816 ( .A1(n7099), .A2(n8293), .ZN(n8480) );
  INV_X1 U8817 ( .A(n6968), .ZN(n6915) );
  NAND2_X1 U8818 ( .A1(n6915), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n6917) );
  AOI22_X1 U8819 ( .A1(n7019), .A2(n8276), .B1(n4967), .B2(n8264), .ZN(n6916)
         );
  OAI211_X1 U8820 ( .C1(n8480), .C2(n8279), .A(n6917), .B(n6916), .ZN(P2_U3172) );
  INV_X1 U8821 ( .A(n6180), .ZN(n6955) );
  INV_X1 U8822 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6918) );
  OAI222_X1 U8823 ( .A1(n9286), .A2(n6955), .B1(P2_U3151), .B2(n8544), .C1(
        n6918), .C2(n9283), .ZN(P2_U3282) );
  AOI211_X1 U8824 ( .C1(n6921), .C2(n6920), .A(n9915), .B(n6919), .ZN(n6929)
         );
  AOI211_X1 U8825 ( .C1(n6924), .C2(n6923), .A(n9928), .B(n6922), .ZN(n6928)
         );
  INV_X1 U8826 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n9079) );
  NAND2_X1 U8827 ( .A1(n9959), .A2(n6925), .ZN(n6926) );
  NAND2_X1 U8828 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n7327) );
  OAI211_X1 U8829 ( .C1(n9079), .C2(n9970), .A(n6926), .B(n7327), .ZN(n6927)
         );
  OR3_X1 U8830 ( .A1(n6929), .A2(n6928), .A3(n6927), .ZN(P1_U3249) );
  AOI211_X1 U8831 ( .C1(n6932), .C2(n6931), .A(n9928), .B(n6930), .ZN(n6941)
         );
  AOI211_X1 U8832 ( .C1(n6935), .C2(n6934), .A(n9915), .B(n6933), .ZN(n6940)
         );
  INV_X1 U8833 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n6938) );
  NAND2_X1 U8834 ( .A1(n9959), .A2(n6936), .ZN(n6937) );
  NAND2_X1 U8835 ( .A1(P1_U3086), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n7430) );
  OAI211_X1 U8836 ( .C1(n6938), .C2(n9970), .A(n6937), .B(n7430), .ZN(n6939)
         );
  OR3_X1 U8837 ( .A1(n6941), .A2(n6940), .A3(n6939), .ZN(P1_U3250) );
  AOI211_X1 U8838 ( .C1(n6944), .C2(n6943), .A(n9928), .B(n6942), .ZN(n6953)
         );
  AOI211_X1 U8839 ( .C1(n6947), .C2(n6946), .A(n9915), .B(n6945), .ZN(n6952)
         );
  INV_X1 U8840 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n6950) );
  NAND2_X1 U8841 ( .A1(n9959), .A2(n6948), .ZN(n6949) );
  NAND2_X1 U8842 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_U3086), .ZN(n7673) );
  OAI211_X1 U8843 ( .C1(n6950), .C2(n9970), .A(n6949), .B(n7673), .ZN(n6951)
         );
  OR3_X1 U8844 ( .A1(n6953), .A2(n6952), .A3(n6951), .ZN(P1_U3251) );
  INV_X1 U8845 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n6956) );
  OAI222_X1 U8846 ( .A1(n7680), .A2(n6956), .B1(n9897), .B2(n6955), .C1(n6954), 
        .C2(P1_U3086), .ZN(P1_U3342) );
  INV_X1 U8847 ( .A(n6957), .ZN(n7022) );
  AOI22_X1 U8848 ( .A1(n9908), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n9894), .ZN(n6958) );
  OAI21_X1 U8849 ( .B1(n7022), .B2(n9897), .A(n6958), .ZN(P1_U3341) );
  OAI21_X1 U8850 ( .B1(n6961), .B2(n6959), .A(n6960), .ZN(n6962) );
  NAND2_X1 U8851 ( .A1(n6962), .A2(n8216), .ZN(n6967) );
  OAI22_X1 U8852 ( .A1(n8266), .A2(n6963), .B1(n6621), .B2(n8285), .ZN(n6964)
         );
  AOI21_X1 U8853 ( .B1(n6965), .B2(n8276), .A(n6964), .ZN(n6966) );
  OAI211_X1 U8854 ( .C1(n6968), .C2(n10166), .A(n6967), .B(n6966), .ZN(
        P2_U3177) );
  INV_X1 U8855 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n6974) );
  AND2_X1 U8856 ( .A1(n7596), .A2(n8911), .ZN(n6972) );
  OR2_X1 U8857 ( .A1(n6963), .A2(n8848), .ZN(n7014) );
  OAI21_X1 U8858 ( .B1(n7396), .B2(n6969), .A(n7014), .ZN(n6970) );
  INV_X1 U8859 ( .A(n6970), .ZN(n6971) );
  OAI21_X1 U8860 ( .B1(n8480), .B2(n6972), .A(n6971), .ZN(n9149) );
  NAND2_X1 U8861 ( .A1(n9149), .A2(n10185), .ZN(n6973) );
  OAI21_X1 U8862 ( .B1(n6974), .B2(n10185), .A(n6973), .ZN(P2_U3390) );
  OR2_X1 U8863 ( .A1(n6976), .A2(n6975), .ZN(n6977) );
  NAND2_X1 U8864 ( .A1(n6978), .A2(n6977), .ZN(n9515) );
  OR2_X1 U8865 ( .A1(n6980), .A2(n6979), .ZN(n7118) );
  AOI22_X1 U8866 ( .A1(n9444), .A2(n10058), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        n7118), .ZN(n6982) );
  NAND2_X1 U8867 ( .A1(n9451), .A2(n7348), .ZN(n6981) );
  OAI211_X1 U8868 ( .C1(n9515), .C2(n9458), .A(n6982), .B(n6981), .ZN(P1_U3232) );
  XNOR2_X1 U8869 ( .A(n6984), .B(n6983), .ZN(n6994) );
  XOR2_X1 U8870 ( .A(n6985), .B(P2_REG1_REG_5__SCAN_IN), .Z(n6992) );
  INV_X1 U8871 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n6990) );
  AND2_X1 U8872 ( .A1(P2_U3151), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n7236) );
  AOI21_X1 U8873 ( .B1(n8631), .B2(n5052), .A(n7236), .ZN(n6989) );
  OAI21_X1 U8874 ( .B1(P2_REG2_REG_5__SCAN_IN), .B2(n4372), .A(n6986), .ZN(
        n6987) );
  NAND2_X1 U8875 ( .A1(n6987), .A2(n8641), .ZN(n6988) );
  OAI211_X1 U8876 ( .C1(n6990), .C2(n8634), .A(n6989), .B(n6988), .ZN(n6991)
         );
  AOI21_X1 U8877 ( .B1(n8541), .B2(n6992), .A(n6991), .ZN(n6993) );
  OAI21_X1 U8878 ( .B1(n6994), .B2(n8626), .A(n6993), .ZN(P2_U3187) );
  NAND2_X1 U8879 ( .A1(n6997), .A2(n6996), .ZN(n6998) );
  AND2_X1 U8880 ( .A1(n10062), .A2(n6998), .ZN(n6999) );
  NAND2_X1 U8881 ( .A1(n6999), .A2(n10063), .ZN(n10053) );
  OR2_X1 U8882 ( .A1(n7000), .A2(n7886), .ZN(n10078) );
  NAND2_X1 U8883 ( .A1(n5896), .A2(n8022), .ZN(n7986) );
  NAND2_X1 U8884 ( .A1(n6602), .A2(n7886), .ZN(n7001) );
  INV_X1 U8885 ( .A(n10058), .ZN(n7642) );
  NAND2_X1 U8886 ( .A1(n7346), .A2(n7642), .ZN(n7902) );
  INV_X1 U8887 ( .A(n7902), .ZN(n7002) );
  OR2_X1 U8888 ( .A1(n7637), .A2(n7002), .ZN(n10064) );
  OAI21_X1 U8889 ( .B1(n10136), .B2(n10013), .A(n10064), .ZN(n7005) );
  NOR2_X1 U8890 ( .A1(n4441), .A2(n10048), .ZN(n10061) );
  NOR2_X1 U8891 ( .A1(n10062), .A2(n7642), .ZN(n7003) );
  NOR2_X1 U8892 ( .A1(n10061), .A2(n7003), .ZN(n7004) );
  AND2_X1 U8893 ( .A1(n7005), .A2(n7004), .ZN(n10077) );
  NAND2_X1 U8894 ( .A1(n10160), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n7006) );
  OAI21_X1 U8895 ( .B1(n10160), .B2(n10077), .A(n7006), .ZN(P1_U3522) );
  NOR2_X1 U8896 ( .A1(n7007), .A2(n5772), .ZN(n7008) );
  OR2_X1 U8897 ( .A1(n7009), .A2(n7008), .ZN(n7010) );
  INV_X1 U8898 ( .A(n7012), .ZN(n7013) );
  NOR3_X1 U8899 ( .A1(n8480), .A2(n7013), .A3(n8998), .ZN(n7016) );
  INV_X1 U8900 ( .A(n7014), .ZN(n7015) );
  OAI21_X1 U8901 ( .B1(n7016), .B2(n7015), .A(n10171), .ZN(n7021) );
  INV_X1 U8902 ( .A(n7017), .ZN(n7018) );
  INV_X1 U8903 ( .A(n10163), .ZN(n8833) );
  NAND2_X1 U8904 ( .A1(n7018), .A2(n8833), .ZN(n8784) );
  AOI22_X1 U8905 ( .A1(n8921), .A2(n7019), .B1(P2_REG3_REG_0__SCAN_IN), .B2(
        n8920), .ZN(n7020) );
  OAI211_X1 U8906 ( .C1(n5134), .C2(n10171), .A(n7021), .B(n7020), .ZN(
        P2_U3233) );
  INV_X1 U8907 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n9119) );
  OAI222_X1 U8908 ( .A1(n9283), .A2(n9119), .B1(n9281), .B2(n7022), .C1(n8557), 
        .C2(P2_U3151), .ZN(P2_U3281) );
  INV_X1 U8909 ( .A(n7023), .ZN(n7027) );
  OAI21_X1 U8910 ( .B1(n7062), .B2(n7025), .A(n7024), .ZN(n7026) );
  NAND3_X1 U8911 ( .A1(n7027), .A2(n7084), .A3(n7026), .ZN(n7045) );
  INV_X1 U8912 ( .A(n7028), .ZN(n7029) );
  OAI21_X1 U8913 ( .B1(n7031), .B2(n7030), .A(n7029), .ZN(n7043) );
  INV_X1 U8914 ( .A(n7032), .ZN(n7034) );
  NAND3_X1 U8915 ( .A1(n7066), .A2(n7034), .A3(n7033), .ZN(n7035) );
  AOI21_X1 U8916 ( .B1(n7036), .B2(n7035), .A(n4586), .ZN(n7042) );
  INV_X1 U8917 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n7040) );
  INV_X1 U8918 ( .A(n7037), .ZN(n7038) );
  AND2_X1 U8919 ( .A1(P2_U3151), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n7162) );
  AOI21_X1 U8920 ( .B1(n8631), .B2(n7038), .A(n7162), .ZN(n7039) );
  OAI21_X1 U8921 ( .B1(n7040), .B2(n8634), .A(n7039), .ZN(n7041) );
  AOI211_X1 U8922 ( .C1(n8541), .C2(n7043), .A(n7042), .B(n7041), .ZN(n7044)
         );
  NAND2_X1 U8923 ( .A1(n7045), .A2(n7044), .ZN(P2_U3186) );
  XNOR2_X1 U8924 ( .A(n7047), .B(n7046), .ZN(n7061) );
  INV_X1 U8925 ( .A(n7083), .ZN(n7052) );
  NOR3_X1 U8926 ( .A1(n7050), .A2(n7049), .A3(n7048), .ZN(n7051) );
  OAI21_X1 U8927 ( .B1(n7052), .B2(n7051), .A(n7084), .ZN(n7060) );
  OAI21_X1 U8928 ( .B1(P2_REG2_REG_7__SCAN_IN), .B2(n7054), .A(n7053), .ZN(
        n7058) );
  INV_X1 U8929 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n7056) );
  AND2_X1 U8930 ( .A1(P2_U3151), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n7446) );
  AOI21_X1 U8931 ( .B1(n8631), .B2(n5065), .A(n7446), .ZN(n7055) );
  OAI21_X1 U8932 ( .B1(n7056), .B2(n8634), .A(n7055), .ZN(n7057) );
  AOI21_X1 U8933 ( .B1(n7058), .B2(n8641), .A(n7057), .ZN(n7059) );
  OAI211_X1 U8934 ( .C1(n7061), .C2(n8645), .A(n7060), .B(n7059), .ZN(P2_U3189) );
  AOI21_X1 U8935 ( .B1(n7064), .B2(n7063), .A(n7062), .ZN(n7076) );
  XNOR2_X1 U8936 ( .A(n7065), .B(P2_REG1_REG_3__SCAN_IN), .ZN(n7074) );
  INV_X1 U8937 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n7072) );
  OAI21_X1 U8938 ( .B1(P2_REG2_REG_3__SCAN_IN), .B2(n7067), .A(n7066), .ZN(
        n7070) );
  NOR2_X1 U8939 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7142), .ZN(n7133) );
  NOR2_X1 U8940 ( .A1(n8615), .A2(n7068), .ZN(n7069) );
  AOI211_X1 U8941 ( .C1(n8641), .C2(n7070), .A(n7133), .B(n7069), .ZN(n7071)
         );
  OAI21_X1 U8942 ( .B1(n8634), .B2(n7072), .A(n7071), .ZN(n7073) );
  AOI21_X1 U8943 ( .B1(n8541), .B2(n7074), .A(n7073), .ZN(n7075) );
  OAI21_X1 U8944 ( .B1(n7076), .B2(n8626), .A(n7075), .ZN(P2_U3185) );
  INV_X1 U8945 ( .A(n7077), .ZN(n7078) );
  AOI21_X1 U8946 ( .B1(n7080), .B2(n7079), .A(n7078), .ZN(n7096) );
  AND3_X1 U8947 ( .A1(n7083), .A2(n7082), .A3(n7081), .ZN(n7085) );
  OAI21_X1 U8948 ( .B1(n7208), .B2(n7085), .A(n7084), .ZN(n7095) );
  NAND2_X1 U8949 ( .A1(P2_U3151), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n8150) );
  OAI21_X1 U8950 ( .B1(n8615), .B2(n7086), .A(n8150), .ZN(n7093) );
  INV_X1 U8951 ( .A(n7087), .ZN(n7089) );
  NAND3_X1 U8952 ( .A1(n7053), .A2(n7089), .A3(n7088), .ZN(n7090) );
  AOI21_X1 U8953 ( .B1(n7091), .B2(n7090), .A(n4586), .ZN(n7092) );
  AOI211_X1 U8954 ( .C1(n8611), .C2(P2_ADDR_REG_8__SCAN_IN), .A(n7093), .B(
        n7092), .ZN(n7094) );
  OAI211_X1 U8955 ( .C1(n7096), .C2(n8645), .A(n7095), .B(n7094), .ZN(P2_U3190) );
  INV_X1 U8956 ( .A(n7097), .ZN(n7098) );
  AOI21_X1 U8957 ( .B1(n7099), .B2(n8484), .A(n7098), .ZN(n7229) );
  XNOR2_X1 U8958 ( .A(n6620), .B(n7100), .ZN(n7101) );
  AOI222_X1 U8959 ( .A1(n8887), .A2(n7101), .B1(n8538), .B2(n8917), .C1(n4937), 
        .C2(n8890), .ZN(n7225) );
  OAI21_X1 U8960 ( .B1(n7596), .B2(n7229), .A(n7225), .ZN(n7154) );
  INV_X1 U8961 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n7102) );
  OAI22_X1 U8962 ( .A1(n7103), .A2(n9264), .B1(n10185), .B2(n7102), .ZN(n7104)
         );
  AOI21_X1 U8963 ( .B1(n7154), .B2(n10185), .A(n7104), .ZN(n7105) );
  INV_X1 U8964 ( .A(n7105), .ZN(P2_U3393) );
  INV_X1 U8965 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n7108) );
  INV_X1 U8966 ( .A(n7106), .ZN(n7109) );
  OAI222_X1 U8967 ( .A1(n7680), .A2(n7108), .B1(n9897), .B2(n7109), .C1(
        P1_U3086), .C2(n7107), .ZN(P1_U3340) );
  INV_X1 U8968 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n7110) );
  OAI222_X1 U8969 ( .A1(n9283), .A2(n7110), .B1(n9281), .B2(n7109), .C1(n8576), 
        .C2(P2_U3151), .ZN(P2_U3280) );
  XOR2_X1 U8970 ( .A(n7112), .B(n7111), .Z(n7115) );
  AOI22_X1 U8971 ( .A1(n9482), .A2(n7346), .B1(n9451), .B2(n7352), .ZN(n7114)
         );
  AOI22_X1 U8972 ( .A1(n9444), .A2(n7903), .B1(P1_REG3_REG_1__SCAN_IN), .B2(
        n7118), .ZN(n7113) );
  OAI211_X1 U8973 ( .C1(n7115), .C2(n9458), .A(n7114), .B(n7113), .ZN(P1_U3222) );
  XOR2_X1 U8974 ( .A(n7117), .B(n7116), .Z(n7121) );
  AOI22_X1 U8975 ( .A1(n9451), .A2(n10011), .B1(n9482), .B2(n7348), .ZN(n7120)
         );
  AOI22_X1 U8976 ( .A1(n9444), .A2(n7353), .B1(P1_REG3_REG_2__SCAN_IN), .B2(
        n7118), .ZN(n7119) );
  OAI211_X1 U8977 ( .C1(n7121), .C2(n9458), .A(n7120), .B(n7119), .ZN(P1_U3237) );
  INV_X1 U8978 ( .A(n7122), .ZN(n7144) );
  AOI22_X1 U8979 ( .A1(n9938), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n9894), .ZN(n7123) );
  OAI21_X1 U8980 ( .B1(n7144), .B2(n9897), .A(n7123), .ZN(P1_U3338) );
  OR2_X1 U8981 ( .A1(n4274), .A2(n8463), .ZN(n7546) );
  NAND2_X1 U8982 ( .A1(n8894), .A2(n7546), .ZN(n7124) );
  NAND2_X1 U8983 ( .A1(n7125), .A2(n7126), .ZN(n7179) );
  XNOR2_X1 U8984 ( .A(n7179), .B(n8481), .ZN(n7173) );
  INV_X1 U8985 ( .A(n7173), .ZN(n7131) );
  XNOR2_X1 U8986 ( .A(n7127), .B(n8481), .ZN(n7128) );
  AOI222_X1 U8987 ( .A1(n8887), .A2(n7128), .B1(n8536), .B2(n8917), .C1(n8538), 
        .C2(n8890), .ZN(n7170) );
  MUX2_X1 U8988 ( .A(n4594), .B(n7170), .S(n10171), .Z(n7130) );
  AOI22_X1 U8989 ( .A1(n8921), .A2(n7132), .B1(n7142), .B2(n8920), .ZN(n7129)
         );
  OAI211_X1 U8990 ( .C1(n8855), .C2(n7131), .A(n7130), .B(n7129), .ZN(P2_U3230) );
  NAND2_X1 U8991 ( .A1(n8276), .A2(n7132), .ZN(n7135) );
  AOI21_X1 U8992 ( .B1(n8283), .B2(n8538), .A(n7133), .ZN(n7134) );
  OAI211_X1 U8993 ( .C1(n7136), .C2(n8285), .A(n7135), .B(n7134), .ZN(n7141)
         );
  AOI211_X1 U8994 ( .C1(n7139), .C2(n7137), .A(n8279), .B(n7138), .ZN(n7140)
         );
  AOI211_X1 U8995 ( .C1(n7142), .C2(n8288), .A(n7141), .B(n7140), .ZN(n7143)
         );
  INV_X1 U8996 ( .A(n7143), .ZN(P2_U3158) );
  OAI222_X1 U8997 ( .A1(n9283), .A2(n7145), .B1(n9281), .B2(n7144), .C1(n8614), 
        .C2(P2_U3151), .ZN(P2_U3278) );
  XOR2_X1 U8998 ( .A(n7146), .B(n7147), .Z(n7153) );
  AOI22_X1 U8999 ( .A1(n9444), .A2(n7493), .B1(n9451), .B2(n9500), .ZN(n7152)
         );
  NAND2_X1 U9000 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_U3086), .ZN(n9532) );
  INV_X1 U9001 ( .A(n9532), .ZN(n7148) );
  AOI21_X1 U9002 ( .B1(n9482), .B2(n7352), .A(n7148), .ZN(n7149) );
  OAI21_X1 U9003 ( .B1(n9479), .B2(P1_REG3_REG_3__SCAN_IN), .A(n7149), .ZN(
        n7150) );
  INV_X1 U9004 ( .A(n7150), .ZN(n7151) );
  OAI211_X1 U9005 ( .C1(n7153), .C2(n9458), .A(n7152), .B(n7151), .ZN(P1_U3218) );
  INV_X1 U9006 ( .A(n7154), .ZN(n7156) );
  INV_X1 U9007 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n9005) );
  AOI22_X1 U9008 ( .A1(n8979), .A2(n7226), .B1(n4269), .B2(
        P2_REG1_REG_1__SCAN_IN), .ZN(n7155) );
  OAI21_X1 U9009 ( .B1(n7156), .B2(n4269), .A(n7155), .ZN(P2_U3460) );
  INV_X1 U9010 ( .A(n7157), .ZN(n7160) );
  OAI222_X1 U9011 ( .A1(n9286), .A2(n7160), .B1(P2_U3151), .B2(n8589), .C1(
        n7158), .C2(n9283), .ZN(P2_U3279) );
  OAI222_X1 U9012 ( .A1(n7680), .A2(n9072), .B1(n9897), .B2(n7160), .C1(n4418), 
        .C2(P1_U3086), .ZN(P1_U3339) );
  OAI21_X1 U9013 ( .B1(n4373), .B2(n7161), .A(n7233), .ZN(n7168) );
  AOI21_X1 U9014 ( .B1(n8537), .B2(n8283), .A(n7162), .ZN(n7166) );
  NAND2_X1 U9015 ( .A1(n8288), .A2(n7218), .ZN(n7165) );
  NAND2_X1 U9016 ( .A1(n8276), .A2(n7219), .ZN(n7164) );
  NAND2_X1 U9017 ( .A1(n8264), .A2(n8535), .ZN(n7163) );
  NAND4_X1 U9018 ( .A1(n7166), .A2(n7165), .A3(n7164), .A4(n7163), .ZN(n7167)
         );
  AOI21_X1 U9019 ( .B1(n7168), .B2(n8216), .A(n7167), .ZN(n7169) );
  INV_X1 U9020 ( .A(n7169), .ZN(P2_U3170) );
  OAI21_X1 U9021 ( .B1(n7171), .B2(n7396), .A(n7170), .ZN(n7172) );
  AOI21_X1 U9022 ( .B1(n7173), .B2(n8999), .A(n7172), .ZN(n10177) );
  INV_X1 U9023 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n7174) );
  OR2_X1 U9024 ( .A1(n9003), .A2(n7174), .ZN(n7175) );
  OAI21_X1 U9025 ( .B1(n10177), .B2(n4269), .A(n7175), .ZN(P2_U3462) );
  NAND2_X1 U9026 ( .A1(n8312), .A2(n8316), .ZN(n8485) );
  INV_X1 U9027 ( .A(n8485), .ZN(n8309) );
  XNOR2_X1 U9028 ( .A(n7176), .B(n8309), .ZN(n7177) );
  OAI222_X1 U9029 ( .A1(n8848), .A2(n7292), .B1(n8905), .B2(n6621), .C1(n8911), 
        .C2(n7177), .ZN(n7215) );
  INV_X1 U9030 ( .A(n7178), .ZN(n8318) );
  AOI21_X1 U9031 ( .B1(n7179), .B2(n8481), .A(n8318), .ZN(n7180) );
  XNOR2_X1 U9032 ( .A(n7180), .B(n8309), .ZN(n7222) );
  OAI22_X1 U9033 ( .A1(n7222), .A2(n7596), .B1(n7181), .B2(n7396), .ZN(n7182)
         );
  NOR2_X1 U9034 ( .A1(n7215), .A2(n7182), .ZN(n10179) );
  NAND2_X1 U9035 ( .A1(n4269), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n7183) );
  OAI21_X1 U9036 ( .B1(n10179), .B2(n4269), .A(n7183), .ZN(P2_U3463) );
  OAI21_X1 U9037 ( .B1(n7184), .B2(n8486), .A(n7125), .ZN(n10169) );
  NOR2_X1 U9038 ( .A1(n10164), .A2(n7396), .ZN(n7189) );
  XNOR2_X1 U9039 ( .A(n7185), .B(n8486), .ZN(n7188) );
  INV_X1 U9040 ( .A(n8894), .ZN(n7392) );
  OAI22_X1 U9041 ( .A1(n6963), .A2(n8905), .B1(n6621), .B2(n8848), .ZN(n7186)
         );
  AOI21_X1 U9042 ( .B1(n10169), .B2(n7392), .A(n7186), .ZN(n7187) );
  OAI21_X1 U9043 ( .B1(n7188), .B2(n8911), .A(n7187), .ZN(n10167) );
  AOI211_X1 U9044 ( .C1(n8993), .C2(n10169), .A(n7189), .B(n10167), .ZN(n10175) );
  NAND2_X1 U9045 ( .A1(n4269), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n7190) );
  OAI21_X1 U9046 ( .B1(n10175), .B2(n4269), .A(n7190), .ZN(P2_U3461) );
  INV_X1 U9047 ( .A(n7191), .ZN(n7224) );
  OAI222_X1 U9048 ( .A1(n9286), .A2(n7224), .B1(P2_U3151), .B2(n8629), .C1(
        n9118), .C2(n9283), .ZN(P2_U3277) );
  XNOR2_X1 U9049 ( .A(n7193), .B(n8478), .ZN(n7197) );
  XNOR2_X1 U9050 ( .A(n7194), .B(n8478), .ZN(n7198) );
  OAI22_X1 U9051 ( .A1(n7390), .A2(n8848), .B1(n7136), .B2(n8905), .ZN(n7195)
         );
  AOI21_X1 U9052 ( .B1(n7198), .B2(n7392), .A(n7195), .ZN(n7196) );
  OAI21_X1 U9053 ( .B1(n7197), .B2(n8911), .A(n7196), .ZN(n7253) );
  INV_X1 U9054 ( .A(n7198), .ZN(n7260) );
  OAI22_X1 U9055 ( .A1(n7260), .A2(n7397), .B1(n7199), .B2(n7396), .ZN(n7200)
         );
  NOR2_X1 U9056 ( .A1(n7253), .A2(n7200), .ZN(n10181) );
  OR2_X1 U9057 ( .A1(n9003), .A2(n5125), .ZN(n7201) );
  OAI21_X1 U9058 ( .B1(n10181), .B2(n4269), .A(n7201), .ZN(P2_U3464) );
  XNOR2_X1 U9059 ( .A(n7202), .B(n8994), .ZN(n7214) );
  OAI21_X1 U9060 ( .B1(P2_REG2_REG_9__SCAN_IN), .B2(n7204), .A(n7203), .ZN(
        n7212) );
  NAND2_X1 U9061 ( .A1(P2_U3151), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n8220) );
  NAND2_X1 U9062 ( .A1(n8611), .A2(P2_ADDR_REG_9__SCAN_IN), .ZN(n7205) );
  OAI211_X1 U9063 ( .C1(n8615), .C2(n4796), .A(n8220), .B(n7205), .ZN(n7211)
         );
  OR3_X1 U9064 ( .A1(n7208), .A2(n7207), .A3(n7206), .ZN(n7209) );
  AOI21_X1 U9065 ( .B1(n7275), .B2(n7209), .A(n8626), .ZN(n7210) );
  AOI211_X1 U9066 ( .C1(n8641), .C2(n7212), .A(n7211), .B(n7210), .ZN(n7213)
         );
  OAI21_X1 U9067 ( .B1(n7214), .B2(n8645), .A(n7213), .ZN(P2_U3191) );
  INV_X1 U9068 ( .A(n7215), .ZN(n7216) );
  MUX2_X1 U9069 ( .A(n7217), .B(n7216), .S(n10171), .Z(n7221) );
  AOI22_X1 U9070 ( .A1(n8921), .A2(n7219), .B1(n8920), .B2(n7218), .ZN(n7220)
         );
  OAI211_X1 U9071 ( .C1(n8855), .C2(n7222), .A(n7221), .B(n7220), .ZN(P2_U3229) );
  INV_X1 U9072 ( .A(n9958), .ZN(n7223) );
  OAI222_X1 U9073 ( .A1(n7680), .A2(n9104), .B1(n9897), .B2(n7224), .C1(n7223), 
        .C2(P1_U3086), .ZN(P1_U3337) );
  MUX2_X1 U9074 ( .A(n4468), .B(n7225), .S(n10171), .Z(n7228) );
  AOI22_X1 U9075 ( .A1(n8921), .A2(n7226), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        n8920), .ZN(n7227) );
  OAI211_X1 U9076 ( .C1(n7229), .C2(n8855), .A(n7228), .B(n7227), .ZN(P2_U3232) );
  INV_X1 U9077 ( .A(n7230), .ZN(n7235) );
  NAND3_X1 U9078 ( .A1(n7233), .A2(n7232), .A3(n7231), .ZN(n7234) );
  AOI21_X1 U9079 ( .B1(n7235), .B2(n7234), .A(n8279), .ZN(n7242) );
  AOI21_X1 U9080 ( .B1(n8536), .B2(n8283), .A(n7236), .ZN(n7240) );
  NAND2_X1 U9081 ( .A1(n8288), .A2(n7256), .ZN(n7239) );
  NAND2_X1 U9082 ( .A1(n8276), .A2(n7257), .ZN(n7238) );
  NAND2_X1 U9083 ( .A1(n8264), .A2(n8534), .ZN(n7237) );
  NAND4_X1 U9084 ( .A1(n7240), .A2(n7239), .A3(n7238), .A4(n7237), .ZN(n7241)
         );
  OR2_X1 U9085 ( .A1(n7242), .A2(n7241), .ZN(P2_U3167) );
  NAND2_X1 U9086 ( .A1(n7243), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n7244) );
  OR2_X1 U9087 ( .A1(n8081), .A2(n7244), .ZN(n7251) );
  INV_X1 U9088 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n7248) );
  NAND2_X1 U9089 ( .A1(n6060), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n7246) );
  NAND2_X1 U9090 ( .A1(n7878), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n7245) );
  OAI211_X1 U9091 ( .C1(n7248), .C2(n7247), .A(n7246), .B(n7245), .ZN(n7249)
         );
  INV_X1 U9092 ( .A(n7249), .ZN(n7250) );
  NAND2_X1 U9093 ( .A1(n9501), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n7252) );
  OAI21_X1 U9094 ( .B1(n9591), .B2(n9501), .A(n7252), .ZN(P1_U3583) );
  INV_X1 U9095 ( .A(n7546), .ZN(n10170) );
  NAND2_X1 U9096 ( .A1(n10171), .A2(n10170), .ZN(n8901) );
  INV_X1 U9097 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n7255) );
  INV_X1 U9098 ( .A(n7253), .ZN(n7254) );
  MUX2_X1 U9099 ( .A(n7255), .B(n7254), .S(n10171), .Z(n7259) );
  AOI22_X1 U9100 ( .A1(n8921), .A2(n7257), .B1(n8920), .B2(n7256), .ZN(n7258)
         );
  OAI211_X1 U9101 ( .C1(n7260), .C2(n8901), .A(n7259), .B(n7258), .ZN(P2_U3228) );
  INV_X1 U9102 ( .A(n7339), .ZN(n7269) );
  INV_X1 U9103 ( .A(n8288), .ZN(n8255) );
  OAI211_X1 U9104 ( .C1(n7263), .C2(n7262), .A(n7261), .B(n8216), .ZN(n7268)
         );
  NAND2_X1 U9105 ( .A1(n8283), .A2(n8535), .ZN(n7264) );
  OAI211_X1 U9106 ( .C1(n8906), .C2(n8285), .A(n7265), .B(n7264), .ZN(n7266)
         );
  AOI21_X1 U9107 ( .B1(n7340), .B2(n8276), .A(n7266), .ZN(n7267) );
  OAI211_X1 U9108 ( .C1(n7269), .C2(n8255), .A(n7268), .B(n7267), .ZN(P2_U3179) );
  XOR2_X1 U9109 ( .A(n7271), .B(n7270), .Z(n7287) );
  NAND2_X1 U9110 ( .A1(P2_U3151), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n8117) );
  OAI21_X1 U9111 ( .B1(n8615), .B2(n7272), .A(n8117), .ZN(n7279) );
  INV_X1 U9112 ( .A(n7480), .ZN(n7277) );
  NAND3_X1 U9113 ( .A1(n7275), .A2(n7274), .A3(n7273), .ZN(n7276) );
  AOI21_X1 U9114 ( .B1(n7277), .B2(n7276), .A(n8626), .ZN(n7278) );
  AOI211_X1 U9115 ( .C1(n8611), .C2(P2_ADDR_REG_10__SCAN_IN), .A(n7279), .B(
        n7278), .ZN(n7286) );
  INV_X1 U9116 ( .A(n7203), .ZN(n7283) );
  INV_X1 U9117 ( .A(n7280), .ZN(n7282) );
  NOR3_X1 U9118 ( .A1(n7283), .A2(n7282), .A3(n7281), .ZN(n7284) );
  OAI21_X1 U9119 ( .B1(n7284), .B2(n4357), .A(n8641), .ZN(n7285) );
  OAI211_X1 U9120 ( .C1(n7287), .C2(n8645), .A(n7286), .B(n7285), .ZN(P2_U3192) );
  INV_X1 U9121 ( .A(n7288), .ZN(n8095) );
  OAI222_X1 U9122 ( .A1(n7680), .A2(n7289), .B1(n9897), .B2(n8095), .C1(n6294), 
        .C2(P1_U3086), .ZN(P1_U3336) );
  INV_X1 U9123 ( .A(n8315), .ZN(n8322) );
  NOR2_X1 U9124 ( .A1(n8321), .A2(n8322), .ZN(n8487) );
  XNOR2_X1 U9125 ( .A(n7290), .B(n8487), .ZN(n7291) );
  OAI222_X1 U9126 ( .A1(n8905), .A2(n7292), .B1(n8848), .B2(n8906), .C1(n7291), 
        .C2(n8911), .ZN(n7336) );
  INV_X1 U9127 ( .A(n8487), .ZN(n7293) );
  XNOR2_X1 U9128 ( .A(n7294), .B(n7293), .ZN(n7343) );
  OAI22_X1 U9129 ( .A1(n7343), .A2(n7596), .B1(n7295), .B2(n7396), .ZN(n7296)
         );
  NOR2_X1 U9130 ( .A1(n7336), .A2(n7296), .ZN(n10183) );
  NAND2_X1 U9131 ( .A1(n4269), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n7297) );
  OAI21_X1 U9132 ( .B1(n10183), .B2(n4269), .A(n7297), .ZN(P2_U3465) );
  OAI21_X1 U9133 ( .B1(n7300), .B2(n7299), .A(n7298), .ZN(n7301) );
  INV_X1 U9134 ( .A(n7301), .ZN(n7311) );
  OAI21_X1 U9135 ( .B1(n7304), .B2(n7303), .A(n7302), .ZN(n7309) );
  INV_X1 U9136 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n7307) );
  NAND2_X1 U9137 ( .A1(n9959), .A2(n7305), .ZN(n7306) );
  NAND2_X1 U9138 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n7699) );
  OAI211_X1 U9139 ( .C1(n7307), .C2(n9970), .A(n7306), .B(n7699), .ZN(n7308)
         );
  AOI21_X1 U9140 ( .B1(n7309), .B2(n9964), .A(n7308), .ZN(n7310) );
  OAI21_X1 U9141 ( .B1(n7311), .B2(n9928), .A(n7310), .ZN(P1_U3255) );
  NAND2_X1 U9142 ( .A1(n7313), .A2(n7312), .ZN(n7315) );
  XNOR2_X1 U9143 ( .A(n7315), .B(n7314), .ZN(n7322) );
  AOI22_X1 U9144 ( .A1(n9444), .A2(n7592), .B1(n9482), .B2(n9500), .ZN(n7321)
         );
  INV_X1 U9145 ( .A(n7316), .ZN(n7317) );
  AOI21_X1 U9146 ( .B1(n9451), .B2(n9499), .A(n7317), .ZN(n7318) );
  OAI21_X1 U9147 ( .B1(n9479), .B2(n7590), .A(n7318), .ZN(n7319) );
  INV_X1 U9148 ( .A(n7319), .ZN(n7320) );
  OAI211_X1 U9149 ( .C1(n7322), .C2(n9458), .A(n7321), .B(n7320), .ZN(P1_U3227) );
  XNOR2_X1 U9150 ( .A(n7325), .B(n7324), .ZN(n7326) );
  XNOR2_X1 U9151 ( .A(n7323), .B(n7326), .ZN(n7333) );
  AOI22_X1 U9152 ( .A1(n9444), .A2(n10001), .B1(n9482), .B2(n7358), .ZN(n7332)
         );
  INV_X1 U9153 ( .A(n7327), .ZN(n7328) );
  AOI21_X1 U9154 ( .B1(n9451), .B2(n9992), .A(n7328), .ZN(n7329) );
  OAI21_X1 U9155 ( .B1(n9479), .B2(n9994), .A(n7329), .ZN(n7330) );
  INV_X1 U9156 ( .A(n7330), .ZN(n7331) );
  OAI211_X1 U9157 ( .C1(n7333), .C2(n9458), .A(n7332), .B(n7331), .ZN(P1_U3239) );
  INV_X1 U9158 ( .A(n7334), .ZN(n7400) );
  OAI222_X1 U9159 ( .A1(n9286), .A2(n7400), .B1(n8503), .B2(P2_U3151), .C1(
        n7335), .C2(n9283), .ZN(P2_U3275) );
  INV_X1 U9160 ( .A(n7336), .ZN(n7337) );
  MUX2_X1 U9161 ( .A(n7338), .B(n7337), .S(n10171), .Z(n7342) );
  AOI22_X1 U9162 ( .A1(n8921), .A2(n7340), .B1(n8920), .B2(n7339), .ZN(n7341)
         );
  OAI211_X1 U9163 ( .C1(n8855), .C2(n7343), .A(n7342), .B(n7341), .ZN(P2_U3227) );
  NAND2_X1 U9164 ( .A1(n10007), .A2(n7906), .ZN(n7488) );
  INV_X1 U9165 ( .A(n7488), .ZN(n7345) );
  OR2_X1 U9166 ( .A1(n10011), .A2(n7493), .ZN(n10019) );
  NAND2_X1 U9167 ( .A1(n7345), .A2(n10019), .ZN(n7355) );
  NAND2_X1 U9168 ( .A1(n10035), .A2(n4441), .ZN(n7347) );
  NAND2_X1 U9169 ( .A1(n7347), .A2(n7903), .ZN(n7351) );
  INV_X1 U9170 ( .A(n10035), .ZN(n7349) );
  NAND2_X1 U9171 ( .A1(n7349), .A2(n7348), .ZN(n7350) );
  XNOR2_X2 U9172 ( .A(n7352), .B(n10086), .ZN(n10045) );
  NAND3_X1 U9173 ( .A1(n7351), .A2(n7350), .A3(n10045), .ZN(n7490) );
  NAND2_X1 U9174 ( .A1(n7356), .A2(n10018), .ZN(n7913) );
  NAND3_X1 U9175 ( .A1(n7355), .A2(n7354), .A3(n10024), .ZN(n7581) );
  NAND2_X1 U9176 ( .A1(n7356), .A2(n10096), .ZN(n7580) );
  NAND2_X1 U9177 ( .A1(n7359), .A2(n10104), .ZN(n9996) );
  AND2_X1 U9178 ( .A1(n7580), .A2(n9996), .ZN(n7357) );
  NAND2_X1 U9179 ( .A1(n7373), .A2(n9996), .ZN(n7361) );
  NAND2_X1 U9180 ( .A1(n7788), .A2(n7794), .ZN(n9999) );
  OR2_X1 U9181 ( .A1(n10001), .A2(n9499), .ZN(n7362) );
  NAND2_X1 U9182 ( .A1(n7363), .A2(n7362), .ZN(n7416) );
  XNOR2_X1 U9183 ( .A(n9975), .B(n7429), .ZN(n7415) );
  INV_X1 U9184 ( .A(n7415), .ZN(n7790) );
  XNOR2_X1 U9185 ( .A(n7416), .B(n7790), .ZN(n10115) );
  NOR2_X1 U9186 ( .A1(n7365), .A2(n7364), .ZN(n7368) );
  INV_X1 U9187 ( .A(n7366), .ZN(n7367) );
  NAND2_X1 U9188 ( .A1(n7368), .A2(n7367), .ZN(n7379) );
  INV_X1 U9189 ( .A(n7420), .ZN(n7369) );
  AND2_X1 U9190 ( .A1(n10070), .A2(n7369), .ZN(n10055) );
  INV_X1 U9191 ( .A(n10055), .ZN(n7644) );
  XNOR2_X2 U9192 ( .A(n10049), .B(n7370), .ZN(n7960) );
  NAND2_X1 U9193 ( .A1(n7352), .A2(n10086), .ZN(n7905) );
  INV_X1 U9194 ( .A(n7407), .ZN(n9991) );
  INV_X1 U9195 ( .A(n7788), .ZN(n7405) );
  AOI21_X1 U9196 ( .B1(n9991), .B2(n7794), .A(n7405), .ZN(n7374) );
  NAND2_X1 U9197 ( .A1(n7374), .A2(n7790), .ZN(n7500) );
  OAI21_X1 U9198 ( .B1(n7374), .B2(n7790), .A(n7500), .ZN(n7375) );
  NAND2_X1 U9199 ( .A1(n7375), .A2(n10013), .ZN(n7377) );
  AOI22_X1 U9200 ( .A1(n10009), .A2(n9498), .B1(n9499), .B2(n10010), .ZN(n7376) );
  OAI211_X1 U9201 ( .C1(n10053), .C2(n10115), .A(n7377), .B(n7376), .ZN(n10118) );
  NAND2_X1 U9202 ( .A1(n10118), .A2(n10070), .ZN(n7383) );
  OAI22_X1 U9203 ( .A1(n10070), .A2(n6579), .B1(n7433), .B2(n10068), .ZN(n7381) );
  INV_X1 U9204 ( .A(n10002), .ZN(n7378) );
  INV_X1 U9205 ( .A(n7429), .ZN(n10117) );
  OAI211_X1 U9206 ( .C1(n7378), .C2(n10117), .A(n10027), .B(n9985), .ZN(n10116) );
  OR2_X1 U9207 ( .A1(n7379), .A2(n6602), .ZN(n9581) );
  NOR2_X1 U9208 ( .A1(n10116), .A2(n9581), .ZN(n7380) );
  AOI211_X1 U9209 ( .C1(n10017), .C2(n7429), .A(n7381), .B(n7380), .ZN(n7382)
         );
  OAI211_X1 U9210 ( .C1(n10115), .C2(n7644), .A(n7383), .B(n7382), .ZN(
        P1_U3286) );
  NOR2_X1 U9211 ( .A1(n7385), .A2(n8479), .ZN(n8907) );
  AOI21_X1 U9212 ( .B1(n8479), .B2(n7385), .A(n8907), .ZN(n7394) );
  INV_X1 U9213 ( .A(n8859), .ZN(n7389) );
  INV_X1 U9214 ( .A(n8479), .ZN(n7388) );
  NAND2_X1 U9215 ( .A1(n8859), .A2(n8479), .ZN(n8903) );
  INV_X1 U9216 ( .A(n8903), .ZN(n7387) );
  AOI21_X1 U9217 ( .B1(n7389), .B2(n7388), .A(n7387), .ZN(n7395) );
  OAI22_X1 U9218 ( .A1(n7390), .A2(n8905), .B1(n8222), .B2(n8848), .ZN(n7391)
         );
  AOI21_X1 U9219 ( .B1(n7395), .B2(n7392), .A(n7391), .ZN(n7393) );
  OAI21_X1 U9220 ( .B1(n7394), .B2(n8911), .A(n7393), .ZN(n7548) );
  INV_X1 U9221 ( .A(n7395), .ZN(n7547) );
  OAI22_X1 U9222 ( .A1(n7547), .A2(n7397), .B1(n7553), .B2(n7396), .ZN(n7398)
         );
  NOR2_X1 U9223 ( .A1(n7548), .A2(n7398), .ZN(n10186) );
  NAND2_X1 U9224 ( .A1(n4269), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n7399) );
  OAI21_X1 U9225 ( .B1(n10186), .B2(n4269), .A(n7399), .ZN(P2_U3466) );
  OAI222_X1 U9226 ( .A1(n7680), .A2(n7401), .B1(P1_U3086), .B2(n6480), .C1(
        n9897), .C2(n7400), .ZN(P1_U3335) );
  OR2_X2 U9227 ( .A1(n9407), .A2(n9974), .ZN(n7818) );
  NAND2_X1 U9228 ( .A1(n7818), .A2(n7502), .ZN(n7808) );
  NAND2_X1 U9229 ( .A1(n9975), .A2(n7429), .ZN(n7499) );
  AND2_X1 U9230 ( .A1(n7807), .A2(n7499), .ZN(n7803) );
  NAND2_X1 U9231 ( .A1(n9407), .A2(n9974), .ZN(n7813) );
  NAND2_X1 U9232 ( .A1(n7402), .A2(n7813), .ZN(n7958) );
  INV_X1 U9233 ( .A(n7794), .ZN(n7403) );
  OR2_X2 U9234 ( .A1(n7958), .A2(n7403), .ZN(n7919) );
  NAND2_X1 U9235 ( .A1(n10117), .A2(n9992), .ZN(n7404) );
  AND2_X1 U9236 ( .A1(n7502), .A2(n7404), .ZN(n7804) );
  NAND2_X1 U9237 ( .A1(n7818), .A2(n7804), .ZN(n7959) );
  NOR2_X1 U9238 ( .A1(n7959), .A2(n7405), .ZN(n7406) );
  OR2_X1 U9239 ( .A1(n7958), .A2(n7406), .ZN(n7918) );
  INV_X1 U9240 ( .A(n7462), .ZN(n7556) );
  NAND2_X1 U9241 ( .A1(n10140), .A2(n9496), .ZN(n7823) );
  NAND2_X1 U9242 ( .A1(n9311), .A2(n7506), .ZN(n7820) );
  NAND2_X1 U9243 ( .A1(n7556), .A2(n7965), .ZN(n7555) );
  NAND2_X1 U9244 ( .A1(n7555), .A2(n7820), .ZN(n7408) );
  INV_X1 U9245 ( .A(n9495), .ZN(n7457) );
  OR2_X1 U9246 ( .A1(n9445), .A2(n7457), .ZN(n7822) );
  XNOR2_X1 U9247 ( .A(n7408), .B(n7968), .ZN(n7410) );
  OAI22_X1 U9248 ( .A1(n10050), .A2(n7506), .B1(n7459), .B2(n10048), .ZN(n7409) );
  AOI21_X1 U9249 ( .B1(n7410), .B2(n10013), .A(n7409), .ZN(n7439) );
  OAI22_X1 U9250 ( .A1(n10070), .A2(n7411), .B1(n9442), .B2(n10068), .ZN(n7414) );
  OAI211_X1 U9251 ( .C1(n7456), .C2(n7562), .A(n7412), .B(n10027), .ZN(n7438)
         );
  NOR2_X1 U9252 ( .A1(n7438), .A2(n9581), .ZN(n7413) );
  AOI211_X1 U9253 ( .C1(n10017), .C2(n9445), .A(n7414), .B(n7413), .ZN(n7423)
         );
  NAND2_X1 U9254 ( .A1(n7416), .A2(n7415), .ZN(n9972) );
  NAND2_X1 U9255 ( .A1(n10117), .A2(n9975), .ZN(n9971) );
  OR2_X1 U9256 ( .A1(n10122), .A2(n9498), .ZN(n7417) );
  AND2_X1 U9257 ( .A1(n9971), .A2(n7417), .ZN(n7419) );
  INV_X1 U9258 ( .A(n7417), .ZN(n7418) );
  NAND2_X1 U9259 ( .A1(n7502), .A2(n7807), .ZN(n9976) );
  NAND2_X1 U9260 ( .A1(n7818), .A2(n7813), .ZN(n7510) );
  XOR2_X1 U9261 ( .A(n7968), .B(n7458), .Z(n7441) );
  NAND2_X1 U9262 ( .A1(n10053), .A2(n7420), .ZN(n7421) );
  NAND2_X1 U9263 ( .A1(n7441), .A2(n10032), .ZN(n7422) );
  OAI211_X1 U9264 ( .C1(n7439), .C2(n4984), .A(n7423), .B(n7422), .ZN(P1_U3282) );
  INV_X1 U9265 ( .A(n7424), .ZN(n7426) );
  NOR2_X1 U9266 ( .A1(n7426), .A2(n7425), .ZN(n7427) );
  XNOR2_X1 U9267 ( .A(n7428), .B(n7427), .ZN(n7437) );
  AOI22_X1 U9268 ( .A1(n9444), .A2(n7429), .B1(n9482), .B2(n9499), .ZN(n7436)
         );
  INV_X1 U9269 ( .A(n7430), .ZN(n7431) );
  AOI21_X1 U9270 ( .B1(n9451), .B2(n9498), .A(n7431), .ZN(n7432) );
  OAI21_X1 U9271 ( .B1(n9479), .B2(n7433), .A(n7432), .ZN(n7434) );
  INV_X1 U9272 ( .A(n7434), .ZN(n7435) );
  OAI211_X1 U9273 ( .C1(n7437), .C2(n9458), .A(n7436), .B(n7435), .ZN(P1_U3213) );
  OAI211_X1 U9274 ( .C1(n7456), .C2(n10139), .A(n7439), .B(n7438), .ZN(n7440)
         );
  AOI21_X1 U9275 ( .B1(n10136), .B2(n7441), .A(n7440), .ZN(n7444) );
  NAND2_X1 U9276 ( .A1(n10160), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n7442) );
  OAI21_X1 U9277 ( .B1(n7444), .B2(n10160), .A(n7442), .ZN(P1_U3533) );
  NAND2_X1 U9278 ( .A1(n10144), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n7443) );
  OAI21_X1 U9279 ( .B1(n7444), .B2(n10144), .A(n7443), .ZN(P1_U3486) );
  NAND2_X1 U9280 ( .A1(n8276), .A2(n7445), .ZN(n7448) );
  AOI21_X1 U9281 ( .B1(n8283), .B2(n8534), .A(n7446), .ZN(n7447) );
  OAI211_X1 U9282 ( .C1(n8222), .C2(n8285), .A(n7448), .B(n7447), .ZN(n7454)
         );
  NAND2_X1 U9283 ( .A1(n7451), .A2(n7450), .ZN(n7452) );
  AOI21_X1 U9284 ( .B1(n7449), .B2(n7452), .A(n8279), .ZN(n7453) );
  AOI211_X1 U9285 ( .C1(n7550), .C2(n8288), .A(n7454), .B(n7453), .ZN(n7455)
         );
  INV_X1 U9286 ( .A(n7455), .ZN(P2_U3153) );
  NAND2_X1 U9287 ( .A1(n7705), .A2(n7459), .ZN(n7923) );
  XNOR2_X1 U9288 ( .A(n7614), .B(n4983), .ZN(n7569) );
  AOI21_X1 U9289 ( .B1(n7412), .B2(n7705), .A(n10039), .ZN(n7460) );
  NAND2_X1 U9290 ( .A1(n7460), .A2(n7617), .ZN(n7573) );
  OAI21_X1 U9291 ( .B1(n7461), .B2(n10139), .A(n7573), .ZN(n7470) );
  AND2_X1 U9292 ( .A1(n7825), .A2(n7820), .ZN(n7921) );
  NAND2_X1 U9293 ( .A1(n7462), .A2(n7921), .ZN(n7466) );
  INV_X1 U9294 ( .A(n7825), .ZN(n7463) );
  NAND2_X1 U9295 ( .A1(n7466), .A2(n7465), .ZN(n7467) );
  OAI211_X1 U9296 ( .C1(n7467), .C2(n4983), .A(n7623), .B(n10013), .ZN(n7469)
         );
  AOI22_X1 U9297 ( .A1(n9493), .A2(n10009), .B1(n10010), .B2(n9495), .ZN(n7468) );
  NAND2_X1 U9298 ( .A1(n7469), .A2(n7468), .ZN(n7575) );
  AOI211_X1 U9299 ( .C1(n7569), .C2(n10136), .A(n7470), .B(n7575), .ZN(n7473)
         );
  NAND2_X1 U9300 ( .A1(n10144), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n7471) );
  OAI21_X1 U9301 ( .B1(n7473), .B2(n10144), .A(n7471), .ZN(P1_U3489) );
  NAND2_X1 U9302 ( .A1(n10160), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n7472) );
  OAI21_X1 U9303 ( .B1(n7473), .B2(n10160), .A(n7472), .ZN(P1_U3534) );
  XNOR2_X1 U9304 ( .A(n7474), .B(P2_REG1_REG_11__SCAN_IN), .ZN(n7486) );
  OAI21_X1 U9305 ( .B1(P2_REG2_REG_11__SCAN_IN), .B2(n4362), .A(n7475), .ZN(
        n7484) );
  NAND2_X1 U9306 ( .A1(n8611), .A2(P2_ADDR_REG_11__SCAN_IN), .ZN(n7476) );
  NAND2_X1 U9307 ( .A1(P2_U3151), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n7630) );
  OAI211_X1 U9308 ( .C1(n8615), .C2(n7477), .A(n7476), .B(n7630), .ZN(n7483)
         );
  OR3_X1 U9309 ( .A1(n7480), .A2(n7479), .A3(n7478), .ZN(n7481) );
  AOI21_X1 U9310 ( .B1(n7524), .B2(n7481), .A(n8626), .ZN(n7482) );
  AOI211_X1 U9311 ( .C1(n8641), .C2(n7484), .A(n7483), .B(n7482), .ZN(n7485)
         );
  OAI21_X1 U9312 ( .B1(n7486), .B2(n8645), .A(n7485), .ZN(P2_U3193) );
  XNOR2_X1 U9313 ( .A(n7487), .B(n10021), .ZN(n7489) );
  AOI222_X1 U9314 ( .A1(n10013), .A2(n7489), .B1(n7352), .B2(n10010), .C1(
        n9500), .C2(n10009), .ZN(n10091) );
  NAND2_X1 U9315 ( .A1(n7490), .A2(n7491), .ZN(n10022) );
  XNOR2_X1 U9316 ( .A(n10021), .B(n10022), .ZN(n10094) );
  OAI211_X1 U9317 ( .C1(n10038), .C2(n10092), .A(n10027), .B(n10025), .ZN(
        n10090) );
  OAI22_X1 U9318 ( .A1(n9581), .A2(n10090), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        n10068), .ZN(n7492) );
  INV_X1 U9319 ( .A(n7492), .ZN(n7495) );
  NAND2_X1 U9320 ( .A1(n10017), .A2(n7493), .ZN(n7494) );
  OAI211_X1 U9321 ( .C1(n10070), .C2(n7496), .A(n7495), .B(n7494), .ZN(n7497)
         );
  AOI21_X1 U9322 ( .B1(n10032), .B2(n10094), .A(n7497), .ZN(n7498) );
  OAI21_X1 U9323 ( .B1(n10091), .B2(n4984), .A(n7498), .ZN(P1_U3290) );
  NAND2_X1 U9324 ( .A1(n7500), .A2(n7499), .ZN(n9977) );
  INV_X1 U9325 ( .A(n7807), .ZN(n7501) );
  AOI21_X1 U9326 ( .B1(n9977), .B2(n7502), .A(n7501), .ZN(n7503) );
  XOR2_X1 U9327 ( .A(n7510), .B(n7503), .Z(n7505) );
  OAI22_X1 U9328 ( .A1(n7505), .A2(n10047), .B1(n7504), .B2(n10050), .ZN(
        n10132) );
  XNOR2_X1 U9329 ( .A(n9984), .B(n9407), .ZN(n7508) );
  NOR2_X1 U9330 ( .A1(n7506), .A2(n10048), .ZN(n7507) );
  AOI21_X1 U9331 ( .B1(n7508), .B2(n10027), .A(n7507), .ZN(n10130) );
  XNOR2_X1 U9332 ( .A(n7509), .B(n7510), .ZN(n10134) );
  NAND2_X1 U9333 ( .A1(n10134), .A2(n10032), .ZN(n7514) );
  OAI22_X1 U9334 ( .A1(n10070), .A2(n7511), .B1(n9408), .B2(n10068), .ZN(n7512) );
  AOI21_X1 U9335 ( .B1(n10017), .B2(n9407), .A(n7512), .ZN(n7513) );
  OAI211_X1 U9336 ( .C1(n10130), .C2(n9581), .A(n7514), .B(n7513), .ZN(n7515)
         );
  AOI21_X1 U9337 ( .B1(n10132), .B2(n10070), .A(n7515), .ZN(n7516) );
  INV_X1 U9338 ( .A(n7516), .ZN(P1_U3284) );
  INV_X1 U9339 ( .A(n7517), .ZN(n7539) );
  OAI222_X1 U9340 ( .A1(n9286), .A2(n7539), .B1(P2_U3151), .B2(n7518), .C1(
        n9007), .C2(n9283), .ZN(P2_U3274) );
  XOR2_X1 U9341 ( .A(n7520), .B(n7519), .Z(n7538) );
  NAND2_X1 U9342 ( .A1(P2_U3151), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n8167) );
  OAI21_X1 U9343 ( .B1(n8615), .B2(n7521), .A(n8167), .ZN(n7528) );
  INV_X1 U9344 ( .A(n8547), .ZN(n7526) );
  NAND3_X1 U9345 ( .A1(n7524), .A2(n7523), .A3(n7522), .ZN(n7525) );
  AOI21_X1 U9346 ( .B1(n7526), .B2(n7525), .A(n8626), .ZN(n7527) );
  AOI211_X1 U9347 ( .C1(n8611), .C2(P2_ADDR_REG_12__SCAN_IN), .A(n7528), .B(
        n7527), .ZN(n7537) );
  INV_X1 U9348 ( .A(n7475), .ZN(n7532) );
  INV_X1 U9349 ( .A(n7529), .ZN(n7531) );
  NOR3_X1 U9350 ( .A1(n7532), .A2(n7531), .A3(n7530), .ZN(n7535) );
  INV_X1 U9351 ( .A(n7533), .ZN(n7534) );
  OAI21_X1 U9352 ( .B1(n7535), .B2(n7534), .A(n8641), .ZN(n7536) );
  OAI211_X1 U9353 ( .C1(n7538), .C2(n8645), .A(n7537), .B(n7536), .ZN(P2_U3194) );
  INV_X1 U9354 ( .A(n7541), .ZN(n7544) );
  OAI222_X1 U9355 ( .A1(n9283), .A2(n7543), .B1(n9281), .B2(n7544), .C1(n7542), 
        .C2(P2_U3151), .ZN(P2_U3273) );
  OAI222_X1 U9356 ( .A1(n7680), .A2(n7545), .B1(n9897), .B2(n7544), .C1(n7985), 
        .C2(P1_U3086), .ZN(P1_U3333) );
  NOR2_X1 U9357 ( .A1(n7547), .A2(n7546), .ZN(n7549) );
  AOI211_X1 U9358 ( .C1(n8920), .C2(n7550), .A(n7549), .B(n7548), .ZN(n7551)
         );
  MUX2_X1 U9359 ( .A(n9074), .B(n7551), .S(n10171), .Z(n7552) );
  OAI21_X1 U9360 ( .B1(n7553), .B2(n8784), .A(n7552), .ZN(P2_U3226) );
  XNOR2_X1 U9361 ( .A(n7554), .B(n7965), .ZN(n10137) );
  INV_X1 U9362 ( .A(n10137), .ZN(n7568) );
  OAI21_X1 U9363 ( .B1(n7965), .B2(n7556), .A(n7555), .ZN(n7557) );
  NAND2_X1 U9364 ( .A1(n7557), .A2(n10013), .ZN(n7559) );
  AOI22_X1 U9365 ( .A1(n10010), .A2(n9497), .B1(n10009), .B2(n9495), .ZN(n7558) );
  NAND2_X1 U9366 ( .A1(n7559), .A2(n7558), .ZN(n10143) );
  OAI21_X1 U9367 ( .B1(n7560), .B2(n10140), .A(n10027), .ZN(n7561) );
  OR2_X1 U9368 ( .A1(n7562), .A2(n7561), .ZN(n10138) );
  OAI22_X1 U9369 ( .A1(n10070), .A2(n7563), .B1(n9312), .B2(n10068), .ZN(n7564) );
  AOI21_X1 U9370 ( .B1(n9311), .B2(n10017), .A(n7564), .ZN(n7565) );
  OAI21_X1 U9371 ( .B1(n10138), .B2(n9581), .A(n7565), .ZN(n7566) );
  AOI21_X1 U9372 ( .B1(n10143), .B2(n10070), .A(n7566), .ZN(n7567) );
  OAI21_X1 U9373 ( .B1(n7568), .B2(n9780), .A(n7567), .ZN(P1_U3283) );
  INV_X1 U9374 ( .A(n7569), .ZN(n7577) );
  OAI22_X1 U9375 ( .A1(n10070), .A2(n7570), .B1(n7703), .B2(n10068), .ZN(n7571) );
  AOI21_X1 U9376 ( .B1(n7705), .B2(n10017), .A(n7571), .ZN(n7572) );
  OAI21_X1 U9377 ( .B1(n7573), .B2(n9581), .A(n7572), .ZN(n7574) );
  AOI21_X1 U9378 ( .B1(n7575), .B2(n10070), .A(n7574), .ZN(n7576) );
  OAI21_X1 U9379 ( .B1(n7577), .B2(n9780), .A(n7576), .ZN(P1_U3281) );
  INV_X1 U9380 ( .A(n7610), .ZN(n7579) );
  AOI21_X1 U9381 ( .B1(P2_DATAO_REG_23__SCAN_IN), .B2(n9894), .A(n8014), .ZN(
        n7578) );
  OAI21_X1 U9382 ( .B1(n7579), .B2(n9897), .A(n7578), .ZN(P1_U3332) );
  AND2_X1 U9383 ( .A1(n7581), .A2(n7580), .ZN(n9997) );
  INV_X1 U9384 ( .A(n7373), .ZN(n7582) );
  XNOR2_X1 U9385 ( .A(n9997), .B(n7582), .ZN(n10102) );
  OAI21_X1 U9386 ( .B1(n7373), .B2(n7583), .A(n7584), .ZN(n7588) );
  NAND2_X1 U9387 ( .A1(n9500), .A2(n10010), .ZN(n7585) );
  OAI21_X1 U9388 ( .B1(n7586), .B2(n10048), .A(n7585), .ZN(n7587) );
  AOI21_X1 U9389 ( .B1(n7588), .B2(n10013), .A(n7587), .ZN(n10108) );
  MUX2_X1 U9390 ( .A(n7589), .B(n10108), .S(n10070), .Z(n7594) );
  OAI211_X1 U9391 ( .C1(n10026), .C2(n10104), .A(n10027), .B(n10000), .ZN(
        n10103) );
  OAI22_X1 U9392 ( .A1(n10103), .A2(n9581), .B1(n7590), .B2(n10068), .ZN(n7591) );
  AOI21_X1 U9393 ( .B1(n10017), .B2(n7592), .A(n7591), .ZN(n7593) );
  OAI211_X1 U9394 ( .C1(n10102), .C2(n9780), .A(n7594), .B(n7593), .ZN(
        P1_U3288) );
  XNOR2_X1 U9395 ( .A(n7595), .B(n8493), .ZN(n7608) );
  INV_X1 U9396 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n9099) );
  XNOR2_X1 U9397 ( .A(n7598), .B(n7597), .ZN(n7599) );
  AOI222_X1 U9398 ( .A1(n8887), .A2(n7599), .B1(n8829), .B2(n8917), .C1(n8889), 
        .C2(n8890), .ZN(n7605) );
  MUX2_X1 U9399 ( .A(n9099), .B(n7605), .S(n10185), .Z(n7601) );
  NAND2_X1 U9400 ( .A1(n8349), .A2(n9247), .ZN(n7600) );
  OAI211_X1 U9401 ( .C1(n7608), .C2(n9255), .A(n7601), .B(n7600), .ZN(P2_U3423) );
  MUX2_X1 U9402 ( .A(n7602), .B(n7605), .S(n9003), .Z(n7604) );
  NAND2_X1 U9403 ( .A1(n8349), .A2(n8979), .ZN(n7603) );
  OAI211_X1 U9404 ( .C1(n8985), .C2(n7608), .A(n7604), .B(n7603), .ZN(P2_U3470) );
  MUX2_X1 U9405 ( .A(n9110), .B(n7605), .S(n10171), .Z(n7607) );
  AOI22_X1 U9406 ( .A1(n8349), .A2(n8921), .B1(n8920), .B2(n7634), .ZN(n7606)
         );
  OAI211_X1 U9407 ( .C1(n7608), .C2(n8855), .A(n7607), .B(n7606), .ZN(P2_U3222) );
  NAND2_X1 U9408 ( .A1(n7610), .A2(n7609), .ZN(n7612) );
  NAND2_X1 U9409 ( .A1(n7611), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8527) );
  OAI211_X1 U9410 ( .C1(n7613), .C2(n9283), .A(n7612), .B(n8527), .ZN(P2_U3272) );
  NAND2_X1 U9411 ( .A1(n7616), .A2(n7615), .ZN(n7650) );
  OAI21_X1 U9412 ( .B1(n7616), .B2(n7615), .A(n7650), .ZN(n7665) );
  NAND2_X1 U9413 ( .A1(n7617), .A2(n9430), .ZN(n7618) );
  NAND2_X1 U9414 ( .A1(n7618), .A2(n10027), .ZN(n7619) );
  OR2_X1 U9415 ( .A1(n7619), .A2(n7651), .ZN(n7662) );
  OAI22_X1 U9416 ( .A1(n10070), .A2(n7620), .B1(n9428), .B2(n10068), .ZN(n7621) );
  AOI21_X1 U9417 ( .B1(n9430), .B2(n10017), .A(n7621), .ZN(n7622) );
  OAI21_X1 U9418 ( .B1(n7662), .B2(n9581), .A(n7622), .ZN(n7628) );
  AND2_X1 U9419 ( .A1(n7623), .A2(n7827), .ZN(n7625) );
  OAI21_X1 U9420 ( .B1(n7625), .B2(n7969), .A(n7655), .ZN(n7626) );
  AOI222_X1 U9421 ( .A1(n10013), .A2(n7626), .B1(n9494), .B2(n10010), .C1(
        n9492), .C2(n10009), .ZN(n7663) );
  NOR2_X1 U9422 ( .A1(n7663), .A2(n4984), .ZN(n7627) );
  AOI211_X1 U9423 ( .C1(n10032), .C2(n7665), .A(n7628), .B(n7627), .ZN(n7629)
         );
  INV_X1 U9424 ( .A(n7629), .ZN(P1_U3280) );
  XNOR2_X1 U9425 ( .A(n8164), .B(n8163), .ZN(n7636) );
  NAND2_X1 U9426 ( .A1(n8283), .A2(n8889), .ZN(n7631) );
  OAI211_X1 U9427 ( .C1(n8355), .C2(n8285), .A(n7631), .B(n7630), .ZN(n7633)
         );
  NOR2_X1 U9428 ( .A1(n8340), .A2(n8291), .ZN(n7632) );
  AOI211_X1 U9429 ( .C1(n7634), .C2(n8288), .A(n7633), .B(n7632), .ZN(n7635)
         );
  OAI21_X1 U9430 ( .B1(n7636), .B2(n8279), .A(n7635), .ZN(P2_U3176) );
  INV_X1 U9431 ( .A(n10053), .ZN(n9981) );
  XNOR2_X1 U9432 ( .A(n7960), .B(n10035), .ZN(n7643) );
  INV_X1 U9433 ( .A(n7643), .ZN(n10083) );
  INV_X1 U9434 ( .A(n7960), .ZN(n10036) );
  XNOR2_X1 U9435 ( .A(n10036), .B(n7637), .ZN(n7639) );
  AOI22_X1 U9436 ( .A1(n10009), .A2(n7352), .B1(n10010), .B2(n7346), .ZN(n7638) );
  OAI21_X1 U9437 ( .B1(n7639), .B2(n10047), .A(n7638), .ZN(n7640) );
  AOI21_X1 U9438 ( .B1(n9981), .B2(n10083), .A(n7640), .ZN(n10080) );
  INV_X1 U9439 ( .A(n7641), .ZN(n10040) );
  OAI211_X1 U9440 ( .C1(n4405), .C2(n7642), .A(n10027), .B(n10040), .ZN(n10079) );
  OAI22_X1 U9441 ( .A1(n9581), .A2(n10079), .B1(n9502), .B2(n10068), .ZN(n7646) );
  OAI22_X1 U9442 ( .A1(n4405), .A2(n9766), .B1(n7644), .B2(n7643), .ZN(n7645)
         );
  AOI211_X1 U9443 ( .C1(P1_REG2_REG_1__SCAN_IN), .C2(n4984), .A(n7646), .B(
        n7645), .ZN(n7647) );
  OAI21_X1 U9444 ( .B1(n4984), .B2(n10080), .A(n7647), .ZN(P1_U3292) );
  NAND2_X1 U9445 ( .A1(n9857), .A2(n9425), .ZN(n7837) );
  NAND2_X1 U9446 ( .A1(n7929), .A2(n7837), .ZN(n7970) );
  INV_X1 U9447 ( .A(n9430), .ZN(n7648) );
  NAND2_X1 U9448 ( .A1(n7648), .A2(n7700), .ZN(n7649) );
  NAND2_X1 U9449 ( .A1(n7650), .A2(n7649), .ZN(n7684) );
  XOR2_X1 U9450 ( .A(n7970), .B(n7684), .Z(n9862) );
  INV_X1 U9451 ( .A(n7651), .ZN(n7652) );
  AOI211_X1 U9452 ( .C1(n9857), .C2(n7652), .A(n10039), .B(n7691), .ZN(n9856)
         );
  INV_X1 U9453 ( .A(n9294), .ZN(n7653) );
  AOI22_X1 U9454 ( .A1(n4984), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n7653), .B2(
        n10015), .ZN(n7654) );
  OAI21_X1 U9455 ( .B1(n7685), .B2(n9766), .A(n7654), .ZN(n7660) );
  AOI211_X1 U9456 ( .C1(n7656), .C2(n7970), .A(n10047), .B(n7687), .ZN(n7658)
         );
  OAI22_X1 U9457 ( .A1(n10050), .A2(n7700), .B1(n9291), .B2(n10048), .ZN(n7657) );
  NOR2_X1 U9458 ( .A1(n7658), .A2(n7657), .ZN(n9860) );
  NOR2_X1 U9459 ( .A1(n9860), .A2(n4984), .ZN(n7659) );
  AOI211_X1 U9460 ( .C1(n9856), .C2(n10031), .A(n7660), .B(n7659), .ZN(n7661)
         );
  OAI21_X1 U9461 ( .B1(n9862), .B2(n9780), .A(n7661), .ZN(P1_U3279) );
  OAI211_X1 U9462 ( .C1(n7648), .C2(n10139), .A(n7663), .B(n7662), .ZN(n7664)
         );
  AOI21_X1 U9463 ( .B1(n10136), .B2(n7665), .A(n7664), .ZN(n7668) );
  NAND2_X1 U9464 ( .A1(n10144), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n7666) );
  OAI21_X1 U9465 ( .B1(n7668), .B2(n10144), .A(n7666), .ZN(P1_U3492) );
  NAND2_X1 U9466 ( .A1(n10160), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n7667) );
  OAI21_X1 U9467 ( .B1(n7668), .B2(n10160), .A(n7667), .ZN(P1_U3535) );
  INV_X1 U9468 ( .A(n7669), .ZN(n7682) );
  OAI222_X1 U9469 ( .A1(n9281), .A2(n7682), .B1(P2_U3151), .B2(n5313), .C1(
        n7670), .C2(n9283), .ZN(P2_U3271) );
  XNOR2_X1 U9470 ( .A(n9401), .B(n9402), .ZN(n7671) );
  NOR2_X1 U9471 ( .A1(n7671), .A2(n7672), .ZN(n9400) );
  AOI21_X1 U9472 ( .B1(n7672), .B2(n7671), .A(n9400), .ZN(n7679) );
  AOI22_X1 U9473 ( .A1(n9444), .A2(n10122), .B1(n9451), .B2(n9497), .ZN(n7678)
         );
  INV_X1 U9474 ( .A(n7673), .ZN(n7674) );
  AOI21_X1 U9475 ( .B1(n9482), .B2(n9992), .A(n7674), .ZN(n7675) );
  OAI21_X1 U9476 ( .B1(n9479), .B2(n9982), .A(n7675), .ZN(n7676) );
  INV_X1 U9477 ( .A(n7676), .ZN(n7677) );
  OAI211_X1 U9478 ( .C1(n7679), .C2(n9458), .A(n7678), .B(n7677), .ZN(P1_U3221) );
  OAI222_X1 U9479 ( .A1(P1_U3086), .A2(n7683), .B1(n9897), .B2(n7682), .C1(
        n7681), .C2(n7680), .ZN(P1_U3331) );
  INV_X1 U9480 ( .A(n9857), .ZN(n7685) );
  NAND2_X1 U9481 ( .A1(n7685), .A2(n9425), .ZN(n7686) );
  XNOR2_X1 U9482 ( .A(n9852), .B(n9491), .ZN(n7972) );
  XNOR2_X1 U9483 ( .A(n7715), .B(n7972), .ZN(n9855) );
  OAI21_X1 U9484 ( .B1(n7688), .B2(n7972), .A(n7716), .ZN(n7689) );
  AOI222_X1 U9485 ( .A1(n10013), .A2(n7689), .B1(n9771), .B2(n10009), .C1(
        n9492), .C2(n10010), .ZN(n9854) );
  OAI22_X1 U9486 ( .A1(n10070), .A2(n9913), .B1(n9478), .B2(n10068), .ZN(n7690) );
  AOI21_X1 U9487 ( .B1(n9852), .B2(n10017), .A(n7690), .ZN(n7694) );
  OR2_X1 U9488 ( .A1(n7691), .A2(n9486), .ZN(n7692) );
  AND3_X1 U9489 ( .A1(n7719), .A2(n7692), .A3(n10027), .ZN(n9851) );
  NAND2_X1 U9490 ( .A1(n9851), .A2(n10031), .ZN(n7693) );
  OAI211_X1 U9491 ( .C1(n9854), .C2(n4984), .A(n7694), .B(n7693), .ZN(n7695)
         );
  INV_X1 U9492 ( .A(n7695), .ZN(n7696) );
  OAI21_X1 U9493 ( .B1(n9780), .B2(n9855), .A(n7696), .ZN(P1_U3278) );
  XOR2_X1 U9494 ( .A(n7697), .B(n7698), .Z(n7707) );
  OAI21_X1 U9495 ( .B1(n9477), .B2(n7700), .A(n7699), .ZN(n7701) );
  AOI21_X1 U9496 ( .B1(n9482), .B2(n9495), .A(n7701), .ZN(n7702) );
  OAI21_X1 U9497 ( .B1(n9479), .B2(n7703), .A(n7702), .ZN(n7704) );
  AOI21_X1 U9498 ( .B1(n7705), .B2(n9444), .A(n7704), .ZN(n7706) );
  OAI21_X1 U9499 ( .B1(n7707), .B2(n9458), .A(n7706), .ZN(P1_U3224) );
  INV_X1 U9500 ( .A(n7708), .ZN(n7713) );
  AOI22_X1 U9501 ( .A1(n7709), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(n9894), .ZN(n7710) );
  OAI21_X1 U9502 ( .B1(n7713), .B2(n9897), .A(n7710), .ZN(P1_U3330) );
  OAI222_X1 U9503 ( .A1(n9281), .A2(n7713), .B1(P2_U3151), .B2(n7712), .C1(
        n7711), .C2(n9283), .ZN(P2_U3270) );
  OR2_X1 U9504 ( .A1(n9848), .A2(n9476), .ZN(n7842) );
  NAND2_X1 U9505 ( .A1(n9848), .A2(n9476), .ZN(n7991) );
  XNOR2_X1 U9506 ( .A(n8058), .B(n8057), .ZN(n9850) );
  NAND2_X1 U9507 ( .A1(n9852), .A2(n9291), .ZN(n7786) );
  NAND2_X1 U9508 ( .A1(n7716), .A2(n7786), .ZN(n7993) );
  XOR2_X1 U9509 ( .A(n8057), .B(n7717), .Z(n7718) );
  OAI222_X1 U9510 ( .A1(n10048), .A2(n9453), .B1(n10050), .B2(n9291), .C1(
        n7718), .C2(n10047), .ZN(n9846) );
  AOI21_X1 U9511 ( .B1(n9848), .B2(n7719), .A(n10039), .ZN(n7720) );
  AND2_X1 U9512 ( .A1(n7720), .A2(n9761), .ZN(n9847) );
  NAND2_X1 U9513 ( .A1(n9847), .A2(n10031), .ZN(n7724) );
  OAI22_X1 U9514 ( .A1(n10070), .A2(n7721), .B1(n9379), .B2(n10068), .ZN(n7722) );
  AOI21_X1 U9515 ( .B1(n9848), .B2(n10017), .A(n7722), .ZN(n7723) );
  NAND2_X1 U9516 ( .A1(n7724), .A2(n7723), .ZN(n7725) );
  AOI21_X1 U9517 ( .B1(n9846), .B2(n10070), .A(n7725), .ZN(n7726) );
  OAI21_X1 U9518 ( .B1(n9850), .B2(n9780), .A(n7726), .ZN(P1_U3277) );
  INV_X1 U9519 ( .A(n7727), .ZN(n7732) );
  AOI22_X1 U9520 ( .A1(n7728), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n9894), .ZN(n7729) );
  OAI21_X1 U9521 ( .B1(n7732), .B2(n9897), .A(n7729), .ZN(P1_U3329) );
  OAI222_X1 U9522 ( .A1(n9286), .A2(n7732), .B1(P2_U3151), .B2(n7731), .C1(
        n7730), .C2(n9283), .ZN(P2_U3269) );
  INV_X1 U9523 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n10196) );
  INV_X1 U9524 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n9952) );
  INV_X1 U9525 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n7733) );
  AOI22_X1 U9526 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .B1(n9952), .B2(n7733), .ZN(n10200) );
  INV_X1 U9527 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n9937) );
  INV_X1 U9528 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n7734) );
  AOI22_X1 U9529 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .B1(n9937), .B2(n7734), .ZN(n10203) );
  NOR2_X1 U9530 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n7735) );
  AOI21_X1 U9531 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n7735), .ZN(n10206) );
  NOR2_X1 U9532 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n7736) );
  AOI21_X1 U9533 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n7736), .ZN(n10209) );
  NOR2_X1 U9534 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n7737) );
  AOI21_X1 U9535 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n7737), .ZN(n10212) );
  NOR2_X1 U9536 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n7738) );
  AOI21_X1 U9537 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n7738), .ZN(n10215) );
  NOR2_X1 U9538 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n7739) );
  AOI21_X1 U9539 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n7739), .ZN(n10218) );
  NOR2_X1 U9540 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n7740) );
  AOI21_X1 U9541 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n7740), .ZN(n10221) );
  NOR2_X1 U9542 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n7741) );
  AOI21_X1 U9543 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(P2_ADDR_REG_9__SCAN_IN), 
        .A(n7741), .ZN(n10230) );
  NOR2_X1 U9544 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n7742) );
  AOI21_X1 U9545 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(P2_ADDR_REG_8__SCAN_IN), 
        .A(n7742), .ZN(n10236) );
  NOR2_X1 U9546 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n7743) );
  AOI21_X1 U9547 ( .B1(P1_ADDR_REG_7__SCAN_IN), .B2(P2_ADDR_REG_7__SCAN_IN), 
        .A(n7743), .ZN(n10233) );
  NOR2_X1 U9548 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(P2_ADDR_REG_6__SCAN_IN), 
        .ZN(n7744) );
  AOI21_X1 U9549 ( .B1(P2_ADDR_REG_6__SCAN_IN), .B2(P1_ADDR_REG_6__SCAN_IN), 
        .A(n7744), .ZN(n10224) );
  NOR2_X1 U9550 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n7745) );
  AOI21_X1 U9551 ( .B1(P1_ADDR_REG_5__SCAN_IN), .B2(P2_ADDR_REG_5__SCAN_IN), 
        .A(n7745), .ZN(n10227) );
  AND2_X1 U9552 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .ZN(n7746) );
  NOR2_X1 U9553 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(n7746), .ZN(n10190) );
  INV_X1 U9554 ( .A(n10190), .ZN(n10191) );
  INV_X1 U9555 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10193) );
  NAND3_X1 U9556 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(P1_ADDR_REG_0__SCAN_IN), 
        .A3(P2_ADDR_REG_0__SCAN_IN), .ZN(n10192) );
  NAND2_X1 U9557 ( .A1(n10193), .A2(n10192), .ZN(n10189) );
  NAND2_X1 U9558 ( .A1(n10191), .A2(n10189), .ZN(n10239) );
  NAND2_X1 U9559 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n7747) );
  OAI21_X1 U9560 ( .B1(P1_ADDR_REG_2__SCAN_IN), .B2(P2_ADDR_REG_2__SCAN_IN), 
        .A(n7747), .ZN(n10238) );
  NOR2_X1 U9561 ( .A1(n10239), .A2(n10238), .ZN(n10237) );
  AOI21_X1 U9562 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(P1_ADDR_REG_2__SCAN_IN), 
        .A(n10237), .ZN(n10242) );
  NAND2_X1 U9563 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n7748) );
  OAI21_X1 U9564 ( .B1(P1_ADDR_REG_3__SCAN_IN), .B2(P2_ADDR_REG_3__SCAN_IN), 
        .A(n7748), .ZN(n10241) );
  NOR2_X1 U9565 ( .A1(n10242), .A2(n10241), .ZN(n10240) );
  AOI21_X1 U9566 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(P1_ADDR_REG_3__SCAN_IN), 
        .A(n10240), .ZN(n10245) );
  NOR2_X1 U9567 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n7749) );
  AOI21_X1 U9568 ( .B1(P2_ADDR_REG_4__SCAN_IN), .B2(P1_ADDR_REG_4__SCAN_IN), 
        .A(n7749), .ZN(n10244) );
  NAND2_X1 U9569 ( .A1(n10245), .A2(n10244), .ZN(n10243) );
  OAI21_X1 U9570 ( .B1(P1_ADDR_REG_4__SCAN_IN), .B2(P2_ADDR_REG_4__SCAN_IN), 
        .A(n10243), .ZN(n10226) );
  NAND2_X1 U9571 ( .A1(n10227), .A2(n10226), .ZN(n10225) );
  OAI21_X1 U9572 ( .B1(P2_ADDR_REG_5__SCAN_IN), .B2(P1_ADDR_REG_5__SCAN_IN), 
        .A(n10225), .ZN(n10223) );
  NAND2_X1 U9573 ( .A1(n10224), .A2(n10223), .ZN(n10222) );
  OAI21_X1 U9574 ( .B1(P1_ADDR_REG_6__SCAN_IN), .B2(P2_ADDR_REG_6__SCAN_IN), 
        .A(n10222), .ZN(n10232) );
  NAND2_X1 U9575 ( .A1(n10233), .A2(n10232), .ZN(n10231) );
  OAI21_X1 U9576 ( .B1(P2_ADDR_REG_7__SCAN_IN), .B2(P1_ADDR_REG_7__SCAN_IN), 
        .A(n10231), .ZN(n10235) );
  NAND2_X1 U9577 ( .A1(n10236), .A2(n10235), .ZN(n10234) );
  OAI21_X1 U9578 ( .B1(P2_ADDR_REG_8__SCAN_IN), .B2(P1_ADDR_REG_8__SCAN_IN), 
        .A(n10234), .ZN(n10229) );
  NAND2_X1 U9579 ( .A1(n10230), .A2(n10229), .ZN(n10228) );
  OAI21_X1 U9580 ( .B1(P2_ADDR_REG_9__SCAN_IN), .B2(P1_ADDR_REG_9__SCAN_IN), 
        .A(n10228), .ZN(n10220) );
  NAND2_X1 U9581 ( .A1(n10221), .A2(n10220), .ZN(n10219) );
  OAI21_X1 U9582 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n10219), .ZN(n10217) );
  NAND2_X1 U9583 ( .A1(n10218), .A2(n10217), .ZN(n10216) );
  OAI21_X1 U9584 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n10216), .ZN(n10214) );
  NAND2_X1 U9585 ( .A1(n10215), .A2(n10214), .ZN(n10213) );
  OAI21_X1 U9586 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10213), .ZN(n10211) );
  NAND2_X1 U9587 ( .A1(n10212), .A2(n10211), .ZN(n10210) );
  OAI21_X1 U9588 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n10210), .ZN(n10208) );
  NAND2_X1 U9589 ( .A1(n10209), .A2(n10208), .ZN(n10207) );
  OAI21_X1 U9590 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10207), .ZN(n10205) );
  NAND2_X1 U9591 ( .A1(n10206), .A2(n10205), .ZN(n10204) );
  OAI21_X1 U9592 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n10204), .ZN(n10202) );
  NAND2_X1 U9593 ( .A1(n10203), .A2(n10202), .ZN(n10201) );
  OAI21_X1 U9594 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n10201), .ZN(n10199) );
  NAND2_X1 U9595 ( .A1(n10200), .A2(n10199), .ZN(n10198) );
  OAI21_X1 U9596 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10198), .ZN(n10195) );
  NAND2_X1 U9597 ( .A1(n10196), .A2(n10195), .ZN(n7750) );
  NOR2_X1 U9598 ( .A1(n10196), .A2(n10195), .ZN(n10194) );
  AOI21_X1 U9599 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(n7750), .A(n10194), .ZN(
        n7752) );
  XNOR2_X1 U9600 ( .A(n4489), .B(P1_ADDR_REG_19__SCAN_IN), .ZN(n7751) );
  XNOR2_X1 U9601 ( .A(n7752), .B(n7751), .ZN(ADD_1068_U4) );
  INV_X1 U9602 ( .A(n7753), .ZN(n7755) );
  NAND2_X1 U9603 ( .A1(n7770), .A2(n7769), .ZN(n9300) );
  NAND2_X1 U9604 ( .A1(n7753), .A2(n7756), .ZN(n9299) );
  INV_X1 U9605 ( .A(n7757), .ZN(n7758) );
  OR2_X1 U9606 ( .A1(n7758), .A2(n7760), .ZN(n9298) );
  NOR3_X1 U9607 ( .A1(n9302), .A2(n7760), .A3(n4698), .ZN(n7762) );
  OAI21_X1 U9608 ( .B1(n7762), .B2(n7761), .A(n9474), .ZN(n7767) );
  INV_X1 U9609 ( .A(n7763), .ZN(n9661) );
  INV_X1 U9610 ( .A(n9687), .ZN(n8067) );
  AOI22_X1 U9611 ( .A1(n9657), .A2(n9451), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3086), .ZN(n7764) );
  OAI21_X1 U9612 ( .B1(n8067), .B2(n9454), .A(n7764), .ZN(n7765) );
  AOI21_X1 U9613 ( .B1(n9661), .B2(n9468), .A(n7765), .ZN(n7766) );
  INV_X1 U9614 ( .A(n9299), .ZN(n7768) );
  NOR2_X1 U9615 ( .A1(n9300), .A2(n7768), .ZN(n7772) );
  AOI21_X1 U9616 ( .B1(n7770), .B2(n9299), .A(n7769), .ZN(n7771) );
  OAI21_X1 U9617 ( .B1(n7772), .B2(n7771), .A(n9474), .ZN(n7776) );
  NOR2_X1 U9618 ( .A1(n9479), .A2(n9691), .ZN(n7774) );
  OAI22_X1 U9619 ( .A1(n8067), .A2(n9477), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9038), .ZN(n7773) );
  AOI211_X1 U9620 ( .C1(n9482), .C2(n9686), .A(n7774), .B(n7773), .ZN(n7775)
         );
  OAI211_X1 U9621 ( .C1(n9695), .C2(n9485), .A(n7776), .B(n7775), .ZN(P1_U3235) );
  NOR2_X1 U9622 ( .A1(n4984), .A2(n7777), .ZN(n9578) );
  NOR2_X1 U9623 ( .A1(n7945), .A2(n9766), .ZN(n7778) );
  AOI211_X1 U9624 ( .C1(n4984), .C2(P1_REG2_REG_30__SCAN_IN), .A(n9578), .B(
        n7778), .ZN(n7779) );
  OAI21_X1 U9625 ( .B1(n9581), .B2(n7780), .A(n7779), .ZN(P1_U3264) );
  NOR2_X1 U9626 ( .A1(n9800), .A2(n8074), .ZN(n7888) );
  NAND2_X1 U9627 ( .A1(n9824), .A2(n8062), .ZN(n7854) );
  INV_X1 U9628 ( .A(n9490), .ZN(n9740) );
  NAND2_X1 U9629 ( .A1(n9829), .A2(n9740), .ZN(n7782) );
  AND2_X1 U9630 ( .A1(n7854), .A2(n7782), .ZN(n7890) );
  INV_X1 U9631 ( .A(n7889), .ZN(n7853) );
  OR2_X1 U9632 ( .A1(n9829), .A2(n9740), .ZN(n9705) );
  MUX2_X1 U9633 ( .A(n7890), .B(n8040), .S(n7877), .Z(n7852) );
  NAND3_X1 U9634 ( .A1(n9705), .A2(n9731), .A3(n7956), .ZN(n7781) );
  OAI21_X1 U9635 ( .B1(n9717), .B2(n7882), .A(n7781), .ZN(n7783) );
  NAND2_X1 U9636 ( .A1(n7783), .A2(n7782), .ZN(n7785) );
  NAND3_X1 U9637 ( .A1(n9705), .A2(n7882), .A3(n7956), .ZN(n7784) );
  NAND2_X1 U9638 ( .A1(n7785), .A2(n7784), .ZN(n7851) );
  NAND2_X1 U9639 ( .A1(n7991), .A2(n7786), .ZN(n7841) );
  INV_X1 U9640 ( .A(n7837), .ZN(n7787) );
  OR2_X1 U9641 ( .A1(n7841), .A2(n7787), .ZN(n7900) );
  NAND3_X1 U9642 ( .A1(n7583), .A2(n7882), .A3(n7798), .ZN(n7802) );
  INV_X1 U9643 ( .A(n7798), .ZN(n7789) );
  NAND3_X1 U9644 ( .A1(n7789), .A2(n7794), .A3(n7877), .ZN(n7791) );
  OAI211_X1 U9645 ( .C1(n7794), .C2(n7877), .A(n7791), .B(n7790), .ZN(n7792)
         );
  INV_X1 U9646 ( .A(n7792), .ZN(n7801) );
  INV_X1 U9647 ( .A(n7793), .ZN(n7796) );
  NAND4_X1 U9648 ( .A1(n7794), .A2(n7913), .A3(n7912), .A4(n7877), .ZN(n7795)
         );
  INV_X1 U9649 ( .A(n7912), .ZN(n7797) );
  NAND3_X1 U9650 ( .A1(n7798), .A2(n7797), .A3(n7882), .ZN(n7799) );
  NAND4_X1 U9651 ( .A1(n7801), .A2(n7802), .A3(n7800), .A4(n7799), .ZN(n7806)
         );
  MUX2_X1 U9652 ( .A(n7804), .B(n7803), .S(n7877), .Z(n7805) );
  NAND2_X1 U9653 ( .A1(n7806), .A2(n7805), .ZN(n7812) );
  NAND2_X1 U9654 ( .A1(n7813), .A2(n7807), .ZN(n7809) );
  MUX2_X1 U9655 ( .A(n7809), .B(n7808), .S(n7877), .Z(n7810) );
  INV_X1 U9656 ( .A(n7810), .ZN(n7811) );
  NAND2_X1 U9657 ( .A1(n7812), .A2(n7811), .ZN(n7819) );
  NAND3_X1 U9658 ( .A1(n7819), .A2(n7921), .A3(n7813), .ZN(n7816) );
  INV_X1 U9659 ( .A(n7823), .ZN(n7814) );
  NAND2_X1 U9660 ( .A1(n7921), .A2(n7814), .ZN(n7815) );
  AND3_X1 U9661 ( .A1(n7827), .A2(n7822), .A3(n7815), .ZN(n7901) );
  NAND2_X1 U9662 ( .A1(n7816), .A2(n7901), .ZN(n7817) );
  NAND2_X1 U9663 ( .A1(n7817), .A2(n7923), .ZN(n7829) );
  NAND2_X1 U9664 ( .A1(n7819), .A2(n7818), .ZN(n7821) );
  NAND2_X1 U9665 ( .A1(n7821), .A2(n7820), .ZN(n7824) );
  INV_X1 U9666 ( .A(n7928), .ZN(n7838) );
  OR2_X1 U9667 ( .A1(n7970), .A2(n7838), .ZN(n7830) );
  AOI21_X1 U9668 ( .B1(n7836), .B2(n7924), .A(n7830), .ZN(n7832) );
  AND2_X1 U9669 ( .A1(n9486), .A2(n9491), .ZN(n7839) );
  NAND2_X1 U9670 ( .A1(n7991), .A2(n7839), .ZN(n7831) );
  AND2_X1 U9671 ( .A1(n7831), .A2(n7842), .ZN(n7930) );
  NAND2_X1 U9672 ( .A1(n9843), .A2(n9453), .ZN(n7957) );
  OR2_X1 U9673 ( .A1(n7834), .A2(n9739), .ZN(n7955) );
  NAND2_X1 U9674 ( .A1(n9834), .A2(n9717), .ZN(n7997) );
  NAND2_X1 U9675 ( .A1(n7834), .A2(n9739), .ZN(n7996) );
  INV_X1 U9676 ( .A(n7839), .ZN(n7840) );
  INV_X1 U9677 ( .A(n7841), .ZN(n7844) );
  INV_X1 U9678 ( .A(n7842), .ZN(n7843) );
  AOI21_X1 U9679 ( .B1(n7845), .B2(n7844), .A(n7843), .ZN(n7850) );
  NAND2_X1 U9680 ( .A1(n7996), .A2(n7957), .ZN(n7934) );
  NAND2_X1 U9681 ( .A1(n7994), .A2(n9739), .ZN(n7848) );
  INV_X1 U9682 ( .A(n9453), .ZN(n9755) );
  NAND3_X1 U9683 ( .A1(n9767), .A2(n9772), .A3(n9755), .ZN(n7846) );
  NAND2_X1 U9684 ( .A1(n7846), .A2(n7877), .ZN(n7847) );
  AOI21_X1 U9685 ( .B1(n9747), .B2(n7848), .A(n7847), .ZN(n7849) );
  MUX2_X1 U9686 ( .A(n7854), .B(n7853), .S(n7882), .Z(n7855) );
  NAND2_X1 U9687 ( .A1(n7858), .A2(n8042), .ZN(n9670) );
  INV_X1 U9688 ( .A(n9670), .ZN(n9668) );
  XNOR2_X1 U9689 ( .A(n9819), .B(n9489), .ZN(n9684) );
  NAND3_X1 U9690 ( .A1(n7856), .A2(n9668), .A3(n9684), .ZN(n7862) );
  NAND2_X1 U9691 ( .A1(n9819), .A2(n9709), .ZN(n7857) );
  NAND2_X1 U9692 ( .A1(n8042), .A2(n7857), .ZN(n7891) );
  NAND2_X1 U9693 ( .A1(n7891), .A2(n7858), .ZN(n7860) );
  NAND2_X1 U9694 ( .A1(n9695), .A2(n9489), .ZN(n8041) );
  NAND2_X1 U9695 ( .A1(n7858), .A2(n8041), .ZN(n7859) );
  NAND2_X1 U9696 ( .A1(n7859), .A2(n8042), .ZN(n7893) );
  MUX2_X1 U9697 ( .A(n7860), .B(n7893), .S(n7882), .Z(n7861) );
  NAND2_X1 U9698 ( .A1(n7862), .A2(n7861), .ZN(n7863) );
  NAND2_X1 U9699 ( .A1(n9809), .A2(n9673), .ZN(n7894) );
  NAND2_X1 U9700 ( .A1(n7863), .A2(n9655), .ZN(n7865) );
  MUX2_X1 U9701 ( .A(n8044), .B(n7894), .S(n7877), .Z(n7864) );
  NAND2_X1 U9702 ( .A1(n9804), .A2(n9630), .ZN(n7954) );
  NAND2_X1 U9703 ( .A1(n7954), .A2(n7882), .ZN(n7866) );
  AND2_X1 U9704 ( .A1(n9800), .A2(n8074), .ZN(n8046) );
  NAND2_X1 U9705 ( .A1(n9788), .A2(n9607), .ZN(n7978) );
  INV_X1 U9706 ( .A(n7952), .ZN(n7867) );
  INV_X1 U9707 ( .A(n7954), .ZN(n7869) );
  INV_X1 U9708 ( .A(n8048), .ZN(n7871) );
  NOR2_X1 U9709 ( .A1(n7872), .A2(n7871), .ZN(n7874) );
  INV_X1 U9710 ( .A(n7953), .ZN(n8047) );
  OAI21_X1 U9711 ( .B1(n7898), .B2(n8047), .A(n8048), .ZN(n7873) );
  NAND2_X1 U9712 ( .A1(n8085), .A2(n9591), .ZN(n7943) );
  MUX2_X1 U9713 ( .A(n7943), .B(n7940), .S(n7877), .Z(n7875) );
  INV_X1 U9714 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n9082) );
  NAND2_X1 U9715 ( .A1(n7878), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n7880) );
  NAND2_X1 U9716 ( .A1(n6486), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n7879) );
  OAI211_X1 U9717 ( .C1(n7881), .C2(n9082), .A(n7880), .B(n7879), .ZN(n9487)
         );
  OAI21_X1 U9718 ( .B1(n7946), .B2(n9487), .A(n8010), .ZN(n7884) );
  NOR2_X1 U9719 ( .A1(n7953), .A2(n7888), .ZN(n7999) );
  INV_X1 U9720 ( .A(n7894), .ZN(n7892) );
  NOR2_X1 U9721 ( .A1(n7890), .A2(n7889), .ZN(n8039) );
  NOR3_X1 U9722 ( .A1(n7892), .A2(n8039), .A3(n7891), .ZN(n7897) );
  NAND2_X1 U9723 ( .A1(n7893), .A2(n8044), .ZN(n7895) );
  NAND2_X1 U9724 ( .A1(n7895), .A2(n7894), .ZN(n7896) );
  NAND2_X1 U9725 ( .A1(n8045), .A2(n7896), .ZN(n7936) );
  OAI21_X1 U9726 ( .B1(n7897), .B2(n7936), .A(n7954), .ZN(n7899) );
  INV_X1 U9727 ( .A(n7900), .ZN(n7933) );
  INV_X1 U9728 ( .A(n7901), .ZN(n7926) );
  OAI211_X1 U9729 ( .C1(n4441), .C2(n7903), .A(n5896), .B(n7902), .ZN(n7904)
         );
  INV_X1 U9730 ( .A(n7904), .ZN(n7907) );
  OAI211_X1 U9731 ( .C1(n7908), .C2(n7907), .A(n7906), .B(n7905), .ZN(n7909)
         );
  NAND2_X1 U9732 ( .A1(n7909), .A2(n10007), .ZN(n7911) );
  NAND2_X1 U9733 ( .A1(n7911), .A2(n7910), .ZN(n7917) );
  AND2_X1 U9734 ( .A1(n7913), .A2(n7912), .ZN(n7916) );
  INV_X1 U9735 ( .A(n7914), .ZN(n7915) );
  AOI21_X1 U9736 ( .B1(n7917), .B2(n7916), .A(n7915), .ZN(n7920) );
  OAI21_X1 U9737 ( .B1(n7920), .B2(n7919), .A(n7918), .ZN(n7922) );
  AND2_X1 U9738 ( .A1(n7922), .A2(n7921), .ZN(n7925) );
  OAI211_X1 U9739 ( .C1(n7926), .C2(n7925), .A(n7924), .B(n7923), .ZN(n7927)
         );
  NAND3_X1 U9740 ( .A1(n7929), .A2(n7928), .A3(n7927), .ZN(n7932) );
  INV_X1 U9741 ( .A(n7994), .ZN(n9749) );
  INV_X1 U9742 ( .A(n7930), .ZN(n7931) );
  AOI211_X1 U9743 ( .C1(n7933), .C2(n7932), .A(n9749), .B(n7931), .ZN(n7935)
         );
  OAI211_X1 U9744 ( .C1(n7935), .C2(n7934), .A(n7955), .B(n7956), .ZN(n7938)
         );
  INV_X1 U9745 ( .A(n7936), .ZN(n7937) );
  NAND2_X1 U9746 ( .A1(n7937), .A2(n8040), .ZN(n7990) );
  AOI21_X1 U9747 ( .B1(n7997), .B2(n7938), .A(n7990), .ZN(n7939) );
  OAI21_X1 U9748 ( .B1(n8046), .B2(n7939), .A(n7999), .ZN(n7941) );
  NAND2_X1 U9749 ( .A1(n7940), .A2(n8048), .ZN(n8003) );
  AOI21_X1 U9750 ( .B1(n8000), .B2(n7941), .A(n8003), .ZN(n7944) );
  INV_X1 U9751 ( .A(n9487), .ZN(n7942) );
  NAND2_X1 U9752 ( .A1(n8004), .A2(n7942), .ZN(n7951) );
  NAND2_X1 U9753 ( .A1(n7951), .A2(n7943), .ZN(n8008) );
  NOR2_X1 U9754 ( .A1(n7944), .A2(n8008), .ZN(n7947) );
  INV_X1 U9755 ( .A(n8016), .ZN(n7984) );
  NAND2_X1 U9756 ( .A1(n7945), .A2(n9487), .ZN(n8009) );
  NAND2_X1 U9757 ( .A1(n7984), .A2(n8009), .ZN(n7950) );
  INV_X1 U9758 ( .A(n8018), .ZN(n7981) );
  OAI21_X1 U9759 ( .B1(n7947), .B2(n7950), .A(n7981), .ZN(n7948) );
  MUX2_X1 U9760 ( .A(n6478), .B(n7949), .S(n7948), .Z(n8030) );
  INV_X1 U9761 ( .A(n8030), .ZN(n8034) );
  INV_X1 U9762 ( .A(n7950), .ZN(n7983) );
  INV_X1 U9763 ( .A(n7951), .ZN(n7980) );
  INV_X1 U9764 ( .A(n9727), .ZN(n9736) );
  XNOR2_X1 U9765 ( .A(n9829), .B(n9490), .ZN(n9712) );
  INV_X1 U9766 ( .A(n7958), .ZN(n7966) );
  INV_X1 U9767 ( .A(n7959), .ZN(n7964) );
  NOR2_X1 U9768 ( .A1(n10064), .A2(n5896), .ZN(n7961) );
  NAND4_X1 U9769 ( .A1(n7961), .A2(n7373), .A3(n7345), .A4(n7960), .ZN(n7962)
         );
  NOR4_X1 U9770 ( .A1(n7962), .A2(n9999), .A3(n10045), .A4(n10024), .ZN(n7963)
         );
  AND4_X1 U9771 ( .A1(n7966), .A2(n7965), .A3(n7964), .A4(n7963), .ZN(n7967)
         );
  NAND4_X1 U9772 ( .A1(n7969), .A2(n4983), .A3(n7968), .A4(n7967), .ZN(n7971)
         );
  NOR2_X1 U9773 ( .A1(n7971), .A2(n7970), .ZN(n7973) );
  AND4_X1 U9774 ( .A1(n8057), .A2(n9769), .A3(n7973), .A4(n7972), .ZN(n7974)
         );
  NAND4_X1 U9775 ( .A1(n9752), .A2(n9736), .A3(n9712), .A4(n7974), .ZN(n7976)
         );
  XNOR2_X1 U9776 ( .A(n9824), .B(n9686), .ZN(n9706) );
  NAND2_X1 U9777 ( .A1(n9706), .A2(n9684), .ZN(n7975) );
  NOR3_X1 U9778 ( .A1(n9670), .A2(n7976), .A3(n7975), .ZN(n7977) );
  NAND4_X1 U9779 ( .A1(n9604), .A2(n9655), .A3(n9639), .A4(n7977), .ZN(n7979)
         );
  NOR4_X1 U9780 ( .A1(n7980), .A2(n7979), .A3(n9629), .A4(n9586), .ZN(n7982)
         );
  NAND4_X1 U9781 ( .A1(n7983), .A2(n8077), .A3(n7982), .A4(n7981), .ZN(n8029)
         );
  NAND4_X1 U9782 ( .A1(n8034), .A2(n6602), .A3(n8014), .A4(n8029), .ZN(n8037)
         );
  NOR2_X1 U9783 ( .A1(n7984), .A2(n6294), .ZN(n7988) );
  NAND2_X1 U9784 ( .A1(n8014), .A2(n7985), .ZN(n8023) );
  AOI211_X1 U9785 ( .C1(n8018), .C2(n6602), .A(n7986), .B(n8023), .ZN(n7987)
         );
  OAI21_X1 U9786 ( .B1(n7989), .B2(n7988), .A(n7987), .ZN(n8036) );
  INV_X1 U9787 ( .A(n7990), .ZN(n7998) );
  INV_X1 U9788 ( .A(n7991), .ZN(n7992) );
  AOI21_X1 U9789 ( .B1(n7998), .B2(n9715), .A(n8046), .ZN(n8002) );
  INV_X1 U9790 ( .A(n7999), .ZN(n8001) );
  OAI21_X1 U9791 ( .B1(n8002), .B2(n8001), .A(n8000), .ZN(n8007) );
  INV_X1 U9792 ( .A(n8003), .ZN(n8006) );
  INV_X1 U9793 ( .A(n8010), .ZN(n8005) );
  AOI22_X1 U9794 ( .A1(n8007), .A2(n8006), .B1(n8005), .B2(n8004), .ZN(n8013)
         );
  INV_X1 U9795 ( .A(n8008), .ZN(n8012) );
  INV_X1 U9796 ( .A(n8009), .ZN(n8011) );
  AOI22_X1 U9797 ( .A1(n8013), .A2(n8012), .B1(n8011), .B2(n8010), .ZN(n8019)
         );
  NAND2_X1 U9798 ( .A1(n6294), .A2(n8014), .ZN(n8028) );
  NOR3_X1 U9799 ( .A1(n8016), .A2(n8015), .A3(n8028), .ZN(n8017) );
  OAI21_X1 U9800 ( .B1(n8019), .B2(n8018), .A(n8017), .ZN(n8020) );
  OAI21_X1 U9801 ( .B1(n8022), .B2(n8021), .A(n8020), .ZN(n8033) );
  INV_X1 U9802 ( .A(n8023), .ZN(n8025) );
  INV_X1 U9803 ( .A(P1_B_REG_SCAN_IN), .ZN(n8024) );
  AOI211_X1 U9804 ( .C1(n8027), .C2(n8026), .A(n8025), .B(n8024), .ZN(n8032)
         );
  NOR3_X1 U9805 ( .A1(n8030), .A2(n8029), .A3(n8028), .ZN(n8031) );
  OAI211_X1 U9806 ( .C1(n8038), .C2(n8037), .A(n8036), .B(n8035), .ZN(P1_U3242) );
  INV_X1 U9807 ( .A(n8042), .ZN(n8043) );
  NAND2_X1 U9808 ( .A1(n9603), .A2(n8047), .ZN(n9585) );
  NAND2_X1 U9809 ( .A1(n9589), .A2(n8048), .ZN(n8050) );
  XNOR2_X1 U9810 ( .A(n8050), .B(n8049), .ZN(n8055) );
  NAND2_X1 U9811 ( .A1(n8051), .A2(n9487), .ZN(n8052) );
  INV_X1 U9812 ( .A(n9848), .ZN(n8056) );
  OAI22_X1 U9813 ( .A1(n8058), .A2(n8057), .B1(n9476), .B2(n8056), .ZN(n9760)
         );
  NOR2_X1 U9814 ( .A1(n9767), .A2(n9453), .ZN(n8059) );
  NOR2_X1 U9815 ( .A1(n7834), .A2(n9772), .ZN(n8060) );
  NAND2_X1 U9816 ( .A1(n9829), .A2(n9490), .ZN(n8061) );
  NAND2_X1 U9817 ( .A1(n8064), .A2(n4977), .ZN(n9682) );
  NOR2_X1 U9818 ( .A1(n9695), .A2(n9709), .ZN(n8066) );
  NAND2_X1 U9819 ( .A1(n9695), .A2(n9709), .ZN(n8065) );
  NOR2_X1 U9820 ( .A1(n9814), .A2(n9687), .ZN(n8068) );
  NAND2_X1 U9821 ( .A1(n9664), .A2(n9673), .ZN(n8070) );
  NOR2_X1 U9822 ( .A1(n9664), .A2(n9673), .ZN(n8069) );
  NAND2_X1 U9823 ( .A1(n9804), .A2(n9657), .ZN(n8071) );
  NAND2_X1 U9824 ( .A1(n9650), .A2(n9630), .ZN(n8072) );
  NOR2_X1 U9825 ( .A1(n9800), .A2(n9642), .ZN(n8075) );
  NAND2_X1 U9826 ( .A1(n9788), .A2(n9488), .ZN(n8076) );
  NAND2_X1 U9827 ( .A1(n9583), .A2(n8076), .ZN(n8078) );
  XNOR2_X1 U9828 ( .A(n8078), .B(n8077), .ZN(n9783) );
  NAND2_X1 U9829 ( .A1(n9783), .A2(n10032), .ZN(n8087) );
  NAND2_X1 U9830 ( .A1(n10015), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n8080) );
  INV_X1 U9831 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n8079) );
  OAI22_X1 U9832 ( .A1(n8081), .A2(n8080), .B1(n8079), .B2(n10070), .ZN(n8084)
         );
  OAI211_X1 U9833 ( .C1(n9595), .C2(n9784), .A(n10027), .B(n8082), .ZN(n9786)
         );
  NOR2_X1 U9834 ( .A1(n9786), .A2(n9581), .ZN(n8083) );
  AOI211_X1 U9835 ( .C1(n10017), .C2(n8085), .A(n8084), .B(n8083), .ZN(n8086)
         );
  OAI211_X1 U9836 ( .C1(n9787), .C2(n4984), .A(n8087), .B(n8086), .ZN(P1_U3356) );
  NOR2_X1 U9837 ( .A1(n8088), .A2(n10165), .ZN(n8649) );
  NOR2_X1 U9838 ( .A1(n8089), .A2(n8784), .ZN(n8090) );
  AOI211_X1 U9839 ( .C1(n10174), .C2(P2_REG2_REG_29__SCAN_IN), .A(n8649), .B(
        n8090), .ZN(n8093) );
  OR2_X1 U9840 ( .A1(n8091), .A2(n8855), .ZN(n8092) );
  OAI211_X1 U9841 ( .C1(n8094), .C2(n10174), .A(n8093), .B(n8092), .ZN(
        P2_U3204) );
  OAI222_X1 U9842 ( .A1(n9283), .A2(n8096), .B1(n9281), .B2(n8095), .C1(n4274), 
        .C2(P2_U3151), .ZN(P2_U3276) );
  XOR2_X1 U9843 ( .A(n8098), .B(n8097), .Z(n8103) );
  NAND2_X1 U9844 ( .A1(n8264), .A2(n8818), .ZN(n8099) );
  NAND2_X1 U9845 ( .A1(P2_U3151), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n8556) );
  OAI211_X1 U9846 ( .C1(n8266), .C2(n8847), .A(n8099), .B(n8556), .ZN(n8101)
         );
  NOR2_X1 U9847 ( .A1(n8361), .A2(n8291), .ZN(n8100) );
  AOI211_X1 U9848 ( .C1(n8821), .C2(n8288), .A(n8101), .B(n8100), .ZN(n8102)
         );
  OAI21_X1 U9849 ( .B1(n8103), .B2(n8279), .A(n8102), .ZN(P2_U3155) );
  XNOR2_X1 U9850 ( .A(n8205), .B(n8206), .ZN(n8207) );
  XNOR2_X1 U9851 ( .A(n8207), .B(n8712), .ZN(n8108) );
  AOI22_X1 U9852 ( .A1(n8724), .A2(n8283), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3151), .ZN(n8105) );
  NAND2_X1 U9853 ( .A1(n8728), .A2(n8288), .ZN(n8104) );
  OAI211_X1 U9854 ( .C1(n8702), .C2(n8285), .A(n8105), .B(n8104), .ZN(n8106)
         );
  AOI21_X1 U9855 ( .B1(n9191), .B2(n8276), .A(n8106), .ZN(n8107) );
  OAI21_X1 U9856 ( .B1(n8108), .B2(n8279), .A(n8107), .ZN(P2_U3156) );
  XOR2_X1 U9857 ( .A(n8110), .B(n8109), .Z(n8148) );
  NOR2_X1 U9858 ( .A1(n8148), .A2(n8891), .ZN(n8147) );
  AOI21_X1 U9859 ( .B1(n4772), .B2(n8110), .A(n8147), .ZN(n8219) );
  XNOR2_X1 U9860 ( .A(n8111), .B(n8916), .ZN(n8218) );
  NAND2_X1 U9861 ( .A1(n8219), .A2(n8218), .ZN(n8217) );
  NAND2_X1 U9862 ( .A1(n8217), .A2(n8112), .ZN(n8115) );
  XNOR2_X1 U9863 ( .A(n8113), .B(n8889), .ZN(n8114) );
  XNOR2_X1 U9864 ( .A(n8115), .B(n8114), .ZN(n8121) );
  NAND2_X1 U9865 ( .A1(n8283), .A2(n8916), .ZN(n8116) );
  OAI211_X1 U9866 ( .C1(n8846), .C2(n8285), .A(n8117), .B(n8116), .ZN(n8119)
         );
  NOR2_X1 U9867 ( .A1(n9260), .A2(n8291), .ZN(n8118) );
  AOI211_X1 U9868 ( .C1(n8874), .C2(n8288), .A(n8119), .B(n8118), .ZN(n8120)
         );
  OAI21_X1 U9869 ( .B1(n8121), .B2(n8279), .A(n8120), .ZN(P2_U3157) );
  INV_X1 U9870 ( .A(n9213), .ZN(n8131) );
  AOI21_X1 U9871 ( .B1(n8123), .B2(n8122), .A(n8279), .ZN(n8125) );
  NAND2_X1 U9872 ( .A1(n8125), .A2(n8124), .ZN(n8130) );
  NAND2_X1 U9873 ( .A1(n8793), .A2(n8283), .ZN(n8126) );
  OAI211_X1 U9874 ( .C1(n8769), .C2(n8285), .A(n8127), .B(n8126), .ZN(n8128)
         );
  AOI21_X1 U9875 ( .B1(n8773), .B2(n8288), .A(n8128), .ZN(n8129) );
  OAI211_X1 U9876 ( .C1(n8131), .C2(n8291), .A(n8130), .B(n8129), .ZN(P2_U3159) );
  XNOR2_X1 U9877 ( .A(n8673), .B(n8132), .ZN(n8133) );
  XNOR2_X1 U9878 ( .A(n9159), .B(n8133), .ZN(n8140) );
  INV_X1 U9879 ( .A(n8140), .ZN(n8134) );
  NAND2_X1 U9880 ( .A1(n8134), .A2(n8216), .ZN(n8146) );
  AOI22_X1 U9881 ( .A1(n8662), .A2(n8288), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3151), .ZN(n8137) );
  NAND2_X1 U9882 ( .A1(n8686), .A2(n8283), .ZN(n8136) );
  OAI211_X1 U9883 ( .C1(n8531), .C2(n8285), .A(n8137), .B(n8136), .ZN(n8142)
         );
  INV_X1 U9884 ( .A(n8138), .ZN(n8139) );
  NOR4_X1 U9885 ( .A1(n8140), .A2(n8139), .A3(n8274), .A4(n8279), .ZN(n8141)
         );
  AOI211_X1 U9886 ( .C1(n9159), .C2(n8276), .A(n8142), .B(n8141), .ZN(n8143)
         );
  OAI211_X1 U9887 ( .C1(n8146), .C2(n8145), .A(n8144), .B(n8143), .ZN(P2_U3160) );
  AOI21_X1 U9888 ( .B1(n8891), .B2(n8148), .A(n8147), .ZN(n8155) );
  NAND2_X1 U9889 ( .A1(n8264), .A2(n8916), .ZN(n8149) );
  OAI211_X1 U9890 ( .C1(n8266), .C2(n8906), .A(n8150), .B(n8149), .ZN(n8153)
         );
  NOR2_X1 U9891 ( .A1(n8291), .A2(n8151), .ZN(n8152) );
  AOI211_X1 U9892 ( .C1(n8919), .C2(n8288), .A(n8153), .B(n8152), .ZN(n8154)
         );
  OAI21_X1 U9893 ( .B1(n8155), .B2(n8279), .A(n8154), .ZN(P2_U3161) );
  XOR2_X1 U9894 ( .A(n8156), .B(n8157), .Z(n8162) );
  AOI22_X1 U9895 ( .A1(n8532), .A2(n8283), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3151), .ZN(n8159) );
  NAND2_X1 U9896 ( .A1(n8748), .A2(n8288), .ZN(n8158) );
  OAI211_X1 U9897 ( .C1(n8747), .C2(n8285), .A(n8159), .B(n8158), .ZN(n8160)
         );
  AOI21_X1 U9898 ( .B1(n8954), .B2(n8276), .A(n8160), .ZN(n8161) );
  OAI21_X1 U9899 ( .B1(n8162), .B2(n8279), .A(n8161), .ZN(P2_U3163) );
  INV_X1 U9900 ( .A(n8846), .ZN(n8869) );
  MUX2_X1 U9901 ( .A(n8869), .B(n8164), .S(n8163), .Z(n8237) );
  NOR2_X1 U9902 ( .A1(n8235), .A2(n8165), .ZN(n8166) );
  XNOR2_X1 U9903 ( .A(n8237), .B(n8166), .ZN(n8173) );
  NAND2_X1 U9904 ( .A1(n8264), .A2(n8819), .ZN(n8168) );
  OAI211_X1 U9905 ( .C1(n8266), .C2(n8846), .A(n8168), .B(n8167), .ZN(n8171)
         );
  NOR2_X1 U9906 ( .A1(n8169), .A2(n8291), .ZN(n8170) );
  AOI211_X1 U9907 ( .C1(n8849), .C2(n8288), .A(n8171), .B(n8170), .ZN(n8172)
         );
  OAI21_X1 U9908 ( .B1(n8173), .B2(n8279), .A(n8172), .ZN(P2_U3164) );
  XOR2_X1 U9909 ( .A(n8175), .B(n8174), .Z(n8181) );
  AOI22_X1 U9910 ( .A1(n8704), .A2(n8288), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3151), .ZN(n8177) );
  NAND2_X1 U9911 ( .A1(n8725), .A2(n8283), .ZN(n8176) );
  OAI211_X1 U9912 ( .C1(n8178), .C2(n8285), .A(n8177), .B(n8176), .ZN(n8179)
         );
  AOI21_X1 U9913 ( .B1(n9178), .B2(n8276), .A(n8179), .ZN(n8180) );
  OAI21_X1 U9914 ( .B1(n8181), .B2(n8279), .A(n8180), .ZN(P2_U3165) );
  NAND2_X1 U9915 ( .A1(n8281), .A2(n8183), .ZN(n8194) );
  XNOR2_X1 U9916 ( .A(n8184), .B(n8286), .ZN(n8185) );
  XNOR2_X1 U9917 ( .A(n8194), .B(n8185), .ZN(n8191) );
  NAND2_X1 U9918 ( .A1(n8283), .A2(n8818), .ZN(n8186) );
  NAND2_X1 U9919 ( .A1(P2_U3151), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8588) );
  OAI211_X1 U9920 ( .C1(n8778), .C2(n8285), .A(n8186), .B(n8588), .ZN(n8189)
         );
  NOR2_X1 U9921 ( .A1(n8187), .A2(n8291), .ZN(n8188) );
  AOI211_X1 U9922 ( .C1(n8805), .C2(n8288), .A(n8189), .B(n8188), .ZN(n8190)
         );
  OAI21_X1 U9923 ( .B1(n8191), .B2(n8279), .A(n8190), .ZN(P2_U3166) );
  NAND2_X1 U9924 ( .A1(n8193), .A2(n8192), .ZN(n8199) );
  NAND2_X1 U9925 ( .A1(n8195), .A2(n8194), .ZN(n8197) );
  NAND2_X1 U9926 ( .A1(n8197), .A2(n8196), .ZN(n8198) );
  XOR2_X1 U9927 ( .A(n8199), .B(n8198), .Z(n8204) );
  NAND2_X1 U9928 ( .A1(n8811), .A2(n8283), .ZN(n8200) );
  NAND2_X1 U9929 ( .A1(P2_U3151), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n8612) );
  OAI211_X1 U9930 ( .C1(n8768), .C2(n8285), .A(n8200), .B(n8612), .ZN(n8201)
         );
  AOI21_X1 U9931 ( .B1(n8796), .B2(n8288), .A(n8201), .ZN(n8203) );
  NAND2_X1 U9932 ( .A1(n9223), .A2(n8276), .ZN(n8202) );
  OAI211_X1 U9933 ( .C1(n8204), .C2(n8279), .A(n8203), .B(n8202), .ZN(P2_U3168) );
  OAI22_X1 U9934 ( .A1(n8207), .A2(n8734), .B1(n8206), .B2(n8205), .ZN(n8210)
         );
  XNOR2_X1 U9935 ( .A(n8208), .B(n8702), .ZN(n8209) );
  XNOR2_X1 U9936 ( .A(n8210), .B(n8209), .ZN(n8215) );
  AOI22_X1 U9937 ( .A1(n8714), .A2(n8288), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3151), .ZN(n8212) );
  NAND2_X1 U9938 ( .A1(n8734), .A2(n8283), .ZN(n8211) );
  OAI211_X1 U9939 ( .C1(n8711), .C2(n8285), .A(n8212), .B(n8211), .ZN(n8213)
         );
  AOI21_X1 U9940 ( .B1(n9185), .B2(n8276), .A(n8213), .ZN(n8214) );
  OAI21_X1 U9941 ( .B1(n8215), .B2(n8279), .A(n8214), .ZN(P2_U3169) );
  INV_X1 U9942 ( .A(n8898), .ZN(n9265) );
  OAI211_X1 U9943 ( .C1(n8219), .C2(n8218), .A(n8217), .B(n8216), .ZN(n8225)
         );
  NAND2_X1 U9944 ( .A1(n8264), .A2(n8889), .ZN(n8221) );
  OAI211_X1 U9945 ( .C1(n8266), .C2(n8222), .A(n8221), .B(n8220), .ZN(n8223)
         );
  AOI21_X1 U9946 ( .B1(n8897), .B2(n8288), .A(n8223), .ZN(n8224) );
  OAI211_X1 U9947 ( .C1(n9265), .C2(n8291), .A(n8225), .B(n8224), .ZN(P2_U3171) );
  INV_X1 U9948 ( .A(n8226), .ZN(n8227) );
  AOI21_X1 U9949 ( .B1(n8229), .B2(n8228), .A(n8227), .ZN(n8234) );
  AOI22_X1 U9950 ( .A1(n8757), .A2(n8283), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3151), .ZN(n8231) );
  NAND2_X1 U9951 ( .A1(n8761), .A2(n8288), .ZN(n8230) );
  OAI211_X1 U9952 ( .C1(n8253), .C2(n8285), .A(n8231), .B(n8230), .ZN(n8232)
         );
  AOI21_X1 U9953 ( .B1(n9207), .B2(n8276), .A(n8232), .ZN(n8233) );
  OAI21_X1 U9954 ( .B1(n8234), .B2(n8279), .A(n8233), .ZN(P2_U3173) );
  AOI21_X1 U9955 ( .B1(n8237), .B2(n8236), .A(n8235), .ZN(n8239) );
  XNOR2_X1 U9956 ( .A(n8239), .B(n8238), .ZN(n8245) );
  NAND2_X1 U9957 ( .A1(n8830), .A2(n8264), .ZN(n8240) );
  NAND2_X1 U9958 ( .A1(P2_U3151), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n8543) );
  OAI211_X1 U9959 ( .C1(n8355), .C2(n8266), .A(n8240), .B(n8543), .ZN(n8243)
         );
  NOR2_X1 U9960 ( .A1(n8241), .A2(n8291), .ZN(n8242) );
  AOI211_X1 U9961 ( .C1(n8832), .C2(n8288), .A(n8243), .B(n8242), .ZN(n8244)
         );
  OAI21_X1 U9962 ( .B1(n8245), .B2(n8279), .A(n8244), .ZN(P2_U3174) );
  NAND2_X1 U9963 ( .A1(n8247), .A2(n8246), .ZN(n8249) );
  AOI21_X1 U9964 ( .B1(n8249), .B2(n8248), .A(n8279), .ZN(n8251) );
  NAND2_X1 U9965 ( .A1(n8251), .A2(n8250), .ZN(n8258) );
  INV_X1 U9966 ( .A(n8252), .ZN(n8736) );
  AOI22_X1 U9967 ( .A1(n8758), .A2(n8283), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3151), .ZN(n8254) );
  OAI21_X1 U9968 ( .B1(n8736), .B2(n8255), .A(n8254), .ZN(n8256) );
  AOI21_X1 U9969 ( .B1(n8264), .B2(n8734), .A(n8256), .ZN(n8257) );
  OAI211_X1 U9970 ( .C1(n8259), .C2(n8291), .A(n8258), .B(n8257), .ZN(P2_U3175) );
  NAND2_X1 U9971 ( .A1(n4765), .A2(n8261), .ZN(n8262) );
  XOR2_X1 U9972 ( .A(n8263), .B(n8262), .Z(n8270) );
  NAND2_X1 U9973 ( .A1(n8757), .A2(n8264), .ZN(n8265) );
  NAND2_X1 U9974 ( .A1(P2_U3151), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8632) );
  OAI211_X1 U9975 ( .C1(n8778), .C2(n8266), .A(n8265), .B(n8632), .ZN(n8268)
         );
  NOR2_X1 U9976 ( .A1(n9220), .A2(n8291), .ZN(n8267) );
  AOI211_X1 U9977 ( .C1(n8782), .C2(n8288), .A(n8268), .B(n8267), .ZN(n8269)
         );
  OAI21_X1 U9978 ( .B1(n8270), .B2(n8279), .A(n8269), .ZN(P2_U3178) );
  XNOR2_X1 U9979 ( .A(n8271), .B(n8699), .ZN(n8278) );
  AOI22_X1 U9980 ( .A1(n8693), .A2(n8288), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3151), .ZN(n8273) );
  NAND2_X1 U9981 ( .A1(n8687), .A2(n8283), .ZN(n8272) );
  OAI211_X1 U9982 ( .C1(n8274), .C2(n8285), .A(n8273), .B(n8272), .ZN(n8275)
         );
  AOI21_X1 U9983 ( .B1(n9171), .B2(n8276), .A(n8275), .ZN(n8277) );
  OAI21_X1 U9984 ( .B1(n8278), .B2(n8279), .A(n8277), .ZN(P2_U3180) );
  AOI21_X1 U9985 ( .B1(n8182), .B2(n8280), .A(n8279), .ZN(n8282) );
  NAND2_X1 U9986 ( .A1(n8282), .A2(n8281), .ZN(n8290) );
  NAND2_X1 U9987 ( .A1(n8830), .A2(n8283), .ZN(n8284) );
  NAND2_X1 U9988 ( .A1(P2_U3151), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8574) );
  OAI211_X1 U9989 ( .C1(n8286), .C2(n8285), .A(n8284), .B(n8574), .ZN(n8287)
         );
  AOI21_X1 U9990 ( .B1(n8814), .B2(n8288), .A(n8287), .ZN(n8289) );
  OAI211_X1 U9991 ( .C1(n8292), .C2(n8291), .A(n8290), .B(n8289), .ZN(P2_U3181) );
  NOR2_X1 U9992 ( .A1(n8733), .A2(n8386), .ZN(n8409) );
  NOR2_X1 U9993 ( .A1(n8484), .A2(n8294), .ZN(n8304) );
  NOR2_X1 U9994 ( .A1(n8294), .A2(n8525), .ZN(n8296) );
  INV_X1 U9995 ( .A(n8300), .ZN(n8303) );
  INV_X1 U9996 ( .A(n8298), .ZN(n8301) );
  NAND2_X1 U9997 ( .A1(n8538), .A2(n10164), .ZN(n8305) );
  NAND2_X1 U9998 ( .A1(n8313), .A2(n8305), .ZN(n8308) );
  INV_X1 U9999 ( .A(n8306), .ZN(n8307) );
  MUX2_X1 U10000 ( .A(n8308), .B(n8307), .S(n8504), .Z(n8310) );
  INV_X1 U10001 ( .A(n8317), .ZN(n8314) );
  OAI211_X1 U10002 ( .C1(n8319), .C2(n8318), .A(n8317), .B(n8316), .ZN(n8324)
         );
  NOR2_X1 U10003 ( .A1(n4910), .A2(n8321), .ZN(n8323) );
  AOI21_X1 U10004 ( .B1(n8324), .B2(n8323), .A(n8322), .ZN(n8325) );
  MUX2_X1 U10005 ( .A(n8326), .B(n8325), .S(n8440), .Z(n8329) );
  MUX2_X1 U10006 ( .A(n8327), .B(n8333), .S(n8504), .Z(n8328) );
  NAND3_X1 U10007 ( .A1(n8329), .A2(n8479), .A3(n8330), .ZN(n8354) );
  OAI21_X1 U10008 ( .B1(n8332), .B2(n8879), .A(n8331), .ZN(n8339) );
  AOI21_X1 U10009 ( .B1(n8334), .B2(n8333), .A(n8332), .ZN(n8337) );
  INV_X1 U10010 ( .A(n8335), .ZN(n8336) );
  AOI211_X1 U10011 ( .C1(n8504), .C2(n8339), .A(n8493), .B(n8338), .ZN(n8353)
         );
  NOR2_X1 U10012 ( .A1(n8869), .A2(n8440), .ZN(n8344) );
  INV_X1 U10013 ( .A(n8344), .ZN(n8342) );
  NAND3_X1 U10014 ( .A1(n8875), .A2(n8345), .A3(n8504), .ZN(n8341) );
  AOI21_X1 U10015 ( .B1(n8342), .B2(n8341), .A(n8340), .ZN(n8352) );
  INV_X1 U10016 ( .A(n8491), .ZN(n8343) );
  NOR2_X1 U10017 ( .A1(n8846), .A2(n8504), .ZN(n8346) );
  AOI21_X1 U10018 ( .B1(n8343), .B2(n8440), .A(n8346), .ZN(n8350) );
  AOI21_X1 U10019 ( .B1(n8345), .B2(n8344), .A(n9260), .ZN(n8348) );
  AOI21_X1 U10020 ( .B1(n8346), .B2(n8889), .A(n8875), .ZN(n8347) );
  OAI22_X1 U10021 ( .A1(n8350), .A2(n8349), .B1(n8348), .B2(n8347), .ZN(n8351)
         );
  NAND2_X1 U10022 ( .A1(n6663), .A2(n8355), .ZN(n8357) );
  MUX2_X1 U10023 ( .A(n8357), .B(n8356), .S(n8440), .Z(n8358) );
  MUX2_X1 U10024 ( .A(n9248), .B(n8819), .S(n8440), .Z(n8359) );
  NOR2_X1 U10025 ( .A1(n8361), .A2(n8830), .ZN(n8363) );
  MUX2_X1 U10026 ( .A(n8363), .B(n8362), .S(n8440), .Z(n8366) );
  INV_X1 U10027 ( .A(n8374), .ZN(n8368) );
  NOR2_X1 U10028 ( .A1(n8368), .A2(n8367), .ZN(n8370) );
  MUX2_X1 U10029 ( .A(n8370), .B(n8369), .S(n8504), .Z(n8372) );
  NAND2_X1 U10030 ( .A1(n8372), .A2(n8371), .ZN(n8373) );
  INV_X1 U10031 ( .A(n8789), .ZN(n8792) );
  NOR2_X1 U10032 ( .A1(n8374), .A2(n8440), .ZN(n8376) );
  INV_X1 U10033 ( .A(n8475), .ZN(n8384) );
  OAI211_X1 U10034 ( .C1(n8378), .C2(n8376), .A(n8384), .B(n8375), .ZN(n8380)
         );
  OAI21_X1 U10035 ( .B1(n8378), .B2(n8377), .A(n8440), .ZN(n8379) );
  AND2_X1 U10036 ( .A1(n8381), .A2(n8440), .ZN(n8382) );
  INV_X1 U10037 ( .A(n8383), .ZN(n8389) );
  NAND3_X1 U10038 ( .A1(n8391), .A2(n8440), .A3(n8384), .ZN(n8385) );
  OAI21_X1 U10039 ( .B1(n8504), .B2(n8390), .A(n8385), .ZN(n8388) );
  NOR3_X1 U10040 ( .A1(n8392), .A2(n8440), .A3(n4948), .ZN(n8393) );
  OAI22_X1 U10041 ( .A1(n8396), .A2(n8395), .B1(n8394), .B2(n8393), .ZN(n8397)
         );
  AOI21_X1 U10042 ( .B1(n8400), .B2(n8398), .A(n8504), .ZN(n8399) );
  INV_X1 U10043 ( .A(n8405), .ZN(n8408) );
  NAND2_X1 U10044 ( .A1(n8473), .A2(n8402), .ZN(n8407) );
  OAI211_X1 U10045 ( .C1(n8405), .C2(n8733), .A(n8715), .B(n8404), .ZN(n8406)
         );
  INV_X1 U10046 ( .A(n8473), .ZN(n8412) );
  NOR3_X1 U10047 ( .A1(n8410), .A2(n8440), .A3(n8471), .ZN(n8411) );
  INV_X1 U10048 ( .A(n8413), .ZN(n8429) );
  INV_X1 U10049 ( .A(n8684), .ZN(n8415) );
  NOR3_X1 U10050 ( .A1(n8415), .A2(n8504), .A3(n8420), .ZN(n8416) );
  AOI211_X1 U10051 ( .C1(n8427), .C2(n8504), .A(n8665), .B(n8416), .ZN(n8422)
         );
  INV_X1 U10052 ( .A(n8472), .ZN(n8424) );
  NAND3_X1 U10053 ( .A1(n8425), .A2(n8504), .A3(n8424), .ZN(n8419) );
  XNOR2_X1 U10054 ( .A(n8417), .B(n8504), .ZN(n8418) );
  OAI211_X1 U10055 ( .C1(n8440), .C2(n8420), .A(n8419), .B(n8418), .ZN(n8421)
         );
  NAND3_X1 U10056 ( .A1(n8425), .A2(n8440), .A3(n8424), .ZN(n8426) );
  MUX2_X1 U10057 ( .A(n8430), .B(n8429), .S(n8504), .Z(n8431) );
  MUX2_X1 U10058 ( .A(n8673), .B(n9159), .S(n8504), .Z(n8442) );
  NOR2_X1 U10059 ( .A1(n9159), .A2(n8504), .ZN(n8434) );
  NOR2_X1 U10060 ( .A1(n8673), .A2(n8440), .ZN(n8443) );
  NOR3_X1 U10061 ( .A1(n8442), .A2(n8434), .A3(n8443), .ZN(n8432) );
  NOR2_X1 U10062 ( .A1(n8466), .A2(n8504), .ZN(n8447) );
  INV_X1 U10063 ( .A(n8500), .ZN(n8441) );
  NOR3_X1 U10064 ( .A1(n8432), .A2(n8447), .A3(n8441), .ZN(n8449) );
  INV_X1 U10065 ( .A(n8466), .ZN(n8433) );
  AOI21_X1 U10066 ( .B1(n8434), .B2(n8442), .A(n8433), .ZN(n8446) );
  NAND2_X1 U10067 ( .A1(n9272), .A2(n8450), .ZN(n8437) );
  OR2_X1 U10068 ( .A1(n8435), .A2(n9274), .ZN(n8436) );
  NAND2_X1 U10069 ( .A1(n9153), .A2(n8438), .ZN(n8467) );
  INV_X1 U10070 ( .A(n8467), .ZN(n8439) );
  INV_X1 U10071 ( .A(n8438), .ZN(n8530) );
  AND2_X1 U10072 ( .A1(n8928), .A2(n8530), .ZN(n8506) );
  AOI211_X1 U10073 ( .C1(n8441), .C2(n8440), .A(n8439), .B(n8506), .ZN(n8445)
         );
  NAND3_X1 U10074 ( .A1(n8500), .A2(n8443), .A3(n8442), .ZN(n8444) );
  OAI211_X1 U10075 ( .C1(n8447), .C2(n8446), .A(n8445), .B(n8444), .ZN(n8448)
         );
  NAND2_X1 U10076 ( .A1(n9267), .A2(n8450), .ZN(n8454) );
  OR2_X1 U10077 ( .A1(n8452), .A2(n8451), .ZN(n8453) );
  NAND2_X1 U10078 ( .A1(n8454), .A2(n8453), .ZN(n8507) );
  NAND2_X1 U10079 ( .A1(n8455), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n8460) );
  NAND2_X1 U10080 ( .A1(n4272), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n8459) );
  NAND2_X1 U10081 ( .A1(n8457), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n8458) );
  AND3_X1 U10082 ( .A1(n8460), .A2(n8459), .A3(n8458), .ZN(n8461) );
  OR2_X1 U10083 ( .A1(n8507), .A2(n8648), .ZN(n8516) );
  INV_X1 U10084 ( .A(n8463), .ZN(n8464) );
  NAND4_X1 U10085 ( .A1(n8516), .A2(n8464), .A3(n8525), .A4(n8467), .ZN(n8519)
         );
  NAND2_X1 U10086 ( .A1(n8465), .A2(n8500), .ZN(n8514) );
  AND2_X1 U10087 ( .A1(n8467), .A2(n8466), .ZN(n8468) );
  NAND2_X1 U10088 ( .A1(n8516), .A2(n8468), .ZN(n8502) );
  AOI211_X1 U10089 ( .C1(n9152), .C2(n9153), .A(n8469), .B(n8502), .ZN(n8513)
         );
  INV_X1 U10090 ( .A(n8764), .ZN(n8767) );
  NOR2_X1 U10091 ( .A1(n8475), .A2(n4953), .ZN(n8781) );
  OR2_X1 U10092 ( .A1(n8477), .A2(n4929), .ZN(n8835) );
  INV_X1 U10093 ( .A(n8881), .ZN(n8885) );
  NAND3_X1 U10094 ( .A1(n8480), .A2(n8479), .A3(n8478), .ZN(n8483) );
  INV_X1 U10095 ( .A(n8481), .ZN(n8482) );
  NOR4_X1 U10096 ( .A1(n8485), .A2(n8484), .A3(n8483), .A4(n8482), .ZN(n8489)
         );
  INV_X1 U10097 ( .A(n8908), .ZN(n8488) );
  NAND4_X1 U10098 ( .A1(n8489), .A2(n8488), .A3(n8487), .A4(n8486), .ZN(n8494)
         );
  INV_X1 U10099 ( .A(n8490), .ZN(n8492) );
  NAND2_X1 U10100 ( .A1(n8492), .A2(n8491), .ZN(n8867) );
  NOR4_X1 U10101 ( .A1(n8885), .A2(n8494), .A3(n8493), .A4(n8867), .ZN(n8495)
         );
  NAND4_X1 U10102 ( .A1(n8835), .A2(n8495), .A3(n8823), .A4(n6630), .ZN(n8496)
         );
  NOR3_X1 U10103 ( .A1(n8496), .A2(n8809), .A3(n8789), .ZN(n8497) );
  AND4_X1 U10104 ( .A1(n8705), .A2(n8717), .A3(n8723), .A4(n8498), .ZN(n8499)
         );
  NAND4_X1 U10105 ( .A1(n8500), .A2(n8684), .A3(n8671), .A4(n8499), .ZN(n8501)
         );
  NOR4_X1 U10106 ( .A1(n8502), .A2(n8506), .A3(n8655), .A4(n8501), .ZN(n8511)
         );
  INV_X1 U10107 ( .A(n8506), .ZN(n8505) );
  INV_X1 U10108 ( .A(n8648), .ZN(n8529) );
  NAND2_X1 U10109 ( .A1(n8504), .A2(n8503), .ZN(n8515) );
  NOR3_X1 U10110 ( .A1(n8505), .A2(n8529), .A3(n8515), .ZN(n8508) );
  OAI22_X1 U10111 ( .A1(n8508), .A2(n8507), .B1(n8506), .B2(n8648), .ZN(n8509)
         );
  OAI21_X1 U10112 ( .B1(n8511), .B2(n8510), .A(n8509), .ZN(n8512) );
  AOI21_X1 U10113 ( .B1(n8514), .B2(n8513), .A(n8512), .ZN(n8518) );
  INV_X1 U10114 ( .A(n8515), .ZN(n8517) );
  XNOR2_X1 U10115 ( .A(n8521), .B(n4274), .ZN(n8528) );
  NAND3_X1 U10116 ( .A1(n8523), .A2(n8522), .A3(n4271), .ZN(n8524) );
  OAI211_X1 U10117 ( .C1(n8525), .C2(n8527), .A(n8524), .B(P2_B_REG_SCAN_IN), 
        .ZN(n8526) );
  OAI21_X1 U10118 ( .B1(n8528), .B2(n8527), .A(n8526), .ZN(P2_U3296) );
  MUX2_X1 U10119 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n8529), .S(P2_U3893), .Z(
        P2_U3522) );
  MUX2_X1 U10120 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n8530), .S(P2_U3893), .Z(
        P2_U3521) );
  INV_X1 U10121 ( .A(n8531), .ZN(n8656) );
  MUX2_X1 U10122 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n8656), .S(P2_U3893), .Z(
        P2_U3520) );
  MUX2_X1 U10123 ( .A(n8673), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8623), .Z(
        P2_U3519) );
  MUX2_X1 U10124 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8686), .S(P2_U3893), .Z(
        P2_U3518) );
  MUX2_X1 U10125 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n8699), .S(P2_U3893), .Z(
        P2_U3517) );
  MUX2_X1 U10126 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8687), .S(P2_U3893), .Z(
        P2_U3516) );
  MUX2_X1 U10127 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n8725), .S(P2_U3893), .Z(
        P2_U3515) );
  MUX2_X1 U10128 ( .A(n8734), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8623), .Z(
        P2_U3514) );
  MUX2_X1 U10129 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8724), .S(P2_U3893), .Z(
        P2_U3513) );
  MUX2_X1 U10130 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8758), .S(P2_U3893), .Z(
        P2_U3512) );
  MUX2_X1 U10131 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8532), .S(P2_U3893), .Z(
        P2_U3511) );
  MUX2_X1 U10132 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8757), .S(P2_U3893), .Z(
        P2_U3510) );
  MUX2_X1 U10133 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n8793), .S(P2_U3893), .Z(
        P2_U3509) );
  MUX2_X1 U10134 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8802), .S(P2_U3893), .Z(
        P2_U3508) );
  MUX2_X1 U10135 ( .A(n8811), .B(P2_DATAO_REG_16__SCAN_IN), .S(n8623), .Z(
        P2_U3507) );
  MUX2_X1 U10136 ( .A(n8818), .B(P2_DATAO_REG_15__SCAN_IN), .S(n8623), .Z(
        P2_U3506) );
  MUX2_X1 U10137 ( .A(n8830), .B(P2_DATAO_REG_14__SCAN_IN), .S(n8623), .Z(
        P2_U3505) );
  MUX2_X1 U10138 ( .A(n8819), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8623), .Z(
        P2_U3504) );
  MUX2_X1 U10139 ( .A(n8829), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8623), .Z(
        P2_U3503) );
  MUX2_X1 U10140 ( .A(n8869), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8623), .Z(
        P2_U3502) );
  MUX2_X1 U10141 ( .A(n8889), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8623), .Z(
        P2_U3501) );
  MUX2_X1 U10142 ( .A(n8916), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8623), .Z(
        P2_U3500) );
  MUX2_X1 U10143 ( .A(n8891), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8623), .Z(
        P2_U3499) );
  MUX2_X1 U10144 ( .A(n8533), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8623), .Z(
        P2_U3498) );
  MUX2_X1 U10145 ( .A(n8534), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8623), .Z(
        P2_U3497) );
  MUX2_X1 U10146 ( .A(n8535), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8623), .Z(
        P2_U3496) );
  MUX2_X1 U10147 ( .A(n8536), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8623), .Z(
        P2_U3495) );
  MUX2_X1 U10148 ( .A(n8537), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8623), .Z(
        P2_U3494) );
  MUX2_X1 U10149 ( .A(n8538), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8623), .Z(
        P2_U3493) );
  MUX2_X1 U10150 ( .A(n4967), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8623), .Z(
        P2_U3492) );
  MUX2_X1 U10151 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n4937), .S(P2_U3893), .Z(
        P2_U3491) );
  AOI21_X1 U10152 ( .B1(n8837), .B2(n8539), .A(n4275), .ZN(n8553) );
  XNOR2_X1 U10153 ( .A(n8540), .B(n9021), .ZN(n8542) );
  NAND2_X1 U10154 ( .A1(n8542), .A2(n8541), .ZN(n8552) );
  OAI21_X1 U10155 ( .B1(n8615), .B2(n8544), .A(n8543), .ZN(n8550) );
  OR3_X1 U10156 ( .A1(n8547), .A2(n8546), .A3(n8545), .ZN(n8548) );
  AOI21_X1 U10157 ( .B1(n8560), .B2(n8548), .A(n8626), .ZN(n8549) );
  AOI211_X1 U10158 ( .C1(n8611), .C2(P2_ADDR_REG_13__SCAN_IN), .A(n8550), .B(
        n8549), .ZN(n8551) );
  OAI211_X1 U10159 ( .C1(n8553), .C2(n4586), .A(n8552), .B(n8551), .ZN(
        P2_U3195) );
  XOR2_X1 U10160 ( .A(n8555), .B(n8554), .Z(n8571) );
  OAI21_X1 U10161 ( .B1(n8615), .B2(n8557), .A(n8556), .ZN(n8564) );
  INV_X1 U10162 ( .A(n8579), .ZN(n8562) );
  NAND3_X1 U10163 ( .A1(n8560), .A2(n8559), .A3(n8558), .ZN(n8561) );
  AOI21_X1 U10164 ( .B1(n8562), .B2(n8561), .A(n8626), .ZN(n8563) );
  AOI211_X1 U10165 ( .C1(n8611), .C2(P2_ADDR_REG_14__SCAN_IN), .A(n8564), .B(
        n8563), .ZN(n8570) );
  INV_X1 U10166 ( .A(n8565), .ZN(n8567) );
  NOR3_X1 U10167 ( .A1(n4275), .A2(n8567), .A3(n8566), .ZN(n8568) );
  OAI21_X1 U10168 ( .B1(n8568), .B2(n4356), .A(n8641), .ZN(n8569) );
  OAI211_X1 U10169 ( .C1(n8571), .C2(n8645), .A(n8570), .B(n8569), .ZN(
        P2_U3196) );
  XNOR2_X1 U10170 ( .A(n8572), .B(P2_REG1_REG_15__SCAN_IN), .ZN(n8585) );
  OAI21_X1 U10171 ( .B1(P2_REG2_REG_15__SCAN_IN), .B2(n8573), .A(n8599), .ZN(
        n8583) );
  NAND2_X1 U10172 ( .A1(n8611), .A2(P2_ADDR_REG_15__SCAN_IN), .ZN(n8575) );
  OAI211_X1 U10173 ( .C1(n8615), .C2(n8576), .A(n8575), .B(n8574), .ZN(n8582)
         );
  OR3_X1 U10174 ( .A1(n8579), .A2(n8578), .A3(n8577), .ZN(n8580) );
  AOI21_X1 U10175 ( .B1(n8592), .B2(n8580), .A(n8626), .ZN(n8581) );
  AOI211_X1 U10176 ( .C1(n8641), .C2(n8583), .A(n8582), .B(n8581), .ZN(n8584)
         );
  OAI21_X1 U10177 ( .B1(n8585), .B2(n8645), .A(n8584), .ZN(P2_U3197) );
  XOR2_X1 U10178 ( .A(n8587), .B(n8586), .Z(n8603) );
  OAI21_X1 U10179 ( .B1(n8615), .B2(n8589), .A(n8588), .ZN(n8596) );
  INV_X1 U10180 ( .A(n8608), .ZN(n8594) );
  NAND3_X1 U10181 ( .A1(n8592), .A2(n8591), .A3(n8590), .ZN(n8593) );
  AOI21_X1 U10182 ( .B1(n8594), .B2(n8593), .A(n8626), .ZN(n8595) );
  AOI211_X1 U10183 ( .C1(n8611), .C2(P2_ADDR_REG_16__SCAN_IN), .A(n8596), .B(
        n8595), .ZN(n8602) );
  AND3_X1 U10184 ( .A1(n8599), .A2(n8598), .A3(n8597), .ZN(n8600) );
  OAI21_X1 U10185 ( .B1(n4352), .B2(n8600), .A(n8641), .ZN(n8601) );
  OAI211_X1 U10186 ( .C1(n8603), .C2(n8645), .A(n8602), .B(n8601), .ZN(
        P2_U3198) );
  XNOR2_X1 U10187 ( .A(n8604), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n8620) );
  OAI21_X1 U10188 ( .B1(P2_REG2_REG_17__SCAN_IN), .B2(n8605), .A(n8640), .ZN(
        n8618) );
  OR3_X1 U10189 ( .A1(n8608), .A2(n8607), .A3(n8606), .ZN(n8609) );
  AOI21_X1 U10190 ( .B1(n8610), .B2(n8609), .A(n8626), .ZN(n8617) );
  NAND2_X1 U10191 ( .A1(n8611), .A2(P2_ADDR_REG_17__SCAN_IN), .ZN(n8613) );
  OAI211_X1 U10192 ( .C1(n8615), .C2(n8614), .A(n8613), .B(n8612), .ZN(n8616)
         );
  AOI211_X1 U10193 ( .C1(n8618), .C2(n8641), .A(n8617), .B(n8616), .ZN(n8619)
         );
  OAI21_X1 U10194 ( .B1(n8620), .B2(n8645), .A(n8619), .ZN(P2_U3199) );
  XOR2_X1 U10195 ( .A(n8622), .B(n8621), .Z(n8646) );
  INV_X1 U10196 ( .A(n8628), .ZN(n8625) );
  NOR3_X1 U10197 ( .A1(n8625), .A2(n8624), .A3(n8623), .ZN(n8637) );
  AOI21_X1 U10198 ( .B1(n8628), .B2(n8627), .A(n8626), .ZN(n8630) );
  INV_X1 U10199 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n8633) );
  OAI21_X1 U10200 ( .B1(n8634), .B2(n8633), .A(n8632), .ZN(n8635) );
  AND3_X1 U10201 ( .A1(n8640), .A2(n8639), .A3(n8638), .ZN(n8642) );
  OAI21_X1 U10202 ( .B1(n8643), .B2(n8642), .A(n8641), .ZN(n8644) );
  AOI21_X1 U10203 ( .B1(n9150), .B2(n10171), .A(n8649), .ZN(n8652) );
  NAND2_X1 U10204 ( .A1(n10174), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n8650) );
  OAI211_X1 U10205 ( .C1(n9152), .C2(n8784), .A(n8652), .B(n8650), .ZN(
        P2_U3202) );
  NAND2_X1 U10206 ( .A1(n10174), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n8651) );
  OAI211_X1 U10207 ( .C1(n8928), .C2(n8784), .A(n8652), .B(n8651), .ZN(
        P2_U3203) );
  INV_X1 U10208 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n8661) );
  XNOR2_X1 U10209 ( .A(n8654), .B(n8655), .ZN(n8660) );
  MUX2_X1 U10210 ( .A(n8661), .B(n9157), .S(n10171), .Z(n8664) );
  AOI22_X1 U10211 ( .A1(n9159), .A2(n8921), .B1(n8920), .B2(n8662), .ZN(n8663)
         );
  OAI211_X1 U10212 ( .C1(n9162), .C2(n8855), .A(n8664), .B(n8663), .ZN(
        P2_U3205) );
  XNOR2_X1 U10213 ( .A(n8666), .B(n8665), .ZN(n9168) );
  INV_X1 U10214 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n8678) );
  NAND2_X1 U10215 ( .A1(n8670), .A2(n8669), .ZN(n8672) );
  MUX2_X1 U10216 ( .A(n8678), .B(n9163), .S(n10171), .Z(n8681) );
  AOI22_X1 U10217 ( .A1(n9165), .A2(n8921), .B1(n8920), .B2(n8679), .ZN(n8680)
         );
  OAI211_X1 U10218 ( .C1(n9168), .C2(n8855), .A(n8681), .B(n8680), .ZN(
        P2_U3206) );
  XNOR2_X1 U10219 ( .A(n8682), .B(n8684), .ZN(n9174) );
  INV_X1 U10220 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n8692) );
  NAND2_X1 U10221 ( .A1(n8696), .A2(n8683), .ZN(n8685) );
  MUX2_X1 U10222 ( .A(n8692), .B(n9169), .S(n10171), .Z(n8695) );
  AOI22_X1 U10223 ( .A1(n9171), .A2(n8921), .B1(n8920), .B2(n8693), .ZN(n8694)
         );
  OAI211_X1 U10224 ( .C1(n9174), .C2(n8855), .A(n8695), .B(n8694), .ZN(
        P2_U3207) );
  INV_X1 U10225 ( .A(n9178), .ZN(n8941) );
  NOR2_X1 U10226 ( .A1(n8941), .A2(n10163), .ZN(n8703) );
  INV_X1 U10227 ( .A(n8667), .ZN(n8698) );
  INV_X1 U10228 ( .A(n8705), .ZN(n8697) );
  OAI211_X1 U10229 ( .C1(n8698), .C2(n8697), .A(n8887), .B(n8696), .ZN(n8701)
         );
  NAND2_X1 U10230 ( .A1(n8699), .A2(n8917), .ZN(n8700) );
  AOI211_X1 U10231 ( .C1(n8920), .C2(n8704), .A(n8703), .B(n9175), .ZN(n8708)
         );
  XNOR2_X1 U10232 ( .A(n8706), .B(n8705), .ZN(n8940) );
  INV_X1 U10233 ( .A(n8855), .ZN(n8786) );
  AOI22_X1 U10234 ( .A1(n8940), .A2(n8786), .B1(P2_REG2_REG_25__SCAN_IN), .B2(
        n10174), .ZN(n8707) );
  OAI21_X1 U10235 ( .B1(n8708), .B2(n10174), .A(n8707), .ZN(P2_U3208) );
  NOR2_X1 U10236 ( .A1(n8945), .A2(n10163), .ZN(n8713) );
  XOR2_X1 U10237 ( .A(n8717), .B(n8709), .Z(n8710) );
  OAI222_X1 U10238 ( .A1(n8905), .A2(n8712), .B1(n8848), .B2(n8711), .C1(n8710), .C2(n8911), .ZN(n9182) );
  AOI211_X1 U10239 ( .C1(n8920), .C2(n8714), .A(n8713), .B(n9182), .ZN(n8720)
         );
  NAND2_X1 U10240 ( .A1(n8716), .A2(n8715), .ZN(n8718) );
  XNOR2_X1 U10241 ( .A(n8718), .B(n8717), .ZN(n8944) );
  AOI22_X1 U10242 ( .A1(n8944), .A2(n8786), .B1(P2_REG2_REG_24__SCAN_IN), .B2(
        n10174), .ZN(n8719) );
  OAI21_X1 U10243 ( .B1(n8720), .B2(n10174), .A(n8719), .ZN(P2_U3209) );
  XOR2_X1 U10244 ( .A(n8721), .B(n8723), .Z(n9194) );
  INV_X1 U10245 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n8727) );
  XOR2_X1 U10246 ( .A(n8723), .B(n8722), .Z(n8726) );
  AOI222_X1 U10247 ( .A1(n8887), .A2(n8726), .B1(n8725), .B2(n8917), .C1(n8724), .C2(n8890), .ZN(n9189) );
  MUX2_X1 U10248 ( .A(n8727), .B(n9189), .S(n10171), .Z(n8730) );
  AOI22_X1 U10249 ( .A1(n9191), .A2(n8921), .B1(n8920), .B2(n8728), .ZN(n8729)
         );
  OAI211_X1 U10250 ( .C1(n9194), .C2(n8855), .A(n8730), .B(n8729), .ZN(
        P2_U3210) );
  XOR2_X1 U10251 ( .A(n8731), .B(n8733), .Z(n9200) );
  XNOR2_X1 U10252 ( .A(n8732), .B(n8733), .ZN(n8735) );
  AOI222_X1 U10253 ( .A1(n8887), .A2(n8735), .B1(n8734), .B2(n8917), .C1(n8758), .C2(n8890), .ZN(n9195) );
  OAI21_X1 U10254 ( .B1(n8736), .B2(n10165), .A(n9195), .ZN(n8737) );
  NAND2_X1 U10255 ( .A1(n8737), .A2(n10171), .ZN(n8739) );
  AOI22_X1 U10256 ( .A1(n9197), .A2(n8921), .B1(P2_REG2_REG_22__SCAN_IN), .B2(
        n10174), .ZN(n8738) );
  OAI211_X1 U10257 ( .C1(n9200), .C2(n8855), .A(n8739), .B(n8738), .ZN(
        P2_U3211) );
  XNOR2_X1 U10258 ( .A(n8740), .B(n8744), .ZN(n9204) );
  AOI21_X1 U10259 ( .B1(n8741), .B2(n8743), .A(n8742), .ZN(n8745) );
  XNOR2_X1 U10260 ( .A(n8745), .B(n8744), .ZN(n8746) );
  OAI222_X1 U10261 ( .A1(n8848), .A2(n8747), .B1(n8905), .B2(n8769), .C1(n8911), .C2(n8746), .ZN(n8953) );
  NAND2_X1 U10262 ( .A1(n8953), .A2(n10171), .ZN(n8752) );
  INV_X1 U10263 ( .A(n8748), .ZN(n8749) );
  OAI22_X1 U10264 ( .A1(n8749), .A2(n10165), .B1(n10171), .B2(n9062), .ZN(
        n8750) );
  AOI21_X1 U10265 ( .B1(n8954), .B2(n8921), .A(n8750), .ZN(n8751) );
  OAI211_X1 U10266 ( .C1(n9204), .C2(n8855), .A(n8752), .B(n8751), .ZN(
        P2_U3212) );
  XOR2_X1 U10267 ( .A(n8755), .B(n8753), .Z(n9210) );
  INV_X1 U10268 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n8760) );
  NOR2_X1 U10269 ( .A1(n8741), .A2(n8767), .ZN(n8766) );
  NOR2_X1 U10270 ( .A1(n8766), .A2(n8754), .ZN(n8756) );
  XNOR2_X1 U10271 ( .A(n8756), .B(n8755), .ZN(n8759) );
  AOI222_X1 U10272 ( .A1(n8887), .A2(n8759), .B1(n8758), .B2(n8917), .C1(n8757), .C2(n8890), .ZN(n9205) );
  MUX2_X1 U10273 ( .A(n8760), .B(n9205), .S(n10171), .Z(n8763) );
  AOI22_X1 U10274 ( .A1(n9207), .A2(n8921), .B1(n8920), .B2(n8761), .ZN(n8762)
         );
  OAI211_X1 U10275 ( .C1(n9210), .C2(n8855), .A(n8763), .B(n8762), .ZN(
        P2_U3213) );
  XNOR2_X1 U10276 ( .A(n8765), .B(n8764), .ZN(n9216) );
  INV_X1 U10277 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n8772) );
  AOI211_X1 U10278 ( .C1(n8767), .C2(n8741), .A(n8911), .B(n8766), .ZN(n8771)
         );
  OAI22_X1 U10279 ( .A1(n8769), .A2(n8848), .B1(n8768), .B2(n8905), .ZN(n8770)
         );
  NOR2_X1 U10280 ( .A1(n8771), .A2(n8770), .ZN(n9211) );
  MUX2_X1 U10281 ( .A(n8772), .B(n9211), .S(n10171), .Z(n8775) );
  AOI22_X1 U10282 ( .A1(n9213), .A2(n8921), .B1(n8920), .B2(n8773), .ZN(n8774)
         );
  OAI211_X1 U10283 ( .C1(n9216), .C2(n8855), .A(n8775), .B(n8774), .ZN(
        P2_U3214) );
  XOR2_X1 U10284 ( .A(n8776), .B(n8781), .Z(n8777) );
  OAI222_X1 U10285 ( .A1(n8848), .A2(n8779), .B1(n8905), .B2(n8778), .C1(n8777), .C2(n8911), .ZN(n8963) );
  INV_X1 U10286 ( .A(n8963), .ZN(n8788) );
  XOR2_X1 U10287 ( .A(n8781), .B(n8780), .Z(n8964) );
  AOI22_X1 U10288 ( .A1(n10174), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n8920), 
        .B2(n8782), .ZN(n8783) );
  OAI21_X1 U10289 ( .B1(n9220), .B2(n8784), .A(n8783), .ZN(n8785) );
  AOI21_X1 U10290 ( .B1(n8964), .B2(n8786), .A(n8785), .ZN(n8787) );
  OAI21_X1 U10291 ( .B1(n8788), .B2(n10174), .A(n8787), .ZN(P2_U3215) );
  XNOR2_X1 U10292 ( .A(n8790), .B(n8789), .ZN(n9226) );
  INV_X1 U10293 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8795) );
  XNOR2_X1 U10294 ( .A(n8791), .B(n8792), .ZN(n8794) );
  AOI222_X1 U10295 ( .A1(n8887), .A2(n8794), .B1(n8793), .B2(n8917), .C1(n8811), .C2(n8890), .ZN(n9221) );
  MUX2_X1 U10296 ( .A(n8795), .B(n9221), .S(n10171), .Z(n8798) );
  AOI22_X1 U10297 ( .A1(n9223), .A2(n8921), .B1(n8920), .B2(n8796), .ZN(n8797)
         );
  OAI211_X1 U10298 ( .C1(n9226), .C2(n8855), .A(n8798), .B(n8797), .ZN(
        P2_U3216) );
  XNOR2_X1 U10299 ( .A(n4470), .B(n8800), .ZN(n9232) );
  XOR2_X1 U10300 ( .A(n8801), .B(n8800), .Z(n8803) );
  AOI222_X1 U10301 ( .A1(n8887), .A2(n8803), .B1(n8802), .B2(n8917), .C1(n8818), .C2(n8890), .ZN(n9227) );
  MUX2_X1 U10302 ( .A(n8804), .B(n9227), .S(n10171), .Z(n8807) );
  AOI22_X1 U10303 ( .A1(n9229), .A2(n8921), .B1(n8920), .B2(n8805), .ZN(n8806)
         );
  OAI211_X1 U10304 ( .C1(n9232), .C2(n8855), .A(n8807), .B(n8806), .ZN(
        P2_U3217) );
  XNOR2_X1 U10305 ( .A(n8808), .B(n8809), .ZN(n9238) );
  XNOR2_X1 U10306 ( .A(n8810), .B(n8809), .ZN(n8812) );
  AOI222_X1 U10307 ( .A1(n8887), .A2(n8812), .B1(n8811), .B2(n8917), .C1(n8830), .C2(n8890), .ZN(n9233) );
  MUX2_X1 U10308 ( .A(n8813), .B(n9233), .S(n10171), .Z(n8816) );
  AOI22_X1 U10309 ( .A1(n9235), .A2(n8921), .B1(n8920), .B2(n8814), .ZN(n8815)
         );
  OAI211_X1 U10310 ( .C1(n9238), .C2(n8855), .A(n8816), .B(n8815), .ZN(
        P2_U3218) );
  XNOR2_X1 U10311 ( .A(n8817), .B(n8823), .ZN(n8820) );
  AOI222_X1 U10312 ( .A1(n8887), .A2(n8820), .B1(n8819), .B2(n8890), .C1(n8818), .C2(n8917), .ZN(n9239) );
  AOI22_X1 U10313 ( .A1(n9241), .A2(n8833), .B1(n8920), .B2(n8821), .ZN(n8822)
         );
  AOI21_X1 U10314 ( .B1(n9239), .B2(n8822), .A(n10174), .ZN(n8827) );
  XNOR2_X1 U10315 ( .A(n8824), .B(n8823), .ZN(n9244) );
  OAI22_X1 U10316 ( .A1(n9244), .A2(n8855), .B1(n8825), .B2(n10171), .ZN(n8826) );
  OR2_X1 U10317 ( .A1(n8827), .A2(n8826), .ZN(P2_U3219) );
  XOR2_X1 U10318 ( .A(n8828), .B(n8835), .Z(n8831) );
  AOI222_X1 U10319 ( .A1(n8887), .A2(n8831), .B1(n8830), .B2(n8917), .C1(n8829), .C2(n8890), .ZN(n9245) );
  AOI22_X1 U10320 ( .A1(n9248), .A2(n8833), .B1(n8920), .B2(n8832), .ZN(n8834)
         );
  AOI21_X1 U10321 ( .B1(n9245), .B2(n8834), .A(n10174), .ZN(n8839) );
  XNOR2_X1 U10322 ( .A(n8836), .B(n8835), .ZN(n9251) );
  OAI22_X1 U10323 ( .A1(n9251), .A2(n8855), .B1(n8837), .B2(n10171), .ZN(n8838) );
  OR2_X1 U10324 ( .A1(n8839), .A2(n8838), .ZN(P2_U3220) );
  NAND2_X1 U10325 ( .A1(n8840), .A2(n8841), .ZN(n8842) );
  NAND2_X1 U10326 ( .A1(n8843), .A2(n8842), .ZN(n9256) );
  XNOR2_X1 U10327 ( .A(n8844), .B(n6630), .ZN(n8845) );
  OAI222_X1 U10328 ( .A1(n8848), .A2(n8847), .B1(n8905), .B2(n8846), .C1(n8911), .C2(n8845), .ZN(n8982) );
  NAND2_X1 U10329 ( .A1(n8982), .A2(n10171), .ZN(n8854) );
  INV_X1 U10330 ( .A(n8849), .ZN(n8850) );
  OAI22_X1 U10331 ( .A1(n10171), .A2(n8851), .B1(n8850), .B2(n10165), .ZN(
        n8852) );
  AOI21_X1 U10332 ( .B1(n6663), .B2(n8921), .A(n8852), .ZN(n8853) );
  OAI211_X1 U10333 ( .C1(n9256), .C2(n8855), .A(n8854), .B(n8853), .ZN(
        P2_U3221) );
  INV_X1 U10334 ( .A(n8879), .ZN(n8858) );
  INV_X1 U10335 ( .A(n8856), .ZN(n8857) );
  OAI21_X1 U10336 ( .B1(n8859), .B2(n8858), .A(n8857), .ZN(n8880) );
  NAND2_X1 U10337 ( .A1(n8880), .A2(n8860), .ZN(n8861) );
  XOR2_X1 U10338 ( .A(n8867), .B(n8861), .Z(n8986) );
  INV_X1 U10339 ( .A(n8883), .ZN(n8863) );
  AOI21_X1 U10340 ( .B1(n7385), .B2(n8863), .A(n8862), .ZN(n8865) );
  NOR2_X1 U10341 ( .A1(n8865), .A2(n8864), .ZN(n8866) );
  XOR2_X1 U10342 ( .A(n8867), .B(n8866), .Z(n8868) );
  NAND2_X1 U10343 ( .A1(n8868), .A2(n8887), .ZN(n8871) );
  AOI22_X1 U10344 ( .A1(n8869), .A2(n8917), .B1(n8890), .B2(n8916), .ZN(n8870)
         );
  OAI211_X1 U10345 ( .C1(n8986), .C2(n8894), .A(n8871), .B(n8870), .ZN(n8987)
         );
  INV_X1 U10346 ( .A(n8987), .ZN(n8872) );
  MUX2_X1 U10347 ( .A(n8873), .B(n8872), .S(n10171), .Z(n8877) );
  AOI22_X1 U10348 ( .A1(n8921), .A2(n8875), .B1(n8920), .B2(n8874), .ZN(n8876)
         );
  OAI211_X1 U10349 ( .C1(n8986), .C2(n8901), .A(n8877), .B(n8876), .ZN(
        P2_U3223) );
  AOI21_X1 U10350 ( .B1(n8903), .B2(n8879), .A(n8878), .ZN(n8882) );
  OAI21_X1 U10351 ( .B1(n8882), .B2(n8881), .A(n8880), .ZN(n8990) );
  NOR2_X1 U10352 ( .A1(n8907), .A2(n8883), .ZN(n8912) );
  NOR2_X1 U10353 ( .A1(n8912), .A2(n8884), .ZN(n8886) );
  XNOR2_X1 U10354 ( .A(n8886), .B(n8885), .ZN(n8888) );
  NAND2_X1 U10355 ( .A1(n8888), .A2(n8887), .ZN(n8893) );
  AOI22_X1 U10356 ( .A1(n8891), .A2(n8890), .B1(n8917), .B2(n8889), .ZN(n8892)
         );
  OAI211_X1 U10357 ( .C1(n8990), .C2(n8894), .A(n8893), .B(n8892), .ZN(n8991)
         );
  INV_X1 U10358 ( .A(n8991), .ZN(n8895) );
  MUX2_X1 U10359 ( .A(n8896), .B(n8895), .S(n10171), .Z(n8900) );
  AOI22_X1 U10360 ( .A1(n8921), .A2(n8898), .B1(n8920), .B2(n8897), .ZN(n8899)
         );
  OAI211_X1 U10361 ( .C1(n8990), .C2(n8901), .A(n8900), .B(n8899), .ZN(
        P2_U3224) );
  NAND2_X1 U10362 ( .A1(n8903), .A2(n8902), .ZN(n8904) );
  XNOR2_X1 U10363 ( .A(n8904), .B(n8908), .ZN(n9000) );
  INV_X1 U10364 ( .A(n9000), .ZN(n8924) );
  NOR2_X1 U10365 ( .A1(n8906), .A2(n8905), .ZN(n8915) );
  INV_X1 U10366 ( .A(n8907), .ZN(n8910) );
  AOI21_X1 U10367 ( .B1(n8910), .B2(n8909), .A(n8908), .ZN(n8913) );
  NOR3_X1 U10368 ( .A1(n8913), .A2(n8912), .A3(n8911), .ZN(n8914) );
  AOI211_X1 U10369 ( .C1(n8917), .C2(n8916), .A(n8915), .B(n8914), .ZN(n9002)
         );
  MUX2_X1 U10370 ( .A(n8918), .B(n9002), .S(n10171), .Z(n8923) );
  AOI22_X1 U10371 ( .A1(n8921), .A2(n8997), .B1(n8920), .B2(n8919), .ZN(n8922)
         );
  OAI211_X1 U10372 ( .C1(n8924), .C2(n8855), .A(n8923), .B(n8922), .ZN(
        P2_U3225) );
  NAND2_X1 U10373 ( .A1(n9150), .A2(n9003), .ZN(n8926) );
  NAND2_X1 U10374 ( .A1(n4269), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n8925) );
  OAI211_X1 U10375 ( .C1(n9152), .C2(n8996), .A(n8926), .B(n8925), .ZN(
        P2_U3490) );
  NAND2_X1 U10376 ( .A1(n4269), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n8927) );
  OAI211_X1 U10377 ( .C1(n8928), .C2(n8996), .A(n8927), .B(n8926), .ZN(
        P2_U3489) );
  INV_X1 U10378 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n8929) );
  NAND2_X1 U10379 ( .A1(n9159), .A2(n8979), .ZN(n8932) );
  OAI211_X1 U10380 ( .C1(n9162), .C2(n8985), .A(n8933), .B(n8932), .ZN(
        P2_U3487) );
  INV_X1 U10381 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n8934) );
  MUX2_X1 U10382 ( .A(n8934), .B(n9163), .S(n9003), .Z(n8936) );
  NAND2_X1 U10383 ( .A1(n9165), .A2(n8979), .ZN(n8935) );
  OAI211_X1 U10384 ( .C1(n9168), .C2(n8985), .A(n8936), .B(n8935), .ZN(
        P2_U3486) );
  INV_X1 U10385 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n8937) );
  MUX2_X1 U10386 ( .A(n8937), .B(n9169), .S(n9003), .Z(n8939) );
  NAND2_X1 U10387 ( .A1(n9171), .A2(n8979), .ZN(n8938) );
  OAI211_X1 U10388 ( .C1(n8985), .C2(n9174), .A(n8939), .B(n8938), .ZN(
        P2_U3485) );
  INV_X1 U10389 ( .A(n8940), .ZN(n9181) );
  OAI22_X1 U10390 ( .A1(n9181), .A2(n8985), .B1(n8941), .B2(n8996), .ZN(n8942)
         );
  OR2_X1 U10391 ( .A1(n8943), .A2(n8942), .ZN(P2_U3484) );
  MUX2_X1 U10392 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n9182), .S(n9003), .Z(n8947) );
  INV_X1 U10393 ( .A(n8944), .ZN(n9188) );
  OAI22_X1 U10394 ( .A1(n9188), .A2(n8985), .B1(n8945), .B2(n8996), .ZN(n8946)
         );
  OR2_X1 U10395 ( .A1(n8947), .A2(n8946), .ZN(P2_U3483) );
  INV_X1 U10396 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n8948) );
  MUX2_X1 U10397 ( .A(n8948), .B(n9189), .S(n9003), .Z(n8950) );
  NAND2_X1 U10398 ( .A1(n9191), .A2(n8979), .ZN(n8949) );
  OAI211_X1 U10399 ( .C1(n9194), .C2(n8985), .A(n8950), .B(n8949), .ZN(
        P2_U3482) );
  MUX2_X1 U10400 ( .A(n9094), .B(n9195), .S(n9003), .Z(n8952) );
  NAND2_X1 U10401 ( .A1(n9197), .A2(n8979), .ZN(n8951) );
  OAI211_X1 U10402 ( .C1(n9200), .C2(n8985), .A(n8952), .B(n8951), .ZN(
        P2_U3481) );
  INV_X1 U10403 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n8955) );
  AOI21_X1 U10404 ( .B1(n8998), .B2(n8954), .A(n8953), .ZN(n9201) );
  MUX2_X1 U10405 ( .A(n8955), .B(n9201), .S(n9003), .Z(n8956) );
  OAI21_X1 U10406 ( .B1(n8985), .B2(n9204), .A(n8956), .ZN(P2_U3480) );
  INV_X1 U10407 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n8957) );
  MUX2_X1 U10408 ( .A(n8957), .B(n9205), .S(n9003), .Z(n8959) );
  NAND2_X1 U10409 ( .A1(n9207), .A2(n8979), .ZN(n8958) );
  OAI211_X1 U10410 ( .C1(n8985), .C2(n9210), .A(n8959), .B(n8958), .ZN(
        P2_U3479) );
  MUX2_X1 U10411 ( .A(n8960), .B(n9211), .S(n9003), .Z(n8962) );
  NAND2_X1 U10412 ( .A1(n9213), .A2(n8979), .ZN(n8961) );
  OAI211_X1 U10413 ( .C1(n9216), .C2(n8985), .A(n8962), .B(n8961), .ZN(
        P2_U3478) );
  AOI21_X1 U10414 ( .B1(n8999), .B2(n8964), .A(n8963), .ZN(n9217) );
  MUX2_X1 U10415 ( .A(n8965), .B(n9217), .S(n9003), .Z(n8966) );
  OAI21_X1 U10416 ( .B1(n9220), .B2(n8996), .A(n8966), .ZN(P2_U3477) );
  MUX2_X1 U10417 ( .A(n8967), .B(n9221), .S(n9003), .Z(n8969) );
  NAND2_X1 U10418 ( .A1(n9223), .A2(n8979), .ZN(n8968) );
  OAI211_X1 U10419 ( .C1(n9226), .C2(n8985), .A(n8969), .B(n8968), .ZN(
        P2_U3476) );
  MUX2_X1 U10420 ( .A(n8970), .B(n9227), .S(n9003), .Z(n8972) );
  NAND2_X1 U10421 ( .A1(n9229), .A2(n8979), .ZN(n8971) );
  OAI211_X1 U10422 ( .C1(n8985), .C2(n9232), .A(n8972), .B(n8971), .ZN(
        P2_U3475) );
  MUX2_X1 U10423 ( .A(n8973), .B(n9233), .S(n9003), .Z(n8975) );
  NAND2_X1 U10424 ( .A1(n9235), .A2(n8979), .ZN(n8974) );
  OAI211_X1 U10425 ( .C1(n8985), .C2(n9238), .A(n8975), .B(n8974), .ZN(
        P2_U3474) );
  MUX2_X1 U10426 ( .A(n8976), .B(n9239), .S(n9003), .Z(n8978) );
  NAND2_X1 U10427 ( .A1(n9241), .A2(n8979), .ZN(n8977) );
  OAI211_X1 U10428 ( .C1(n8985), .C2(n9244), .A(n8978), .B(n8977), .ZN(
        P2_U3473) );
  MUX2_X1 U10429 ( .A(n9021), .B(n9245), .S(n9003), .Z(n8981) );
  NAND2_X1 U10430 ( .A1(n9248), .A2(n8979), .ZN(n8980) );
  OAI211_X1 U10431 ( .C1(n8985), .C2(n9251), .A(n8981), .B(n8980), .ZN(
        P2_U3472) );
  AOI21_X1 U10432 ( .B1(n8998), .B2(n6663), .A(n8982), .ZN(n9252) );
  MUX2_X1 U10433 ( .A(n8983), .B(n9252), .S(n9003), .Z(n8984) );
  OAI21_X1 U10434 ( .B1(n8985), .B2(n9256), .A(n8984), .ZN(P2_U3471) );
  INV_X1 U10435 ( .A(n8986), .ZN(n8988) );
  AOI21_X1 U10436 ( .B1(n8993), .B2(n8988), .A(n8987), .ZN(n9257) );
  MUX2_X1 U10437 ( .A(n9024), .B(n9257), .S(n9003), .Z(n8989) );
  OAI21_X1 U10438 ( .B1(n9260), .B2(n8996), .A(n8989), .ZN(P2_U3469) );
  INV_X1 U10439 ( .A(n8990), .ZN(n8992) );
  AOI21_X1 U10440 ( .B1(n8993), .B2(n8992), .A(n8991), .ZN(n9261) );
  MUX2_X1 U10441 ( .A(n8994), .B(n9261), .S(n9003), .Z(n8995) );
  OAI21_X1 U10442 ( .B1(n9265), .B2(n8996), .A(n8995), .ZN(P2_U3468) );
  AOI22_X1 U10443 ( .A1(n9000), .A2(n8999), .B1(n8998), .B2(n8997), .ZN(n9001)
         );
  NAND2_X1 U10444 ( .A1(n9002), .A2(n9001), .ZN(n9266) );
  MUX2_X1 U10445 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n9266), .S(n9003), .Z(n9147)
         );
  AOI22_X1 U10446 ( .A1(n9005), .A2(keyinput27), .B1(n9115), .B2(keyinput39), 
        .ZN(n9004) );
  OAI221_X1 U10447 ( .B1(n9005), .B2(keyinput27), .C1(n9115), .C2(keyinput39), 
        .A(n9004), .ZN(n9019) );
  AOI22_X1 U10448 ( .A1(n9008), .A2(keyinput46), .B1(n9007), .B2(keyinput5), 
        .ZN(n9006) );
  OAI221_X1 U10449 ( .B1(n9008), .B2(keyinput46), .C1(n9007), .C2(keyinput5), 
        .A(n9006), .ZN(n9018) );
  INV_X1 U10450 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n10187) );
  XOR2_X1 U10451 ( .A(n10187), .B(keyinput13), .Z(n9011) );
  XNOR2_X1 U10452 ( .A(P1_IR_REG_17__SCAN_IN), .B(keyinput51), .ZN(n9010) );
  XNOR2_X1 U10453 ( .A(P1_IR_REG_20__SCAN_IN), .B(keyinput0), .ZN(n9009) );
  NAND3_X1 U10454 ( .A1(n9011), .A2(n9010), .A3(n9009), .ZN(n9017) );
  XNOR2_X1 U10455 ( .A(P1_IR_REG_19__SCAN_IN), .B(keyinput45), .ZN(n9015) );
  XNOR2_X1 U10456 ( .A(P2_IR_REG_2__SCAN_IN), .B(keyinput12), .ZN(n9014) );
  XNOR2_X1 U10457 ( .A(P1_ADDR_REG_19__SCAN_IN), .B(keyinput60), .ZN(n9013) );
  XNOR2_X1 U10458 ( .A(P2_REG0_REG_12__SCAN_IN), .B(keyinput32), .ZN(n9012) );
  NAND4_X1 U10459 ( .A1(n9015), .A2(n9014), .A3(n9013), .A4(n9012), .ZN(n9016)
         );
  NOR4_X1 U10460 ( .A1(n9019), .A2(n9018), .A3(n9017), .A4(n9016), .ZN(n9058)
         );
  AOI22_X1 U10461 ( .A1(n9022), .A2(keyinput62), .B1(keyinput9), .B2(n9021), 
        .ZN(n9020) );
  OAI221_X1 U10462 ( .B1(n9022), .B2(keyinput62), .C1(n9021), .C2(keyinput9), 
        .A(n9020), .ZN(n9028) );
  AOI22_X1 U10463 ( .A1(n9113), .A2(keyinput2), .B1(keyinput49), .B2(n9024), 
        .ZN(n9023) );
  OAI221_X1 U10464 ( .B1(n9113), .B2(keyinput2), .C1(n9024), .C2(keyinput49), 
        .A(n9023), .ZN(n9027) );
  XNOR2_X1 U10465 ( .A(n9025), .B(keyinput53), .ZN(n9026) );
  NOR3_X1 U10466 ( .A1(n9028), .A2(n9027), .A3(n9026), .ZN(n9057) );
  INV_X1 U10467 ( .A(SI_14_), .ZN(n9030) );
  AOI22_X1 U10468 ( .A1(n9030), .A2(keyinput33), .B1(keyinput21), .B2(n9114), 
        .ZN(n9029) );
  OAI221_X1 U10469 ( .B1(n9030), .B2(keyinput33), .C1(n9114), .C2(keyinput21), 
        .A(n9029), .ZN(n9036) );
  AOI22_X1 U10470 ( .A1(n9702), .A2(keyinput28), .B1(n9032), .B2(keyinput56), 
        .ZN(n9031) );
  OAI221_X1 U10471 ( .B1(n9702), .B2(keyinput28), .C1(n9032), .C2(keyinput56), 
        .A(n9031), .ZN(n9035) );
  XNOR2_X1 U10472 ( .A(n9033), .B(keyinput17), .ZN(n9034) );
  NOR3_X1 U10473 ( .A1(n9036), .A2(n9035), .A3(n9034), .ZN(n9056) );
  AOI22_X1 U10474 ( .A1(n7589), .A2(keyinput59), .B1(n9038), .B2(keyinput58), 
        .ZN(n9037) );
  OAI221_X1 U10475 ( .B1(n7589), .B2(keyinput59), .C1(n9038), .C2(keyinput58), 
        .A(n9037), .ZN(n9054) );
  XOR2_X1 U10476 ( .A(n7046), .B(keyinput26), .Z(n9042) );
  XNOR2_X1 U10477 ( .A(P1_IR_REG_14__SCAN_IN), .B(keyinput37), .ZN(n9041) );
  XNOR2_X1 U10478 ( .A(P1_REG0_REG_18__SCAN_IN), .B(keyinput6), .ZN(n9040) );
  XNOR2_X1 U10479 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(keyinput4), .ZN(n9039) );
  NAND4_X1 U10480 ( .A1(n9042), .A2(n9041), .A3(n9040), .A4(n9039), .ZN(n9053)
         );
  XNOR2_X1 U10481 ( .A(P2_REG0_REG_31__SCAN_IN), .B(keyinput30), .ZN(n9046) );
  XNOR2_X1 U10482 ( .A(n9109), .B(keyinput42), .ZN(n9045) );
  XNOR2_X1 U10483 ( .A(P1_REG3_REG_7__SCAN_IN), .B(keyinput47), .ZN(n9044) );
  XNOR2_X1 U10484 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(keyinput19), .ZN(n9043)
         );
  NAND4_X1 U10485 ( .A1(n9046), .A2(n9045), .A3(n9044), .A4(n9043), .ZN(n9052)
         );
  XNOR2_X1 U10486 ( .A(P1_IR_REG_24__SCAN_IN), .B(keyinput29), .ZN(n9050) );
  XNOR2_X1 U10487 ( .A(P1_IR_REG_7__SCAN_IN), .B(keyinput55), .ZN(n9049) );
  XNOR2_X1 U10488 ( .A(P1_REG3_REG_15__SCAN_IN), .B(keyinput24), .ZN(n9048) );
  XNOR2_X1 U10489 ( .A(P1_IR_REG_31__SCAN_IN), .B(keyinput10), .ZN(n9047) );
  NAND4_X1 U10490 ( .A1(n9050), .A2(n9049), .A3(n9048), .A4(n9047), .ZN(n9051)
         );
  NOR4_X1 U10491 ( .A1(n9054), .A2(n9053), .A3(n9052), .A4(n9051), .ZN(n9055)
         );
  AND4_X1 U10492 ( .A1(n9058), .A2(n9057), .A3(n9056), .A4(n9055), .ZN(n9090)
         );
  INV_X1 U10493 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n10176) );
  INV_X1 U10494 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n10075) );
  AOI22_X1 U10495 ( .A1(n10176), .A2(keyinput8), .B1(n10075), .B2(keyinput16), 
        .ZN(n9059) );
  OAI221_X1 U10496 ( .B1(n10176), .B2(keyinput8), .C1(n10075), .C2(keyinput16), 
        .A(n9059), .ZN(n9068) );
  AOI22_X1 U10497 ( .A1(n9062), .A2(keyinput22), .B1(n9061), .B2(keyinput14), 
        .ZN(n9060) );
  OAI221_X1 U10498 ( .B1(n9062), .B2(keyinput22), .C1(n9061), .C2(keyinput14), 
        .A(n9060), .ZN(n9067) );
  INV_X1 U10499 ( .A(P1_D_REG_28__SCAN_IN), .ZN(n10072) );
  AOI22_X1 U10500 ( .A1(n9105), .A2(keyinput50), .B1(n10072), .B2(keyinput31), 
        .ZN(n9063) );
  OAI221_X1 U10501 ( .B1(n9105), .B2(keyinput50), .C1(n10072), .C2(keyinput31), 
        .A(n9063), .ZN(n9066) );
  AOI22_X1 U10502 ( .A1(n9952), .A2(keyinput57), .B1(n5953), .B2(keyinput18), 
        .ZN(n9064) );
  OAI221_X1 U10503 ( .B1(n9952), .B2(keyinput57), .C1(n5953), .C2(keyinput18), 
        .A(n9064), .ZN(n9065) );
  NOR4_X1 U10504 ( .A1(n9068), .A2(n9067), .A3(n9066), .A4(n9065), .ZN(n9089)
         );
  INV_X1 U10505 ( .A(P1_D_REG_13__SCAN_IN), .ZN(n10073) );
  AOI22_X1 U10506 ( .A1(n5973), .A2(keyinput15), .B1(n10073), .B2(keyinput36), 
        .ZN(n9069) );
  OAI221_X1 U10507 ( .B1(n5973), .B2(keyinput15), .C1(n10073), .C2(keyinput36), 
        .A(n9069), .ZN(n9077) );
  AOI22_X1 U10508 ( .A1(n9072), .A2(keyinput54), .B1(keyinput52), .B2(n9071), 
        .ZN(n9070) );
  OAI221_X1 U10509 ( .B1(n9072), .B2(keyinput54), .C1(n9071), .C2(keyinput52), 
        .A(n9070), .ZN(n9076) );
  AOI22_X1 U10510 ( .A1(n9074), .A2(keyinput48), .B1(n9104), .B2(keyinput43), 
        .ZN(n9073) );
  OAI221_X1 U10511 ( .B1(n9074), .B2(keyinput48), .C1(n9104), .C2(keyinput43), 
        .A(n9073), .ZN(n9075) );
  NOR3_X1 U10512 ( .A1(n9077), .A2(n9076), .A3(n9075), .ZN(n9088) );
  AOI22_X1 U10513 ( .A1(n9137), .A2(keyinput20), .B1(keyinput7), .B2(n9079), 
        .ZN(n9078) );
  OAI221_X1 U10514 ( .B1(n9137), .B2(keyinput20), .C1(n9079), .C2(keyinput7), 
        .A(n9078), .ZN(n9086) );
  INV_X1 U10515 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n9246) );
  AOI22_X1 U10516 ( .A1(n9119), .A2(keyinput40), .B1(keyinput63), .B2(n9246), 
        .ZN(n9080) );
  OAI221_X1 U10517 ( .B1(n9119), .B2(keyinput40), .C1(n9246), .C2(keyinput63), 
        .A(n9080), .ZN(n9085) );
  INV_X1 U10518 ( .A(SI_12_), .ZN(n9083) );
  AOI22_X1 U10519 ( .A1(n9083), .A2(keyinput34), .B1(keyinput61), .B2(n9082), 
        .ZN(n9081) );
  OAI221_X1 U10520 ( .B1(n9083), .B2(keyinput34), .C1(n9082), .C2(keyinput61), 
        .A(n9081), .ZN(n9084) );
  NOR3_X1 U10521 ( .A1(n9086), .A2(n9085), .A3(n9084), .ZN(n9087) );
  AND4_X1 U10522 ( .A1(n9090), .A2(n9089), .A3(n9088), .A4(n9087), .ZN(n9145)
         );
  AOI22_X1 U10523 ( .A1(n9092), .A2(keyinput1), .B1(keyinput38), .B2(n9110), 
        .ZN(n9091) );
  OAI221_X1 U10524 ( .B1(n9092), .B2(keyinput1), .C1(n9110), .C2(keyinput38), 
        .A(n9091), .ZN(n9103) );
  AOI22_X1 U10525 ( .A1(n9095), .A2(keyinput11), .B1(keyinput3), .B2(n9094), 
        .ZN(n9093) );
  OAI221_X1 U10526 ( .B1(n9095), .B2(keyinput11), .C1(n9094), .C2(keyinput3), 
        .A(n9093), .ZN(n9102) );
  AOI22_X1 U10527 ( .A1(n5123), .A2(keyinput35), .B1(n9097), .B2(keyinput25), 
        .ZN(n9096) );
  OAI221_X1 U10528 ( .B1(n5123), .B2(keyinput35), .C1(n9097), .C2(keyinput25), 
        .A(n9096), .ZN(n9101) );
  AOI22_X1 U10529 ( .A1(n9118), .A2(keyinput41), .B1(keyinput44), .B2(n9099), 
        .ZN(n9098) );
  OAI221_X1 U10530 ( .B1(n9118), .B2(keyinput41), .C1(n9099), .C2(keyinput44), 
        .A(n9098), .ZN(n9100) );
  NOR4_X1 U10531 ( .A1(n9103), .A2(n9102), .A3(n9101), .A4(n9100), .ZN(n9144)
         );
  NOR4_X1 U10532 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_REG0_REG_28__SCAN_IN), 
        .A3(n9104), .A4(n7046), .ZN(n9106) );
  NAND4_X1 U10533 ( .A1(n9107), .A2(P1_ADDR_REG_6__SCAN_IN), .A3(n9106), .A4(
        n9105), .ZN(n9136) );
  NOR4_X1 U10534 ( .A1(n9108), .A2(P1_IR_REG_14__SCAN_IN), .A3(
        P1_REG3_REG_12__SCAN_IN), .A4(P1_REG3_REG_7__SCAN_IN), .ZN(n9127) );
  INV_X1 U10535 ( .A(n9109), .ZN(n9125) );
  NAND4_X1 U10536 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P2_DATAO_REG_16__SCAN_IN), 
        .A3(P2_REG1_REG_13__SCAN_IN), .A4(P2_REG1_REG_10__SCAN_IN), .ZN(n9112)
         );
  NAND4_X1 U10537 ( .A1(P2_REG1_REG_22__SCAN_IN), .A2(P1_REG0_REG_20__SCAN_IN), 
        .A3(n9110), .A4(n5123), .ZN(n9111) );
  NOR2_X1 U10538 ( .A1(n9112), .A2(n9111), .ZN(n9123) );
  NAND4_X1 U10539 ( .A1(P1_REG3_REG_22__SCAN_IN), .A2(n7589), .A3(n9114), .A4(
        n9113), .ZN(n9117) );
  NAND4_X1 U10540 ( .A1(P1_REG2_REG_21__SCAN_IN), .A2(P2_REG0_REG_13__SCAN_IN), 
        .A3(P2_REG1_REG_1__SCAN_IN), .A4(n9115), .ZN(n9116) );
  NOR2_X1 U10541 ( .A1(n9117), .A2(n9116), .ZN(n9122) );
  NOR4_X1 U10542 ( .A1(P2_REG2_REG_21__SCAN_IN), .A2(P1_REG1_REG_21__SCAN_IN), 
        .A3(P2_REG0_REG_11__SCAN_IN), .A4(n9118), .ZN(n9121) );
  INV_X1 U10543 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n9253) );
  AND4_X1 U10544 ( .A1(P1_IR_REG_24__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), 
        .A3(n9119), .A4(n9253), .ZN(n9120) );
  NAND4_X1 U10545 ( .A1(n9123), .A2(n9122), .A3(n9121), .A4(n9120), .ZN(n9124)
         );
  NOR2_X1 U10546 ( .A1(n9125), .A2(n9124), .ZN(n9126) );
  NAND4_X1 U10547 ( .A1(n9127), .A2(SI_14_), .A3(n9126), .A4(n9276), .ZN(n9135) );
  NAND4_X1 U10548 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), 
        .A3(P2_D_REG_25__SCAN_IN), .A4(n9128), .ZN(n9134) );
  NAND4_X1 U10549 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(P1_REG0_REG_3__SCAN_IN), 
        .A3(P2_REG0_REG_31__SCAN_IN), .A4(n10073), .ZN(n9132) );
  NAND4_X1 U10550 ( .A1(P1_D_REG_28__SCAN_IN), .A2(P1_ADDR_REG_19__SCAN_IN), 
        .A3(P2_REG2_REG_7__SCAN_IN), .A4(P2_REG0_REG_7__SCAN_IN), .ZN(n9131)
         );
  NAND4_X1 U10551 ( .A1(n9129), .A2(P1_REG0_REG_25__SCAN_IN), .A3(
        P1_REG0_REG_2__SCAN_IN), .A4(P1_ADDR_REG_17__SCAN_IN), .ZN(n9130) );
  OR3_X1 U10552 ( .A1(n9132), .A2(n9131), .A3(n9130), .ZN(n9133) );
  NOR4_X1 U10553 ( .A1(n9136), .A2(n9135), .A3(n9134), .A4(n9133), .ZN(n9141)
         );
  NAND2_X1 U10554 ( .A1(SI_12_), .A2(P2_D_REG_28__SCAN_IN), .ZN(n9139) );
  NAND4_X1 U10555 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P2_REG0_REG_2__SCAN_IN), 
        .A3(P1_REG0_REG_30__SCAN_IN), .A4(n9137), .ZN(n9138) );
  NOR4_X1 U10556 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .A3(
        n9139), .A4(n9138), .ZN(n9140) );
  AOI21_X1 U10557 ( .B1(n9141), .B2(n9140), .A(keyinput23), .ZN(n9142) );
  MUX2_X1 U10558 ( .A(keyinput23), .B(n9142), .S(n4495), .Z(n9143) );
  NAND3_X1 U10559 ( .A1(n9145), .A2(n9144), .A3(n9143), .ZN(n9146) );
  XNOR2_X1 U10560 ( .A(n9147), .B(n9146), .ZN(P2_U3467) );
  MUX2_X1 U10561 ( .A(n9149), .B(P2_REG1_REG_0__SCAN_IN), .S(n4269), .Z(
        P2_U3459) );
  NAND2_X1 U10562 ( .A1(n9150), .A2(n10185), .ZN(n9154) );
  NAND2_X1 U10563 ( .A1(n10188), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n9151) );
  OAI211_X1 U10564 ( .C1(n9152), .C2(n9264), .A(n9154), .B(n9151), .ZN(
        P2_U3458) );
  NAND2_X1 U10565 ( .A1(n9153), .A2(n9247), .ZN(n9155) );
  OAI211_X1 U10566 ( .C1(n10185), .C2(n9156), .A(n9155), .B(n9154), .ZN(
        P2_U3457) );
  MUX2_X1 U10567 ( .A(n9158), .B(n9157), .S(n10185), .Z(n9161) );
  NAND2_X1 U10568 ( .A1(n9159), .A2(n9247), .ZN(n9160) );
  OAI211_X1 U10569 ( .C1(n9162), .C2(n9255), .A(n9161), .B(n9160), .ZN(
        P2_U3455) );
  MUX2_X1 U10570 ( .A(n9164), .B(n9163), .S(n10185), .Z(n9167) );
  NAND2_X1 U10571 ( .A1(n9165), .A2(n9247), .ZN(n9166) );
  OAI211_X1 U10572 ( .C1(n9168), .C2(n9255), .A(n9167), .B(n9166), .ZN(
        P2_U3454) );
  MUX2_X1 U10573 ( .A(n9170), .B(n9169), .S(n10185), .Z(n9173) );
  NAND2_X1 U10574 ( .A1(n9171), .A2(n9247), .ZN(n9172) );
  OAI211_X1 U10575 ( .C1(n9174), .C2(n9255), .A(n9173), .B(n9172), .ZN(
        P2_U3453) );
  INV_X1 U10576 ( .A(n9175), .ZN(n9176) );
  MUX2_X1 U10577 ( .A(n9177), .B(n9176), .S(n10185), .Z(n9180) );
  NAND2_X1 U10578 ( .A1(n9178), .A2(n9247), .ZN(n9179) );
  OAI211_X1 U10579 ( .C1(n9181), .C2(n9255), .A(n9180), .B(n9179), .ZN(
        P2_U3452) );
  INV_X1 U10580 ( .A(n9182), .ZN(n9183) );
  MUX2_X1 U10581 ( .A(n9184), .B(n9183), .S(n10185), .Z(n9187) );
  NAND2_X1 U10582 ( .A1(n9185), .A2(n9247), .ZN(n9186) );
  OAI211_X1 U10583 ( .C1(n9188), .C2(n9255), .A(n9187), .B(n9186), .ZN(
        P2_U3451) );
  MUX2_X1 U10584 ( .A(n9190), .B(n9189), .S(n10185), .Z(n9193) );
  NAND2_X1 U10585 ( .A1(n9191), .A2(n9247), .ZN(n9192) );
  OAI211_X1 U10586 ( .C1(n9194), .C2(n9255), .A(n9193), .B(n9192), .ZN(
        P2_U3450) );
  INV_X1 U10587 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n9196) );
  MUX2_X1 U10588 ( .A(n9196), .B(n9195), .S(n10185), .Z(n9199) );
  NAND2_X1 U10589 ( .A1(n9197), .A2(n9247), .ZN(n9198) );
  OAI211_X1 U10590 ( .C1(n9200), .C2(n9255), .A(n9199), .B(n9198), .ZN(
        P2_U3449) );
  INV_X1 U10591 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n9202) );
  MUX2_X1 U10592 ( .A(n9202), .B(n9201), .S(n10185), .Z(n9203) );
  OAI21_X1 U10593 ( .B1(n9204), .B2(n9255), .A(n9203), .ZN(P2_U3448) );
  MUX2_X1 U10594 ( .A(n9206), .B(n9205), .S(n10185), .Z(n9209) );
  NAND2_X1 U10595 ( .A1(n9207), .A2(n9247), .ZN(n9208) );
  OAI211_X1 U10596 ( .C1(n9210), .C2(n9255), .A(n9209), .B(n9208), .ZN(
        P2_U3447) );
  INV_X1 U10597 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n9212) );
  MUX2_X1 U10598 ( .A(n9212), .B(n9211), .S(n10185), .Z(n9215) );
  NAND2_X1 U10599 ( .A1(n9213), .A2(n9247), .ZN(n9214) );
  OAI211_X1 U10600 ( .C1(n9216), .C2(n9255), .A(n9215), .B(n9214), .ZN(
        P2_U3446) );
  INV_X1 U10601 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n9218) );
  MUX2_X1 U10602 ( .A(n9218), .B(n9217), .S(n10185), .Z(n9219) );
  OAI21_X1 U10603 ( .B1(n9220), .B2(n9264), .A(n9219), .ZN(P2_U3444) );
  INV_X1 U10604 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n9222) );
  MUX2_X1 U10605 ( .A(n9222), .B(n9221), .S(n10185), .Z(n9225) );
  NAND2_X1 U10606 ( .A1(n9223), .A2(n9247), .ZN(n9224) );
  OAI211_X1 U10607 ( .C1(n9226), .C2(n9255), .A(n9225), .B(n9224), .ZN(
        P2_U3441) );
  INV_X1 U10608 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n9228) );
  MUX2_X1 U10609 ( .A(n9228), .B(n9227), .S(n10185), .Z(n9231) );
  NAND2_X1 U10610 ( .A1(n9229), .A2(n9247), .ZN(n9230) );
  OAI211_X1 U10611 ( .C1(n9232), .C2(n9255), .A(n9231), .B(n9230), .ZN(
        P2_U3438) );
  INV_X1 U10612 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n9234) );
  MUX2_X1 U10613 ( .A(n9234), .B(n9233), .S(n10185), .Z(n9237) );
  NAND2_X1 U10614 ( .A1(n9235), .A2(n9247), .ZN(n9236) );
  OAI211_X1 U10615 ( .C1(n9238), .C2(n9255), .A(n9237), .B(n9236), .ZN(
        P2_U3435) );
  INV_X1 U10616 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n9240) );
  MUX2_X1 U10617 ( .A(n9240), .B(n9239), .S(n10185), .Z(n9243) );
  NAND2_X1 U10618 ( .A1(n9241), .A2(n9247), .ZN(n9242) );
  OAI211_X1 U10619 ( .C1(n9244), .C2(n9255), .A(n9243), .B(n9242), .ZN(
        P2_U3432) );
  MUX2_X1 U10620 ( .A(n9246), .B(n9245), .S(n10185), .Z(n9250) );
  NAND2_X1 U10621 ( .A1(n9248), .A2(n9247), .ZN(n9249) );
  OAI211_X1 U10622 ( .C1(n9251), .C2(n9255), .A(n9250), .B(n9249), .ZN(
        P2_U3429) );
  MUX2_X1 U10623 ( .A(n9253), .B(n9252), .S(n10185), .Z(n9254) );
  OAI21_X1 U10624 ( .B1(n9256), .B2(n9255), .A(n9254), .ZN(P2_U3426) );
  INV_X1 U10625 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n9258) );
  MUX2_X1 U10626 ( .A(n9258), .B(n9257), .S(n10185), .Z(n9259) );
  OAI21_X1 U10627 ( .B1(n9260), .B2(n9264), .A(n9259), .ZN(P2_U3420) );
  INV_X1 U10628 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n9262) );
  MUX2_X1 U10629 ( .A(n9262), .B(n9261), .S(n10185), .Z(n9263) );
  OAI21_X1 U10630 ( .B1(n9265), .B2(n9264), .A(n9263), .ZN(P2_U3417) );
  MUX2_X1 U10631 ( .A(P2_REG0_REG_8__SCAN_IN), .B(n9266), .S(n10185), .Z(
        P2_U3414) );
  INV_X1 U10632 ( .A(n9267), .ZN(n9884) );
  NOR4_X1 U10633 ( .A1(n9269), .A2(P2_IR_REG_30__SCAN_IN), .A3(P2_U3151), .A4(
        n5023), .ZN(n9270) );
  AOI21_X1 U10634 ( .B1(n9279), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n9270), .ZN(
        n9271) );
  OAI21_X1 U10635 ( .B1(n9884), .B2(n9281), .A(n9271), .ZN(P2_U3264) );
  INV_X1 U10636 ( .A(n9272), .ZN(n9887) );
  OAI222_X1 U10637 ( .A1(n9283), .A2(n9274), .B1(n9281), .B2(n9887), .C1(
        P2_U3151), .C2(n9273), .ZN(P2_U3265) );
  INV_X1 U10638 ( .A(n9275), .ZN(n9890) );
  OAI222_X1 U10639 ( .A1(n9286), .A2(n9890), .B1(n9277), .B2(P2_U3151), .C1(
        n9276), .C2(n9283), .ZN(P2_U3266) );
  INV_X1 U10640 ( .A(n9278), .ZN(n9893) );
  AOI21_X1 U10641 ( .B1(P1_DATAO_REG_28__SCAN_IN), .B2(n9279), .A(n4364), .ZN(
        n9280) );
  OAI21_X1 U10642 ( .B1(n9893), .B2(n9281), .A(n9280), .ZN(P2_U3267) );
  INV_X1 U10643 ( .A(n9282), .ZN(n9898) );
  OAI222_X1 U10644 ( .A1(n9286), .A2(n9898), .B1(P2_U3151), .B2(n4270), .C1(
        n9284), .C2(n9283), .ZN(P2_U3268) );
  INV_X1 U10645 ( .A(n9287), .ZN(n9288) );
  MUX2_X1 U10646 ( .A(n9288), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  XOR2_X1 U10647 ( .A(n9366), .B(n9368), .Z(n9290) );
  NOR2_X1 U10648 ( .A1(n9290), .A2(n9289), .ZN(n9367) );
  AOI21_X1 U10649 ( .B1(n9290), .B2(n9289), .A(n9367), .ZN(n9297) );
  NAND2_X1 U10650 ( .A1(P1_U3086), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n9909) );
  OAI21_X1 U10651 ( .B1(n9477), .B2(n9291), .A(n9909), .ZN(n9292) );
  AOI21_X1 U10652 ( .B1(n9482), .B2(n9493), .A(n9292), .ZN(n9293) );
  OAI21_X1 U10653 ( .B1(n9479), .B2(n9294), .A(n9293), .ZN(n9295) );
  AOI21_X1 U10654 ( .B1(n9857), .B2(n9444), .A(n9295), .ZN(n9296) );
  OAI21_X1 U10655 ( .B1(n9297), .B2(n9458), .A(n9296), .ZN(P1_U3215) );
  AND3_X1 U10656 ( .A1(n9300), .A2(n9299), .A3(n9298), .ZN(n9301) );
  OAI21_X1 U10657 ( .B1(n9302), .B2(n9301), .A(n9474), .ZN(n9306) );
  AOI22_X1 U10658 ( .A1(n9641), .A2(n9451), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        P1_U3086), .ZN(n9303) );
  OAI21_X1 U10659 ( .B1(n9709), .B2(n9454), .A(n9303), .ZN(n9304) );
  AOI21_X1 U10660 ( .B1(n9676), .B2(n9468), .A(n9304), .ZN(n9305) );
  OAI211_X1 U10661 ( .C1(n9679), .C2(n9485), .A(n9306), .B(n9305), .ZN(
        P1_U3216) );
  XNOR2_X1 U10662 ( .A(n9308), .B(n9434), .ZN(n9310) );
  NOR2_X1 U10663 ( .A1(n9310), .A2(n9309), .ZN(n9433) );
  AOI21_X1 U10664 ( .B1(n9310), .B2(n9309), .A(n9433), .ZN(n9317) );
  AOI22_X1 U10665 ( .A1(n9444), .A2(n9311), .B1(n9482), .B2(n9497), .ZN(n9316)
         );
  NOR2_X1 U10666 ( .A1(n9479), .A2(n9312), .ZN(n9313) );
  AOI211_X1 U10667 ( .C1(n9451), .C2(n9495), .A(n9314), .B(n9313), .ZN(n9315)
         );
  OAI211_X1 U10668 ( .C1(n9317), .C2(n9458), .A(n9316), .B(n9315), .ZN(
        P1_U3217) );
  INV_X1 U10669 ( .A(n9318), .ZN(n9320) );
  NAND2_X1 U10670 ( .A1(n9320), .A2(n9319), .ZN(n9321) );
  OAI21_X1 U10671 ( .B1(n9320), .B2(n9319), .A(n9321), .ZN(n9449) );
  NOR2_X1 U10672 ( .A1(n9449), .A2(n9450), .ZN(n9448) );
  INV_X1 U10673 ( .A(n9321), .ZN(n9322) );
  NOR2_X1 U10674 ( .A1(n9448), .A2(n9322), .ZN(n9327) );
  INV_X1 U10675 ( .A(n9323), .ZN(n9325) );
  NOR2_X1 U10676 ( .A1(n9325), .A2(n9324), .ZN(n9326) );
  XNOR2_X1 U10677 ( .A(n9327), .B(n9326), .ZN(n9333) );
  OAI21_X1 U10678 ( .B1(n9477), .B2(n9740), .A(n9328), .ZN(n9329) );
  AOI21_X1 U10679 ( .B1(n9482), .B2(n9772), .A(n9329), .ZN(n9330) );
  OAI21_X1 U10680 ( .B1(n9479), .B2(n9732), .A(n9330), .ZN(n9331) );
  AOI21_X1 U10681 ( .B1(n9834), .B2(n9444), .A(n9331), .ZN(n9332) );
  OAI21_X1 U10682 ( .B1(n9333), .B2(n9458), .A(n9332), .ZN(P1_U3219) );
  OAI22_X1 U10683 ( .A1(n9599), .A2(n9334), .B1(n9607), .B2(n6389), .ZN(n9336)
         );
  XNOR2_X1 U10684 ( .A(n9336), .B(n9335), .ZN(n9339) );
  OAI22_X1 U10685 ( .A1(n9599), .A2(n6389), .B1(n9607), .B2(n4423), .ZN(n9338)
         );
  XNOR2_X1 U10686 ( .A(n9339), .B(n9338), .ZN(n9340) );
  INV_X1 U10687 ( .A(n9340), .ZN(n9346) );
  NAND3_X1 U10688 ( .A1(n9346), .A2(n9474), .A3(n9345), .ZN(n9351) );
  NAND3_X1 U10689 ( .A1(n9352), .A2(n9474), .A3(n9340), .ZN(n9350) );
  INV_X1 U10690 ( .A(n9596), .ZN(n9344) );
  INV_X1 U10691 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n9341) );
  OAI22_X1 U10692 ( .A1(n9591), .A2(n9477), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9341), .ZN(n9342) );
  AOI21_X1 U10693 ( .B1(n9482), .B2(n9590), .A(n9342), .ZN(n9343) );
  OAI21_X1 U10694 ( .B1(n9479), .B2(n9344), .A(n9343), .ZN(n9348) );
  NOR3_X1 U10695 ( .A1(n9346), .A2(n9345), .A3(n9458), .ZN(n9347) );
  AOI211_X1 U10696 ( .C1(n9788), .C2(n9444), .A(n9348), .B(n9347), .ZN(n9349)
         );
  OAI211_X1 U10697 ( .C1(n9352), .C2(n9351), .A(n9350), .B(n9349), .ZN(
        P1_U3220) );
  XOR2_X1 U10698 ( .A(n9353), .B(n9354), .Z(n9359) );
  AOI22_X1 U10699 ( .A1(n9489), .A2(n9451), .B1(P1_REG3_REG_21__SCAN_IN), .B2(
        P1_U3086), .ZN(n9356) );
  NAND2_X1 U10700 ( .A1(n9482), .A2(n9490), .ZN(n9355) );
  OAI211_X1 U10701 ( .C1(n9479), .C2(n9701), .A(n9356), .B(n9355), .ZN(n9357)
         );
  AOI21_X1 U10702 ( .B1(n9824), .B2(n9444), .A(n9357), .ZN(n9358) );
  OAI21_X1 U10703 ( .B1(n9359), .B2(n9458), .A(n9358), .ZN(P1_U3223) );
  AOI21_X1 U10704 ( .B1(n4315), .B2(n9360), .A(n9463), .ZN(n9365) );
  AOI22_X1 U10705 ( .A1(n9642), .A2(n9451), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3086), .ZN(n9362) );
  NAND2_X1 U10706 ( .A1(n9641), .A2(n9482), .ZN(n9361) );
  OAI211_X1 U10707 ( .C1(n9479), .C2(n9646), .A(n9362), .B(n9361), .ZN(n9363)
         );
  AOI21_X1 U10708 ( .B1(n9804), .B2(n9444), .A(n9363), .ZN(n9364) );
  OAI21_X1 U10709 ( .B1(n9365), .B2(n9458), .A(n9364), .ZN(P1_U3225) );
  INV_X1 U10710 ( .A(n9366), .ZN(n9369) );
  AOI21_X1 U10711 ( .B1(n9369), .B2(n9368), .A(n9367), .ZN(n9372) );
  XNOR2_X1 U10712 ( .A(n9372), .B(n9370), .ZN(n9472) );
  NAND2_X1 U10713 ( .A1(n9472), .A2(n9473), .ZN(n9471) );
  OAI21_X1 U10714 ( .B1(n9372), .B2(n9371), .A(n9471), .ZN(n9376) );
  XNOR2_X1 U10715 ( .A(n9374), .B(n9373), .ZN(n9375) );
  XNOR2_X1 U10716 ( .A(n9376), .B(n9375), .ZN(n9382) );
  NAND2_X1 U10717 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9935) );
  OAI21_X1 U10718 ( .B1(n9477), .B2(n9453), .A(n9935), .ZN(n9377) );
  AOI21_X1 U10719 ( .B1(n9482), .B2(n9491), .A(n9377), .ZN(n9378) );
  OAI21_X1 U10720 ( .B1(n9479), .B2(n9379), .A(n9378), .ZN(n9380) );
  AOI21_X1 U10721 ( .B1(n9848), .B2(n9444), .A(n9380), .ZN(n9381) );
  OAI21_X1 U10722 ( .B1(n9382), .B2(n9458), .A(n9381), .ZN(P1_U3226) );
  XNOR2_X1 U10723 ( .A(n9384), .B(n9383), .ZN(n9385) );
  XNOR2_X1 U10724 ( .A(n9386), .B(n9385), .ZN(n9391) );
  NAND2_X1 U10725 ( .A1(n9482), .A2(n9771), .ZN(n9387) );
  NAND2_X1 U10726 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9950) );
  OAI211_X1 U10727 ( .C1(n9477), .C2(n9739), .A(n9387), .B(n9950), .ZN(n9389)
         );
  NOR2_X1 U10728 ( .A1(n9767), .A2(n9485), .ZN(n9388) );
  AOI211_X1 U10729 ( .C1(n9775), .C2(n9468), .A(n9389), .B(n9388), .ZN(n9390)
         );
  OAI21_X1 U10730 ( .B1(n9391), .B2(n9458), .A(n9390), .ZN(P1_U3228) );
  AOI21_X1 U10731 ( .B1(n9392), .B2(n9393), .A(n9458), .ZN(n9395) );
  NAND2_X1 U10732 ( .A1(n9395), .A2(n9394), .ZN(n9399) );
  AOI22_X1 U10733 ( .A1(n9444), .A2(n10018), .B1(n9451), .B2(n7358), .ZN(n9398) );
  AND2_X1 U10734 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_U3086), .ZN(n9545) );
  AOI21_X1 U10735 ( .B1(n9482), .B2(n10011), .A(n9545), .ZN(n9397) );
  OR2_X1 U10736 ( .A1(n9479), .A2(n10014), .ZN(n9396) );
  NAND4_X1 U10737 ( .A1(n9399), .A2(n9398), .A3(n9397), .A4(n9396), .ZN(
        P1_U3230) );
  AOI21_X1 U10738 ( .B1(n9402), .B2(n9401), .A(n9400), .ZN(n9406) );
  XNOR2_X1 U10739 ( .A(n9404), .B(n9403), .ZN(n9405) );
  XNOR2_X1 U10740 ( .A(n9406), .B(n9405), .ZN(n9412) );
  AOI22_X1 U10741 ( .A1(n9444), .A2(n9407), .B1(n9482), .B2(n9498), .ZN(n9411)
         );
  AND2_X1 U10742 ( .A1(P1_U3086), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n9571) );
  NOR2_X1 U10743 ( .A1(n9479), .A2(n9408), .ZN(n9409) );
  AOI211_X1 U10744 ( .C1(n9451), .C2(n9496), .A(n9571), .B(n9409), .ZN(n9410)
         );
  OAI211_X1 U10745 ( .C1(n9412), .C2(n9458), .A(n9411), .B(n9410), .ZN(
        P1_U3231) );
  XNOR2_X1 U10746 ( .A(n9414), .B(n9413), .ZN(n9415) );
  XNOR2_X1 U10747 ( .A(n9416), .B(n9415), .ZN(n9421) );
  NAND2_X1 U10748 ( .A1(n9468), .A2(n9721), .ZN(n9418) );
  AOI22_X1 U10749 ( .A1(n9451), .A2(n9686), .B1(P1_REG3_REG_20__SCAN_IN), .B2(
        P1_U3086), .ZN(n9417) );
  OAI211_X1 U10750 ( .C1(n9717), .C2(n9454), .A(n9418), .B(n9417), .ZN(n9419)
         );
  AOI21_X1 U10751 ( .B1(n9829), .B2(n9444), .A(n9419), .ZN(n9420) );
  OAI21_X1 U10752 ( .B1(n9421), .B2(n9458), .A(n9420), .ZN(P1_U3233) );
  XOR2_X1 U10753 ( .A(n9422), .B(n9423), .Z(n9432) );
  OAI21_X1 U10754 ( .B1(n9477), .B2(n9425), .A(n9424), .ZN(n9426) );
  AOI21_X1 U10755 ( .B1(n9482), .B2(n9494), .A(n9426), .ZN(n9427) );
  OAI21_X1 U10756 ( .B1(n9479), .B2(n9428), .A(n9427), .ZN(n9429) );
  AOI21_X1 U10757 ( .B1(n9430), .B2(n9444), .A(n9429), .ZN(n9431) );
  OAI21_X1 U10758 ( .B1(n9432), .B2(n9458), .A(n9431), .ZN(P1_U3234) );
  AOI21_X1 U10759 ( .B1(n9434), .B2(n9308), .A(n9433), .ZN(n9438) );
  XNOR2_X1 U10760 ( .A(n9436), .B(n9435), .ZN(n9437) );
  XNOR2_X1 U10761 ( .A(n9438), .B(n9437), .ZN(n9447) );
  AOI21_X1 U10762 ( .B1(n9482), .B2(n9496), .A(n9439), .ZN(n9441) );
  NAND2_X1 U10763 ( .A1(n9451), .A2(n9494), .ZN(n9440) );
  OAI211_X1 U10764 ( .C1(n9479), .C2(n9442), .A(n9441), .B(n9440), .ZN(n9443)
         );
  AOI21_X1 U10765 ( .B1(n9445), .B2(n9444), .A(n9443), .ZN(n9446) );
  OAI21_X1 U10766 ( .B1(n9447), .B2(n9458), .A(n9446), .ZN(P1_U3236) );
  AOI21_X1 U10767 ( .B1(n9450), .B2(n9449), .A(n9448), .ZN(n9459) );
  NAND2_X1 U10768 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9968) );
  NAND2_X1 U10769 ( .A1(n9451), .A2(n9754), .ZN(n9452) );
  OAI211_X1 U10770 ( .C1(n9454), .C2(n9453), .A(n9968), .B(n9452), .ZN(n9456)
         );
  NOR2_X1 U10771 ( .A1(n9747), .A2(n9485), .ZN(n9455) );
  AOI211_X1 U10772 ( .C1(n9745), .C2(n9468), .A(n9456), .B(n9455), .ZN(n9457)
         );
  OAI21_X1 U10773 ( .B1(n9459), .B2(n9458), .A(n9457), .ZN(P1_U3238) );
  OAI21_X1 U10774 ( .B1(n9463), .B2(n9462), .A(n9461), .ZN(n9464) );
  NAND3_X1 U10775 ( .A1(n9465), .A2(n9474), .A3(n9464), .ZN(n9470) );
  AOI22_X1 U10776 ( .A1(n9657), .A2(n9482), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3086), .ZN(n9466) );
  OAI21_X1 U10777 ( .B1(n9631), .B2(n9477), .A(n9466), .ZN(n9467) );
  AOI21_X1 U10778 ( .B1(n9632), .B2(n9468), .A(n9467), .ZN(n9469) );
  OAI211_X1 U10779 ( .C1(n9626), .C2(n9485), .A(n9470), .B(n9469), .ZN(
        P1_U3240) );
  OAI21_X1 U10780 ( .B1(n9473), .B2(n9472), .A(n9471), .ZN(n9475) );
  NAND2_X1 U10781 ( .A1(n9475), .A2(n9474), .ZN(n9484) );
  NAND2_X1 U10782 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9922) );
  OAI21_X1 U10783 ( .B1(n9477), .B2(n9476), .A(n9922), .ZN(n9481) );
  NOR2_X1 U10784 ( .A1(n9479), .A2(n9478), .ZN(n9480) );
  AOI211_X1 U10785 ( .C1(n9482), .C2(n9492), .A(n9481), .B(n9480), .ZN(n9483)
         );
  OAI211_X1 U10786 ( .C1(n9486), .C2(n9485), .A(n9484), .B(n9483), .ZN(
        P1_U3241) );
  MUX2_X1 U10787 ( .A(n9487), .B(P1_DATAO_REG_30__SCAN_IN), .S(n9501), .Z(
        P1_U3584) );
  MUX2_X1 U10788 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9488), .S(P1_U3973), .Z(
        P1_U3582) );
  MUX2_X1 U10789 ( .A(n9590), .B(P1_DATAO_REG_27__SCAN_IN), .S(n9501), .Z(
        P1_U3581) );
  MUX2_X1 U10790 ( .A(n9642), .B(P1_DATAO_REG_26__SCAN_IN), .S(n9501), .Z(
        P1_U3580) );
  MUX2_X1 U10791 ( .A(n9657), .B(P1_DATAO_REG_25__SCAN_IN), .S(n9501), .Z(
        P1_U3579) );
  MUX2_X1 U10792 ( .A(n9641), .B(P1_DATAO_REG_24__SCAN_IN), .S(n9501), .Z(
        P1_U3578) );
  MUX2_X1 U10793 ( .A(n9687), .B(P1_DATAO_REG_23__SCAN_IN), .S(n9501), .Z(
        P1_U3577) );
  MUX2_X1 U10794 ( .A(n9489), .B(P1_DATAO_REG_22__SCAN_IN), .S(n9501), .Z(
        P1_U3576) );
  MUX2_X1 U10795 ( .A(n9686), .B(P1_DATAO_REG_21__SCAN_IN), .S(n9501), .Z(
        P1_U3575) );
  MUX2_X1 U10796 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9490), .S(P1_U3973), .Z(
        P1_U3574) );
  MUX2_X1 U10797 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9754), .S(P1_U3973), .Z(
        P1_U3573) );
  MUX2_X1 U10798 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9772), .S(P1_U3973), .Z(
        P1_U3572) );
  MUX2_X1 U10799 ( .A(n9755), .B(P1_DATAO_REG_17__SCAN_IN), .S(n9501), .Z(
        P1_U3571) );
  MUX2_X1 U10800 ( .A(n9771), .B(P1_DATAO_REG_16__SCAN_IN), .S(n9501), .Z(
        P1_U3570) );
  MUX2_X1 U10801 ( .A(n9491), .B(P1_DATAO_REG_15__SCAN_IN), .S(n9501), .Z(
        P1_U3569) );
  MUX2_X1 U10802 ( .A(n9492), .B(P1_DATAO_REG_14__SCAN_IN), .S(n9501), .Z(
        P1_U3568) );
  MUX2_X1 U10803 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9493), .S(P1_U3973), .Z(
        P1_U3567) );
  MUX2_X1 U10804 ( .A(n9494), .B(P1_DATAO_REG_12__SCAN_IN), .S(n9501), .Z(
        P1_U3566) );
  MUX2_X1 U10805 ( .A(n9495), .B(P1_DATAO_REG_11__SCAN_IN), .S(n9501), .Z(
        P1_U3565) );
  MUX2_X1 U10806 ( .A(n9496), .B(P1_DATAO_REG_10__SCAN_IN), .S(n9501), .Z(
        P1_U3564) );
  MUX2_X1 U10807 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n9497), .S(P1_U3973), .Z(
        P1_U3563) );
  MUX2_X1 U10808 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9498), .S(P1_U3973), .Z(
        P1_U3562) );
  MUX2_X1 U10809 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n9992), .S(P1_U3973), .Z(
        P1_U3561) );
  MUX2_X1 U10810 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n9499), .S(P1_U3973), .Z(
        P1_U3560) );
  MUX2_X1 U10811 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n7358), .S(P1_U3973), .Z(
        P1_U3559) );
  MUX2_X1 U10812 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n9500), .S(P1_U3973), .Z(
        P1_U3558) );
  MUX2_X1 U10813 ( .A(n10011), .B(P1_DATAO_REG_3__SCAN_IN), .S(n9501), .Z(
        P1_U3557) );
  MUX2_X1 U10814 ( .A(n7352), .B(P1_DATAO_REG_2__SCAN_IN), .S(n9501), .Z(
        P1_U3556) );
  MUX2_X1 U10815 ( .A(n7346), .B(P1_DATAO_REG_0__SCAN_IN), .S(n9501), .Z(
        P1_U3554) );
  INV_X1 U10816 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n9503) );
  OAI22_X1 U10817 ( .A1(n9970), .A2(n9503), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9502), .ZN(n9504) );
  AOI21_X1 U10818 ( .B1(n9505), .B2(n9959), .A(n9504), .ZN(n9513) );
  OAI211_X1 U10819 ( .C1(n9514), .C2(n9507), .A(n9957), .B(n9506), .ZN(n9512)
         );
  OAI211_X1 U10820 ( .C1(n9510), .C2(n9509), .A(n9964), .B(n9508), .ZN(n9511)
         );
  NAND3_X1 U10821 ( .A1(n9513), .A2(n9512), .A3(n9511), .ZN(P1_U3244) );
  MUX2_X1 U10822 ( .A(n9515), .B(n9514), .S(n9895), .Z(n9518) );
  OAI21_X1 U10823 ( .B1(P1_IR_REG_0__SCAN_IN), .B2(n9516), .A(P1_U3973), .ZN(
        n9517) );
  AOI21_X1 U10824 ( .B1(n9518), .B2(n9891), .A(n9517), .ZN(n9519) );
  INV_X1 U10825 ( .A(n9519), .ZN(n9560) );
  INV_X1 U10826 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n9520) );
  OAI22_X1 U10827 ( .A1(n9970), .A2(n9520), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10043), .ZN(n9521) );
  AOI21_X1 U10828 ( .B1(n4431), .B2(n9959), .A(n9521), .ZN(n9531) );
  OAI211_X1 U10829 ( .C1(n9525), .C2(n9524), .A(n9964), .B(n9523), .ZN(n9530)
         );
  OAI211_X1 U10830 ( .C1(n9528), .C2(n9527), .A(n9957), .B(n9526), .ZN(n9529)
         );
  NAND4_X1 U10831 ( .A1(n9560), .A2(n9531), .A3(n9530), .A4(n9529), .ZN(
        P1_U3245) );
  INV_X1 U10832 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n9533) );
  OAI21_X1 U10833 ( .B1(n9970), .B2(n9533), .A(n9532), .ZN(n9534) );
  AOI21_X1 U10834 ( .B1(n9535), .B2(n9959), .A(n9534), .ZN(n9544) );
  OAI211_X1 U10835 ( .C1(n9538), .C2(n9537), .A(n9964), .B(n9536), .ZN(n9543)
         );
  OAI211_X1 U10836 ( .C1(n9541), .C2(n9540), .A(n9957), .B(n9539), .ZN(n9542)
         );
  NAND3_X1 U10837 ( .A1(n9544), .A2(n9543), .A3(n9542), .ZN(P1_U3246) );
  AOI21_X1 U10838 ( .B1(n9546), .B2(P1_ADDR_REG_4__SCAN_IN), .A(n9545), .ZN(
        n9559) );
  NOR2_X1 U10839 ( .A1(n9548), .A2(n9547), .ZN(n9549) );
  NOR2_X1 U10840 ( .A1(n9550), .A2(n9549), .ZN(n9551) );
  AOI22_X1 U10841 ( .A1(n4422), .A2(n9959), .B1(n9957), .B2(n9551), .ZN(n9558)
         );
  INV_X1 U10842 ( .A(n9553), .ZN(n9554) );
  OAI211_X1 U10843 ( .C1(n9556), .C2(n9555), .A(n9964), .B(n9554), .ZN(n9557)
         );
  NAND4_X1 U10844 ( .A1(n9560), .A2(n9559), .A3(n9558), .A4(n9557), .ZN(
        P1_U3247) );
  OAI21_X1 U10845 ( .B1(n9563), .B2(n9562), .A(n9561), .ZN(n9564) );
  NAND2_X1 U10846 ( .A1(n9564), .A2(n9957), .ZN(n9575) );
  OAI21_X1 U10847 ( .B1(n9567), .B2(n9566), .A(n9565), .ZN(n9568) );
  NAND2_X1 U10848 ( .A1(n9568), .A2(n9964), .ZN(n9574) );
  INV_X1 U10849 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n9569) );
  NOR2_X1 U10850 ( .A1(n9970), .A2(n9569), .ZN(n9570) );
  AOI211_X1 U10851 ( .C1(n9572), .C2(n9959), .A(n9571), .B(n9570), .ZN(n9573)
         );
  NAND3_X1 U10852 ( .A1(n9575), .A2(n9574), .A3(n9573), .ZN(P1_U3252) );
  NOR2_X1 U10853 ( .A1(n10070), .A2(n9576), .ZN(n9577) );
  AOI211_X1 U10854 ( .C1(n9579), .C2(n10017), .A(n9578), .B(n9577), .ZN(n9580)
         );
  OAI21_X1 U10855 ( .B1(n9582), .B2(n9581), .A(n9580), .ZN(P1_U3263) );
  INV_X1 U10856 ( .A(n9585), .ZN(n9587) );
  NAND3_X1 U10857 ( .A1(n9589), .A2(n10013), .A3(n9588), .ZN(n9594) );
  NAND2_X1 U10858 ( .A1(n9590), .A2(n10010), .ZN(n9592) );
  AOI211_X1 U10859 ( .C1(n9788), .C2(n9612), .A(n10039), .B(n9595), .ZN(n9789)
         );
  NAND2_X1 U10860 ( .A1(n9789), .A2(n10031), .ZN(n9598) );
  AOI22_X1 U10861 ( .A1(n9596), .A2(n10015), .B1(P1_REG2_REG_28__SCAN_IN), 
        .B2(n4984), .ZN(n9597) );
  OAI211_X1 U10862 ( .C1(n9599), .C2(n9766), .A(n9598), .B(n9597), .ZN(n9600)
         );
  AOI21_X1 U10863 ( .B1(n9790), .B2(n10070), .A(n9600), .ZN(n9601) );
  OAI21_X1 U10864 ( .B1(n9793), .B2(n9780), .A(n9601), .ZN(P1_U3265) );
  NAND2_X1 U10865 ( .A1(n9642), .A2(n10010), .ZN(n9606) );
  OAI21_X1 U10866 ( .B1(n9607), .B2(n10048), .A(n9606), .ZN(n9608) );
  INV_X1 U10867 ( .A(n9608), .ZN(n9609) );
  INV_X1 U10868 ( .A(n9624), .ZN(n9614) );
  INV_X1 U10869 ( .A(n9612), .ZN(n9613) );
  AOI211_X1 U10870 ( .C1(n9796), .C2(n9614), .A(n10039), .B(n9613), .ZN(n9795)
         );
  NAND2_X1 U10871 ( .A1(n9795), .A2(n10031), .ZN(n9618) );
  INV_X1 U10872 ( .A(n9615), .ZN(n9616) );
  AOI22_X1 U10873 ( .A1(n9616), .A2(n10015), .B1(P1_REG2_REG_27__SCAN_IN), 
        .B2(n4984), .ZN(n9617) );
  OAI211_X1 U10874 ( .C1(n9619), .C2(n9766), .A(n9618), .B(n9617), .ZN(n9620)
         );
  AOI21_X1 U10875 ( .B1(n9794), .B2(n10070), .A(n9620), .ZN(n9621) );
  OAI21_X1 U10876 ( .B1(n9798), .B2(n9780), .A(n9621), .ZN(P1_U3266) );
  XOR2_X1 U10877 ( .A(n9622), .B(n9629), .Z(n9801) );
  NOR2_X1 U10878 ( .A1(n9626), .A2(n9645), .ZN(n9623) );
  OAI22_X1 U10879 ( .A1(n9626), .A2(n9766), .B1(n9625), .B2(n10070), .ZN(n9635) );
  NOR2_X1 U10880 ( .A1(n9633), .A2(n4984), .ZN(n9634) );
  AOI211_X1 U10881 ( .C1(n10031), .C2(n4973), .A(n9635), .B(n9634), .ZN(n9636)
         );
  OAI21_X1 U10882 ( .B1(n9780), .B2(n9801), .A(n9636), .ZN(P1_U3267) );
  XNOR2_X1 U10883 ( .A(n9637), .B(n9639), .ZN(n9806) );
  OAI211_X1 U10884 ( .C1(n9640), .C2(n9639), .A(n9638), .B(n10013), .ZN(n9644)
         );
  AOI22_X1 U10885 ( .A1(n9642), .A2(n10009), .B1(n10010), .B2(n9641), .ZN(
        n9643) );
  NAND2_X1 U10886 ( .A1(n9644), .A2(n9643), .ZN(n9802) );
  AOI211_X1 U10887 ( .C1(n9804), .C2(n9660), .A(n10039), .B(n9645), .ZN(n9803)
         );
  NAND2_X1 U10888 ( .A1(n9803), .A2(n10031), .ZN(n9649) );
  INV_X1 U10889 ( .A(n9646), .ZN(n9647) );
  AOI22_X1 U10890 ( .A1(n9647), .A2(n10015), .B1(P1_REG2_REG_25__SCAN_IN), 
        .B2(n4984), .ZN(n9648) );
  OAI211_X1 U10891 ( .C1(n9650), .C2(n9766), .A(n9649), .B(n9648), .ZN(n9651)
         );
  AOI21_X1 U10892 ( .B1(n9802), .B2(n10070), .A(n9651), .ZN(n9652) );
  OAI21_X1 U10893 ( .B1(n9806), .B2(n9780), .A(n9652), .ZN(P1_U3268) );
  XOR2_X1 U10894 ( .A(n9655), .B(n9653), .Z(n9811) );
  OAI211_X1 U10895 ( .C1(n9656), .C2(n9655), .A(n9654), .B(n10013), .ZN(n9659)
         );
  AOI22_X1 U10896 ( .A1(n9657), .A2(n10009), .B1(n10010), .B2(n9687), .ZN(
        n9658) );
  NAND2_X1 U10897 ( .A1(n9659), .A2(n9658), .ZN(n9807) );
  AOI211_X1 U10898 ( .C1(n9809), .C2(n9674), .A(n10039), .B(n6523), .ZN(n9808)
         );
  NAND2_X1 U10899 ( .A1(n9808), .A2(n10031), .ZN(n9663) );
  AOI22_X1 U10900 ( .A1(n9661), .A2(n10015), .B1(P1_REG2_REG_24__SCAN_IN), 
        .B2(n4984), .ZN(n9662) );
  OAI211_X1 U10901 ( .C1(n9664), .C2(n9766), .A(n9663), .B(n9662), .ZN(n9665)
         );
  AOI21_X1 U10902 ( .B1(n9807), .B2(n10070), .A(n9665), .ZN(n9666) );
  OAI21_X1 U10903 ( .B1(n9811), .B2(n9780), .A(n9666), .ZN(P1_U3269) );
  XNOR2_X1 U10904 ( .A(n9667), .B(n9668), .ZN(n9816) );
  AOI21_X1 U10905 ( .B1(n9671), .B2(n9670), .A(n9669), .ZN(n9672) );
  OAI222_X1 U10906 ( .A1(n10050), .A2(n9709), .B1(n10048), .B2(n9673), .C1(
        n10047), .C2(n9672), .ZN(n9812) );
  INV_X1 U10907 ( .A(n9674), .ZN(n9675) );
  AOI211_X1 U10908 ( .C1(n9814), .C2(n4898), .A(n10039), .B(n9675), .ZN(n9813)
         );
  NAND2_X1 U10909 ( .A1(n9813), .A2(n10031), .ZN(n9678) );
  AOI22_X1 U10910 ( .A1(n9676), .A2(n10015), .B1(P1_REG2_REG_23__SCAN_IN), 
        .B2(n4984), .ZN(n9677) );
  OAI211_X1 U10911 ( .C1(n9679), .C2(n9766), .A(n9678), .B(n9677), .ZN(n9680)
         );
  AOI21_X1 U10912 ( .B1(n9812), .B2(n10070), .A(n9680), .ZN(n9681) );
  OAI21_X1 U10913 ( .B1(n9816), .B2(n9780), .A(n9681), .ZN(P1_U3270) );
  XOR2_X1 U10914 ( .A(n9682), .B(n9684), .Z(n9821) );
  OAI211_X1 U10915 ( .C1(n9685), .C2(n9684), .A(n9683), .B(n10013), .ZN(n9689)
         );
  AOI22_X1 U10916 ( .A1(n9687), .A2(n10009), .B1(n10010), .B2(n9686), .ZN(
        n9688) );
  NAND2_X1 U10917 ( .A1(n9689), .A2(n9688), .ZN(n9817) );
  AOI211_X1 U10918 ( .C1(n9819), .C2(n9699), .A(n10039), .B(n9690), .ZN(n9818)
         );
  NAND2_X1 U10919 ( .A1(n9818), .A2(n10031), .ZN(n9694) );
  INV_X1 U10920 ( .A(n9691), .ZN(n9692) );
  AOI22_X1 U10921 ( .A1(n9692), .A2(n10015), .B1(n4984), .B2(
        P1_REG2_REG_22__SCAN_IN), .ZN(n9693) );
  OAI211_X1 U10922 ( .C1(n9695), .C2(n9766), .A(n9694), .B(n9693), .ZN(n9696)
         );
  AOI21_X1 U10923 ( .B1(n9817), .B2(n10070), .A(n9696), .ZN(n9697) );
  OAI21_X1 U10924 ( .B1(n9821), .B2(n9780), .A(n9697), .ZN(P1_U3271) );
  XOR2_X1 U10925 ( .A(n9698), .B(n9706), .Z(n9826) );
  INV_X1 U10926 ( .A(n9699), .ZN(n9700) );
  AOI211_X1 U10927 ( .C1(n9824), .C2(n9718), .A(n10039), .B(n9700), .ZN(n9823)
         );
  NOR2_X1 U10928 ( .A1(n8063), .A2(n9766), .ZN(n9704) );
  OAI22_X1 U10929 ( .A1(n10070), .A2(n9702), .B1(n9701), .B2(n10068), .ZN(
        n9703) );
  AOI211_X1 U10930 ( .C1(n9823), .C2(n10031), .A(n9704), .B(n9703), .ZN(n9711)
         );
  INV_X1 U10931 ( .A(n9712), .ZN(n9714) );
  OAI21_X1 U10932 ( .B1(n9715), .B2(n9714), .A(n9705), .ZN(n9707) );
  XNOR2_X1 U10933 ( .A(n9707), .B(n9706), .ZN(n9708) );
  OAI222_X1 U10934 ( .A1(n10048), .A2(n9709), .B1(n10050), .B2(n9740), .C1(
        n9708), .C2(n10047), .ZN(n9822) );
  NAND2_X1 U10935 ( .A1(n9822), .A2(n10070), .ZN(n9710) );
  OAI211_X1 U10936 ( .C1(n9826), .C2(n9780), .A(n9711), .B(n9710), .ZN(
        P1_U3272) );
  XNOR2_X1 U10937 ( .A(n9713), .B(n9712), .ZN(n9831) );
  XNOR2_X1 U10938 ( .A(n9715), .B(n9714), .ZN(n9716) );
  OAI222_X1 U10939 ( .A1(n10048), .A2(n8062), .B1(n10050), .B2(n9717), .C1(
        n10047), .C2(n9716), .ZN(n9827) );
  INV_X1 U10940 ( .A(n9729), .ZN(n9720) );
  INV_X1 U10941 ( .A(n9718), .ZN(n9719) );
  AOI211_X1 U10942 ( .C1(n9829), .C2(n9720), .A(n10039), .B(n9719), .ZN(n9828)
         );
  NAND2_X1 U10943 ( .A1(n9828), .A2(n10031), .ZN(n9723) );
  AOI22_X1 U10944 ( .A1(n4984), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9721), .B2(
        n10015), .ZN(n9722) );
  OAI211_X1 U10945 ( .C1(n9724), .C2(n9766), .A(n9723), .B(n9722), .ZN(n9725)
         );
  AOI21_X1 U10946 ( .B1(n9827), .B2(n10070), .A(n9725), .ZN(n9726) );
  OAI21_X1 U10947 ( .B1(n9831), .B2(n9780), .A(n9726), .ZN(P1_U3273) );
  XNOR2_X1 U10948 ( .A(n9728), .B(n9727), .ZN(n9836) );
  INV_X1 U10949 ( .A(n9744), .ZN(n9730) );
  AOI211_X1 U10950 ( .C1(n9834), .C2(n9730), .A(n10039), .B(n9729), .ZN(n9833)
         );
  NOR2_X1 U10951 ( .A1(n9731), .A2(n9766), .ZN(n9735) );
  OAI22_X1 U10952 ( .A1(n10070), .A2(n9733), .B1(n9732), .B2(n10068), .ZN(
        n9734) );
  AOI211_X1 U10953 ( .C1(n9833), .C2(n10031), .A(n9735), .B(n9734), .ZN(n9742)
         );
  XNOR2_X1 U10954 ( .A(n9737), .B(n9736), .ZN(n9738) );
  OAI222_X1 U10955 ( .A1(n10048), .A2(n9740), .B1(n10050), .B2(n9739), .C1(
        n9738), .C2(n10047), .ZN(n9832) );
  NAND2_X1 U10956 ( .A1(n9832), .A2(n10070), .ZN(n9741) );
  OAI211_X1 U10957 ( .C1(n9836), .C2(n9780), .A(n9742), .B(n9741), .ZN(
        P1_U3274) );
  XNOR2_X1 U10958 ( .A(n9743), .B(n9752), .ZN(n9840) );
  AOI211_X1 U10959 ( .C1(n7834), .C2(n4895), .A(n10039), .B(n9744), .ZN(n9837)
         );
  AOI22_X1 U10960 ( .A1(n4984), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9745), .B2(
        n10015), .ZN(n9746) );
  OAI21_X1 U10961 ( .B1(n9747), .B2(n9766), .A(n9746), .ZN(n9758) );
  INV_X1 U10962 ( .A(n9768), .ZN(n9750) );
  NOR2_X1 U10963 ( .A1(n9750), .A2(n9749), .ZN(n9753) );
  OAI21_X1 U10964 ( .B1(n9753), .B2(n9752), .A(n4404), .ZN(n9756) );
  AOI222_X1 U10965 ( .A1(n10013), .A2(n9756), .B1(n9755), .B2(n10010), .C1(
        n9754), .C2(n10009), .ZN(n9839) );
  NOR2_X1 U10966 ( .A1(n9839), .A2(n4984), .ZN(n9757) );
  AOI211_X1 U10967 ( .C1(n9837), .C2(n10031), .A(n9758), .B(n9757), .ZN(n9759)
         );
  OAI21_X1 U10968 ( .B1(n9840), .B2(n9780), .A(n9759), .ZN(P1_U3275) );
  XOR2_X1 U10969 ( .A(n9769), .B(n9760), .Z(n9845) );
  NAND2_X1 U10970 ( .A1(n9761), .A2(n9843), .ZN(n9762) );
  NAND2_X1 U10971 ( .A1(n9762), .A2(n10027), .ZN(n9763) );
  NOR2_X1 U10972 ( .A1(n9764), .A2(n9763), .ZN(n9842) );
  OAI22_X1 U10973 ( .A1(n9767), .A2(n9766), .B1(n9765), .B2(n10070), .ZN(n9778) );
  OAI211_X1 U10974 ( .C1(n9770), .C2(n9769), .A(n9768), .B(n10013), .ZN(n9774)
         );
  AOI22_X1 U10975 ( .A1(n9772), .A2(n10009), .B1(n9771), .B2(n10010), .ZN(
        n9773) );
  NAND2_X1 U10976 ( .A1(n9774), .A2(n9773), .ZN(n9841) );
  AOI21_X1 U10977 ( .B1(n9775), .B2(n10015), .A(n9841), .ZN(n9776) );
  NOR2_X1 U10978 ( .A1(n9776), .A2(n4984), .ZN(n9777) );
  AOI211_X1 U10979 ( .C1(n9842), .C2(n10031), .A(n9778), .B(n9777), .ZN(n9779)
         );
  OAI21_X1 U10980 ( .B1(n9780), .B2(n9845), .A(n9779), .ZN(P1_U3276) );
  MUX2_X1 U10981 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n9781), .S(n10162), .Z(
        P1_U3553) );
  MUX2_X1 U10982 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n9782), .S(n10162), .Z(
        P1_U3552) );
  MUX2_X1 U10983 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9864), .S(n10162), .Z(
        P1_U3550) );
  OAI21_X1 U10984 ( .B1(n9798), .B2(n9861), .A(n9797), .ZN(n9865) );
  MUX2_X1 U10985 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9865), .S(n10162), .Z(
        P1_U3549) );
  MUX2_X1 U10986 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9866), .S(n10162), .Z(
        P1_U3548) );
  AOI211_X1 U10987 ( .C1(n9858), .C2(n9804), .A(n9803), .B(n9802), .ZN(n9805)
         );
  OAI21_X1 U10988 ( .B1(n9806), .B2(n9861), .A(n9805), .ZN(n9867) );
  MUX2_X1 U10989 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9867), .S(n10162), .Z(
        P1_U3547) );
  AOI211_X1 U10990 ( .C1(n9858), .C2(n9809), .A(n9808), .B(n9807), .ZN(n9810)
         );
  OAI21_X1 U10991 ( .B1(n9811), .B2(n9861), .A(n9810), .ZN(n9868) );
  MUX2_X1 U10992 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9868), .S(n10162), .Z(
        P1_U3546) );
  AOI211_X1 U10993 ( .C1(n9858), .C2(n9814), .A(n9813), .B(n9812), .ZN(n9815)
         );
  OAI21_X1 U10994 ( .B1(n9861), .B2(n9816), .A(n9815), .ZN(n9869) );
  MUX2_X1 U10995 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9869), .S(n10162), .Z(
        P1_U3545) );
  AOI211_X1 U10996 ( .C1(n9858), .C2(n9819), .A(n9818), .B(n9817), .ZN(n9820)
         );
  OAI21_X1 U10997 ( .B1(n9821), .B2(n9861), .A(n9820), .ZN(n9870) );
  MUX2_X1 U10998 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9870), .S(n10162), .Z(
        P1_U3544) );
  AOI211_X1 U10999 ( .C1(n9858), .C2(n9824), .A(n9823), .B(n9822), .ZN(n9825)
         );
  OAI21_X1 U11000 ( .B1(n9826), .B2(n9861), .A(n9825), .ZN(n9871) );
  MUX2_X1 U11001 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9871), .S(n10162), .Z(
        P1_U3543) );
  AOI211_X1 U11002 ( .C1(n9858), .C2(n9829), .A(n9828), .B(n9827), .ZN(n9830)
         );
  OAI21_X1 U11003 ( .B1(n9861), .B2(n9831), .A(n9830), .ZN(n9872) );
  MUX2_X1 U11004 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9872), .S(n10162), .Z(
        P1_U3542) );
  AOI211_X1 U11005 ( .C1(n9858), .C2(n9834), .A(n9833), .B(n9832), .ZN(n9835)
         );
  OAI21_X1 U11006 ( .B1(n9836), .B2(n9861), .A(n9835), .ZN(n9873) );
  MUX2_X1 U11007 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9873), .S(n10162), .Z(
        P1_U3541) );
  AOI21_X1 U11008 ( .B1(n9858), .B2(n7834), .A(n9837), .ZN(n9838) );
  OAI211_X1 U11009 ( .C1(n9840), .C2(n9861), .A(n9839), .B(n9838), .ZN(n9874)
         );
  MUX2_X1 U11010 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9874), .S(n10162), .Z(
        P1_U3540) );
  AOI211_X1 U11011 ( .C1(n9858), .C2(n9843), .A(n9842), .B(n9841), .ZN(n9844)
         );
  OAI21_X1 U11012 ( .B1(n9845), .B2(n9861), .A(n9844), .ZN(n9875) );
  MUX2_X1 U11013 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9875), .S(n10162), .Z(
        P1_U3539) );
  AOI211_X1 U11014 ( .C1(n9858), .C2(n9848), .A(n9847), .B(n9846), .ZN(n9849)
         );
  OAI21_X1 U11015 ( .B1(n9861), .B2(n9850), .A(n9849), .ZN(n9876) );
  MUX2_X1 U11016 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9876), .S(n10162), .Z(
        P1_U3538) );
  AOI21_X1 U11017 ( .B1(n9858), .B2(n9852), .A(n9851), .ZN(n9853) );
  OAI211_X1 U11018 ( .C1(n9861), .C2(n9855), .A(n9854), .B(n9853), .ZN(n9877)
         );
  MUX2_X1 U11019 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n9877), .S(n10162), .Z(
        P1_U3537) );
  AOI21_X1 U11020 ( .B1(n9858), .B2(n9857), .A(n9856), .ZN(n9859) );
  OAI211_X1 U11021 ( .C1(n9862), .C2(n9861), .A(n9860), .B(n9859), .ZN(n9878)
         );
  MUX2_X1 U11022 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n9878), .S(n10162), .Z(
        P1_U3536) );
  MUX2_X1 U11023 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n9864), .S(n10145), .Z(
        P1_U3518) );
  MUX2_X1 U11024 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9865), .S(n10145), .Z(
        P1_U3517) );
  MUX2_X1 U11025 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9866), .S(n10145), .Z(
        P1_U3516) );
  MUX2_X1 U11026 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9867), .S(n10145), .Z(
        P1_U3515) );
  MUX2_X1 U11027 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9868), .S(n10145), .Z(
        P1_U3514) );
  MUX2_X1 U11028 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9869), .S(n10145), .Z(
        P1_U3513) );
  MUX2_X1 U11029 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9870), .S(n10145), .Z(
        P1_U3512) );
  MUX2_X1 U11030 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9871), .S(n10145), .Z(
        P1_U3511) );
  MUX2_X1 U11031 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9872), .S(n10145), .Z(
        P1_U3510) );
  MUX2_X1 U11032 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9873), .S(n10145), .Z(
        P1_U3509) );
  MUX2_X1 U11033 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9874), .S(n10145), .Z(
        P1_U3507) );
  MUX2_X1 U11034 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9875), .S(n10145), .Z(
        P1_U3504) );
  MUX2_X1 U11035 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n9876), .S(n10145), .Z(
        P1_U3501) );
  MUX2_X1 U11036 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n9877), .S(n10145), .Z(
        P1_U3498) );
  MUX2_X1 U11037 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n9878), .S(n10145), .Z(
        P1_U3495) );
  MUX2_X1 U11038 ( .A(P1_D_REG_1__SCAN_IN), .B(n9879), .S(n10076), .Z(P1_U3440) );
  NOR4_X1 U11039 ( .A1(n9881), .A2(P1_IR_REG_30__SCAN_IN), .A3(n5884), .A4(
        P1_U3086), .ZN(n9882) );
  AOI21_X1 U11040 ( .B1(n9894), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9882), .ZN(
        n9883) );
  OAI21_X1 U11041 ( .B1(n9884), .B2(n9897), .A(n9883), .ZN(P1_U3324) );
  AOI22_X1 U11042 ( .A1(n9885), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_30__SCAN_IN), .B2(n9894), .ZN(n9886) );
  OAI21_X1 U11043 ( .B1(n9887), .B2(n9897), .A(n9886), .ZN(P1_U3325) );
  AOI22_X1 U11044 ( .A1(n9888), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n9894), .ZN(n9889) );
  OAI21_X1 U11045 ( .B1(n9890), .B2(n9897), .A(n9889), .ZN(P1_U3326) );
  AOI22_X1 U11046 ( .A1(n9891), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(n9894), .ZN(n9892) );
  OAI21_X1 U11047 ( .B1(n9893), .B2(n9897), .A(n9892), .ZN(P1_U3327) );
  AOI22_X1 U11048 ( .A1(n9895), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(n9894), .ZN(n9896) );
  OAI21_X1 U11049 ( .B1(n9898), .B2(n9897), .A(n9896), .ZN(P1_U3328) );
  MUX2_X1 U11050 ( .A(n9899), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  XNOR2_X1 U11051 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U11052 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  INV_X1 U11053 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n9911) );
  AOI211_X1 U11054 ( .C1(n9902), .C2(n9901), .A(n9928), .B(n9900), .ZN(n9907)
         );
  AOI211_X1 U11055 ( .C1(n9905), .C2(n9904), .A(n9915), .B(n9903), .ZN(n9906)
         );
  AOI211_X1 U11056 ( .C1(n9959), .C2(n9908), .A(n9907), .B(n9906), .ZN(n9910)
         );
  OAI211_X1 U11057 ( .C1(n9970), .C2(n9911), .A(n9910), .B(n9909), .ZN(
        P1_U3257) );
  INV_X1 U11058 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n9924) );
  AOI211_X1 U11059 ( .C1(n9914), .C2(n9913), .A(n9912), .B(n9928), .ZN(n9920)
         );
  AOI211_X1 U11060 ( .C1(n9918), .C2(n9917), .A(n9916), .B(n9915), .ZN(n9919)
         );
  AOI211_X1 U11061 ( .C1(n9959), .C2(n9921), .A(n9920), .B(n9919), .ZN(n9923)
         );
  OAI211_X1 U11062 ( .C1(n9970), .C2(n9924), .A(n9923), .B(n9922), .ZN(
        P1_U3258) );
  OAI21_X1 U11063 ( .B1(n9927), .B2(n9926), .A(n9925), .ZN(n9934) );
  NOR2_X1 U11064 ( .A1(n9948), .A2(n4418), .ZN(n9933) );
  AOI211_X1 U11065 ( .C1(n9931), .C2(n9930), .A(n9929), .B(n9928), .ZN(n9932)
         );
  AOI211_X1 U11066 ( .C1(n9964), .C2(n9934), .A(n9933), .B(n9932), .ZN(n9936)
         );
  OAI211_X1 U11067 ( .C1(n9970), .C2(n9937), .A(n9936), .B(n9935), .ZN(
        P1_U3259) );
  INV_X1 U11068 ( .A(n9938), .ZN(n9947) );
  XNOR2_X1 U11069 ( .A(n9940), .B(n9939), .ZN(n9941) );
  NAND2_X1 U11070 ( .A1(n9957), .A2(n9941), .ZN(n9946) );
  XNOR2_X1 U11071 ( .A(n9943), .B(n9942), .ZN(n9944) );
  NAND2_X1 U11072 ( .A1(n9964), .A2(n9944), .ZN(n9945) );
  OAI211_X1 U11073 ( .C1(n9948), .C2(n9947), .A(n9946), .B(n9945), .ZN(n9949)
         );
  INV_X1 U11074 ( .A(n9949), .ZN(n9951) );
  OAI211_X1 U11075 ( .C1(n9952), .C2(n9970), .A(n9951), .B(n9950), .ZN(
        P1_U3260) );
  NAND2_X1 U11076 ( .A1(n9954), .A2(n9953), .ZN(n9955) );
  NAND3_X1 U11077 ( .A1(n9957), .A2(n9956), .A3(n9955), .ZN(n9967) );
  NAND2_X1 U11078 ( .A1(n9959), .A2(n9958), .ZN(n9966) );
  NAND2_X1 U11079 ( .A1(n9961), .A2(n9960), .ZN(n9962) );
  NAND3_X1 U11080 ( .A1(n9964), .A2(n9963), .A3(n9962), .ZN(n9965) );
  OAI211_X1 U11081 ( .C1(n9970), .C2(n10196), .A(n9969), .B(n9968), .ZN(
        P1_U3261) );
  NAND2_X1 U11082 ( .A1(n9972), .A2(n9971), .ZN(n9973) );
  XNOR2_X1 U11083 ( .A(n9973), .B(n9976), .ZN(n10128) );
  OAI22_X1 U11084 ( .A1(n10050), .A2(n9975), .B1(n9974), .B2(n10048), .ZN(
        n9980) );
  XNOR2_X1 U11085 ( .A(n9977), .B(n9976), .ZN(n9978) );
  NOR2_X1 U11086 ( .A1(n9978), .A2(n10047), .ZN(n9979) );
  AOI211_X1 U11087 ( .C1(n9981), .C2(n10128), .A(n9980), .B(n9979), .ZN(n10125) );
  INV_X1 U11088 ( .A(n9982), .ZN(n9983) );
  AOI222_X1 U11089 ( .A1(n10122), .A2(n10017), .B1(P1_REG2_REG_8__SCAN_IN), 
        .B2(n4984), .C1(n9983), .C2(n10015), .ZN(n9990) );
  INV_X1 U11090 ( .A(n9984), .ZN(n9987) );
  AOI21_X1 U11091 ( .B1(n9985), .B2(n10122), .A(n10039), .ZN(n9986) );
  NAND2_X1 U11092 ( .A1(n9987), .A2(n9986), .ZN(n10123) );
  INV_X1 U11093 ( .A(n10123), .ZN(n9988) );
  AOI22_X1 U11094 ( .A1(n10031), .A2(n9988), .B1(n10128), .B2(n10055), .ZN(
        n9989) );
  OAI211_X1 U11095 ( .C1(n4984), .C2(n10125), .A(n9990), .B(n9989), .ZN(
        P1_U3285) );
  XNOR2_X1 U11096 ( .A(n9999), .B(n9991), .ZN(n9993) );
  AOI222_X1 U11097 ( .A1(n10013), .A2(n9993), .B1(n9992), .B2(n10009), .C1(
        n7358), .C2(n10010), .ZN(n10110) );
  INV_X1 U11098 ( .A(n9994), .ZN(n9995) );
  AOI222_X1 U11099 ( .A1(n10001), .A2(n10017), .B1(P1_REG2_REG_6__SCAN_IN), 
        .B2(n4984), .C1(n10015), .C2(n9995), .ZN(n10006) );
  OAI21_X1 U11100 ( .B1(n9997), .B2(n7373), .A(n9996), .ZN(n9998) );
  XNOR2_X1 U11101 ( .A(n9999), .B(n9998), .ZN(n10113) );
  INV_X1 U11102 ( .A(n10000), .ZN(n10003) );
  OAI211_X1 U11103 ( .C1(n10003), .C2(n7360), .A(n10027), .B(n10002), .ZN(
        n10109) );
  INV_X1 U11104 ( .A(n10109), .ZN(n10004) );
  AOI22_X1 U11105 ( .A1(n10113), .A2(n10032), .B1(n10031), .B2(n10004), .ZN(
        n10005) );
  OAI211_X1 U11106 ( .C1(n4984), .C2(n10110), .A(n10006), .B(n10005), .ZN(
        P1_U3287) );
  OAI21_X1 U11107 ( .B1(n7487), .B2(n10021), .A(n10007), .ZN(n10008) );
  XOR2_X1 U11108 ( .A(n10024), .B(n10008), .Z(n10012) );
  AOI222_X1 U11109 ( .A1(n10013), .A2(n10012), .B1(n10011), .B2(n10010), .C1(
        n7358), .C2(n10009), .ZN(n10097) );
  INV_X1 U11110 ( .A(n10014), .ZN(n10016) );
  AOI222_X1 U11111 ( .A1(n10018), .A2(n10017), .B1(P1_REG2_REG_4__SCAN_IN), 
        .B2(n4984), .C1(n10016), .C2(n10015), .ZN(n10034) );
  INV_X1 U11112 ( .A(n10019), .ZN(n10020) );
  AOI21_X1 U11113 ( .B1(n10022), .B2(n10021), .A(n10020), .ZN(n10023) );
  XOR2_X1 U11114 ( .A(n10024), .B(n10023), .Z(n10100) );
  INV_X1 U11115 ( .A(n10025), .ZN(n10029) );
  INV_X1 U11116 ( .A(n10026), .ZN(n10028) );
  OAI211_X1 U11117 ( .C1(n10096), .C2(n10029), .A(n10028), .B(n10027), .ZN(
        n10095) );
  INV_X1 U11118 ( .A(n10095), .ZN(n10030) );
  AOI22_X1 U11119 ( .A1(n10100), .A2(n10032), .B1(n10031), .B2(n10030), .ZN(
        n10033) );
  OAI211_X1 U11120 ( .C1(n4984), .C2(n10097), .A(n10034), .B(n10033), .ZN(
        P1_U3289) );
  AOI22_X1 U11121 ( .A1(n10036), .A2(n10035), .B1(n4441), .B2(n4405), .ZN(
        n10037) );
  XNOR2_X1 U11122 ( .A(n10045), .B(n10037), .ZN(n10054) );
  AOI211_X1 U11123 ( .C1(n7353), .C2(n10040), .A(n10039), .B(n10038), .ZN(
        n10084) );
  INV_X1 U11124 ( .A(n10041), .ZN(n10042) );
  OAI22_X1 U11125 ( .A1(n10068), .A2(n10043), .B1(n10042), .B2(n10086), .ZN(
        n10051) );
  XNOR2_X1 U11126 ( .A(n10044), .B(n10045), .ZN(n10046) );
  OAI222_X1 U11127 ( .A1(n10050), .A2(n4441), .B1(n10048), .B2(n7344), .C1(
        n10047), .C2(n10046), .ZN(n10087) );
  AOI211_X1 U11128 ( .C1(n10084), .C2(n6294), .A(n10051), .B(n10087), .ZN(
        n10052) );
  OAI21_X1 U11129 ( .B1(n10053), .B2(n10054), .A(n10052), .ZN(n10056) );
  INV_X1 U11130 ( .A(n10054), .ZN(n10089) );
  AOI22_X1 U11131 ( .A1(n10056), .A2(n10070), .B1(n10089), .B2(n10055), .ZN(
        n10057) );
  OAI21_X1 U11132 ( .B1(n5952), .B2(n10070), .A(n10057), .ZN(P1_U3291) );
  NAND2_X1 U11133 ( .A1(n7000), .A2(n10058), .ZN(n10059) );
  NOR2_X1 U11134 ( .A1(n10062), .A2(n10059), .ZN(n10060) );
  NOR2_X1 U11135 ( .A1(n10061), .A2(n10060), .ZN(n10066) );
  NAND3_X1 U11136 ( .A1(n10064), .A2(n10063), .A3(n10062), .ZN(n10065) );
  OAI211_X1 U11137 ( .C1(n10068), .C2(n10067), .A(n10066), .B(n10065), .ZN(
        n10069) );
  INV_X1 U11138 ( .A(n10069), .ZN(n10071) );
  AOI22_X1 U11139 ( .A1(n4984), .A2(n5921), .B1(n10071), .B2(n10070), .ZN(
        P1_U3293) );
  AND2_X1 U11140 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n10074), .ZN(P1_U3294) );
  AND2_X1 U11141 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n10074), .ZN(P1_U3295) );
  AND2_X1 U11142 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n10074), .ZN(P1_U3296) );
  NOR2_X1 U11143 ( .A1(n10076), .A2(n10072), .ZN(P1_U3297) );
  AND2_X1 U11144 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n10074), .ZN(P1_U3298) );
  AND2_X1 U11145 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n10074), .ZN(P1_U3299) );
  AND2_X1 U11146 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n10074), .ZN(P1_U3300) );
  AND2_X1 U11147 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n10074), .ZN(P1_U3301) );
  AND2_X1 U11148 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n10074), .ZN(P1_U3302) );
  AND2_X1 U11149 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n10074), .ZN(P1_U3303) );
  AND2_X1 U11150 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n10074), .ZN(P1_U3304) );
  AND2_X1 U11151 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n10074), .ZN(P1_U3305) );
  AND2_X1 U11152 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n10074), .ZN(P1_U3306) );
  AND2_X1 U11153 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n10074), .ZN(P1_U3307) );
  AND2_X1 U11154 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n10074), .ZN(P1_U3308) );
  AND2_X1 U11155 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n10074), .ZN(P1_U3309) );
  AND2_X1 U11156 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n10074), .ZN(P1_U3310) );
  AND2_X1 U11157 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n10074), .ZN(P1_U3311) );
  NOR2_X1 U11158 ( .A1(n10076), .A2(n10073), .ZN(P1_U3312) );
  AND2_X1 U11159 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n10074), .ZN(P1_U3313) );
  AND2_X1 U11160 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n10074), .ZN(P1_U3314) );
  AND2_X1 U11161 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n10074), .ZN(P1_U3315) );
  AND2_X1 U11162 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n10074), .ZN(P1_U3316) );
  AND2_X1 U11163 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n10074), .ZN(P1_U3317) );
  AND2_X1 U11164 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n10074), .ZN(P1_U3318) );
  AND2_X1 U11165 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n10074), .ZN(P1_U3319) );
  AND2_X1 U11166 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n10074), .ZN(P1_U3320) );
  AND2_X1 U11167 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n10074), .ZN(P1_U3321) );
  AND2_X1 U11168 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n10074), .ZN(P1_U3322) );
  NOR2_X1 U11169 ( .A1(n10076), .A2(n10075), .ZN(P1_U3323) );
  AOI22_X1 U11170 ( .A1(n10145), .A2(n10077), .B1(n5922), .B2(n10144), .ZN(
        P1_U3453) );
  INV_X1 U11171 ( .A(n10078), .ZN(n10129) );
  OAI21_X1 U11172 ( .B1(n4405), .B2(n10139), .A(n10079), .ZN(n10082) );
  INV_X1 U11173 ( .A(n10080), .ZN(n10081) );
  AOI211_X1 U11174 ( .C1(n10129), .C2(n10083), .A(n10082), .B(n10081), .ZN(
        n10147) );
  AOI22_X1 U11175 ( .A1(n10145), .A2(n10147), .B1(n5914), .B2(n10144), .ZN(
        P1_U3456) );
  INV_X1 U11176 ( .A(n10084), .ZN(n10085) );
  OAI21_X1 U11177 ( .B1(n10086), .B2(n10139), .A(n10085), .ZN(n10088) );
  AOI211_X1 U11178 ( .C1(n10089), .C2(n10136), .A(n10088), .B(n10087), .ZN(
        n10149) );
  AOI22_X1 U11179 ( .A1(n10145), .A2(n10149), .B1(n5953), .B2(n10144), .ZN(
        P1_U3459) );
  OAI211_X1 U11180 ( .C1(n10092), .C2(n10139), .A(n10091), .B(n10090), .ZN(
        n10093) );
  AOI21_X1 U11181 ( .B1(n10136), .B2(n10094), .A(n10093), .ZN(n10150) );
  AOI22_X1 U11182 ( .A1(n10145), .A2(n10150), .B1(n5973), .B2(n10144), .ZN(
        P1_U3462) );
  OAI21_X1 U11183 ( .B1(n10096), .B2(n10139), .A(n10095), .ZN(n10099) );
  INV_X1 U11184 ( .A(n10097), .ZN(n10098) );
  AOI211_X1 U11185 ( .C1(n10136), .C2(n10100), .A(n10099), .B(n10098), .ZN(
        n10152) );
  INV_X1 U11186 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n10101) );
  AOI22_X1 U11187 ( .A1(n10145), .A2(n10152), .B1(n10101), .B2(n10144), .ZN(
        P1_U3465) );
  INV_X1 U11188 ( .A(n10102), .ZN(n10106) );
  OAI21_X1 U11189 ( .B1(n10104), .B2(n10139), .A(n10103), .ZN(n10105) );
  AOI21_X1 U11190 ( .B1(n10106), .B2(n10136), .A(n10105), .ZN(n10107) );
  AND2_X1 U11191 ( .A1(n10108), .A2(n10107), .ZN(n10154) );
  AOI22_X1 U11192 ( .A1(n10145), .A2(n10154), .B1(n6012), .B2(n10144), .ZN(
        P1_U3468) );
  OAI21_X1 U11193 ( .B1(n7360), .B2(n10139), .A(n10109), .ZN(n10112) );
  INV_X1 U11194 ( .A(n10110), .ZN(n10111) );
  AOI211_X1 U11195 ( .C1(n10136), .C2(n10113), .A(n10112), .B(n10111), .ZN(
        n10155) );
  INV_X1 U11196 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n10114) );
  AOI22_X1 U11197 ( .A1(n10145), .A2(n10155), .B1(n10114), .B2(n10144), .ZN(
        P1_U3471) );
  INV_X1 U11198 ( .A(n10115), .ZN(n10120) );
  OAI21_X1 U11199 ( .B1(n10117), .B2(n10139), .A(n10116), .ZN(n10119) );
  AOI211_X1 U11200 ( .C1(n10129), .C2(n10120), .A(n10119), .B(n10118), .ZN(
        n10156) );
  INV_X1 U11201 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n10121) );
  AOI22_X1 U11202 ( .A1(n10145), .A2(n10156), .B1(n10121), .B2(n10144), .ZN(
        P1_U3474) );
  INV_X1 U11203 ( .A(n10122), .ZN(n10124) );
  OAI21_X1 U11204 ( .B1(n10124), .B2(n10139), .A(n10123), .ZN(n10127) );
  INV_X1 U11205 ( .A(n10125), .ZN(n10126) );
  AOI211_X1 U11206 ( .C1(n10129), .C2(n10128), .A(n10127), .B(n10126), .ZN(
        n10158) );
  AOI22_X1 U11207 ( .A1(n10145), .A2(n10158), .B1(n6101), .B2(n10144), .ZN(
        P1_U3477) );
  OAI21_X1 U11208 ( .B1(n10131), .B2(n10139), .A(n10130), .ZN(n10133) );
  AOI211_X1 U11209 ( .C1(n10136), .C2(n10134), .A(n10133), .B(n10132), .ZN(
        n10159) );
  INV_X1 U11210 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n10135) );
  AOI22_X1 U11211 ( .A1(n10145), .A2(n10159), .B1(n10135), .B2(n10144), .ZN(
        P1_U3480) );
  AND2_X1 U11212 ( .A1(n10137), .A2(n10136), .ZN(n10142) );
  OAI21_X1 U11213 ( .B1(n10140), .B2(n10139), .A(n10138), .ZN(n10141) );
  NOR3_X1 U11214 ( .A1(n10143), .A2(n10142), .A3(n10141), .ZN(n10161) );
  AOI22_X1 U11215 ( .A1(n10145), .A2(n10161), .B1(n6143), .B2(n10144), .ZN(
        P1_U3483) );
  INV_X1 U11216 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n10146) );
  AOI22_X1 U11217 ( .A1(n10162), .A2(n10147), .B1(n10146), .B2(n10160), .ZN(
        P1_U3523) );
  AOI22_X1 U11218 ( .A1(n10162), .A2(n10149), .B1(n10148), .B2(n10160), .ZN(
        P1_U3524) );
  AOI22_X1 U11219 ( .A1(n10162), .A2(n10150), .B1(n6589), .B2(n10160), .ZN(
        P1_U3525) );
  AOI22_X1 U11220 ( .A1(n10162), .A2(n10152), .B1(n10151), .B2(n10160), .ZN(
        P1_U3526) );
  INV_X1 U11221 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n10153) );
  AOI22_X1 U11222 ( .A1(n10162), .A2(n10154), .B1(n10153), .B2(n10160), .ZN(
        P1_U3527) );
  AOI22_X1 U11223 ( .A1(n10162), .A2(n10155), .B1(n6042), .B2(n10160), .ZN(
        P1_U3528) );
  AOI22_X1 U11224 ( .A1(n10162), .A2(n10156), .B1(n6591), .B2(n10160), .ZN(
        P1_U3529) );
  INV_X1 U11225 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n10157) );
  AOI22_X1 U11226 ( .A1(n10162), .A2(n10158), .B1(n10157), .B2(n10160), .ZN(
        P1_U3530) );
  AOI22_X1 U11227 ( .A1(n10162), .A2(n10159), .B1(n6592), .B2(n10160), .ZN(
        P1_U3531) );
  AOI22_X1 U11228 ( .A1(n10162), .A2(n10161), .B1(n6593), .B2(n10160), .ZN(
        P1_U3532) );
  OAI22_X1 U11229 ( .A1(n10166), .A2(n10165), .B1(n10164), .B2(n10163), .ZN(
        n10168) );
  AOI211_X1 U11230 ( .C1(n10170), .C2(n10169), .A(n10168), .B(n10167), .ZN(
        n10172) );
  AOI22_X1 U11231 ( .A1(n10174), .A2(n10173), .B1(n10172), .B2(n10171), .ZN(
        P2_U3231) );
  AOI22_X1 U11232 ( .A1(n10188), .A2(n10176), .B1(n10175), .B2(n10185), .ZN(
        P2_U3396) );
  INV_X1 U11233 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n10178) );
  AOI22_X1 U11234 ( .A1(n10188), .A2(n10178), .B1(n10177), .B2(n10185), .ZN(
        P2_U3399) );
  INV_X1 U11235 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n10180) );
  AOI22_X1 U11236 ( .A1(n10188), .A2(n10180), .B1(n10179), .B2(n10185), .ZN(
        P2_U3402) );
  INV_X1 U11237 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n10182) );
  AOI22_X1 U11238 ( .A1(n10188), .A2(n10182), .B1(n10181), .B2(n10185), .ZN(
        P2_U3405) );
  INV_X1 U11239 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10184) );
  AOI22_X1 U11240 ( .A1(n10188), .A2(n10184), .B1(n10183), .B2(n10185), .ZN(
        P2_U3408) );
  AOI22_X1 U11241 ( .A1(n10188), .A2(n10187), .B1(n10186), .B2(n10185), .ZN(
        P2_U3411) );
  OAI222_X1 U11242 ( .A1(n10193), .A2(n10192), .B1(n10193), .B2(n10191), .C1(
        n10190), .C2(n10189), .ZN(ADD_1068_U5) );
  XOR2_X1 U11243 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1068_U46) );
  AOI21_X1 U11244 ( .B1(n10196), .B2(n10195), .A(n10194), .ZN(n10197) );
  XOR2_X1 U11245 ( .A(P2_ADDR_REG_18__SCAN_IN), .B(n10197), .Z(ADD_1068_U55)
         );
  OAI21_X1 U11246 ( .B1(n10200), .B2(n10199), .A(n10198), .ZN(ADD_1068_U56) );
  OAI21_X1 U11247 ( .B1(n10203), .B2(n10202), .A(n10201), .ZN(ADD_1068_U57) );
  OAI21_X1 U11248 ( .B1(n10206), .B2(n10205), .A(n10204), .ZN(ADD_1068_U58) );
  OAI21_X1 U11249 ( .B1(n10209), .B2(n10208), .A(n10207), .ZN(ADD_1068_U59) );
  OAI21_X1 U11250 ( .B1(n10212), .B2(n10211), .A(n10210), .ZN(ADD_1068_U60) );
  OAI21_X1 U11251 ( .B1(n10215), .B2(n10214), .A(n10213), .ZN(ADD_1068_U61) );
  OAI21_X1 U11252 ( .B1(n10218), .B2(n10217), .A(n10216), .ZN(ADD_1068_U62) );
  OAI21_X1 U11253 ( .B1(n10221), .B2(n10220), .A(n10219), .ZN(ADD_1068_U63) );
  OAI21_X1 U11254 ( .B1(n10224), .B2(n10223), .A(n10222), .ZN(ADD_1068_U50) );
  OAI21_X1 U11255 ( .B1(n10227), .B2(n10226), .A(n10225), .ZN(ADD_1068_U51) );
  OAI21_X1 U11256 ( .B1(n10230), .B2(n10229), .A(n10228), .ZN(ADD_1068_U47) );
  OAI21_X1 U11257 ( .B1(n10233), .B2(n10232), .A(n10231), .ZN(ADD_1068_U49) );
  OAI21_X1 U11258 ( .B1(n10236), .B2(n10235), .A(n10234), .ZN(ADD_1068_U48) );
  AOI21_X1 U11259 ( .B1(n10239), .B2(n10238), .A(n10237), .ZN(ADD_1068_U54) );
  AOI21_X1 U11260 ( .B1(n10242), .B2(n10241), .A(n10240), .ZN(ADD_1068_U53) );
  OAI21_X1 U11261 ( .B1(n10245), .B2(n10244), .A(n10243), .ZN(ADD_1068_U52) );
  BUF_X2 U5027 ( .A(n5992), .Z(n6442) );
  INV_X1 U7804 ( .A(n7586), .ZN(n9499) );
  CLKBUF_X1 U4789 ( .A(n5835), .Z(n5860) );
  CLKBUF_X1 U4812 ( .A(n5387), .Z(n8452) );
  CLKBUF_X1 U4813 ( .A(n9751), .Z(n4404) );
  OR2_X2 U4834 ( .A1(n10002), .A2(n7429), .ZN(n9985) );
  CLKBUF_X1 U4846 ( .A(P2_IR_REG_8__SCAN_IN), .Z(n9109) );
  NAND2_X1 U4851 ( .A1(n5035), .A2(n4938), .ZN(n5034) );
  CLKBUF_X1 U4892 ( .A(n9337), .Z(n4423) );
  INV_X1 U5214 ( .A(n6041), .ZN(n7247) );
  CLKBUF_X1 U5291 ( .A(n6041), .Z(n6323) );
  OR2_X2 U5357 ( .A1(n9885), .A2(n9888), .ZN(n5991) );
  CLKBUF_X1 U5785 ( .A(n6484), .Z(n6828) );
  CLKBUF_X1 U6575 ( .A(n8799), .Z(n4470) );
  CLKBUF_X1 U6687 ( .A(n5307), .Z(n6778) );
  NAND2_X1 U7177 ( .A1(n5855), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5852) );
  CLKBUF_X1 U7677 ( .A(n5312), .Z(n4274) );
endmodule

