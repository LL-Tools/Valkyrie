

module b21_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, P2_WR_REG_SCAN_IN, SI_31_, 
        SI_30_, SI_29_, SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, 
        SI_21_, SI_20_, SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, 
        SI_12_, SI_11_, SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, 
        SI_3_, SI_2_, SI_1_, SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, 
        ADD_1071_U57, ADD_1071_U58, ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, 
        ADD_1071_U62, ADD_1071_U63, ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, 
        ADD_1071_U50, ADD_1071_U51, ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, 
        ADD_1071_U5, ADD_1071_U46, U126, U123, P1_U3353, P1_U3352, P1_U3351, 
        P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, 
        P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, 
        P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, 
        P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, 
        P1_U3322, P1_U3440, P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, 
        P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, 
        P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, 
        P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, 
        P1_U3296, P1_U3295, P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, 
        P1_U3460, P1_U3463, P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, 
        P1_U3481, P1_U3484, P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, 
        P1_U3502, P1_U3505, P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, 
        P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, 
        P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, 
        P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, 
        P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, 
        P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, 
        P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, 
        P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, 
        P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, 
        P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, 
        P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, 
        P1_U3355, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, 
        P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, 
        P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, 
        P1_U3242, P1_U3241, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, 
        P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, 
        P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, 
        P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, 
        P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, 
        P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, 
        P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, 
        P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, 
        P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, 
        P1_U3211, P1_U3084, P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, 
        P2_U3355, P2_U3354, P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, 
        P2_U3348, P2_U3347, P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, 
        P2_U3341, P2_U3340, P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, 
        P2_U3334, P2_U3333, P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, 
        P2_U3327, P2_U3437, P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, 
        P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, 
        P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, 
        P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, 
        P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, 
        P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, 
        P2_U3478, P2_U3481, P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, 
        P2_U3499, P2_U3502, P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, 
        P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, 
        P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, 
        P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, 
        P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, 
        P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, 
        P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, 
        P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, 
        P2_U3564, P2_U3565, P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, 
        P2_U3571, P2_U3572, P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, 
        P2_U3578, P2_U3579, P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, 
        P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3152, P2_U3151, P2_U3966 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_,
         SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_,
         SI_20_, SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_,
         SI_12_, SI_11_, SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_,
         SI_3_, SI_2_, SI_1_, SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_REG3_REG_7__SCAN_IN, P2_REG3_REG_27__SCAN_IN,
         P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_23__SCAN_IN,
         P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_3__SCAN_IN,
         P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_28__SCAN_IN,
         P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_1__SCAN_IN,
         P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_12__SCAN_IN,
         P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_16__SCAN_IN,
         P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_17__SCAN_IN,
         P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_4__SCAN_IN,
         P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN,
         P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN,
         P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN,
         P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN,
         P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN,
         P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4848, n4849, n4850, n4851, n4852, n4854, n4855, n4856, n4857, n4858,
         n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868,
         n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878,
         n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888,
         n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898,
         n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908,
         n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918,
         n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928,
         n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938,
         n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948,
         n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958,
         n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968,
         n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978,
         n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988,
         n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998,
         n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008,
         n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018,
         n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028,
         n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038,
         n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048,
         n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058,
         n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068,
         n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078,
         n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088,
         n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098,
         n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108,
         n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118,
         n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128,
         n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138,
         n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148,
         n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158,
         n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168,
         n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178,
         n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188,
         n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198,
         n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208,
         n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218,
         n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228,
         n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238,
         n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248,
         n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258,
         n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268,
         n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278,
         n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288,
         n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298,
         n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308,
         n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318,
         n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328,
         n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338,
         n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348,
         n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358,
         n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368,
         n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378,
         n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388,
         n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398,
         n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408,
         n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418,
         n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428,
         n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438,
         n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448,
         n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458,
         n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468,
         n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478,
         n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488,
         n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498,
         n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508,
         n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518,
         n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528,
         n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538,
         n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548,
         n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558,
         n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568,
         n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578,
         n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588,
         n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598,
         n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608,
         n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618,
         n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628,
         n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638,
         n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648,
         n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658,
         n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668,
         n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678,
         n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688,
         n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698,
         n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708,
         n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718,
         n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728,
         n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738,
         n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748,
         n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758,
         n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768,
         n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778,
         n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788,
         n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798,
         n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808,
         n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818,
         n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828,
         n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838,
         n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848,
         n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858,
         n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868,
         n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878,
         n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888,
         n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898,
         n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908,
         n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918,
         n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928,
         n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938,
         n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948,
         n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958,
         n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968,
         n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978,
         n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988,
         n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998,
         n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008,
         n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018,
         n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028,
         n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038,
         n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048,
         n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058,
         n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068,
         n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078,
         n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088,
         n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098,
         n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108,
         n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118,
         n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128,
         n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138,
         n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148,
         n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158,
         n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168,
         n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178,
         n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188,
         n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198,
         n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208,
         n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218,
         n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228,
         n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238,
         n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248,
         n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258,
         n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268,
         n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278,
         n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288,
         n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298,
         n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308,
         n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318,
         n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328,
         n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338,
         n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348,
         n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358,
         n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368,
         n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378,
         n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388,
         n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398,
         n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408,
         n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418,
         n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428,
         n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438,
         n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448,
         n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458,
         n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468,
         n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478,
         n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488,
         n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498,
         n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508,
         n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518,
         n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528,
         n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538,
         n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548,
         n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558,
         n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568,
         n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578,
         n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588,
         n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598,
         n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608,
         n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618,
         n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628,
         n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638,
         n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648,
         n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658,
         n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668,
         n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678,
         n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688,
         n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698,
         n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708,
         n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718,
         n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728,
         n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738,
         n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748,
         n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758,
         n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768,
         n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778,
         n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788,
         n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798,
         n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808,
         n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818,
         n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828,
         n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838,
         n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848,
         n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858,
         n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868,
         n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878,
         n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888,
         n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898,
         n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908,
         n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918,
         n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928,
         n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938,
         n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948,
         n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958,
         n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968,
         n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978,
         n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988,
         n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998,
         n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008,
         n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018,
         n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028,
         n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038,
         n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048,
         n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058,
         n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068,
         n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078,
         n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088,
         n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098,
         n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108,
         n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118,
         n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128,
         n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138,
         n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148,
         n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158,
         n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168,
         n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178,
         n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188,
         n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198,
         n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208,
         n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218,
         n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228,
         n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238,
         n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248,
         n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258,
         n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268,
         n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278,
         n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288,
         n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298,
         n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308,
         n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318,
         n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328,
         n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338,
         n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348,
         n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358,
         n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368,
         n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378,
         n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388,
         n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398,
         n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408,
         n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418,
         n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428,
         n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438,
         n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448,
         n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458,
         n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468,
         n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478,
         n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488,
         n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498,
         n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508,
         n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518,
         n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528,
         n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538,
         n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548,
         n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558,
         n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568,
         n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578,
         n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588,
         n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598,
         n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608,
         n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618,
         n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628,
         n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638,
         n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648,
         n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658,
         n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668,
         n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678,
         n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688,
         n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698,
         n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708,
         n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718,
         n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728,
         n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738,
         n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748,
         n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758,
         n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768,
         n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778,
         n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788,
         n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798,
         n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808,
         n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818,
         n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828,
         n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838,
         n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848,
         n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858,
         n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868,
         n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878,
         n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888,
         n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898,
         n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908,
         n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918,
         n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928,
         n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938,
         n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948,
         n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958,
         n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968,
         n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978,
         n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988,
         n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998,
         n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008,
         n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018,
         n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028,
         n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038,
         n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048,
         n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058,
         n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068,
         n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078,
         n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088,
         n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098,
         n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108,
         n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118,
         n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128,
         n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138,
         n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148,
         n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158,
         n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168,
         n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178,
         n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188,
         n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198,
         n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208,
         n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218,
         n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228,
         n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238,
         n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248,
         n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258,
         n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268,
         n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278,
         n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288,
         n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298,
         n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308,
         n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318,
         n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328,
         n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338,
         n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348,
         n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358,
         n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368,
         n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378,
         n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388,
         n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398,
         n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408,
         n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418,
         n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428,
         n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438,
         n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448,
         n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458,
         n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468,
         n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478,
         n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488,
         n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498,
         n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508,
         n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518,
         n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528,
         n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538,
         n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548,
         n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558,
         n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568,
         n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578,
         n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588,
         n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598,
         n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608,
         n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618,
         n8619, n8620, n8621, n8622, n8623, n8625, n8626, n8627, n8628, n8629,
         n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639,
         n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649,
         n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659,
         n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669,
         n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679,
         n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689,
         n8690, n8691, n8692, n8693, n8694, n8696, n8697, n8698, n8699, n8700,
         n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710,
         n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720,
         n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730,
         n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740,
         n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750,
         n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760,
         n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770,
         n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780,
         n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790,
         n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800,
         n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810,
         n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820,
         n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830,
         n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840,
         n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850,
         n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860,
         n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870,
         n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880,
         n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890,
         n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900,
         n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910,
         n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920,
         n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930,
         n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940,
         n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950,
         n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960,
         n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970,
         n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980,
         n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990,
         n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000,
         n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010,
         n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020,
         n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030,
         n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040,
         n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050,
         n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060,
         n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070,
         n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080,
         n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090,
         n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100,
         n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110,
         n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120,
         n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130,
         n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140,
         n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150,
         n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160,
         n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170,
         n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180,
         n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190,
         n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200,
         n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210,
         n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220,
         n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230,
         n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240,
         n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250,
         n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260,
         n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270,
         n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280,
         n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290,
         n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300,
         n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310,
         n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320,
         n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330,
         n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340,
         n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350,
         n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360,
         n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370,
         n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380,
         n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390,
         n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400,
         n9401, n9402, n9403, n9405, n9406, n9407, n9408, n9409, n9410, n9411,
         n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421,
         n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431,
         n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441,
         n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451,
         n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461,
         n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471,
         n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481,
         n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491,
         n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501,
         n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511,
         n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521,
         n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531,
         n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541,
         n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551,
         n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561,
         n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571,
         n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581,
         n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591,
         n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601,
         n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611,
         n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621,
         n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631,
         n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641,
         n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651,
         n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661,
         n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671,
         n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681,
         n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691,
         n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701,
         n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711,
         n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721,
         n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731,
         n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741,
         n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751,
         n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761,
         n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771,
         n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781,
         n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791,
         n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801,
         n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811,
         n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821,
         n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831,
         n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841,
         n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851,
         n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861,
         n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871,
         n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881,
         n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891,
         n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901,
         n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911,
         n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921,
         n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931,
         n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941,
         n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951,
         n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961,
         n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971,
         n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981,
         n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991,
         n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
         n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
         n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296,
         n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304,
         n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
         n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320,
         n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328,
         n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336,
         n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344,
         n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352,
         n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360,
         n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368,
         n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376,
         n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384,
         n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392,
         n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400,
         n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408,
         n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416,
         n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424,
         n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432,
         n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440,
         n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448,
         n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456,
         n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464,
         n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472,
         n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480,
         n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488,
         n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496,
         n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504,
         n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512,
         n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520,
         n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528,
         n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536,
         n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544,
         n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552,
         n10553, n10554, n10555, n10556, n10557;

  AND2_X1 U4913 ( .A1(n5807), .A2(n9305), .ZN(n5830) );
  NAND2_X2 U4914 ( .A1(n9571), .A2(n9569), .ZN(n9889) );
  AND3_X1 U4915 ( .A1(n7907), .A2(n5623), .A3(n5622), .ZN(n5626) );
  NAND2_X1 U4916 ( .A1(n9551), .A2(n9553), .ZN(n9670) );
  CLKBUF_X2 U4917 ( .A(n7068), .Z(n8543) );
  INV_X2 U4918 ( .A(n6081), .ZN(n6765) );
  OR2_X1 U4919 ( .A1(n5814), .A2(n5813), .ZN(n5815) );
  NOR2_X2 U4920 ( .A1(n9658), .A2(n9459), .ZN(n6150) );
  NAND4_X1 U4921 ( .A1(n5508), .A2(n5507), .A3(n5506), .A4(n5505), .ZN(n9717)
         );
  INV_X1 U4922 ( .A(n6348), .ZN(n7304) );
  INV_X1 U4923 ( .A(n10411), .ZN(n9856) );
  INV_X1 U4924 ( .A(n7139), .ZN(n7138) );
  CLKBUF_X2 U4925 ( .A(n5473), .Z(n7139) );
  NOR2_X1 U4926 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n6289) );
  OR2_X1 U4927 ( .A1(n6157), .A2(n9978), .ZN(n9556) );
  NOR2_X1 U4928 ( .A1(n7045), .A2(n8542), .ZN(n7047) );
  INV_X1 U4929 ( .A(n7658), .ZN(n7231) );
  INV_X1 U4930 ( .A(n6762), .ZN(n6767) );
  NAND2_X1 U4931 ( .A1(n5124), .A2(n5123), .ZN(n8804) );
  AND2_X1 U4932 ( .A1(n6710), .A2(n8008), .ZN(n7130) );
  INV_X1 U4933 ( .A(n6762), .ZN(n6062) );
  INV_X1 U4934 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n5409) );
  AND2_X1 U4935 ( .A1(n6320), .A2(n6319), .ZN(n8840) );
  INV_X1 U4936 ( .A(n5435), .ZN(n6762) );
  XNOR2_X1 U4937 ( .A(n5393), .B(P1_IR_REG_28__SCAN_IN), .ZN(n6129) );
  INV_X1 U4938 ( .A(n10062), .ZN(n9959) );
  INV_X1 U4939 ( .A(n7876), .ZN(n4989) );
  INV_X2 U4940 ( .A(n7138), .ZN(n7142) );
  NAND2_X2 U4941 ( .A1(n6505), .A2(n6504), .ZN(n9267) );
  INV_X2 U4942 ( .A(n8542), .ZN(n7288) );
  AND2_X1 U4943 ( .A1(n5272), .A2(n4866), .ZN(n8857) );
  INV_X1 U4944 ( .A(n10536), .ZN(n10550) );
  NAND2_X1 U4945 ( .A1(n5814), .A2(n5813), .ZN(n5835) );
  INV_X2 U4946 ( .A(n8810), .ZN(n10466) );
  INV_X2 U4948 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  OR3_X1 U4949 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), .A3(
        P1_IR_REG_21__SCAN_IN), .ZN(n4848) );
  XOR2_X1 U4950 ( .A(n5493), .B(n5492), .Z(n4849) );
  NAND2_X2 U4951 ( .A1(n5815), .A2(n5835), .ZN(n7686) );
  OR2_X2 U4952 ( .A1(n5858), .A2(n5857), .ZN(n5899) );
  OAI22_X2 U4953 ( .A1(n7487), .A2(n5050), .B1(n5052), .B2(n5049), .ZN(n7818)
         );
  NOR3_X2 U4954 ( .A1(n9923), .A2(n9905), .A3(n9908), .ZN(n6159) );
  NAND2_X2 U4955 ( .A1(n5149), .A2(n5147), .ZN(n9923) );
  INV_X1 U4956 ( .A(n9622), .ZN(n8218) );
  NAND2_X4 U4957 ( .A1(n6570), .A2(n6569), .ZN(n9242) );
  NOR2_X2 U4958 ( .A1(n6936), .A2(n5308), .ZN(n5307) );
  OAI22_X2 U4959 ( .A1(n7309), .A2(n7308), .B1(n7060), .B2(n7061), .ZN(n7346)
         );
  NAND2_X1 U4960 ( .A1(n7297), .A2(n7059), .ZN(n7309) );
  INV_X1 U4961 ( .A(n5671), .ZN(n4850) );
  INV_X2 U4962 ( .A(n5671), .ZN(n4851) );
  AND2_X1 U4963 ( .A1(n4996), .A2(n8604), .ZN(n5864) );
  INV_X1 U4964 ( .A(n4849), .ZN(n4852) );
  XNOR2_X2 U4965 ( .A(n9267), .B(n8691), .ZN(n8242) );
  XNOR2_X2 U4966 ( .A(n10408), .B(n9718), .ZN(n10395) );
  NAND2_X2 U4967 ( .A1(n6494), .A2(n6493), .ZN(n8139) );
  OAI21_X2 U4968 ( .B1(n7346), .B2(n5061), .A(n5058), .ZN(n7488) );
  AOI21_X1 U4969 ( .B1(n9753), .B2(n10397), .A(n9752), .ZN(n10001) );
  AND2_X1 U4970 ( .A1(n5146), .A2(n9636), .ZN(n6268) );
  AOI21_X1 U4971 ( .B1(n6803), .B2(n8937), .A(n6802), .ZN(n8963) );
  NAND2_X1 U4972 ( .A1(n9767), .A2(n9770), .ZN(n9766) );
  AOI211_X1 U4973 ( .C1(n10550), .C2(n10549), .A(n10548), .B(n10547), .ZN(
        n10556) );
  AND2_X1 U4974 ( .A1(n5330), .A2(n5329), .ZN(n5066) );
  OAI21_X1 U4975 ( .B1(n8831), .B2(n5313), .A(n5310), .ZN(n5309) );
  NAND2_X1 U4976 ( .A1(n5267), .A2(n4882), .ZN(n9838) );
  NAND2_X1 U4977 ( .A1(n8833), .A2(n8832), .ZN(n8831) );
  AND2_X1 U4978 ( .A1(n5226), .A2(n5224), .ZN(n9389) );
  OAI21_X1 U4979 ( .B1(n5257), .B2(n4961), .A(n4958), .ZN(n5226) );
  NAND2_X1 U4980 ( .A1(n6832), .A2(n6831), .ZN(n8602) );
  AND2_X1 U4981 ( .A1(n5216), .A2(n6734), .ZN(n5215) );
  AND2_X1 U4982 ( .A1(n5233), .A2(n9875), .ZN(n4936) );
  CLKBUF_X1 U4983 ( .A(n9880), .Z(n4935) );
  AND2_X1 U4984 ( .A1(n5344), .A2(n5343), .ZN(n8645) );
  NOR2_X2 U4985 ( .A1(n6838), .A2(n5220), .ZN(n5219) );
  NAND2_X1 U4986 ( .A1(n5046), .A2(n5045), .ZN(n8443) );
  NAND2_X1 U4987 ( .A1(n6010), .A2(n6009), .ZN(n10014) );
  NAND2_X1 U4988 ( .A1(n5965), .A2(n5964), .ZN(n9835) );
  NAND2_X1 U4989 ( .A1(n5948), .A2(n5947), .ZN(n10030) );
  OAI21_X1 U4990 ( .B1(n7921), .B2(n5039), .A(n5037), .ZN(n8207) );
  NAND2_X1 U4991 ( .A1(n6584), .A2(n6583), .ZN(n9232) );
  INV_X1 U4992 ( .A(n8453), .ZN(n9249) );
  NAND2_X1 U4993 ( .A1(n5863), .A2(n5862), .ZN(n10049) );
  NAND2_X1 U4994 ( .A1(n6520), .A2(n6519), .ZN(n9262) );
  NAND2_X1 U4995 ( .A1(n5191), .A2(n5190), .ZN(n8127) );
  AND2_X1 U4996 ( .A1(n8046), .A2(n6459), .ZN(n7985) );
  NAND2_X2 U4997 ( .A1(n9556), .A2(n9554), .ZN(n9671) );
  NAND2_X1 U4998 ( .A1(n6724), .A2(n6902), .ZN(n7987) );
  NAND2_X2 U4999 ( .A1(n9546), .A2(n9537), .ZN(n9658) );
  OR2_X1 U5000 ( .A1(n8184), .A2(n8155), .ZN(n9546) );
  AOI21_X1 U5001 ( .B1(n7764), .B2(n6391), .A(n5382), .ZN(n7688) );
  AND2_X1 U5002 ( .A1(n7476), .A2(n6876), .ZN(n7753) );
  AOI21_X1 U5003 ( .B1(n5211), .B2(n5209), .A(n5208), .ZN(n5207) );
  NAND2_X1 U5004 ( .A1(n5641), .A2(n5640), .ZN(n8155) );
  NAND2_X1 U5005 ( .A1(n5463), .A2(n7460), .ZN(n8588) );
  NAND2_X1 U5006 ( .A1(n5593), .A2(n5592), .ZN(n8162) );
  NAND2_X1 U5007 ( .A1(n5667), .A2(n5666), .ZN(n10490) );
  NOR2_X1 U5008 ( .A1(n7052), .A2(n7049), .ZN(n7258) );
  AND2_X1 U5009 ( .A1(n6394), .A2(n6393), .ZN(n10456) );
  INV_X1 U5010 ( .A(n9712), .ZN(n8276) );
  NAND4_X2 U5011 ( .A1(n5523), .A2(n5522), .A3(n5521), .A4(n5520), .ZN(n9716)
         );
  NAND4_X1 U5012 ( .A1(n6389), .A2(n6388), .A3(n6387), .A4(n6386), .ZN(n8698)
         );
  NAND2_X1 U5013 ( .A1(n6371), .A2(n5189), .ZN(n7665) );
  NOR2_X2 U5014 ( .A1(n6205), .A2(n7365), .ZN(n10396) );
  AND3_X1 U5015 ( .A1(n5375), .A2(n6368), .A3(n6367), .ZN(n7830) );
  NAND2_X1 U5016 ( .A1(n7046), .A2(n5073), .ZN(n7068) );
  AND2_X2 U5017 ( .A1(n5454), .A2(n5453), .ZN(n6083) );
  INV_X1 U5019 ( .A(n6379), .ZN(n6534) );
  INV_X2 U5020 ( .A(n5529), .ZN(n8558) );
  AND2_X1 U5021 ( .A1(n9299), .A2(n8519), .ZN(n6382) );
  NAND2_X2 U5023 ( .A1(n7043), .A2(n7142), .ZN(n5529) );
  NAND2_X1 U5024 ( .A1(n4998), .A2(n4997), .ZN(n10111) );
  INV_X1 U5025 ( .A(n6703), .ZN(n8008) );
  XNOR2_X1 U5026 ( .A(n6707), .B(n6706), .ZN(n6712) );
  NAND2_X2 U5027 ( .A1(n6348), .A2(n7138), .ZN(n6537) );
  OR2_X1 U5028 ( .A1(n9685), .A2(n9622), .ZN(n5443) );
  INV_X1 U5029 ( .A(n8519), .ZN(n6306) );
  NAND2_X2 U5030 ( .A1(n6129), .A2(n9695), .ZN(n7043) );
  XNOR2_X1 U5031 ( .A(n6301), .B(P2_IR_REG_30__SCAN_IN), .ZN(n6307) );
  INV_X1 U5032 ( .A(n6871), .ZN(n8221) );
  NAND2_X1 U5033 ( .A1(n5068), .A2(n5067), .ZN(n6702) );
  XNOR2_X1 U5034 ( .A(n6705), .B(P2_IR_REG_21__SCAN_IN), .ZN(n6871) );
  NAND2_X1 U5035 ( .A1(n9295), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6301) );
  NAND2_X1 U5036 ( .A1(n10104), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5425) );
  NAND2_X1 U5037 ( .A1(n5414), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5410) );
  AND2_X1 U5038 ( .A1(n5471), .A2(n5399), .ZN(n5400) );
  NAND2_X1 U5039 ( .A1(n6314), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6316) );
  NAND2_X1 U5040 ( .A1(n5412), .A2(n5411), .ZN(n5414) );
  XNOR2_X1 U5041 ( .A(n5420), .B(P1_IR_REG_20__SCAN_IN), .ZN(n9622) );
  OR2_X1 U5042 ( .A1(n5412), .A2(n5411), .ZN(n5413) );
  OR2_X1 U5043 ( .A1(n6668), .A2(n9294), .ZN(n6582) );
  AND2_X1 U5044 ( .A1(n6547), .A2(n6568), .ZN(n6668) );
  NAND2_X2 U5045 ( .A1(n7138), .A2(P2_U3152), .ZN(n8219) );
  NOR2_X1 U5046 ( .A1(n6545), .A2(P2_IR_REG_16__SCAN_IN), .ZN(n6547) );
  NOR2_X1 U5047 ( .A1(n5261), .A2(n5035), .ZN(n5260) );
  AND4_X1 U5048 ( .A1(n6299), .A2(n5374), .A3(n6298), .A4(n6297), .ZN(n6300)
         );
  AND2_X1 U5049 ( .A1(n4971), .A2(n4970), .ZN(n5384) );
  AND2_X1 U5050 ( .A1(n5492), .A2(n5126), .ZN(n5524) );
  NOR2_X1 U5051 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n6286) );
  INV_X1 U5052 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n6516) );
  INV_X1 U5053 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5383) );
  NOR2_X1 U5054 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_5__SCAN_IN), .ZN(
        n6290) );
  NOR2_X2 U5055 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .ZN(
        n5127) );
  NOR2_X2 U5056 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n5468) );
  INV_X1 U5057 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5126) );
  INV_X4 U5058 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  INV_X1 U5059 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n9735) );
  INV_X1 U5060 ( .A(P2_RD_REG_SCAN_IN), .ZN(n5327) );
  INV_X1 U5061 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n6678) );
  NOR2_X2 U5062 ( .A1(n8336), .A2(n9262), .ZN(n8411) );
  NAND2_X1 U5063 ( .A1(n9802), .A2(n9801), .ZN(n9800) );
  AOI21_X2 U5064 ( .B1(n9814), .B2(n6243), .A(n5366), .ZN(n9802) );
  NOR2_X2 U5065 ( .A1(n8939), .A2(n7105), .ZN(n8942) );
  AND2_X1 U5066 ( .A1(n7209), .A2(n7734), .ZN(n4856) );
  AND3_X2 U5067 ( .A1(n6356), .A2(n6286), .A3(n6287), .ZN(n6377) );
  NOR2_X4 U5068 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n6356) );
  XNOR2_X2 U5069 ( .A(n6316), .B(n6315), .ZN(n6741) );
  AND2_X1 U5070 ( .A1(n6886), .A2(n6722), .ZN(n5211) );
  OR2_X1 U5071 ( .A1(n6715), .A2(n8221), .ZN(n7046) );
  OR2_X1 U5072 ( .A1(n5996), .A2(n5995), .ZN(n6005) );
  NAND2_X1 U5073 ( .A1(n5743), .A2(SI_12_), .ZN(n5353) );
  INV_X1 U5074 ( .A(n5311), .ZN(n5310) );
  NAND2_X1 U5075 ( .A1(n9506), .A2(n9805), .ZN(n5006) );
  INV_X1 U5076 ( .A(SI_26_), .ZN(n9133) );
  OAI211_X1 U5077 ( .C1(n7686), .C2(n5364), .A(n5362), .B(n5361), .ZN(n7100)
         );
  NAND2_X1 U5078 ( .A1(n8543), .A2(n6833), .ZN(n5364) );
  AND2_X1 U5079 ( .A1(n5363), .A2(n5365), .ZN(n5362) );
  NAND2_X1 U5080 ( .A1(n8818), .A2(n8686), .ZN(n5323) );
  OR2_X1 U5081 ( .A1(n8801), .A2(n8627), .ZN(n6986) );
  OR2_X1 U5082 ( .A1(n8139), .A2(n8211), .ZN(n6858) );
  NAND2_X1 U5083 ( .A1(n8139), .A2(n8211), .ZN(n6860) );
  NAND2_X1 U5084 ( .A1(n6669), .A2(n6296), .ZN(n6676) );
  INV_X1 U5085 ( .A(n6704), .ZN(n6669) );
  NAND2_X1 U5086 ( .A1(n6676), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6707) );
  INV_X1 U5087 ( .A(n9378), .ZN(n5231) );
  NAND2_X1 U5088 ( .A1(n4870), .A2(n4964), .ZN(n4963) );
  INV_X1 U5089 ( .A(n9399), .ZN(n4964) );
  NAND2_X1 U5090 ( .A1(n9881), .A2(n9882), .ZN(n9880) );
  OAI21_X1 U5091 ( .B1(n6228), .B2(n5245), .A(n9929), .ZN(n5244) );
  OR2_X1 U5092 ( .A1(n10080), .A2(n6153), .ZN(n9551) );
  NAND2_X1 U5093 ( .A1(n10080), .A2(n6153), .ZN(n9553) );
  NAND2_X1 U5094 ( .A1(n5384), .A2(n5385), .ZN(n5261) );
  INV_X1 U5095 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5385) );
  NAND2_X1 U5096 ( .A1(n9847), .A2(n9846), .ZN(n5267) );
  NOR2_X1 U5097 ( .A1(n4848), .A2(P1_IR_REG_19__SCAN_IN), .ZN(n5159) );
  NAND2_X1 U5098 ( .A1(n6005), .A2(n6003), .ZN(n6032) );
  AND2_X1 U5099 ( .A1(n6004), .A2(n6002), .ZN(n6003) );
  AOI21_X1 U5100 ( .B1(n5409), .B2(n5418), .A(n5409), .ZN(n4941) );
  INV_X1 U5101 ( .A(n5111), .ZN(n5110) );
  OAI21_X1 U5102 ( .B1(n5372), .B2(n5898), .A(n5112), .ZN(n5111) );
  INV_X1 U5103 ( .A(n5915), .ZN(n5112) );
  NAND3_X1 U5104 ( .A1(n6699), .A2(n10328), .A3(n10327), .ZN(n7039) );
  OR2_X1 U5105 ( .A1(n8522), .A2(n8521), .ZN(n8523) );
  NOR2_X1 U5106 ( .A1(n7071), .A2(n7577), .ZN(n5055) );
  NAND2_X1 U5107 ( .A1(n8008), .A2(n5072), .ZN(n5073) );
  AND2_X1 U5108 ( .A1(n8425), .A2(n5048), .ZN(n5047) );
  OR2_X1 U5109 ( .A1(n8373), .A2(n7102), .ZN(n5048) );
  NAND2_X1 U5110 ( .A1(n6606), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6619) );
  AOI21_X1 U5111 ( .B1(n7005), .B2(n6710), .A(n6871), .ZN(n7006) );
  AND4_X1 U5112 ( .A1(n6474), .A2(n6473), .A3(n6472), .A4(n6471), .ZN(n7922)
         );
  OR2_X1 U5114 ( .A1(n10345), .A2(n10346), .ZN(n5165) );
  AOI22_X1 U5115 ( .A1(n8312), .A2(P2_REG1_REG_14__SCAN_IN), .B1(n8031), .B2(
        n8030), .ZN(n8701) );
  NOR2_X1 U5116 ( .A1(n8998), .A2(n6626), .ZN(n8833) );
  OAI22_X1 U5117 ( .A1(n8857), .A2(n8862), .B1(n8999), .B2(n8871), .ZN(n8846)
         );
  OR2_X1 U5118 ( .A1(n8999), .A2(n8617), .ZN(n6962) );
  OR2_X1 U5119 ( .A1(n8651), .A2(n8687), .ZN(n5371) );
  INV_X1 U5120 ( .A(n6534), .ZN(n6820) );
  NAND2_X1 U5121 ( .A1(n5206), .A2(n5204), .ZN(n6723) );
  AOI21_X1 U5122 ( .B1(n5207), .B2(n5210), .A(n5205), .ZN(n5204) );
  INV_X1 U5123 ( .A(n8673), .ZN(n8916) );
  OR2_X1 U5124 ( .A1(n7587), .A2(n6537), .ZN(n6520) );
  AND2_X1 U5125 ( .A1(n6712), .A2(n8221), .ZN(n10378) );
  AND2_X1 U5126 ( .A1(n7039), .A2(n10331), .ZN(n10155) );
  AND2_X1 U5127 ( .A1(n6067), .A2(n5250), .ZN(n5249) );
  NAND2_X1 U5128 ( .A1(n9344), .A2(n5251), .ZN(n5250) );
  INV_X1 U5129 ( .A(n6030), .ZN(n5251) );
  NAND2_X1 U5130 ( .A1(n4872), .A2(n5017), .ZN(n5016) );
  NOR2_X1 U5131 ( .A1(n9691), .A2(n9692), .ZN(n5017) );
  OAI21_X1 U5132 ( .B1(n9526), .B2(n9527), .A(n5019), .ZN(n5018) );
  NAND2_X1 U5133 ( .A1(n5020), .A2(n9477), .ZN(n5019) );
  OAI21_X1 U5134 ( .B1(n9766), .B2(n5145), .A(n5141), .ZN(n6191) );
  AOI21_X1 U5135 ( .B1(n5144), .B2(n5143), .A(n5142), .ZN(n5141) );
  INV_X1 U5136 ( .A(n9616), .ZN(n5142) );
  AND2_X1 U5137 ( .A1(n9498), .A2(n9499), .ZN(n9850) );
  AOI21_X1 U5138 ( .B1(n9869), .B2(n5132), .A(n9497), .ZN(n5131) );
  INV_X1 U5139 ( .A(n9572), .ZN(n5132) );
  AND2_X1 U5140 ( .A1(n9558), .A2(n9559), .ZN(n5153) );
  INV_X1 U5141 ( .A(n9929), .ZN(n5151) );
  AOI21_X1 U5142 ( .B1(n8273), .B2(n9470), .A(n6218), .ZN(n8323) );
  INV_X2 U5143 ( .A(n5528), .ZN(n6072) );
  NAND2_X1 U5144 ( .A1(n5442), .A2(n9696), .ZN(n10401) );
  NAND2_X1 U5145 ( .A1(n6192), .A2(n9442), .ZN(n10397) );
  AND2_X1 U5146 ( .A1(n5718), .A2(n5716), .ZN(n5332) );
  INV_X1 U5147 ( .A(n5719), .ZN(n5718) );
  NAND2_X1 U5148 ( .A1(n7395), .A2(n7394), .ZN(n10357) );
  XNOR2_X1 U5149 ( .A(n5439), .B(P1_IR_REG_22__SCAN_IN), .ZN(n9441) );
  NAND2_X1 U5150 ( .A1(n5438), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5439) );
  XNOR2_X1 U5151 ( .A(n6251), .B(n9650), .ZN(n9996) );
  NAND2_X1 U5152 ( .A1(n6265), .A2(n4877), .ZN(n6251) );
  NOR2_X1 U5153 ( .A1(n6915), .A2(n8128), .ZN(n4934) );
  AOI21_X1 U5154 ( .B1(n9488), .B2(n4910), .A(n5025), .ZN(n5024) );
  NAND2_X1 U5155 ( .A1(n5238), .A2(n5022), .ZN(n5021) );
  NAND2_X1 U5156 ( .A1(n4898), .A2(n5023), .ZN(n5022) );
  INV_X1 U5157 ( .A(n9491), .ZN(n5023) );
  AND2_X1 U5158 ( .A1(n5004), .A2(n4904), .ZN(n5003) );
  OR2_X1 U5159 ( .A1(n5006), .A2(n4903), .ZN(n5004) );
  NAND2_X1 U5160 ( .A1(n7719), .A2(n5285), .ZN(n5284) );
  INV_X1 U5161 ( .A(n5100), .ZN(n5099) );
  OAI21_X1 U5162 ( .B1(n5102), .B2(n5101), .A(n6068), .ZN(n5100) );
  INV_X1 U5163 ( .A(n4914), .ZN(n5101) );
  INV_X1 U5164 ( .A(SI_20_), .ZN(n9020) );
  AND2_X1 U5165 ( .A1(n5334), .A2(n5082), .ZN(n5081) );
  NOR2_X1 U5166 ( .A1(n5660), .A2(n5335), .ZN(n5334) );
  NAND2_X1 U5167 ( .A1(n5587), .A2(n5083), .ZN(n5082) );
  INV_X1 U5168 ( .A(n5634), .ZN(n5335) );
  INV_X1 U5169 ( .A(n5587), .ZN(n5084) );
  INV_X1 U5170 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n5075) );
  NOR2_X1 U5171 ( .A1(n6599), .A2(n9084), .ZN(n6321) );
  AND2_X1 U5172 ( .A1(n6837), .A2(n6999), .ZN(n7022) );
  NAND2_X1 U5173 ( .A1(n8768), .A2(n8684), .ZN(n6837) );
  OR2_X1 U5174 ( .A1(n6395), .A2(n7667), .ZN(n6366) );
  NAND2_X1 U5175 ( .A1(n5118), .A2(n6757), .ZN(n5117) );
  INV_X1 U5176 ( .A(n8862), .ZN(n5217) );
  NAND2_X1 U5177 ( .A1(n5185), .A2(n5187), .ZN(n5183) );
  AND2_X1 U5178 ( .A1(n6953), .A2(n6955), .ZN(n6847) );
  AND2_X1 U5179 ( .A1(n6952), .A2(n6949), .ZN(n6944) );
  INV_X1 U5180 ( .A(n6557), .ZN(n5308) );
  AND2_X1 U5181 ( .A1(n6940), .A2(n6939), .ZN(n6936) );
  OR2_X1 U5182 ( .A1(n7105), .A2(n7104), .ZN(n6933) );
  AND2_X1 U5183 ( .A1(n6922), .A2(n6726), .ZN(n5214) );
  INV_X1 U5184 ( .A(n5202), .ZN(n5201) );
  OAI21_X1 U5185 ( .B1(n7787), .B2(n5203), .A(n7805), .ZN(n5202) );
  INV_X1 U5186 ( .A(n6896), .ZN(n5203) );
  NAND2_X1 U5187 ( .A1(n7296), .A2(n7310), .ZN(n6877) );
  NAND2_X1 U5188 ( .A1(n7830), .A2(n7665), .ZN(n6876) );
  NOR2_X1 U5189 ( .A1(n8801), .A2(n8982), .ZN(n5123) );
  NAND2_X1 U5190 ( .A1(n5279), .A2(n5284), .ZN(n5278) );
  NAND2_X1 U5191 ( .A1(n7785), .A2(n6417), .ZN(n5279) );
  OAI21_X1 U5192 ( .B1(n5283), .B2(n5276), .A(n5275), .ZN(n7804) );
  INV_X1 U5193 ( .A(n5278), .ZN(n5276) );
  AOI21_X1 U5194 ( .B1(n5278), .B2(n5281), .A(n7805), .ZN(n5275) );
  INV_X1 U5195 ( .A(n4955), .ZN(n4950) );
  OR2_X1 U5196 ( .A1(n8362), .A2(n4954), .ZN(n4953) );
  NAND2_X1 U5197 ( .A1(n5758), .A2(n4957), .ZN(n4954) );
  NAND2_X1 U5198 ( .A1(n8249), .A2(n5738), .ZN(n4947) );
  NOR2_X1 U5199 ( .A1(n8362), .A2(n4956), .ZN(n4955) );
  INV_X1 U5200 ( .A(n4957), .ZN(n4956) );
  OR2_X1 U5201 ( .A1(n9994), .A2(n7368), .ZN(n9519) );
  OR2_X1 U5202 ( .A1(n9998), .A2(n10003), .ZN(n4984) );
  OR2_X1 U5203 ( .A1(n9820), .A2(n9831), .ZN(n9633) );
  OR2_X1 U5204 ( .A1(n9896), .A2(n9907), .ZN(n6234) );
  NAND2_X1 U5205 ( .A1(n9959), .A2(n4994), .ZN(n4993) );
  OR2_X1 U5206 ( .A1(n10068), .A2(n9707), .ZN(n6223) );
  NAND2_X1 U5207 ( .A1(n9671), .A2(n8468), .ZN(n6222) );
  NOR2_X1 U5208 ( .A1(n10068), .A2(n6157), .ZN(n4994) );
  NAND2_X1 U5209 ( .A1(n4896), .A2(n6216), .ZN(n5254) );
  AND2_X1 U5210 ( .A1(n9658), .A2(n6215), .ZN(n5255) );
  AND2_X1 U5211 ( .A1(n9457), .A2(n9454), .ZN(n9452) );
  NAND2_X1 U5212 ( .A1(n4989), .A2(n7936), .ZN(n4988) );
  NAND2_X1 U5213 ( .A1(n6147), .A2(n5008), .ZN(n9625) );
  INV_X1 U5214 ( .A(n9596), .ZN(n5009) );
  NAND2_X1 U5215 ( .A1(n9592), .A2(n10408), .ZN(n4995) );
  NAND2_X1 U5216 ( .A1(n6182), .A2(n6181), .ZN(n6826) );
  INV_X1 U5217 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5427) );
  INV_X1 U5218 ( .A(n5937), .ZN(n5108) );
  AOI21_X1 U5219 ( .B1(n5110), .B2(n5372), .A(n4912), .ZN(n5109) );
  OR2_X1 U5220 ( .A1(n5836), .A2(P1_IR_REG_15__SCAN_IN), .ZN(n5860) );
  INV_X1 U5221 ( .A(SI_15_), .ZN(n9121) );
  NAND2_X1 U5222 ( .A1(n5759), .A2(n5354), .ZN(n5352) );
  INV_X1 U5223 ( .A(n5781), .ZN(n5354) );
  INV_X1 U5224 ( .A(SI_10_), .ZN(n9155) );
  AND2_X1 U5225 ( .A1(n5499), .A2(n5536), .ZN(n5337) );
  INV_X1 U5226 ( .A(n5530), .ZN(n5340) );
  AND2_X1 U5227 ( .A1(n8120), .A2(n5043), .ZN(n5040) );
  NAND2_X1 U5228 ( .A1(n8528), .A2(n5331), .ZN(n5330) );
  OR2_X1 U5229 ( .A1(n8372), .A2(n7102), .ZN(n5044) );
  XNOR2_X1 U5230 ( .A(n8528), .B(n8529), .ZN(n8634) );
  OAI21_X1 U5231 ( .B1(n5055), .B2(n5054), .A(n7717), .ZN(n5053) );
  NAND2_X1 U5232 ( .A1(n7076), .A2(n7077), .ZN(n5056) );
  NAND2_X1 U5233 ( .A1(n8486), .A2(n5348), .ZN(n5341) );
  NAND2_X1 U5234 ( .A1(n8439), .A2(n8440), .ZN(n5348) );
  AND2_X1 U5235 ( .A1(n7332), .A2(n7288), .ZN(n7056) );
  OR2_X1 U5236 ( .A1(n7112), .A2(n7111), .ZN(n5350) );
  NAND2_X1 U5237 ( .A1(n8372), .A2(n8373), .ZN(n8371) );
  AND4_X1 U5238 ( .A1(n6416), .A2(n6415), .A3(n6414), .A4(n6413), .ZN(n7579)
         );
  AND2_X1 U5239 ( .A1(n5165), .A2(n5164), .ZN(n10360) );
  NOR2_X1 U5240 ( .A1(n10360), .A2(n10359), .ZN(n10358) );
  AOI21_X1 U5241 ( .B1(P2_REG1_REG_8__SCAN_IN), .B2(n7520), .A(n7568), .ZN(
        n7522) );
  AND2_X1 U5242 ( .A1(n7014), .A2(n7010), .ZN(n6994) );
  AOI21_X1 U5243 ( .B1(n5316), .B2(n5315), .A(n4894), .ZN(n5314) );
  INV_X1 U5244 ( .A(n5321), .ZN(n5315) );
  INV_X1 U5245 ( .A(n8795), .ZN(n5318) );
  AND2_X1 U5246 ( .A1(n5323), .A2(n5322), .ZN(n5321) );
  NAND2_X1 U5247 ( .A1(n8813), .A2(n5323), .ZN(n5320) );
  NAND2_X1 U5248 ( .A1(n8840), .A2(n8629), .ZN(n5322) );
  NOR2_X1 U5249 ( .A1(n8882), .A2(n5274), .ZN(n5273) );
  INV_X1 U5250 ( .A(n5371), .ZN(n5274) );
  AND2_X1 U5251 ( .A1(n6960), .A2(n6956), .ZN(n8882) );
  INV_X1 U5252 ( .A(n6949), .ZN(n5187) );
  INV_X1 U5253 ( .A(n5186), .ZN(n5185) );
  OAI21_X1 U5254 ( .B1(n6731), .B2(n5187), .A(n6952), .ZN(n5186) );
  INV_X1 U5255 ( .A(n6847), .ZN(n8896) );
  INV_X1 U5256 ( .A(n6944), .ZN(n8903) );
  NAND2_X1 U5257 ( .A1(n6929), .A2(n6928), .ZN(n8419) );
  NAND2_X1 U5258 ( .A1(n6727), .A2(n5214), .ZN(n8344) );
  AOI21_X1 U5259 ( .B1(n8132), .B2(n5293), .A(n4862), .ZN(n5292) );
  OR2_X1 U5260 ( .A1(n7330), .A2(n6537), .ZN(n6494) );
  AOI21_X1 U5261 ( .B1(n5193), .B2(n5196), .A(n6857), .ZN(n5190) );
  INV_X1 U5262 ( .A(n6909), .ZN(n5196) );
  AOI21_X1 U5263 ( .B1(n5297), .B2(n5300), .A(n4874), .ZN(n5295) );
  INV_X1 U5264 ( .A(n6475), .ZN(n5300) );
  AND2_X1 U5265 ( .A1(n6912), .A2(n6910), .ZN(n8091) );
  NAND2_X1 U5266 ( .A1(n7985), .A2(n7988), .ZN(n7984) );
  INV_X1 U5267 ( .A(n6885), .ZN(n5208) );
  INV_X1 U5268 ( .A(n7767), .ZN(n5209) );
  INV_X1 U5269 ( .A(n5211), .ZN(n5210) );
  AND2_X1 U5270 ( .A1(n6886), .A2(n6885), .ZN(n7689) );
  NAND2_X1 U5271 ( .A1(n7753), .A2(n7767), .ZN(n7752) );
  OR2_X1 U5272 ( .A1(n7371), .A2(n6748), .ZN(n8673) );
  INV_X1 U5273 ( .A(n8768), .ZN(n8957) );
  NAND2_X1 U5274 ( .A1(n6595), .A2(n6594), .ZN(n9011) );
  NAND2_X1 U5275 ( .A1(n6710), .A2(n10378), .ZN(n10545) );
  NAND2_X1 U5276 ( .A1(n6677), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6708) );
  NAND2_X1 U5277 ( .A1(n6300), .A2(n6547), .ZN(n6674) );
  NOR2_X1 U5278 ( .A1(P2_IR_REG_27__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), .ZN(
        n5324) );
  NOR2_X1 U5279 ( .A1(n6676), .A2(n6671), .ZN(n6681) );
  NAND2_X1 U5280 ( .A1(n6704), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6705) );
  AOI21_X1 U5281 ( .B1(n5070), .B2(n9294), .A(n9294), .ZN(n5067) );
  XNOR2_X1 U5282 ( .A(n6701), .B(P2_IR_REG_19__SCAN_IN), .ZN(n6703) );
  NAND2_X1 U5283 ( .A1(n4900), .A2(n5231), .ZN(n5228) );
  AOI21_X1 U5284 ( .B1(n4899), .B2(n4963), .A(n4959), .ZN(n4958) );
  AND2_X1 U5285 ( .A1(n4960), .A2(n9400), .ZN(n4959) );
  INV_X1 U5286 ( .A(n5256), .ZN(n4960) );
  NOR2_X1 U5287 ( .A1(n4963), .A2(n9400), .ZN(n4961) );
  AND2_X1 U5288 ( .A1(n9410), .A2(n6030), .ZN(n4944) );
  AOI21_X1 U5289 ( .B1(n4941), .B2(P1_IR_REG_20__SCAN_IN), .A(
        P1_IR_REG_21__SCAN_IN), .ZN(n4939) );
  INV_X1 U5290 ( .A(n4941), .ZN(n4940) );
  NOR2_X1 U5291 ( .A1(n8604), .A2(n10111), .ZN(n5548) );
  NAND2_X1 U5292 ( .A1(n8560), .A2(n8559), .ZN(n9742) );
  OR2_X1 U5293 ( .A1(n9789), .A2(n4984), .ZN(n9761) );
  NOR2_X1 U5294 ( .A1(n9789), .A2(n4981), .ZN(n6273) );
  AND2_X1 U5295 ( .A1(n9513), .A2(n9616), .ZN(n9678) );
  OR2_X1 U5296 ( .A1(n6263), .A2(n9678), .ZN(n6265) );
  AND2_X1 U5297 ( .A1(n6187), .A2(n6136), .ZN(n8594) );
  NAND2_X1 U5298 ( .A1(n6249), .A2(n6248), .ZN(n9755) );
  INV_X1 U5299 ( .A(n9754), .ZN(n9748) );
  AND2_X1 U5300 ( .A1(n9610), .A2(n9747), .ZN(n9770) );
  INV_X1 U5301 ( .A(n9704), .ZN(n9768) );
  NAND2_X1 U5302 ( .A1(n9800), .A2(n4881), .ZN(n9793) );
  INV_X1 U5303 ( .A(n9796), .ZN(n6245) );
  AND2_X1 U5304 ( .A1(n9609), .A2(n9607), .ZN(n9796) );
  AND2_X1 U5305 ( .A1(n9579), .A2(n9575), .ZN(n9841) );
  NAND2_X1 U5306 ( .A1(n5130), .A2(n5128), .ZN(n9848) );
  AND2_X1 U5307 ( .A1(n9850), .A2(n5129), .ZN(n5128) );
  NAND2_X1 U5308 ( .A1(n5131), .A2(n5133), .ZN(n5129) );
  NAND2_X1 U5309 ( .A1(n6239), .A2(n6238), .ZN(n9847) );
  INV_X1 U5310 ( .A(n9850), .ZN(n9846) );
  NAND2_X1 U5311 ( .A1(n10039), .A2(n9405), .ZN(n9572) );
  AND2_X1 U5312 ( .A1(n9573), .A2(n9572), .ZN(n9882) );
  INV_X1 U5313 ( .A(n6234), .ZN(n5239) );
  NAND2_X1 U5314 ( .A1(n6233), .A2(n6232), .ZN(n9890) );
  NOR2_X1 U5315 ( .A1(n10049), .A2(n9936), .ZN(n9914) );
  NAND2_X1 U5316 ( .A1(n5240), .A2(n5243), .ZN(n9928) );
  INV_X1 U5317 ( .A(n5244), .ZN(n5243) );
  NOR2_X1 U5318 ( .A1(n5242), .A2(n5245), .ZN(n5241) );
  OAI21_X1 U5319 ( .B1(n5150), .B2(n5148), .A(n5151), .ZN(n5147) );
  AND2_X1 U5320 ( .A1(n5153), .A2(n9973), .ZN(n5150) );
  NAND2_X1 U5321 ( .A1(n8381), .A2(n6221), .ZN(n9943) );
  NAND2_X1 U5322 ( .A1(n9943), .A2(n6228), .ZN(n9944) );
  NOR2_X1 U5323 ( .A1(n9974), .A2(n9973), .ZN(n9971) );
  AND2_X1 U5324 ( .A1(n8328), .A2(n10521), .ZN(n8388) );
  NAND2_X1 U5325 ( .A1(n8112), .A2(n5255), .ZN(n8144) );
  OR2_X1 U5326 ( .A1(n8152), .A2(n8155), .ZN(n8190) );
  NOR2_X1 U5327 ( .A1(n9452), .A2(n5266), .ZN(n5265) );
  INV_X1 U5328 ( .A(n6214), .ZN(n5266) );
  INV_X1 U5329 ( .A(n9452), .ZN(n9656) );
  AND2_X1 U5330 ( .A1(n7871), .A2(n6211), .ZN(n7938) );
  NAND2_X1 U5331 ( .A1(n7938), .A2(n6213), .ZN(n7937) );
  NAND2_X1 U5332 ( .A1(n7621), .A2(n6196), .ZN(n9977) );
  NOR2_X1 U5333 ( .A1(n10408), .A2(n10385), .ZN(n10388) );
  OR2_X1 U5334 ( .A1(n6117), .A2(n9693), .ZN(n9696) );
  INV_X1 U5335 ( .A(n9975), .ZN(n10391) );
  OR2_X1 U5336 ( .A1(n7330), .A2(n5529), .ZN(n5747) );
  NAND2_X1 U5337 ( .A1(n5694), .A2(n5693), .ZN(n10501) );
  AND2_X1 U5338 ( .A1(n6097), .A2(n6096), .ZN(n10121) );
  AND2_X1 U5339 ( .A1(n8397), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7037) );
  NOR2_X1 U5340 ( .A1(n4889), .A2(n5270), .ZN(n5269) );
  XNOR2_X1 U5341 ( .A(n6819), .B(n6818), .ZN(n9293) );
  AND2_X1 U5342 ( .A1(n6815), .A2(n6827), .ZN(n6819) );
  NAND2_X1 U5343 ( .A1(n5098), .A2(n4914), .ZN(n6069) );
  NAND2_X1 U5344 ( .A1(n6032), .A2(n5102), .ZN(n5098) );
  NAND2_X1 U5345 ( .A1(n6032), .A2(n6031), .ZN(n6047) );
  INV_X1 U5346 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n6115) );
  XNOR2_X1 U5347 ( .A(n5981), .B(n5992), .ZN(n8396) );
  OR2_X1 U5348 ( .A1(n5996), .A2(n5994), .ZN(n5980) );
  OR2_X1 U5349 ( .A1(n5790), .A2(P1_IR_REG_14__SCAN_IN), .ZN(n5836) );
  NAND2_X1 U5350 ( .A1(n5353), .A2(n5089), .ZN(n5088) );
  INV_X1 U5351 ( .A(n5352), .ZN(n5089) );
  NOR2_X1 U5352 ( .A1(n5742), .A2(n5105), .ZN(n5104) );
  INV_X1 U5353 ( .A(n5739), .ZN(n5105) );
  INV_X1 U5354 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n4971) );
  NAND2_X1 U5355 ( .A1(n5400), .A2(n5401), .ZN(n5472) );
  AND2_X1 U5356 ( .A1(n4876), .A2(n4861), .ZN(n5258) );
  NAND2_X1 U5357 ( .A1(n6654), .A2(n6653), .ZN(n8965) );
  AND2_X1 U5358 ( .A1(n6614), .A2(n6613), .ZN(n8617) );
  AOI21_X1 U5359 ( .B1(n5047), .B2(n7102), .A(n7108), .ZN(n5045) );
  AND2_X1 U5360 ( .A1(n6625), .A2(n6624), .ZN(n8661) );
  AND2_X1 U5361 ( .A1(n6591), .A2(n6590), .ZN(n8492) );
  AND2_X1 U5362 ( .A1(n7256), .A2(n7129), .ZN(n8641) );
  NAND2_X1 U5363 ( .A1(n7133), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8678) );
  INV_X1 U5364 ( .A(n8669), .ZN(n8657) );
  OR3_X1 U5365 ( .A1(n6543), .A2(n6542), .A3(n6541), .ZN(n8308) );
  INV_X1 U5366 ( .A(n7579), .ZN(n7789) );
  AND2_X1 U5367 ( .A1(n5163), .A2(n5162), .ZN(n7599) );
  NAND2_X1 U5368 ( .A1(n7602), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n5162) );
  AND2_X1 U5369 ( .A1(n6531), .A2(n6518), .ZN(n8312) );
  AND2_X1 U5370 ( .A1(n7395), .A2(n6741), .ZN(n10364) );
  AOI21_X1 U5371 ( .B1(n10352), .B2(P2_ADDR_REG_19__SCAN_IN), .A(n8764), .ZN(
        n5177) );
  INV_X1 U5372 ( .A(n5181), .ZN(n5180) );
  AOI21_X1 U5373 ( .B1(n8961), .B2(n8926), .A(n6807), .ZN(n6808) );
  OR2_X1 U5374 ( .A1(n8968), .A2(n10466), .ZN(n6760) );
  NAND2_X1 U5375 ( .A1(n8810), .A2(n10452), .ZN(n8930) );
  NAND2_X1 U5376 ( .A1(n8810), .A2(n10463), .ZN(n8952) );
  INV_X1 U5377 ( .A(n8777), .ZN(n8926) );
  NAND2_X1 U5378 ( .A1(n5248), .A2(n5246), .ZN(n6786) );
  AND2_X1 U5379 ( .A1(n6091), .A2(n5247), .ZN(n5246) );
  AND2_X1 U5380 ( .A1(n6092), .A2(n6093), .ZN(n6091) );
  NAND2_X1 U5381 ( .A1(n5725), .A2(n5724), .ZN(n9446) );
  OR2_X1 U5382 ( .A1(n7686), .A2(n5529), .ZN(n5819) );
  OAI21_X1 U5383 ( .B1(n5018), .B2(n4857), .A(n5015), .ZN(n5014) );
  AOI21_X1 U5384 ( .B1(n5018), .B2(n9528), .A(n5016), .ZN(n5015) );
  INV_X1 U5385 ( .A(n9701), .ZN(n5013) );
  AOI21_X1 U5386 ( .B1(n9995), .B2(n10368), .A(n6259), .ZN(n6260) );
  NAND2_X1 U5387 ( .A1(n6200), .A2(n4917), .ZN(n5139) );
  OR2_X1 U5388 ( .A1(n10419), .A2(n10406), .ZN(n9969) );
  OR2_X1 U5389 ( .A1(n10419), .A2(n7735), .ZN(n9779) );
  NAND2_X1 U5390 ( .A1(n6203), .A2(n6278), .ZN(n10376) );
  NAND2_X1 U5391 ( .A1(n9995), .A2(n10386), .ZN(n4976) );
  OR2_X1 U5392 ( .A1(n9996), .A2(n10436), .ZN(n4977) );
  AOI21_X1 U5393 ( .B1(n5007), .B2(n9653), .A(n9453), .ZN(n9460) );
  XNOR2_X1 U5394 ( .A(n9451), .B(n9477), .ZN(n5007) );
  NAND2_X1 U5395 ( .A1(n5034), .A2(n6151), .ZN(n5033) );
  OAI21_X1 U5396 ( .B1(n9467), .B2(n9658), .A(n9466), .ZN(n5034) );
  NOR2_X1 U5397 ( .A1(n9470), .A2(n9471), .ZN(n5032) );
  NAND2_X1 U5398 ( .A1(n9476), .A2(n9475), .ZN(n5028) );
  AND2_X1 U5399 ( .A1(n9473), .A2(n9474), .ZN(n5030) );
  AOI21_X1 U5400 ( .B1(n5031), .B2(n5029), .A(n5027), .ZN(n9482) );
  NOR2_X1 U5401 ( .A1(n5030), .A2(n9472), .ZN(n5029) );
  NAND2_X1 U5402 ( .A1(n6154), .A2(n5028), .ZN(n5027) );
  NAND2_X1 U5403 ( .A1(n5033), .A2(n5032), .ZN(n5031) );
  OR2_X1 U5404 ( .A1(n9489), .A2(n9556), .ZN(n5026) );
  AND2_X1 U5405 ( .A1(n5002), .A2(n4905), .ZN(n5001) );
  NAND2_X1 U5406 ( .A1(n5003), .A2(n5005), .ZN(n5002) );
  OAI211_X1 U5407 ( .C1(n5024), .C2(n5021), .A(n9492), .B(n9882), .ZN(n9494)
         );
  INV_X1 U5408 ( .A(n5582), .ZN(n5083) );
  OR2_X1 U5409 ( .A1(n6536), .A2(n8537), .ZN(n5365) );
  NAND2_X1 U5410 ( .A1(n4873), .A2(n6537), .ZN(n5363) );
  NOR2_X1 U5411 ( .A1(n7017), .A2(n4932), .ZN(n4931) );
  INV_X1 U5412 ( .A(n6999), .ZN(n4932) );
  NAND2_X1 U5413 ( .A1(n7472), .A2(n7054), .ZN(n6720) );
  INV_X1 U5414 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n6700) );
  INV_X1 U5415 ( .A(n5229), .ZN(n5227) );
  INV_X1 U5416 ( .A(n5370), .ZN(n5010) );
  NOR2_X1 U5417 ( .A1(n5095), .A2(n5092), .ZN(n5091) );
  INV_X1 U5418 ( .A(n6168), .ZN(n5092) );
  INV_X1 U5419 ( .A(n6181), .ZN(n5095) );
  NAND2_X1 U5420 ( .A1(n6181), .A2(n5094), .ZN(n5093) );
  INV_X1 U5421 ( .A(n6175), .ZN(n5094) );
  INV_X1 U5422 ( .A(SI_23_), .ZN(n5990) );
  INV_X1 U5423 ( .A(SI_9_), .ZN(n9161) );
  OAI21_X1 U5424 ( .B1(n5314), .B2(n5312), .A(n4864), .ZN(n5311) );
  OR2_X1 U5425 ( .A1(n8993), .A2(n8661), .ZN(n6965) );
  INV_X1 U5426 ( .A(n6962), .ZN(n5220) );
  OR2_X1 U5427 ( .A1(n9232), .A2(n8492), .ZN(n6952) );
  AND2_X1 U5428 ( .A1(n6562), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n6571) );
  NOR2_X1 U5429 ( .A1(n6523), .A2(n6522), .ZN(n6521) );
  AND2_X1 U5430 ( .A1(n6912), .A2(n5194), .ZN(n5193) );
  NAND2_X1 U5431 ( .A1(n5195), .A2(n6909), .ZN(n5194) );
  INV_X1 U5432 ( .A(n6911), .ZN(n5195) );
  AND2_X1 U5433 ( .A1(n8089), .A2(n5298), .ZN(n5297) );
  NAND2_X1 U5434 ( .A1(n5299), .A2(n6475), .ZN(n5298) );
  INV_X1 U5435 ( .A(n7988), .ZN(n5299) );
  NOR2_X1 U5436 ( .A1(n7809), .A2(n7849), .ZN(n5122) );
  NOR2_X1 U5437 ( .A1(n7768), .A2(n8698), .ZN(n6881) );
  NAND2_X1 U5438 ( .A1(n6717), .A2(n7286), .ZN(n6719) );
  NOR2_X1 U5439 ( .A1(n7693), .A2(n7681), .ZN(n7794) );
  OAI21_X1 U5440 ( .B1(n6698), .B2(n6697), .A(n6696), .ZN(n7120) );
  OAI21_X1 U5441 ( .B1(P2_D_REG_1__SCAN_IN), .B2(n10154), .A(n10153), .ZN(
        n7223) );
  INV_X1 U5442 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n6670) );
  INV_X1 U5443 ( .A(n5071), .ZN(n5070) );
  OAI21_X1 U5444 ( .B1(n6581), .B2(n9294), .A(n6700), .ZN(n5071) );
  INV_X1 U5445 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n6581) );
  INV_X1 U5446 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n6288) );
  INV_X1 U5447 ( .A(n4870), .ZN(n4965) );
  INV_X1 U5448 ( .A(n9649), .ZN(n5020) );
  INV_X1 U5449 ( .A(n9647), .ZN(n9684) );
  NAND2_X1 U5450 ( .A1(n4983), .A2(n4982), .ZN(n4981) );
  INV_X1 U5451 ( .A(n4984), .ZN(n4983) );
  NOR2_X1 U5452 ( .A1(n5239), .A2(n5235), .ZN(n5234) );
  INV_X1 U5453 ( .A(n6232), .ZN(n5235) );
  NAND2_X1 U5454 ( .A1(n5238), .A2(n6234), .ZN(n5237) );
  INV_X1 U5455 ( .A(n6221), .ZN(n5242) );
  INV_X1 U5456 ( .A(n6229), .ZN(n5245) );
  NAND2_X1 U5457 ( .A1(n7739), .A2(n9717), .ZN(n9598) );
  AND2_X1 U5458 ( .A1(n8218), .A2(n9856), .ZN(n6124) );
  NAND2_X1 U5459 ( .A1(n6115), .A2(n5271), .ZN(n5270) );
  NAND2_X1 U5460 ( .A1(n6176), .A2(n6175), .ZN(n6182) );
  NAND2_X1 U5461 ( .A1(n5391), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5394) );
  AOI21_X1 U5462 ( .B1(n5099), .B2(n5101), .A(n4919), .ZN(n5097) );
  NOR2_X1 U5463 ( .A1(n6046), .A2(n5103), .ZN(n5102) );
  INV_X1 U5464 ( .A(n6031), .ZN(n5103) );
  AND3_X1 U5465 ( .A1(n5260), .A2(n5636), .A3(n5158), .ZN(n5422) );
  AND2_X1 U5466 ( .A1(n5159), .A2(n5268), .ZN(n5158) );
  INV_X1 U5467 ( .A(n5270), .ZN(n5268) );
  AOI21_X1 U5468 ( .B1(n5081), .B2(n5084), .A(n4895), .ZN(n5079) );
  INV_X1 U5469 ( .A(SI_5_), .ZN(n9165) );
  INV_X1 U5470 ( .A(P1_RD_REG_SCAN_IN), .ZN(n5076) );
  NAND2_X1 U5471 ( .A1(n6571), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n6597) );
  OR2_X1 U5472 ( .A1(n6597), .A2(n6596), .ZN(n6599) );
  NAND2_X1 U5473 ( .A1(n7346), .A2(n7343), .ZN(n5064) );
  AOI21_X1 U5474 ( .B1(n8120), .B2(n5038), .A(n7090), .ZN(n5037) );
  INV_X1 U5475 ( .A(n5040), .ZN(n5039) );
  NOR2_X1 U5476 ( .A1(n7920), .A2(n5042), .ZN(n5038) );
  NAND2_X1 U5477 ( .A1(n6871), .A2(n5072), .ZN(n7371) );
  INV_X1 U5478 ( .A(n7344), .ZN(n5063) );
  OR2_X1 U5479 ( .A1(n8531), .A2(n8530), .ZN(n8532) );
  NAND2_X1 U5480 ( .A1(n5066), .A2(n8636), .ZN(n8623) );
  INV_X1 U5481 ( .A(n8626), .ZN(n5329) );
  AOI21_X1 U5482 ( .B1(n8816), .B2(n6747), .A(n6634), .ZN(n8686) );
  INV_X1 U5483 ( .A(n6384), .ZN(n6747) );
  AND4_X1 U5484 ( .A1(n6456), .A2(n6455), .A3(n6454), .A4(n6453), .ZN(n7902)
         );
  AND2_X1 U5485 ( .A1(n6366), .A2(n6365), .ZN(n6367) );
  OR2_X1 U5486 ( .A1(n6384), .A2(n7294), .ZN(n6345) );
  AOI21_X1 U5487 ( .B1(n7441), .B2(P2_REG1_REG_3__SCAN_IN), .A(n7429), .ZN(
        n7401) );
  OR2_X1 U5488 ( .A1(n7402), .A2(n7401), .ZN(n7404) );
  OR2_X1 U5489 ( .A1(n7517), .A2(n7516), .ZN(n5163) );
  AOI21_X1 U5490 ( .B1(n7892), .B2(P2_REG1_REG_11__SCAN_IN), .A(n7883), .ZN(
        n7886) );
  NOR2_X1 U5491 ( .A1(n8036), .A2(n5168), .ZN(n8040) );
  AND2_X1 U5492 ( .A1(n8037), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n5168) );
  NAND2_X1 U5493 ( .A1(n8040), .A2(n8039), .ZN(n8311) );
  AOI21_X1 U5494 ( .B1(P2_REG1_REG_17__SCAN_IN), .B2(n8738), .A(n8737), .ZN(
        n8750) );
  NAND2_X1 U5495 ( .A1(n5171), .A2(n5170), .ZN(n8759) );
  INV_X1 U5496 ( .A(n8748), .ZN(n5170) );
  NAND2_X1 U5497 ( .A1(n8746), .A2(n5172), .ZN(n5171) );
  INV_X1 U5498 ( .A(n8747), .ZN(n5172) );
  INV_X1 U5499 ( .A(n5117), .ZN(n5115) );
  NAND2_X1 U5500 ( .A1(n8786), .A2(n5116), .ZN(n8771) );
  NOR2_X1 U5501 ( .A1(n10549), .A2(n5117), .ZN(n5116) );
  AND2_X1 U5502 ( .A1(n6665), .A2(n6664), .ZN(n8609) );
  OR2_X1 U5503 ( .A1(n8965), .A2(n8609), .ZN(n7011) );
  AND2_X1 U5504 ( .A1(n6657), .A2(n6656), .ZN(n6805) );
  NAND2_X1 U5505 ( .A1(n6636), .A2(n6635), .ZN(n8801) );
  AND2_X2 U5506 ( .A1(n6965), .A2(n8826), .ZN(n8845) );
  NAND2_X1 U5507 ( .A1(n8863), .A2(n8862), .ZN(n5221) );
  NAND2_X1 U5508 ( .A1(n5219), .A2(n5221), .ZN(n5367) );
  AND2_X1 U5509 ( .A1(n6962), .A2(n6964), .ZN(n8862) );
  NAND2_X1 U5510 ( .A1(n6732), .A2(n6953), .ZN(n8869) );
  AND2_X1 U5511 ( .A1(n6847), .A2(n5183), .ZN(n5182) );
  AOI21_X1 U5512 ( .B1(n5307), .B2(n5305), .A(n4865), .ZN(n5304) );
  INV_X1 U5513 ( .A(n8950), .ZN(n5305) );
  INV_X1 U5514 ( .A(n5307), .ZN(n5306) );
  OR2_X1 U5515 ( .A1(n6552), .A2(n6551), .ZN(n6563) );
  NAND2_X1 U5516 ( .A1(n8942), .A2(n8453), .ZN(n8923) );
  OR2_X1 U5517 ( .A1(n5214), .A2(n5213), .ZN(n5212) );
  NAND2_X1 U5518 ( .A1(n6929), .A2(n6728), .ZN(n5213) );
  NAND2_X1 U5519 ( .A1(n8411), .A2(n7099), .ZN(n8939) );
  OAI21_X1 U5520 ( .B1(n8131), .B2(n5288), .A(n5287), .ZN(n8420) );
  INV_X1 U5521 ( .A(n5289), .ZN(n5288) );
  AOI21_X1 U5522 ( .B1(n5289), .B2(n5286), .A(n4890), .ZN(n5287) );
  AND2_X1 U5523 ( .A1(n5292), .A2(n5290), .ZN(n5289) );
  OR2_X1 U5524 ( .A1(n6496), .A2(n6495), .ZN(n6506) );
  INV_X1 U5525 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n9210) );
  OR2_X1 U5526 ( .A1(n6506), .A2(n9210), .ZN(n6523) );
  NAND2_X1 U5527 ( .A1(n8133), .A2(n6750), .ZN(n8336) );
  NOR2_X1 U5528 ( .A1(n8054), .A2(n10512), .ZN(n8095) );
  NAND2_X1 U5529 ( .A1(n8095), .A2(n8174), .ZN(n8134) );
  INV_X1 U5530 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n6449) );
  INV_X1 U5531 ( .A(n6901), .ZN(n5198) );
  AND2_X1 U5532 ( .A1(n6900), .A2(n6902), .ZN(n8049) );
  NAND2_X1 U5533 ( .A1(n5122), .A2(n5121), .ZN(n8054) );
  INV_X1 U5534 ( .A(n5122), .ZN(n8056) );
  NAND2_X1 U5535 ( .A1(n7046), .A2(n6712), .ZN(n5074) );
  NAND2_X1 U5536 ( .A1(n7759), .A2(n10456), .ZN(n7693) );
  NAND2_X1 U5537 ( .A1(n6605), .A2(n6604), .ZN(n8999) );
  OAI21_X1 U5538 ( .B1(n7686), .B2(n6537), .A(n6536), .ZN(n9257) );
  NAND2_X1 U5539 ( .A1(n5283), .A2(n5280), .ZN(n5277) );
  INV_X1 U5540 ( .A(n10545), .ZN(n10429) );
  INV_X1 U5541 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n6303) );
  INV_X1 U5542 ( .A(n6547), .ZN(n6558) );
  OR2_X1 U5543 ( .A1(n6418), .A2(P2_IR_REG_6__SCAN_IN), .ZN(n6429) );
  OR2_X1 U5544 ( .A1(n4952), .A2(n4947), .ZN(n4946) );
  AOI21_X1 U5545 ( .B1(n4951), .B2(n4950), .A(n4908), .ZN(n4949) );
  NAND2_X1 U5546 ( .A1(n8355), .A2(n4955), .ZN(n4948) );
  OR2_X1 U5547 ( .A1(n5669), .A2(n5668), .ZN(n5696) );
  NAND2_X1 U5548 ( .A1(n5249), .A2(n5252), .ZN(n5247) );
  NAND2_X1 U5549 ( .A1(n5231), .A2(n5230), .ZN(n5229) );
  INV_X1 U5550 ( .A(n9325), .ZN(n5230) );
  AND2_X1 U5551 ( .A1(n5840), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n5865) );
  AND2_X1 U5552 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n5549) );
  OR2_X1 U5553 ( .A1(n9422), .A2(n9351), .ZN(n5259) );
  NOR2_X1 U5554 ( .A1(n5984), .A2(n9317), .ZN(n6011) );
  AOI21_X1 U5555 ( .B1(n9716), .B2(n6083), .A(n5544), .ZN(n7610) );
  NOR2_X1 U5556 ( .A1(n5903), .A2(n5902), .ZN(n5922) );
  OR2_X1 U5557 ( .A1(n9324), .A2(n9325), .ZN(n5232) );
  OR2_X1 U5558 ( .A1(n8352), .A2(n8353), .ZN(n4957) );
  NOR2_X1 U5559 ( .A1(n5949), .A2(n9335), .ZN(n5966) );
  AND2_X1 U5560 ( .A1(n5865), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n5888) );
  NOR2_X1 U5561 ( .A1(n6123), .A2(n10242), .ZN(n6128) );
  AND2_X1 U5562 ( .A1(n9440), .A2(n9702), .ZN(n9647) );
  INV_X1 U5563 ( .A(n5261), .ZN(n5262) );
  CLKBUF_X1 U5564 ( .A(n6129), .Z(n6130) );
  NOR3_X1 U5565 ( .A1(n9789), .A2(n9994), .A3(n4981), .ZN(n9741) );
  NAND2_X1 U5566 ( .A1(n9766), .A2(n6161), .ZN(n5146) );
  NOR2_X1 U5567 ( .A1(n10014), .A2(n9816), .ZN(n9808) );
  AND2_X1 U5568 ( .A1(n9631), .A2(n9606), .ZN(n9805) );
  AND2_X1 U5569 ( .A1(n9633), .A2(n9581), .ZN(n9823) );
  NAND2_X1 U5570 ( .A1(n9838), .A2(n6242), .ZN(n9814) );
  NAND2_X1 U5571 ( .A1(n9914), .A2(n4885), .ZN(n9853) );
  INV_X1 U5572 ( .A(n10030), .ZN(n4978) );
  NOR2_X1 U5573 ( .A1(n9835), .A2(n9853), .ZN(n9833) );
  NAND2_X1 U5574 ( .A1(n9914), .A2(n4860), .ZN(n9862) );
  NAND2_X1 U5575 ( .A1(n9914), .A2(n9896), .ZN(n9891) );
  NOR2_X1 U5576 ( .A1(n10058), .A2(n4993), .ZN(n4991) );
  NAND2_X1 U5577 ( .A1(n5377), .A2(n6226), .ZN(n9942) );
  INV_X1 U5578 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n8082) );
  NOR2_X1 U5579 ( .A1(n8477), .A2(n4992), .ZN(n9966) );
  INV_X1 U5580 ( .A(n4994), .ZN(n4992) );
  OR2_X1 U5581 ( .A1(n8470), .A2(n8472), .ZN(n9963) );
  INV_X1 U5582 ( .A(n6124), .ZN(n9693) );
  INV_X1 U5583 ( .A(n9671), .ZN(n8472) );
  NOR2_X1 U5584 ( .A1(n8190), .A2(n10490), .ZN(n8277) );
  AND2_X1 U5585 ( .A1(n8277), .A2(n8282), .ZN(n8328) );
  OR2_X1 U5586 ( .A1(n5255), .A2(n5254), .ZN(n5253) );
  AND2_X1 U5587 ( .A1(n9547), .A2(n9534), .ZN(n9667) );
  INV_X1 U5588 ( .A(n7043), .ZN(n10246) );
  NAND2_X1 U5589 ( .A1(n8145), .A2(n6150), .ZN(n8147) );
  NOR2_X1 U5590 ( .A1(n4988), .A2(n8162), .ZN(n4985) );
  NAND2_X1 U5591 ( .A1(n5157), .A2(n9661), .ZN(n8145) );
  AOI21_X1 U5592 ( .B1(n9653), .B2(n5265), .A(n4863), .ZN(n5263) );
  INV_X1 U5593 ( .A(n5265), .ZN(n5264) );
  NAND2_X1 U5594 ( .A1(n10467), .A2(n4987), .ZN(n8107) );
  NOR2_X1 U5595 ( .A1(n4988), .A2(n7873), .ZN(n4987) );
  NOR2_X1 U5596 ( .A1(n7873), .A2(n7876), .ZN(n7931) );
  NOR2_X1 U5597 ( .A1(n7873), .A2(n4988), .ZN(n7949) );
  NAND2_X1 U5598 ( .A1(n7730), .A2(n7729), .ZN(n7728) );
  NAND2_X1 U5599 ( .A1(n9596), .A2(n9598), .ZN(n7729) );
  INV_X1 U5600 ( .A(n4995), .ZN(n5136) );
  INV_X1 U5601 ( .A(n7729), .ZN(n9652) );
  NAND2_X1 U5602 ( .A1(n8572), .A2(n8579), .ZN(n8571) );
  NAND2_X1 U5603 ( .A1(n10395), .A2(n10396), .ZN(n10394) );
  INV_X1 U5604 ( .A(n10242), .ZN(n6203) );
  NAND2_X1 U5605 ( .A1(n8557), .A2(n8556), .ZN(n9986) );
  AOI21_X1 U5606 ( .B1(n9994), .B2(n10502), .A(n6199), .ZN(n4975) );
  NAND2_X1 U5607 ( .A1(n6034), .A2(n6033), .ZN(n10008) );
  NAND2_X1 U5608 ( .A1(n5267), .A2(n6240), .ZN(n9840) );
  AND2_X1 U5609 ( .A1(n10401), .A2(n10504), .ZN(n10436) );
  OR2_X1 U5610 ( .A1(n7364), .A2(n9622), .ZN(n10522) );
  OR2_X1 U5611 ( .A1(n7364), .A2(n6124), .ZN(n10520) );
  OR2_X1 U5612 ( .A1(n6830), .A2(n6829), .ZN(n6831) );
  INV_X1 U5613 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5411) );
  AND2_X1 U5614 ( .A1(n6032), .A2(n6008), .ZN(n8402) );
  XNOR2_X1 U5615 ( .A(n6116), .B(n6115), .ZN(n8397) );
  AND2_X1 U5616 ( .A1(n5419), .A2(n5438), .ZN(n9591) );
  OAI21_X1 U5617 ( .B1(n5109), .B2(n5108), .A(n4911), .ZN(n5107) );
  NAND2_X1 U5618 ( .A1(n5106), .A2(n5109), .ZN(n5938) );
  NAND2_X1 U5619 ( .A1(n5899), .A2(n5110), .ZN(n5106) );
  AOI21_X1 U5620 ( .B1(n5899), .B2(n5898), .A(n5372), .ZN(n5916) );
  NAND2_X1 U5621 ( .A1(n4927), .A2(n5896), .ZN(n5880) );
  OR2_X1 U5622 ( .A1(n5860), .A2(P1_IR_REG_16__SCAN_IN), .ZN(n5861) );
  AND2_X1 U5623 ( .A1(n5859), .A2(n5899), .ZN(n7916) );
  INV_X1 U5624 ( .A(n5808), .ZN(n5086) );
  AND2_X1 U5625 ( .A1(n5834), .A2(n5812), .ZN(n5813) );
  AND2_X1 U5626 ( .A1(n5791), .A2(n5836), .ZN(n8077) );
  XNOR2_X1 U5627 ( .A(n5659), .B(n5660), .ZN(n7161) );
  NAND2_X1 U5628 ( .A1(n5635), .A2(n5634), .ZN(n5659) );
  NAND2_X1 U5629 ( .A1(n5614), .A2(n5582), .ZN(n5588) );
  NAND2_X1 U5630 ( .A1(n5588), .A2(n5587), .ZN(n5635) );
  AOI21_X1 U5631 ( .B1(n5536), .B2(n5340), .A(n5339), .ZN(n5338) );
  INV_X1 U5632 ( .A(n5556), .ZN(n5339) );
  XNOR2_X1 U5633 ( .A(n6708), .B(P2_IR_REG_23__SCAN_IN), .ZN(n7040) );
  NOR2_X1 U5634 ( .A1(n7039), .A2(P2_U3152), .ZN(n7372) );
  AND4_X1 U5635 ( .A1(n6486), .A2(n6485), .A3(n6484), .A4(n6483), .ZN(n8130)
         );
  NAND2_X1 U5636 ( .A1(n5346), .A2(n5345), .ZN(n8505) );
  NAND2_X1 U5637 ( .A1(n5051), .A2(n5057), .ZN(n7718) );
  NAND2_X1 U5638 ( .A1(n7487), .A2(n5055), .ZN(n5051) );
  NOR2_X1 U5639 ( .A1(n8644), .A2(n7117), .ZN(n7127) );
  NAND2_X1 U5640 ( .A1(n5041), .A2(n5040), .ZN(n8119) );
  NAND2_X1 U5641 ( .A1(n7921), .A2(n7920), .ZN(n5041) );
  NAND2_X1 U5642 ( .A1(n6628), .A2(n6627), .ZN(n8982) );
  NAND2_X1 U5643 ( .A1(n8371), .A2(n7103), .ZN(n8424) );
  NAND2_X1 U5644 ( .A1(n5044), .A2(n5047), .ZN(n8423) );
  AND2_X1 U5645 ( .A1(n5064), .A2(n5063), .ZN(n7353) );
  NAND2_X1 U5646 ( .A1(n5064), .A2(n5062), .ZN(n7352) );
  INV_X1 U5647 ( .A(n5061), .ZN(n5062) );
  INV_X1 U5648 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n8444) );
  CLKBUF_X1 U5649 ( .A(n8634), .Z(n8635) );
  NAND2_X1 U5650 ( .A1(n5057), .A2(n5056), .ZN(n5050) );
  INV_X1 U5651 ( .A(n5056), .ZN(n5049) );
  INV_X1 U5652 ( .A(n5053), .ZN(n5052) );
  OR2_X1 U5653 ( .A1(n7113), .A2(n5349), .ZN(n5343) );
  NAND2_X1 U5654 ( .A1(n7113), .A2(n5349), .ZN(n5342) );
  NAND2_X1 U5655 ( .A1(n8520), .A2(n7116), .ZN(n5358) );
  AND2_X1 U5656 ( .A1(n6617), .A2(n6608), .ZN(n8859) );
  NAND2_X1 U5657 ( .A1(n5036), .A2(n7053), .ZN(n7298) );
  AND2_X1 U5658 ( .A1(n7056), .A2(n7055), .ZN(n7057) );
  NAND2_X1 U5659 ( .A1(n8680), .A2(n8916), .ZN(n8662) );
  NAND2_X1 U5660 ( .A1(n5347), .A2(n8440), .ZN(n8490) );
  OR2_X1 U5661 ( .A1(n8443), .A2(n8439), .ZN(n5347) );
  INV_X1 U5662 ( .A(n9257), .ZN(n7099) );
  NAND2_X1 U5663 ( .A1(n6715), .A2(n6871), .ZN(n5188) );
  NAND2_X1 U5664 ( .A1(n5369), .A2(n7006), .ZN(n7025) );
  INV_X1 U5665 ( .A(n8609), .ZN(n8781) );
  INV_X1 U5666 ( .A(n8627), .ZN(n8821) );
  INV_X1 U5667 ( .A(n5165), .ZN(n10344) );
  NOR2_X1 U5668 ( .A1(n10341), .A2(n4869), .ZN(n10356) );
  NOR2_X1 U5669 ( .A1(n10358), .A2(n4888), .ZN(n7438) );
  NOR2_X1 U5670 ( .A1(n7512), .A2(n5167), .ZN(n7565) );
  AND2_X1 U5671 ( .A1(n7513), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n5167) );
  NOR2_X1 U5672 ( .A1(n7565), .A2(n7564), .ZN(n7563) );
  NOR2_X1 U5673 ( .A1(n7563), .A2(n5166), .ZN(n7535) );
  AND2_X1 U5674 ( .A1(n7520), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n5166) );
  NOR2_X1 U5675 ( .A1(n7535), .A2(n7534), .ZN(n7533) );
  INV_X1 U5676 ( .A(n5163), .ZN(n7597) );
  NOR2_X1 U5677 ( .A1(n7523), .A2(n7536), .ZN(n7526) );
  NAND2_X1 U5678 ( .A1(n7599), .A2(n7598), .ZN(n7891) );
  NAND2_X1 U5679 ( .A1(n7891), .A2(n5161), .ZN(n7893) );
  OR2_X1 U5680 ( .A1(n7892), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n5161) );
  NOR2_X1 U5681 ( .A1(n7966), .A2(n7967), .ZN(n8036) );
  NOR2_X1 U5682 ( .A1(n7963), .A2(n5169), .ZN(n7967) );
  AND2_X1 U5683 ( .A1(n7964), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n5169) );
  NOR2_X1 U5684 ( .A1(n8703), .A2(n8702), .ZN(n8717) );
  AOI21_X1 U5685 ( .B1(P2_REG2_REG_16__SCAN_IN), .B2(n8723), .A(n8722), .ZN(
        n8726) );
  NOR2_X1 U5686 ( .A1(n8733), .A2(n5173), .ZN(n8746) );
  NOR2_X1 U5687 ( .A1(n5174), .A2(n8455), .ZN(n5173) );
  INV_X1 U5688 ( .A(n8738), .ZN(n5174) );
  AND2_X1 U5689 ( .A1(n5113), .A2(n4921), .ZN(n8768) );
  NAND2_X1 U5690 ( .A1(n9293), .A2(n6833), .ZN(n5113) );
  NAND2_X1 U5691 ( .A1(n8771), .A2(n5119), .ZN(n10546) );
  NAND2_X1 U5692 ( .A1(n5120), .A2(n10549), .ZN(n5119) );
  OAI21_X1 U5693 ( .B1(n8831), .B2(n5317), .A(n5314), .ZN(n8784) );
  NAND2_X1 U5694 ( .A1(n5319), .A2(n5320), .ZN(n8794) );
  NAND2_X1 U5695 ( .A1(n8831), .A2(n5321), .ZN(n5319) );
  NAND2_X1 U5696 ( .A1(n8831), .A2(n5322), .ZN(n8814) );
  NAND2_X1 U5697 ( .A1(n9009), .A2(n5371), .ZN(n8881) );
  INV_X1 U5698 ( .A(n5272), .ZN(n8880) );
  NAND2_X1 U5699 ( .A1(n8897), .A2(n8896), .ZN(n9009) );
  OAI21_X1 U5700 ( .B1(n8912), .B2(n5187), .A(n5185), .ZN(n8886) );
  NAND2_X1 U5701 ( .A1(n8912), .A2(n6731), .ZN(n8900) );
  NAND2_X1 U5702 ( .A1(n8949), .A2(n6557), .ZN(n8450) );
  NAND2_X1 U5703 ( .A1(n8344), .A2(n6728), .ZN(n8408) );
  NAND2_X1 U5704 ( .A1(n6727), .A2(n6726), .ZN(n8341) );
  NAND2_X1 U5705 ( .A1(n5291), .A2(n5292), .ZN(n8335) );
  NAND2_X1 U5706 ( .A1(n8131), .A2(n5293), .ZN(n5291) );
  NAND2_X1 U5707 ( .A1(n5294), .A2(n5293), .ZN(n8234) );
  NAND2_X1 U5708 ( .A1(n6502), .A2(n8128), .ZN(n5294) );
  NAND2_X1 U5709 ( .A1(n7984), .A2(n6475), .ZN(n8090) );
  NAND2_X1 U5710 ( .A1(n5192), .A2(n6909), .ZN(n8092) );
  NAND2_X1 U5711 ( .A1(n7987), .A2(n6911), .ZN(n5192) );
  NAND2_X1 U5712 ( .A1(n5200), .A2(n6896), .ZN(n7806) );
  NAND2_X1 U5713 ( .A1(n7788), .A2(n7787), .ZN(n5200) );
  NAND2_X1 U5714 ( .A1(n5282), .A2(n6417), .ZN(n7786) );
  NAND2_X1 U5715 ( .A1(n5283), .A2(n4858), .ZN(n5282) );
  OAI21_X1 U5716 ( .B1(n7753), .B2(n5210), .A(n5207), .ZN(n7673) );
  NAND2_X1 U5717 ( .A1(n7752), .A2(n6722), .ZN(n7691) );
  AOI22_X1 U5718 ( .A1(n7304), .A2(n7441), .B1(P1_DATAO_REG_3__SCAN_IN), .B2(
        n6379), .ZN(n5189) );
  NAND2_X1 U5719 ( .A1(n10155), .A2(n6711), .ZN(n10454) );
  OR2_X1 U5720 ( .A1(n6754), .A2(n7288), .ZN(n8777) );
  INV_X1 U5721 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n9222) );
  XNOR2_X1 U5722 ( .A(n6680), .B(P2_IR_REG_24__SCAN_IN), .ZN(n10327) );
  NAND2_X1 U5723 ( .A1(n6679), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6680) );
  AND2_X1 U5724 ( .A1(n6675), .A2(n6674), .ZN(n10328) );
  INV_X1 U5725 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n6315) );
  NAND2_X1 U5726 ( .A1(n6674), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6317) );
  OR2_X1 U5727 ( .A1(n6685), .A2(n6684), .ZN(n8435) );
  CLKBUF_X1 U5728 ( .A(n6712), .Z(n8350) );
  AND2_X1 U5729 ( .A1(n6476), .A2(n6463), .ZN(n7602) );
  AND2_X1 U5730 ( .A1(n6356), .A2(n6286), .ZN(n6375) );
  NAND2_X1 U5731 ( .A1(n4967), .A2(n4966), .ZN(n9324) );
  NAND2_X1 U5732 ( .A1(n4962), .A2(n9399), .ZN(n4966) );
  NAND2_X1 U5733 ( .A1(n9402), .A2(n9400), .ZN(n4967) );
  NAND2_X1 U5734 ( .A1(n5257), .A2(n4968), .ZN(n4962) );
  OR2_X1 U5735 ( .A1(n5529), .A2(n7143), .ZN(n5408) );
  INV_X1 U5736 ( .A(n5406), .ZN(n5407) );
  NAND2_X1 U5737 ( .A1(n5223), .A2(n5228), .ZN(n9334) );
  OR2_X1 U5738 ( .A1(n9324), .A2(n5229), .ZN(n5223) );
  INV_X1 U5739 ( .A(n9708), .ZN(n9978) );
  INV_X1 U5740 ( .A(n9710), .ZN(n8387) );
  NAND2_X1 U5741 ( .A1(n9343), .A2(n9344), .ZN(n9411) );
  INV_X1 U5742 ( .A(n9705), .ZN(n9947) );
  AND2_X1 U5743 ( .A1(n5259), .A2(n4861), .ZN(n9360) );
  AND2_X1 U5744 ( .A1(n5232), .A2(n5914), .ZN(n9381) );
  OAI21_X1 U5745 ( .B1(n8355), .B2(n5758), .A(n4957), .ZN(n8365) );
  AOI21_X1 U5746 ( .B1(n5225), .B2(n9331), .A(n9330), .ZN(n5224) );
  INV_X1 U5747 ( .A(n5228), .ZN(n5225) );
  NAND2_X1 U5748 ( .A1(n7336), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9392) );
  NAND2_X1 U5749 ( .A1(n6131), .A2(n7621), .ZN(n9431) );
  NAND2_X1 U5750 ( .A1(n6049), .A2(n6048), .ZN(n10003) );
  INV_X1 U5751 ( .A(n9431), .ZN(n9417) );
  AND2_X1 U5752 ( .A1(n6053), .A2(n6135), .ZN(n9776) );
  NAND2_X1 U5753 ( .A1(n4943), .A2(n4942), .ZN(n9415) );
  NAND2_X1 U5754 ( .A1(n5252), .A2(n9410), .ZN(n4942) );
  INV_X1 U5755 ( .A(n9409), .ZN(n9435) );
  AND2_X1 U5756 ( .A1(n6189), .A2(n6188), .ZN(n7368) );
  NAND2_X1 U5757 ( .A1(n5864), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5433) );
  XNOR2_X1 U5758 ( .A(n9986), .B(n9989), .ZN(n9988) );
  INV_X1 U5759 ( .A(n9742), .ZN(n9993) );
  INV_X1 U5760 ( .A(n9751), .ZN(n9752) );
  XNOR2_X1 U5761 ( .A(n9749), .B(n9748), .ZN(n9753) );
  AOI22_X1 U5762 ( .A1(n9750), .A2(n10391), .B1(n10393), .B2(n9785), .ZN(n9751) );
  AOI211_X1 U5763 ( .C1(n9774), .C2(n10397), .A(n9773), .B(n9772), .ZN(n10006)
         );
  NAND2_X1 U5764 ( .A1(n9800), .A2(n6244), .ZN(n9795) );
  AND2_X1 U5765 ( .A1(n5983), .A2(n5982), .ZN(n9820) );
  OAI21_X1 U5766 ( .B1(n4935), .B2(n5133), .A(n5131), .ZN(n9849) );
  NAND2_X1 U5767 ( .A1(n9868), .A2(n9869), .ZN(n9867) );
  NAND2_X1 U5768 ( .A1(n4935), .A2(n9572), .ZN(n9868) );
  INV_X1 U5769 ( .A(n5236), .ZN(n9876) );
  AOI21_X1 U5770 ( .B1(n9890), .B2(n9889), .A(n5239), .ZN(n5236) );
  NAND2_X1 U5771 ( .A1(n9944), .A2(n6229), .ZN(n9930) );
  NAND2_X1 U5772 ( .A1(n5152), .A2(n5153), .ZN(n9924) );
  AND2_X1 U5773 ( .A1(n4913), .A2(n8478), .ZN(n10073) );
  NAND2_X1 U5774 ( .A1(n8144), .A2(n6216), .ZN(n8181) );
  NAND2_X1 U5775 ( .A1(n7937), .A2(n5265), .ZN(n7944) );
  INV_X1 U5776 ( .A(n10368), .ZN(n9918) );
  INV_X1 U5777 ( .A(n10376), .ZN(n10409) );
  NAND2_X2 U5778 ( .A1(n5481), .A2(n5480), .ZN(n8590) );
  OR2_X1 U5779 ( .A1(n5529), .A2(n7149), .ZN(n5480) );
  INV_X1 U5780 ( .A(n5470), .ZN(n5481) );
  INV_X1 U5781 ( .A(n9969), .ZN(n10367) );
  NAND2_X1 U5782 ( .A1(n5260), .A2(n5636), .ZN(n5440) );
  INV_X1 U5783 ( .A(n10531), .ZN(n10529) );
  AOI21_X1 U5784 ( .B1(n10121), .B2(n6100), .A(n6099), .ZN(n10103) );
  NAND2_X1 U5785 ( .A1(n5424), .A2(n5423), .ZN(n10104) );
  NOR2_X1 U5786 ( .A1(P1_IR_REG_29__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), .ZN(
        n5423) );
  INV_X1 U5787 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n10105) );
  NAND2_X1 U5788 ( .A1(n5429), .A2(P1_IR_REG_29__SCAN_IN), .ZN(n4997) );
  NAND2_X1 U5789 ( .A1(n5430), .A2(n4999), .ZN(n4998) );
  INV_X1 U5790 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n4999) );
  AND2_X1 U5791 ( .A1(n7142), .A2(P1_U3084), .ZN(n10114) );
  INV_X1 U5792 ( .A(n9441), .ZN(n8515) );
  INV_X1 U5793 ( .A(n9591), .ZN(n9685) );
  NAND2_X1 U5794 ( .A1(n5088), .A2(n5087), .ZN(n5809) );
  NAND2_X1 U5795 ( .A1(n5759), .A2(n5351), .ZN(n5760) );
  NAND2_X1 U5796 ( .A1(n5333), .A2(n5716), .ZN(n5720) );
  AND2_X1 U5797 ( .A1(n5636), .A2(n5384), .ZN(n5691) );
  NAND2_X1 U5798 ( .A1(n5537), .A2(n5536), .ZN(n5557) );
  NAND2_X1 U5799 ( .A1(n5531), .A2(n5530), .ZN(n5537) );
  NOR2_X1 U5800 ( .A1(n10216), .A2(n10215), .ZN(n10218) );
  AOI21_X1 U5801 ( .B1(n5258), .B2(n9351), .A(n4897), .ZN(n5256) );
  NAND2_X1 U5802 ( .A1(n7487), .A2(n7072), .ZN(n7578) );
  AOI211_X1 U5803 ( .C1(n8993), .C2(n8641), .A(n8619), .B(n8618), .ZN(n8620)
         );
  AOI21_X1 U5804 ( .B1(n8763), .B2(n8008), .A(n5176), .ZN(n5175) );
  NAND2_X1 U5805 ( .A1(n5179), .A2(n10461), .ZN(n5178) );
  INV_X1 U5806 ( .A(n5177), .ZN(n5176) );
  INV_X1 U5807 ( .A(n6809), .ZN(n6810) );
  OAI21_X1 U5808 ( .B1(n8963), .B2(n10466), .A(n6808), .ZN(n6809) );
  NAND2_X1 U5809 ( .A1(n5380), .A2(n5373), .ZN(P2_U3268) );
  AND2_X1 U5810 ( .A1(n6760), .A2(n6759), .ZN(n5373) );
  OAI21_X1 U5811 ( .B1(n6772), .B2(n6119), .A(n9413), .ZN(n6145) );
  NAND2_X1 U5812 ( .A1(n5012), .A2(n5011), .ZN(P1_U3240) );
  OR2_X1 U5813 ( .A1(n9700), .A2(n9699), .ZN(n5011) );
  NAND2_X1 U5814 ( .A1(n5014), .A2(n5013), .ZN(n5012) );
  NAND2_X1 U5815 ( .A1(n5139), .A2(n5138), .ZN(n6262) );
  OR2_X1 U5816 ( .A1(n5140), .A2(n10419), .ZN(n5138) );
  AOI211_X1 U5817 ( .C1(n10368), .C2(n8599), .A(n8598), .B(n8597), .ZN(n8600)
         );
  OR2_X1 U5818 ( .A1(n10531), .A2(n4973), .ZN(n4972) );
  NAND2_X1 U5819 ( .A1(n10086), .A2(n10531), .ZN(n4974) );
  INV_X1 U5820 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n4973) );
  NAND2_X1 U5821 ( .A1(n5257), .A2(n5256), .ZN(n9402) );
  INV_X1 U5822 ( .A(n5286), .ZN(n5293) );
  OR3_X1 U5823 ( .A1(n9647), .A2(n6117), .A3(n9689), .ZN(n4857) );
  OR2_X1 U5824 ( .A1(n7681), .A2(n7789), .ZN(n4858) );
  AND2_X1 U5825 ( .A1(n6330), .A2(n6329), .ZN(n8879) );
  INV_X1 U5826 ( .A(n8879), .ZN(n9004) );
  AND2_X1 U5827 ( .A1(n9896), .A2(n4979), .ZN(n4859) );
  INV_X1 U5828 ( .A(n7859), .ZN(n5285) );
  AND2_X1 U5829 ( .A1(n9866), .A2(n4859), .ZN(n4860) );
  AND2_X1 U5830 ( .A1(n9495), .A2(n9496), .ZN(n9869) );
  INV_X1 U5831 ( .A(n9869), .ZN(n5133) );
  NAND2_X1 U5832 ( .A1(n5852), .A2(n5851), .ZN(n4861) );
  NAND2_X1 U5833 ( .A1(n8623), .A2(n4887), .ZN(n8671) );
  NAND2_X1 U5834 ( .A1(n6646), .A2(n6645), .ZN(n8970) );
  INV_X1 U5835 ( .A(n5353), .ZN(n5351) );
  AND2_X1 U5836 ( .A1(n9267), .A2(n8691), .ZN(n4862) );
  INV_X1 U5837 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5418) );
  AND2_X1 U5838 ( .A1(n7979), .A2(n10467), .ZN(n4863) );
  INV_X1 U5839 ( .A(n5644), .ZN(n5822) );
  INV_X2 U5840 ( .A(n5822), .ZN(n8561) );
  AND2_X1 U5841 ( .A1(n10111), .A2(n8604), .ZN(n5644) );
  OR2_X1 U5842 ( .A1(n8685), .A2(n8970), .ZN(n4864) );
  INV_X1 U5843 ( .A(n8840), .ZN(n8987) );
  AND2_X1 U5844 ( .A1(n8453), .A2(n8428), .ZN(n4865) );
  OR2_X1 U5845 ( .A1(n9004), .A2(n8887), .ZN(n4866) );
  AND2_X1 U5846 ( .A1(n5253), .A2(n6217), .ZN(n4867) );
  NAND2_X1 U5847 ( .A1(n6858), .A2(n6860), .ZN(n8128) );
  INV_X1 U5848 ( .A(n9344), .ZN(n5252) );
  INV_X1 U5849 ( .A(n5454), .ZN(n5987) );
  AND2_X1 U5850 ( .A1(n7209), .A2(n5443), .ZN(n5454) );
  AND3_X1 U5851 ( .A1(n5260), .A2(n5636), .A3(n5160), .ZN(n4868) );
  AND2_X1 U5852 ( .A1(n10349), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n4869) );
  INV_X1 U5853 ( .A(n6382), .ZN(n6433) );
  NAND2_X1 U5854 ( .A1(n6836), .A2(n6835), .ZN(n10549) );
  INV_X1 U5855 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n9294) );
  NAND2_X1 U5856 ( .A1(n6877), .A2(n6876), .ZN(n6721) );
  NAND2_X1 U5857 ( .A1(n8235), .A2(n4915), .ZN(n5286) );
  NAND2_X1 U5858 ( .A1(n5318), .A2(n5320), .ZN(n5317) );
  AND2_X1 U5859 ( .A1(n5227), .A2(n9331), .ZN(n4870) );
  NAND2_X1 U5860 ( .A1(n6186), .A2(n6185), .ZN(n9994) );
  AND3_X1 U5861 ( .A1(n6354), .A2(n6353), .A3(n6352), .ZN(n4871) );
  NAND2_X1 U5862 ( .A1(n8614), .A2(n8527), .ZN(n8528) );
  OR3_X1 U5863 ( .A1(n9687), .A2(n10411), .A3(n9688), .ZN(n4872) );
  OR2_X1 U5864 ( .A1(n9998), .A2(n9768), .ZN(n9636) );
  INV_X1 U5865 ( .A(n5043), .ZN(n5042) );
  NAND2_X1 U5866 ( .A1(n7086), .A2(n7087), .ZN(n5043) );
  AND2_X1 U5867 ( .A1(n6536), .A2(n8537), .ZN(n4873) );
  NAND2_X1 U5868 ( .A1(n6172), .A2(n6171), .ZN(n6781) );
  INV_X1 U5869 ( .A(n6781), .ZN(n4982) );
  AND2_X1 U5870 ( .A1(n8098), .A2(n7986), .ZN(n4874) );
  OR3_X1 U5871 ( .A1(n7029), .A2(n6715), .A3(n10378), .ZN(n4875) );
  NAND2_X1 U5872 ( .A1(n8636), .A2(n5330), .ZN(n8622) );
  NAND2_X1 U5873 ( .A1(n6074), .A2(n6073), .ZN(n9998) );
  INV_X1 U5874 ( .A(n5065), .ZN(n8644) );
  OR2_X1 U5875 ( .A1(n9358), .A2(n5876), .ZN(n4876) );
  NAND2_X1 U5876 ( .A1(n8623), .A2(n8532), .ZN(n8668) );
  NAND2_X1 U5877 ( .A1(n8634), .A2(n8637), .ZN(n8636) );
  OR2_X1 U5878 ( .A1(n4982), .A2(n9703), .ZN(n4877) );
  NOR2_X1 U5879 ( .A1(n7127), .A2(n7126), .ZN(n4878) );
  NAND2_X1 U5880 ( .A1(n9367), .A2(n6030), .ZN(n9343) );
  AND2_X1 U5881 ( .A1(n4951), .A2(n5738), .ZN(n4879) );
  NAND2_X1 U5882 ( .A1(n8849), .A2(n8840), .ZN(n8834) );
  INV_X1 U5883 ( .A(n8834), .ZN(n5124) );
  AND2_X1 U5884 ( .A1(n5221), .A2(n6962), .ZN(n4880) );
  NAND2_X1 U5885 ( .A1(n5069), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6701) );
  NAND3_X1 U5886 ( .A1(n9368), .A2(n9370), .A3(n9369), .ZN(n9367) );
  AND2_X1 U5887 ( .A1(n6245), .A2(n6244), .ZN(n4881) );
  AND2_X1 U5888 ( .A1(n6241), .A2(n6240), .ZN(n4882) );
  INV_X1 U5889 ( .A(n5281), .ZN(n5280) );
  NAND2_X1 U5890 ( .A1(n4858), .A2(n5284), .ZN(n5281) );
  AND2_X1 U5891 ( .A1(n4938), .A2(n4941), .ZN(n4883) );
  NAND2_X1 U5892 ( .A1(n7611), .A2(n7610), .ZN(n4884) );
  AND2_X1 U5893 ( .A1(n4860), .A2(n4978), .ZN(n4885) );
  AND2_X1 U5894 ( .A1(n5359), .A2(n8655), .ZN(n4886) );
  AND2_X1 U5895 ( .A1(n8535), .A2(n8532), .ZN(n4887) );
  AND2_X1 U5896 ( .A1(n10363), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n4888) );
  INV_X1 U5897 ( .A(n5125), .ZN(n8858) );
  NOR2_X1 U5898 ( .A1(n8874), .A2(n8999), .ZN(n5125) );
  NAND2_X1 U5899 ( .A1(n5376), .A2(n5421), .ZN(n4889) );
  NOR2_X1 U5900 ( .A1(n9262), .A2(n8409), .ZN(n4890) );
  INV_X1 U5901 ( .A(n5356), .ZN(n5355) );
  NOR2_X1 U5902 ( .A1(n5780), .A2(SI_13_), .ZN(n5356) );
  AND2_X1 U5903 ( .A1(n5212), .A2(n6928), .ZN(n4891) );
  AND2_X1 U5904 ( .A1(n7030), .A2(n4875), .ZN(n4892) );
  AND2_X1 U5905 ( .A1(n9455), .A2(n9624), .ZN(n9653) );
  INV_X1 U5906 ( .A(n4969), .ZN(n4968) );
  AND2_X1 U5907 ( .A1(n4948), .A2(n4951), .ZN(n4893) );
  NOR2_X1 U5908 ( .A1(n8801), .A2(n8821), .ZN(n4894) );
  INV_X1 U5909 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5160) );
  INV_X1 U5910 ( .A(n5145), .ZN(n5144) );
  NAND2_X1 U5911 ( .A1(n9678), .A2(n9636), .ZN(n5145) );
  AND2_X1 U5912 ( .A1(n5663), .A2(n5662), .ZN(n4895) );
  AND4_X1 U5913 ( .A1(n6428), .A2(n6427), .A3(n6426), .A4(n6425), .ZN(n7719)
         );
  NAND2_X1 U5914 ( .A1(n10490), .A2(n9712), .ZN(n4896) );
  AND2_X1 U5915 ( .A1(n9358), .A2(n5876), .ZN(n4897) );
  NAND2_X1 U5916 ( .A1(n9673), .A2(n9443), .ZN(n4898) );
  OR2_X1 U5917 ( .A1(n4965), .A2(n4969), .ZN(n4899) );
  INV_X1 U5918 ( .A(n5057), .ZN(n5054) );
  NAND2_X1 U5919 ( .A1(n7073), .A2(n7074), .ZN(n5057) );
  NAND2_X1 U5920 ( .A1(n9377), .A2(n5914), .ZN(n4900) );
  NAND2_X1 U5921 ( .A1(n5921), .A2(n5920), .ZN(n10035) );
  INV_X1 U5922 ( .A(n6891), .ZN(n5205) );
  AND2_X1 U5923 ( .A1(n5110), .A2(n5937), .ZN(n4901) );
  INV_X1 U5924 ( .A(n10111), .ZN(n4996) );
  AND2_X1 U5925 ( .A1(n6151), .A2(n9546), .ZN(n4902) );
  NOR2_X1 U5926 ( .A1(n5356), .A2(n5784), .ZN(n5087) );
  AND2_X1 U5927 ( .A1(n9823), .A2(n9503), .ZN(n4903) );
  AND2_X1 U5928 ( .A1(n9507), .A2(n9796), .ZN(n4904) );
  INV_X1 U5929 ( .A(n4952), .ZN(n4951) );
  NAND2_X1 U5930 ( .A1(n4953), .A2(n8361), .ZN(n4952) );
  AND2_X1 U5931 ( .A1(n9508), .A2(n9770), .ZN(n4905) );
  AND2_X1 U5932 ( .A1(n5137), .A2(n4975), .ZN(n4906) );
  AND2_X1 U5933 ( .A1(n5151), .A2(n5153), .ZN(n4907) );
  INV_X1 U5934 ( .A(n5317), .ZN(n5316) );
  AND2_X2 U5935 ( .A1(n7209), .A2(n7734), .ZN(n5435) );
  NAND2_X1 U5936 ( .A1(n5636), .A2(n5262), .ZN(n5722) );
  AND2_X1 U5937 ( .A1(n6652), .A2(n6651), .ZN(n8674) );
  INV_X1 U5938 ( .A(n8674), .ZN(n8685) );
  XOR2_X1 U5939 ( .A(n5804), .B(n6765), .Z(n4908) );
  INV_X1 U5940 ( .A(n7068), .ZN(n8537) );
  INV_X1 U5941 ( .A(n9922), .ZN(n5148) );
  AND2_X1 U5942 ( .A1(n5294), .A2(n4915), .ZN(n4909) );
  NAND2_X1 U5943 ( .A1(n8951), .A2(n8950), .ZN(n8949) );
  NAND2_X1 U5944 ( .A1(n6791), .A2(n6790), .ZN(n8960) );
  INV_X1 U5945 ( .A(n8960), .ZN(n5118) );
  AND2_X1 U5946 ( .A1(n5026), .A2(n9950), .ZN(n4910) );
  NAND2_X1 U5947 ( .A1(n9914), .A2(n4859), .ZN(n4980) );
  INV_X1 U5948 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n4970) );
  INV_X1 U5949 ( .A(SI_12_), .ZN(n9153) );
  OR2_X1 U5950 ( .A1(n5936), .A2(SI_20_), .ZN(n4911) );
  AND2_X1 U5951 ( .A1(n5919), .A2(n5918), .ZN(n4912) );
  INV_X1 U5952 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5271) );
  XNOR2_X1 U5953 ( .A(n5410), .B(P1_IR_REG_26__SCAN_IN), .ZN(n6096) );
  NAND2_X1 U5954 ( .A1(n9441), .A2(n9591), .ZN(n6117) );
  INV_X1 U5955 ( .A(n7671), .ZN(n5283) );
  INV_X1 U5956 ( .A(n6922), .ZN(n5290) );
  INV_X1 U5957 ( .A(n6712), .ZN(n5072) );
  OR2_X1 U5958 ( .A1(n8477), .A2(n6157), .ZN(n4913) );
  OR2_X1 U5959 ( .A1(n6045), .A2(SI_25_), .ZN(n4914) );
  OR2_X1 U5960 ( .A1(n8139), .A2(n8244), .ZN(n4915) );
  NAND2_X1 U5961 ( .A1(n5296), .A2(n5295), .ZN(n8131) );
  INV_X1 U5962 ( .A(n10039), .ZN(n4979) );
  NAND2_X1 U5963 ( .A1(n5414), .A2(n5413), .ZN(n6094) );
  NOR3_X1 U5964 ( .A1(n10274), .A2(n10273), .A3(n10272), .ZN(n4916) );
  NAND2_X1 U5965 ( .A1(n5277), .A2(n5278), .ZN(n7803) );
  AND2_X1 U5966 ( .A1(n9940), .A2(n10397), .ZN(n4917) );
  AND2_X1 U5967 ( .A1(n7937), .A2(n6214), .ZN(n4918) );
  AND2_X1 U5968 ( .A1(n6071), .A2(n9133), .ZN(n4919) );
  INV_X1 U5969 ( .A(n9940), .ZN(n10419) );
  AND2_X1 U5970 ( .A1(n8112), .A2(n6215), .ZN(n4920) );
  NAND2_X1 U5971 ( .A1(n6820), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n4921) );
  AND2_X1 U5972 ( .A1(n8147), .A2(n9546), .ZN(n4922) );
  AND2_X1 U5973 ( .A1(n5041), .A2(n5043), .ZN(n4923) );
  AND2_X1 U5974 ( .A1(n5093), .A2(n6812), .ZN(n4924) );
  INV_X1 U5975 ( .A(n8196), .ZN(n5121) );
  NAND4_X1 U5976 ( .A1(n6346), .A2(n6345), .A3(n6344), .A4(n6343), .ZN(n8700)
         );
  INV_X1 U5977 ( .A(n8700), .ZN(n4928) );
  INV_X1 U5978 ( .A(n7343), .ZN(n5060) );
  AND2_X1 U5979 ( .A1(n5074), .A2(n8008), .ZN(n4925) );
  INV_X1 U5980 ( .A(n6307), .ZN(n9299) );
  INV_X1 U5981 ( .A(n8783), .ZN(n5312) );
  NAND2_X1 U5982 ( .A1(n5316), .A2(n8783), .ZN(n5313) );
  NOR4_X1 U5983 ( .A1(n6853), .A2(n6852), .A3(n8783), .A4(n6851), .ZN(n6854)
         );
  NOR2_X1 U5984 ( .A1(n7142), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10107) );
  OR2_X2 U5985 ( .A1(n7209), .A2(n7038), .ZN(n9719) );
  NAND2_X1 U5986 ( .A1(n6096), .A2(n5417), .ZN(n7209) );
  NAND2_X1 U5987 ( .A1(n5612), .A2(n5611), .ZN(n5614) );
  NAND2_X1 U5988 ( .A1(n5333), .A2(n5332), .ZN(n5740) );
  AOI21_X1 U5989 ( .B1(n5352), .B2(n5087), .A(n5086), .ZN(n4926) );
  OAI21_X1 U5990 ( .B1(n9755), .B2(n9748), .A(n6250), .ZN(n6263) );
  NAND2_X1 U5991 ( .A1(n5080), .A2(n5079), .ZN(n5686) );
  NAND2_X1 U5992 ( .A1(n5237), .A2(n4936), .ZN(n6236) );
  OAI22_X1 U5993 ( .A1(n5855), .A2(n5854), .B1(SI_16_), .B2(n5853), .ZN(n5858)
         );
  NAND2_X1 U5994 ( .A1(n5713), .A2(n5712), .ZN(n5333) );
  NAND2_X1 U5995 ( .A1(n6740), .A2(n6739), .ZN(n7009) );
  AOI21_X2 U5996 ( .B1(n8820), .B2(n8813), .A(n6736), .ZN(n8796) );
  AOI21_X1 U5997 ( .B1(n5899), .B2(n4901), .A(n5107), .ZN(n5943) );
  NAND2_X1 U5998 ( .A1(n5336), .A2(n5338), .ZN(n5562) );
  NAND2_X1 U5999 ( .A1(n4926), .A2(n5085), .ZN(n5814) );
  NAND2_X1 U6000 ( .A1(n4974), .A2(n4972), .ZN(P1_U3552) );
  INV_X1 U6001 ( .A(n5878), .ZN(n4927) );
  AND2_X1 U6002 ( .A1(n5899), .A2(n5894), .ZN(n5878) );
  MUX2_X2 U6004 ( .A(n6997), .B(n6868), .S(n6869), .Z(n6875) );
  NAND2_X1 U6005 ( .A1(n4929), .A2(n6900), .ZN(n6906) );
  NAND3_X1 U6006 ( .A1(n6899), .A2(n6898), .A3(n7805), .ZN(n4929) );
  AOI21_X2 U6007 ( .B1(n4930), .B2(n7004), .A(n7003), .ZN(n7028) );
  NAND3_X1 U6008 ( .A1(n7000), .A2(n6998), .A3(n4931), .ZN(n4930) );
  NAND3_X1 U6010 ( .A1(n4933), .A2(n6956), .A3(n6964), .ZN(n6959) );
  NAND3_X1 U6011 ( .A1(n6948), .A2(n8882), .A3(n6953), .ZN(n4933) );
  OAI21_X1 U6012 ( .B1(n6907), .B2(n6908), .A(n4934), .ZN(n6916) );
  OAI211_X1 U6013 ( .C1(n5188), .C2(n7024), .A(n4892), .B(n7025), .ZN(n5078)
         );
  NAND2_X1 U6014 ( .A1(n5156), .A2(n4902), .ZN(n5155) );
  AOI21_X1 U6015 ( .B1(n6269), .B2(n10397), .A(n6270), .ZN(n6271) );
  AOI21_X2 U6016 ( .B1(n8274), .B2(n9667), .A(n9447), .ZN(n8324) );
  NOR2_X1 U6017 ( .A1(n6159), .A2(n9444), .ZN(n9898) );
  OAI21_X1 U6018 ( .B1(n8473), .B2(n9671), .A(n9554), .ZN(n9974) );
  NAND2_X1 U6019 ( .A1(n8913), .A2(n5302), .ZN(n8912) );
  NAND2_X1 U6020 ( .A1(n5088), .A2(n5355), .ZN(n5785) );
  OAI21_X1 U6021 ( .B1(n8863), .B2(n5218), .A(n5215), .ZN(n6735) );
  AOI21_X1 U6022 ( .B1(n7023), .B2(n7022), .A(n7021), .ZN(n7026) );
  NOR2_X1 U6023 ( .A1(n10356), .A2(n10355), .ZN(n10354) );
  NAND2_X1 U6024 ( .A1(n8761), .A2(n5180), .ZN(n5179) );
  OAI21_X1 U6025 ( .B1(n8762), .B2(n10353), .A(n10335), .ZN(n5181) );
  NAND2_X1 U6026 ( .A1(n5178), .A2(n5175), .ZN(P2_U3264) );
  NAND2_X1 U6027 ( .A1(n5690), .A2(n5689), .ZN(n5713) );
  INV_X1 U6028 ( .A(n5309), .ZN(n6789) );
  INV_X1 U6029 ( .A(n8921), .ZN(n5302) );
  NAND2_X1 U6030 ( .A1(n5303), .A2(n5301), .ZN(n8920) );
  INV_X1 U6031 ( .A(n9451), .ZN(n9450) );
  NOR2_X1 U6032 ( .A1(n5010), .A2(n5009), .ZN(n5008) );
  INV_X1 U6033 ( .A(n5154), .ZN(n8182) );
  NAND2_X1 U6034 ( .A1(n9793), .A2(n6246), .ZN(n9771) );
  INV_X1 U6035 ( .A(n9889), .ZN(n5238) );
  NAND2_X2 U6036 ( .A1(n5741), .A2(n5742), .ZN(n5759) );
  NAND2_X4 U6037 ( .A1(n10401), .A2(n5443), .ZN(n6081) );
  XNOR2_X1 U6038 ( .A(n5543), .B(n6765), .ZN(n7611) );
  OR2_X1 U6039 ( .A1(n4868), .A2(n4940), .ZN(n4937) );
  NAND2_X1 U6040 ( .A1(n4868), .A2(n5418), .ZN(n4938) );
  NAND2_X1 U6041 ( .A1(n4937), .A2(n4939), .ZN(n5438) );
  OR2_X1 U6042 ( .A1(n4868), .A2(n5409), .ZN(n5420) );
  NAND2_X1 U6043 ( .A1(n9367), .A2(n4944), .ZN(n4943) );
  NAND3_X1 U6044 ( .A1(n4946), .A2(n4945), .A3(n4949), .ZN(n9304) );
  NAND2_X1 U6045 ( .A1(n8248), .A2(n4879), .ZN(n4945) );
  OAI21_X2 U6046 ( .B1(n8248), .B2(n8249), .A(n5738), .ZN(n8355) );
  NAND2_X1 U6047 ( .A1(n5256), .A2(n5893), .ZN(n4969) );
  NAND3_X1 U6048 ( .A1(n4977), .A2(n4976), .A3(n4906), .ZN(n10086) );
  INV_X1 U6049 ( .A(n4980), .ZN(n9877) );
  NOR2_X1 U6050 ( .A1(n9789), .A2(n10003), .ZN(n9759) );
  INV_X1 U6051 ( .A(n7873), .ZN(n4986) );
  NAND3_X1 U6052 ( .A1(n4986), .A2(n10467), .A3(n4985), .ZN(n8152) );
  INV_X1 U6053 ( .A(n8477), .ZN(n4990) );
  NAND2_X1 U6054 ( .A1(n4990), .A2(n4991), .ZN(n9936) );
  NOR2_X1 U6055 ( .A1(n8477), .A2(n4993), .ZN(n9954) );
  NAND2_X1 U6056 ( .A1(n5135), .A2(n4995), .ZN(n5134) );
  NAND2_X1 U6057 ( .A1(n10394), .A2(n4995), .ZN(n9588) );
  XNOR2_X2 U6058 ( .A(n5425), .B(n10105), .ZN(n8604) );
  NAND2_X1 U6059 ( .A1(n5000), .A2(n5001), .ZN(n9510) );
  NAND2_X1 U6060 ( .A1(n9505), .A2(n5003), .ZN(n5000) );
  OR2_X1 U6061 ( .A1(n5006), .A2(n9504), .ZN(n5005) );
  AND2_X2 U6062 ( .A1(n9625), .A2(n9623), .ZN(n9451) );
  NAND3_X1 U6063 ( .A1(n9673), .A2(n9490), .A3(n5151), .ZN(n5025) );
  AND3_X2 U6064 ( .A1(n5636), .A2(n5260), .A3(n5159), .ZN(n6113) );
  NAND4_X1 U6065 ( .A1(n5386), .A2(n5387), .A3(n5388), .A4(n5389), .ZN(n5035)
         );
  OAI21_X1 U6066 ( .B1(n7257), .B2(n7258), .A(n5036), .ZN(n7260) );
  NAND2_X1 U6067 ( .A1(n7258), .A2(n7257), .ZN(n5036) );
  OAI22_X2 U6068 ( .A1(n7900), .A2(n7901), .B1(n7085), .B2(n7084), .ZN(n7921)
         );
  NAND2_X1 U6069 ( .A1(n8372), .A2(n5047), .ZN(n5046) );
  NAND2_X1 U6070 ( .A1(n7818), .A2(n7817), .ZN(n7816) );
  NAND3_X1 U6071 ( .A1(n5063), .A2(n5060), .A3(n7354), .ZN(n5059) );
  AND2_X1 U6072 ( .A1(n5059), .A2(n7067), .ZN(n5058) );
  NAND2_X1 U6073 ( .A1(n5063), .A2(n7354), .ZN(n5061) );
  OAI21_X2 U6074 ( .B1(n5065), .B2(n7126), .A(n4886), .ZN(n8654) );
  OR2_X2 U6075 ( .A1(n8645), .A2(n8646), .ZN(n5065) );
  NAND2_X1 U6076 ( .A1(n6582), .A2(n5070), .ZN(n5068) );
  NAND2_X1 U6077 ( .A1(n6582), .A2(n6581), .ZN(n5069) );
  NAND3_X1 U6078 ( .A1(n9735), .A2(n5076), .A3(n5075), .ZN(n5328) );
  NAND2_X1 U6079 ( .A1(n5077), .A2(n7036), .ZN(P2_U3244) );
  NAND2_X1 U6080 ( .A1(n5078), .A2(n7031), .ZN(n5077) );
  NAND2_X1 U6081 ( .A1(n5614), .A2(n5081), .ZN(n5080) );
  NAND2_X1 U6082 ( .A1(n5351), .A2(n5087), .ZN(n5085) );
  NAND2_X1 U6083 ( .A1(n6169), .A2(n6168), .ZN(n6176) );
  NAND2_X1 U6084 ( .A1(n5090), .A2(n4924), .ZN(n6815) );
  NAND2_X1 U6085 ( .A1(n6169), .A2(n5091), .ZN(n5090) );
  NAND2_X1 U6086 ( .A1(n6032), .A2(n5099), .ZN(n5096) );
  NAND2_X1 U6087 ( .A1(n5096), .A2(n5097), .ZN(n6163) );
  NAND2_X1 U6088 ( .A1(n5740), .A2(n5104), .ZN(n5743) );
  NAND2_X1 U6089 ( .A1(n5740), .A2(n5739), .ZN(n5741) );
  OAI211_X2 U6090 ( .C1(n6537), .C2(n7143), .A(n6333), .B(n5114), .ZN(n7658)
         );
  NAND2_X1 U6091 ( .A1(n6379), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n5114) );
  AND2_X2 U6092 ( .A1(n6348), .A2(n7139), .ZN(n6379) );
  AND2_X2 U6094 ( .A1(n7757), .A2(n10445), .ZN(n7759) );
  NOR2_X2 U6095 ( .A1(n7842), .A2(n7665), .ZN(n7757) );
  NAND2_X1 U6096 ( .A1(n8786), .A2(n5115), .ZN(n5120) );
  NAND2_X1 U6097 ( .A1(n8786), .A2(n6757), .ZN(n6804) );
  INV_X1 U6098 ( .A(n5120), .ZN(n8772) );
  NOR2_X2 U6099 ( .A1(n8993), .A2(n8858), .ZN(n8849) );
  NAND4_X2 U6100 ( .A1(n5524), .A2(n5468), .A3(n5127), .A4(n5383), .ZN(n5590)
         );
  NAND3_X1 U6101 ( .A1(n5524), .A2(n5468), .A3(n5127), .ZN(n5608) );
  NAND2_X1 U6102 ( .A1(n9880), .A2(n5131), .ZN(n5130) );
  OAI211_X1 U6103 ( .C1(n10395), .C2(n5136), .A(n9659), .B(n5134), .ZN(n6146)
         );
  INV_X1 U6104 ( .A(n10396), .ZN(n5135) );
  NAND2_X1 U6105 ( .A1(n6200), .A2(n10397), .ZN(n5137) );
  INV_X1 U6106 ( .A(n6199), .ZN(n5140) );
  INV_X1 U6107 ( .A(n6161), .ZN(n5143) );
  NAND2_X1 U6108 ( .A1(n5146), .A2(n5144), .ZN(n6267) );
  NAND2_X1 U6109 ( .A1(n4907), .A2(n9974), .ZN(n5149) );
  NOR2_X1 U6110 ( .A1(n9971), .A2(n6158), .ZN(n9949) );
  INV_X1 U6111 ( .A(n9971), .ZN(n5152) );
  AOI21_X1 U6112 ( .B1(n8104), .B2(n6150), .A(n5155), .ZN(n5154) );
  NAND2_X1 U6113 ( .A1(n6150), .A2(n8113), .ZN(n5156) );
  INV_X1 U6114 ( .A(n8104), .ZN(n5157) );
  NOR2_X4 U6115 ( .A1(n5590), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n5636) );
  NAND2_X1 U6116 ( .A1(n10349), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n5164) );
  NAND2_X1 U6117 ( .A1(n8912), .A2(n5185), .ZN(n5184) );
  NAND2_X1 U6118 ( .A1(n5184), .A2(n5182), .ZN(n6732) );
  NAND2_X1 U6119 ( .A1(n7987), .A2(n5193), .ZN(n5191) );
  NAND2_X1 U6120 ( .A1(n7788), .A2(n5201), .ZN(n5199) );
  NAND2_X1 U6121 ( .A1(n5199), .A2(n5197), .ZN(n8045) );
  AOI21_X1 U6122 ( .B1(n5201), .B2(n5203), .A(n5198), .ZN(n5197) );
  NAND2_X1 U6123 ( .A1(n7753), .A2(n5207), .ZN(n5206) );
  OAI21_X2 U6124 ( .B1(n6727), .B2(n5213), .A(n4891), .ZN(n8935) );
  NAND2_X1 U6125 ( .A1(n5219), .A2(n5217), .ZN(n5216) );
  INV_X1 U6126 ( .A(n5219), .ZN(n5218) );
  NAND2_X1 U6127 ( .A1(n5517), .A2(n5516), .ZN(n7613) );
  NAND2_X1 U6128 ( .A1(n5222), .A2(n5547), .ZN(n7743) );
  NAND3_X1 U6129 ( .A1(n5517), .A2(n5516), .A3(n4884), .ZN(n5222) );
  INV_X1 U6130 ( .A(n5232), .ZN(n9323) );
  NAND2_X1 U6131 ( .A1(n6233), .A2(n5234), .ZN(n5233) );
  NAND2_X1 U6132 ( .A1(n8381), .A2(n5241), .ZN(n5240) );
  OAI21_X1 U6133 ( .B1(n9367), .B2(n5252), .A(n5249), .ZN(n9412) );
  NAND2_X1 U6134 ( .A1(n9367), .A2(n5249), .ZN(n5248) );
  OAI21_X1 U6135 ( .B1(n8112), .B2(n5254), .A(n4867), .ZN(n8273) );
  NAND2_X2 U6136 ( .A1(n9422), .A2(n5258), .ZN(n5257) );
  INV_X1 U6137 ( .A(n5259), .ZN(n9350) );
  OAI21_X1 U6138 ( .B1(n7938), .B2(n5264), .A(n5263), .ZN(n8114) );
  NAND2_X1 U6139 ( .A1(n8580), .A2(n7776), .ZN(n9596) );
  NAND2_X1 U6140 ( .A1(n6113), .A2(n5269), .ZN(n5426) );
  NAND2_X1 U6141 ( .A1(n6113), .A2(n6115), .ZN(n5415) );
  INV_X1 U6142 ( .A(n5426), .ZN(n5428) );
  NAND2_X1 U6143 ( .A1(n9009), .A2(n5273), .ZN(n5272) );
  NAND2_X1 U6144 ( .A1(n7985), .A2(n5297), .ZN(n5296) );
  NAND2_X1 U6145 ( .A1(n8951), .A2(n5304), .ZN(n5303) );
  OAI21_X1 U6146 ( .B1(n8951), .B2(n5306), .A(n5304), .ZN(n8922) );
  AOI21_X1 U6147 ( .B1(n5304), .B2(n5306), .A(n5302), .ZN(n5301) );
  INV_X1 U6148 ( .A(n6545), .ZN(n5325) );
  NAND2_X2 U6149 ( .A1(n5328), .A2(n5326), .ZN(n5473) );
  NAND3_X1 U6150 ( .A1(n5327), .A2(P2_ADDR_REG_19__SCAN_IN), .A3(
        P1_ADDR_REG_19__SCAN_IN), .ZN(n5326) );
  INV_X1 U6151 ( .A(n8529), .ZN(n5331) );
  NAND2_X1 U6152 ( .A1(n5500), .A2(n5499), .ZN(n5531) );
  NAND2_X1 U6153 ( .A1(n5500), .A2(n5337), .ZN(n5336) );
  NAND3_X1 U6154 ( .A1(n5346), .A2(n5342), .A3(n5345), .ZN(n5344) );
  NAND2_X1 U6155 ( .A1(n5341), .A2(n5350), .ZN(n5345) );
  NAND3_X1 U6156 ( .A1(n8443), .A2(n8440), .A3(n5350), .ZN(n5346) );
  INV_X1 U6157 ( .A(n5350), .ZN(n8488) );
  INV_X1 U6158 ( .A(n8502), .ZN(n5349) );
  NAND2_X1 U6159 ( .A1(n5353), .A2(n5759), .ZN(n5782) );
  NAND2_X1 U6160 ( .A1(n5743), .A2(n5759), .ZN(n5744) );
  OAI21_X1 U6161 ( .B1(n8644), .B2(n5358), .A(n5357), .ZN(n8656) );
  NAND2_X1 U6162 ( .A1(n7126), .A2(n8520), .ZN(n5357) );
  INV_X1 U6163 ( .A(n5360), .ZN(n5359) );
  OAI21_X1 U6164 ( .B1(n7126), .B2(n7116), .A(n8520), .ZN(n5360) );
  NAND2_X1 U6165 ( .A1(n7686), .A2(n4873), .ZN(n5361) );
  INV_X1 U6166 ( .A(n6275), .ZN(n6276) );
  NAND2_X1 U6167 ( .A1(n6265), .A2(n6264), .ZN(n8596) );
  OR2_X1 U6168 ( .A1(n9481), .A2(n8382), .ZN(n6155) );
  OAI21_X1 U6169 ( .B1(n8596), .B2(n10504), .A(n6274), .ZN(n6275) );
  OR2_X1 U6170 ( .A1(n6262), .A2(n6261), .ZN(P1_U3355) );
  NAND2_X1 U6171 ( .A1(n9997), .A2(n10535), .ZN(n6284) );
  NAND2_X1 U6172 ( .A1(n8601), .A2(n6276), .ZN(n9997) );
  INV_X1 U6173 ( .A(n6272), .ZN(n8601) );
  NAND2_X1 U6174 ( .A1(n7209), .A2(n7037), .ZN(n10242) );
  OR2_X1 U6175 ( .A1(n7587), .A2(n5529), .ZN(n5793) );
  AND2_X1 U6176 ( .A1(n5446), .A2(n5381), .ZN(n5452) );
  NOR2_X1 U6177 ( .A1(n8134), .A2(n8139), .ZN(n8133) );
  NAND2_X1 U6178 ( .A1(n8616), .A2(n8615), .ZN(n8614) );
  XNOR2_X1 U6179 ( .A(n8526), .B(n8524), .ZN(n8616) );
  INV_X1 U6180 ( .A(n6083), .ZN(n6769) );
  AOI21_X1 U6181 ( .B1(n10392), .B2(n6083), .A(n5485), .ZN(n5487) );
  CLKBUF_X1 U6182 ( .A(n6340), .Z(n8699) );
  OR2_X1 U6183 ( .A1(n6744), .A2(n7380), .ZN(n6368) );
  OR2_X1 U6184 ( .A1(n6744), .A2(n6334), .ZN(n6339) );
  NAND3_X1 U6185 ( .A1(n6339), .A2(n6338), .A3(n6337), .ZN(n6340) );
  AND2_X1 U6186 ( .A1(n6336), .A2(n6335), .ZN(n6338) );
  MUX2_X1 U6187 ( .A(P1_IR_REG_0__SCAN_IN), .B(n10120), .S(n7043), .Z(n10385)
         );
  OAI22_X1 U6188 ( .A1(n5528), .A2(n7144), .B1(n7043), .B2(n7279), .ZN(n5406)
         );
  OAI22_X1 U6189 ( .A1(n5528), .A2(n5469), .B1(n7043), .B2(n7647), .ZN(n5470)
         );
  XNOR2_X1 U6190 ( .A(n5782), .B(n5781), .ZN(n7543) );
  NAND2_X1 U6191 ( .A1(n6723), .A2(n6890), .ZN(n7788) );
  OR2_X1 U6192 ( .A1(n5422), .A2(n5409), .ZN(n5412) );
  NAND2_X1 U6193 ( .A1(n5835), .A2(n5834), .ZN(n5855) );
  OR2_X1 U6194 ( .A1(n6302), .A2(n9294), .ZN(n6304) );
  OAI21_X1 U6195 ( .B1(n9996), .B2(n9985), .A(n6260), .ZN(n6261) );
  OAI211_X1 U6196 ( .C1(n5473), .C2(P1_DATAO_REG_0__SCAN_IN), .A(n5396), .B(
        SI_0_), .ZN(n5398) );
  NAND2_X1 U6197 ( .A1(n5473), .A2(n5395), .ZN(n5396) );
  OAI21_X1 U6198 ( .B1(n8458), .B2(n8459), .A(n6940), .ZN(n8913) );
  NAND2_X1 U6199 ( .A1(n7868), .A2(n9596), .ZN(n7869) );
  XNOR2_X2 U6200 ( .A(n6331), .B(P2_IR_REG_1__SCAN_IN), .ZN(n10349) );
  INV_X1 U6201 ( .A(n8400), .ZN(n7031) );
  NAND2_X1 U6202 ( .A1(n7251), .A2(n7250), .ZN(n10551) );
  INV_X2 U6203 ( .A(n10551), .ZN(n10553) );
  NAND2_X1 U6204 ( .A1(n7250), .A2(n7224), .ZN(n10554) );
  INV_X2 U6205 ( .A(n10554), .ZN(n10557) );
  AND2_X1 U6206 ( .A1(n9820), .A2(n9394), .ZN(n5366) );
  OR4_X1 U6207 ( .A1(n7033), .A2(n8512), .A3(n7032), .A4(n8675), .ZN(n5368) );
  XOR2_X1 U6208 ( .A(n6854), .B(n10461), .Z(n5369) );
  OR2_X1 U6209 ( .A1(n9716), .A2(n4989), .ZN(n5370) );
  NOR2_X1 U6210 ( .A1(n5897), .A2(n5896), .ZN(n5372) );
  AND4_X1 U6211 ( .A1(n6706), .A2(n6296), .A3(n6678), .A4(n6670), .ZN(n5374)
         );
  NAND2_X1 U6212 ( .A1(n7933), .A2(n10376), .ZN(n9940) );
  OR2_X1 U6213 ( .A1(n6384), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n5375) );
  AND2_X2 U6214 ( .A1(n7372), .A2(n7041), .ZN(P2_U3966) );
  AND2_X1 U6215 ( .A1(n5411), .A2(n5390), .ZN(n5376) );
  INV_X1 U6216 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n6434) );
  NAND2_X1 U6217 ( .A1(n6225), .A2(n6224), .ZN(n5377) );
  OR2_X1 U6218 ( .A1(n8964), .A2(n8952), .ZN(n5378) );
  INV_X1 U6219 ( .A(n9267), .ZN(n6750) );
  INV_X1 U6220 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n6184) );
  INV_X1 U6221 ( .A(n9759), .ZN(n9775) );
  OR2_X1 U6222 ( .A1(n10003), .A2(n9785), .ZN(n5379) );
  OR2_X1 U6223 ( .A1(n8969), .A2(n8952), .ZN(n5380) );
  INV_X1 U6224 ( .A(n9664), .ZN(n6151) );
  INV_X1 U6225 ( .A(n10401), .ZN(n6266) );
  OR2_X1 U6226 ( .A1(n7209), .A2(n10250), .ZN(n5381) );
  INV_X1 U6227 ( .A(n9413), .ZN(n9438) );
  AND2_X1 U6228 ( .A1(n6128), .A2(n6118), .ZN(n9413) );
  AND2_X1 U6229 ( .A1(n6878), .A2(n7767), .ZN(n5382) );
  NAND2_X1 U6230 ( .A1(n5830), .A2(n5831), .ZN(n9423) );
  INV_X1 U6231 ( .A(n7805), .ZN(n6442) );
  INV_X1 U6232 ( .A(n8419), .ZN(n6927) );
  INV_X1 U6233 ( .A(n6721), .ZN(n6874) );
  INV_X1 U6234 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n6292) );
  INV_X1 U6236 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n5390) );
  INV_X1 U6237 ( .A(n6222), .ZN(n6219) );
  INV_X1 U6238 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5421) );
  INV_X1 U6239 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n6551) );
  AND2_X1 U6240 ( .A1(n8828), .A2(n8826), .ZN(n6734) );
  INV_X1 U6241 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n6287) );
  NAND2_X1 U6242 ( .A1(n8590), .A2(n5454), .ZN(n5482) );
  OR2_X1 U6243 ( .A1(n9998), .A2(n9704), .ZN(n6250) );
  INV_X1 U6244 ( .A(SI_29_), .ZN(n9125) );
  INV_X1 U6245 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n6522) );
  INV_X1 U6246 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n6495) );
  INV_X1 U6247 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n6596) );
  NOR2_X1 U6248 ( .A1(n6563), .A2(n8444), .ZN(n6562) );
  AND2_X1 U6249 ( .A1(n6448), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n6466) );
  INV_X1 U6250 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n5668) );
  INV_X1 U6251 ( .A(n9653), .ZN(n6213) );
  OR2_X1 U6252 ( .A1(n6117), .A2(n6124), .ZN(n6201) );
  INV_X1 U6253 ( .A(SI_21_), .ZN(n9144) );
  NOR2_X1 U6254 ( .A1(n6637), .A2(n9114), .ZN(n6657) );
  AND2_X1 U6255 ( .A1(n7048), .A2(n7047), .ZN(n7049) );
  OR2_X1 U6256 ( .A1(n6619), .A2(n8638), .ZN(n6629) );
  AND2_X1 U6257 ( .A1(n6321), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6606) );
  OR2_X1 U6258 ( .A1(n6629), .A2(n9197), .ZN(n6637) );
  AND2_X1 U6259 ( .A1(n8993), .A2(n8864), .ZN(n6626) );
  NAND2_X1 U6260 ( .A1(n9257), .A2(n8427), .ZN(n6928) );
  INV_X1 U6261 ( .A(n8049), .ZN(n6457) );
  OR2_X1 U6262 ( .A1(n6435), .A2(n6434), .ZN(n6450) );
  INV_X1 U6263 ( .A(n7220), .ZN(n6711) );
  INV_X2 U6264 ( .A(n6534), .ZN(n6834) );
  OR2_X1 U6265 ( .A1(n10545), .A2(n8008), .ZN(n7220) );
  INV_X1 U6266 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n6672) );
  OR2_X1 U6267 ( .A1(n6491), .A2(n6490), .ZN(n6503) );
  INV_X1 U6268 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n5794) );
  AND2_X1 U6269 ( .A1(n5726), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5748) );
  INV_X1 U6270 ( .A(n9841), .ZN(n6241) );
  INV_X1 U6271 ( .A(n9667), .ZN(n9470) );
  INV_X1 U6272 ( .A(n9650), .ZN(n6190) );
  NAND2_X1 U6273 ( .A1(n6247), .A2(n5379), .ZN(n6249) );
  AND2_X1 U6274 ( .A1(n6825), .A2(n6180), .ZN(n6181) );
  INV_X1 U6275 ( .A(n6657), .ZN(n6655) );
  NOR2_X1 U6276 ( .A1(n7057), .A2(n7058), .ZN(n7299) );
  INV_X1 U6277 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n9114) );
  AND2_X1 U6278 ( .A1(n6637), .A2(n6630), .ZN(n8816) );
  AND4_X1 U6279 ( .A1(n6501), .A2(n6500), .A3(n6499), .A4(n6498), .ZN(n8211)
         );
  AND2_X1 U6280 ( .A1(n7221), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7255) );
  INV_X1 U6281 ( .A(n8873), .ZN(n8891) );
  INV_X1 U6282 ( .A(n8133), .ZN(n8237) );
  OR2_X1 U6284 ( .A1(n6348), .A2(n6332), .ZN(n6333) );
  INV_X1 U6285 ( .A(n8128), .ZN(n8132) );
  OR2_X1 U6286 ( .A1(n7371), .A2(n6741), .ZN(n8675) );
  OR2_X1 U6287 ( .A1(n7130), .A2(n7124), .ZN(n10536) );
  AND3_X1 U6288 ( .A1(n7221), .A2(P2_STATE_REG_SCAN_IN), .A3(n7220), .ZN(n7222) );
  OR3_X1 U6289 ( .A1(n5796), .A2(n5795), .A3(n5794), .ZN(n5820) );
  NAND2_X1 U6290 ( .A1(n6773), .A2(n9413), .ZN(n6774) );
  AND2_X1 U6291 ( .A1(n9414), .A2(n9410), .ZN(n6067) );
  NOR2_X1 U6292 ( .A1(n5820), .A2(n8082), .ZN(n5840) );
  AND3_X1 U6293 ( .A1(n6195), .A2(n6194), .A3(n6193), .ZN(n9618) );
  INV_X1 U6294 ( .A(n10008), .ZN(n9792) );
  AND2_X1 U6295 ( .A1(n9550), .A2(n9533), .ZN(n9668) );
  INV_X1 U6296 ( .A(n10522), .ZN(n10386) );
  INV_X1 U6297 ( .A(n10520), .ZN(n10502) );
  NAND2_X1 U6298 ( .A1(n6130), .A2(n6196), .ZN(n9975) );
  INV_X1 U6299 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n9084) );
  AND2_X1 U6300 ( .A1(n7132), .A2(n7131), .ZN(n8680) );
  INV_X1 U6301 ( .A(n7034), .ZN(n7035) );
  AND2_X1 U6302 ( .A1(n6644), .A2(n6643), .ZN(n8627) );
  AND2_X1 U6303 ( .A1(n7307), .A2(n7306), .ZN(n8741) );
  INV_X1 U6304 ( .A(n10353), .ZN(n10333) );
  INV_X1 U6305 ( .A(n10549), .ZN(n8773) );
  AND2_X1 U6306 ( .A1(n6986), .A2(n8778), .ZN(n8795) );
  INV_X1 U6307 ( .A(n6936), .ZN(n8459) );
  INV_X1 U6308 ( .A(n8675), .ZN(n8915) );
  INV_X1 U6309 ( .A(n8952), .ZN(n8933) );
  NOR2_X1 U6310 ( .A1(n7122), .A2(n7121), .ZN(n7251) );
  AND2_X1 U6311 ( .A1(n8051), .A2(n10510), .ZN(n9271) );
  INV_X1 U6312 ( .A(n9271), .ZN(n10541) );
  NAND2_X1 U6313 ( .A1(n10328), .A2(n6687), .ZN(n10154) );
  AND2_X1 U6314 ( .A1(n7139), .A2(P2_U3152), .ZN(n9297) );
  NAND2_X1 U6315 ( .A1(n6783), .A2(n6782), .ZN(n6784) );
  AOI21_X1 U6316 ( .B1(n9718), .B2(n6083), .A(n5458), .ZN(n7461) );
  INV_X1 U6317 ( .A(n9430), .ZN(n9416) );
  AND2_X1 U6318 ( .A1(n6138), .A2(n6137), .ZN(n9703) );
  AND2_X1 U6319 ( .A1(n5986), .A2(n5985), .ZN(n9394) );
  AND2_X1 U6320 ( .A1(n5891), .A2(n5890), .ZN(n9907) );
  NAND2_X1 U6321 ( .A1(n5548), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n5467) );
  INV_X1 U6322 ( .A(n10298), .ZN(n10318) );
  INV_X1 U6323 ( .A(n9736), .ZN(n10313) );
  AND2_X1 U6324 ( .A1(n7211), .A2(n6130), .ZN(n10312) );
  OAI21_X1 U6325 ( .B1(n8596), .B2(n10401), .A(n6271), .ZN(n6272) );
  INV_X1 U6326 ( .A(n9882), .ZN(n9875) );
  INV_X1 U6327 ( .A(n9977), .ZN(n10393) );
  NOR2_X1 U6328 ( .A1(n10504), .A2(n9591), .ZN(n6278) );
  NAND2_X1 U6329 ( .A1(n8515), .A2(n9685), .ZN(n7364) );
  OR2_X1 U6330 ( .A1(n9449), .A2(n9622), .ZN(n10504) );
  AND2_X1 U6331 ( .A1(n10240), .A2(n6280), .ZN(n7775) );
  AOI21_X1 U6332 ( .B1(n10121), .B2(n10241), .A(n6102), .ZN(n6277) );
  INV_X1 U6333 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n6100) );
  AND2_X1 U6334 ( .A1(n5639), .A2(n5664), .ZN(n7321) );
  INV_X1 U6335 ( .A(n8741), .ZN(n10352) );
  NAND2_X1 U6336 ( .A1(n8680), .A2(n8915), .ZN(n8660) );
  NAND2_X1 U6337 ( .A1(n7132), .A2(n7125), .ZN(n8669) );
  AND3_X1 U6338 ( .A1(n6799), .A2(n6798), .A3(n6797), .ZN(n7174) );
  INV_X1 U6339 ( .A(P2_U3966), .ZN(n8688) );
  NAND2_X1 U6340 ( .A1(n7377), .A2(n7376), .ZN(n10353) );
  INV_X1 U6341 ( .A(n10364), .ZN(n10335) );
  AND2_X1 U6342 ( .A1(n8919), .A2(n8918), .ZN(n9245) );
  AND3_X1 U6343 ( .A1(n7838), .A2(n7837), .A3(n7836), .ZN(n10432) );
  NAND2_X1 U6344 ( .A1(n10155), .A2(n10154), .ZN(n10329) );
  NOR2_X1 U6345 ( .A1(n7040), .A2(P2_U3152), .ZN(n10331) );
  INV_X1 U6346 ( .A(n8312), .ZN(n8038) );
  INV_X1 U6347 ( .A(n6143), .ZN(n6144) );
  AOI21_X1 U6348 ( .B1(n6786), .B2(n6785), .A(n6784), .ZN(n6787) );
  AND2_X1 U6349 ( .A1(n6121), .A2(n10376), .ZN(n9409) );
  INV_X1 U6350 ( .A(n9394), .ZN(n9831) );
  INV_X1 U6351 ( .A(n9907), .ZN(n9884) );
  OR2_X1 U6352 ( .A1(P1_U3083), .A2(n7210), .ZN(n9736) );
  OR2_X1 U6353 ( .A1(n10274), .A2(n6130), .ZN(n10298) );
  OR3_X1 U6354 ( .A1(n10116), .A2(n10245), .A3(n10247), .ZN(n10269) );
  OR2_X1 U6355 ( .A1(n10419), .A2(n6253), .ZN(n9985) );
  AND2_X2 U6356 ( .A1(n7775), .A2(n10103), .ZN(n10531) );
  OR2_X1 U6357 ( .A1(n10535), .A2(n6282), .ZN(n6283) );
  OR2_X1 U6358 ( .A1(n10077), .A2(n10076), .ZN(n10101) );
  INV_X1 U6359 ( .A(n10535), .ZN(n10532) );
  AND2_X2 U6360 ( .A1(n7775), .A2(n6281), .ZN(n10535) );
  INV_X1 U6361 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n8603) );
  XNOR2_X1 U6362 ( .A(n5416), .B(n5271), .ZN(n8404) );
  INV_X1 U6363 ( .A(n8077), .ZN(n7712) );
  NOR2_X1 U6364 ( .A1(n10212), .A2(n10211), .ZN(n10214) );
  NAND2_X1 U6365 ( .A1(n5378), .A2(n6810), .ZN(P2_U3267) );
  INV_X1 U6366 ( .A(n9719), .ZN(P1_U4006) );
  NAND2_X1 U6367 ( .A1(n6284), .A2(n6283), .ZN(P1_U3519) );
  NOR2_X1 U6368 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n5389) );
  NOR2_X1 U6369 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n5388) );
  NOR2_X1 U6370 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .ZN(
        n5387) );
  NOR2_X1 U6371 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n5386) );
  NAND2_X1 U6372 ( .A1(n5422), .A2(n5376), .ZN(n5391) );
  NAND2_X1 U6373 ( .A1(P1_IR_REG_27__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), 
        .ZN(n5392) );
  NAND2_X1 U6374 ( .A1(n5394), .A2(n5392), .ZN(n5393) );
  XNOR2_X2 U6375 ( .A(n5394), .B(n5427), .ZN(n9695) );
  INV_X1 U6376 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5395) );
  INV_X1 U6377 ( .A(n5398), .ZN(n5397) );
  NAND2_X1 U6378 ( .A1(n5397), .A2(SI_1_), .ZN(n5471) );
  INV_X1 U6379 ( .A(SI_1_), .ZN(n9172) );
  NAND2_X1 U6380 ( .A1(n5398), .A2(n9172), .ZN(n5399) );
  MUX2_X1 U6381 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .S(n5473), .Z(n5401) );
  INV_X1 U6382 ( .A(n5400), .ZN(n5403) );
  INV_X1 U6383 ( .A(n5401), .ZN(n5402) );
  NAND2_X1 U6384 ( .A1(n5403), .A2(n5402), .ZN(n5404) );
  NAND2_X1 U6385 ( .A1(n5472), .A2(n5404), .ZN(n7143) );
  NAND2_X2 U6386 ( .A1(n7043), .A2(n7138), .ZN(n5528) );
  INV_X1 U6387 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n7144) );
  NAND2_X1 U6388 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5405) );
  XNOR2_X1 U6389 ( .A(n5405), .B(P1_IR_REG_1__SCAN_IN), .ZN(n7201) );
  INV_X1 U6390 ( .A(n7201), .ZN(n7279) );
  NAND2_X4 U6391 ( .A1(n5408), .A2(n5407), .ZN(n10408) );
  NAND2_X1 U6392 ( .A1(n5415), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5416) );
  NOR2_X1 U6393 ( .A1(n6094), .A2(n8404), .ZN(n5417) );
  NAND2_X1 U6394 ( .A1(n4883), .A2(P1_IR_REG_21__SCAN_IN), .ZN(n5419) );
  NAND2_X1 U6395 ( .A1(n10408), .A2(n5454), .ZN(n5437) );
  INV_X1 U6396 ( .A(n5426), .ZN(n5424) );
  AOI21_X1 U6397 ( .B1(n5428), .B2(n5427), .A(n5409), .ZN(n5429) );
  INV_X1 U6398 ( .A(n5429), .ZN(n5430) );
  NAND2_X1 U6399 ( .A1(n5548), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n5434) );
  NAND2_X1 U6400 ( .A1(n5644), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n5432) );
  NOR2_X2 U6401 ( .A1(n4996), .A2(n8604), .ZN(n5519) );
  NAND2_X1 U6402 ( .A1(n5519), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5431) );
  NAND4_X2 U6403 ( .A1(n5434), .A2(n5433), .A3(n5432), .A4(n5431), .ZN(n9718)
         );
  INV_X1 U6404 ( .A(n5443), .ZN(n7734) );
  NAND2_X1 U6405 ( .A1(n9718), .A2(n5435), .ZN(n5436) );
  NAND2_X1 U6406 ( .A1(n5437), .A2(n5436), .ZN(n5444) );
  NAND2_X1 U6407 ( .A1(n5440), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5441) );
  XNOR2_X2 U6408 ( .A(n5441), .B(P1_IR_REG_19__SCAN_IN), .ZN(n10411) );
  OAI22_X1 U6409 ( .A1(n8515), .A2(n10411), .B1(n9693), .B2(n9685), .ZN(n5442)
         );
  XNOR2_X1 U6410 ( .A(n5444), .B(n6081), .ZN(n5460) );
  NAND2_X1 U6411 ( .A1(n7142), .A2(SI_0_), .ZN(n5445) );
  XNOR2_X1 U6412 ( .A(n5445), .B(P2_DATAO_REG_0__SCAN_IN), .ZN(n10120) );
  NAND2_X1 U6413 ( .A1(n10385), .A2(n5454), .ZN(n5446) );
  INV_X1 U6414 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n10250) );
  NAND2_X1 U6415 ( .A1(n5644), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5450) );
  NAND2_X1 U6416 ( .A1(n5864), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5449) );
  NAND2_X1 U6417 ( .A1(n5548), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n5448) );
  NAND2_X1 U6418 ( .A1(n5519), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n5447) );
  NAND4_X1 U6419 ( .A1(n5450), .A2(n5449), .A3(n5448), .A4(n5447), .ZN(n6205)
         );
  NAND2_X1 U6420 ( .A1(n6205), .A2(n5435), .ZN(n5451) );
  NAND2_X1 U6421 ( .A1(n5452), .A2(n5451), .ZN(n7335) );
  INV_X1 U6422 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n10253) );
  NAND2_X1 U6423 ( .A1(n8515), .A2(n6124), .ZN(n5453) );
  NAND2_X1 U6424 ( .A1(n6205), .A2(n6083), .ZN(n5456) );
  NAND2_X1 U6425 ( .A1(n10385), .A2(n4856), .ZN(n5455) );
  OAI211_X1 U6426 ( .C1(n7209), .C2(n10253), .A(n5456), .B(n5455), .ZN(n7334)
         );
  NAND2_X1 U6427 ( .A1(n7335), .A2(n7334), .ZN(n5457) );
  OAI21_X1 U6428 ( .B1(n7335), .B2(n6081), .A(n5457), .ZN(n5459) );
  NAND2_X1 U6429 ( .A1(n5460), .A2(n5459), .ZN(n7459) );
  AND2_X1 U6430 ( .A1(n10408), .A2(n5435), .ZN(n5458) );
  NAND2_X1 U6431 ( .A1(n7459), .A2(n7461), .ZN(n5463) );
  INV_X1 U6432 ( .A(n5459), .ZN(n5462) );
  INV_X1 U6433 ( .A(n5460), .ZN(n5461) );
  NAND2_X1 U6434 ( .A1(n5462), .A2(n5461), .ZN(n7460) );
  NAND2_X1 U6435 ( .A1(n5864), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5466) );
  NAND2_X1 U6436 ( .A1(n5644), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5465) );
  NAND2_X1 U6437 ( .A1(n5519), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5464) );
  NAND4_X2 U6438 ( .A1(n5467), .A2(n5466), .A3(n5465), .A4(n5464), .ZN(n10392)
         );
  NAND2_X1 U6439 ( .A1(n10392), .A2(n4856), .ZN(n5483) );
  INV_X1 U6440 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n5469) );
  OR2_X1 U6441 ( .A1(n5468), .A2(n5409), .ZN(n5526) );
  NAND2_X1 U6442 ( .A1(n5526), .A2(n5126), .ZN(n5491) );
  OAI21_X1 U6443 ( .B1(n5526), .B2(n5126), .A(n5491), .ZN(n7647) );
  NAND2_X1 U6444 ( .A1(n5472), .A2(n5471), .ZN(n5478) );
  INV_X1 U6445 ( .A(n5478), .ZN(n5475) );
  MUX2_X1 U6446 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .S(n5473), .Z(n5474) );
  NAND2_X1 U6447 ( .A1(n5474), .A2(SI_2_), .ZN(n5494) );
  OAI21_X1 U6448 ( .B1(n5474), .B2(SI_2_), .A(n5494), .ZN(n5476) );
  NAND2_X1 U6449 ( .A1(n5475), .A2(n5476), .ZN(n5479) );
  INV_X1 U6450 ( .A(n5476), .ZN(n5477) );
  NAND2_X1 U6451 ( .A1(n5478), .A2(n5477), .ZN(n5495) );
  NAND2_X1 U6452 ( .A1(n5479), .A2(n5495), .ZN(n7149) );
  NAND2_X1 U6453 ( .A1(n5483), .A2(n5482), .ZN(n5484) );
  XNOR2_X1 U6454 ( .A(n5484), .B(n6081), .ZN(n5486) );
  AND2_X1 U6455 ( .A1(n8590), .A2(n5435), .ZN(n5485) );
  XNOR2_X1 U6456 ( .A(n5486), .B(n5487), .ZN(n8587) );
  NAND2_X1 U6457 ( .A1(n8588), .A2(n8587), .ZN(n5490) );
  INV_X1 U6458 ( .A(n5486), .ZN(n5488) );
  NAND2_X1 U6459 ( .A1(n5488), .A2(n5487), .ZN(n5489) );
  NAND2_X1 U6460 ( .A1(n5490), .A2(n5489), .ZN(n7589) );
  NAND2_X1 U6461 ( .A1(n5491), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5493) );
  INV_X1 U6462 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n5492) );
  NAND2_X1 U6463 ( .A1(n5495), .A2(n5494), .ZN(n5500) );
  MUX2_X1 U6464 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .S(n5473), .Z(n5496) );
  NAND2_X1 U6465 ( .A1(n5496), .A2(SI_3_), .ZN(n5530) );
  INV_X1 U6466 ( .A(n5496), .ZN(n5497) );
  INV_X1 U6467 ( .A(SI_3_), .ZN(n9056) );
  NAND2_X1 U6468 ( .A1(n5497), .A2(n9056), .ZN(n5498) );
  AND2_X1 U6469 ( .A1(n5530), .A2(n5498), .ZN(n5499) );
  OR2_X1 U6470 ( .A1(n5500), .A2(n5499), .ZN(n5501) );
  NAND2_X1 U6471 ( .A1(n5531), .A2(n5501), .ZN(n7146) );
  OR2_X1 U6472 ( .A1(n5529), .A2(n7146), .ZN(n5504) );
  INV_X1 U6473 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n5502) );
  OR2_X1 U6474 ( .A1(n5528), .A2(n5502), .ZN(n5503) );
  OAI211_X1 U6475 ( .C1(n7043), .C2(n4852), .A(n5504), .B(n5503), .ZN(n7776)
         );
  INV_X2 U6476 ( .A(n5987), .ZN(n6761) );
  NAND2_X1 U6477 ( .A1(n7776), .A2(n6761), .ZN(n5510) );
  INV_X1 U6478 ( .A(n5864), .ZN(n5671) );
  NAND2_X1 U6479 ( .A1(n4851), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n5508) );
  INV_X1 U6480 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n7736) );
  NAND2_X1 U6481 ( .A1(n5548), .A2(n7736), .ZN(n5507) );
  NAND2_X1 U6482 ( .A1(n5644), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5506) );
  NAND2_X1 U6483 ( .A1(n4854), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5505) );
  NAND2_X1 U6484 ( .A1(n9717), .A2(n5435), .ZN(n5509) );
  NAND2_X1 U6485 ( .A1(n5510), .A2(n5509), .ZN(n5511) );
  XNOR2_X1 U6486 ( .A(n5511), .B(n6081), .ZN(n5513) );
  AND2_X1 U6487 ( .A1(n7776), .A2(n4856), .ZN(n5512) );
  AOI21_X1 U6488 ( .B1(n9717), .B2(n6083), .A(n5512), .ZN(n5514) );
  XNOR2_X1 U6489 ( .A(n5513), .B(n5514), .ZN(n7590) );
  NAND2_X1 U6490 ( .A1(n7589), .A2(n7590), .ZN(n5517) );
  INV_X1 U6491 ( .A(n5513), .ZN(n5515) );
  NAND2_X1 U6492 ( .A1(n5515), .A2(n5514), .ZN(n5516) );
  NAND2_X1 U6493 ( .A1(n4851), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5523) );
  NOR2_X1 U6494 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n5518) );
  NOR2_X1 U6495 ( .A1(n5549), .A2(n5518), .ZN(n7875) );
  NAND2_X1 U6496 ( .A1(n4855), .A2(n7875), .ZN(n5522) );
  NAND2_X1 U6497 ( .A1(n8561), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5521) );
  NAND2_X1 U6498 ( .A1(n4854), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n5520) );
  NAND2_X1 U6499 ( .A1(n9716), .A2(n6062), .ZN(n5542) );
  OR2_X1 U6500 ( .A1(n5524), .A2(n5409), .ZN(n5525) );
  NAND2_X1 U6501 ( .A1(n5526), .A2(n5525), .ZN(n5554) );
  INV_X1 U6502 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5527) );
  XNOR2_X1 U6503 ( .A(n5554), .B(n5527), .ZN(n7204) );
  INV_X1 U6504 ( .A(n7204), .ZN(n7636) );
  INV_X1 U6505 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n7148) );
  OR2_X1 U6506 ( .A1(n5528), .A2(n7148), .ZN(n5540) );
  MUX2_X1 U6507 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .S(n5473), .Z(n5532) );
  NAND2_X1 U6508 ( .A1(n5532), .A2(SI_4_), .ZN(n5556) );
  INV_X1 U6509 ( .A(n5532), .ZN(n5534) );
  INV_X1 U6510 ( .A(SI_4_), .ZN(n5533) );
  NAND2_X1 U6511 ( .A1(n5534), .A2(n5533), .ZN(n5535) );
  AND2_X1 U6512 ( .A1(n5556), .A2(n5535), .ZN(n5536) );
  OR2_X1 U6513 ( .A1(n5537), .A2(n5536), .ZN(n5538) );
  NAND2_X1 U6514 ( .A1(n5557), .A2(n5538), .ZN(n7147) );
  OR2_X1 U6515 ( .A1(n5529), .A2(n7147), .ZN(n5539) );
  OAI211_X1 U6516 ( .C1(n7636), .C2(n7043), .A(n5540), .B(n5539), .ZN(n7876)
         );
  NAND2_X1 U6517 ( .A1(n7876), .A2(n6761), .ZN(n5541) );
  NAND2_X1 U6518 ( .A1(n5542), .A2(n5541), .ZN(n5543) );
  AND2_X1 U6519 ( .A1(n7876), .A2(n6062), .ZN(n5544) );
  INV_X1 U6520 ( .A(n7611), .ZN(n5546) );
  INV_X1 U6521 ( .A(n7610), .ZN(n5545) );
  NAND2_X1 U6522 ( .A1(n5546), .A2(n5545), .ZN(n5547) );
  NAND2_X1 U6523 ( .A1(n4851), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5553) );
  NAND2_X1 U6524 ( .A1(n5549), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n5603) );
  OAI21_X1 U6525 ( .B1(n5549), .B2(P1_REG3_REG_5__SCAN_IN), .A(n5603), .ZN(
        n7747) );
  INV_X1 U6526 ( .A(n7747), .ZN(n7934) );
  NAND2_X1 U6527 ( .A1(n4855), .A2(n7934), .ZN(n5552) );
  NAND2_X1 U6528 ( .A1(n5644), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n5551) );
  NAND2_X1 U6529 ( .A1(n4854), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n5550) );
  NAND4_X1 U6530 ( .A1(n5553), .A2(n5552), .A3(n5551), .A4(n5550), .ZN(n9715)
         );
  NAND2_X1 U6531 ( .A1(n9715), .A2(n6062), .ZN(n5567) );
  OAI21_X1 U6532 ( .B1(n5554), .B2(P1_IR_REG_4__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5555) );
  XNOR2_X1 U6533 ( .A(n5555), .B(P1_IR_REG_5__SCAN_IN), .ZN(n10311) );
  INV_X1 U6534 ( .A(n10311), .ZN(n7152) );
  MUX2_X1 U6535 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n7139), .Z(n5558) );
  NAND2_X1 U6536 ( .A1(n5558), .A2(SI_5_), .ZN(n5576) );
  INV_X1 U6537 ( .A(n5558), .ZN(n5559) );
  NAND2_X1 U6538 ( .A1(n5559), .A2(n9165), .ZN(n5560) );
  AND2_X1 U6539 ( .A1(n5576), .A2(n5560), .ZN(n5561) );
  NAND2_X1 U6540 ( .A1(n5562), .A2(n5561), .ZN(n5577) );
  OR2_X1 U6541 ( .A1(n5562), .A2(n5561), .ZN(n5563) );
  NAND2_X1 U6542 ( .A1(n5577), .A2(n5563), .ZN(n7153) );
  OR2_X1 U6543 ( .A1(n5529), .A2(n7153), .ZN(n5565) );
  INV_X1 U6544 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n7154) );
  OR2_X1 U6545 ( .A1(n5528), .A2(n7154), .ZN(n5564) );
  OAI211_X1 U6546 ( .C1(n7043), .C2(n7152), .A(n5565), .B(n5564), .ZN(n8065)
         );
  NAND2_X1 U6547 ( .A1(n8065), .A2(n6761), .ZN(n5566) );
  NAND2_X1 U6548 ( .A1(n5567), .A2(n5566), .ZN(n5568) );
  XNOR2_X1 U6549 ( .A(n5568), .B(n6081), .ZN(n7744) );
  NAND2_X1 U6550 ( .A1(n7743), .A2(n7744), .ZN(n7907) );
  INV_X1 U6551 ( .A(n5603), .ZN(n5569) );
  AOI21_X1 U6552 ( .B1(n5569), .B2(P1_REG3_REG_6__SCAN_IN), .A(
        P1_REG3_REG_7__SCAN_IN), .ZN(n5571) );
  NAND2_X1 U6553 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_REG3_REG_7__SCAN_IN), 
        .ZN(n5570) );
  NOR2_X1 U6554 ( .A1(n5603), .A2(n5570), .ZN(n5642) );
  OR2_X1 U6555 ( .A1(n5571), .A2(n5642), .ZN(n7978) );
  INV_X1 U6556 ( .A(n7978), .ZN(n8109) );
  NAND2_X1 U6557 ( .A1(n4855), .A2(n8109), .ZN(n5575) );
  NAND2_X1 U6558 ( .A1(n4851), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5574) );
  NAND2_X1 U6559 ( .A1(n8561), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5573) );
  NAND2_X1 U6560 ( .A1(n4854), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n5572) );
  NAND4_X1 U6561 ( .A1(n5575), .A2(n5574), .A3(n5573), .A4(n5572), .ZN(n9713)
         );
  NAND2_X1 U6562 ( .A1(n9713), .A2(n6767), .ZN(n5595) );
  NAND2_X1 U6563 ( .A1(n5577), .A2(n5576), .ZN(n5612) );
  MUX2_X1 U6564 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n7139), .Z(n5578) );
  NAND2_X1 U6565 ( .A1(n5578), .A2(SI_6_), .ZN(n5582) );
  INV_X1 U6566 ( .A(n5578), .ZN(n5580) );
  INV_X1 U6567 ( .A(SI_6_), .ZN(n5579) );
  NAND2_X1 U6568 ( .A1(n5580), .A2(n5579), .ZN(n5581) );
  AND2_X1 U6569 ( .A1(n5582), .A2(n5581), .ZN(n5611) );
  MUX2_X1 U6570 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n7139), .Z(n5583) );
  NAND2_X1 U6571 ( .A1(n5583), .A2(SI_7_), .ZN(n5634) );
  INV_X1 U6572 ( .A(n5583), .ZN(n5585) );
  INV_X1 U6573 ( .A(SI_7_), .ZN(n5584) );
  NAND2_X1 U6574 ( .A1(n5585), .A2(n5584), .ZN(n5586) );
  AND2_X1 U6575 ( .A1(n5634), .A2(n5586), .ZN(n5587) );
  OR2_X1 U6576 ( .A1(n5588), .A2(n5587), .ZN(n5589) );
  NAND2_X1 U6577 ( .A1(n5635), .A2(n5589), .ZN(n7159) );
  OR2_X1 U6578 ( .A1(n7159), .A2(n5529), .ZN(n5593) );
  NAND2_X1 U6579 ( .A1(n5590), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5591) );
  XNOR2_X1 U6580 ( .A(n5591), .B(P1_IR_REG_7__SCAN_IN), .ZN(n7246) );
  AOI22_X1 U6581 ( .A1(n6072), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n10246), .B2(
        n7246), .ZN(n5592) );
  NAND2_X1 U6582 ( .A1(n8162), .A2(n6761), .ZN(n5594) );
  NAND2_X1 U6583 ( .A1(n5595), .A2(n5594), .ZN(n5596) );
  XNOR2_X1 U6584 ( .A(n5596), .B(n6765), .ZN(n5601) );
  NAND2_X1 U6585 ( .A1(n9713), .A2(n6083), .ZN(n5598) );
  NAND2_X1 U6586 ( .A1(n8162), .A2(n6767), .ZN(n5597) );
  NAND2_X1 U6587 ( .A1(n5598), .A2(n5597), .ZN(n5600) );
  INV_X1 U6588 ( .A(n5600), .ZN(n5599) );
  NAND2_X1 U6589 ( .A1(n5601), .A2(n5599), .ZN(n5631) );
  INV_X1 U6590 ( .A(n5631), .ZN(n5602) );
  XNOR2_X1 U6591 ( .A(n5601), .B(n5600), .ZN(n7976) );
  NOR2_X1 U6592 ( .A1(n5602), .A2(n7976), .ZN(n5633) );
  INV_X1 U6593 ( .A(n5633), .ZN(n5623) );
  XNOR2_X1 U6594 ( .A(n5603), .B(P1_REG3_REG_6__SCAN_IN), .ZN(n7951) );
  NAND2_X1 U6595 ( .A1(n4855), .A2(n7951), .ZN(n5607) );
  NAND2_X1 U6596 ( .A1(n4851), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n5606) );
  NAND2_X1 U6597 ( .A1(n8561), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5605) );
  NAND2_X1 U6598 ( .A1(n4854), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n5604) );
  NAND4_X1 U6599 ( .A1(n5607), .A2(n5606), .A3(n5605), .A4(n5604), .ZN(n9714)
         );
  NAND2_X1 U6600 ( .A1(n9714), .A2(n6062), .ZN(n5618) );
  NAND2_X1 U6601 ( .A1(n5608), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5609) );
  XNOR2_X1 U6602 ( .A(n5609), .B(P1_IR_REG_6__SCAN_IN), .ZN(n10256) );
  INV_X1 U6603 ( .A(n10256), .ZN(n7157) );
  INV_X1 U6604 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n5610) );
  OR2_X1 U6605 ( .A1(n5528), .A2(n5610), .ZN(n5616) );
  OR2_X1 U6606 ( .A1(n5612), .A2(n5611), .ZN(n5613) );
  NAND2_X1 U6607 ( .A1(n5614), .A2(n5613), .ZN(n7156) );
  OR2_X1 U6608 ( .A1(n5529), .A2(n7156), .ZN(n5615) );
  OAI211_X1 U6609 ( .C1(n7043), .C2(n7157), .A(n5616), .B(n5615), .ZN(n7952)
         );
  NAND2_X1 U6610 ( .A1(n7952), .A2(n6761), .ZN(n5617) );
  NAND2_X1 U6611 ( .A1(n5618), .A2(n5617), .ZN(n5619) );
  XNOR2_X1 U6612 ( .A(n5619), .B(n6081), .ZN(n5627) );
  NAND2_X1 U6613 ( .A1(n9714), .A2(n6083), .ZN(n5621) );
  NAND2_X1 U6614 ( .A1(n7952), .A2(n6062), .ZN(n5620) );
  NAND2_X1 U6615 ( .A1(n5621), .A2(n5620), .ZN(n5628) );
  AND2_X1 U6616 ( .A1(n5627), .A2(n5628), .ZN(n7971) );
  INV_X1 U6617 ( .A(n7971), .ZN(n5622) );
  NAND2_X1 U6618 ( .A1(n9715), .A2(n6083), .ZN(n5625) );
  NAND2_X1 U6619 ( .A1(n8065), .A2(n6062), .ZN(n5624) );
  NAND2_X1 U6620 ( .A1(n5625), .A2(n5624), .ZN(n7745) );
  OAI21_X1 U6621 ( .B1(n7743), .B2(n7744), .A(n7745), .ZN(n7908) );
  NAND2_X1 U6622 ( .A1(n5626), .A2(n7908), .ZN(n5654) );
  INV_X1 U6623 ( .A(n5627), .ZN(n5630) );
  INV_X1 U6624 ( .A(n5628), .ZN(n5629) );
  NAND2_X1 U6625 ( .A1(n5630), .A2(n5629), .ZN(n7973) );
  AND2_X1 U6626 ( .A1(n7973), .A2(n5631), .ZN(n5632) );
  OR2_X1 U6627 ( .A1(n5633), .A2(n5632), .ZN(n5652) );
  NAND2_X1 U6628 ( .A1(n5654), .A2(n5652), .ZN(n5649) );
  MUX2_X1 U6629 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .S(n7139), .Z(n5661) );
  XNOR2_X1 U6630 ( .A(n5661), .B(SI_8_), .ZN(n5660) );
  NAND2_X1 U6631 ( .A1(n7161), .A2(n8558), .ZN(n5641) );
  NOR2_X1 U6632 ( .A1(n5636), .A2(n5409), .ZN(n5637) );
  NAND2_X1 U6633 ( .A1(n5637), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n5639) );
  INV_X1 U6634 ( .A(n5637), .ZN(n5638) );
  NAND2_X1 U6635 ( .A1(n5638), .A2(n4970), .ZN(n5664) );
  AOI22_X1 U6636 ( .A1(n6072), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n10246), .B2(
        n7321), .ZN(n5640) );
  NAND2_X1 U6637 ( .A1(n5864), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5648) );
  NAND2_X1 U6638 ( .A1(n5642), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5669) );
  OR2_X1 U6639 ( .A1(n5642), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5643) );
  AND2_X1 U6640 ( .A1(n5669), .A2(n5643), .ZN(n8154) );
  NAND2_X1 U6641 ( .A1(n4855), .A2(n8154), .ZN(n5647) );
  NAND2_X1 U6642 ( .A1(n5644), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n5646) );
  NAND2_X1 U6643 ( .A1(n4854), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n5645) );
  NAND4_X1 U6644 ( .A1(n5648), .A2(n5647), .A3(n5646), .A4(n5645), .ZN(n8105)
         );
  AOI22_X1 U6645 ( .A1(n8155), .A2(n6767), .B1(n6083), .B2(n8105), .ZN(n5650)
         );
  NAND2_X1 U6646 ( .A1(n5649), .A2(n5650), .ZN(n8017) );
  INV_X1 U6647 ( .A(n5650), .ZN(n5651) );
  AND2_X1 U6648 ( .A1(n5652), .A2(n5651), .ZN(n5653) );
  NAND2_X1 U6649 ( .A1(n5654), .A2(n5653), .ZN(n8016) );
  NAND2_X1 U6650 ( .A1(n8155), .A2(n6761), .ZN(n5656) );
  NAND2_X1 U6651 ( .A1(n8105), .A2(n6062), .ZN(n5655) );
  NAND2_X1 U6652 ( .A1(n5656), .A2(n5655), .ZN(n5657) );
  XNOR2_X1 U6653 ( .A(n5657), .B(n6765), .ZN(n8018) );
  NAND2_X1 U6654 ( .A1(n8016), .A2(n8018), .ZN(n5658) );
  NAND2_X1 U6655 ( .A1(n8017), .A2(n5658), .ZN(n7999) );
  INV_X1 U6656 ( .A(n5661), .ZN(n5663) );
  INV_X1 U6657 ( .A(SI_8_), .ZN(n5662) );
  MUX2_X1 U6658 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(P2_DATAO_REG_9__SCAN_IN), 
        .S(n7139), .Z(n5687) );
  XNOR2_X1 U6659 ( .A(n5687), .B(n9161), .ZN(n5685) );
  XNOR2_X1 U6660 ( .A(n5686), .B(n5685), .ZN(n7169) );
  NAND2_X1 U6661 ( .A1(n7169), .A2(n8558), .ZN(n5667) );
  NAND2_X1 U6662 ( .A1(n5664), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5665) );
  XNOR2_X1 U6663 ( .A(n5665), .B(P1_IR_REG_9__SCAN_IN), .ZN(n7502) );
  AOI22_X1 U6664 ( .A1(n6072), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n10246), .B2(
        n7502), .ZN(n5666) );
  NAND2_X1 U6665 ( .A1(n10490), .A2(n6761), .ZN(n5677) );
  NAND2_X1 U6666 ( .A1(n5669), .A2(n5668), .ZN(n5670) );
  AND2_X1 U6667 ( .A1(n5696), .A2(n5670), .ZN(n8001) );
  NAND2_X1 U6668 ( .A1(n4855), .A2(n8001), .ZN(n5675) );
  NAND2_X1 U6669 ( .A1(n4850), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n5674) );
  NAND2_X1 U6670 ( .A1(n5644), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5673) );
  NAND2_X1 U6671 ( .A1(n4854), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5672) );
  NAND4_X1 U6672 ( .A1(n5675), .A2(n5674), .A3(n5673), .A4(n5672), .ZN(n9712)
         );
  NAND2_X1 U6673 ( .A1(n9712), .A2(n6767), .ZN(n5676) );
  NAND2_X1 U6674 ( .A1(n5677), .A2(n5676), .ZN(n5678) );
  XNOR2_X1 U6675 ( .A(n5678), .B(n6081), .ZN(n5680) );
  AND2_X1 U6676 ( .A1(n9712), .A2(n6083), .ZN(n5679) );
  AOI21_X1 U6677 ( .B1(n10490), .B2(n6062), .A(n5679), .ZN(n5681) );
  XNOR2_X1 U6678 ( .A(n5680), .B(n5681), .ZN(n8000) );
  NAND2_X1 U6679 ( .A1(n7999), .A2(n8000), .ZN(n5684) );
  INV_X1 U6680 ( .A(n5680), .ZN(n5682) );
  NAND2_X1 U6681 ( .A1(n5682), .A2(n5681), .ZN(n5683) );
  NAND2_X1 U6682 ( .A1(n5684), .A2(n5683), .ZN(n5707) );
  NAND2_X1 U6683 ( .A1(n5686), .A2(n5685), .ZN(n5690) );
  INV_X1 U6684 ( .A(n5687), .ZN(n5688) );
  NAND2_X1 U6685 ( .A1(n5688), .A2(n9161), .ZN(n5689) );
  MUX2_X1 U6686 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .S(n7139), .Z(n5714) );
  XNOR2_X1 U6687 ( .A(n5714), .B(n9155), .ZN(n5712) );
  XNOR2_X1 U6688 ( .A(n5713), .B(n5712), .ZN(n7175) );
  NAND2_X1 U6689 ( .A1(n7175), .A2(n8558), .ZN(n5694) );
  OR2_X1 U6690 ( .A1(n5691), .A2(n5409), .ZN(n5692) );
  XNOR2_X1 U6691 ( .A(n5692), .B(P1_IR_REG_10__SCAN_IN), .ZN(n7556) );
  AOI22_X1 U6692 ( .A1(n6072), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n10246), 
        .B2(n7556), .ZN(n5693) );
  NAND2_X1 U6693 ( .A1(n10501), .A2(n6761), .ZN(n5703) );
  NAND2_X1 U6694 ( .A1(n4850), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n5701) );
  INV_X1 U6695 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n5695) );
  NOR2_X1 U6696 ( .A1(n5696), .A2(n5695), .ZN(n5726) );
  AND2_X1 U6697 ( .A1(n5696), .A2(n5695), .ZN(n5697) );
  NOR2_X1 U6698 ( .A1(n5726), .A2(n5697), .ZN(n8279) );
  NAND2_X1 U6699 ( .A1(n4855), .A2(n8279), .ZN(n5700) );
  NAND2_X1 U6700 ( .A1(n8561), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5699) );
  NAND2_X1 U6701 ( .A1(n4854), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n5698) );
  NAND4_X1 U6702 ( .A1(n5701), .A2(n5700), .A3(n5699), .A4(n5698), .ZN(n9711)
         );
  NAND2_X1 U6703 ( .A1(n9711), .A2(n6062), .ZN(n5702) );
  NAND2_X1 U6704 ( .A1(n5703), .A2(n5702), .ZN(n5704) );
  XNOR2_X1 U6705 ( .A(n5704), .B(n6765), .ZN(n5708) );
  NAND2_X1 U6706 ( .A1(n5707), .A2(n5708), .ZN(n8223) );
  NAND2_X1 U6707 ( .A1(n10501), .A2(n6767), .ZN(n5706) );
  NAND2_X1 U6708 ( .A1(n9711), .A2(n6083), .ZN(n5705) );
  NAND2_X1 U6709 ( .A1(n5706), .A2(n5705), .ZN(n8225) );
  NAND2_X1 U6710 ( .A1(n8223), .A2(n8225), .ZN(n5711) );
  INV_X1 U6711 ( .A(n5707), .ZN(n5710) );
  INV_X1 U6712 ( .A(n5708), .ZN(n5709) );
  NAND2_X1 U6713 ( .A1(n5710), .A2(n5709), .ZN(n8224) );
  NAND2_X1 U6714 ( .A1(n5711), .A2(n8224), .ZN(n8248) );
  INV_X1 U6715 ( .A(n5714), .ZN(n5715) );
  NAND2_X1 U6716 ( .A1(n5715), .A2(n9155), .ZN(n5716) );
  MUX2_X1 U6717 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .S(n7139), .Z(n5717) );
  NAND2_X1 U6718 ( .A1(n5717), .A2(SI_11_), .ZN(n5739) );
  OAI21_X1 U6719 ( .B1(n5717), .B2(SI_11_), .A(n5739), .ZN(n5719) );
  NAND2_X1 U6720 ( .A1(n5720), .A2(n5719), .ZN(n5721) );
  NAND2_X1 U6721 ( .A1(n5740), .A2(n5721), .ZN(n7180) );
  OR2_X1 U6722 ( .A1(n7180), .A2(n5529), .ZN(n5725) );
  NAND2_X1 U6723 ( .A1(n5722), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5723) );
  XNOR2_X1 U6724 ( .A(n5723), .B(P1_IR_REG_11__SCAN_IN), .ZN(n10268) );
  AOI22_X1 U6725 ( .A1(n6072), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n10246), 
        .B2(n10268), .ZN(n5724) );
  NAND2_X1 U6726 ( .A1(n9446), .A2(n6761), .ZN(n5733) );
  NAND2_X1 U6727 ( .A1(n4851), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n5731) );
  NOR2_X1 U6728 ( .A1(n5726), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5727) );
  OR2_X1 U6729 ( .A1(n5748), .A2(n5727), .ZN(n8251) );
  INV_X1 U6730 ( .A(n8251), .ZN(n8330) );
  NAND2_X1 U6731 ( .A1(n4855), .A2(n8330), .ZN(n5730) );
  NAND2_X1 U6732 ( .A1(n8561), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5729) );
  NAND2_X1 U6733 ( .A1(n4854), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n5728) );
  NAND4_X1 U6734 ( .A1(n5731), .A2(n5730), .A3(n5729), .A4(n5728), .ZN(n9710)
         );
  NAND2_X1 U6735 ( .A1(n9710), .A2(n6767), .ZN(n5732) );
  NAND2_X1 U6736 ( .A1(n5733), .A2(n5732), .ZN(n5734) );
  XNOR2_X1 U6737 ( .A(n5734), .B(n6765), .ZN(n5737) );
  AND2_X1 U6738 ( .A1(n9710), .A2(n6083), .ZN(n5735) );
  AOI21_X1 U6739 ( .B1(n9446), .B2(n6062), .A(n5735), .ZN(n5736) );
  XNOR2_X1 U6740 ( .A(n5737), .B(n5736), .ZN(n8249) );
  NAND2_X1 U6741 ( .A1(n5737), .A2(n5736), .ZN(n5738) );
  MUX2_X1 U6742 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .S(n7142), .Z(n5742) );
  NAND2_X1 U6743 ( .A1(n5744), .A2(n9153), .ZN(n5745) );
  NAND2_X1 U6744 ( .A1(n5760), .A2(n5745), .ZN(n7330) );
  NOR2_X1 U6745 ( .A1(n5722), .A2(P1_IR_REG_11__SCAN_IN), .ZN(n5788) );
  OR2_X1 U6746 ( .A1(n5788), .A2(n5409), .ZN(n5762) );
  XNOR2_X1 U6747 ( .A(n5762), .B(P1_IR_REG_12__SCAN_IN), .ZN(n7709) );
  AOI22_X1 U6748 ( .A1(n6072), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n10246), 
        .B2(n7709), .ZN(n5746) );
  NAND2_X2 U6749 ( .A1(n5747), .A2(n5746), .ZN(n10080) );
  NAND2_X1 U6750 ( .A1(n10080), .A2(n6761), .ZN(n5755) );
  NAND2_X1 U6751 ( .A1(n4850), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n5753) );
  NAND2_X1 U6752 ( .A1(n5748), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n5796) );
  OR2_X1 U6753 ( .A1(n5748), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n5749) );
  AND2_X1 U6754 ( .A1(n5796), .A2(n5749), .ZN(n8390) );
  NAND2_X1 U6755 ( .A1(n4855), .A2(n8390), .ZN(n5752) );
  NAND2_X1 U6756 ( .A1(n5644), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5751) );
  NAND2_X1 U6757 ( .A1(n4854), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n5750) );
  NAND4_X1 U6758 ( .A1(n5753), .A2(n5752), .A3(n5751), .A4(n5750), .ZN(n9709)
         );
  NAND2_X1 U6759 ( .A1(n9709), .A2(n6767), .ZN(n5754) );
  NAND2_X1 U6760 ( .A1(n5755), .A2(n5754), .ZN(n5756) );
  XNOR2_X1 U6761 ( .A(n5756), .B(n6765), .ZN(n8352) );
  AND2_X1 U6762 ( .A1(n9709), .A2(n6083), .ZN(n5757) );
  AOI21_X1 U6763 ( .B1(n10080), .B2(n6767), .A(n5757), .ZN(n8353) );
  AND2_X1 U6764 ( .A1(n8352), .A2(n8353), .ZN(n5758) );
  MUX2_X1 U6765 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n7142), .Z(n5780) );
  XNOR2_X1 U6766 ( .A(n5780), .B(SI_13_), .ZN(n5781) );
  NAND2_X1 U6767 ( .A1(n7543), .A2(n8558), .ZN(n5766) );
  INV_X1 U6768 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n5761) );
  NAND2_X1 U6769 ( .A1(n5762), .A2(n5761), .ZN(n5763) );
  NAND2_X1 U6770 ( .A1(n5763), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5764) );
  XNOR2_X1 U6771 ( .A(n5764), .B(P1_IR_REG_13__SCAN_IN), .ZN(n10293) );
  AOI22_X1 U6772 ( .A1(n6072), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n10246), 
        .B2(n10293), .ZN(n5765) );
  NAND2_X2 U6773 ( .A1(n5766), .A2(n5765), .ZN(n6157) );
  NAND2_X1 U6774 ( .A1(n6157), .A2(n6761), .ZN(n5772) );
  NAND2_X1 U6775 ( .A1(n4851), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n5770) );
  XNOR2_X1 U6776 ( .A(n5796), .B(P1_REG3_REG_13__SCAN_IN), .ZN(n8479) );
  NAND2_X1 U6777 ( .A1(n4855), .A2(n8479), .ZN(n5769) );
  NAND2_X1 U6778 ( .A1(n8561), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n5768) );
  NAND2_X1 U6779 ( .A1(n4854), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n5767) );
  NAND4_X1 U6780 ( .A1(n5770), .A2(n5769), .A3(n5768), .A4(n5767), .ZN(n9708)
         );
  NAND2_X1 U6781 ( .A1(n9708), .A2(n6062), .ZN(n5771) );
  NAND2_X1 U6782 ( .A1(n5772), .A2(n5771), .ZN(n5773) );
  XNOR2_X1 U6783 ( .A(n5773), .B(n6081), .ZN(n5776) );
  NAND2_X1 U6784 ( .A1(n6157), .A2(n6062), .ZN(n5775) );
  NAND2_X1 U6785 ( .A1(n9708), .A2(n6083), .ZN(n5774) );
  NAND2_X1 U6786 ( .A1(n5775), .A2(n5774), .ZN(n5777) );
  AND2_X1 U6787 ( .A1(n5776), .A2(n5777), .ZN(n8362) );
  INV_X1 U6788 ( .A(n5776), .ZN(n5779) );
  INV_X1 U6789 ( .A(n5777), .ZN(n5778) );
  NAND2_X1 U6790 ( .A1(n5779), .A2(n5778), .ZN(n8361) );
  MUX2_X1 U6791 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n7142), .Z(n5783) );
  NAND2_X1 U6792 ( .A1(n5783), .A2(SI_14_), .ZN(n5808) );
  OAI21_X1 U6793 ( .B1(n5783), .B2(SI_14_), .A(n5808), .ZN(n5784) );
  NAND2_X1 U6794 ( .A1(n5785), .A2(n5784), .ZN(n5786) );
  NAND2_X1 U6795 ( .A1(n5786), .A2(n5809), .ZN(n7587) );
  NOR2_X1 U6796 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n5787) );
  NAND2_X1 U6797 ( .A1(n5788), .A2(n5787), .ZN(n5790) );
  NAND2_X1 U6798 ( .A1(n5790), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5789) );
  MUX2_X1 U6799 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5789), .S(
        P1_IR_REG_14__SCAN_IN), .Z(n5791) );
  AOI22_X1 U6800 ( .A1(n6072), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n10246), 
        .B2(n8077), .ZN(n5792) );
  NAND2_X2 U6801 ( .A1(n5793), .A2(n5792), .ZN(n10068) );
  NAND2_X1 U6802 ( .A1(n10068), .A2(n6761), .ZN(n5803) );
  INV_X1 U6803 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n5795) );
  OAI21_X1 U6804 ( .B1(n5796), .B2(n5795), .A(n5794), .ZN(n5797) );
  AND2_X1 U6805 ( .A1(n5797), .A2(n5820), .ZN(n9967) );
  NAND2_X1 U6806 ( .A1(n4855), .A2(n9967), .ZN(n5801) );
  NAND2_X1 U6807 ( .A1(n4851), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n5800) );
  NAND2_X1 U6808 ( .A1(n8561), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5799) );
  NAND2_X1 U6809 ( .A1(n4854), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n5798) );
  NAND4_X1 U6810 ( .A1(n5801), .A2(n5800), .A3(n5799), .A4(n5798), .ZN(n9707)
         );
  NAND2_X1 U6811 ( .A1(n9707), .A2(n4856), .ZN(n5802) );
  NAND2_X1 U6812 ( .A1(n5803), .A2(n5802), .ZN(n5804) );
  NAND2_X1 U6813 ( .A1(n10068), .A2(n5435), .ZN(n5806) );
  NAND2_X1 U6814 ( .A1(n9707), .A2(n6083), .ZN(n5805) );
  NAND2_X1 U6815 ( .A1(n5806), .A2(n5805), .ZN(n9307) );
  NAND2_X1 U6816 ( .A1(n9304), .A2(n9307), .ZN(n5807) );
  NAND2_X1 U6817 ( .A1(n4893), .A2(n4908), .ZN(n9305) );
  MUX2_X1 U6818 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .S(n7142), .Z(n5810) );
  NAND2_X1 U6819 ( .A1(n5810), .A2(SI_15_), .ZN(n5834) );
  INV_X1 U6820 ( .A(n5810), .ZN(n5811) );
  NAND2_X1 U6821 ( .A1(n5811), .A2(n9121), .ZN(n5812) );
  NAND2_X1 U6822 ( .A1(n5836), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5817) );
  INV_X1 U6823 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n5816) );
  XNOR2_X1 U6824 ( .A(n5817), .B(n5816), .ZN(n8261) );
  INV_X1 U6825 ( .A(n8261), .ZN(n8083) );
  AOI22_X1 U6826 ( .A1(n6072), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n10246), 
        .B2(n8083), .ZN(n5818) );
  NAND2_X2 U6827 ( .A1(n5819), .A2(n5818), .ZN(n10062) );
  NAND2_X1 U6828 ( .A1(n10062), .A2(n6761), .ZN(n5828) );
  NAND2_X1 U6829 ( .A1(n4850), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n5826) );
  AND2_X1 U6830 ( .A1(n5820), .A2(n8082), .ZN(n5821) );
  NOR2_X1 U6831 ( .A1(n5840), .A2(n5821), .ZN(n9956) );
  NAND2_X1 U6832 ( .A1(n4855), .A2(n9956), .ZN(n5825) );
  NAND2_X1 U6833 ( .A1(n8561), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n5824) );
  NAND2_X1 U6834 ( .A1(n4854), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n5823) );
  NAND4_X1 U6835 ( .A1(n5826), .A2(n5825), .A3(n5824), .A4(n5823), .ZN(n9706)
         );
  NAND2_X1 U6836 ( .A1(n9706), .A2(n4856), .ZN(n5827) );
  NAND2_X1 U6837 ( .A1(n5828), .A2(n5827), .ZN(n5829) );
  XNOR2_X1 U6838 ( .A(n5829), .B(n6765), .ZN(n5831) );
  INV_X1 U6839 ( .A(n9706), .ZN(n9976) );
  OAI22_X1 U6840 ( .A1(n9959), .A2(n6762), .B1(n9976), .B2(n6769), .ZN(n9427)
         );
  NAND2_X2 U6841 ( .A1(n9423), .A2(n9427), .ZN(n9424) );
  INV_X1 U6842 ( .A(n5830), .ZN(n5833) );
  INV_X1 U6843 ( .A(n5831), .ZN(n5832) );
  NAND2_X1 U6844 ( .A1(n5833), .A2(n5832), .ZN(n9425) );
  NAND2_X2 U6845 ( .A1(n9424), .A2(n9425), .ZN(n9422) );
  MUX2_X1 U6846 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(P2_DATAO_REG_16__SCAN_IN), 
        .S(n7142), .Z(n5853) );
  XNOR2_X1 U6847 ( .A(n5853), .B(SI_16_), .ZN(n5854) );
  XNOR2_X1 U6848 ( .A(n5855), .B(n5854), .ZN(n7801) );
  NAND2_X1 U6849 ( .A1(n7801), .A2(n8558), .ZN(n5839) );
  NAND2_X1 U6850 ( .A1(n5860), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5837) );
  XNOR2_X1 U6851 ( .A(n5837), .B(P1_IR_REG_16__SCAN_IN), .ZN(n8295) );
  AOI22_X1 U6852 ( .A1(n6072), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n10246), 
        .B2(n8295), .ZN(n5838) );
  NAND2_X2 U6853 ( .A1(n5839), .A2(n5838), .ZN(n10058) );
  NOR2_X1 U6854 ( .A1(n5840), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n5841) );
  OR2_X1 U6855 ( .A1(n5865), .A2(n5841), .ZN(n9932) );
  INV_X1 U6856 ( .A(n9932), .ZN(n5842) );
  NAND2_X1 U6857 ( .A1(n4855), .A2(n5842), .ZN(n5846) );
  NAND2_X1 U6858 ( .A1(n4851), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n5845) );
  NAND2_X1 U6859 ( .A1(n8561), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n5844) );
  NAND2_X1 U6860 ( .A1(n4854), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n5843) );
  NAND4_X1 U6861 ( .A1(n5846), .A2(n5845), .A3(n5844), .A4(n5843), .ZN(n9705)
         );
  AOI22_X1 U6862 ( .A1(n10058), .A2(n4856), .B1(n6083), .B2(n9705), .ZN(n5851)
         );
  NAND2_X1 U6863 ( .A1(n10058), .A2(n6761), .ZN(n5848) );
  NAND2_X1 U6864 ( .A1(n9705), .A2(n6767), .ZN(n5847) );
  NAND2_X1 U6865 ( .A1(n5848), .A2(n5847), .ZN(n5849) );
  XNOR2_X1 U6866 ( .A(n5849), .B(n6081), .ZN(n5850) );
  XOR2_X1 U6867 ( .A(n5851), .B(n5850), .Z(n9351) );
  INV_X1 U6868 ( .A(n5850), .ZN(n5852) );
  MUX2_X1 U6869 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(P2_DATAO_REG_17__SCAN_IN), 
        .S(n7142), .Z(n5856) );
  NAND2_X1 U6870 ( .A1(n5856), .A2(SI_17_), .ZN(n5894) );
  OAI21_X1 U6871 ( .B1(n5856), .B2(SI_17_), .A(n5894), .ZN(n5857) );
  NAND2_X1 U6872 ( .A1(n5858), .A2(n5857), .ZN(n5859) );
  NAND2_X1 U6873 ( .A1(n7916), .A2(n8558), .ZN(n5863) );
  NAND2_X1 U6874 ( .A1(n5861), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5883) );
  XNOR2_X1 U6875 ( .A(n5883), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9727) );
  AOI22_X1 U6876 ( .A1(n6072), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n10246), 
        .B2(n9727), .ZN(n5862) );
  NAND2_X1 U6877 ( .A1(n10049), .A2(n6761), .ZN(n5872) );
  NAND2_X1 U6878 ( .A1(n4851), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n5870) );
  NOR2_X1 U6879 ( .A1(n5865), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n5866) );
  OR2_X1 U6880 ( .A1(n5888), .A2(n5866), .ZN(n9362) );
  INV_X1 U6881 ( .A(n9362), .ZN(n9915) );
  NAND2_X1 U6882 ( .A1(n4855), .A2(n9915), .ZN(n5869) );
  NAND2_X1 U6883 ( .A1(n8561), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n5868) );
  NAND2_X1 U6884 ( .A1(n4854), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n5867) );
  NAND4_X1 U6885 ( .A1(n5870), .A2(n5869), .A3(n5868), .A4(n5867), .ZN(n9899)
         );
  NAND2_X1 U6886 ( .A1(n9899), .A2(n6767), .ZN(n5871) );
  NAND2_X1 U6887 ( .A1(n5872), .A2(n5871), .ZN(n5873) );
  XNOR2_X1 U6888 ( .A(n5873), .B(n6081), .ZN(n9358) );
  NAND2_X1 U6889 ( .A1(n10049), .A2(n6767), .ZN(n5875) );
  NAND2_X1 U6890 ( .A1(n9899), .A2(n6083), .ZN(n5874) );
  NAND2_X1 U6891 ( .A1(n5875), .A2(n5874), .ZN(n5876) );
  INV_X1 U6892 ( .A(n5876), .ZN(n9357) );
  MUX2_X1 U6893 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n7142), .Z(n5877) );
  NAND2_X1 U6894 ( .A1(n5877), .A2(SI_18_), .ZN(n5895) );
  OAI21_X1 U6895 ( .B1(n5877), .B2(SI_18_), .A(n5895), .ZN(n5879) );
  NAND2_X1 U6896 ( .A1(n5878), .A2(n5879), .ZN(n5881) );
  INV_X1 U6897 ( .A(n5879), .ZN(n5896) );
  AND2_X2 U6898 ( .A1(n5881), .A2(n5880), .ZN(n8012) );
  NAND2_X1 U6899 ( .A1(n8012), .A2(n8558), .ZN(n5887) );
  INV_X1 U6900 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5882) );
  NAND2_X1 U6901 ( .A1(n5883), .A2(n5882), .ZN(n5884) );
  NAND2_X1 U6902 ( .A1(n5884), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5885) );
  XNOR2_X1 U6903 ( .A(n5885), .B(P1_IR_REG_18__SCAN_IN), .ZN(n10304) );
  AOI22_X1 U6904 ( .A1(n6072), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n10246), 
        .B2(n10304), .ZN(n5886) );
  AND2_X2 U6905 ( .A1(n5887), .A2(n5886), .ZN(n9896) );
  AOI22_X1 U6906 ( .A1(n4850), .A2(P1_REG1_REG_18__SCAN_IN), .B1(n8561), .B2(
        P1_REG0_REG_18__SCAN_IN), .ZN(n5891) );
  NAND2_X1 U6907 ( .A1(n5888), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n5903) );
  OR2_X1 U6908 ( .A1(n5888), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n5889) );
  AND2_X1 U6909 ( .A1(n5903), .A2(n5889), .ZN(n9894) );
  AOI22_X1 U6910 ( .A1(n4855), .A2(n9894), .B1(n4854), .B2(
        P1_REG2_REG_18__SCAN_IN), .ZN(n5890) );
  OAI22_X1 U6911 ( .A1(n9896), .A2(n5987), .B1(n9907), .B2(n6762), .ZN(n5892)
         );
  XNOR2_X1 U6912 ( .A(n5892), .B(n6081), .ZN(n9400) );
  INV_X1 U6913 ( .A(n9400), .ZN(n5893) );
  OAI22_X1 U6914 ( .A1(n9896), .A2(n6762), .B1(n9907), .B2(n6769), .ZN(n9399)
         );
  AND2_X1 U6915 ( .A1(n5894), .A2(n5895), .ZN(n5898) );
  INV_X1 U6916 ( .A(n5895), .ZN(n5897) );
  MUX2_X1 U6917 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(P2_DATAO_REG_19__SCAN_IN), 
        .S(n7142), .Z(n5917) );
  XNOR2_X1 U6918 ( .A(n5917), .B(SI_19_), .ZN(n5915) );
  XNOR2_X1 U6919 ( .A(n5916), .B(n5915), .ZN(n8007) );
  NAND2_X1 U6920 ( .A1(n8007), .A2(n8558), .ZN(n5901) );
  AOI22_X1 U6921 ( .A1(n6072), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n10246), 
        .B2(n10411), .ZN(n5900) );
  NAND2_X2 U6922 ( .A1(n5901), .A2(n5900), .ZN(n10039) );
  NAND2_X1 U6923 ( .A1(n10039), .A2(n6761), .ZN(n5909) );
  NAND2_X1 U6924 ( .A1(n4850), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n5907) );
  INV_X1 U6925 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n5902) );
  AOI21_X1 U6926 ( .B1(n5903), .B2(n5902), .A(n5922), .ZN(n9878) );
  NAND2_X1 U6927 ( .A1(n4855), .A2(n9878), .ZN(n5906) );
  NAND2_X1 U6928 ( .A1(n8561), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n5905) );
  NAND2_X1 U6929 ( .A1(n4854), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n5904) );
  NAND4_X1 U6930 ( .A1(n5907), .A2(n5906), .A3(n5905), .A4(n5904), .ZN(n9900)
         );
  NAND2_X1 U6931 ( .A1(n9900), .A2(n6062), .ZN(n5908) );
  NAND2_X1 U6932 ( .A1(n5909), .A2(n5908), .ZN(n5910) );
  XNOR2_X1 U6933 ( .A(n5910), .B(n6765), .ZN(n5913) );
  AND2_X1 U6934 ( .A1(n9900), .A2(n6083), .ZN(n5911) );
  AOI21_X1 U6935 ( .B1(n10039), .B2(n5435), .A(n5911), .ZN(n5912) );
  NAND2_X1 U6936 ( .A1(n5913), .A2(n5912), .ZN(n5914) );
  OAI21_X1 U6937 ( .B1(n5913), .B2(n5912), .A(n5914), .ZN(n9325) );
  INV_X1 U6938 ( .A(n5917), .ZN(n5919) );
  INV_X1 U6939 ( .A(SI_19_), .ZN(n5918) );
  MUX2_X1 U6940 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(P2_DATAO_REG_20__SCAN_IN), 
        .S(n7142), .Z(n5936) );
  XNOR2_X1 U6941 ( .A(n5936), .B(n9020), .ZN(n5937) );
  XNOR2_X1 U6942 ( .A(n5938), .B(n5937), .ZN(n8216) );
  NAND2_X1 U6943 ( .A1(n8216), .A2(n8558), .ZN(n5921) );
  NAND2_X1 U6944 ( .A1(n6072), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n5920) );
  NAND2_X1 U6945 ( .A1(n10035), .A2(n6761), .ZN(n5928) );
  NAND2_X1 U6946 ( .A1(n4851), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n5926) );
  NAND2_X1 U6947 ( .A1(n5922), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n5949) );
  OAI21_X1 U6948 ( .B1(P1_REG3_REG_20__SCAN_IN), .B2(n5922), .A(n5949), .ZN(
        n9383) );
  INV_X1 U6949 ( .A(n9383), .ZN(n9864) );
  NAND2_X1 U6950 ( .A1(n4855), .A2(n9864), .ZN(n5925) );
  NAND2_X1 U6951 ( .A1(n8561), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n5924) );
  NAND2_X1 U6952 ( .A1(n4854), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n5923) );
  NAND4_X1 U6953 ( .A1(n5926), .A2(n5925), .A3(n5924), .A4(n5923), .ZN(n9883)
         );
  NAND2_X1 U6954 ( .A1(n9883), .A2(n6062), .ZN(n5927) );
  NAND2_X1 U6955 ( .A1(n5928), .A2(n5927), .ZN(n5929) );
  XNOR2_X1 U6956 ( .A(n5929), .B(n6081), .ZN(n5935) );
  INV_X1 U6957 ( .A(n5935), .ZN(n5933) );
  NAND2_X1 U6958 ( .A1(n10035), .A2(n5435), .ZN(n5931) );
  NAND2_X1 U6959 ( .A1(n9883), .A2(n6083), .ZN(n5930) );
  NAND2_X1 U6960 ( .A1(n5931), .A2(n5930), .ZN(n5934) );
  INV_X1 U6961 ( .A(n5934), .ZN(n5932) );
  NAND2_X1 U6962 ( .A1(n5933), .A2(n5932), .ZN(n9377) );
  AND2_X1 U6963 ( .A1(n5935), .A2(n5934), .ZN(n9378) );
  MUX2_X1 U6964 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(P2_DATAO_REG_21__SCAN_IN), 
        .S(n7142), .Z(n5939) );
  NAND2_X1 U6965 ( .A1(n5939), .A2(SI_21_), .ZN(n5962) );
  INV_X1 U6966 ( .A(n5939), .ZN(n5940) );
  NAND2_X1 U6967 ( .A1(n5940), .A2(n9144), .ZN(n5941) );
  NAND2_X1 U6968 ( .A1(n5962), .A2(n5941), .ZN(n5944) );
  INV_X1 U6969 ( .A(n5944), .ZN(n5942) );
  NAND2_X1 U6970 ( .A1(n5943), .A2(n5942), .ZN(n5963) );
  INV_X1 U6971 ( .A(n5943), .ZN(n5945) );
  NAND2_X1 U6972 ( .A1(n5945), .A2(n5944), .ZN(n5946) );
  NAND2_X1 U6973 ( .A1(n5963), .A2(n5946), .ZN(n8220) );
  OR2_X1 U6974 ( .A1(n8220), .A2(n5529), .ZN(n5948) );
  NAND2_X1 U6975 ( .A1(n6072), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n5947) );
  NAND2_X1 U6976 ( .A1(n10030), .A2(n6761), .ZN(n5955) );
  INV_X1 U6977 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n9335) );
  AOI21_X1 U6978 ( .B1(n9335), .B2(n5949), .A(n5966), .ZN(n9855) );
  NAND2_X1 U6979 ( .A1(n4855), .A2(n9855), .ZN(n5953) );
  NAND2_X1 U6980 ( .A1(n4850), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n5952) );
  NAND2_X1 U6981 ( .A1(n8561), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n5951) );
  NAND2_X1 U6982 ( .A1(n4854), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n5950) );
  NAND4_X1 U6983 ( .A1(n5953), .A2(n5952), .A3(n5951), .A4(n5950), .ZN(n9870)
         );
  NAND2_X1 U6984 ( .A1(n9870), .A2(n4856), .ZN(n5954) );
  NAND2_X1 U6985 ( .A1(n5955), .A2(n5954), .ZN(n5956) );
  XNOR2_X1 U6986 ( .A(n5956), .B(n6765), .ZN(n5961) );
  INV_X1 U6987 ( .A(n5961), .ZN(n5959) );
  AND2_X1 U6988 ( .A1(n9870), .A2(n6083), .ZN(n5957) );
  AOI21_X1 U6989 ( .B1(n10030), .B2(n5435), .A(n5957), .ZN(n5960) );
  INV_X1 U6990 ( .A(n5960), .ZN(n5958) );
  NAND2_X1 U6991 ( .A1(n5959), .A2(n5958), .ZN(n9331) );
  AND2_X1 U6992 ( .A1(n5961), .A2(n5960), .ZN(n9330) );
  NAND2_X1 U6993 ( .A1(n5963), .A2(n5962), .ZN(n5996) );
  MUX2_X1 U6994 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(P2_DATAO_REG_22__SCAN_IN), 
        .S(n7142), .Z(n5977) );
  XNOR2_X1 U6995 ( .A(n5977), .B(SI_22_), .ZN(n5994) );
  XNOR2_X1 U6996 ( .A(n5996), .B(n5994), .ZN(n8349) );
  NAND2_X1 U6997 ( .A1(n8349), .A2(n8558), .ZN(n5965) );
  NAND2_X1 U6998 ( .A1(n6072), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n5964) );
  NAND2_X1 U6999 ( .A1(n5966), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n5984) );
  OAI21_X1 U7000 ( .B1(P1_REG3_REG_22__SCAN_IN), .B2(n5966), .A(n5984), .ZN(
        n9391) );
  INV_X1 U7001 ( .A(n9391), .ZN(n9836) );
  NAND2_X1 U7002 ( .A1(n4855), .A2(n9836), .ZN(n5970) );
  NAND2_X1 U7003 ( .A1(n4851), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n5969) );
  NAND2_X1 U7004 ( .A1(n8561), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n5968) );
  NAND2_X1 U7005 ( .A1(n4854), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n5967) );
  NAND4_X1 U7006 ( .A1(n5970), .A2(n5969), .A3(n5968), .A4(n5967), .ZN(n9851)
         );
  AOI22_X1 U7007 ( .A1(n9835), .A2(n4856), .B1(n6083), .B2(n9851), .ZN(n5974)
         );
  NAND2_X1 U7008 ( .A1(n9835), .A2(n6761), .ZN(n5972) );
  NAND2_X1 U7009 ( .A1(n9851), .A2(n5435), .ZN(n5971) );
  NAND2_X1 U7010 ( .A1(n5972), .A2(n5971), .ZN(n5973) );
  XNOR2_X1 U7011 ( .A(n5973), .B(n6081), .ZN(n5976) );
  XOR2_X1 U7012 ( .A(n5974), .B(n5976), .Z(n9388) );
  INV_X1 U7013 ( .A(n5974), .ZN(n5975) );
  OAI22_X1 U7014 ( .A1(n9389), .A2(n9388), .B1(n5976), .B2(n5975), .ZN(n6026)
         );
  INV_X1 U7015 ( .A(n5977), .ZN(n5979) );
  INV_X1 U7016 ( .A(SI_22_), .ZN(n5978) );
  NAND2_X1 U7017 ( .A1(n5979), .A2(n5978), .ZN(n5998) );
  NAND2_X1 U7018 ( .A1(n5980), .A2(n5998), .ZN(n5981) );
  MUX2_X1 U7019 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(P2_DATAO_REG_23__SCAN_IN), 
        .S(n7142), .Z(n5989) );
  XNOR2_X1 U7020 ( .A(n5989), .B(n5990), .ZN(n5992) );
  NAND2_X1 U7021 ( .A1(n8396), .A2(n8558), .ZN(n5983) );
  NAND2_X1 U7022 ( .A1(n6072), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n5982) );
  AOI22_X1 U7023 ( .A1(n4851), .A2(P1_REG1_REG_23__SCAN_IN), .B1(n8561), .B2(
        P1_REG0_REG_23__SCAN_IN), .ZN(n5986) );
  INV_X1 U7024 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n9317) );
  AOI21_X1 U7025 ( .B1(n9317), .B2(n5984), .A(n6011), .ZN(n9316) );
  AOI22_X1 U7026 ( .A1(n4855), .A2(n9316), .B1(n4854), .B2(
        P1_REG2_REG_23__SCAN_IN), .ZN(n5985) );
  OAI22_X1 U7027 ( .A1(n9820), .A2(n5987), .B1(n9394), .B2(n6762), .ZN(n5988)
         );
  XOR2_X1 U7028 ( .A(n6081), .B(n5988), .Z(n6027) );
  NAND2_X1 U7029 ( .A1(n6026), .A2(n6027), .ZN(n9313) );
  OAI22_X1 U7030 ( .A1(n9820), .A2(n6762), .B1(n9394), .B2(n6769), .ZN(n9315)
         );
  NAND2_X1 U7031 ( .A1(n9313), .A2(n9315), .ZN(n9368) );
  INV_X1 U7032 ( .A(n5989), .ZN(n5991) );
  NAND2_X1 U7033 ( .A1(n5991), .A2(n5990), .ZN(n5997) );
  INV_X1 U7034 ( .A(n5997), .ZN(n5993) );
  NOR2_X1 U7035 ( .A1(n5993), .A2(n5992), .ZN(n6000) );
  OR2_X1 U7036 ( .A1(n5994), .A2(n6000), .ZN(n5995) );
  AND2_X1 U7037 ( .A1(n5998), .A2(n5997), .ZN(n5999) );
  OR2_X1 U7038 ( .A1(n6000), .A2(n5999), .ZN(n6004) );
  MUX2_X1 U7039 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(P2_DATAO_REG_24__SCAN_IN), 
        .S(n7142), .Z(n6001) );
  NAND2_X1 U7040 ( .A1(n6001), .A2(SI_24_), .ZN(n6031) );
  OAI21_X1 U7041 ( .B1(n6001), .B2(SI_24_), .A(n6031), .ZN(n6006) );
  INV_X1 U7042 ( .A(n6006), .ZN(n6002) );
  NAND2_X1 U7043 ( .A1(n6005), .A2(n6004), .ZN(n6007) );
  NAND2_X1 U7044 ( .A1(n6007), .A2(n6006), .ZN(n6008) );
  NAND2_X1 U7045 ( .A1(n8402), .A2(n8558), .ZN(n6010) );
  NAND2_X1 U7046 ( .A1(n6072), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n6009) );
  NAND2_X1 U7047 ( .A1(n10014), .A2(n6761), .ZN(n6018) );
  NAND2_X1 U7048 ( .A1(n6011), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n6036) );
  OAI21_X1 U7049 ( .B1(n6011), .B2(P1_REG3_REG_24__SCAN_IN), .A(n6036), .ZN(
        n6012) );
  INV_X1 U7050 ( .A(n6012), .ZN(n9809) );
  NAND2_X1 U7051 ( .A1(n4855), .A2(n9809), .ZN(n6016) );
  NAND2_X1 U7052 ( .A1(n4850), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n6015) );
  NAND2_X1 U7053 ( .A1(n8561), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n6014) );
  NAND2_X1 U7054 ( .A1(n4854), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n6013) );
  NAND4_X1 U7055 ( .A1(n6016), .A2(n6015), .A3(n6014), .A4(n6013), .ZN(n9824)
         );
  NAND2_X1 U7056 ( .A1(n9824), .A2(n4856), .ZN(n6017) );
  NAND2_X1 U7057 ( .A1(n6018), .A2(n6017), .ZN(n6019) );
  XNOR2_X1 U7058 ( .A(n6019), .B(n6765), .ZN(n6021) );
  AND2_X1 U7059 ( .A1(n9824), .A2(n6083), .ZN(n6020) );
  AOI21_X1 U7060 ( .B1(n10014), .B2(n4856), .A(n6020), .ZN(n6022) );
  NAND2_X1 U7061 ( .A1(n6021), .A2(n6022), .ZN(n6030) );
  INV_X1 U7062 ( .A(n6021), .ZN(n6024) );
  INV_X1 U7063 ( .A(n6022), .ZN(n6023) );
  NAND2_X1 U7064 ( .A1(n6024), .A2(n6023), .ZN(n6025) );
  AND2_X1 U7065 ( .A1(n6030), .A2(n6025), .ZN(n9369) );
  INV_X1 U7066 ( .A(n6026), .ZN(n6029) );
  INV_X1 U7067 ( .A(n6027), .ZN(n6028) );
  NAND2_X1 U7068 ( .A1(n6029), .A2(n6028), .ZN(n9370) );
  MUX2_X1 U7069 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(P2_DATAO_REG_25__SCAN_IN), 
        .S(n7142), .Z(n6045) );
  XNOR2_X1 U7070 ( .A(n6045), .B(SI_25_), .ZN(n6046) );
  XNOR2_X1 U7071 ( .A(n6047), .B(n6046), .ZN(n8434) );
  NAND2_X1 U7072 ( .A1(n8434), .A2(n8558), .ZN(n6034) );
  NAND2_X1 U7073 ( .A1(n6072), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n6033) );
  NAND2_X1 U7074 ( .A1(n4850), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n6041) );
  INV_X1 U7075 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n6037) );
  INV_X1 U7076 ( .A(n6036), .ZN(n6035) );
  NAND2_X1 U7077 ( .A1(n6035), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n6050) );
  INV_X1 U7078 ( .A(n6050), .ZN(n6052) );
  AOI21_X1 U7079 ( .B1(n6037), .B2(n6036), .A(n6052), .ZN(n9790) );
  NAND2_X1 U7080 ( .A1(n4855), .A2(n9790), .ZN(n6040) );
  NAND2_X1 U7081 ( .A1(n8561), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n6039) );
  NAND2_X1 U7082 ( .A1(n4854), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n6038) );
  NAND4_X1 U7083 ( .A1(n6041), .A2(n6040), .A3(n6039), .A4(n6038), .ZN(n9806)
         );
  INV_X1 U7084 ( .A(n9806), .ZN(n9769) );
  OAI22_X1 U7085 ( .A1(n9792), .A2(n6762), .B1(n9769), .B2(n6769), .ZN(n6064)
         );
  NAND2_X1 U7086 ( .A1(n10008), .A2(n6761), .ZN(n6043) );
  NAND2_X1 U7087 ( .A1(n9806), .A2(n4856), .ZN(n6042) );
  NAND2_X1 U7088 ( .A1(n6043), .A2(n6042), .ZN(n6044) );
  XNOR2_X1 U7089 ( .A(n6044), .B(n6081), .ZN(n6063) );
  XOR2_X1 U7090 ( .A(n6064), .B(n6063), .Z(n9344) );
  MUX2_X1 U7091 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(P2_DATAO_REG_26__SCAN_IN), 
        .S(n7142), .Z(n6070) );
  XNOR2_X1 U7092 ( .A(n6070), .B(n9133), .ZN(n6068) );
  XNOR2_X1 U7093 ( .A(n6069), .B(n6068), .ZN(n8465) );
  NAND2_X1 U7094 ( .A1(n8465), .A2(n8558), .ZN(n6049) );
  NAND2_X1 U7095 ( .A1(n6072), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n6048) );
  NAND2_X1 U7096 ( .A1(n10003), .A2(n6761), .ZN(n6059) );
  NAND2_X1 U7097 ( .A1(n4851), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n6057) );
  INV_X1 U7098 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n6051) );
  NAND2_X1 U7099 ( .A1(n6051), .A2(n6050), .ZN(n6053) );
  NAND2_X1 U7100 ( .A1(P1_REG3_REG_26__SCAN_IN), .A2(n6052), .ZN(n6135) );
  NAND2_X1 U7101 ( .A1(n4855), .A2(n9776), .ZN(n6056) );
  NAND2_X1 U7102 ( .A1(n8561), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n6055) );
  NAND2_X1 U7103 ( .A1(n4854), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n6054) );
  NAND4_X1 U7104 ( .A1(n6057), .A2(n6056), .A3(n6055), .A4(n6054), .ZN(n9785)
         );
  NAND2_X1 U7105 ( .A1(n9785), .A2(n5435), .ZN(n6058) );
  NAND2_X1 U7106 ( .A1(n6059), .A2(n6058), .ZN(n6060) );
  XNOR2_X1 U7107 ( .A(n6060), .B(n6081), .ZN(n6090) );
  AND2_X1 U7108 ( .A1(n9785), .A2(n6083), .ZN(n6061) );
  AOI21_X1 U7109 ( .B1(n10003), .B2(n5435), .A(n6061), .ZN(n6088) );
  XNOR2_X1 U7110 ( .A(n6090), .B(n6088), .ZN(n9414) );
  INV_X1 U7111 ( .A(n6063), .ZN(n6066) );
  INV_X1 U7112 ( .A(n6064), .ZN(n6065) );
  NAND2_X1 U7113 ( .A1(n6066), .A2(n6065), .ZN(n9410) );
  INV_X1 U7114 ( .A(n6070), .ZN(n6071) );
  MUX2_X1 U7115 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(P2_DATAO_REG_27__SCAN_IN), 
        .S(n7142), .Z(n6164) );
  INV_X1 U7116 ( .A(SI_27_), .ZN(n9130) );
  XNOR2_X1 U7117 ( .A(n6164), .B(n9130), .ZN(n6162) );
  XNOR2_X1 U7118 ( .A(n6163), .B(n6162), .ZN(n8499) );
  NAND2_X1 U7119 ( .A1(n8499), .A2(n8558), .ZN(n6074) );
  NAND2_X1 U7120 ( .A1(n6072), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n6073) );
  NAND2_X1 U7121 ( .A1(n9998), .A2(n6761), .ZN(n6080) );
  NAND2_X1 U7122 ( .A1(n4851), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n6078) );
  XNOR2_X1 U7123 ( .A(n6135), .B(P1_REG3_REG_27__SCAN_IN), .ZN(n6127) );
  NAND2_X1 U7124 ( .A1(n4855), .A2(n6127), .ZN(n6077) );
  NAND2_X1 U7125 ( .A1(n8561), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n6076) );
  NAND2_X1 U7126 ( .A1(n4854), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n6075) );
  NAND4_X1 U7127 ( .A1(n6078), .A2(n6077), .A3(n6076), .A4(n6075), .ZN(n9704)
         );
  NAND2_X1 U7128 ( .A1(n9704), .A2(n4856), .ZN(n6079) );
  NAND2_X1 U7129 ( .A1(n6080), .A2(n6079), .ZN(n6082) );
  XNOR2_X1 U7130 ( .A(n6082), .B(n6081), .ZN(n6087) );
  NAND2_X1 U7131 ( .A1(n9998), .A2(n5435), .ZN(n6085) );
  NAND2_X1 U7132 ( .A1(n9704), .A2(n6083), .ZN(n6084) );
  NAND2_X1 U7133 ( .A1(n6085), .A2(n6084), .ZN(n6086) );
  NOR2_X1 U7134 ( .A1(n6087), .A2(n6086), .ZN(n6775) );
  AOI21_X1 U7135 ( .B1(n6087), .B2(n6086), .A(n6775), .ZN(n6092) );
  INV_X1 U7136 ( .A(n6088), .ZN(n6089) );
  NAND2_X1 U7137 ( .A1(n6090), .A2(n6089), .ZN(n6093) );
  INV_X1 U7138 ( .A(n6786), .ZN(n6772) );
  AOI21_X1 U7139 ( .B1(n9412), .B2(n6093), .A(n6092), .ZN(n6119) );
  NAND2_X1 U7140 ( .A1(n6094), .A2(P1_B_REG_SCAN_IN), .ZN(n6095) );
  MUX2_X1 U7141 ( .A(P1_B_REG_SCAN_IN), .B(n6095), .S(n8404), .Z(n6097) );
  INV_X1 U7142 ( .A(n8404), .ZN(n6098) );
  NOR2_X1 U7143 ( .A1(n6096), .A2(n6098), .ZN(n6099) );
  INV_X1 U7144 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n10241) );
  INV_X1 U7145 ( .A(n6094), .ZN(n6101) );
  NOR2_X1 U7146 ( .A1(n6096), .A2(n6101), .ZN(n6102) );
  NOR2_X1 U7147 ( .A1(P1_D_REG_31__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .ZN(
        n6106) );
  NOR4_X1 U7148 ( .A1(P1_D_REG_4__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        P1_D_REG_29__SCAN_IN), .A4(P1_D_REG_28__SCAN_IN), .ZN(n6105) );
  NOR4_X1 U7149 ( .A1(P1_D_REG_23__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_21__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n6104) );
  NOR4_X1 U7150 ( .A1(P1_D_REG_27__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_25__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n6103) );
  NAND4_X1 U7151 ( .A1(n6106), .A2(n6105), .A3(n6104), .A4(n6103), .ZN(n6112)
         );
  NOR4_X1 U7152 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_13__SCAN_IN), .A4(P1_D_REG_12__SCAN_IN), .ZN(n6110) );
  NOR4_X1 U7153 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_18__SCAN_IN), .A4(P1_D_REG_16__SCAN_IN), .ZN(n6109) );
  NOR4_X1 U7154 ( .A1(P1_D_REG_7__SCAN_IN), .A2(P1_D_REG_6__SCAN_IN), .A3(
        P1_D_REG_5__SCAN_IN), .A4(P1_D_REG_2__SCAN_IN), .ZN(n6108) );
  NOR4_X1 U7155 ( .A1(P1_D_REG_11__SCAN_IN), .A2(P1_D_REG_10__SCAN_IN), .A3(
        P1_D_REG_9__SCAN_IN), .A4(P1_D_REG_8__SCAN_IN), .ZN(n6107) );
  NAND4_X1 U7156 ( .A1(n6110), .A2(n6109), .A3(n6108), .A4(n6107), .ZN(n6111)
         );
  OAI21_X1 U7157 ( .B1(n6112), .B2(n6111), .A(n10121), .ZN(n6202) );
  NAND3_X1 U7158 ( .A1(n10103), .A2(n6277), .A3(n6202), .ZN(n6123) );
  INV_X1 U7159 ( .A(n6113), .ZN(n6114) );
  NAND2_X1 U7160 ( .A1(n6114), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6116) );
  AND2_X1 U7161 ( .A1(n10520), .A2(n6117), .ZN(n6118) );
  INV_X1 U7162 ( .A(n9998), .ZN(n6142) );
  INV_X1 U7163 ( .A(n6128), .ZN(n6120) );
  OR2_X1 U7164 ( .A1(n7364), .A2(n8218), .ZN(n10406) );
  OR2_X1 U7165 ( .A1(n6120), .A2(n10406), .ZN(n6121) );
  NAND2_X1 U7166 ( .A1(n8515), .A2(n10411), .ZN(n9449) );
  INV_X1 U7167 ( .A(n6278), .ZN(n6122) );
  NAND2_X1 U7168 ( .A1(n6123), .A2(n6122), .ZN(n6126) );
  AND3_X1 U7169 ( .A1(n7209), .A2(n8397), .A3(n6201), .ZN(n6125) );
  NAND2_X1 U7170 ( .A1(n6126), .A2(n6125), .ZN(n7336) );
  INV_X1 U7171 ( .A(n6127), .ZN(n9757) );
  NOR2_X1 U7172 ( .A1(n9392), .A2(n9757), .ZN(n6140) );
  INV_X1 U7173 ( .A(n9785), .ZN(n6160) );
  INV_X1 U7174 ( .A(n9696), .ZN(n6252) );
  AND2_X1 U7175 ( .A1(n6128), .A2(n6252), .ZN(n6131) );
  INV_X1 U7176 ( .A(n6130), .ZN(n7621) );
  NAND2_X1 U7177 ( .A1(n6131), .A2(n6130), .ZN(n9430) );
  AOI22_X1 U7178 ( .A1(n4851), .A2(P1_REG1_REG_28__SCAN_IN), .B1(n8561), .B2(
        P1_REG0_REG_28__SCAN_IN), .ZN(n6138) );
  INV_X1 U7179 ( .A(n6135), .ZN(n6133) );
  AND2_X1 U7180 ( .A1(P1_REG3_REG_28__SCAN_IN), .A2(P1_REG3_REG_27__SCAN_IN), 
        .ZN(n6132) );
  NAND2_X1 U7181 ( .A1(n6133), .A2(n6132), .ZN(n6187) );
  INV_X1 U7182 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n6134) );
  INV_X1 U7183 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n6777) );
  OAI21_X1 U7184 ( .B1(n6135), .B2(n6134), .A(n6777), .ZN(n6136) );
  AOI22_X1 U7185 ( .A1(n4855), .A2(n8594), .B1(n4854), .B2(
        P1_REG2_REG_28__SCAN_IN), .ZN(n6137) );
  OAI22_X1 U7186 ( .A1(n6160), .A2(n9431), .B1(n9430), .B2(n9703), .ZN(n6139)
         );
  AOI211_X1 U7187 ( .C1(P1_REG3_REG_27__SCAN_IN), .C2(P1_U3084), .A(n6140), 
        .B(n6139), .ZN(n6141) );
  OAI21_X1 U7188 ( .B1(n6142), .B2(n9409), .A(n6141), .ZN(n6143) );
  NAND2_X1 U7189 ( .A1(n6145), .A2(n6144), .ZN(P1_U3212) );
  INV_X1 U7190 ( .A(n10385), .ZN(n7365) );
  INV_X1 U7191 ( .A(n9718), .ZN(n9592) );
  XNOR2_X1 U7192 ( .A(n10392), .B(n8590), .ZN(n9659) );
  INV_X1 U7193 ( .A(n10392), .ZN(n6208) );
  NAND2_X1 U7194 ( .A1(n6208), .A2(n8590), .ZN(n9594) );
  NAND2_X1 U7195 ( .A1(n6146), .A2(n9594), .ZN(n7727) );
  INV_X1 U7196 ( .A(n7776), .ZN(n7739) );
  NAND2_X1 U7197 ( .A1(n7727), .A2(n9598), .ZN(n6147) );
  INV_X1 U7198 ( .A(n9717), .ZN(n8580) );
  NAND2_X1 U7199 ( .A1(n9716), .A2(n4989), .ZN(n9623) );
  INV_X1 U7200 ( .A(n9714), .ZN(n7979) );
  NAND2_X1 U7201 ( .A1(n7979), .A2(n7952), .ZN(n9457) );
  INV_X1 U7202 ( .A(n9715), .ZN(n7945) );
  NAND2_X1 U7203 ( .A1(n7945), .A2(n8065), .ZN(n9455) );
  AND2_X1 U7204 ( .A1(n9457), .A2(n9455), .ZN(n9627) );
  NAND2_X1 U7205 ( .A1(n9450), .A2(n9627), .ZN(n6149) );
  INV_X1 U7206 ( .A(n8065), .ZN(n7936) );
  AND2_X1 U7207 ( .A1(n9715), .A2(n7936), .ZN(n6212) );
  NAND2_X1 U7208 ( .A1(n9457), .A2(n6212), .ZN(n9603) );
  INV_X1 U7209 ( .A(n7952), .ZN(n10467) );
  NAND2_X1 U7210 ( .A1(n9714), .A2(n10467), .ZN(n9454) );
  AND2_X1 U7211 ( .A1(n9603), .A2(n9454), .ZN(n6148) );
  NAND2_X1 U7212 ( .A1(n6149), .A2(n6148), .ZN(n8104) );
  INV_X1 U7213 ( .A(n9713), .ZN(n8020) );
  NAND2_X1 U7214 ( .A1(n8020), .A2(n8162), .ZN(n9536) );
  INV_X1 U7215 ( .A(n8162), .ZN(n8111) );
  NAND2_X1 U7216 ( .A1(n8111), .A2(n9713), .ZN(n9461) );
  NAND2_X1 U7217 ( .A1(n9536), .A2(n9461), .ZN(n8113) );
  INV_X1 U7218 ( .A(n8105), .ZN(n8184) );
  NAND2_X1 U7219 ( .A1(n8155), .A2(n8184), .ZN(n9537) );
  INV_X1 U7220 ( .A(n9536), .ZN(n9459) );
  OR2_X1 U7221 ( .A1(n10490), .A2(n8276), .ZN(n9545) );
  NAND2_X1 U7222 ( .A1(n10490), .A2(n8276), .ZN(n9468) );
  NAND2_X1 U7223 ( .A1(n9545), .A2(n9468), .ZN(n9664) );
  NAND2_X1 U7224 ( .A1(n8182), .A2(n9468), .ZN(n8274) );
  INV_X1 U7225 ( .A(n9711), .ZN(n8183) );
  OR2_X1 U7226 ( .A1(n10501), .A2(n8183), .ZN(n9547) );
  NAND2_X1 U7227 ( .A1(n10501), .A2(n8183), .ZN(n9534) );
  INV_X1 U7228 ( .A(n9534), .ZN(n9447) );
  OR2_X1 U7229 ( .A1(n9446), .A2(n8387), .ZN(n9550) );
  NAND2_X1 U7230 ( .A1(n9446), .A2(n8387), .ZN(n9533) );
  INV_X1 U7231 ( .A(n9709), .ZN(n6153) );
  AND2_X1 U7232 ( .A1(n9668), .A2(n9553), .ZN(n6152) );
  NAND2_X1 U7233 ( .A1(n8324), .A2(n6152), .ZN(n6156) );
  INV_X1 U7234 ( .A(n9553), .ZN(n9481) );
  INV_X1 U7235 ( .A(n9670), .ZN(n6154) );
  AND2_X1 U7236 ( .A1(n6154), .A2(n9550), .ZN(n8382) );
  NAND2_X1 U7237 ( .A1(n6156), .A2(n6155), .ZN(n8473) );
  INV_X1 U7239 ( .A(n9707), .ZN(n9948) );
  OR2_X1 U7240 ( .A1(n10068), .A2(n9948), .ZN(n9558) );
  NAND2_X1 U7241 ( .A1(n10068), .A2(n9948), .ZN(n9530) );
  NAND2_X1 U7242 ( .A1(n9558), .A2(n9530), .ZN(n9973) );
  INV_X1 U7243 ( .A(n9558), .ZN(n6158) );
  NAND2_X1 U7244 ( .A1(n9959), .A2(n9706), .ZN(n9559) );
  NAND2_X1 U7245 ( .A1(n10062), .A2(n9976), .ZN(n9922) );
  OR2_X1 U7246 ( .A1(n10058), .A2(n9947), .ZN(n9564) );
  NAND2_X1 U7247 ( .A1(n10058), .A2(n9947), .ZN(n9562) );
  NAND2_X1 U7248 ( .A1(n9564), .A2(n9562), .ZN(n9929) );
  INV_X1 U7249 ( .A(n9562), .ZN(n9905) );
  INV_X1 U7250 ( .A(n9899), .ZN(n9927) );
  OR2_X1 U7251 ( .A1(n10049), .A2(n9927), .ZN(n9568) );
  NAND2_X1 U7252 ( .A1(n10049), .A2(n9927), .ZN(n9567) );
  NAND2_X1 U7253 ( .A1(n9568), .A2(n9567), .ZN(n9908) );
  INV_X1 U7254 ( .A(n9568), .ZN(n9444) );
  OR2_X2 U7255 ( .A1(n9896), .A2(n9884), .ZN(n9571) );
  NAND2_X1 U7256 ( .A1(n9896), .A2(n9884), .ZN(n9569) );
  NAND2_X1 U7257 ( .A1(n9898), .A2(n5238), .ZN(n9897) );
  NAND2_X1 U7258 ( .A1(n9897), .A2(n9571), .ZN(n9881) );
  INV_X1 U7259 ( .A(n9900), .ZN(n9405) );
  OR2_X1 U7260 ( .A1(n10039), .A2(n9405), .ZN(n9573) );
  INV_X1 U7261 ( .A(n9883), .ZN(n9338) );
  OR2_X1 U7262 ( .A1(n10035), .A2(n9338), .ZN(n9495) );
  NAND2_X1 U7263 ( .A1(n10035), .A2(n9338), .ZN(n9496) );
  INV_X1 U7264 ( .A(n9870), .ZN(n9393) );
  OR2_X1 U7265 ( .A1(n10030), .A2(n9393), .ZN(n9498) );
  NAND2_X1 U7266 ( .A1(n10030), .A2(n9393), .ZN(n9499) );
  NAND2_X1 U7267 ( .A1(n9848), .A2(n9499), .ZN(n9830) );
  INV_X1 U7268 ( .A(n9851), .ZN(n9337) );
  OR2_X1 U7269 ( .A1(n9835), .A2(n9337), .ZN(n9579) );
  NAND2_X1 U7270 ( .A1(n9835), .A2(n9337), .ZN(n9575) );
  NAND2_X1 U7271 ( .A1(n9830), .A2(n9841), .ZN(n9829) );
  NAND2_X1 U7272 ( .A1(n9829), .A2(n9575), .ZN(n9822) );
  NAND2_X1 U7273 ( .A1(n9820), .A2(n9831), .ZN(n9581) );
  NAND2_X1 U7274 ( .A1(n9822), .A2(n9823), .ZN(n9821) );
  NAND2_X1 U7275 ( .A1(n9821), .A2(n9633), .ZN(n9804) );
  INV_X1 U7276 ( .A(n9824), .ZN(n9318) );
  OR2_X1 U7277 ( .A1(n10014), .A2(n9318), .ZN(n9631) );
  NAND2_X1 U7278 ( .A1(n10014), .A2(n9318), .ZN(n9606) );
  NAND2_X1 U7279 ( .A1(n9804), .A2(n9805), .ZN(n9803) );
  NAND2_X1 U7280 ( .A1(n9803), .A2(n9606), .ZN(n9784) );
  OR2_X1 U7281 ( .A1(n10008), .A2(n9769), .ZN(n9609) );
  NAND2_X1 U7282 ( .A1(n10008), .A2(n9769), .ZN(n9607) );
  NAND2_X1 U7283 ( .A1(n9784), .A2(n9796), .ZN(n9783) );
  NAND2_X1 U7284 ( .A1(n9783), .A2(n9607), .ZN(n9767) );
  OR2_X1 U7285 ( .A1(n10003), .A2(n6160), .ZN(n9610) );
  NAND2_X1 U7286 ( .A1(n10003), .A2(n6160), .ZN(n9747) );
  NAND2_X1 U7287 ( .A1(n9998), .A2(n9768), .ZN(n9615) );
  NAND2_X1 U7288 ( .A1(n9636), .A2(n9615), .ZN(n9754) );
  INV_X1 U7289 ( .A(n9747), .ZN(n9613) );
  NOR2_X1 U7290 ( .A1(n9754), .A2(n9613), .ZN(n6161) );
  NAND2_X1 U7291 ( .A1(n6163), .A2(n6162), .ZN(n6167) );
  INV_X1 U7292 ( .A(n6164), .ZN(n6165) );
  NAND2_X1 U7293 ( .A1(n6165), .A2(n9130), .ZN(n6166) );
  NAND2_X1 U7294 ( .A1(n6167), .A2(n6166), .ZN(n6169) );
  MUX2_X1 U7295 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(P2_DATAO_REG_28__SCAN_IN), 
        .S(n7142), .Z(n6173) );
  INV_X1 U7296 ( .A(SI_28_), .ZN(n9027) );
  XNOR2_X1 U7297 ( .A(n6173), .B(n9027), .ZN(n6168) );
  OR2_X1 U7298 ( .A1(n6169), .A2(n6168), .ZN(n6170) );
  NAND2_X1 U7299 ( .A1(n6176), .A2(n6170), .ZN(n10115) );
  NAND2_X1 U7300 ( .A1(n10115), .A2(n8558), .ZN(n6172) );
  INV_X1 U7301 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n10118) );
  OR2_X1 U7302 ( .A1(n5528), .A2(n10118), .ZN(n6171) );
  OR2_X1 U7303 ( .A1(n6781), .A2(n9703), .ZN(n9513) );
  NAND2_X1 U7304 ( .A1(n6781), .A2(n9703), .ZN(n9616) );
  INV_X1 U7305 ( .A(n6173), .ZN(n6174) );
  NAND2_X1 U7306 ( .A1(n6174), .A2(n9027), .ZN(n6175) );
  INV_X1 U7307 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n6177) );
  MUX2_X1 U7308 ( .A(n6177), .B(n6184), .S(n7142), .Z(n6178) );
  NAND2_X1 U7309 ( .A1(n6178), .A2(n9125), .ZN(n6825) );
  INV_X1 U7310 ( .A(n6178), .ZN(n6179) );
  NAND2_X1 U7311 ( .A1(n6179), .A2(SI_29_), .ZN(n6180) );
  OR2_X1 U7312 ( .A1(n6182), .A2(n6181), .ZN(n6183) );
  NAND2_X1 U7313 ( .A1(n6183), .A2(n6826), .ZN(n8518) );
  NAND2_X1 U7314 ( .A1(n8518), .A2(n8558), .ZN(n6186) );
  OR2_X1 U7315 ( .A1(n5528), .A2(n6184), .ZN(n6185) );
  AOI22_X1 U7316 ( .A1(n4851), .A2(P1_REG1_REG_29__SCAN_IN), .B1(n8561), .B2(
        P1_REG0_REG_29__SCAN_IN), .ZN(n6189) );
  INV_X1 U7317 ( .A(n6187), .ZN(n6256) );
  AOI22_X1 U7318 ( .A1(n4855), .A2(n6256), .B1(n4854), .B2(
        P1_REG2_REG_29__SCAN_IN), .ZN(n6188) );
  NAND2_X1 U7319 ( .A1(n9994), .A2(n7368), .ZN(n9643) );
  NAND2_X1 U7320 ( .A1(n9519), .A2(n9643), .ZN(n9650) );
  XNOR2_X1 U7321 ( .A(n6191), .B(n6190), .ZN(n6200) );
  OR2_X1 U7322 ( .A1(n8515), .A2(n9856), .ZN(n6192) );
  NAND2_X1 U7323 ( .A1(n9591), .A2(n9622), .ZN(n9442) );
  INV_X1 U7324 ( .A(n6117), .ZN(n6196) );
  NAND2_X1 U7325 ( .A1(n4850), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n6195) );
  NAND2_X1 U7326 ( .A1(n4854), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n6194) );
  NAND2_X1 U7327 ( .A1(n8561), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n6193) );
  INV_X1 U7328 ( .A(P1_B_REG_SCAN_IN), .ZN(n6197) );
  NOR2_X1 U7329 ( .A1(n9695), .A2(n6197), .ZN(n6198) );
  OR2_X1 U7330 ( .A1(n9975), .A2(n6198), .ZN(n8565) );
  OAI22_X1 U7331 ( .A1(n9703), .A2(n9977), .B1(n9618), .B2(n8565), .ZN(n6199)
         );
  INV_X1 U7332 ( .A(n10103), .ZN(n6281) );
  NAND2_X1 U7333 ( .A1(n6202), .A2(n6201), .ZN(n6279) );
  INV_X1 U7334 ( .A(n6279), .ZN(n6204) );
  NAND4_X1 U7335 ( .A1(n6281), .A2(n6204), .A3(n6203), .A4(n6277), .ZN(n7933)
         );
  AND2_X1 U7336 ( .A1(n6205), .A2(n10385), .ZN(n10384) );
  OAI21_X1 U7337 ( .B1(n9718), .B2(n10408), .A(n10384), .ZN(n6207) );
  NAND2_X1 U7338 ( .A1(n9718), .A2(n10408), .ZN(n6206) );
  AND2_X1 U7339 ( .A1(n6207), .A2(n6206), .ZN(n8572) );
  INV_X1 U7340 ( .A(n9659), .ZN(n8579) );
  INV_X1 U7341 ( .A(n8590), .ZN(n10420) );
  NAND2_X1 U7342 ( .A1(n6208), .A2(n10420), .ZN(n6209) );
  NAND2_X1 U7343 ( .A1(n8571), .A2(n6209), .ZN(n7730) );
  NAND2_X1 U7344 ( .A1(n8580), .A2(n7739), .ZN(n6210) );
  NAND2_X1 U7345 ( .A1(n7728), .A2(n6210), .ZN(n7872) );
  NAND2_X1 U7346 ( .A1(n5370), .A2(n9623), .ZN(n9651) );
  NAND2_X1 U7347 ( .A1(n7872), .A2(n9651), .ZN(n7871) );
  INV_X1 U7348 ( .A(n9716), .ZN(n7592) );
  NAND2_X1 U7349 ( .A1(n7592), .A2(n4989), .ZN(n6211) );
  INV_X1 U7350 ( .A(n6212), .ZN(n9624) );
  NAND2_X1 U7351 ( .A1(n9715), .A2(n8065), .ZN(n6214) );
  NAND2_X1 U7352 ( .A1(n8114), .A2(n8113), .ZN(n8112) );
  NAND2_X1 U7353 ( .A1(n8020), .A2(n8111), .ZN(n6215) );
  NAND2_X1 U7354 ( .A1(n8155), .A2(n8105), .ZN(n6216) );
  OR2_X1 U7355 ( .A1(n10490), .A2(n9712), .ZN(n6217) );
  NOR2_X1 U7356 ( .A1(n10501), .A2(n9711), .ZN(n6218) );
  OR2_X1 U7357 ( .A1(n9446), .A2(n9710), .ZN(n9475) );
  NAND2_X1 U7358 ( .A1(n8323), .A2(n9475), .ZN(n8381) );
  NAND2_X1 U7359 ( .A1(n9446), .A2(n9710), .ZN(n9474) );
  NAND2_X1 U7360 ( .A1(n10080), .A2(n9709), .ZN(n8468) );
  AND2_X1 U7361 ( .A1(n9474), .A2(n6219), .ZN(n6220) );
  NAND2_X1 U7362 ( .A1(n10068), .A2(n9707), .ZN(n6226) );
  AND2_X1 U7363 ( .A1(n6220), .A2(n6226), .ZN(n6221) );
  AND2_X2 U7364 ( .A1(n9559), .A2(n9922), .ZN(n9950) );
  INV_X1 U7365 ( .A(n9950), .ZN(n6227) );
  OR2_X1 U7366 ( .A1(n6222), .A2(n9670), .ZN(n6225) );
  OR2_X1 U7367 ( .A1(n6157), .A2(n9708), .ZN(n9962) );
  AND2_X1 U7368 ( .A1(n9962), .A2(n6223), .ZN(n6224) );
  AND2_X2 U7369 ( .A1(n6227), .A2(n9942), .ZN(n6228) );
  NAND2_X1 U7370 ( .A1(n10062), .A2(n9706), .ZN(n6229) );
  NAND2_X1 U7371 ( .A1(n10058), .A2(n9705), .ZN(n6230) );
  NAND2_X1 U7372 ( .A1(n9928), .A2(n6230), .ZN(n9909) );
  OR2_X1 U7373 ( .A1(n10049), .A2(n9899), .ZN(n6231) );
  NAND2_X1 U7374 ( .A1(n9909), .A2(n6231), .ZN(n6233) );
  NAND2_X1 U7375 ( .A1(n10049), .A2(n9899), .ZN(n6232) );
  NAND2_X1 U7376 ( .A1(n10039), .A2(n9900), .ZN(n6235) );
  NAND2_X1 U7377 ( .A1(n6236), .A2(n6235), .ZN(n9861) );
  OR2_X1 U7378 ( .A1(n10035), .A2(n9883), .ZN(n6237) );
  NAND2_X1 U7379 ( .A1(n9861), .A2(n6237), .ZN(n6239) );
  NAND2_X1 U7380 ( .A1(n10035), .A2(n9883), .ZN(n6238) );
  NAND2_X1 U7381 ( .A1(n10030), .A2(n9870), .ZN(n6240) );
  OR2_X1 U7382 ( .A1(n9835), .A2(n9851), .ZN(n6242) );
  OR2_X1 U7383 ( .A1(n9820), .A2(n9394), .ZN(n6243) );
  NAND2_X1 U7384 ( .A1(n10014), .A2(n9824), .ZN(n6244) );
  OR2_X1 U7385 ( .A1(n10008), .A2(n9806), .ZN(n6246) );
  INV_X1 U7386 ( .A(n9771), .ZN(n6247) );
  NAND2_X1 U7387 ( .A1(n10003), .A2(n9785), .ZN(n6248) );
  OR2_X1 U7388 ( .A1(n6765), .A2(n6252), .ZN(n6253) );
  INV_X1 U7389 ( .A(n10035), .ZN(n9866) );
  INV_X1 U7390 ( .A(n10058), .ZN(n9934) );
  NAND2_X1 U7391 ( .A1(n10388), .A2(n10420), .ZN(n8576) );
  OR2_X1 U7392 ( .A1(n8576), .A2(n7776), .ZN(n7873) );
  INV_X1 U7393 ( .A(n10501), .ZN(n8282) );
  INV_X1 U7394 ( .A(n9446), .ZN(n10521) );
  INV_X1 U7395 ( .A(n10080), .ZN(n8393) );
  NAND2_X1 U7396 ( .A1(n8388), .A2(n8393), .ZN(n8477) );
  NAND2_X1 U7397 ( .A1(n9820), .A2(n9833), .ZN(n9816) );
  NAND2_X1 U7398 ( .A1(n9792), .A2(n9808), .ZN(n9789) );
  INV_X1 U7399 ( .A(n6273), .ZN(n6254) );
  INV_X1 U7400 ( .A(n9994), .ZN(n6258) );
  AOI21_X1 U7401 ( .B1(n9994), .B2(n6254), .A(n9741), .ZN(n9995) );
  INV_X2 U7402 ( .A(n9940), .ZN(n10371) );
  OR2_X1 U7403 ( .A1(n7364), .A2(n9693), .ZN(n6255) );
  NOR2_X2 U7404 ( .A1(n10371), .A2(n6255), .ZN(n10368) );
  AOI22_X1 U7405 ( .A1(n10371), .A2(P1_REG2_REG_29__SCAN_IN), .B1(n6256), .B2(
        n10409), .ZN(n6257) );
  OAI21_X1 U7406 ( .B1(n6258), .B2(n9969), .A(n6257), .ZN(n6259) );
  NAND2_X1 U7407 ( .A1(n6263), .A2(n9678), .ZN(n6264) );
  OAI21_X1 U7408 ( .B1(n9678), .B2(n6268), .A(n6267), .ZN(n6269) );
  OAI22_X1 U7409 ( .A1(n9768), .A2(n9977), .B1(n7368), .B2(n9975), .ZN(n6270)
         );
  AOI21_X1 U7410 ( .B1(n6781), .B2(n9761), .A(n6273), .ZN(n8599) );
  AOI22_X1 U7411 ( .A1(n8599), .A2(n10386), .B1(n10502), .B2(n6781), .ZN(n6274) );
  NOR2_X1 U7412 ( .A1(n6277), .A2(n10242), .ZN(n10240) );
  NOR2_X1 U7413 ( .A1(n6279), .A2(n6278), .ZN(n6280) );
  INV_X1 U7414 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n6282) );
  AND2_X1 U7415 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n6383) );
  NAND2_X1 U7416 ( .A1(n6383), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n6410) );
  NOR2_X1 U7417 ( .A1(n6410), .A2(n9222), .ZN(n6409) );
  NAND2_X1 U7418 ( .A1(n6409), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n6435) );
  NOR2_X1 U7419 ( .A1(n6450), .A2(n6449), .ZN(n6448) );
  NAND2_X1 U7420 ( .A1(n6466), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6496) );
  NAND2_X1 U7421 ( .A1(n6521), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n6552) );
  INV_X1 U7422 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n8638) );
  NAND2_X1 U7423 ( .A1(n6619), .A2(n8638), .ZN(n6285) );
  NAND2_X1 U7424 ( .A1(n6629), .A2(n6285), .ZN(n8836) );
  NOR2_X1 U7425 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .ZN(
        n6291) );
  NAND4_X1 U7426 ( .A1(n6291), .A2(n6290), .A3(n6289), .A4(n6288), .ZN(n6294)
         );
  INV_X2 U7427 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n6489) );
  INV_X2 U7428 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n6488) );
  NAND4_X1 U7429 ( .A1(n6489), .A2(n6516), .A3(n6488), .A4(n6292), .ZN(n6293)
         );
  NOR2_X1 U7430 ( .A1(n6294), .A2(n6293), .ZN(n6295) );
  NAND2_X1 U7431 ( .A1(n6377), .A2(n6295), .ZN(n6545) );
  NAND2_X1 U7432 ( .A1(n6700), .A2(n6581), .ZN(n6666) );
  INV_X1 U7433 ( .A(n6666), .ZN(n6299) );
  INV_X1 U7434 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n6296) );
  INV_X2 U7435 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n6706) );
  NOR2_X1 U7436 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(P2_IR_REG_26__SCAN_IN), .ZN(
        n6298) );
  NOR2_X1 U7437 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), .ZN(
        n6297) );
  NOR2_X2 U7438 ( .A1(n6314), .A2(P2_IR_REG_28__SCAN_IN), .ZN(n6302) );
  NAND2_X1 U7439 ( .A1(n6302), .A2(n6303), .ZN(n9295) );
  XNOR2_X2 U7440 ( .A(n6304), .B(n6303), .ZN(n8519) );
  NAND2_X2 U7441 ( .A1(n6305), .A2(n6306), .ZN(n6384) );
  OR2_X1 U7442 ( .A1(n8836), .A2(n6384), .ZN(n6313) );
  INV_X1 U7443 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n6310) );
  NAND2_X4 U7444 ( .A1(n9299), .A2(n6306), .ZN(n6744) );
  INV_X2 U7445 ( .A(n6433), .ZN(n6796) );
  NAND2_X1 U7446 ( .A1(n6796), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n6309) );
  NAND2_X2 U7447 ( .A1(n6307), .A2(n8519), .ZN(n6395) );
  INV_X4 U7448 ( .A(n6395), .ZN(n6821) );
  NAND2_X1 U7449 ( .A1(n6821), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n6308) );
  OAI211_X1 U7450 ( .C1(n6310), .C2(n6744), .A(n6309), .B(n6308), .ZN(n6311)
         );
  INV_X1 U7451 ( .A(n6311), .ZN(n6312) );
  NAND2_X1 U7452 ( .A1(n6313), .A2(n6312), .ZN(n8843) );
  MUX2_X1 U7453 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6317), .S(
        P2_IR_REG_27__SCAN_IN), .Z(n6318) );
  INV_X2 U7455 ( .A(n6537), .ZN(n6833) );
  NAND2_X1 U7456 ( .A1(n8402), .A2(n6833), .ZN(n6320) );
  NAND2_X1 U7457 ( .A1(n6820), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n6319) );
  INV_X1 U7458 ( .A(n6321), .ZN(n6607) );
  NAND2_X1 U7459 ( .A1(n6599), .A2(n9084), .ZN(n6322) );
  NAND2_X1 U7460 ( .A1(n6607), .A2(n6322), .ZN(n8876) );
  OR2_X1 U7461 ( .A1(n8876), .A2(n6384), .ZN(n6328) );
  INV_X1 U7462 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n6325) );
  NAND2_X1 U7463 ( .A1(n6796), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n6324) );
  NAND2_X1 U7464 ( .A1(n6821), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n6323) );
  OAI211_X1 U7465 ( .C1(n6325), .C2(n6744), .A(n6324), .B(n6323), .ZN(n6326)
         );
  INV_X1 U7466 ( .A(n6326), .ZN(n6327) );
  NAND2_X1 U7467 ( .A1(n6328), .A2(n6327), .ZN(n8887) );
  INV_X1 U7468 ( .A(n8887), .ZN(n8659) );
  OR2_X1 U7469 ( .A1(n8220), .A2(n6537), .ZN(n6330) );
  NAND2_X1 U7470 ( .A1(n6820), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n6329) );
  NAND2_X1 U7471 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n6331) );
  INV_X1 U7472 ( .A(n10349), .ZN(n6332) );
  INV_X1 U7473 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n6334) );
  NAND2_X1 U7474 ( .A1(n6821), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n6336) );
  NAND2_X1 U7475 ( .A1(n6382), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n6335) );
  INV_X1 U7476 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n7653) );
  OR2_X1 U7477 ( .A1(n6384), .A2(n7653), .ZN(n6337) );
  NAND2_X1 U7478 ( .A1(n7231), .A2(n8699), .ZN(n6718) );
  INV_X1 U7479 ( .A(n6340), .ZN(n7045) );
  NAND2_X1 U7480 ( .A1(n7045), .A2(n7658), .ZN(n6717) );
  NAND2_X1 U7481 ( .A1(n6718), .A2(n6717), .ZN(n6839) );
  NAND2_X1 U7482 ( .A1(n6382), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n6346) );
  INV_X1 U7483 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n7294) );
  INV_X1 U7484 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n6341) );
  OR2_X1 U7485 ( .A1(n6395), .A2(n6341), .ZN(n6344) );
  INV_X1 U7486 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n6342) );
  OR2_X1 U7487 ( .A1(n6744), .A2(n6342), .ZN(n6343) );
  INV_X1 U7488 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n6349) );
  NOR2_X1 U7489 ( .A1(n7142), .A2(n9173), .ZN(n6347) );
  XNOR2_X1 U7490 ( .A(n6347), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n9302) );
  MUX2_X1 U7491 ( .A(n6349), .B(n9302), .S(n6348), .Z(n7050) );
  INV_X1 U7492 ( .A(n7050), .ZN(n10377) );
  AND2_X1 U7493 ( .A1(n8700), .A2(n10377), .ZN(n7226) );
  NAND2_X1 U7494 ( .A1(n6839), .A2(n7226), .ZN(n7228) );
  OR2_X1 U7495 ( .A1(n7045), .A2(n7231), .ZN(n6350) );
  NAND2_X1 U7496 ( .A1(n7228), .A2(n6350), .ZN(n7827) );
  INV_X1 U7497 ( .A(n7827), .ZN(n6363) );
  INV_X1 U7498 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n9219) );
  OR2_X1 U7499 ( .A1(n6384), .A2(n9219), .ZN(n6354) );
  INV_X1 U7500 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n6351) );
  OR2_X1 U7501 ( .A1(n6433), .A2(n6351), .ZN(n6353) );
  NAND2_X1 U7502 ( .A1(n6821), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6352) );
  INV_X1 U7503 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n7379) );
  OR2_X1 U7504 ( .A1(n6744), .A2(n7379), .ZN(n6355) );
  NAND2_X1 U7505 ( .A1(n4871), .A2(n6355), .ZN(n7332) );
  INV_X1 U7506 ( .A(n7332), .ZN(n7472) );
  INV_X1 U7507 ( .A(n6356), .ZN(n6357) );
  NAND2_X1 U7508 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n6357), .ZN(n6358) );
  MUX2_X1 U7509 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6358), .S(
        P2_IR_REG_2__SCAN_IN), .Z(n6360) );
  INV_X1 U7510 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n6359) );
  NAND2_X1 U7511 ( .A1(n6359), .A2(n6356), .ZN(n6369) );
  NAND2_X1 U7512 ( .A1(n6360), .A2(n6369), .ZN(n7389) );
  OR2_X1 U7513 ( .A1(n6537), .A2(n7149), .ZN(n6362) );
  NAND2_X1 U7514 ( .A1(n6379), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n6361) );
  OAI211_X1 U7515 ( .C1(n6348), .C2(n7389), .A(n6362), .B(n6361), .ZN(n7054)
         );
  INV_X1 U7516 ( .A(n7054), .ZN(n6364) );
  NAND2_X1 U7517 ( .A1(n6364), .A2(n7332), .ZN(n6869) );
  NAND2_X1 U7518 ( .A1(n6720), .A2(n6869), .ZN(n7826) );
  NAND2_X1 U7519 ( .A1(n6363), .A2(n7826), .ZN(n7468) );
  NAND2_X1 U7520 ( .A1(n7472), .A2(n6364), .ZN(n7469) );
  INV_X1 U7521 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n7380) );
  INV_X1 U7522 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n7667) );
  NAND2_X1 U7523 ( .A1(n6382), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n6365) );
  OR2_X1 U7524 ( .A1(n7146), .A2(n6537), .ZN(n6371) );
  NAND2_X1 U7525 ( .A1(n6369), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6370) );
  XNOR2_X1 U7526 ( .A(n6370), .B(P2_IR_REG_3__SCAN_IN), .ZN(n7441) );
  INV_X1 U7527 ( .A(n7665), .ZN(n7310) );
  NAND2_X1 U7528 ( .A1(n7830), .A2(n7310), .ZN(n6373) );
  AND2_X1 U7529 ( .A1(n7469), .A2(n6373), .ZN(n6372) );
  NAND2_X1 U7530 ( .A1(n7468), .A2(n6372), .ZN(n7764) );
  INV_X1 U7531 ( .A(n6373), .ZN(n6374) );
  INV_X1 U7532 ( .A(n7830), .ZN(n7296) );
  OR2_X1 U7533 ( .A1(n6374), .A2(n6721), .ZN(n7763) );
  OR2_X1 U7534 ( .A1(n7147), .A2(n6537), .ZN(n6381) );
  NOR2_X1 U7535 ( .A1(n6375), .A2(n9294), .ZN(n6376) );
  MUX2_X1 U7536 ( .A(n9294), .B(n6376), .S(P2_IR_REG_4__SCAN_IN), .Z(n6378) );
  NOR2_X1 U7537 ( .A1(n6378), .A2(n6377), .ZN(n7414) );
  AOI22_X1 U7538 ( .A1(n6379), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n7304), .B2(
        n7414), .ZN(n6380) );
  NAND2_X1 U7539 ( .A1(n6381), .A2(n6380), .ZN(n7768) );
  NAND2_X1 U7540 ( .A1(n6796), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n6389) );
  INV_X1 U7541 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n7756) );
  OR2_X1 U7542 ( .A1(n6395), .A2(n7756), .ZN(n6388) );
  INV_X1 U7543 ( .A(n6383), .ZN(n6397) );
  OAI21_X1 U7544 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(P2_REG3_REG_3__SCAN_IN), 
        .A(n6397), .ZN(n7760) );
  OR2_X1 U7545 ( .A1(n6384), .A2(n7760), .ZN(n6387) );
  INV_X1 U7546 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6385) );
  OR2_X1 U7547 ( .A1(n6744), .A2(n6385), .ZN(n6386) );
  NAND2_X1 U7548 ( .A1(n7768), .A2(n8698), .ZN(n6878) );
  AND2_X1 U7549 ( .A1(n7763), .A2(n6878), .ZN(n6391) );
  INV_X1 U7550 ( .A(n6881), .ZN(n6390) );
  NAND2_X2 U7551 ( .A1(n6390), .A2(n6878), .ZN(n7767) );
  OR2_X1 U7552 ( .A1(n7153), .A2(n6537), .ZN(n6394) );
  OR2_X1 U7553 ( .A1(n6377), .A2(n9294), .ZN(n6392) );
  XNOR2_X1 U7554 ( .A(n6392), .B(P2_IR_REG_5__SCAN_IN), .ZN(n7427) );
  AOI22_X1 U7555 ( .A1(n6834), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n7304), .B2(
        n7427), .ZN(n6393) );
  NAND2_X1 U7556 ( .A1(n6382), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n6403) );
  INV_X1 U7557 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n6396) );
  OR2_X1 U7558 ( .A1(n6395), .A2(n6396), .ZN(n6402) );
  INV_X1 U7559 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n9092) );
  NAND2_X1 U7560 ( .A1(n6397), .A2(n9092), .ZN(n6398) );
  NAND2_X1 U7561 ( .A1(n6410), .A2(n6398), .ZN(n10453) );
  OR2_X1 U7562 ( .A1(n6384), .A2(n10453), .ZN(n6401) );
  INV_X1 U7563 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n6399) );
  OR2_X1 U7564 ( .A1(n6744), .A2(n6399), .ZN(n6400) );
  NAND4_X1 U7565 ( .A1(n6403), .A2(n6402), .A3(n6401), .A4(n6400), .ZN(n8697)
         );
  INV_X1 U7566 ( .A(n8697), .ZN(n7675) );
  NOR2_X1 U7567 ( .A1(n10456), .A2(n7675), .ZN(n6404) );
  INV_X1 U7568 ( .A(n10456), .ZN(n7355) );
  OAI22_X1 U7569 ( .A1(n7688), .A2(n6404), .B1(n7355), .B2(n8697), .ZN(n7671)
         );
  OR2_X1 U7570 ( .A1(n7156), .A2(n6537), .ZN(n6408) );
  INV_X1 U7571 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n6405) );
  NAND2_X1 U7572 ( .A1(n6377), .A2(n6405), .ZN(n6418) );
  NAND2_X1 U7573 ( .A1(n6418), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6406) );
  XNOR2_X1 U7574 ( .A(n6406), .B(P2_IR_REG_6__SCAN_IN), .ZN(n7452) );
  AOI22_X1 U7575 ( .A1(n6834), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n7304), .B2(
        n7452), .ZN(n6407) );
  NAND2_X1 U7576 ( .A1(n6408), .A2(n6407), .ZN(n7681) );
  NAND2_X1 U7577 ( .A1(n6796), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n6416) );
  INV_X1 U7578 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n7393) );
  OR2_X1 U7579 ( .A1(n6395), .A2(n7393), .ZN(n6415) );
  INV_X1 U7580 ( .A(n6409), .ZN(n6422) );
  NAND2_X1 U7581 ( .A1(n6410), .A2(n9222), .ZN(n6411) );
  NAND2_X1 U7582 ( .A1(n6422), .A2(n6411), .ZN(n7678) );
  OR2_X1 U7583 ( .A1(n6384), .A2(n7678), .ZN(n6414) );
  INV_X1 U7584 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n6412) );
  OR2_X1 U7585 ( .A1(n6744), .A2(n6412), .ZN(n6413) );
  NAND2_X1 U7586 ( .A1(n7681), .A2(n7789), .ZN(n6417) );
  OR2_X1 U7587 ( .A1(n7159), .A2(n6537), .ZN(n6421) );
  NAND2_X1 U7588 ( .A1(n6429), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6419) );
  XNOR2_X1 U7589 ( .A(n6419), .B(P2_IR_REG_7__SCAN_IN), .ZN(n7513) );
  AOI22_X1 U7590 ( .A1(n6834), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n7304), .B2(
        n7513), .ZN(n6420) );
  NAND2_X1 U7591 ( .A1(n6421), .A2(n6420), .ZN(n7859) );
  NAND2_X1 U7592 ( .A1(n6796), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n6428) );
  INV_X1 U7593 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n7792) );
  OR2_X1 U7594 ( .A1(n6395), .A2(n7792), .ZN(n6427) );
  INV_X1 U7595 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n7580) );
  NAND2_X1 U7596 ( .A1(n6422), .A2(n7580), .ZN(n6423) );
  NAND2_X1 U7597 ( .A1(n6435), .A2(n6423), .ZN(n7791) );
  OR2_X1 U7598 ( .A1(n6384), .A2(n7791), .ZN(n6426) );
  INV_X1 U7599 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n6424) );
  OR2_X1 U7600 ( .A1(n6744), .A2(n6424), .ZN(n6425) );
  OR2_X1 U7601 ( .A1(n7859), .A2(n7719), .ZN(n6897) );
  NAND2_X1 U7602 ( .A1(n7859), .A2(n7719), .ZN(n6896) );
  NAND2_X1 U7603 ( .A1(n6897), .A2(n6896), .ZN(n7785) );
  INV_X1 U7604 ( .A(n7785), .ZN(n7787) );
  INV_X1 U7605 ( .A(n7719), .ZN(n8696) );
  NAND2_X1 U7606 ( .A1(n7161), .A2(n6833), .ZN(n6432) );
  NOR2_X1 U7607 ( .A1(n6429), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n6445) );
  OR2_X1 U7608 ( .A1(n6445), .A2(n9294), .ZN(n6430) );
  XNOR2_X1 U7609 ( .A(n6430), .B(P2_IR_REG_8__SCAN_IN), .ZN(n7520) );
  AOI22_X1 U7610 ( .A1(n6834), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n7304), .B2(
        n7520), .ZN(n6431) );
  NAND2_X1 U7611 ( .A1(n6432), .A2(n6431), .ZN(n7849) );
  NAND2_X1 U7612 ( .A1(n6796), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n6441) );
  INV_X1 U7613 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7852) );
  OR2_X1 U7614 ( .A1(n6395), .A2(n7852), .ZN(n6440) );
  NAND2_X1 U7615 ( .A1(n6435), .A2(n6434), .ZN(n6436) );
  NAND2_X1 U7616 ( .A1(n6450), .A2(n6436), .ZN(n7851) );
  OR2_X1 U7617 ( .A1(n6384), .A2(n7851), .ZN(n6439) );
  INV_X1 U7618 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n6437) );
  OR2_X1 U7619 ( .A1(n6744), .A2(n6437), .ZN(n6438) );
  NAND4_X1 U7620 ( .A1(n6441), .A2(n6440), .A3(n6439), .A4(n6438), .ZN(n8694)
         );
  XNOR2_X1 U7621 ( .A(n7849), .B(n8694), .ZN(n7805) );
  NAND2_X1 U7622 ( .A1(n7849), .A2(n8694), .ZN(n6443) );
  NAND2_X1 U7623 ( .A1(n7804), .A2(n6443), .ZN(n8048) );
  INV_X1 U7624 ( .A(n8048), .ZN(n6458) );
  NAND2_X1 U7625 ( .A1(n7169), .A2(n6833), .ZN(n6447) );
  INV_X1 U7626 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n6444) );
  NAND2_X1 U7627 ( .A1(n6445), .A2(n6444), .ZN(n6491) );
  NAND2_X1 U7628 ( .A1(n6491), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6460) );
  XNOR2_X1 U7629 ( .A(n6460), .B(n6489), .ZN(n7521) );
  INV_X1 U7630 ( .A(n7521), .ZN(n7538) );
  AOI22_X1 U7631 ( .A1(n6834), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n7304), .B2(
        n7538), .ZN(n6446) );
  NAND2_X1 U7632 ( .A1(n6447), .A2(n6446), .ZN(n8196) );
  NAND2_X1 U7633 ( .A1(n6796), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n6456) );
  INV_X1 U7634 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n8058) );
  OR2_X1 U7635 ( .A1(n6395), .A2(n8058), .ZN(n6455) );
  INV_X1 U7636 ( .A(n6448), .ZN(n6468) );
  NAND2_X1 U7637 ( .A1(n6450), .A2(n6449), .ZN(n6451) );
  NAND2_X1 U7638 ( .A1(n6468), .A2(n6451), .ZN(n8057) );
  OR2_X1 U7639 ( .A1(n6384), .A2(n8057), .ZN(n6454) );
  INV_X1 U7640 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n6452) );
  OR2_X1 U7641 ( .A1(n6744), .A2(n6452), .ZN(n6453) );
  NOR2_X1 U7642 ( .A1(n8196), .A2(n7902), .ZN(n6864) );
  INV_X1 U7643 ( .A(n6864), .ZN(n6900) );
  NAND2_X1 U7644 ( .A1(n8196), .A2(n7902), .ZN(n6902) );
  NAND2_X1 U7645 ( .A1(n6458), .A2(n6457), .ZN(n8046) );
  INV_X1 U7646 ( .A(n7902), .ZN(n8693) );
  OR2_X1 U7647 ( .A1(n8196), .A2(n8693), .ZN(n6459) );
  NAND2_X1 U7648 ( .A1(n7175), .A2(n6833), .ZN(n6465) );
  NAND2_X1 U7649 ( .A1(n6460), .A2(n6489), .ZN(n6461) );
  NAND2_X1 U7650 ( .A1(n6461), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6462) );
  NAND2_X1 U7651 ( .A1(n6462), .A2(n6488), .ZN(n6476) );
  OR2_X1 U7652 ( .A1(n6462), .A2(n6488), .ZN(n6463) );
  AOI22_X1 U7653 ( .A1(n6834), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n7602), .B2(
        n7304), .ZN(n6464) );
  NAND2_X1 U7654 ( .A1(n6465), .A2(n6464), .ZN(n10512) );
  INV_X1 U7655 ( .A(n6744), .ZN(n6795) );
  NAND2_X1 U7656 ( .A1(n6795), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n6474) );
  INV_X1 U7657 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7993) );
  OR2_X1 U7658 ( .A1(n6395), .A2(n7993), .ZN(n6473) );
  INV_X1 U7659 ( .A(n6466), .ZN(n6481) );
  INV_X1 U7660 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n6467) );
  NAND2_X1 U7661 ( .A1(n6468), .A2(n6467), .ZN(n6469) );
  NAND2_X1 U7662 ( .A1(n6481), .A2(n6469), .ZN(n7992) );
  OR2_X1 U7663 ( .A1(n6384), .A2(n7992), .ZN(n6472) );
  INV_X1 U7664 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n6470) );
  OR2_X1 U7665 ( .A1(n6433), .A2(n6470), .ZN(n6471) );
  OR2_X1 U7666 ( .A1(n10512), .A2(n7922), .ZN(n6911) );
  NAND2_X1 U7667 ( .A1(n10512), .A2(n7922), .ZN(n6909) );
  NAND2_X1 U7668 ( .A1(n6911), .A2(n6909), .ZN(n7988) );
  INV_X1 U7669 ( .A(n7922), .ZN(n8692) );
  NAND2_X1 U7670 ( .A1(n10512), .A2(n8692), .ZN(n6475) );
  OR2_X1 U7671 ( .A1(n7180), .A2(n6537), .ZN(n6479) );
  NAND2_X1 U7672 ( .A1(n6476), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6477) );
  XNOR2_X1 U7673 ( .A(n6477), .B(P2_IR_REG_11__SCAN_IN), .ZN(n7892) );
  AOI22_X1 U7674 ( .A1(n7892), .A2(n7304), .B1(n6834), .B2(
        P1_DATAO_REG_11__SCAN_IN), .ZN(n6478) );
  NAND2_X1 U7675 ( .A1(n6479), .A2(n6478), .ZN(n8098) );
  NAND2_X1 U7676 ( .A1(n6796), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n6486) );
  INV_X1 U7677 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n6480) );
  OR2_X1 U7678 ( .A1(n6395), .A2(n6480), .ZN(n6485) );
  INV_X1 U7679 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n9215) );
  NAND2_X1 U7680 ( .A1(n6481), .A2(n9215), .ZN(n6482) );
  NAND2_X1 U7681 ( .A1(n6496), .A2(n6482), .ZN(n8171) );
  OR2_X1 U7682 ( .A1(n6384), .A2(n8171), .ZN(n6484) );
  INV_X1 U7683 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n7603) );
  OR2_X1 U7684 ( .A1(n6744), .A2(n7603), .ZN(n6483) );
  OR2_X1 U7685 ( .A1(n8098), .A2(n8130), .ZN(n6912) );
  AND2_X1 U7686 ( .A1(n8098), .A2(n8130), .ZN(n6857) );
  INV_X1 U7687 ( .A(n6857), .ZN(n6910) );
  INV_X1 U7688 ( .A(n8091), .ZN(n8089) );
  INV_X1 U7689 ( .A(n8130), .ZN(n7986) );
  INV_X1 U7690 ( .A(n8131), .ZN(n6502) );
  INV_X1 U7691 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n6487) );
  NAND3_X1 U7692 ( .A1(n6489), .A2(n6488), .A3(n6487), .ZN(n6490) );
  NAND2_X1 U7693 ( .A1(n6503), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6492) );
  XNOR2_X1 U7694 ( .A(n6492), .B(P2_IR_REG_12__SCAN_IN), .ZN(n7964) );
  AOI22_X1 U7695 ( .A1(n6834), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n7304), .B2(
        n7964), .ZN(n6493) );
  NAND2_X1 U7696 ( .A1(n6796), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n6501) );
  INV_X1 U7697 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n8137) );
  OR2_X1 U7698 ( .A1(n6395), .A2(n8137), .ZN(n6500) );
  NAND2_X1 U7699 ( .A1(n6496), .A2(n6495), .ZN(n6497) );
  NAND2_X1 U7700 ( .A1(n6506), .A2(n6497), .ZN(n8136) );
  OR2_X1 U7701 ( .A1(n6384), .A2(n8136), .ZN(n6499) );
  INV_X1 U7702 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n7884) );
  OR2_X1 U7703 ( .A1(n6744), .A2(n7884), .ZN(n6498) );
  INV_X1 U7704 ( .A(n8211), .ZN(n8244) );
  NAND2_X1 U7705 ( .A1(n7543), .A2(n6833), .ZN(n6505) );
  OAI21_X1 U7706 ( .B1(n6503), .B2(P2_IR_REG_12__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n6514) );
  XNOR2_X1 U7707 ( .A(n6514), .B(P2_IR_REG_13__SCAN_IN), .ZN(n8037) );
  AOI22_X1 U7708 ( .A1(n7304), .A2(n8037), .B1(n6834), .B2(
        P1_DATAO_REG_13__SCAN_IN), .ZN(n6504) );
  NAND2_X1 U7709 ( .A1(n6796), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n6512) );
  INV_X1 U7710 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n8239) );
  OR2_X1 U7711 ( .A1(n6395), .A2(n8239), .ZN(n6511) );
  NAND2_X1 U7712 ( .A1(n6506), .A2(n9210), .ZN(n6507) );
  NAND2_X1 U7713 ( .A1(n6523), .A2(n6507), .ZN(n8238) );
  OR2_X1 U7714 ( .A1(n6384), .A2(n8238), .ZN(n6510) );
  INV_X1 U7715 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n6508) );
  OR2_X1 U7716 ( .A1(n6744), .A2(n6508), .ZN(n6509) );
  NAND4_X1 U7717 ( .A1(n6512), .A2(n6511), .A3(n6510), .A4(n6509), .ZN(n8691)
         );
  INV_X1 U7718 ( .A(n8242), .ZN(n8235) );
  INV_X1 U7719 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n6513) );
  NAND2_X1 U7720 ( .A1(n6514), .A2(n6513), .ZN(n6515) );
  NAND2_X1 U7721 ( .A1(n6515), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6517) );
  NAND2_X1 U7722 ( .A1(n6517), .A2(n6516), .ZN(n6531) );
  OR2_X1 U7723 ( .A1(n6517), .A2(n6516), .ZN(n6518) );
  AOI22_X1 U7724 ( .A1(n8312), .A2(n7304), .B1(n6834), .B2(
        P1_DATAO_REG_14__SCAN_IN), .ZN(n6519) );
  INV_X1 U7725 ( .A(n6521), .ZN(n6539) );
  NAND2_X1 U7726 ( .A1(n6523), .A2(n6522), .ZN(n6524) );
  NAND2_X1 U7727 ( .A1(n6539), .A2(n6524), .ZN(n8337) );
  OR2_X1 U7728 ( .A1(n6384), .A2(n8337), .ZN(n6530) );
  INV_X1 U7729 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n6525) );
  OR2_X1 U7730 ( .A1(n6433), .A2(n6525), .ZN(n6529) );
  INV_X1 U7731 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n6526) );
  OR2_X1 U7732 ( .A1(n6395), .A2(n6526), .ZN(n6528) );
  INV_X1 U7733 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n8029) );
  OR2_X1 U7734 ( .A1(n6744), .A2(n8029), .ZN(n6527) );
  NAND4_X1 U7735 ( .A1(n6530), .A2(n6529), .A3(n6528), .A4(n6527), .ZN(n8409)
         );
  XNOR2_X1 U7736 ( .A(n9262), .B(n8409), .ZN(n6922) );
  NAND2_X1 U7737 ( .A1(n6531), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6533) );
  INV_X1 U7738 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n6532) );
  XNOR2_X1 U7739 ( .A(n6533), .B(n6532), .ZN(n8708) );
  INV_X1 U7740 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n7687) );
  OAI22_X1 U7741 ( .A1(n8708), .A2(n6348), .B1(n6534), .B2(n7687), .ZN(n6535)
         );
  INV_X1 U7742 ( .A(n6535), .ZN(n6536) );
  INV_X1 U7743 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n8415) );
  NAND2_X1 U7744 ( .A1(n6796), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n6538) );
  OAI21_X1 U7745 ( .B1(n8415), .B2(n6395), .A(n6538), .ZN(n6543) );
  INV_X1 U7746 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n9112) );
  NAND2_X1 U7747 ( .A1(n6539), .A2(n9112), .ZN(n6540) );
  NAND2_X1 U7748 ( .A1(n6552), .A2(n6540), .ZN(n8414) );
  NOR2_X1 U7749 ( .A1(n8414), .A2(n6384), .ZN(n6542) );
  INV_X1 U7750 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n8317) );
  NOR2_X1 U7751 ( .A1(n6744), .A2(n8317), .ZN(n6541) );
  NAND2_X1 U7752 ( .A1(n7099), .A2(n8308), .ZN(n6929) );
  INV_X1 U7753 ( .A(n8308), .ZN(n8427) );
  NAND2_X1 U7754 ( .A1(n8420), .A2(n8419), .ZN(n8418) );
  NAND2_X1 U7755 ( .A1(n7099), .A2(n8427), .ZN(n6544) );
  AND2_X2 U7756 ( .A1(n8418), .A2(n6544), .ZN(n8951) );
  NAND2_X1 U7757 ( .A1(n7801), .A2(n6833), .ZN(n6550) );
  NAND2_X1 U7758 ( .A1(n6545), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6546) );
  MUX2_X1 U7759 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6546), .S(
        P2_IR_REG_16__SCAN_IN), .Z(n6548) );
  AND2_X1 U7760 ( .A1(n6548), .A2(n6558), .ZN(n8723) );
  AOI22_X1 U7761 ( .A1(n6834), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n7304), .B2(
        n8723), .ZN(n6549) );
  NAND2_X1 U7762 ( .A1(n6550), .A2(n6549), .ZN(n7105) );
  NAND2_X1 U7763 ( .A1(n6552), .A2(n6551), .ZN(n6553) );
  AND2_X1 U7764 ( .A1(n6563), .A2(n6553), .ZN(n8944) );
  NAND2_X1 U7765 ( .A1(n8944), .A2(n6747), .ZN(n6556) );
  AOI22_X1 U7766 ( .A1(n6821), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n6796), .B2(
        P2_REG0_REG_16__SCAN_IN), .ZN(n6555) );
  NAND2_X1 U7767 ( .A1(n6795), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n6554) );
  AND3_X1 U7768 ( .A1(n6556), .A2(n6555), .A3(n6554), .ZN(n7104) );
  NAND2_X1 U7769 ( .A1(n7105), .A2(n7104), .ZN(n6932) );
  NAND2_X1 U7770 ( .A1(n6933), .A2(n6932), .ZN(n8950) );
  INV_X1 U7771 ( .A(n7104), .ZN(n8690) );
  NAND2_X1 U7772 ( .A1(n7105), .A2(n8690), .ZN(n6557) );
  NAND2_X1 U7773 ( .A1(n7916), .A2(n6833), .ZN(n6561) );
  NAND2_X1 U7774 ( .A1(n6558), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6559) );
  XNOR2_X1 U7775 ( .A(n6559), .B(P2_IR_REG_17__SCAN_IN), .ZN(n8738) );
  AOI22_X1 U7776 ( .A1(n6834), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n7304), .B2(
        n8738), .ZN(n6560) );
  AND2_X2 U7777 ( .A1(n6561), .A2(n6560), .ZN(n8453) );
  INV_X1 U7778 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n6567) );
  INV_X1 U7779 ( .A(n6562), .ZN(n6573) );
  NAND2_X1 U7780 ( .A1(n6563), .A2(n8444), .ZN(n6564) );
  NAND2_X1 U7781 ( .A1(n6573), .A2(n6564), .ZN(n8454) );
  OR2_X1 U7782 ( .A1(n8454), .A2(n6384), .ZN(n6566) );
  AOI22_X1 U7783 ( .A1(n6821), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n6796), .B2(
        P2_REG0_REG_17__SCAN_IN), .ZN(n6565) );
  OAI211_X1 U7784 ( .C1(n6744), .C2(n6567), .A(n6566), .B(n6565), .ZN(n8914)
         );
  NAND2_X1 U7785 ( .A1(n8453), .A2(n8914), .ZN(n6940) );
  INV_X1 U7786 ( .A(n8914), .ZN(n8428) );
  NAND2_X1 U7787 ( .A1(n9249), .A2(n8428), .ZN(n6939) );
  NAND2_X1 U7788 ( .A1(n8012), .A2(n6833), .ZN(n6570) );
  INV_X1 U7789 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n6568) );
  XNOR2_X1 U7790 ( .A(n6582), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8736) );
  AOI22_X1 U7791 ( .A1(n6834), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n7304), .B2(
        n8736), .ZN(n6569) );
  INV_X1 U7792 ( .A(n6571), .ZN(n6585) );
  INV_X1 U7793 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n6572) );
  NAND2_X1 U7794 ( .A1(n6573), .A2(n6572), .ZN(n6574) );
  AND2_X1 U7795 ( .A1(n6585), .A2(n6574), .ZN(n8927) );
  NAND2_X1 U7796 ( .A1(n8927), .A2(n6747), .ZN(n6579) );
  INV_X1 U7797 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8752) );
  NAND2_X1 U7798 ( .A1(n6796), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n6576) );
  NAND2_X1 U7799 ( .A1(n6821), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n6575) );
  OAI211_X1 U7800 ( .C1(n8752), .C2(n6744), .A(n6576), .B(n6575), .ZN(n6577)
         );
  INV_X1 U7801 ( .A(n6577), .ZN(n6578) );
  NAND2_X1 U7802 ( .A1(n6579), .A2(n6578), .ZN(n8689) );
  INV_X1 U7803 ( .A(n8689), .ZN(n6730) );
  XNOR2_X1 U7804 ( .A(n9242), .B(n6730), .ZN(n8921) );
  OR2_X1 U7805 ( .A1(n9242), .A2(n8689), .ZN(n6580) );
  NAND2_X1 U7806 ( .A1(n8920), .A2(n6580), .ZN(n8904) );
  NAND2_X1 U7807 ( .A1(n8007), .A2(n6833), .ZN(n6584) );
  AOI22_X1 U7808 ( .A1(n6820), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n10461), 
        .B2(n7304), .ZN(n6583) );
  INV_X1 U7809 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n9118) );
  NAND2_X1 U7810 ( .A1(n6585), .A2(n9118), .ZN(n6586) );
  NAND2_X1 U7811 ( .A1(n6597), .A2(n6586), .ZN(n8906) );
  OR2_X1 U7812 ( .A1(n8906), .A2(n6384), .ZN(n6591) );
  INV_X1 U7813 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n9238) );
  NAND2_X1 U7814 ( .A1(n6796), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n6588) );
  NAND2_X1 U7815 ( .A1(n6821), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n6587) );
  OAI211_X1 U7816 ( .C1(n9238), .C2(n6744), .A(n6588), .B(n6587), .ZN(n6589)
         );
  INV_X1 U7817 ( .A(n6589), .ZN(n6590) );
  INV_X1 U7818 ( .A(n8492), .ZN(n8917) );
  NAND2_X1 U7819 ( .A1(n9232), .A2(n8917), .ZN(n6593) );
  INV_X1 U7820 ( .A(n9232), .ZN(n6592) );
  AOI22_X1 U7821 ( .A1(n8904), .A2(n6593), .B1(n8492), .B2(n6592), .ZN(n8897)
         );
  NAND2_X1 U7822 ( .A1(n8216), .A2(n6833), .ZN(n6595) );
  NAND2_X1 U7823 ( .A1(n6820), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n6594) );
  NAND2_X1 U7824 ( .A1(n6597), .A2(n6596), .ZN(n6598) );
  AND2_X1 U7825 ( .A1(n6599), .A2(n6598), .ZN(n8892) );
  INV_X1 U7826 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n6602) );
  NAND2_X1 U7827 ( .A1(n6796), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n6601) );
  NAND2_X1 U7828 ( .A1(n6821), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n6600) );
  OAI211_X1 U7829 ( .C1(n6602), .C2(n6744), .A(n6601), .B(n6600), .ZN(n6603)
         );
  AOI21_X1 U7830 ( .B1(n8892), .B2(n6747), .A(n6603), .ZN(n8687) );
  OR2_X1 U7831 ( .A1(n9011), .A2(n8687), .ZN(n6953) );
  NAND2_X1 U7832 ( .A1(n9011), .A2(n8687), .ZN(n6955) );
  INV_X1 U7833 ( .A(n9011), .ZN(n8651) );
  NAND2_X1 U7834 ( .A1(n8879), .A2(n8887), .ZN(n6960) );
  NAND2_X1 U7835 ( .A1(n9004), .A2(n8659), .ZN(n6956) );
  NAND2_X1 U7836 ( .A1(n8349), .A2(n6833), .ZN(n6605) );
  NAND2_X1 U7837 ( .A1(n6820), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n6604) );
  INV_X1 U7838 ( .A(n6606), .ZN(n6617) );
  INV_X1 U7839 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n9209) );
  NAND2_X1 U7840 ( .A1(n6607), .A2(n9209), .ZN(n6608) );
  NAND2_X1 U7841 ( .A1(n8859), .A2(n6747), .ZN(n6614) );
  INV_X1 U7842 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n6611) );
  NAND2_X1 U7843 ( .A1(n6821), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n6610) );
  NAND2_X1 U7844 ( .A1(n6796), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n6609) );
  OAI211_X1 U7845 ( .C1(n6744), .C2(n6611), .A(n6610), .B(n6609), .ZN(n6612)
         );
  INV_X1 U7846 ( .A(n6612), .ZN(n6613) );
  NAND2_X1 U7847 ( .A1(n8999), .A2(n8617), .ZN(n6964) );
  INV_X1 U7848 ( .A(n8617), .ZN(n8871) );
  NAND2_X1 U7849 ( .A1(n8396), .A2(n6833), .ZN(n6616) );
  NAND2_X1 U7850 ( .A1(n6820), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n6615) );
  NAND2_X2 U7851 ( .A1(n6616), .A2(n6615), .ZN(n8993) );
  INV_X1 U7852 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n9184) );
  NAND2_X1 U7853 ( .A1(n6617), .A2(n9184), .ZN(n6618) );
  NAND2_X1 U7854 ( .A1(n6619), .A2(n6618), .ZN(n8850) );
  OR2_X1 U7855 ( .A1(n8850), .A2(n6384), .ZN(n6625) );
  INV_X1 U7856 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n6622) );
  NAND2_X1 U7857 ( .A1(n6821), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n6621) );
  NAND2_X1 U7858 ( .A1(n6796), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n6620) );
  OAI211_X1 U7859 ( .C1(n6622), .C2(n6744), .A(n6621), .B(n6620), .ZN(n6623)
         );
  INV_X1 U7860 ( .A(n6623), .ZN(n6624) );
  NAND2_X1 U7861 ( .A1(n8993), .A2(n8661), .ZN(n8826) );
  NOR2_X1 U7862 ( .A1(n8846), .A2(n8845), .ZN(n8998) );
  INV_X1 U7863 ( .A(n8661), .ZN(n8864) );
  NAND2_X1 U7864 ( .A1(n8840), .A2(n8843), .ZN(n6974) );
  INV_X1 U7865 ( .A(n8843), .ZN(n8629) );
  NAND2_X1 U7866 ( .A1(n8987), .A2(n8629), .ZN(n6966) );
  NAND2_X1 U7867 ( .A1(n6974), .A2(n6966), .ZN(n8832) );
  NAND2_X1 U7868 ( .A1(n8434), .A2(n6833), .ZN(n6628) );
  NAND2_X1 U7869 ( .A1(n6820), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n6627) );
  INV_X1 U7870 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n9197) );
  NAND2_X1 U7871 ( .A1(n6629), .A2(n9197), .ZN(n6630) );
  INV_X1 U7872 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n6633) );
  NAND2_X1 U7873 ( .A1(n6796), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n6632) );
  NAND2_X1 U7874 ( .A1(n6821), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n6631) );
  OAI211_X1 U7875 ( .C1(n6633), .C2(n6744), .A(n6632), .B(n6631), .ZN(n6634)
         );
  OR2_X1 U7876 ( .A1(n8982), .A2(n8686), .ZN(n6980) );
  NAND2_X1 U7877 ( .A1(n8982), .A2(n8686), .ZN(n6979) );
  NAND2_X1 U7878 ( .A1(n6980), .A2(n6979), .ZN(n8819) );
  INV_X1 U7879 ( .A(n8982), .ZN(n8818) );
  NAND2_X1 U7880 ( .A1(n8465), .A2(n6833), .ZN(n6636) );
  NAND2_X1 U7881 ( .A1(n6820), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n6635) );
  NAND2_X1 U7882 ( .A1(n6637), .A2(n9114), .ZN(n6638) );
  NAND2_X1 U7883 ( .A1(n6655), .A2(n6638), .ZN(n8798) );
  OR2_X1 U7884 ( .A1(n8798), .A2(n6384), .ZN(n6644) );
  INV_X1 U7885 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n6641) );
  NAND2_X1 U7886 ( .A1(n6796), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n6640) );
  NAND2_X1 U7887 ( .A1(n6821), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n6639) );
  OAI211_X1 U7888 ( .C1(n6641), .C2(n6744), .A(n6640), .B(n6639), .ZN(n6642)
         );
  INV_X1 U7889 ( .A(n6642), .ZN(n6643) );
  NAND2_X1 U7890 ( .A1(n8801), .A2(n8627), .ZN(n8778) );
  NAND2_X1 U7891 ( .A1(n8499), .A2(n6833), .ZN(n6646) );
  NAND2_X1 U7892 ( .A1(n6834), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n6645) );
  XNOR2_X1 U7893 ( .A(n6655), .B(P2_REG3_REG_27__SCAN_IN), .ZN(n8787) );
  NAND2_X1 U7894 ( .A1(n8787), .A2(n6747), .ZN(n6652) );
  INV_X1 U7895 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n6649) );
  NAND2_X1 U7896 ( .A1(n6821), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n6648) );
  NAND2_X1 U7897 ( .A1(n6796), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n6647) );
  OAI211_X1 U7898 ( .C1(n6649), .C2(n6744), .A(n6648), .B(n6647), .ZN(n6650)
         );
  INV_X1 U7899 ( .A(n6650), .ZN(n6651) );
  XNOR2_X1 U7900 ( .A(n8970), .B(n8674), .ZN(n8783) );
  INV_X1 U7901 ( .A(n8970), .ZN(n8790) );
  NAND2_X1 U7902 ( .A1(n10115), .A2(n6833), .ZN(n6654) );
  NAND2_X1 U7903 ( .A1(n6820), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n6653) );
  INV_X1 U7904 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n8608) );
  INV_X1 U7905 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n8548) );
  OAI21_X1 U7906 ( .B1(n6655), .B2(n8608), .A(n8548), .ZN(n6659) );
  AND2_X1 U7907 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(P2_REG3_REG_28__SCAN_IN), 
        .ZN(n6656) );
  INV_X1 U7908 ( .A(n6805), .ZN(n6658) );
  NAND2_X1 U7909 ( .A1(n6659), .A2(n6658), .ZN(n8550) );
  OR2_X1 U7910 ( .A1(n8550), .A2(n6384), .ZN(n6665) );
  INV_X1 U7911 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n6662) );
  NAND2_X1 U7912 ( .A1(n6821), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n6661) );
  NAND2_X1 U7913 ( .A1(n6796), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n6660) );
  OAI211_X1 U7914 ( .C1(n6744), .C2(n6662), .A(n6661), .B(n6660), .ZN(n6663)
         );
  INV_X1 U7915 ( .A(n6663), .ZN(n6664) );
  NAND2_X1 U7916 ( .A1(n8965), .A2(n8609), .ZN(n7007) );
  NAND2_X1 U7917 ( .A1(n7011), .A2(n7007), .ZN(n6992) );
  XNOR2_X1 U7918 ( .A(n6789), .B(n6992), .ZN(n8969) );
  NOR2_X1 U7919 ( .A1(n6666), .A2(P2_IR_REG_20__SCAN_IN), .ZN(n6667) );
  NAND2_X1 U7920 ( .A1(n6668), .A2(n6667), .ZN(n6704) );
  NAND3_X1 U7921 ( .A1(n6706), .A2(n6678), .A3(n6670), .ZN(n6671) );
  NAND2_X1 U7922 ( .A1(n6681), .A2(n6672), .ZN(n6683) );
  NAND2_X1 U7923 ( .A1(n6683), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6673) );
  MUX2_X1 U7924 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6673), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n6675) );
  NAND2_X1 U7925 ( .A1(n6707), .A2(n6706), .ZN(n6677) );
  NAND2_X1 U7926 ( .A1(n6708), .A2(n6678), .ZN(n6679) );
  INV_X1 U7927 ( .A(n10327), .ZN(n8407) );
  INV_X1 U7928 ( .A(P2_B_REG_SCAN_IN), .ZN(n6686) );
  NOR2_X1 U7929 ( .A1(n6681), .A2(n9294), .ZN(n6682) );
  MUX2_X1 U7930 ( .A(n9294), .B(n6682), .S(P2_IR_REG_25__SCAN_IN), .Z(n6685)
         );
  INV_X1 U7931 ( .A(n6683), .ZN(n6684) );
  OAI221_X1 U7932 ( .B1(n10327), .B2(P2_B_REG_SCAN_IN), .C1(n8407), .C2(n6686), 
        .A(n8435), .ZN(n6687) );
  INV_X1 U7933 ( .A(n10328), .ZN(n8498) );
  NAND2_X1 U7934 ( .A1(n8498), .A2(n8435), .ZN(n10153) );
  INV_X1 U7935 ( .A(n7223), .ZN(n7123) );
  OAI22_X1 U7936 ( .A1(n10154), .A2(P2_D_REG_0__SCAN_IN), .B1(n10327), .B2(
        n10328), .ZN(n7121) );
  NOR4_X1 U7937 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n6691) );
  NOR4_X1 U7938 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_18__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n6690) );
  NOR4_X1 U7939 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n6689) );
  NOR4_X1 U7940 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n6688) );
  NAND4_X1 U7941 ( .A1(n6691), .A2(n6690), .A3(n6689), .A4(n6688), .ZN(n6698)
         );
  NOR2_X1 U7942 ( .A1(P2_D_REG_31__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .ZN(
        n6695) );
  NOR4_X1 U7943 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_29__SCAN_IN), .A4(P2_D_REG_28__SCAN_IN), .ZN(n6694) );
  NOR4_X1 U7944 ( .A1(P2_D_REG_23__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n6693) );
  NOR4_X1 U7945 ( .A1(P2_D_REG_27__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_25__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n6692) );
  NAND4_X1 U7946 ( .A1(n6695), .A2(n6694), .A3(n6693), .A4(n6692), .ZN(n6697)
         );
  INV_X1 U7947 ( .A(n10154), .ZN(n6696) );
  AND2_X1 U7948 ( .A1(n7121), .A2(n7120), .ZN(n7224) );
  INV_X1 U7949 ( .A(n8435), .ZN(n6699) );
  XNOR2_X2 U7950 ( .A(n6702), .B(P2_IR_REG_20__SCAN_IN), .ZN(n6715) );
  INV_X1 U7951 ( .A(n6715), .ZN(n6710) );
  INV_X1 U7952 ( .A(n7130), .ZN(n7032) );
  INV_X1 U7953 ( .A(n7371), .ZN(n7305) );
  AOI21_X1 U7954 ( .B1(n7032), .B2(n7305), .A(n7040), .ZN(n6709) );
  AND2_X1 U7955 ( .A1(n7039), .A2(n6709), .ZN(n7221) );
  NAND3_X1 U7956 ( .A1(n7123), .A2(n7224), .A3(n7255), .ZN(n6754) );
  NAND2_X2 U7957 ( .A1(n6754), .A2(n10454), .ZN(n8810) );
  INV_X1 U7958 ( .A(n7046), .ZN(n6714) );
  NAND2_X1 U7959 ( .A1(n6714), .A2(n5072), .ZN(n6713) );
  NAND2_X1 U7960 ( .A1(n4925), .A2(n6713), .ZN(n8051) );
  NAND2_X1 U7961 ( .A1(n6714), .A2(n10461), .ZN(n7662) );
  NAND2_X1 U7962 ( .A1(n8051), .A2(n7662), .ZN(n10463) );
  NAND2_X1 U7963 ( .A1(n6715), .A2(n6871), .ZN(n6716) );
  NAND2_X1 U7964 ( .A1(n5072), .A2(n10461), .ZN(n7027) );
  NAND2_X2 U7965 ( .A1(n6716), .A2(n7027), .ZN(n8937) );
  NAND2_X1 U7966 ( .A1(n6719), .A2(n6718), .ZN(n7832) );
  NAND2_X2 U7967 ( .A1(n7832), .A2(n6720), .ZN(n6866) );
  NAND2_X1 U7968 ( .A1(n6866), .A2(n6869), .ZN(n7474) );
  OR2_X1 U7969 ( .A1(n7474), .A2(n6721), .ZN(n7476) );
  INV_X1 U7970 ( .A(n7768), .ZN(n10445) );
  NAND2_X1 U7971 ( .A1(n10445), .A2(n8698), .ZN(n6722) );
  NAND2_X1 U7972 ( .A1(n10456), .A2(n8697), .ZN(n6886) );
  NAND2_X1 U7973 ( .A1(n7355), .A2(n7675), .ZN(n6885) );
  OR2_X1 U7974 ( .A1(n7681), .A2(n7579), .ZN(n6891) );
  NAND2_X1 U7975 ( .A1(n7681), .A2(n7579), .ZN(n6890) );
  INV_X1 U7976 ( .A(n8694), .ZN(n7821) );
  NAND2_X1 U7977 ( .A1(n7849), .A2(n7821), .ZN(n6901) );
  NAND2_X1 U7978 ( .A1(n8045), .A2(n8049), .ZN(n6724) );
  NAND2_X1 U7979 ( .A1(n8127), .A2(n8132), .ZN(n6725) );
  NAND2_X1 U7980 ( .A1(n6725), .A2(n6860), .ZN(n8243) );
  NAND2_X1 U7981 ( .A1(n8243), .A2(n8242), .ZN(n6727) );
  INV_X1 U7982 ( .A(n8691), .ZN(n8342) );
  NAND2_X1 U7983 ( .A1(n9267), .A2(n8342), .ZN(n6726) );
  INV_X1 U7984 ( .A(n8409), .ZN(n8376) );
  OR2_X1 U7985 ( .A1(n9262), .A2(n8376), .ZN(n6728) );
  NAND2_X1 U7986 ( .A1(n8935), .A2(n6933), .ZN(n6729) );
  NAND2_X1 U7987 ( .A1(n6729), .A2(n6932), .ZN(n8458) );
  OR2_X1 U7988 ( .A1(n9242), .A2(n6730), .ZN(n6731) );
  NAND2_X1 U7989 ( .A1(n9232), .A2(n8492), .ZN(n6949) );
  NAND2_X1 U7990 ( .A1(n8869), .A2(n8882), .ZN(n6733) );
  NAND2_X1 U7991 ( .A1(n6733), .A2(n6960), .ZN(n8863) );
  INV_X1 U7992 ( .A(n8845), .ZN(n6838) );
  INV_X1 U7993 ( .A(n8832), .ZN(n8828) );
  NAND2_X1 U7994 ( .A1(n6735), .A2(n6974), .ZN(n8820) );
  INV_X1 U7995 ( .A(n8819), .ZN(n8813) );
  INV_X1 U7996 ( .A(n6980), .ZN(n6736) );
  NAND2_X1 U7997 ( .A1(n8796), .A2(n6986), .ZN(n8779) );
  INV_X1 U7998 ( .A(n8778), .ZN(n6737) );
  NOR2_X1 U7999 ( .A1(n8783), .A2(n6737), .ZN(n6738) );
  NAND2_X1 U8000 ( .A1(n8779), .A2(n6738), .ZN(n6740) );
  OR2_X1 U8001 ( .A1(n8970), .A2(n8674), .ZN(n6739) );
  XNOR2_X1 U8002 ( .A(n7009), .B(n6992), .ZN(n6749) );
  INV_X1 U8003 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n6745) );
  NAND2_X1 U8004 ( .A1(n6796), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n6743) );
  NAND2_X1 U8005 ( .A1(n6821), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n6742) );
  OAI211_X1 U8006 ( .C1(n6745), .C2(n6744), .A(n6743), .B(n6742), .ZN(n6746)
         );
  AOI21_X1 U8007 ( .B1(n6805), .B2(n6747), .A(n6746), .ZN(n8549) );
  INV_X1 U8008 ( .A(n8549), .ZN(n7466) );
  INV_X1 U8009 ( .A(n6741), .ZN(n6748) );
  AOI222_X1 U8010 ( .A1(n8937), .A2(n6749), .B1(n8685), .B2(n8915), .C1(n7466), 
        .C2(n8916), .ZN(n8968) );
  INV_X1 U8011 ( .A(n9242), .ZN(n8931) );
  INV_X1 U8012 ( .A(n8098), .ZN(n8174) );
  NAND2_X1 U8013 ( .A1(n7231), .A2(n7050), .ZN(n7840) );
  OR2_X1 U8014 ( .A1(n7840), .A2(n7054), .ZN(n7842) );
  NAND2_X1 U8015 ( .A1(n5285), .A2(n7794), .ZN(n7809) );
  NOR2_X1 U8016 ( .A1(n8923), .A2(n9232), .ZN(n6751) );
  NAND2_X1 U8017 ( .A1(n8931), .A2(n6751), .ZN(n8889) );
  NOR2_X2 U8018 ( .A1(n8889), .A2(n9011), .ZN(n8873) );
  NAND2_X1 U8019 ( .A1(n8879), .A2(n8873), .ZN(n8874) );
  NOR2_X4 U8020 ( .A1(n8970), .A2(n8804), .ZN(n8786) );
  INV_X1 U8021 ( .A(n8786), .ZN(n6753) );
  INV_X1 U8022 ( .A(n8965), .ZN(n6757) );
  INV_X1 U8023 ( .A(n6804), .ZN(n6752) );
  AOI21_X1 U8024 ( .B1(n8965), .B2(n6753), .A(n6752), .ZN(n8966) );
  AND2_X4 U8025 ( .A1(n7130), .A2(n10378), .ZN(n8542) );
  AND2_X1 U8026 ( .A1(n10378), .A2(n6715), .ZN(n10452) );
  INV_X1 U8027 ( .A(n8550), .ZN(n6755) );
  INV_X1 U8028 ( .A(n10454), .ZN(n8945) );
  AOI22_X1 U8029 ( .A1(n6755), .A2(n8945), .B1(P2_REG2_REG_28__SCAN_IN), .B2(
        n10466), .ZN(n6756) );
  OAI21_X1 U8030 ( .B1(n6757), .B2(n8930), .A(n6756), .ZN(n6758) );
  AOI21_X1 U8031 ( .B1(n8966), .B2(n8926), .A(n6758), .ZN(n6759) );
  NAND2_X1 U8032 ( .A1(n6781), .A2(n6761), .ZN(n6764) );
  OR2_X1 U8033 ( .A1(n9703), .A2(n6762), .ZN(n6763) );
  NAND2_X1 U8034 ( .A1(n6764), .A2(n6763), .ZN(n6766) );
  XNOR2_X1 U8035 ( .A(n6766), .B(n6765), .ZN(n6771) );
  NAND2_X1 U8036 ( .A1(n6781), .A2(n4856), .ZN(n6768) );
  OAI21_X1 U8037 ( .B1(n9703), .B2(n6769), .A(n6768), .ZN(n6770) );
  XNOR2_X1 U8038 ( .A(n6771), .B(n6770), .ZN(n6776) );
  NAND3_X1 U8039 ( .A1(n6772), .A2(n9413), .A3(n6776), .ZN(n6788) );
  INV_X1 U8040 ( .A(n6775), .ZN(n6773) );
  NOR2_X1 U8041 ( .A1(n6776), .A2(n6774), .ZN(n6785) );
  NAND3_X1 U8042 ( .A1(n6776), .A2(n9413), .A3(n6775), .ZN(n6783) );
  INV_X1 U8043 ( .A(n8594), .ZN(n6778) );
  OAI22_X1 U8044 ( .A1(n9392), .A2(n6778), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n6777), .ZN(n6780) );
  OAI22_X1 U8045 ( .A1(n9768), .A2(n9431), .B1(n9430), .B2(n7368), .ZN(n6779)
         );
  AOI211_X1 U8046 ( .C1(n6781), .C2(n9435), .A(n6780), .B(n6779), .ZN(n6782)
         );
  NAND2_X1 U8047 ( .A1(n6788), .A2(n6787), .ZN(P1_U3218) );
  INV_X1 U8048 ( .A(n6992), .ZN(n6850) );
  OAI22_X1 U8049 ( .A1(n6789), .A2(n6850), .B1(n8965), .B2(n8781), .ZN(n6792)
         );
  NAND2_X1 U8050 ( .A1(n8518), .A2(n6833), .ZN(n6791) );
  NAND2_X1 U8051 ( .A1(n6820), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n6790) );
  OR2_X1 U8052 ( .A1(n8960), .A2(n8549), .ZN(n7014) );
  NAND2_X1 U8053 ( .A1(n8960), .A2(n8549), .ZN(n7010) );
  XNOR2_X1 U8054 ( .A(n6792), .B(n6994), .ZN(n8964) );
  NAND2_X1 U8055 ( .A1(n7009), .A2(n7007), .ZN(n6793) );
  NAND2_X1 U8056 ( .A1(n6793), .A2(n7011), .ZN(n6794) );
  XOR2_X1 U8057 ( .A(n6994), .B(n6794), .Z(n6803) );
  NAND2_X1 U8058 ( .A1(n6795), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n6799) );
  NAND2_X1 U8059 ( .A1(n6821), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n6798) );
  NAND2_X1 U8060 ( .A1(n6796), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n6797) );
  INV_X1 U8061 ( .A(n8512), .ZN(n6800) );
  NAND2_X1 U8062 ( .A1(n6800), .A2(P2_B_REG_SCAN_IN), .ZN(n6801) );
  NAND2_X1 U8063 ( .A1(n8916), .A2(n6801), .ZN(n8765) );
  OAI22_X1 U8064 ( .A1(n8609), .A2(n8675), .B1(n7174), .B2(n8765), .ZN(n6802)
         );
  AOI21_X1 U8065 ( .B1(n8960), .B2(n6804), .A(n8772), .ZN(n8961) );
  AOI22_X1 U8066 ( .A1(n6805), .A2(n8945), .B1(P2_REG2_REG_29__SCAN_IN), .B2(
        n10466), .ZN(n6806) );
  OAI21_X1 U8067 ( .B1(n5118), .B2(n8930), .A(n6806), .ZN(n6807) );
  INV_X1 U8068 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n6811) );
  MUX2_X1 U8069 ( .A(n6811), .B(n8603), .S(n7142), .Z(n6813) );
  INV_X1 U8070 ( .A(SI_30_), .ZN(n9023) );
  NAND2_X1 U8071 ( .A1(n6813), .A2(n9023), .ZN(n6828) );
  AND2_X1 U8072 ( .A1(n6825), .A2(n6828), .ZN(n6812) );
  INV_X1 U8073 ( .A(n6813), .ZN(n6814) );
  NAND2_X1 U8074 ( .A1(n6814), .A2(SI_30_), .ZN(n6827) );
  MUX2_X1 U8075 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .S(n7142), .Z(n6817) );
  INV_X1 U8076 ( .A(SI_31_), .ZN(n6816) );
  XNOR2_X1 U8077 ( .A(n6817), .B(n6816), .ZN(n6818) );
  INV_X1 U8078 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n6824) );
  NAND2_X1 U8079 ( .A1(n6821), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n6823) );
  NAND2_X1 U8080 ( .A1(n6796), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n6822) );
  OAI211_X1 U8081 ( .C1(n6744), .C2(n6824), .A(n6823), .B(n6822), .ZN(n8684)
         );
  NOR2_X1 U8082 ( .A1(n8768), .A2(n8684), .ZN(n7021) );
  NAND2_X1 U8083 ( .A1(n6826), .A2(n6825), .ZN(n6830) );
  AND2_X1 U8084 ( .A1(n6828), .A2(n6827), .ZN(n6829) );
  NAND2_X1 U8085 ( .A1(n6830), .A2(n6829), .ZN(n6832) );
  NAND2_X1 U8086 ( .A1(n8602), .A2(n6833), .ZN(n6836) );
  NAND2_X1 U8087 ( .A1(n6834), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n6835) );
  NOR2_X1 U8088 ( .A1(n10549), .A2(n7174), .ZN(n7017) );
  NOR2_X1 U8089 ( .A1(n7021), .A2(n7017), .ZN(n6855) );
  INV_X1 U8090 ( .A(n6855), .ZN(n6853) );
  INV_X1 U8091 ( .A(n8684), .ZN(n8766) );
  NAND2_X1 U8092 ( .A1(n10549), .A2(n7174), .ZN(n6999) );
  INV_X1 U8093 ( .A(n7022), .ZN(n6852) );
  AND2_X1 U8094 ( .A1(n6891), .A2(n6890), .ZN(n6888) );
  INV_X1 U8095 ( .A(n6888), .ZN(n7672) );
  INV_X1 U8096 ( .A(n7689), .ZN(n7690) );
  NAND2_X1 U8097 ( .A1(n8700), .A2(n7050), .ZN(n7287) );
  NAND2_X1 U8098 ( .A1(n7286), .A2(n7287), .ZN(n10379) );
  NOR4_X1 U8099 ( .A1(n7826), .A2(n6839), .A3(n10379), .A4(n6710), .ZN(n6840)
         );
  NAND3_X1 U8100 ( .A1(n6840), .A2(n7767), .A3(n6874), .ZN(n6841) );
  NOR4_X1 U8101 ( .A1(n7785), .A2(n7672), .A3(n7690), .A4(n6841), .ZN(n6842)
         );
  NAND4_X1 U8102 ( .A1(n8091), .A2(n8049), .A3(n6842), .A4(n7805), .ZN(n6843)
         );
  NOR4_X1 U8103 ( .A1(n8419), .A2(n8128), .A3(n7988), .A4(n6843), .ZN(n6844)
         );
  NAND4_X1 U8104 ( .A1(n6936), .A2(n6844), .A3(n6922), .A4(n8242), .ZN(n6845)
         );
  NOR4_X1 U8105 ( .A1(n8903), .A2(n8921), .A3(n6845), .A4(n8950), .ZN(n6846)
         );
  NAND4_X1 U8106 ( .A1(n8862), .A2(n6847), .A3(n8882), .A4(n6846), .ZN(n6848)
         );
  NOR4_X1 U8107 ( .A1(n8819), .A2(n8832), .A3(n6838), .A4(n6848), .ZN(n6849)
         );
  NAND4_X1 U8108 ( .A1(n6994), .A2(n6850), .A3(n8795), .A4(n6849), .ZN(n6851)
         );
  NAND3_X1 U8109 ( .A1(n8350), .A2(n10461), .A3(n6871), .ZN(n6865) );
  MUX2_X1 U8110 ( .A(n7022), .B(n6855), .S(n7001), .Z(n7004) );
  NAND2_X1 U8111 ( .A1(n6858), .A2(n6912), .ZN(n6856) );
  NAND2_X1 U8112 ( .A1(n6856), .A2(n6860), .ZN(n6862) );
  NAND2_X1 U8113 ( .A1(n6858), .A2(n6857), .ZN(n6859) );
  AND2_X1 U8114 ( .A1(n6860), .A2(n6859), .ZN(n6861) );
  MUX2_X1 U8115 ( .A(n6862), .B(n6861), .S(n7001), .Z(n6917) );
  NAND2_X1 U8116 ( .A1(n6909), .A2(n6902), .ZN(n6863) );
  MUX2_X1 U8117 ( .A(n6864), .B(n6863), .S(n7001), .Z(n6908) );
  INV_X1 U8118 ( .A(n6865), .ZN(n6997) );
  AND2_X1 U8119 ( .A1(n6718), .A2(n7287), .ZN(n6867) );
  OAI21_X1 U8120 ( .B1(n6866), .B2(n6867), .A(n6997), .ZN(n6868) );
  INV_X1 U8121 ( .A(n6869), .ZN(n6870) );
  NOR2_X1 U8122 ( .A1(n6866), .A2(n6870), .ZN(n7835) );
  NAND3_X1 U8123 ( .A1(n6718), .A2(n7287), .A3(n6871), .ZN(n6872) );
  NAND3_X1 U8124 ( .A1(n7835), .A2(n7001), .A3(n6872), .ZN(n6873) );
  NAND3_X1 U8125 ( .A1(n6875), .A2(n6874), .A3(n6873), .ZN(n6880) );
  MUX2_X1 U8126 ( .A(n6877), .B(n6876), .S(n7001), .Z(n6879) );
  MUX2_X1 U8127 ( .A(n7768), .B(n8698), .S(n7001), .Z(n6882) );
  AOI22_X1 U8128 ( .A1(n6880), .A2(n6879), .B1(n6878), .B2(n6882), .ZN(n6884)
         );
  NOR2_X1 U8129 ( .A1(n6882), .A2(n6881), .ZN(n6883) );
  OAI21_X1 U8130 ( .B1(n6884), .B2(n6883), .A(n7689), .ZN(n6889) );
  MUX2_X1 U8131 ( .A(n6886), .B(n6885), .S(n7001), .Z(n6887) );
  NAND3_X1 U8132 ( .A1(n6889), .A2(n6888), .A3(n6887), .ZN(n6895) );
  INV_X1 U8133 ( .A(n6890), .ZN(n6892) );
  MUX2_X1 U8134 ( .A(n6892), .B(n5205), .S(n7001), .Z(n6893) );
  NOR2_X1 U8135 ( .A1(n7785), .A2(n6893), .ZN(n6894) );
  NAND2_X1 U8136 ( .A1(n6895), .A2(n6894), .ZN(n6899) );
  MUX2_X1 U8137 ( .A(n6897), .B(n6896), .S(n7001), .Z(n6898) );
  NOR2_X1 U8138 ( .A1(n7849), .A2(n7821), .ZN(n6904) );
  NAND2_X1 U8139 ( .A1(n6902), .A2(n6901), .ZN(n6903) );
  MUX2_X1 U8140 ( .A(n6904), .B(n6903), .S(n6997), .Z(n6905) );
  OAI21_X1 U8141 ( .B1(n6906), .B2(n6905), .A(n6911), .ZN(n6907) );
  NAND2_X1 U8142 ( .A1(n6910), .A2(n6909), .ZN(n6914) );
  NAND2_X1 U8143 ( .A1(n6912), .A2(n6911), .ZN(n6913) );
  MUX2_X1 U8144 ( .A(n6914), .B(n6913), .S(n7001), .Z(n6915) );
  NAND3_X1 U8145 ( .A1(n6917), .A2(n8242), .A3(n6916), .ZN(n6921) );
  NAND2_X1 U8146 ( .A1(n9267), .A2(n6997), .ZN(n6919) );
  OR2_X1 U8147 ( .A1(n9267), .A2(n6997), .ZN(n6918) );
  MUX2_X1 U8148 ( .A(n6919), .B(n6918), .S(n8691), .Z(n6920) );
  NAND3_X1 U8149 ( .A1(n6922), .A2(n6921), .A3(n6920), .ZN(n6926) );
  NAND2_X1 U8150 ( .A1(n8409), .A2(n6997), .ZN(n6924) );
  NAND2_X1 U8151 ( .A1(n8376), .A2(n7001), .ZN(n6923) );
  MUX2_X1 U8152 ( .A(n6924), .B(n6923), .S(n9262), .Z(n6925) );
  NAND3_X1 U8153 ( .A1(n6927), .A2(n6926), .A3(n6925), .ZN(n6931) );
  MUX2_X1 U8154 ( .A(n6929), .B(n6928), .S(n6997), .Z(n6930) );
  AOI21_X1 U8155 ( .B1(n6931), .B2(n6930), .A(n8950), .ZN(n6938) );
  INV_X1 U8156 ( .A(n6932), .ZN(n6935) );
  INV_X1 U8157 ( .A(n6933), .ZN(n6934) );
  MUX2_X1 U8158 ( .A(n6935), .B(n6934), .S(n7001), .Z(n6937) );
  OAI21_X1 U8159 ( .B1(n6938), .B2(n6937), .A(n6936), .ZN(n6942) );
  MUX2_X1 U8160 ( .A(n6940), .B(n6939), .S(n6997), .Z(n6941) );
  NAND2_X1 U8161 ( .A1(n6942), .A2(n6941), .ZN(n6946) );
  MUX2_X1 U8162 ( .A(n9242), .B(n8689), .S(n7001), .Z(n6945) );
  NOR2_X1 U8163 ( .A1(n6946), .A2(n6945), .ZN(n6943) );
  NAND2_X1 U8164 ( .A1(n6944), .A2(n6943), .ZN(n6954) );
  NAND2_X1 U8165 ( .A1(n6946), .A2(n6945), .ZN(n6950) );
  NAND3_X1 U8166 ( .A1(n6950), .A2(n9242), .A3(n6952), .ZN(n6947) );
  NAND4_X1 U8167 ( .A1(n6954), .A2(n6955), .A3(n6949), .A4(n6947), .ZN(n6948)
         );
  NAND3_X1 U8168 ( .A1(n6950), .A2(n8689), .A3(n6949), .ZN(n6951) );
  NAND4_X1 U8169 ( .A1(n6954), .A2(n6953), .A3(n6952), .A4(n6951), .ZN(n6957)
         );
  AND3_X1 U8170 ( .A1(n6957), .A2(n6956), .A3(n6955), .ZN(n6958) );
  MUX2_X1 U8171 ( .A(n6959), .B(n6958), .S(n6997), .Z(n6963) );
  AOI21_X1 U8172 ( .B1(n6962), .B2(n6960), .A(n7001), .ZN(n6961) );
  AOI21_X1 U8173 ( .B1(n6963), .B2(n6962), .A(n6961), .ZN(n6972) );
  AOI22_X1 U8174 ( .A1(n8845), .A2(n6964), .B1(n6965), .B2(n7001), .ZN(n6971)
         );
  NAND2_X1 U8175 ( .A1(n6974), .A2(n6965), .ZN(n6968) );
  NAND2_X1 U8176 ( .A1(n6966), .A2(n8826), .ZN(n6967) );
  MUX2_X1 U8177 ( .A(n6968), .B(n6967), .S(n7001), .Z(n6969) );
  INV_X1 U8178 ( .A(n6969), .ZN(n6970) );
  OAI21_X1 U8179 ( .B1(n6972), .B2(n6971), .A(n6970), .ZN(n6973) );
  AOI21_X1 U8180 ( .B1(n6973), .B2(n8840), .A(n8819), .ZN(n6978) );
  AND2_X1 U8181 ( .A1(n6979), .A2(n7001), .ZN(n6977) );
  INV_X1 U8182 ( .A(n6973), .ZN(n6976) );
  OAI21_X1 U8183 ( .B1(n8843), .B2(n7001), .A(n6974), .ZN(n6975) );
  OAI22_X1 U8184 ( .A1(n6978), .A2(n6977), .B1(n6976), .B2(n6975), .ZN(n6985)
         );
  NAND2_X1 U8185 ( .A1(n8778), .A2(n6979), .ZN(n6982) );
  NAND2_X1 U8186 ( .A1(n6986), .A2(n6980), .ZN(n6981) );
  MUX2_X1 U8187 ( .A(n6982), .B(n6981), .S(n7001), .Z(n6983) );
  INV_X1 U8188 ( .A(n6983), .ZN(n6984) );
  NAND2_X1 U8189 ( .A1(n6985), .A2(n6984), .ZN(n6988) );
  MUX2_X1 U8190 ( .A(n8778), .B(n6986), .S(n6997), .Z(n6987) );
  AOI21_X1 U8191 ( .B1(n6988), .B2(n6987), .A(n8783), .ZN(n6996) );
  AND2_X1 U8192 ( .A1(n8685), .A2(n6997), .ZN(n6990) );
  NOR2_X1 U8193 ( .A1(n8685), .A2(n6997), .ZN(n6989) );
  MUX2_X1 U8194 ( .A(n6990), .B(n6989), .S(n8970), .Z(n6991) );
  OR2_X1 U8195 ( .A1(n6992), .A2(n6991), .ZN(n6995) );
  MUX2_X1 U8196 ( .A(n7007), .B(n7011), .S(n7001), .Z(n6993) );
  OAI211_X1 U8197 ( .C1(n6996), .C2(n6995), .A(n6994), .B(n6993), .ZN(n7000)
         );
  MUX2_X1 U8198 ( .A(n7010), .B(n7014), .S(n6997), .Z(n6998) );
  MUX2_X1 U8199 ( .A(n8684), .B(n8957), .S(n7001), .Z(n7002) );
  AOI21_X1 U8200 ( .B1(n8768), .B2(n8766), .A(n7002), .ZN(n7003) );
  INV_X1 U8201 ( .A(n7028), .ZN(n7005) );
  AND2_X1 U8202 ( .A1(n7007), .A2(n7010), .ZN(n7008) );
  NAND2_X1 U8203 ( .A1(n7009), .A2(n7008), .ZN(n7016) );
  INV_X1 U8204 ( .A(n7010), .ZN(n7012) );
  OR2_X1 U8205 ( .A1(n7012), .A2(n7011), .ZN(n7013) );
  AND2_X1 U8206 ( .A1(n7014), .A2(n7013), .ZN(n7015) );
  NAND2_X1 U8207 ( .A1(n7016), .A2(n7015), .ZN(n7018) );
  INV_X1 U8208 ( .A(n7018), .ZN(n7020) );
  OAI22_X1 U8209 ( .A1(n7018), .A2(n7017), .B1(n8221), .B2(n8684), .ZN(n7019)
         );
  OAI21_X1 U8210 ( .B1(n7020), .B2(n10549), .A(n7019), .ZN(n7023) );
  XNOR2_X1 U8211 ( .A(n7026), .B(n10461), .ZN(n7024) );
  NAND2_X1 U8212 ( .A1(n7026), .A2(n8542), .ZN(n7030) );
  XNOR2_X1 U8213 ( .A(n7028), .B(n7027), .ZN(n7029) );
  NAND2_X1 U8214 ( .A1(n7040), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8400) );
  INV_X1 U8215 ( .A(n10155), .ZN(n7033) );
  OAI21_X1 U8216 ( .B1(n8400), .B2(n5072), .A(P2_B_REG_SCAN_IN), .ZN(n7034) );
  NAND2_X1 U8217 ( .A1(n5368), .A2(n7035), .ZN(n7036) );
  INV_X1 U8218 ( .A(n7037), .ZN(n7038) );
  INV_X1 U8219 ( .A(n7040), .ZN(n7041) );
  NAND2_X1 U8220 ( .A1(n7209), .A2(n6117), .ZN(n7042) );
  NAND2_X1 U8221 ( .A1(n7042), .A2(n8397), .ZN(n7196) );
  NAND2_X1 U8222 ( .A1(n7196), .A2(n7043), .ZN(n7044) );
  NAND2_X1 U8223 ( .A1(n7044), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U3083) );
  XNOR2_X1 U8224 ( .A(n7068), .B(n7658), .ZN(n7048) );
  NOR2_X1 U8225 ( .A1(n7047), .A2(n7048), .ZN(n7052) );
  NAND2_X1 U8226 ( .A1(n8700), .A2(n7288), .ZN(n7051) );
  MUX2_X1 U8227 ( .A(n7051), .B(n7068), .S(n7050), .Z(n7257) );
  INV_X1 U8228 ( .A(n7052), .ZN(n7053) );
  XNOR2_X1 U8229 ( .A(n7068), .B(n7054), .ZN(n7055) );
  NOR2_X1 U8230 ( .A1(n7056), .A2(n7055), .ZN(n7058) );
  NAND2_X1 U8231 ( .A1(n7298), .A2(n7299), .ZN(n7297) );
  INV_X1 U8232 ( .A(n7058), .ZN(n7059) );
  XNOR2_X1 U8233 ( .A(n8537), .B(n7665), .ZN(n7061) );
  OR2_X1 U8234 ( .A1(n7830), .A2(n8542), .ZN(n7060) );
  XNOR2_X1 U8235 ( .A(n7061), .B(n7060), .ZN(n7308) );
  XNOR2_X1 U8236 ( .A(n7768), .B(n8537), .ZN(n7063) );
  NAND2_X1 U8237 ( .A1(n8698), .A2(n7288), .ZN(n7062) );
  NAND2_X1 U8238 ( .A1(n7063), .A2(n7062), .ZN(n7343) );
  NOR2_X1 U8239 ( .A1(n7063), .A2(n7062), .ZN(n7344) );
  AND2_X1 U8240 ( .A1(n8697), .A2(n7288), .ZN(n7065) );
  XNOR2_X1 U8241 ( .A(n10456), .B(n8537), .ZN(n7064) );
  NOR2_X1 U8242 ( .A1(n7064), .A2(n7065), .ZN(n7066) );
  AOI21_X1 U8243 ( .B1(n7065), .B2(n7064), .A(n7066), .ZN(n7354) );
  INV_X1 U8244 ( .A(n7066), .ZN(n7067) );
  NOR2_X1 U8245 ( .A1(n7579), .A2(n8542), .ZN(n7070) );
  XNOR2_X1 U8246 ( .A(n7681), .B(n8543), .ZN(n7069) );
  NOR2_X1 U8247 ( .A1(n7069), .A2(n7070), .ZN(n7071) );
  AOI21_X1 U8248 ( .B1(n7070), .B2(n7069), .A(n7071), .ZN(n7489) );
  NAND2_X1 U8249 ( .A1(n7488), .A2(n7489), .ZN(n7487) );
  INV_X1 U8250 ( .A(n7071), .ZN(n7072) );
  XNOR2_X1 U8251 ( .A(n7859), .B(n8543), .ZN(n7073) );
  NOR2_X1 U8252 ( .A1(n7719), .A2(n8542), .ZN(n7074) );
  XNOR2_X1 U8253 ( .A(n7073), .B(n7074), .ZN(n7577) );
  XNOR2_X1 U8254 ( .A(n7849), .B(n8543), .ZN(n7076) );
  NAND2_X1 U8255 ( .A1(n8694), .A2(n7288), .ZN(n7075) );
  XNOR2_X1 U8256 ( .A(n7076), .B(n7075), .ZN(n7717) );
  INV_X1 U8257 ( .A(n7075), .ZN(n7077) );
  NOR2_X1 U8258 ( .A1(n7902), .A2(n8542), .ZN(n7079) );
  XNOR2_X1 U8259 ( .A(n8196), .B(n8543), .ZN(n7078) );
  NOR2_X1 U8260 ( .A1(n7078), .A2(n7079), .ZN(n7080) );
  AOI21_X1 U8261 ( .B1(n7079), .B2(n7078), .A(n7080), .ZN(n7817) );
  INV_X1 U8262 ( .A(n7080), .ZN(n7081) );
  NAND2_X1 U8263 ( .A1(n7816), .A2(n7081), .ZN(n7900) );
  XNOR2_X1 U8264 ( .A(n10512), .B(n8543), .ZN(n7082) );
  NOR2_X1 U8265 ( .A1(n7922), .A2(n8542), .ZN(n7083) );
  XNOR2_X1 U8266 ( .A(n7082), .B(n7083), .ZN(n7901) );
  INV_X1 U8267 ( .A(n7082), .ZN(n7085) );
  INV_X1 U8268 ( .A(n7083), .ZN(n7084) );
  NOR2_X1 U8269 ( .A1(n8130), .A2(n8542), .ZN(n7087) );
  XNOR2_X1 U8270 ( .A(n8098), .B(n8543), .ZN(n7086) );
  XOR2_X1 U8271 ( .A(n7087), .B(n7086), .Z(n7920) );
  NOR2_X1 U8272 ( .A1(n8211), .A2(n8542), .ZN(n7089) );
  XNOR2_X1 U8273 ( .A(n8139), .B(n8543), .ZN(n7088) );
  NOR2_X1 U8274 ( .A1(n7088), .A2(n7089), .ZN(n7090) );
  AOI21_X1 U8275 ( .B1(n7089), .B2(n7088), .A(n7090), .ZN(n8120) );
  AND2_X1 U8276 ( .A1(n8691), .A2(n7288), .ZN(n7092) );
  XNOR2_X1 U8277 ( .A(n9267), .B(n8543), .ZN(n7091) );
  NOR2_X1 U8278 ( .A1(n7091), .A2(n7092), .ZN(n7093) );
  AOI21_X1 U8279 ( .B1(n7092), .B2(n7091), .A(n7093), .ZN(n8208) );
  NAND2_X1 U8280 ( .A1(n8207), .A2(n8208), .ZN(n8206) );
  INV_X1 U8281 ( .A(n7093), .ZN(n7094) );
  NAND2_X1 U8282 ( .A1(n8206), .A2(n7094), .ZN(n8303) );
  AND2_X1 U8283 ( .A1(n8409), .A2(n7288), .ZN(n7096) );
  XNOR2_X1 U8284 ( .A(n9262), .B(n8543), .ZN(n7095) );
  NOR2_X1 U8285 ( .A1(n7095), .A2(n7096), .ZN(n7097) );
  AOI21_X1 U8286 ( .B1(n7096), .B2(n7095), .A(n7097), .ZN(n8304) );
  NAND2_X1 U8287 ( .A1(n8303), .A2(n8304), .ZN(n8302) );
  INV_X1 U8288 ( .A(n7097), .ZN(n7098) );
  NAND2_X1 U8289 ( .A1(n8302), .A2(n7098), .ZN(n8372) );
  AND2_X1 U8290 ( .A1(n8308), .A2(n7288), .ZN(n7101) );
  NOR2_X1 U8291 ( .A1(n7100), .A2(n7101), .ZN(n7102) );
  AOI21_X1 U8292 ( .B1(n7101), .B2(n7100), .A(n7102), .ZN(n8373) );
  INV_X1 U8293 ( .A(n7102), .ZN(n7103) );
  NOR2_X1 U8294 ( .A1(n7104), .A2(n8542), .ZN(n7107) );
  XNOR2_X1 U8295 ( .A(n7105), .B(n8543), .ZN(n7106) );
  NOR2_X1 U8296 ( .A1(n7106), .A2(n7107), .ZN(n7108) );
  AOI21_X1 U8297 ( .B1(n7107), .B2(n7106), .A(n7108), .ZN(n8425) );
  XNOR2_X1 U8298 ( .A(n8453), .B(n8537), .ZN(n7110) );
  AND2_X1 U8299 ( .A1(n8914), .A2(n7288), .ZN(n7109) );
  NOR2_X1 U8300 ( .A1(n7110), .A2(n7109), .ZN(n8439) );
  NAND2_X1 U8301 ( .A1(n7110), .A2(n7109), .ZN(n8440) );
  XNOR2_X1 U8302 ( .A(n9242), .B(n8537), .ZN(n7112) );
  NAND2_X1 U8303 ( .A1(n8689), .A2(n7288), .ZN(n7111) );
  NAND2_X1 U8304 ( .A1(n7112), .A2(n7111), .ZN(n8486) );
  XOR2_X1 U8305 ( .A(n8543), .B(n9232), .Z(n7113) );
  NOR2_X1 U8306 ( .A1(n8492), .A2(n8542), .ZN(n8502) );
  INV_X1 U8307 ( .A(n7113), .ZN(n8503) );
  XNOR2_X1 U8308 ( .A(n9011), .B(n8543), .ZN(n7115) );
  NOR2_X1 U8309 ( .A1(n8687), .A2(n8542), .ZN(n7114) );
  NAND2_X1 U8310 ( .A1(n7115), .A2(n7114), .ZN(n7116) );
  OAI21_X1 U8311 ( .B1(n7115), .B2(n7114), .A(n7116), .ZN(n8646) );
  INV_X1 U8312 ( .A(n7116), .ZN(n7117) );
  XNOR2_X1 U8313 ( .A(n8879), .B(n8537), .ZN(n7119) );
  AND2_X1 U8314 ( .A1(n8887), .A2(n7288), .ZN(n7118) );
  NAND2_X1 U8315 ( .A1(n7119), .A2(n7118), .ZN(n8520) );
  OAI21_X1 U8316 ( .B1(n7119), .B2(n7118), .A(n8520), .ZN(n7126) );
  INV_X1 U8317 ( .A(n7120), .ZN(n7122) );
  NAND2_X1 U8318 ( .A1(n7251), .A2(n7123), .ZN(n7128) );
  INV_X1 U8319 ( .A(n7128), .ZN(n7132) );
  INV_X1 U8320 ( .A(n10378), .ZN(n7124) );
  AND3_X1 U8321 ( .A1(n10155), .A2(n7371), .A3(n10536), .ZN(n7125) );
  AOI211_X1 U8322 ( .C1(n7127), .C2(n7126), .A(n8669), .B(n4878), .ZN(n7137)
         );
  NAND2_X1 U8323 ( .A1(n7128), .A2(n7220), .ZN(n7256) );
  AND2_X1 U8324 ( .A1(n10155), .A2(n10550), .ZN(n7129) );
  INV_X1 U8325 ( .A(n8641), .ZN(n8683) );
  NOR2_X1 U8326 ( .A1(n8879), .A2(n8683), .ZN(n7136) );
  AND2_X1 U8327 ( .A1(n10155), .A2(n7130), .ZN(n7131) );
  OAI22_X1 U8328 ( .A1(n8662), .A2(n8617), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9084), .ZN(n7135) );
  NAND2_X1 U8329 ( .A1(n7256), .A2(n7221), .ZN(n7133) );
  OAI22_X1 U8330 ( .A1(n8876), .A2(n8678), .B1(n8660), .B2(n8687), .ZN(n7134)
         );
  OR4_X1 U8331 ( .A1(n7137), .A2(n7136), .A3(n7135), .A4(n7134), .ZN(P2_U3225)
         );
  AOI22_X1 U8332 ( .A1(n9297), .A2(P1_DATAO_REG_1__SCAN_IN), .B1(n10349), .B2(
        P2_STATE_REG_SCAN_IN), .ZN(n7140) );
  OAI21_X1 U8333 ( .B1(n7143), .B2(n8219), .A(n7140), .ZN(P2_U3357) );
  AOI22_X1 U8334 ( .A1(n9297), .A2(P1_DATAO_REG_3__SCAN_IN), .B1(n7441), .B2(
        P2_STATE_REG_SCAN_IN), .ZN(n7141) );
  OAI21_X1 U8335 ( .B1(n7146), .B2(n8219), .A(n7141), .ZN(P2_U3355) );
  INV_X1 U8336 ( .A(n10107), .ZN(n10119) );
  INV_X2 U8337 ( .A(n10114), .ZN(n10113) );
  OAI222_X1 U8338 ( .A1(n10119), .A2(n7144), .B1(n10113), .B2(n7143), .C1(
        n7279), .C2(P1_U3084), .ZN(P1_U3352) );
  AOI22_X1 U8339 ( .A1(n7414), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_4__SCAN_IN), .B2(n9297), .ZN(n7145) );
  OAI21_X1 U8340 ( .B1(n7147), .B2(n8219), .A(n7145), .ZN(P2_U3354) );
  OAI222_X1 U8341 ( .A1(P1_U3084), .A2(n4852), .B1(n10119), .B2(n5502), .C1(
        n7146), .C2(n10113), .ZN(P1_U3350) );
  OAI222_X1 U8342 ( .A1(P1_U3084), .A2(n7647), .B1(n10119), .B2(n5469), .C1(
        n7149), .C2(n10113), .ZN(P1_U3351) );
  OAI222_X1 U8343 ( .A1(n10119), .A2(n7148), .B1(P1_U3084), .B2(n7636), .C1(
        n7147), .C2(n10113), .ZN(P1_U3349) );
  INV_X1 U8344 ( .A(n9297), .ZN(n9300) );
  INV_X1 U8345 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n7150) );
  OAI222_X1 U8346 ( .A1(n9300), .A2(n7150), .B1(n8219), .B2(n7149), .C1(n7389), 
        .C2(P2_U3152), .ZN(P2_U3356) );
  AOI22_X1 U8347 ( .A1(n7427), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_5__SCAN_IN), .B2(n9297), .ZN(n7151) );
  OAI21_X1 U8348 ( .B1(n7153), .B2(n8219), .A(n7151), .ZN(P2_U3353) );
  OAI222_X1 U8349 ( .A1(n10119), .A2(n7154), .B1(n10113), .B2(n7153), .C1(
        n7152), .C2(P1_U3084), .ZN(P1_U3348) );
  AOI22_X1 U8350 ( .A1(n7452), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_6__SCAN_IN), .B2(n9297), .ZN(n7155) );
  OAI21_X1 U8351 ( .B1(n7156), .B2(n8219), .A(n7155), .ZN(P2_U3352) );
  OAI222_X1 U8352 ( .A1(P1_U3084), .A2(n7157), .B1(n10119), .B2(n5610), .C1(
        n7156), .C2(n10113), .ZN(P1_U3347) );
  AOI22_X1 U8353 ( .A1(n7513), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_7__SCAN_IN), .B2(n9297), .ZN(n7158) );
  OAI21_X1 U8354 ( .B1(n7159), .B2(n8219), .A(n7158), .ZN(P2_U3351) );
  INV_X1 U8355 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n7160) );
  INV_X1 U8356 ( .A(n7246), .ZN(n7192) );
  OAI222_X1 U8357 ( .A1(n10119), .A2(n7160), .B1(n10113), .B2(n7159), .C1(
        n7192), .C2(P1_U3084), .ZN(P1_U3346) );
  INV_X1 U8358 ( .A(n7520), .ZN(n7574) );
  INV_X1 U8359 ( .A(n7161), .ZN(n7162) );
  INV_X1 U8360 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n7183) );
  OAI222_X1 U8361 ( .A1(P2_U3152), .A2(n7574), .B1(n8219), .B2(n7162), .C1(
        n9300), .C2(n7183), .ZN(P2_U3350) );
  INV_X1 U8362 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n7163) );
  INV_X1 U8363 ( .A(n7321), .ZN(n7316) );
  OAI222_X1 U8364 ( .A1(n10119), .A2(n7163), .B1(n10113), .B2(n7162), .C1(
        P1_U3084), .C2(n7316), .ZN(P1_U3345) );
  INV_X1 U8365 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n7181) );
  NAND2_X1 U8366 ( .A1(P2_U3966), .A2(n7986), .ZN(n7164) );
  OAI21_X1 U8367 ( .B1(P2_U3966), .B2(n7181), .A(n7164), .ZN(P2_U3563) );
  NAND2_X1 U8368 ( .A1(P2_U3966), .A2(n7789), .ZN(n7165) );
  OAI21_X1 U8369 ( .B1(P2_U3966), .B2(n5610), .A(n7165), .ZN(P2_U3558) );
  INV_X1 U8370 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n7331) );
  NAND2_X1 U8371 ( .A1(P2_U3966), .A2(n8244), .ZN(n7166) );
  OAI21_X1 U8372 ( .B1(P2_U3966), .B2(n7331), .A(n7166), .ZN(P2_U3564) );
  INV_X1 U8373 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n7588) );
  NAND2_X1 U8374 ( .A1(P2_U3966), .A2(n8409), .ZN(n7167) );
  OAI21_X1 U8375 ( .B1(P2_U3966), .B2(n7588), .A(n7167), .ZN(P2_U3566) );
  INV_X1 U8376 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n7685) );
  NAND2_X1 U8377 ( .A1(P2_U3966), .A2(n8308), .ZN(n7168) );
  OAI21_X1 U8378 ( .B1(P2_U3966), .B2(n7685), .A(n7168), .ZN(P2_U3567) );
  INV_X1 U8379 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n7170) );
  INV_X1 U8380 ( .A(n7169), .ZN(n7171) );
  INV_X1 U8381 ( .A(n7502), .ZN(n7319) );
  OAI222_X1 U8382 ( .A1(n10119), .A2(n7170), .B1(n10113), .B2(n7171), .C1(
        n7319), .C2(P1_U3084), .ZN(P1_U3344) );
  INV_X1 U8383 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n7172) );
  OAI222_X1 U8384 ( .A1(n9300), .A2(n7172), .B1(n8219), .B2(n7171), .C1(n7521), 
        .C2(P2_U3152), .ZN(P2_U3349) );
  NAND2_X1 U8385 ( .A1(n8688), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n7173) );
  OAI21_X1 U8386 ( .B1(n8688), .B2(n7174), .A(n7173), .ZN(P2_U3582) );
  INV_X1 U8387 ( .A(n7175), .ZN(n7178) );
  AOI22_X1 U8388 ( .A1(n7556), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n10107), .ZN(n7176) );
  OAI21_X1 U8389 ( .B1(n7178), .B2(n10113), .A(n7176), .ZN(P1_U3343) );
  AOI22_X1 U8390 ( .A1(n7602), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_10__SCAN_IN), .B2(n9297), .ZN(n7177) );
  OAI21_X1 U8391 ( .B1(n7178), .B2(n8219), .A(n7177), .ZN(P2_U3348) );
  INV_X1 U8392 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n7179) );
  INV_X1 U8393 ( .A(n7892), .ZN(n7609) );
  OAI222_X1 U8394 ( .A1(n9300), .A2(n7179), .B1(n8219), .B2(n7180), .C1(n7609), 
        .C2(P2_U3152), .ZN(P2_U3347) );
  INV_X1 U8395 ( .A(n10268), .ZN(n10278) );
  OAI222_X1 U8396 ( .A1(P1_U3084), .A2(n10278), .B1(n10119), .B2(n7181), .C1(
        n7180), .C2(n10113), .ZN(P1_U3342) );
  NAND2_X1 U8397 ( .A1(n8105), .A2(P1_U4006), .ZN(n7182) );
  OAI21_X1 U8398 ( .B1(P1_U4006), .B2(n7183), .A(n7182), .ZN(P1_U3563) );
  NOR2_X1 U8399 ( .A1(n7246), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n7193) );
  NAND2_X1 U8400 ( .A1(n10256), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n7191) );
  INV_X1 U8401 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n7184) );
  MUX2_X1 U8402 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n7184), .S(n10256), .Z(n10262) );
  NAND2_X1 U8403 ( .A1(P1_REG1_REG_5__SCAN_IN), .A2(n10311), .ZN(n7190) );
  NOR2_X1 U8404 ( .A1(n7204), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n7188) );
  INV_X1 U8405 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n7187) );
  NAND2_X1 U8406 ( .A1(P1_REG1_REG_1__SCAN_IN), .A2(n7201), .ZN(n7186) );
  INV_X1 U8407 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n7185) );
  MUX2_X1 U8408 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n7185), .S(n7201), .Z(n7275)
         );
  NAND3_X1 U8409 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .A3(n7275), .ZN(n7274) );
  NAND2_X1 U8410 ( .A1(n7186), .A2(n7274), .ZN(n7643) );
  XNOR2_X1 U8411 ( .A(n7647), .B(P1_REG1_REG_2__SCAN_IN), .ZN(n7644) );
  INV_X1 U8412 ( .A(n7647), .ZN(n7202) );
  AOI22_X1 U8413 ( .A1(n7643), .A2(n7644), .B1(n7202), .B2(
        P1_REG1_REG_2__SCAN_IN), .ZN(n7264) );
  MUX2_X1 U8414 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n7187), .S(n4852), .Z(n7263)
         );
  OR2_X1 U8415 ( .A1(n7264), .A2(n7263), .ZN(n7266) );
  OAI21_X1 U8416 ( .B1(n7187), .B2(n4852), .A(n7266), .ZN(n7627) );
  INV_X1 U8417 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n10442) );
  AOI22_X1 U8418 ( .A1(n7204), .A2(n10442), .B1(P1_REG1_REG_4__SCAN_IN), .B2(
        n7636), .ZN(n7626) );
  NOR2_X1 U8419 ( .A1(n7627), .A2(n7626), .ZN(n7625) );
  NOR2_X1 U8420 ( .A1(n7188), .A2(n7625), .ZN(n10322) );
  INV_X1 U8421 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n7189) );
  MUX2_X1 U8422 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n7189), .S(n10311), .Z(n10321) );
  NAND2_X1 U8423 ( .A1(n10322), .A2(n10321), .ZN(n10319) );
  NAND2_X1 U8424 ( .A1(n7190), .A2(n10319), .ZN(n10263) );
  NAND2_X1 U8425 ( .A1(n10262), .A2(n10263), .ZN(n10261) );
  NAND2_X1 U8426 ( .A1(n7191), .A2(n10261), .ZN(n7241) );
  INV_X1 U8427 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n8167) );
  AOI22_X1 U8428 ( .A1(n7246), .A2(n8167), .B1(P1_REG1_REG_7__SCAN_IN), .B2(
        n7192), .ZN(n7240) );
  NOR2_X1 U8429 ( .A1(n7241), .A2(n7240), .ZN(n7239) );
  NOR2_X1 U8430 ( .A1(n7193), .A2(n7239), .ZN(n7195) );
  INV_X1 U8431 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n10486) );
  AOI22_X1 U8432 ( .A1(P1_REG1_REG_8__SCAN_IN), .A2(n7316), .B1(n7321), .B2(
        n10486), .ZN(n7194) );
  NOR2_X1 U8433 ( .A1(n7195), .A2(n7194), .ZN(n7315) );
  AOI21_X1 U8434 ( .B1(n7195), .B2(n7194), .A(n7315), .ZN(n7219) );
  NAND2_X1 U8435 ( .A1(n7621), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10116) );
  INV_X1 U8436 ( .A(n9695), .ZN(n10245) );
  INV_X1 U8437 ( .A(n7196), .ZN(n10247) );
  NOR2_X1 U8438 ( .A1(n9695), .A2(P1_U3084), .ZN(n8500) );
  NAND2_X1 U8439 ( .A1(n7196), .A2(n8500), .ZN(n10274) );
  INV_X1 U8440 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n7197) );
  AOI22_X1 U8441 ( .A1(P1_REG2_REG_8__SCAN_IN), .A2(n7321), .B1(n7316), .B2(
        n7197), .ZN(n7207) );
  NAND2_X1 U8442 ( .A1(n10256), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n7198) );
  OAI21_X1 U8443 ( .B1(n10256), .B2(P1_REG2_REG_6__SCAN_IN), .A(n7198), .ZN(
        n10259) );
  NOR2_X1 U8444 ( .A1(P1_REG2_REG_5__SCAN_IN), .A2(n10311), .ZN(n7199) );
  AOI21_X1 U8445 ( .B1(n10311), .B2(P1_REG2_REG_5__SCAN_IN), .A(n7199), .ZN(
        n10315) );
  INV_X1 U8446 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n8574) );
  XNOR2_X1 U8447 ( .A(n7647), .B(n8574), .ZN(n7641) );
  NAND2_X1 U8448 ( .A1(P1_REG2_REG_1__SCAN_IN), .A2(n7201), .ZN(n7200) );
  OAI21_X1 U8449 ( .B1(n7201), .B2(P1_REG2_REG_1__SCAN_IN), .A(n7200), .ZN(
        n7281) );
  NAND2_X1 U8450 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n7282) );
  NOR2_X1 U8451 ( .A1(n7281), .A2(n7282), .ZN(n7280) );
  AOI21_X1 U8452 ( .B1(n7201), .B2(P1_REG2_REG_1__SCAN_IN), .A(n7280), .ZN(
        n7642) );
  NOR2_X1 U8453 ( .A1(n7641), .A2(n7642), .ZN(n7640) );
  AOI21_X1 U8454 ( .B1(P1_REG2_REG_2__SCAN_IN), .B2(n7202), .A(n7640), .ZN(
        n7270) );
  XOR2_X1 U8455 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n4852), .Z(n7269) );
  NOR2_X1 U8456 ( .A1(n7270), .A2(n7269), .ZN(n7268) );
  AOI21_X1 U8457 ( .B1(P1_REG2_REG_3__SCAN_IN), .B2(n4849), .A(n7268), .ZN(
        n7630) );
  NOR2_X1 U8458 ( .A1(n7204), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n7203) );
  AOI21_X1 U8459 ( .B1(n7204), .B2(P1_REG2_REG_4__SCAN_IN), .A(n7203), .ZN(
        n7629) );
  NAND2_X1 U8460 ( .A1(n7630), .A2(n7629), .ZN(n7628) );
  OAI21_X1 U8461 ( .B1(n7204), .B2(P1_REG2_REG_4__SCAN_IN), .A(n7628), .ZN(
        n10316) );
  NAND2_X1 U8462 ( .A1(n10315), .A2(n10316), .ZN(n10314) );
  OAI21_X1 U8463 ( .B1(P1_REG2_REG_5__SCAN_IN), .B2(n10311), .A(n10314), .ZN(
        n10258) );
  NOR2_X1 U8464 ( .A1(n10259), .A2(n10258), .ZN(n10257) );
  AOI21_X1 U8465 ( .B1(P1_REG2_REG_6__SCAN_IN), .B2(n10256), .A(n10257), .ZN(
        n7238) );
  NOR2_X1 U8466 ( .A1(n7246), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n7205) );
  AOI21_X1 U8467 ( .B1(P1_REG2_REG_7__SCAN_IN), .B2(n7246), .A(n7205), .ZN(
        n7237) );
  NAND2_X1 U8468 ( .A1(n7238), .A2(n7237), .ZN(n7236) );
  OAI21_X1 U8469 ( .B1(n7246), .B2(P1_REG2_REG_7__SCAN_IN), .A(n7236), .ZN(
        n7206) );
  NAND2_X1 U8470 ( .A1(n7207), .A2(n7206), .ZN(n7320) );
  OAI21_X1 U8471 ( .B1(n7207), .B2(n7206), .A(n7320), .ZN(n7217) );
  INV_X1 U8472 ( .A(n8397), .ZN(n7208) );
  NOR2_X1 U8473 ( .A1(n7209), .A2(n7208), .ZN(n7210) );
  INV_X1 U8474 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n7215) );
  INV_X1 U8475 ( .A(n10274), .ZN(n7211) );
  NAND2_X1 U8476 ( .A1(n10312), .A2(n7321), .ZN(n7214) );
  INV_X1 U8477 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n7212) );
  NOR2_X1 U8478 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7212), .ZN(n8022) );
  INV_X1 U8479 ( .A(n8022), .ZN(n7213) );
  OAI211_X1 U8480 ( .C1(n9736), .C2(n7215), .A(n7214), .B(n7213), .ZN(n7216)
         );
  AOI21_X1 U8481 ( .B1(n10318), .B2(n7217), .A(n7216), .ZN(n7218) );
  OAI21_X1 U8482 ( .B1(n7219), .B2(n10269), .A(n7218), .ZN(P1_U3249) );
  AND2_X1 U8483 ( .A1(n7223), .A2(n7222), .ZN(n7250) );
  INV_X1 U8484 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n7235) );
  NAND2_X1 U8485 ( .A1(n8350), .A2(n10461), .ZN(n7225) );
  OR2_X1 U8486 ( .A1(n6715), .A2(n7225), .ZN(n10510) );
  OR2_X1 U8487 ( .A1(n6839), .A2(n7226), .ZN(n7227) );
  NAND2_X1 U8488 ( .A1(n7228), .A2(n7227), .ZN(n7661) );
  XNOR2_X1 U8489 ( .A(n6839), .B(n7286), .ZN(n7229) );
  OAI22_X1 U8490 ( .A1(n4928), .A2(n8675), .B1(n7472), .B2(n8673), .ZN(n7259)
         );
  AOI21_X1 U8491 ( .B1(n7229), .B2(n8937), .A(n7259), .ZN(n7655) );
  NAND2_X1 U8492 ( .A1(n10377), .A2(n7658), .ZN(n7230) );
  NAND2_X1 U8493 ( .A1(n7840), .A2(n7230), .ZN(n7654) );
  OAI22_X1 U8494 ( .A1(n7654), .A2(n10545), .B1(n7231), .B2(n10536), .ZN(n7232) );
  INV_X1 U8495 ( .A(n7232), .ZN(n7233) );
  OAI211_X1 U8496 ( .C1(n9271), .C2(n7661), .A(n7655), .B(n7233), .ZN(n7252)
         );
  NAND2_X1 U8497 ( .A1(n10557), .A2(n7252), .ZN(n7234) );
  OAI21_X1 U8498 ( .B1(n10557), .B2(n7235), .A(n7234), .ZN(P2_U3454) );
  INV_X1 U8499 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n7249) );
  OAI21_X1 U8500 ( .B1(n7238), .B2(n7237), .A(n7236), .ZN(n7244) );
  AOI21_X1 U8501 ( .B1(n7241), .B2(n7240), .A(n7239), .ZN(n7242) );
  NOR2_X1 U8502 ( .A1(n7242), .A2(n10269), .ZN(n7243) );
  AOI21_X1 U8503 ( .B1(n10318), .B2(n7244), .A(n7243), .ZN(n7248) );
  NAND2_X1 U8504 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3084), .ZN(n7977) );
  INV_X1 U8505 ( .A(n7977), .ZN(n7245) );
  AOI21_X1 U8506 ( .B1(n10312), .B2(n7246), .A(n7245), .ZN(n7247) );
  OAI211_X1 U8507 ( .C1(n7249), .C2(n9736), .A(n7248), .B(n7247), .ZN(P1_U3248) );
  NAND2_X1 U8508 ( .A1(n10553), .A2(n7252), .ZN(n7253) );
  OAI21_X1 U8509 ( .B1(n10553), .B2(n6334), .A(n7253), .ZN(P2_U3521) );
  INV_X1 U8510 ( .A(n9618), .ZN(n9515) );
  NAND2_X1 U8511 ( .A1(n9515), .A2(P1_U4006), .ZN(n7254) );
  OAI21_X1 U8512 ( .B1(n6811), .B2(P1_U4006), .A(n7254), .ZN(P1_U3585) );
  NAND2_X1 U8513 ( .A1(n7256), .A2(n7255), .ZN(n7300) );
  INV_X1 U8514 ( .A(n7300), .ZN(n7295) );
  AOI22_X1 U8515 ( .A1(n8657), .A2(n7260), .B1(n8680), .B2(n7259), .ZN(n7262)
         );
  NAND2_X1 U8516 ( .A1(n8641), .A2(n7658), .ZN(n7261) );
  OAI211_X1 U8517 ( .C1(n7295), .C2(n7653), .A(n7262), .B(n7261), .ZN(P2_U3224) );
  INV_X1 U8518 ( .A(n10312), .ZN(n8269) );
  NAND2_X1 U8519 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_U3084), .ZN(n7591) );
  INV_X1 U8520 ( .A(n10269), .ZN(n10320) );
  NAND2_X1 U8521 ( .A1(n7264), .A2(n7263), .ZN(n7265) );
  NAND3_X1 U8522 ( .A1(n10320), .A2(n7266), .A3(n7265), .ZN(n7267) );
  OAI211_X1 U8523 ( .C1(n8269), .C2(n4852), .A(n7591), .B(n7267), .ZN(n7272)
         );
  AOI211_X1 U8524 ( .C1(n7270), .C2(n7269), .A(n7268), .B(n10298), .ZN(n7271)
         );
  AOI211_X1 U8525 ( .C1(n10313), .C2(P1_ADDR_REG_3__SCAN_IN), .A(n7272), .B(
        n7271), .ZN(n7273) );
  INV_X1 U8526 ( .A(n7273), .ZN(P1_U3244) );
  NAND2_X1 U8527 ( .A1(P1_U3084), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n7278) );
  NOR2_X1 U8528 ( .A1(n10253), .A2(n10250), .ZN(n7276) );
  OAI211_X1 U8529 ( .C1(n7276), .C2(n7275), .A(n10320), .B(n7274), .ZN(n7277)
         );
  OAI211_X1 U8530 ( .C1(n8269), .C2(n7279), .A(n7278), .B(n7277), .ZN(n7284)
         );
  AOI211_X1 U8531 ( .C1(n7282), .C2(n7281), .A(n7280), .B(n10298), .ZN(n7283)
         );
  AOI211_X1 U8532 ( .C1(n10313), .C2(P1_ADDR_REG_1__SCAN_IN), .A(n7284), .B(
        n7283), .ZN(n7285) );
  INV_X1 U8533 ( .A(n7285), .ZN(P1_U3242) );
  INV_X1 U8534 ( .A(n8662), .ZN(n8647) );
  AOI22_X1 U8535 ( .A1(n8647), .A2(n8699), .B1(n8641), .B2(n10377), .ZN(n7293)
         );
  INV_X1 U8536 ( .A(n7286), .ZN(n7291) );
  INV_X1 U8537 ( .A(n7287), .ZN(n7289) );
  MUX2_X1 U8538 ( .A(n10377), .B(n7289), .S(n7288), .Z(n7290) );
  OAI21_X1 U8539 ( .B1(n7291), .B2(n7290), .A(n8657), .ZN(n7292) );
  OAI211_X1 U8540 ( .C1(n7295), .C2(n7294), .A(n7293), .B(n7292), .ZN(P2_U3234) );
  AOI22_X1 U8541 ( .A1(n8647), .A2(n7296), .B1(n8641), .B2(n7054), .ZN(n7303)
         );
  OAI21_X1 U8542 ( .B1(n7299), .B2(n7298), .A(n7297), .ZN(n7301) );
  AOI22_X1 U8543 ( .A1(n8657), .A2(n7301), .B1(n7300), .B2(
        P2_REG3_REG_2__SCAN_IN), .ZN(n7302) );
  OAI211_X1 U8544 ( .C1(n7045), .C2(n8660), .A(n7303), .B(n7302), .ZN(P2_U3239) );
  OAI21_X1 U8545 ( .B1(n10155), .B2(n7031), .A(n7304), .ZN(n7307) );
  NAND2_X1 U8546 ( .A1(n10155), .A2(n7305), .ZN(n7306) );
  NOR2_X1 U8547 ( .A1(n10352), .A2(P2_U3966), .ZN(P2_U3151) );
  XNOR2_X1 U8548 ( .A(n7309), .B(n7308), .ZN(n7314) );
  INV_X1 U8549 ( .A(n8660), .ZN(n8648) );
  INV_X1 U8550 ( .A(n8698), .ZN(n7473) );
  OAI22_X1 U8551 ( .A1(n8683), .A2(n7310), .B1(n8662), .B2(n7473), .ZN(n7311)
         );
  AOI21_X1 U8552 ( .B1(n8648), .B2(n7332), .A(n7311), .ZN(n7313) );
  MUX2_X1 U8553 ( .A(n8678), .B(P2_STATE_REG_SCAN_IN), .S(
        P2_REG3_REG_3__SCAN_IN), .Z(n7312) );
  OAI211_X1 U8554 ( .C1(n7314), .C2(n8669), .A(n7313), .B(n7312), .ZN(P2_U3220) );
  AOI21_X1 U8555 ( .B1(n10486), .B2(n7316), .A(n7315), .ZN(n7318) );
  INV_X1 U8556 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n10496) );
  AOI22_X1 U8557 ( .A1(n7502), .A2(n10496), .B1(P1_REG1_REG_9__SCAN_IN), .B2(
        n7319), .ZN(n7317) );
  NOR2_X1 U8558 ( .A1(n7318), .A2(n7317), .ZN(n7497) );
  AOI21_X1 U8559 ( .B1(n7318), .B2(n7317), .A(n7497), .ZN(n7328) );
  NAND2_X1 U8560 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_U3084), .ZN(n8002) );
  OAI21_X1 U8561 ( .B1(n8269), .B2(n7319), .A(n8002), .ZN(n7326) );
  OAI21_X1 U8562 ( .B1(P1_REG2_REG_8__SCAN_IN), .B2(n7321), .A(n7320), .ZN(
        n7324) );
  NAND2_X1 U8563 ( .A1(n7502), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n7322) );
  OAI21_X1 U8564 ( .B1(n7502), .B2(P1_REG2_REG_9__SCAN_IN), .A(n7322), .ZN(
        n7323) );
  NOR2_X1 U8565 ( .A1(n7323), .A2(n7324), .ZN(n7501) );
  AOI211_X1 U8566 ( .C1(n7324), .C2(n7323), .A(n7501), .B(n10298), .ZN(n7325)
         );
  AOI211_X1 U8567 ( .C1(n10313), .C2(P1_ADDR_REG_9__SCAN_IN), .A(n7326), .B(
        n7325), .ZN(n7327) );
  OAI21_X1 U8568 ( .B1(n7328), .B2(n10269), .A(n7327), .ZN(P1_U3250) );
  AOI22_X1 U8569 ( .A1(n7964), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_12__SCAN_IN), .B2(n9297), .ZN(n7329) );
  OAI21_X1 U8570 ( .B1(n7330), .B2(n8219), .A(n7329), .ZN(P2_U3346) );
  INV_X1 U8571 ( .A(n7709), .ZN(n7552) );
  OAI222_X1 U8572 ( .A1(P1_U3084), .A2(n7552), .B1(n10119), .B2(n7331), .C1(
        n7330), .C2(n10113), .ZN(P1_U3341) );
  NAND2_X1 U8573 ( .A1(P2_U3966), .A2(n7332), .ZN(n7333) );
  OAI21_X1 U8574 ( .B1(P2_U3966), .B2(n5469), .A(n7333), .ZN(P2_U3554) );
  XOR2_X1 U8575 ( .A(n7335), .B(n7334), .Z(n7622) );
  NAND2_X1 U8576 ( .A1(n7622), .A2(n9413), .ZN(n7338) );
  OR2_X1 U8577 ( .A1(n7336), .A2(P1_U3084), .ZN(n8589) );
  AOI22_X1 U8578 ( .A1(n9435), .A2(n10385), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        n8589), .ZN(n7337) );
  OAI211_X1 U8579 ( .C1(n9592), .C2(n9430), .A(n7338), .B(n7337), .ZN(P1_U3230) );
  INV_X1 U8580 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n7340) );
  NAND2_X1 U8581 ( .A1(n8864), .A2(P2_U3966), .ZN(n7339) );
  OAI21_X1 U8582 ( .B1(P2_U3966), .B2(n7340), .A(n7339), .ZN(P2_U3575) );
  INV_X1 U8583 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n8403) );
  NAND2_X1 U8584 ( .A1(n8843), .A2(P2_U3966), .ZN(n7341) );
  OAI21_X1 U8585 ( .B1(n8403), .B2(P2_U3966), .A(n7341), .ZN(P2_U3576) );
  NAND2_X1 U8586 ( .A1(P2_U3966), .A2(n7296), .ZN(n7342) );
  OAI21_X1 U8587 ( .B1(P2_U3966), .B2(n5502), .A(n7342), .ZN(P2_U3555) );
  NOR2_X1 U8588 ( .A1(n7344), .A2(n5060), .ZN(n7345) );
  XNOR2_X1 U8589 ( .A(n7346), .B(n7345), .ZN(n7351) );
  INV_X1 U8590 ( .A(n7760), .ZN(n7349) );
  INV_X1 U8591 ( .A(n8678), .ZN(n8665) );
  OAI22_X1 U8592 ( .A1(n7830), .A2(n8660), .B1(n8662), .B2(n7675), .ZN(n7348)
         );
  INV_X1 U8593 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n9202) );
  OAI22_X1 U8594 ( .A1(n8683), .A2(n10445), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9202), .ZN(n7347) );
  AOI211_X1 U8595 ( .C1(n7349), .C2(n8665), .A(n7348), .B(n7347), .ZN(n7350)
         );
  OAI21_X1 U8596 ( .B1(n7351), .B2(n8669), .A(n7350), .ZN(P2_U3232) );
  OAI21_X1 U8597 ( .B1(n7354), .B2(n7353), .A(n7352), .ZN(n7359) );
  OAI22_X1 U8598 ( .A1(n7473), .A2(n8660), .B1(n8662), .B2(n7579), .ZN(n7358)
         );
  NAND2_X1 U8599 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(P2_U3152), .ZN(n7419) );
  NAND2_X1 U8600 ( .A1(n8641), .A2(n7355), .ZN(n7356) );
  OAI211_X1 U8601 ( .C1(n8678), .C2(n10453), .A(n7419), .B(n7356), .ZN(n7357)
         );
  AOI211_X1 U8602 ( .C1(n7359), .C2(n8657), .A(n7358), .B(n7357), .ZN(n7360)
         );
  INV_X1 U8603 ( .A(n7360), .ZN(P2_U3229) );
  INV_X1 U8604 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n7367) );
  AND2_X1 U8605 ( .A1(n6205), .A2(n7365), .ZN(n9589) );
  NOR2_X1 U8606 ( .A1(n10396), .A2(n9589), .ZN(n9655) );
  NAND2_X1 U8607 ( .A1(n9696), .A2(n7364), .ZN(n7361) );
  OR2_X1 U8608 ( .A1(n9655), .A2(n7361), .ZN(n7363) );
  NAND2_X1 U8609 ( .A1(n9718), .A2(n10391), .ZN(n7362) );
  AND2_X1 U8610 ( .A1(n7363), .A2(n7362), .ZN(n10372) );
  OAI21_X1 U8611 ( .B1(n7365), .B2(n7364), .A(n10372), .ZN(n10083) );
  NAND2_X1 U8612 ( .A1(n10083), .A2(n10535), .ZN(n7366) );
  OAI21_X1 U8613 ( .B1(n10535), .B2(n7367), .A(n7366), .ZN(P1_U3454) );
  INV_X1 U8614 ( .A(n7368), .ZN(n7369) );
  NAND2_X1 U8615 ( .A1(n7369), .A2(P1_U4006), .ZN(n7370) );
  OAI21_X1 U8616 ( .B1(n6177), .B2(P1_U4006), .A(n7370), .ZN(P1_U3584) );
  NAND2_X1 U8617 ( .A1(n10155), .A2(n7371), .ZN(n7374) );
  INV_X1 U8618 ( .A(n7372), .ZN(n7373) );
  NAND3_X1 U8619 ( .A1(n7374), .A2(n8400), .A3(n7373), .ZN(n7377) );
  NAND2_X1 U8620 ( .A1(n7377), .A2(n6348), .ZN(n7375) );
  NAND2_X1 U8621 ( .A1(n7375), .A2(n8688), .ZN(n7395) );
  AND2_X1 U8622 ( .A1(n6348), .A2(n8512), .ZN(n7376) );
  MUX2_X1 U8623 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n6412), .S(n7452), .Z(n7385)
         );
  XNOR2_X1 U8624 ( .A(n7414), .B(P2_REG1_REG_4__SCAN_IN), .ZN(n7402) );
  INV_X1 U8625 ( .A(n7389), .ZN(n10363) );
  NAND2_X1 U8626 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n10343) );
  NAND2_X1 U8627 ( .A1(n10349), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n7378) );
  OAI21_X1 U8628 ( .B1(n10349), .B2(P2_REG1_REG_1__SCAN_IN), .A(n7378), .ZN(
        n10342) );
  NOR2_X1 U8629 ( .A1(n10343), .A2(n10342), .ZN(n10341) );
  MUX2_X1 U8630 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n7379), .S(n7389), .Z(n10355)
         );
  AOI21_X1 U8631 ( .B1(n10363), .B2(P2_REG1_REG_2__SCAN_IN), .A(n10354), .ZN(
        n7430) );
  MUX2_X1 U8632 ( .A(n7380), .B(P2_REG1_REG_3__SCAN_IN), .S(n7441), .Z(n7431)
         );
  NOR2_X1 U8633 ( .A1(n7430), .A2(n7431), .ZN(n7429) );
  NAND2_X1 U8634 ( .A1(n7414), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n7381) );
  NAND2_X1 U8635 ( .A1(n7404), .A2(n7381), .ZN(n7417) );
  NAND2_X1 U8636 ( .A1(n7427), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n7383) );
  OAI21_X1 U8637 ( .B1(n7427), .B2(P2_REG1_REG_5__SCAN_IN), .A(n7383), .ZN(
        n7382) );
  INV_X1 U8638 ( .A(n7382), .ZN(n7418) );
  NAND2_X1 U8639 ( .A1(n7417), .A2(n7418), .ZN(n7416) );
  NAND2_X1 U8640 ( .A1(n7416), .A2(n7383), .ZN(n7384) );
  NAND2_X1 U8641 ( .A1(n7384), .A2(n7385), .ZN(n7445) );
  OAI21_X1 U8642 ( .B1(n7385), .B2(n7384), .A(n7445), .ZN(n7387) );
  INV_X1 U8643 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n10181) );
  OR2_X1 U8644 ( .A1(n8741), .A2(n10181), .ZN(n7386) );
  NAND2_X1 U8645 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3152), .ZN(n7491) );
  OAI211_X1 U8646 ( .C1(n10353), .C2(n7387), .A(n7386), .B(n7491), .ZN(n7399)
         );
  XNOR2_X1 U8647 ( .A(n7414), .B(P2_REG2_REG_4__SCAN_IN), .ZN(n7410) );
  NAND2_X1 U8648 ( .A1(n10349), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n7388) );
  OAI21_X1 U8649 ( .B1(n10349), .B2(P2_REG2_REG_1__SCAN_IN), .A(n7388), .ZN(
        n10345) );
  NAND2_X1 U8650 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n10346) );
  INV_X1 U8651 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n7390) );
  MUX2_X1 U8652 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n7390), .S(n7389), .Z(n10359)
         );
  MUX2_X1 U8653 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n7667), .S(n7441), .Z(n7391)
         );
  INV_X1 U8654 ( .A(n7391), .ZN(n7437) );
  NOR2_X1 U8655 ( .A1(n7438), .A2(n7437), .ZN(n7436) );
  AOI21_X1 U8656 ( .B1(n7441), .B2(P2_REG2_REG_3__SCAN_IN), .A(n7436), .ZN(
        n7411) );
  NOR2_X1 U8657 ( .A1(n7410), .A2(n7411), .ZN(n7409) );
  AOI21_X1 U8658 ( .B1(P2_REG2_REG_4__SCAN_IN), .B2(n7414), .A(n7409), .ZN(
        n7424) );
  NAND2_X1 U8659 ( .A1(n7427), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n7392) );
  OAI21_X1 U8660 ( .B1(n7427), .B2(P2_REG2_REG_5__SCAN_IN), .A(n7392), .ZN(
        n7423) );
  NOR2_X1 U8661 ( .A1(n7424), .A2(n7423), .ZN(n7422) );
  AOI21_X1 U8662 ( .B1(P2_REG2_REG_5__SCAN_IN), .B2(n7427), .A(n7422), .ZN(
        n7397) );
  MUX2_X1 U8663 ( .A(n7393), .B(P2_REG2_REG_6__SCAN_IN), .S(n7452), .Z(n7396)
         );
  NOR2_X1 U8664 ( .A1(n7397), .A2(n7396), .ZN(n7451) );
  NOR2_X1 U8665 ( .A1(n6741), .A2(n8512), .ZN(n7394) );
  AOI211_X1 U8666 ( .C1(n7397), .C2(n7396), .A(n7451), .B(n10357), .ZN(n7398)
         );
  AOI211_X1 U8667 ( .C1(n10364), .C2(n7452), .A(n7399), .B(n7398), .ZN(n7400)
         );
  INV_X1 U8668 ( .A(n7400), .ZN(P2_U3251) );
  NAND2_X1 U8669 ( .A1(n7402), .A2(n7401), .ZN(n7403) );
  NAND2_X1 U8670 ( .A1(n7404), .A2(n7403), .ZN(n7408) );
  INV_X1 U8671 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n7405) );
  OR2_X1 U8672 ( .A1(n8741), .A2(n7405), .ZN(n7407) );
  NAND2_X1 U8673 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3152), .ZN(n7406) );
  OAI211_X1 U8674 ( .C1(n7408), .C2(n10353), .A(n7407), .B(n7406), .ZN(n7413)
         );
  AOI211_X1 U8675 ( .C1(n7411), .C2(n7410), .A(n7409), .B(n10357), .ZN(n7412)
         );
  AOI211_X1 U8676 ( .C1(n10364), .C2(n7414), .A(n7413), .B(n7412), .ZN(n7415)
         );
  INV_X1 U8677 ( .A(n7415), .ZN(P2_U3249) );
  OAI21_X1 U8678 ( .B1(n7418), .B2(n7417), .A(n7416), .ZN(n7421) );
  INV_X1 U8679 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n10176) );
  OR2_X1 U8680 ( .A1(n8741), .A2(n10176), .ZN(n7420) );
  OAI211_X1 U8681 ( .C1(n10353), .C2(n7421), .A(n7420), .B(n7419), .ZN(n7426)
         );
  AOI211_X1 U8682 ( .C1(n7424), .C2(n7423), .A(n7422), .B(n10357), .ZN(n7425)
         );
  AOI211_X1 U8683 ( .C1(n10364), .C2(n7427), .A(n7426), .B(n7425), .ZN(n7428)
         );
  INV_X1 U8684 ( .A(n7428), .ZN(P2_U3250) );
  INV_X1 U8685 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n7435) );
  AOI21_X1 U8686 ( .B1(n7431), .B2(n7430), .A(n7429), .ZN(n7432) );
  NAND2_X1 U8687 ( .A1(n10333), .A2(n7432), .ZN(n7434) );
  NAND2_X1 U8688 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_U3152), .ZN(n7433) );
  OAI211_X1 U8689 ( .C1(n8741), .C2(n7435), .A(n7434), .B(n7433), .ZN(n7440)
         );
  AOI211_X1 U8690 ( .C1(n7438), .C2(n7437), .A(n7436), .B(n10357), .ZN(n7439)
         );
  AOI211_X1 U8691 ( .C1(n10364), .C2(n7441), .A(n7440), .B(n7439), .ZN(n7442)
         );
  INV_X1 U8692 ( .A(n7442), .ZN(P2_U3248) );
  NAND2_X1 U8693 ( .A1(n7513), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n7518) );
  OAI21_X1 U8694 ( .B1(n7513), .B2(P2_REG1_REG_7__SCAN_IN), .A(n7518), .ZN(
        n7443) );
  INV_X1 U8695 ( .A(n7443), .ZN(n7447) );
  NAND2_X1 U8696 ( .A1(n7452), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n7444) );
  NAND2_X1 U8697 ( .A1(n7445), .A2(n7444), .ZN(n7446) );
  NAND2_X1 U8698 ( .A1(n7446), .A2(n7447), .ZN(n7519) );
  OAI21_X1 U8699 ( .B1(n7447), .B2(n7446), .A(n7519), .ZN(n7450) );
  INV_X1 U8700 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n10186) );
  OR2_X1 U8701 ( .A1(n8741), .A2(n10186), .ZN(n7449) );
  NAND2_X1 U8702 ( .A1(P2_REG3_REG_7__SCAN_IN), .A2(P2_U3152), .ZN(n7448) );
  OAI211_X1 U8703 ( .C1(n10353), .C2(n7450), .A(n7449), .B(n7448), .ZN(n7457)
         );
  AOI21_X1 U8704 ( .B1(P2_REG2_REG_6__SCAN_IN), .B2(n7452), .A(n7451), .ZN(
        n7455) );
  NAND2_X1 U8705 ( .A1(n7513), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n7453) );
  OAI21_X1 U8706 ( .B1(n7513), .B2(P2_REG2_REG_7__SCAN_IN), .A(n7453), .ZN(
        n7454) );
  NOR2_X1 U8707 ( .A1(n7455), .A2(n7454), .ZN(n7512) );
  AOI211_X1 U8708 ( .C1(n7455), .C2(n7454), .A(n10357), .B(n7512), .ZN(n7456)
         );
  AOI211_X1 U8709 ( .C1(n10364), .C2(n7513), .A(n7457), .B(n7456), .ZN(n7458)
         );
  INV_X1 U8710 ( .A(n7458), .ZN(P2_U3252) );
  NAND2_X1 U8711 ( .A1(n7459), .A2(n7460), .ZN(n7462) );
  XNOR2_X1 U8712 ( .A(n7462), .B(n7461), .ZN(n7465) );
  AOI22_X1 U8713 ( .A1(n9435), .A2(n10408), .B1(P1_REG3_REG_1__SCAN_IN), .B2(
        n8589), .ZN(n7464) );
  AOI22_X1 U8714 ( .A1(n9417), .A2(n6205), .B1(n9416), .B2(n10392), .ZN(n7463)
         );
  OAI211_X1 U8715 ( .C1(n7465), .C2(n9438), .A(n7464), .B(n7463), .ZN(P1_U3220) );
  NAND2_X1 U8716 ( .A1(n7466), .A2(P2_U3966), .ZN(n7467) );
  OAI21_X1 U8717 ( .B1(n6184), .B2(P2_U3966), .A(n7467), .ZN(P2_U3581) );
  INV_X1 U8718 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n7484) );
  NAND2_X1 U8719 ( .A1(n7468), .A2(n7469), .ZN(n7471) );
  NAND2_X1 U8720 ( .A1(n7471), .A2(n6721), .ZN(n7470) );
  OAI21_X1 U8721 ( .B1(n7471), .B2(n6721), .A(n7470), .ZN(n7479) );
  INV_X1 U8722 ( .A(n7479), .ZN(n7670) );
  INV_X1 U8723 ( .A(n8051), .ZN(n7829) );
  OAI22_X1 U8724 ( .A1(n7473), .A2(n8673), .B1(n7472), .B2(n8675), .ZN(n7478)
         );
  NAND2_X1 U8725 ( .A1(n7474), .A2(n6721), .ZN(n7475) );
  INV_X1 U8726 ( .A(n8937), .ZN(n8461) );
  AOI21_X1 U8727 ( .B1(n7476), .B2(n7475), .A(n8461), .ZN(n7477) );
  AOI211_X1 U8728 ( .C1(n7829), .C2(n7479), .A(n7478), .B(n7477), .ZN(n7666)
         );
  AND2_X1 U8729 ( .A1(n7842), .A2(n7665), .ZN(n7480) );
  OR2_X1 U8730 ( .A1(n7480), .A2(n7757), .ZN(n7663) );
  INV_X1 U8731 ( .A(n7663), .ZN(n7481) );
  AOI22_X1 U8732 ( .A1(n7481), .A2(n10429), .B1(n10550), .B2(n7665), .ZN(n7482) );
  OAI211_X1 U8733 ( .C1(n7670), .C2(n10510), .A(n7666), .B(n7482), .ZN(n7485)
         );
  NAND2_X1 U8734 ( .A1(n7485), .A2(n10557), .ZN(n7483) );
  OAI21_X1 U8735 ( .B1(n10557), .B2(n7484), .A(n7483), .ZN(P2_U3460) );
  NAND2_X1 U8736 ( .A1(n7485), .A2(n10553), .ZN(n7486) );
  OAI21_X1 U8737 ( .B1(n10553), .B2(n7380), .A(n7486), .ZN(P2_U3523) );
  OAI21_X1 U8738 ( .B1(n7489), .B2(n7488), .A(n7487), .ZN(n7494) );
  OAI22_X1 U8739 ( .A1(n7675), .A2(n8660), .B1(n8662), .B2(n7719), .ZN(n7493)
         );
  NAND2_X1 U8740 ( .A1(n8641), .A2(n7681), .ZN(n7490) );
  OAI211_X1 U8741 ( .C1(n8678), .C2(n7678), .A(n7491), .B(n7490), .ZN(n7492)
         );
  AOI211_X1 U8742 ( .C1(n7494), .C2(n8657), .A(n7493), .B(n7492), .ZN(n7495)
         );
  INV_X1 U8743 ( .A(n7495), .ZN(P2_U3241) );
  NOR2_X1 U8744 ( .A1(n7502), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n7496) );
  NOR2_X1 U8745 ( .A1(n7497), .A2(n7496), .ZN(n7500) );
  INV_X1 U8746 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n7498) );
  MUX2_X1 U8747 ( .A(n7498), .B(P1_REG1_REG_10__SCAN_IN), .S(n7556), .Z(n7499)
         );
  NOR2_X1 U8748 ( .A1(n7500), .A2(n7499), .ZN(n7547) );
  AOI21_X1 U8749 ( .B1(n7500), .B2(n7499), .A(n7547), .ZN(n7511) );
  AND2_X1 U8750 ( .A1(P1_U3084), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n8229) );
  INV_X1 U8751 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n7508) );
  AOI21_X1 U8752 ( .B1(n7502), .B2(P1_REG2_REG_9__SCAN_IN), .A(n7501), .ZN(
        n7505) );
  NAND2_X1 U8753 ( .A1(P1_REG2_REG_10__SCAN_IN), .A2(n7556), .ZN(n7503) );
  OAI21_X1 U8754 ( .B1(n7556), .B2(P1_REG2_REG_10__SCAN_IN), .A(n7503), .ZN(
        n7504) );
  NOR2_X1 U8755 ( .A1(n7505), .A2(n7504), .ZN(n7555) );
  AOI211_X1 U8756 ( .C1(n7505), .C2(n7504), .A(n7555), .B(n10298), .ZN(n7506)
         );
  INV_X1 U8757 ( .A(n7506), .ZN(n7507) );
  OAI21_X1 U8758 ( .B1(n7508), .B2(n9736), .A(n7507), .ZN(n7509) );
  AOI211_X1 U8759 ( .C1(n10312), .C2(n7556), .A(n8229), .B(n7509), .ZN(n7510)
         );
  OAI21_X1 U8760 ( .B1(n7511), .B2(n10269), .A(n7510), .ZN(P1_U3251) );
  XNOR2_X1 U8761 ( .A(n7520), .B(P2_REG2_REG_8__SCAN_IN), .ZN(n7564) );
  MUX2_X1 U8762 ( .A(n8058), .B(P2_REG2_REG_9__SCAN_IN), .S(n7521), .Z(n7514)
         );
  INV_X1 U8763 ( .A(n7514), .ZN(n7534) );
  AOI21_X1 U8764 ( .B1(P2_REG2_REG_9__SCAN_IN), .B2(n7538), .A(n7533), .ZN(
        n7517) );
  MUX2_X1 U8765 ( .A(P2_REG2_REG_10__SCAN_IN), .B(n7993), .S(n7602), .Z(n7515)
         );
  INV_X1 U8766 ( .A(n7515), .ZN(n7516) );
  AOI211_X1 U8767 ( .C1(n7517), .C2(n7516), .A(n7597), .B(n10357), .ZN(n7532)
         );
  NAND2_X1 U8768 ( .A1(n7519), .A2(n7518), .ZN(n7570) );
  MUX2_X1 U8769 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n6437), .S(n7520), .Z(n7571)
         );
  AND2_X1 U8770 ( .A1(n7570), .A2(n7571), .ZN(n7568) );
  NOR2_X1 U8771 ( .A1(n7522), .A2(n7521), .ZN(n7523) );
  XNOR2_X1 U8772 ( .A(n7522), .B(n7521), .ZN(n7537) );
  NOR2_X1 U8773 ( .A1(n6452), .A2(n7537), .ZN(n7536) );
  INV_X1 U8774 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n7524) );
  MUX2_X1 U8775 ( .A(n7524), .B(P2_REG1_REG_10__SCAN_IN), .S(n7602), .Z(n7525)
         );
  NOR2_X1 U8776 ( .A1(n7526), .A2(n7525), .ZN(n7601) );
  AOI211_X1 U8777 ( .C1(n7526), .C2(n7525), .A(n7601), .B(n10353), .ZN(n7531)
         );
  INV_X1 U8778 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n7529) );
  NAND2_X1 U8779 ( .A1(n10364), .A2(n7602), .ZN(n7528) );
  NAND2_X1 U8780 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3152), .ZN(n7527) );
  OAI211_X1 U8781 ( .C1(n8741), .C2(n7529), .A(n7528), .B(n7527), .ZN(n7530)
         );
  OR3_X1 U8782 ( .A1(n7532), .A2(n7531), .A3(n7530), .ZN(P2_U3255) );
  AOI211_X1 U8783 ( .C1(n7535), .C2(n7534), .A(n10357), .B(n7533), .ZN(n7542)
         );
  AOI211_X1 U8784 ( .C1(n7537), .C2(n6452), .A(n7536), .B(n10353), .ZN(n7541)
         );
  INV_X1 U8785 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n10196) );
  NAND2_X1 U8786 ( .A1(n10364), .A2(n7538), .ZN(n7539) );
  NAND2_X1 U8787 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3152), .ZN(n7820) );
  OAI211_X1 U8788 ( .C1(n8741), .C2(n10196), .A(n7539), .B(n7820), .ZN(n7540)
         );
  OR3_X1 U8789 ( .A1(n7542), .A2(n7541), .A3(n7540), .ZN(P2_U3254) );
  INV_X1 U8790 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n7544) );
  INV_X1 U8791 ( .A(n7543), .ZN(n7545) );
  INV_X1 U8792 ( .A(n8037), .ZN(n8028) );
  OAI222_X1 U8793 ( .A1(n9300), .A2(n7544), .B1(n8219), .B2(n7545), .C1(
        P2_U3152), .C2(n8028), .ZN(P2_U3345) );
  INV_X1 U8794 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n7546) );
  INV_X1 U8795 ( .A(n10293), .ZN(n7707) );
  OAI222_X1 U8796 ( .A1(n10119), .A2(n7546), .B1(n10113), .B2(n7545), .C1(
        P1_U3084), .C2(n7707), .ZN(P1_U3340) );
  INV_X1 U8797 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n7562) );
  XNOR2_X1 U8798 ( .A(n7552), .B(P1_REG1_REG_12__SCAN_IN), .ZN(n7551) );
  OR2_X1 U8799 ( .A1(n7556), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n7549) );
  INV_X1 U8800 ( .A(n7547), .ZN(n7548) );
  NAND2_X1 U8801 ( .A1(n7549), .A2(n7548), .ZN(n10279) );
  INV_X1 U8802 ( .A(n10279), .ZN(n10277) );
  INV_X1 U8803 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n10530) );
  OAI21_X1 U8804 ( .B1(n10279), .B2(n10530), .A(n10278), .ZN(n7550) );
  OAI21_X1 U8805 ( .B1(n10277), .B2(P1_REG1_REG_11__SCAN_IN), .A(n7550), .ZN(
        n10281) );
  NAND2_X1 U8806 ( .A1(n10281), .A2(n7551), .ZN(n7708) );
  OAI21_X1 U8807 ( .B1(n7551), .B2(n10281), .A(n7708), .ZN(n7554) );
  AND2_X1 U8808 ( .A1(P1_U3084), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n8358) );
  NOR2_X1 U8809 ( .A1(n8269), .A2(n7552), .ZN(n7553) );
  AOI211_X1 U8810 ( .C1(n10320), .C2(n7554), .A(n8358), .B(n7553), .ZN(n7561)
         );
  NOR2_X1 U8811 ( .A1(n10268), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n10271) );
  AOI21_X1 U8812 ( .B1(n7556), .B2(P1_REG2_REG_10__SCAN_IN), .A(n7555), .ZN(
        n10273) );
  NAND2_X1 U8813 ( .A1(n10268), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n10272) );
  OAI21_X1 U8814 ( .B1(n10271), .B2(n10273), .A(n10272), .ZN(n10270) );
  INV_X1 U8815 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n7557) );
  MUX2_X1 U8816 ( .A(n7557), .B(P1_REG2_REG_12__SCAN_IN), .S(n7709), .Z(n7558)
         );
  INV_X1 U8817 ( .A(n7558), .ZN(n7559) );
  NAND2_X1 U8818 ( .A1(n7559), .A2(n10270), .ZN(n7701) );
  OAI211_X1 U8819 ( .C1(n10270), .C2(n7559), .A(n10318), .B(n7701), .ZN(n7560)
         );
  OAI211_X1 U8820 ( .C1(n7562), .C2(n9736), .A(n7561), .B(n7560), .ZN(P1_U3253) );
  AOI211_X1 U8821 ( .C1(n7565), .C2(n7564), .A(n10357), .B(n7563), .ZN(n7576)
         );
  INV_X1 U8822 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n10191) );
  NAND2_X1 U8823 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3152), .ZN(n7566) );
  OAI21_X1 U8824 ( .B1(n8741), .B2(n10191), .A(n7566), .ZN(n7567) );
  INV_X1 U8825 ( .A(n7567), .ZN(n7573) );
  INV_X1 U8826 ( .A(n7568), .ZN(n7569) );
  OAI211_X1 U8827 ( .C1(n7571), .C2(n7570), .A(n10333), .B(n7569), .ZN(n7572)
         );
  OAI211_X1 U8828 ( .C1(n10335), .C2(n7574), .A(n7573), .B(n7572), .ZN(n7575)
         );
  OR2_X1 U8829 ( .A1(n7576), .A2(n7575), .ZN(P2_U3253) );
  XNOR2_X1 U8830 ( .A(n7578), .B(n7577), .ZN(n7585) );
  INV_X1 U8831 ( .A(n7791), .ZN(n7583) );
  OAI22_X1 U8832 ( .A1(n7579), .A2(n8660), .B1(n8662), .B2(n7821), .ZN(n7582)
         );
  OAI22_X1 U8833 ( .A1(n8683), .A2(n5285), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7580), .ZN(n7581) );
  AOI211_X1 U8834 ( .C1(n7583), .C2(n8665), .A(n7582), .B(n7581), .ZN(n7584)
         );
  OAI21_X1 U8835 ( .B1(n7585), .B2(n8669), .A(n7584), .ZN(P2_U3215) );
  INV_X1 U8836 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n7586) );
  OAI222_X1 U8837 ( .A1(n9300), .A2(n7586), .B1(n8219), .B2(n7587), .C1(n8038), 
        .C2(P2_U3152), .ZN(P2_U3344) );
  OAI222_X1 U8838 ( .A1(P1_U3084), .A2(n7712), .B1(n10119), .B2(n7588), .C1(
        n7587), .C2(n10113), .ZN(P1_U3339) );
  XOR2_X1 U8839 ( .A(n7590), .B(n7589), .Z(n7596) );
  OAI21_X1 U8840 ( .B1(n9392), .B2(P1_REG3_REG_3__SCAN_IN), .A(n7591), .ZN(
        n7594) );
  OAI22_X1 U8841 ( .A1(n9430), .A2(n7592), .B1(n9409), .B2(n7739), .ZN(n7593)
         );
  AOI211_X1 U8842 ( .C1(n9417), .C2(n10392), .A(n7594), .B(n7593), .ZN(n7595)
         );
  OAI21_X1 U8843 ( .B1(n7596), .B2(n9438), .A(n7595), .ZN(P1_U3216) );
  AOI22_X1 U8844 ( .A1(n7892), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n6480), .B2(
        n7609), .ZN(n7598) );
  OAI21_X1 U8845 ( .B1(n7599), .B2(n7598), .A(n7891), .ZN(n7600) );
  INV_X1 U8846 ( .A(n10357), .ZN(n10334) );
  NAND2_X1 U8847 ( .A1(n7600), .A2(n10334), .ZN(n7608) );
  NOR2_X1 U8848 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9215), .ZN(n7925) );
  AOI21_X1 U8849 ( .B1(n7602), .B2(P2_REG1_REG_10__SCAN_IN), .A(n7601), .ZN(
        n7605) );
  MUX2_X1 U8850 ( .A(n7603), .B(P2_REG1_REG_11__SCAN_IN), .S(n7892), .Z(n7604)
         );
  NOR2_X1 U8851 ( .A1(n7605), .A2(n7604), .ZN(n7883) );
  AOI211_X1 U8852 ( .C1(n7605), .C2(n7604), .A(n7883), .B(n10353), .ZN(n7606)
         );
  AOI211_X1 U8853 ( .C1(P2_ADDR_REG_11__SCAN_IN), .C2(n10352), .A(n7925), .B(
        n7606), .ZN(n7607) );
  OAI211_X1 U8854 ( .C1(n10335), .C2(n7609), .A(n7608), .B(n7607), .ZN(
        P2_U3256) );
  XNOR2_X1 U8855 ( .A(n7611), .B(n7610), .ZN(n7612) );
  XNOR2_X1 U8856 ( .A(n7613), .B(n7612), .ZN(n7618) );
  INV_X1 U8857 ( .A(n7875), .ZN(n7614) );
  NAND2_X1 U8858 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_U3084), .ZN(n7632) );
  OAI21_X1 U8859 ( .B1(n9392), .B2(n7614), .A(n7632), .ZN(n7616) );
  OAI22_X1 U8860 ( .A1(n9430), .A2(n7945), .B1(n9409), .B2(n4989), .ZN(n7615)
         );
  AOI211_X1 U8861 ( .C1(n9417), .C2(n9717), .A(n7616), .B(n7615), .ZN(n7617)
         );
  OAI21_X1 U8862 ( .B1(n7618), .B2(n9438), .A(n7617), .ZN(P1_U3228) );
  INV_X1 U8863 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n7619) );
  NAND2_X1 U8864 ( .A1(n10245), .A2(n7619), .ZN(n7620) );
  NAND2_X1 U8865 ( .A1(n7621), .A2(n7620), .ZN(n10243) );
  NOR2_X1 U8866 ( .A1(n7622), .A2(n10243), .ZN(n7623) );
  NOR2_X1 U8867 ( .A1(n10243), .A2(n10253), .ZN(n10248) );
  MUX2_X1 U8868 ( .A(n7623), .B(n10248), .S(n10245), .Z(n7624) );
  AOI211_X1 U8869 ( .C1(n10253), .C2(n10243), .A(n9719), .B(n7624), .ZN(n7651)
         );
  AOI21_X1 U8870 ( .B1(n7627), .B2(n7626), .A(n7625), .ZN(n7634) );
  OAI21_X1 U8871 ( .B1(n7630), .B2(n7629), .A(n7628), .ZN(n7631) );
  NAND2_X1 U8872 ( .A1(n10318), .A2(n7631), .ZN(n7633) );
  OAI211_X1 U8873 ( .C1(n7634), .C2(n10269), .A(n7633), .B(n7632), .ZN(n7638)
         );
  INV_X1 U8874 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n7635) );
  OAI22_X1 U8875 ( .A1(n8269), .A2(n7636), .B1(n7635), .B2(n9736), .ZN(n7637)
         );
  OR3_X1 U8876 ( .A1(n7651), .A2(n7638), .A3(n7637), .ZN(P1_U3245) );
  INV_X1 U8877 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n7639) );
  NOR2_X1 U8878 ( .A1(n9736), .A2(n7639), .ZN(n7650) );
  AOI211_X1 U8879 ( .C1(n7642), .C2(n7641), .A(n7640), .B(n10298), .ZN(n7649)
         );
  XOR2_X1 U8880 ( .A(n7644), .B(n7643), .Z(n7645) );
  AOI22_X1 U8881 ( .A1(n10320), .A2(n7645), .B1(P1_U3084), .B2(
        P1_REG3_REG_2__SCAN_IN), .ZN(n7646) );
  OAI21_X1 U8882 ( .B1(n8269), .B2(n7647), .A(n7646), .ZN(n7648) );
  OR4_X1 U8883 ( .A1(n7651), .A2(n7650), .A3(n7649), .A4(n7648), .ZN(P1_U3243)
         );
  NAND2_X1 U8884 ( .A1(n8781), .A2(P2_U3966), .ZN(n7652) );
  OAI21_X1 U8885 ( .B1(P2_U3966), .B2(n10118), .A(n7652), .ZN(P2_U3580) );
  OAI22_X1 U8886 ( .A1(n8777), .A2(n7654), .B1(n7653), .B2(n10454), .ZN(n7657)
         );
  NOR2_X1 U8887 ( .A1(n10466), .A2(n7655), .ZN(n7656) );
  AOI211_X1 U8888 ( .C1(n10466), .C2(P2_REG2_REG_1__SCAN_IN), .A(n7657), .B(
        n7656), .ZN(n7660) );
  INV_X1 U8889 ( .A(n8930), .ZN(n8943) );
  NAND2_X1 U8890 ( .A1(n8943), .A2(n7658), .ZN(n7659) );
  OAI211_X1 U8891 ( .C1(n8952), .C2(n7661), .A(n7660), .B(n7659), .ZN(P2_U3295) );
  OR2_X1 U8892 ( .A1(n10466), .A2(n7662), .ZN(n8061) );
  OAI22_X1 U8893 ( .A1(n8777), .A2(n7663), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        n10454), .ZN(n7664) );
  AOI21_X1 U8894 ( .B1(n8943), .B2(n7665), .A(n7664), .ZN(n7669) );
  MUX2_X1 U8895 ( .A(n7667), .B(n7666), .S(n8810), .Z(n7668) );
  OAI211_X1 U8896 ( .C1(n7670), .C2(n8061), .A(n7669), .B(n7668), .ZN(P2_U3293) );
  XNOR2_X1 U8897 ( .A(n7671), .B(n7672), .ZN(n10478) );
  INV_X1 U8898 ( .A(n10478), .ZN(n7684) );
  XNOR2_X1 U8899 ( .A(n7673), .B(n7672), .ZN(n7674) );
  OAI222_X1 U8900 ( .A1(n8673), .A2(n7719), .B1(n8675), .B2(n7675), .C1(n7674), 
        .C2(n8461), .ZN(n10476) );
  NAND2_X1 U8901 ( .A1(n10476), .A2(n8810), .ZN(n7683) );
  NOR2_X1 U8902 ( .A1(n8810), .A2(n7393), .ZN(n7680) );
  INV_X1 U8903 ( .A(n7681), .ZN(n10474) );
  INV_X1 U8904 ( .A(n7693), .ZN(n7677) );
  INV_X1 U8905 ( .A(n7794), .ZN(n7676) );
  OAI21_X1 U8906 ( .B1(n10474), .B2(n7677), .A(n7676), .ZN(n10475) );
  OAI22_X1 U8907 ( .A1(n8777), .A2(n10475), .B1(n7678), .B2(n10454), .ZN(n7679) );
  AOI211_X1 U8908 ( .C1(n8943), .C2(n7681), .A(n7680), .B(n7679), .ZN(n7682)
         );
  OAI211_X1 U8909 ( .C1(n7684), .C2(n8952), .A(n7683), .B(n7682), .ZN(P2_U3290) );
  OAI222_X1 U8910 ( .A1(P1_U3084), .A2(n8261), .B1(n10119), .B2(n7685), .C1(
        n7686), .C2(n10113), .ZN(P1_U3338) );
  OAI222_X1 U8911 ( .A1(n9300), .A2(n7687), .B1(n8219), .B2(n7686), .C1(n8708), 
        .C2(P2_U3152), .ZN(P2_U3343) );
  XNOR2_X1 U8912 ( .A(n7688), .B(n7689), .ZN(n10464) );
  XNOR2_X1 U8913 ( .A(n7691), .B(n7690), .ZN(n7692) );
  AOI222_X1 U8914 ( .A1(n8937), .A2(n7692), .B1(n7789), .B2(n8916), .C1(n8698), 
        .C2(n8915), .ZN(n10459) );
  OAI211_X1 U8915 ( .C1(n7759), .C2(n10456), .A(n10429), .B(n7693), .ZN(n10460) );
  OAI211_X1 U8916 ( .C1(n10456), .C2(n10536), .A(n10459), .B(n10460), .ZN(
        n7694) );
  AOI21_X1 U8917 ( .B1(n10464), .B2(n10541), .A(n7694), .ZN(n7698) );
  OR2_X1 U8918 ( .A1(n10553), .A2(n6399), .ZN(n7695) );
  OAI21_X1 U8919 ( .B1(n7698), .B2(n10551), .A(n7695), .ZN(P2_U3525) );
  INV_X1 U8920 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n7696) );
  OR2_X1 U8921 ( .A1(n10557), .A2(n7696), .ZN(n7697) );
  OAI21_X1 U8922 ( .B1(n7698), .B2(n10554), .A(n7697), .ZN(P2_U3466) );
  NAND2_X1 U8923 ( .A1(P1_REG2_REG_13__SCAN_IN), .A2(n10293), .ZN(n7703) );
  INV_X1 U8924 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n7699) );
  MUX2_X1 U8925 ( .A(n7699), .B(P1_REG2_REG_13__SCAN_IN), .S(n10293), .Z(n7700) );
  INV_X1 U8926 ( .A(n7700), .ZN(n10291) );
  NAND2_X1 U8927 ( .A1(P1_REG2_REG_12__SCAN_IN), .A2(n7709), .ZN(n7702) );
  NAND2_X1 U8928 ( .A1(n7702), .A2(n7701), .ZN(n10292) );
  NAND2_X1 U8929 ( .A1(n10291), .A2(n10292), .ZN(n10290) );
  NAND2_X1 U8930 ( .A1(n7703), .A2(n10290), .ZN(n8079) );
  INV_X1 U8931 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n7704) );
  NOR2_X1 U8932 ( .A1(n7712), .A2(n7704), .ZN(n8078) );
  AOI21_X1 U8933 ( .B1(n7704), .B2(n7712), .A(n8078), .ZN(n7705) );
  XNOR2_X1 U8934 ( .A(n8079), .B(n7705), .ZN(n7716) );
  INV_X1 U8935 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n7706) );
  AOI22_X1 U8936 ( .A1(P1_REG1_REG_13__SCAN_IN), .A2(n10293), .B1(n7707), .B2(
        n7706), .ZN(n10288) );
  OAI21_X1 U8937 ( .B1(P1_REG1_REG_12__SCAN_IN), .B2(n7709), .A(n7708), .ZN(
        n10287) );
  NAND2_X1 U8938 ( .A1(n10288), .A2(n10287), .ZN(n10286) );
  OAI21_X1 U8939 ( .B1(P1_REG1_REG_13__SCAN_IN), .B2(n10293), .A(n10286), .ZN(
        n7710) );
  INV_X1 U8940 ( .A(n7710), .ZN(n8074) );
  XNOR2_X1 U8941 ( .A(n8077), .B(P1_REG1_REG_14__SCAN_IN), .ZN(n8073) );
  XNOR2_X1 U8942 ( .A(n8074), .B(n8073), .ZN(n7711) );
  NAND2_X1 U8943 ( .A1(n7711), .A2(n10320), .ZN(n7715) );
  AND2_X1 U8944 ( .A1(P1_U3084), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n9309) );
  NOR2_X1 U8945 ( .A1(n8269), .A2(n7712), .ZN(n7713) );
  AOI211_X1 U8946 ( .C1(n10313), .C2(P1_ADDR_REG_14__SCAN_IN), .A(n9309), .B(
        n7713), .ZN(n7714) );
  OAI211_X1 U8947 ( .C1(n10298), .C2(n7716), .A(n7715), .B(n7714), .ZN(
        P1_U3255) );
  XOR2_X1 U8948 ( .A(n7718), .B(n7717), .Z(n7725) );
  OR2_X1 U8949 ( .A1(n7902), .A2(n8673), .ZN(n7721) );
  OR2_X1 U8950 ( .A1(n7719), .A2(n8675), .ZN(n7720) );
  NAND2_X1 U8951 ( .A1(n7721), .A2(n7720), .ZN(n7807) );
  AOI22_X1 U8952 ( .A1(n8680), .A2(n7807), .B1(P2_REG3_REG_8__SCAN_IN), .B2(
        P2_U3152), .ZN(n7723) );
  NAND2_X1 U8953 ( .A1(n8641), .A2(n7849), .ZN(n7722) );
  OAI211_X1 U8954 ( .C1(n8678), .C2(n7851), .A(n7723), .B(n7722), .ZN(n7724)
         );
  AOI21_X1 U8955 ( .B1(n7725), .B2(n8657), .A(n7724), .ZN(n7726) );
  INV_X1 U8956 ( .A(n7726), .ZN(P2_U3223) );
  NAND2_X1 U8957 ( .A1(n7727), .A2(n9652), .ZN(n7868) );
  OAI21_X1 U8958 ( .B1(n9652), .B2(n7727), .A(n7868), .ZN(n7733) );
  OAI21_X1 U8959 ( .B1(n7730), .B2(n7729), .A(n7728), .ZN(n7741) );
  INV_X1 U8960 ( .A(n7741), .ZN(n7780) );
  AOI22_X1 U8961 ( .A1(n10393), .A2(n10392), .B1(n9716), .B2(n10391), .ZN(
        n7731) );
  OAI21_X1 U8962 ( .B1(n7780), .B2(n10401), .A(n7731), .ZN(n7732) );
  AOI21_X1 U8963 ( .B1(n10397), .B2(n7733), .A(n7732), .ZN(n7779) );
  NAND2_X1 U8964 ( .A1(n7734), .A2(n10411), .ZN(n7735) );
  INV_X1 U8965 ( .A(n9779), .ZN(n10415) );
  AOI21_X1 U8966 ( .B1(n7776), .B2(n8576), .A(n4986), .ZN(n7777) );
  NAND2_X1 U8967 ( .A1(n7777), .A2(n10368), .ZN(n7738) );
  AOI22_X1 U8968 ( .A1(n10371), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n10409), .B2(
        n7736), .ZN(n7737) );
  OAI211_X1 U8969 ( .C1(n7739), .C2(n9969), .A(n7738), .B(n7737), .ZN(n7740)
         );
  AOI21_X1 U8970 ( .B1(n10415), .B2(n7741), .A(n7740), .ZN(n7742) );
  OAI21_X1 U8971 ( .B1(n7779), .B2(n10371), .A(n7742), .ZN(P1_U3288) );
  XOR2_X1 U8972 ( .A(n7745), .B(n7744), .Z(n7746) );
  XNOR2_X1 U8973 ( .A(n7743), .B(n7746), .ZN(n7751) );
  NAND2_X1 U8974 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3084), .ZN(n10325) );
  OAI21_X1 U8975 ( .B1(n9392), .B2(n7747), .A(n10325), .ZN(n7749) );
  OAI22_X1 U8976 ( .A1(n9430), .A2(n7979), .B1(n9409), .B2(n7936), .ZN(n7748)
         );
  AOI211_X1 U8977 ( .C1(n9417), .C2(n9716), .A(n7749), .B(n7748), .ZN(n7750)
         );
  OAI21_X1 U8978 ( .B1(n7751), .B2(n9438), .A(n7750), .ZN(P1_U3225) );
  OAI211_X1 U8979 ( .C1(n7753), .C2(n7767), .A(n7752), .B(n8937), .ZN(n7755)
         );
  AOI22_X1 U8980 ( .A1(n7296), .A2(n8915), .B1(n8916), .B2(n8697), .ZN(n7754)
         );
  NAND2_X1 U8981 ( .A1(n7755), .A2(n7754), .ZN(n10448) );
  NOR2_X1 U8982 ( .A1(n8810), .A2(n7756), .ZN(n7762) );
  NOR2_X1 U8983 ( .A1(n7757), .A2(n10445), .ZN(n7758) );
  OR2_X1 U8984 ( .A1(n7759), .A2(n7758), .ZN(n10446) );
  OAI22_X1 U8985 ( .A1(n8777), .A2(n10446), .B1(n7760), .B2(n10454), .ZN(n7761) );
  AOI211_X1 U8986 ( .C1(n8810), .C2(n10448), .A(n7762), .B(n7761), .ZN(n7770)
         );
  AND2_X1 U8987 ( .A1(n7764), .A2(n7763), .ZN(n7766) );
  NOR2_X1 U8988 ( .A1(n7766), .A2(n7767), .ZN(n7765) );
  AOI21_X1 U8989 ( .B1(n7767), .B2(n7766), .A(n7765), .ZN(n10449) );
  AOI22_X1 U8990 ( .A1(n10449), .A2(n8933), .B1(n8943), .B2(n7768), .ZN(n7769)
         );
  NAND2_X1 U8991 ( .A1(n7770), .A2(n7769), .ZN(P2_U3292) );
  INV_X1 U8992 ( .A(n10379), .ZN(n7774) );
  AOI22_X1 U8993 ( .A1(n10379), .A2(n8937), .B1(n8699), .B2(n8916), .ZN(n10381) );
  OAI22_X1 U8994 ( .A1(n10466), .A2(n10381), .B1(n7294), .B2(n10454), .ZN(
        n7771) );
  AOI21_X1 U8995 ( .B1(P2_REG2_REG_0__SCAN_IN), .B2(n10466), .A(n7771), .ZN(
        n7773) );
  OAI21_X1 U8996 ( .B1(n8943), .B2(n8926), .A(n10377), .ZN(n7772) );
  OAI211_X1 U8997 ( .C1(n7774), .C2(n8952), .A(n7773), .B(n7772), .ZN(P2_U3296) );
  AOI22_X1 U8998 ( .A1(n7777), .A2(n10386), .B1(n10502), .B2(n7776), .ZN(n7778) );
  OAI211_X1 U8999 ( .C1(n7780), .C2(n10504), .A(n7779), .B(n7778), .ZN(n7782)
         );
  NAND2_X1 U9000 ( .A1(n7782), .A2(n10531), .ZN(n7781) );
  OAI21_X1 U9001 ( .B1(n10531), .B2(n7187), .A(n7781), .ZN(P1_U3526) );
  INV_X1 U9002 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n7784) );
  NAND2_X1 U9003 ( .A1(n7782), .A2(n10535), .ZN(n7783) );
  OAI21_X1 U9004 ( .B1(n10535), .B2(n7784), .A(n7783), .ZN(P1_U3463) );
  XNOR2_X1 U9005 ( .A(n7786), .B(n7785), .ZN(n7863) );
  XNOR2_X1 U9006 ( .A(n7788), .B(n7787), .ZN(n7790) );
  AOI222_X1 U9007 ( .A1(n8937), .A2(n7790), .B1(n8694), .B2(n8916), .C1(n7789), 
        .C2(n8915), .ZN(n7862) );
  INV_X1 U9008 ( .A(n7862), .ZN(n7799) );
  OAI22_X1 U9009 ( .A1(n8810), .A2(n7792), .B1(n7791), .B2(n10454), .ZN(n7793)
         );
  INV_X1 U9010 ( .A(n7793), .ZN(n7797) );
  OR2_X1 U9011 ( .A1(n5285), .A2(n7794), .ZN(n7795) );
  AND2_X1 U9012 ( .A1(n7809), .A2(n7795), .ZN(n7860) );
  NAND2_X1 U9013 ( .A1(n8926), .A2(n7860), .ZN(n7796) );
  OAI211_X1 U9014 ( .C1(n5285), .C2(n8930), .A(n7797), .B(n7796), .ZN(n7798)
         );
  AOI21_X1 U9015 ( .B1(n7799), .B2(n8810), .A(n7798), .ZN(n7800) );
  OAI21_X1 U9016 ( .B1(n8952), .B2(n7863), .A(n7800), .ZN(P2_U3289) );
  INV_X1 U9017 ( .A(n7801), .ZN(n7898) );
  AOI22_X1 U9018 ( .A1(n8723), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_16__SCAN_IN), .B2(n9297), .ZN(n7802) );
  OAI21_X1 U9019 ( .B1(n7898), .B2(n8219), .A(n7802), .ZN(P2_U3342) );
  INV_X1 U9020 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n7813) );
  OAI21_X1 U9021 ( .B1(n7803), .B2(n6442), .A(n7804), .ZN(n7846) );
  XNOR2_X1 U9022 ( .A(n7806), .B(n7805), .ZN(n7808) );
  AOI21_X1 U9023 ( .B1(n7808), .B2(n8937), .A(n7807), .ZN(n7858) );
  AOI21_X1 U9024 ( .B1(n7849), .B2(n7809), .A(n10545), .ZN(n7810) );
  AND2_X1 U9025 ( .A1(n7810), .A2(n8056), .ZN(n7847) );
  AOI21_X1 U9026 ( .B1(n10550), .B2(n7849), .A(n7847), .ZN(n7811) );
  OAI211_X1 U9027 ( .C1(n7846), .C2(n9271), .A(n7858), .B(n7811), .ZN(n7814)
         );
  NAND2_X1 U9028 ( .A1(n7814), .A2(n10557), .ZN(n7812) );
  OAI21_X1 U9029 ( .B1(n10557), .B2(n7813), .A(n7812), .ZN(P2_U3475) );
  NAND2_X1 U9030 ( .A1(n7814), .A2(n10553), .ZN(n7815) );
  OAI21_X1 U9031 ( .B1(n10553), .B2(n6437), .A(n7815), .ZN(P2_U3528) );
  OAI21_X1 U9032 ( .B1(n7818), .B2(n7817), .A(n7816), .ZN(n7819) );
  NAND2_X1 U9033 ( .A1(n7819), .A2(n8657), .ZN(n7825) );
  INV_X1 U9034 ( .A(n7820), .ZN(n7823) );
  OAI22_X1 U9035 ( .A1(n8057), .A2(n8678), .B1(n8660), .B2(n7821), .ZN(n7822)
         );
  AOI211_X1 U9036 ( .C1(n8647), .C2(n8692), .A(n7823), .B(n7822), .ZN(n7824)
         );
  OAI211_X1 U9037 ( .C1(n5121), .C2(n8683), .A(n7825), .B(n7824), .ZN(P2_U3233) );
  INV_X1 U9038 ( .A(n7826), .ZN(n7833) );
  NAND2_X1 U9039 ( .A1(n7827), .A2(n7833), .ZN(n7828) );
  NAND2_X1 U9040 ( .A1(n7468), .A2(n7828), .ZN(n10428) );
  NAND2_X1 U9041 ( .A1(n10428), .A2(n7829), .ZN(n7838) );
  OAI22_X1 U9042 ( .A1(n7045), .A2(n8675), .B1(n7830), .B2(n8673), .ZN(n7831)
         );
  INV_X1 U9043 ( .A(n7831), .ZN(n7837) );
  OAI21_X1 U9044 ( .B1(n7833), .B2(n7832), .A(n8937), .ZN(n7834) );
  OR2_X1 U9045 ( .A1(n7835), .A2(n7834), .ZN(n7836) );
  INV_X1 U9046 ( .A(n8061), .ZN(n7839) );
  AOI22_X1 U9047 ( .A1(n7839), .A2(n10428), .B1(n8943), .B2(n7054), .ZN(n7845)
         );
  NAND2_X1 U9048 ( .A1(n7840), .A2(n7054), .ZN(n7841) );
  AND2_X1 U9049 ( .A1(n7842), .A2(n7841), .ZN(n10430) );
  OAI22_X1 U9050 ( .A1(n7390), .A2(n8810), .B1(n9219), .B2(n10454), .ZN(n7843)
         );
  AOI21_X1 U9051 ( .B1(n8926), .B2(n10430), .A(n7843), .ZN(n7844) );
  OAI211_X1 U9052 ( .C1(n10466), .C2(n10432), .A(n7845), .B(n7844), .ZN(
        P2_U3294) );
  NOR2_X1 U9053 ( .A1(n7846), .A2(n8952), .ZN(n7856) );
  INV_X1 U9054 ( .A(n7847), .ZN(n7848) );
  NAND2_X1 U9055 ( .A1(n8810), .A2(n8008), .ZN(n8909) );
  NOR2_X1 U9056 ( .A1(n7848), .A2(n8909), .ZN(n7855) );
  INV_X1 U9057 ( .A(n7849), .ZN(n7850) );
  NOR2_X1 U9058 ( .A1(n8930), .A2(n7850), .ZN(n7854) );
  OAI22_X1 U9059 ( .A1(n8810), .A2(n7852), .B1(n7851), .B2(n10454), .ZN(n7853)
         );
  NOR4_X1 U9060 ( .A1(n7856), .A2(n7855), .A3(n7854), .A4(n7853), .ZN(n7857)
         );
  OAI21_X1 U9061 ( .B1(n10466), .B2(n7858), .A(n7857), .ZN(P2_U3288) );
  INV_X1 U9062 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n7865) );
  AOI22_X1 U9063 ( .A1(n7860), .A2(n10429), .B1(n10550), .B2(n7859), .ZN(n7861) );
  OAI211_X1 U9064 ( .C1(n9271), .C2(n7863), .A(n7862), .B(n7861), .ZN(n7866)
         );
  NAND2_X1 U9065 ( .A1(n7866), .A2(n10557), .ZN(n7864) );
  OAI21_X1 U9066 ( .B1(n10557), .B2(n7865), .A(n7864), .ZN(P2_U3472) );
  NAND2_X1 U9067 ( .A1(n7866), .A2(n10553), .ZN(n7867) );
  OAI21_X1 U9068 ( .B1(n10553), .B2(n6424), .A(n7867), .ZN(P2_U3527) );
  XNOR2_X1 U9069 ( .A(n7869), .B(n9651), .ZN(n7870) );
  INV_X1 U9070 ( .A(n10397), .ZN(n9972) );
  OAI222_X1 U9071 ( .A1(n9975), .A2(n7945), .B1(n9977), .B2(n8580), .C1(n7870), 
        .C2(n9972), .ZN(n10438) );
  INV_X1 U9072 ( .A(n10438), .ZN(n7882) );
  OAI21_X1 U9073 ( .B1(n7872), .B2(n9651), .A(n7871), .ZN(n10440) );
  INV_X1 U9074 ( .A(n9985), .ZN(n7880) );
  AND2_X1 U9075 ( .A1(n7873), .A2(n7876), .ZN(n7874) );
  OR2_X1 U9076 ( .A1(n7874), .A2(n7931), .ZN(n10437) );
  AOI22_X1 U9077 ( .A1(n10371), .A2(P1_REG2_REG_4__SCAN_IN), .B1(n7875), .B2(
        n10409), .ZN(n7878) );
  NAND2_X1 U9078 ( .A1(n10367), .A2(n7876), .ZN(n7877) );
  OAI211_X1 U9079 ( .C1(n10437), .C2(n9918), .A(n7878), .B(n7877), .ZN(n7879)
         );
  AOI21_X1 U9080 ( .B1(n10440), .B2(n7880), .A(n7879), .ZN(n7881) );
  OAI21_X1 U9081 ( .B1(n7882), .B2(n10371), .A(n7881), .ZN(P1_U3287) );
  INV_X1 U9082 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n7889) );
  MUX2_X1 U9083 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n7884), .S(n7964), .Z(n7885)
         );
  NAND2_X1 U9084 ( .A1(n7886), .A2(n7885), .ZN(n7958) );
  OAI21_X1 U9085 ( .B1(n7886), .B2(n7885), .A(n7958), .ZN(n7887) );
  NAND2_X1 U9086 ( .A1(n10333), .A2(n7887), .ZN(n7888) );
  NAND2_X1 U9087 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3152), .ZN(n8122) );
  OAI211_X1 U9088 ( .C1(n8741), .C2(n7889), .A(n7888), .B(n8122), .ZN(n7896)
         );
  MUX2_X1 U9089 ( .A(P2_REG2_REG_12__SCAN_IN), .B(n8137), .S(n7964), .Z(n7890)
         );
  INV_X1 U9090 ( .A(n7890), .ZN(n7894) );
  NOR2_X1 U9091 ( .A1(n7893), .A2(n7894), .ZN(n7963) );
  AOI211_X1 U9092 ( .C1(n7894), .C2(n7893), .A(n10357), .B(n7963), .ZN(n7895)
         );
  AOI211_X1 U9093 ( .C1(n10364), .C2(n7964), .A(n7896), .B(n7895), .ZN(n7897)
         );
  INV_X1 U9094 ( .A(n7897), .ZN(P2_U3257) );
  INV_X1 U9095 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n7899) );
  INV_X1 U9096 ( .A(n8295), .ZN(n8268) );
  OAI222_X1 U9097 ( .A1(n10119), .A2(n7899), .B1(n10113), .B2(n7898), .C1(
        P1_U3084), .C2(n8268), .ZN(P1_U3337) );
  XNOR2_X1 U9098 ( .A(n7900), .B(n7901), .ZN(n7906) );
  OAI22_X1 U9099 ( .A1(n8662), .A2(n8130), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6467), .ZN(n7904) );
  OAI22_X1 U9100 ( .A1(n7992), .A2(n8678), .B1(n8660), .B2(n7902), .ZN(n7903)
         );
  AOI211_X1 U9101 ( .C1(n8641), .C2(n10512), .A(n7904), .B(n7903), .ZN(n7905)
         );
  OAI21_X1 U9102 ( .B1(n7906), .B2(n8669), .A(n7905), .ZN(P2_U3219) );
  NAND2_X1 U9103 ( .A1(n7908), .A2(n7907), .ZN(n7972) );
  INV_X1 U9104 ( .A(n7973), .ZN(n7909) );
  NOR2_X1 U9105 ( .A1(n7909), .A2(n7971), .ZN(n7910) );
  XNOR2_X1 U9106 ( .A(n7972), .B(n7910), .ZN(n7915) );
  AOI22_X1 U9107 ( .A1(n9416), .A2(n9713), .B1(n9435), .B2(n7952), .ZN(n7914)
         );
  INV_X1 U9108 ( .A(n9392), .ZN(n9434) );
  NAND2_X1 U9109 ( .A1(P1_U3084), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n10266) );
  INV_X1 U9110 ( .A(n10266), .ZN(n7912) );
  NOR2_X1 U9111 ( .A1(n9431), .A2(n7945), .ZN(n7911) );
  AOI211_X1 U9112 ( .C1(n9434), .C2(n7951), .A(n7912), .B(n7911), .ZN(n7913)
         );
  OAI211_X1 U9113 ( .C1(n7915), .C2(n9438), .A(n7914), .B(n7913), .ZN(P1_U3237) );
  INV_X1 U9114 ( .A(n7916), .ZN(n7919) );
  AOI22_X1 U9115 ( .A1(n8738), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_17__SCAN_IN), .B2(n9297), .ZN(n7917) );
  OAI21_X1 U9116 ( .B1(n7919), .B2(n8219), .A(n7917), .ZN(P2_U3341) );
  AOI22_X1 U9117 ( .A1(n9727), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n10107), .ZN(n7918) );
  OAI21_X1 U9118 ( .B1(n7919), .B2(n10113), .A(n7918), .ZN(P1_U3336) );
  XNOR2_X1 U9119 ( .A(n7921), .B(n7920), .ZN(n7929) );
  OR2_X1 U9120 ( .A1(n8211), .A2(n8673), .ZN(n7924) );
  OR2_X1 U9121 ( .A1(n7922), .A2(n8675), .ZN(n7923) );
  NAND2_X1 U9122 ( .A1(n7924), .A2(n7923), .ZN(n8093) );
  AOI21_X1 U9123 ( .B1(n8680), .B2(n8093), .A(n7925), .ZN(n7926) );
  OAI21_X1 U9124 ( .B1(n8678), .B2(n8171), .A(n7926), .ZN(n7927) );
  AOI21_X1 U9125 ( .B1(n8641), .B2(n8098), .A(n7927), .ZN(n7928) );
  OAI21_X1 U9126 ( .B1(n7929), .B2(n8669), .A(n7928), .ZN(P2_U3238) );
  NAND2_X1 U9127 ( .A1(n9451), .A2(n9653), .ZN(n7942) );
  OAI21_X1 U9128 ( .B1(n9653), .B2(n9451), .A(n7942), .ZN(n7930) );
  AOI222_X1 U9129 ( .A1(n10397), .A2(n7930), .B1(n9714), .B2(n10391), .C1(
        n9716), .C2(n10393), .ZN(n8067) );
  INV_X1 U9130 ( .A(n7931), .ZN(n7932) );
  AOI211_X1 U9131 ( .C1(n8065), .C2(n7932), .A(n10522), .B(n7949), .ZN(n8064)
         );
  NOR2_X1 U9132 ( .A1(n7933), .A2(n10411), .ZN(n9983) );
  AOI22_X1 U9133 ( .A1(n10371), .A2(P1_REG2_REG_5__SCAN_IN), .B1(n7934), .B2(
        n10409), .ZN(n7935) );
  OAI21_X1 U9134 ( .B1(n9969), .B2(n7936), .A(n7935), .ZN(n7940) );
  OAI21_X1 U9135 ( .B1(n7938), .B2(n6213), .A(n7937), .ZN(n8068) );
  NOR2_X1 U9136 ( .A1(n8068), .A2(n9985), .ZN(n7939) );
  AOI211_X1 U9137 ( .C1(n8064), .C2(n9983), .A(n7940), .B(n7939), .ZN(n7941)
         );
  OAI21_X1 U9138 ( .B1(n8067), .B2(n10371), .A(n7941), .ZN(P1_U3286) );
  NAND2_X1 U9139 ( .A1(n7942), .A2(n9455), .ZN(n7943) );
  XNOR2_X1 U9140 ( .A(n7943), .B(n9656), .ZN(n7948) );
  OAI21_X1 U9141 ( .B1(n4918), .B2(n9656), .A(n7944), .ZN(n10471) );
  OAI22_X1 U9142 ( .A1(n7945), .A2(n9977), .B1(n8020), .B2(n9975), .ZN(n7946)
         );
  AOI21_X1 U9143 ( .B1(n10471), .B2(n6266), .A(n7946), .ZN(n7947) );
  OAI21_X1 U9144 ( .B1(n9972), .B2(n7948), .A(n7947), .ZN(n10469) );
  INV_X1 U9145 ( .A(n10469), .ZN(n7957) );
  OR2_X1 U9146 ( .A1(n7949), .A2(n10467), .ZN(n7950) );
  NAND2_X1 U9147 ( .A1(n8107), .A2(n7950), .ZN(n10468) );
  AOI22_X1 U9148 ( .A1(n10371), .A2(P1_REG2_REG_6__SCAN_IN), .B1(n7951), .B2(
        n10409), .ZN(n7954) );
  NAND2_X1 U9149 ( .A1(n10367), .A2(n7952), .ZN(n7953) );
  OAI211_X1 U9150 ( .C1(n10468), .C2(n9918), .A(n7954), .B(n7953), .ZN(n7955)
         );
  AOI21_X1 U9151 ( .B1(n10471), .B2(n10415), .A(n7955), .ZN(n7956) );
  OAI21_X1 U9152 ( .B1(n7957), .B2(n10371), .A(n7956), .ZN(P1_U3285) );
  INV_X1 U9153 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n7962) );
  NAND2_X1 U9154 ( .A1(n8037), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n8027) );
  OAI21_X1 U9155 ( .B1(n8037), .B2(P2_REG1_REG_13__SCAN_IN), .A(n8027), .ZN(
        n7959) );
  OAI21_X1 U9156 ( .B1(n7964), .B2(P2_REG1_REG_12__SCAN_IN), .A(n7958), .ZN(
        n8026) );
  XOR2_X1 U9157 ( .A(n7959), .B(n8026), .Z(n7960) );
  NAND2_X1 U9158 ( .A1(n10333), .A2(n7960), .ZN(n7961) );
  NAND2_X1 U9159 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(P2_U3152), .ZN(n8210) );
  OAI211_X1 U9160 ( .C1(n8741), .C2(n7962), .A(n7961), .B(n8210), .ZN(n7969)
         );
  MUX2_X1 U9161 ( .A(P2_REG2_REG_13__SCAN_IN), .B(n8239), .S(n8037), .Z(n7965)
         );
  INV_X1 U9162 ( .A(n7965), .ZN(n7966) );
  AOI211_X1 U9163 ( .C1(n7967), .C2(n7966), .A(n10357), .B(n8036), .ZN(n7968)
         );
  AOI211_X1 U9164 ( .C1(n10364), .C2(n8037), .A(n7969), .B(n7968), .ZN(n7970)
         );
  INV_X1 U9165 ( .A(n7970), .ZN(P2_U3258) );
  OR2_X1 U9166 ( .A1(n7972), .A2(n7971), .ZN(n7974) );
  NAND2_X1 U9167 ( .A1(n7974), .A2(n7973), .ZN(n7975) );
  XOR2_X1 U9168 ( .A(n7976), .B(n7975), .Z(n7983) );
  OAI21_X1 U9169 ( .B1(n9392), .B2(n7978), .A(n7977), .ZN(n7981) );
  OAI22_X1 U9170 ( .A1(n7979), .A2(n9431), .B1(n9430), .B2(n8184), .ZN(n7980)
         );
  AOI211_X1 U9171 ( .C1(n8162), .C2(n9435), .A(n7981), .B(n7980), .ZN(n7982)
         );
  OAI21_X1 U9172 ( .B1(n7983), .B2(n9438), .A(n7982), .ZN(P1_U3211) );
  OAI21_X1 U9173 ( .B1(n7985), .B2(n7988), .A(n7984), .ZN(n10511) );
  AOI22_X1 U9174 ( .A1(n8915), .A2(n8693), .B1(n7986), .B2(n8916), .ZN(n7991)
         );
  XOR2_X1 U9175 ( .A(n7988), .B(n7987), .Z(n7989) );
  NAND2_X1 U9176 ( .A1(n7989), .A2(n8937), .ZN(n7990) );
  OAI211_X1 U9177 ( .C1(n10511), .C2(n8051), .A(n7991), .B(n7990), .ZN(n10515)
         );
  NAND2_X1 U9178 ( .A1(n10515), .A2(n8810), .ZN(n7998) );
  OAI22_X1 U9179 ( .A1(n8810), .A2(n7993), .B1(n7992), .B2(n10454), .ZN(n7996)
         );
  AND2_X1 U9180 ( .A1(n10512), .A2(n8054), .ZN(n7994) );
  OR2_X1 U9181 ( .A1(n8095), .A2(n7994), .ZN(n10514) );
  NOR2_X1 U9182 ( .A1(n10514), .A2(n8777), .ZN(n7995) );
  AOI211_X1 U9183 ( .C1(n8943), .C2(n10512), .A(n7996), .B(n7995), .ZN(n7997)
         );
  OAI211_X1 U9184 ( .C1(n10511), .C2(n8061), .A(n7998), .B(n7997), .ZN(
        P2_U3286) );
  XOR2_X1 U9185 ( .A(n7999), .B(n8000), .Z(n8006) );
  INV_X1 U9186 ( .A(n8001), .ZN(n8188) );
  AOI22_X1 U9187 ( .A1(n9417), .A2(n8105), .B1(n9416), .B2(n9711), .ZN(n8003)
         );
  OAI211_X1 U9188 ( .C1(n8188), .C2(n9392), .A(n8003), .B(n8002), .ZN(n8004)
         );
  AOI21_X1 U9189 ( .B1(n10490), .B2(n9435), .A(n8004), .ZN(n8005) );
  OAI21_X1 U9190 ( .B1(n8006), .B2(n9438), .A(n8005), .ZN(P1_U3229) );
  INV_X1 U9191 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n8009) );
  INV_X1 U9192 ( .A(n8007), .ZN(n8010) );
  OAI222_X1 U9193 ( .A1(n9300), .A2(n8009), .B1(n8219), .B2(n8010), .C1(n8008), 
        .C2(P2_U3152), .ZN(P2_U3339) );
  INV_X1 U9194 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n8011) );
  OAI222_X1 U9195 ( .A1(n10119), .A2(n8011), .B1(n10113), .B2(n8010), .C1(
        P1_U3084), .C2(n9856), .ZN(P1_U3334) );
  INV_X1 U9196 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n8013) );
  INV_X1 U9197 ( .A(n8012), .ZN(n8014) );
  INV_X1 U9198 ( .A(n10304), .ZN(n9721) );
  OAI222_X1 U9199 ( .A1(n10119), .A2(n8013), .B1(n10113), .B2(n8014), .C1(
        n9721), .C2(P1_U3084), .ZN(P1_U3335) );
  INV_X1 U9200 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n8015) );
  INV_X1 U9201 ( .A(n8736), .ZN(n8753) );
  OAI222_X1 U9202 ( .A1(n9300), .A2(n8015), .B1(n8219), .B2(n8014), .C1(n8753), 
        .C2(P2_U3152), .ZN(P2_U3340) );
  NAND2_X1 U9203 ( .A1(n8016), .A2(n8017), .ZN(n8019) );
  XNOR2_X1 U9204 ( .A(n8019), .B(n8018), .ZN(n8025) );
  OAI22_X1 U9205 ( .A1(n8020), .A2(n9431), .B1(n9430), .B2(n8276), .ZN(n8021)
         );
  AOI211_X1 U9206 ( .C1(n9434), .C2(n8154), .A(n8022), .B(n8021), .ZN(n8024)
         );
  NAND2_X1 U9207 ( .A1(n9435), .A2(n8155), .ZN(n8023) );
  OAI211_X1 U9208 ( .C1(n8025), .C2(n9438), .A(n8024), .B(n8023), .ZN(P1_U3219) );
  AOI22_X1 U9209 ( .A1(n8028), .A2(n6508), .B1(n8027), .B2(n8026), .ZN(n8031)
         );
  NAND2_X1 U9210 ( .A1(n8038), .A2(n8029), .ZN(n8030) );
  OAI21_X1 U9211 ( .B1(n8031), .B2(n8030), .A(n8701), .ZN(n8033) );
  NAND3_X1 U9212 ( .A1(n8312), .A2(P2_REG1_REG_14__SCAN_IN), .A3(n8031), .ZN(
        n8032) );
  AND2_X1 U9213 ( .A1(n8033), .A2(n8032), .ZN(n8044) );
  NOR2_X1 U9214 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6522), .ZN(n8307) );
  INV_X1 U9215 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n8034) );
  NOR2_X1 U9216 ( .A1(n8741), .A2(n8034), .ZN(n8035) );
  AOI211_X1 U9217 ( .C1(n8312), .C2(n10364), .A(n8307), .B(n8035), .ZN(n8043)
         );
  AOI22_X1 U9218 ( .A1(n8312), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n6526), .B2(
        n8038), .ZN(n8039) );
  OAI21_X1 U9219 ( .B1(n8040), .B2(n8039), .A(n8311), .ZN(n8041) );
  NAND2_X1 U9220 ( .A1(n8041), .A2(n10334), .ZN(n8042) );
  OAI211_X1 U9221 ( .C1(n8044), .C2(n10353), .A(n8043), .B(n8042), .ZN(
        P2_U3259) );
  XNOR2_X1 U9222 ( .A(n8045), .B(n8049), .ZN(n8053) );
  INV_X1 U9223 ( .A(n8046), .ZN(n8047) );
  AOI21_X1 U9224 ( .B1(n8049), .B2(n8048), .A(n8047), .ZN(n8200) );
  AOI22_X1 U9225 ( .A1(n8692), .A2(n8916), .B1(n8915), .B2(n8694), .ZN(n8050)
         );
  OAI21_X1 U9226 ( .B1(n8200), .B2(n8051), .A(n8050), .ZN(n8052) );
  AOI21_X1 U9227 ( .B1(n8053), .B2(n8937), .A(n8052), .ZN(n8199) );
  INV_X1 U9228 ( .A(n8054), .ZN(n8055) );
  AOI21_X1 U9229 ( .B1(n8196), .B2(n8056), .A(n8055), .ZN(n8197) );
  OAI22_X1 U9230 ( .A1(n8810), .A2(n8058), .B1(n8057), .B2(n10454), .ZN(n8060)
         );
  NOR2_X1 U9231 ( .A1(n8930), .A2(n5121), .ZN(n8059) );
  AOI211_X1 U9232 ( .C1(n8197), .C2(n8926), .A(n8060), .B(n8059), .ZN(n8063)
         );
  OR2_X1 U9233 ( .A1(n8200), .A2(n8061), .ZN(n8062) );
  OAI211_X1 U9234 ( .C1(n8199), .C2(n10466), .A(n8063), .B(n8062), .ZN(
        P2_U3287) );
  AOI21_X1 U9235 ( .B1(n10502), .B2(n8065), .A(n8064), .ZN(n8066) );
  OAI211_X1 U9236 ( .C1(n10436), .C2(n8068), .A(n8067), .B(n8066), .ZN(n8070)
         );
  NAND2_X1 U9237 ( .A1(n8070), .A2(n10531), .ZN(n8069) );
  OAI21_X1 U9238 ( .B1(n10531), .B2(n7189), .A(n8069), .ZN(P1_U3528) );
  INV_X1 U9239 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n8072) );
  NAND2_X1 U9240 ( .A1(n8070), .A2(n10535), .ZN(n8071) );
  OAI21_X1 U9241 ( .B1(n10535), .B2(n8072), .A(n8071), .ZN(P1_U3469) );
  OAI22_X1 U9242 ( .A1(n8074), .A2(n8073), .B1(P1_REG1_REG_14__SCAN_IN), .B2(
        n8077), .ZN(n8255) );
  XNOR2_X1 U9243 ( .A(n8255), .B(n8261), .ZN(n8076) );
  INV_X1 U9244 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n8075) );
  NOR2_X1 U9245 ( .A1(n8075), .A2(n8076), .ZN(n8256) );
  AOI211_X1 U9246 ( .C1(n8076), .C2(n8075), .A(n8256), .B(n10269), .ZN(n8088)
         );
  OAI22_X1 U9247 ( .A1(n8079), .A2(n8078), .B1(P1_REG2_REG_14__SCAN_IN), .B2(
        n8077), .ZN(n8260) );
  XNOR2_X1 U9248 ( .A(n8260), .B(n8261), .ZN(n8081) );
  INV_X1 U9249 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n8080) );
  NOR2_X1 U9250 ( .A1(n8080), .A2(n8081), .ZN(n8262) );
  AOI211_X1 U9251 ( .C1(n8081), .C2(n8080), .A(n8262), .B(n10298), .ZN(n8087)
         );
  INV_X1 U9252 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n8085) );
  NOR2_X1 U9253 ( .A1(n8082), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9433) );
  AOI21_X1 U9254 ( .B1(n10312), .B2(n8083), .A(n9433), .ZN(n8084) );
  OAI21_X1 U9255 ( .B1(n9736), .B2(n8085), .A(n8084), .ZN(n8086) );
  OR3_X1 U9256 ( .A1(n8088), .A2(n8087), .A3(n8086), .ZN(P1_U3256) );
  INV_X1 U9257 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n8101) );
  XNOR2_X1 U9258 ( .A(n8090), .B(n8089), .ZN(n8175) );
  XNOR2_X1 U9259 ( .A(n8092), .B(n8091), .ZN(n8094) );
  AOI21_X1 U9260 ( .B1(n8094), .B2(n8937), .A(n8093), .ZN(n8180) );
  INV_X1 U9261 ( .A(n8095), .ZN(n8097) );
  INV_X1 U9262 ( .A(n8134), .ZN(n8096) );
  AOI211_X1 U9263 ( .C1(n8098), .C2(n8097), .A(n10545), .B(n8096), .ZN(n8178)
         );
  AOI21_X1 U9264 ( .B1(n10550), .B2(n8098), .A(n8178), .ZN(n8099) );
  OAI211_X1 U9265 ( .C1(n8175), .C2(n9271), .A(n8180), .B(n8099), .ZN(n8102)
         );
  NAND2_X1 U9266 ( .A1(n8102), .A2(n10557), .ZN(n8100) );
  OAI21_X1 U9267 ( .B1(n10557), .B2(n8101), .A(n8100), .ZN(P2_U3484) );
  NAND2_X1 U9268 ( .A1(n8102), .A2(n10553), .ZN(n8103) );
  OAI21_X1 U9269 ( .B1(n10553), .B2(n7603), .A(n8103), .ZN(P2_U3531) );
  INV_X1 U9270 ( .A(n8113), .ZN(n9661) );
  OAI21_X1 U9271 ( .B1(n5157), .B2(n9661), .A(n8145), .ZN(n8106) );
  AOI222_X1 U9272 ( .A1(n10397), .A2(n8106), .B1(n8105), .B2(n10391), .C1(
        n9714), .C2(n10393), .ZN(n8164) );
  AOI21_X1 U9273 ( .B1(n8107), .B2(n8162), .A(n10522), .ZN(n8108) );
  AND2_X1 U9274 ( .A1(n8108), .A2(n8152), .ZN(n8161) );
  AOI22_X1 U9275 ( .A1(n10371), .A2(P1_REG2_REG_7__SCAN_IN), .B1(n8109), .B2(
        n10409), .ZN(n8110) );
  OAI21_X1 U9276 ( .B1(n9969), .B2(n8111), .A(n8110), .ZN(n8117) );
  OAI21_X1 U9277 ( .B1(n8114), .B2(n8113), .A(n8112), .ZN(n8115) );
  INV_X1 U9278 ( .A(n8115), .ZN(n8165) );
  NOR2_X1 U9279 ( .A1(n8165), .A2(n9985), .ZN(n8116) );
  AOI211_X1 U9280 ( .C1(n8161), .C2(n9983), .A(n8117), .B(n8116), .ZN(n8118)
         );
  OAI21_X1 U9281 ( .B1(n10419), .B2(n8164), .A(n8118), .ZN(P1_U3284) );
  INV_X1 U9282 ( .A(n8139), .ZN(n10537) );
  OAI21_X1 U9283 ( .B1(n8120), .B2(n4923), .A(n8119), .ZN(n8121) );
  NAND2_X1 U9284 ( .A1(n8121), .A2(n8657), .ZN(n8126) );
  INV_X1 U9285 ( .A(n8122), .ZN(n8124) );
  OAI22_X1 U9286 ( .A1(n8136), .A2(n8678), .B1(n8660), .B2(n8130), .ZN(n8123)
         );
  AOI211_X1 U9287 ( .C1(n8647), .C2(n8691), .A(n8124), .B(n8123), .ZN(n8125)
         );
  OAI211_X1 U9288 ( .C1(n10537), .C2(n8683), .A(n8126), .B(n8125), .ZN(
        P2_U3226) );
  XNOR2_X1 U9289 ( .A(n8128), .B(n8127), .ZN(n8129) );
  OAI222_X1 U9290 ( .A1(n8673), .A2(n8342), .B1(n8675), .B2(n8130), .C1(n8129), 
        .C2(n8461), .ZN(n10539) );
  INV_X1 U9291 ( .A(n10539), .ZN(n8143) );
  XNOR2_X1 U9292 ( .A(n8131), .B(n8132), .ZN(n10542) );
  NAND2_X1 U9293 ( .A1(n8139), .A2(n8134), .ZN(n8135) );
  NAND2_X1 U9294 ( .A1(n8237), .A2(n8135), .ZN(n10538) );
  OAI22_X1 U9295 ( .A1(n8810), .A2(n8137), .B1(n8136), .B2(n10454), .ZN(n8138)
         );
  AOI21_X1 U9296 ( .B1(n8139), .B2(n8943), .A(n8138), .ZN(n8140) );
  OAI21_X1 U9297 ( .B1(n10538), .B2(n8777), .A(n8140), .ZN(n8141) );
  AOI21_X1 U9298 ( .B1(n10542), .B2(n8933), .A(n8141), .ZN(n8142) );
  OAI21_X1 U9299 ( .B1(n8143), .B2(n10466), .A(n8142), .ZN(P2_U3284) );
  OAI21_X1 U9300 ( .B1(n4920), .B2(n9658), .A(n8144), .ZN(n8151) );
  AOI22_X1 U9301 ( .A1(n10393), .A2(n9713), .B1(n9712), .B2(n10391), .ZN(n8150) );
  INV_X1 U9302 ( .A(n8145), .ZN(n8146) );
  OAI21_X1 U9303 ( .B1(n8146), .B2(n9459), .A(n9658), .ZN(n8148) );
  NAND3_X1 U9304 ( .A1(n8148), .A2(n10397), .A3(n8147), .ZN(n8149) );
  OAI211_X1 U9305 ( .C1(n8151), .C2(n10401), .A(n8150), .B(n8149), .ZN(n10483)
         );
  INV_X1 U9306 ( .A(n10483), .ZN(n8160) );
  INV_X1 U9307 ( .A(n8151), .ZN(n10485) );
  INV_X1 U9308 ( .A(n8152), .ZN(n8153) );
  INV_X1 U9309 ( .A(n8155), .ZN(n10481) );
  OAI21_X1 U9310 ( .B1(n8153), .B2(n10481), .A(n8190), .ZN(n10482) );
  AOI22_X1 U9311 ( .A1(n10371), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n8154), .B2(
        n10409), .ZN(n8157) );
  NAND2_X1 U9312 ( .A1(n10367), .A2(n8155), .ZN(n8156) );
  OAI211_X1 U9313 ( .C1(n10482), .C2(n9918), .A(n8157), .B(n8156), .ZN(n8158)
         );
  AOI21_X1 U9314 ( .B1(n10485), .B2(n10415), .A(n8158), .ZN(n8159) );
  OAI21_X1 U9315 ( .B1(n8160), .B2(n10419), .A(n8159), .ZN(P1_U3283) );
  AOI21_X1 U9316 ( .B1(n10502), .B2(n8162), .A(n8161), .ZN(n8163) );
  OAI211_X1 U9317 ( .C1(n10436), .C2(n8165), .A(n8164), .B(n8163), .ZN(n8168)
         );
  NAND2_X1 U9318 ( .A1(n8168), .A2(n10531), .ZN(n8166) );
  OAI21_X1 U9319 ( .B1(n10531), .B2(n8167), .A(n8166), .ZN(P1_U3530) );
  INV_X1 U9320 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n8170) );
  NAND2_X1 U9321 ( .A1(n8168), .A2(n10535), .ZN(n8169) );
  OAI21_X1 U9322 ( .B1(n10535), .B2(n8170), .A(n8169), .ZN(P1_U3475) );
  INV_X1 U9323 ( .A(n8909), .ZN(n8955) );
  INV_X1 U9324 ( .A(n8171), .ZN(n8172) );
  AOI22_X1 U9325 ( .A1(n10466), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n8172), .B2(
        n8945), .ZN(n8173) );
  OAI21_X1 U9326 ( .B1(n8174), .B2(n8930), .A(n8173), .ZN(n8177) );
  NOR2_X1 U9327 ( .A1(n8175), .A2(n8952), .ZN(n8176) );
  AOI211_X1 U9328 ( .C1(n8178), .C2(n8955), .A(n8177), .B(n8176), .ZN(n8179)
         );
  OAI21_X1 U9329 ( .B1(n10466), .B2(n8180), .A(n8179), .ZN(P2_U3285) );
  XNOR2_X1 U9330 ( .A(n8181), .B(n9664), .ZN(n10489) );
  OAI21_X1 U9331 ( .B1(n4922), .B2(n6151), .A(n8182), .ZN(n8186) );
  OAI22_X1 U9332 ( .A1(n8184), .A2(n9977), .B1(n8183), .B2(n9975), .ZN(n8185)
         );
  AOI21_X1 U9333 ( .B1(n8186), .B2(n10397), .A(n8185), .ZN(n8187) );
  OAI21_X1 U9334 ( .B1(n10489), .B2(n10401), .A(n8187), .ZN(n10493) );
  NAND2_X1 U9335 ( .A1(n10493), .A2(n9940), .ZN(n8195) );
  INV_X1 U9336 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n8189) );
  OAI22_X1 U9337 ( .A1(n9940), .A2(n8189), .B1(n8188), .B2(n10376), .ZN(n8193)
         );
  AND2_X1 U9338 ( .A1(n8190), .A2(n10490), .ZN(n8191) );
  OR2_X1 U9339 ( .A1(n8191), .A2(n8277), .ZN(n10492) );
  NOR2_X1 U9340 ( .A1(n10492), .A2(n9918), .ZN(n8192) );
  AOI211_X1 U9341 ( .C1(n10367), .C2(n10490), .A(n8193), .B(n8192), .ZN(n8194)
         );
  OAI211_X1 U9342 ( .C1(n10489), .C2(n9779), .A(n8195), .B(n8194), .ZN(
        P1_U3282) );
  AOI22_X1 U9343 ( .A1(n8197), .A2(n10429), .B1(n10550), .B2(n8196), .ZN(n8198) );
  OAI211_X1 U9344 ( .C1(n8200), .C2(n10510), .A(n8199), .B(n8198), .ZN(n8202)
         );
  NAND2_X1 U9345 ( .A1(n8202), .A2(n10553), .ZN(n8201) );
  OAI21_X1 U9346 ( .B1(n10553), .B2(n6452), .A(n8201), .ZN(P2_U3529) );
  INV_X1 U9347 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n8204) );
  NAND2_X1 U9348 ( .A1(n8202), .A2(n10557), .ZN(n8203) );
  OAI21_X1 U9349 ( .B1(n10557), .B2(n8204), .A(n8203), .ZN(P2_U3478) );
  INV_X1 U9350 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n8205) );
  OAI222_X1 U9351 ( .A1(P1_U3084), .A2(n9685), .B1(n10113), .B2(n8220), .C1(
        n8205), .C2(n10119), .ZN(P1_U3332) );
  OAI21_X1 U9352 ( .B1(n8208), .B2(n8207), .A(n8206), .ZN(n8209) );
  NAND2_X1 U9353 ( .A1(n8209), .A2(n8657), .ZN(n8215) );
  INV_X1 U9354 ( .A(n8210), .ZN(n8213) );
  OAI22_X1 U9355 ( .A1(n8238), .A2(n8678), .B1(n8660), .B2(n8211), .ZN(n8212)
         );
  AOI211_X1 U9356 ( .C1(n8647), .C2(n8409), .A(n8213), .B(n8212), .ZN(n8214)
         );
  OAI211_X1 U9357 ( .C1(n6750), .C2(n8683), .A(n8215), .B(n8214), .ZN(P2_U3236) );
  INV_X1 U9358 ( .A(n8216), .ZN(n8232) );
  INV_X1 U9359 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n8217) );
  OAI222_X1 U9360 ( .A1(P1_U3084), .A2(n8218), .B1(n10113), .B2(n8232), .C1(
        n8217), .C2(n10119), .ZN(P1_U3333) );
  INV_X1 U9361 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n8222) );
  OAI222_X1 U9362 ( .A1(n9300), .A2(n8222), .B1(P2_U3152), .B2(n8221), .C1(
        n8219), .C2(n8220), .ZN(P2_U3337) );
  NAND2_X1 U9363 ( .A1(n8224), .A2(n8223), .ZN(n8226) );
  XNOR2_X1 U9364 ( .A(n8226), .B(n8225), .ZN(n8227) );
  NAND2_X1 U9365 ( .A1(n8227), .A2(n9413), .ZN(n8231) );
  OAI22_X1 U9366 ( .A1(n8276), .A2(n9431), .B1(n9430), .B2(n8387), .ZN(n8228)
         );
  AOI211_X1 U9367 ( .C1(n9434), .C2(n8279), .A(n8229), .B(n8228), .ZN(n8230)
         );
  OAI211_X1 U9368 ( .C1(n8282), .C2(n9409), .A(n8231), .B(n8230), .ZN(P1_U3215) );
  INV_X1 U9369 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n8233) );
  OAI222_X1 U9370 ( .A1(n9300), .A2(n8233), .B1(P2_U3152), .B2(n6710), .C1(
        n8219), .C2(n8232), .ZN(P2_U3338) );
  OAI21_X1 U9371 ( .B1(n4909), .B2(n8235), .A(n8234), .ZN(n9272) );
  INV_X1 U9372 ( .A(n8336), .ZN(n8236) );
  AOI21_X1 U9373 ( .B1(n9267), .B2(n8237), .A(n8236), .ZN(n9268) );
  NOR2_X1 U9374 ( .A1(n6750), .A2(n8930), .ZN(n8241) );
  OAI22_X1 U9375 ( .A1(n8810), .A2(n8239), .B1(n8238), .B2(n10454), .ZN(n8240)
         );
  AOI211_X1 U9376 ( .C1(n9268), .C2(n8926), .A(n8241), .B(n8240), .ZN(n8247)
         );
  XNOR2_X1 U9377 ( .A(n8243), .B(n8242), .ZN(n8245) );
  AOI222_X1 U9378 ( .A1(n8937), .A2(n8245), .B1(n8409), .B2(n8916), .C1(n8244), 
        .C2(n8915), .ZN(n9270) );
  OR2_X1 U9379 ( .A1(n9270), .A2(n10466), .ZN(n8246) );
  OAI211_X1 U9380 ( .C1(n9272), .C2(n8952), .A(n8247), .B(n8246), .ZN(P2_U3283) );
  XOR2_X1 U9381 ( .A(n8249), .B(n8248), .Z(n8254) );
  AOI22_X1 U9382 ( .A1(n9417), .A2(n9711), .B1(n9416), .B2(n9709), .ZN(n8250)
         );
  NAND2_X1 U9383 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3084), .ZN(n10283) );
  OAI211_X1 U9384 ( .C1(n8251), .C2(n9392), .A(n8250), .B(n10283), .ZN(n8252)
         );
  AOI21_X1 U9385 ( .B1(n9446), .B2(n9435), .A(n8252), .ZN(n8253) );
  OAI21_X1 U9386 ( .B1(n8254), .B2(n9438), .A(n8253), .ZN(P1_U3234) );
  NOR2_X1 U9387 ( .A1(n8261), .A2(n8255), .ZN(n8257) );
  NOR2_X1 U9388 ( .A1(n8257), .A2(n8256), .ZN(n8259) );
  XNOR2_X1 U9389 ( .A(n8295), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n8258) );
  NOR2_X1 U9390 ( .A1(n8259), .A2(n8258), .ZN(n8294) );
  AOI211_X1 U9391 ( .C1(n8259), .C2(n8258), .A(n10269), .B(n8294), .ZN(n8272)
         );
  NOR2_X1 U9392 ( .A1(n8261), .A2(n8260), .ZN(n8263) );
  NOR2_X1 U9393 ( .A1(n8263), .A2(n8262), .ZN(n8266) );
  XNOR2_X1 U9394 ( .A(n8295), .B(P1_REG2_REG_16__SCAN_IN), .ZN(n8265) );
  OR2_X1 U9395 ( .A1(n8266), .A2(n8265), .ZN(n8286) );
  INV_X1 U9396 ( .A(n8286), .ZN(n8264) );
  AOI211_X1 U9397 ( .C1(n8266), .C2(n8265), .A(n10298), .B(n8264), .ZN(n8271)
         );
  NAND2_X1 U9398 ( .A1(P1_U3084), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9352) );
  NAND2_X1 U9399 ( .A1(n10313), .A2(P1_ADDR_REG_16__SCAN_IN), .ZN(n8267) );
  OAI211_X1 U9400 ( .C1(n8269), .C2(n8268), .A(n9352), .B(n8267), .ZN(n8270)
         );
  OR3_X1 U9401 ( .A1(n8272), .A2(n8271), .A3(n8270), .ZN(P1_U3257) );
  XNOR2_X1 U9402 ( .A(n8273), .B(n9667), .ZN(n10505) );
  XNOR2_X1 U9403 ( .A(n8274), .B(n9470), .ZN(n8275) );
  OAI222_X1 U9404 ( .A1(n9975), .A2(n8387), .B1(n9977), .B2(n8276), .C1(n8275), 
        .C2(n9972), .ZN(n10499) );
  INV_X1 U9405 ( .A(n8277), .ZN(n8278) );
  AOI211_X1 U9406 ( .C1(n10501), .C2(n8278), .A(n10522), .B(n8328), .ZN(n10500) );
  NAND2_X1 U9407 ( .A1(n10500), .A2(n9983), .ZN(n8281) );
  AOI22_X1 U9408 ( .A1(n10371), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n8279), .B2(
        n10409), .ZN(n8280) );
  OAI211_X1 U9409 ( .C1(n8282), .C2(n9969), .A(n8281), .B(n8280), .ZN(n8283)
         );
  AOI21_X1 U9410 ( .B1(n10499), .B2(n9940), .A(n8283), .ZN(n8284) );
  OAI21_X1 U9411 ( .B1(n9985), .B2(n10505), .A(n8284), .ZN(P1_U3281) );
  NAND2_X1 U9412 ( .A1(n8295), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n8285) );
  NAND2_X1 U9413 ( .A1(n8286), .A2(n8285), .ZN(n8291) );
  INV_X1 U9414 ( .A(n8291), .ZN(n8288) );
  NAND2_X1 U9415 ( .A1(n9727), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n8287) );
  OAI21_X1 U9416 ( .B1(n9727), .B2(P1_REG2_REG_17__SCAN_IN), .A(n8287), .ZN(
        n8289) );
  AOI21_X1 U9417 ( .B1(n8288), .B2(n8289), .A(n10298), .ZN(n8300) );
  INV_X1 U9418 ( .A(n8289), .ZN(n8290) );
  NAND2_X1 U9419 ( .A1(n8291), .A2(n8290), .ZN(n9725) );
  INV_X1 U9420 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n8293) );
  NAND2_X1 U9421 ( .A1(n10312), .A2(n9727), .ZN(n8292) );
  NAND2_X1 U9422 ( .A1(P1_U3084), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9361) );
  OAI211_X1 U9423 ( .C1(n9736), .C2(n8293), .A(n8292), .B(n9361), .ZN(n8299)
         );
  AOI21_X1 U9424 ( .B1(P1_REG1_REG_16__SCAN_IN), .B2(n8295), .A(n8294), .ZN(
        n8297) );
  XNOR2_X1 U9425 ( .A(n9727), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n8296) );
  NOR2_X1 U9426 ( .A1(n8297), .A2(n8296), .ZN(n9720) );
  AOI211_X1 U9427 ( .C1(n8297), .C2(n8296), .A(n10269), .B(n9720), .ZN(n8298)
         );
  AOI211_X1 U9428 ( .C1(n8300), .C2(n9725), .A(n8299), .B(n8298), .ZN(n8301)
         );
  INV_X1 U9429 ( .A(n8301), .ZN(P1_U3258) );
  INV_X1 U9430 ( .A(n9262), .ZN(n8340) );
  OAI21_X1 U9431 ( .B1(n8304), .B2(n8303), .A(n8302), .ZN(n8305) );
  NAND2_X1 U9432 ( .A1(n8305), .A2(n8657), .ZN(n8310) );
  OAI22_X1 U9433 ( .A1(n8337), .A2(n8678), .B1(n8660), .B2(n8342), .ZN(n8306)
         );
  AOI211_X1 U9434 ( .C1(n8647), .C2(n8308), .A(n8307), .B(n8306), .ZN(n8309)
         );
  OAI211_X1 U9435 ( .C1(n8340), .C2(n8683), .A(n8310), .B(n8309), .ZN(P2_U3217) );
  OAI21_X1 U9436 ( .B1(n8312), .B2(P2_REG2_REG_14__SCAN_IN), .A(n8311), .ZN(
        n8707) );
  XOR2_X1 U9437 ( .A(n8708), .B(n8707), .Z(n8313) );
  NAND2_X1 U9438 ( .A1(n8313), .A2(n8415), .ZN(n8709) );
  OAI21_X1 U9439 ( .B1(n8313), .B2(n8415), .A(n8709), .ZN(n8321) );
  INV_X1 U9440 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n8316) );
  INV_X1 U9441 ( .A(n8708), .ZN(n8314) );
  NAND2_X1 U9442 ( .A1(n10364), .A2(n8314), .ZN(n8315) );
  NAND2_X1 U9443 ( .A1(P2_REG3_REG_15__SCAN_IN), .A2(P2_U3152), .ZN(n8375) );
  OAI211_X1 U9444 ( .C1(n8741), .C2(n8316), .A(n8315), .B(n8375), .ZN(n8320)
         );
  XNOR2_X1 U9445 ( .A(n8701), .B(n8708), .ZN(n8318) );
  NOR2_X1 U9446 ( .A1(n8317), .A2(n8318), .ZN(n8702) );
  AOI211_X1 U9447 ( .C1(n8318), .C2(n8317), .A(n8702), .B(n10353), .ZN(n8319)
         );
  AOI211_X1 U9448 ( .C1(n10334), .C2(n8321), .A(n8320), .B(n8319), .ZN(n8322)
         );
  INV_X1 U9449 ( .A(n8322), .ZN(P2_U3260) );
  XNOR2_X1 U9450 ( .A(n8323), .B(n9668), .ZN(n10526) );
  NAND2_X1 U9451 ( .A1(n8324), .A2(n9668), .ZN(n8383) );
  OAI211_X1 U9452 ( .C1(n8324), .C2(n9668), .A(n8383), .B(n10397), .ZN(n8326)
         );
  AOI22_X1 U9453 ( .A1(n10393), .A2(n9711), .B1(n9709), .B2(n10391), .ZN(n8325) );
  NAND2_X1 U9454 ( .A1(n8326), .A2(n8325), .ZN(n8327) );
  AOI21_X1 U9455 ( .B1(n10526), .B2(n6266), .A(n8327), .ZN(n10528) );
  NOR2_X1 U9456 ( .A1(n8328), .A2(n10521), .ZN(n8329) );
  OR2_X1 U9457 ( .A1(n8388), .A2(n8329), .ZN(n10523) );
  AOI22_X1 U9458 ( .A1(n10419), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n8330), .B2(
        n10409), .ZN(n8332) );
  NAND2_X1 U9459 ( .A1(n9446), .A2(n10367), .ZN(n8331) );
  OAI211_X1 U9460 ( .C1(n10523), .C2(n9918), .A(n8332), .B(n8331), .ZN(n8333)
         );
  AOI21_X1 U9461 ( .B1(n10526), .B2(n10415), .A(n8333), .ZN(n8334) );
  OAI21_X1 U9462 ( .B1(n10528), .B2(n10371), .A(n8334), .ZN(P1_U3280) );
  XNOR2_X1 U9463 ( .A(n8335), .B(n5290), .ZN(n9266) );
  AOI21_X1 U9464 ( .B1(n9262), .B2(n8336), .A(n8411), .ZN(n9263) );
  INV_X1 U9465 ( .A(n8337), .ZN(n8338) );
  AOI22_X1 U9466 ( .A1(n10466), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n8338), .B2(
        n8945), .ZN(n8339) );
  OAI21_X1 U9467 ( .B1(n8340), .B2(n8930), .A(n8339), .ZN(n8347) );
  AOI21_X1 U9468 ( .B1(n5290), .B2(n8341), .A(n8461), .ZN(n8345) );
  OAI22_X1 U9469 ( .A1(n8427), .A2(n8673), .B1(n8342), .B2(n8675), .ZN(n8343)
         );
  AOI21_X1 U9470 ( .B1(n8345), .B2(n8344), .A(n8343), .ZN(n9265) );
  NOR2_X1 U9471 ( .A1(n9265), .A2(n10466), .ZN(n8346) );
  AOI211_X1 U9472 ( .C1(n9263), .C2(n8926), .A(n8347), .B(n8346), .ZN(n8348)
         );
  OAI21_X1 U9473 ( .B1(n9266), .B2(n8952), .A(n8348), .ZN(P2_U3282) );
  INV_X1 U9474 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n8351) );
  INV_X1 U9475 ( .A(n8349), .ZN(n8516) );
  OAI222_X1 U9476 ( .A1(n9300), .A2(n8351), .B1(n8219), .B2(n8516), .C1(n8350), 
        .C2(P2_U3152), .ZN(P2_U3336) );
  XOR2_X1 U9477 ( .A(n8353), .B(n8352), .Z(n8354) );
  XNOR2_X1 U9478 ( .A(n8355), .B(n8354), .ZN(n8356) );
  NAND2_X1 U9479 ( .A1(n8356), .A2(n9413), .ZN(n8360) );
  OAI22_X1 U9480 ( .A1(n8387), .A2(n9431), .B1(n9430), .B2(n9978), .ZN(n8357)
         );
  AOI211_X1 U9481 ( .C1(n9434), .C2(n8390), .A(n8358), .B(n8357), .ZN(n8359)
         );
  OAI211_X1 U9482 ( .C1(n8393), .C2(n9409), .A(n8360), .B(n8359), .ZN(P1_U3222) );
  INV_X1 U9483 ( .A(n8361), .ZN(n8363) );
  NOR2_X1 U9484 ( .A1(n8363), .A2(n8362), .ZN(n8364) );
  XNOR2_X1 U9485 ( .A(n8365), .B(n8364), .ZN(n8370) );
  INV_X1 U9486 ( .A(n8479), .ZN(n8367) );
  AOI22_X1 U9487 ( .A1(n9416), .A2(n9707), .B1(n9417), .B2(n9709), .ZN(n8366)
         );
  NAND2_X1 U9488 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3084), .ZN(n10296) );
  OAI211_X1 U9489 ( .C1(n8367), .C2(n9392), .A(n8366), .B(n10296), .ZN(n8368)
         );
  AOI21_X1 U9490 ( .B1(n6157), .B2(n9435), .A(n8368), .ZN(n8369) );
  OAI21_X1 U9491 ( .B1(n8370), .B2(n9438), .A(n8369), .ZN(P1_U3232) );
  OAI21_X1 U9492 ( .B1(n8373), .B2(n8372), .A(n8371), .ZN(n8374) );
  NAND2_X1 U9493 ( .A1(n8374), .A2(n8657), .ZN(n8380) );
  INV_X1 U9494 ( .A(n8375), .ZN(n8378) );
  OAI22_X1 U9495 ( .A1(n8414), .A2(n8678), .B1(n8660), .B2(n8376), .ZN(n8377)
         );
  AOI211_X1 U9496 ( .C1(n8647), .C2(n8690), .A(n8378), .B(n8377), .ZN(n8379)
         );
  OAI211_X1 U9497 ( .C1(n7099), .C2(n8683), .A(n8380), .B(n8379), .ZN(P2_U3243) );
  NAND2_X1 U9498 ( .A1(n8381), .A2(n9474), .ZN(n8467) );
  XNOR2_X1 U9499 ( .A(n8467), .B(n9670), .ZN(n10082) );
  NAND2_X1 U9500 ( .A1(n8383), .A2(n9550), .ZN(n8385) );
  AND2_X1 U9501 ( .A1(n8383), .A2(n8382), .ZN(n8384) );
  AOI21_X1 U9502 ( .B1(n9670), .B2(n8385), .A(n8384), .ZN(n8386) );
  OAI222_X1 U9503 ( .A1(n9975), .A2(n9978), .B1(n9977), .B2(n8387), .C1(n9972), 
        .C2(n8386), .ZN(n10078) );
  INV_X1 U9504 ( .A(n8388), .ZN(n8389) );
  AOI211_X1 U9505 ( .C1(n10080), .C2(n8389), .A(n10522), .B(n4990), .ZN(n10079) );
  NAND2_X1 U9506 ( .A1(n10079), .A2(n9983), .ZN(n8392) );
  AOI22_X1 U9507 ( .A1(n10371), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n8390), .B2(
        n10409), .ZN(n8391) );
  OAI211_X1 U9508 ( .C1(n8393), .C2(n9969), .A(n8392), .B(n8391), .ZN(n8394)
         );
  AOI21_X1 U9509 ( .B1(n10078), .B2(n9940), .A(n8394), .ZN(n8395) );
  OAI21_X1 U9510 ( .B1(n9985), .B2(n10082), .A(n8395), .ZN(P1_U3279) );
  INV_X1 U9511 ( .A(n8396), .ZN(n8401) );
  NOR2_X1 U9512 ( .A1(n8397), .A2(P1_U3084), .ZN(n9697) );
  AOI21_X1 U9513 ( .B1(P2_DATAO_REG_23__SCAN_IN), .B2(n10107), .A(n9697), .ZN(
        n8398) );
  OAI21_X1 U9514 ( .B1(n8401), .B2(n10113), .A(n8398), .ZN(P1_U3330) );
  NAND2_X1 U9515 ( .A1(n9297), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n8399) );
  OAI211_X1 U9516 ( .C1(n8401), .C2(n8219), .A(n8400), .B(n8399), .ZN(P2_U3335) );
  INV_X1 U9517 ( .A(n8402), .ZN(n8406) );
  OAI222_X1 U9518 ( .A1(P1_U3084), .A2(n8404), .B1(n10119), .B2(n8403), .C1(
        n8406), .C2(n10113), .ZN(P1_U3329) );
  INV_X1 U9519 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n8405) );
  OAI222_X1 U9520 ( .A1(P2_U3152), .A2(n8407), .B1(n8219), .B2(n8406), .C1(
        n8405), .C2(n9300), .ZN(P2_U3334) );
  XNOR2_X1 U9521 ( .A(n8419), .B(n8408), .ZN(n8410) );
  AOI222_X1 U9522 ( .A1(n8937), .A2(n8410), .B1(n8690), .B2(n8916), .C1(n8409), 
        .C2(n8915), .ZN(n9260) );
  INV_X1 U9523 ( .A(n8411), .ZN(n8413) );
  INV_X1 U9524 ( .A(n8939), .ZN(n8412) );
  AOI21_X1 U9525 ( .B1(n9257), .B2(n8413), .A(n8412), .ZN(n9258) );
  NOR2_X1 U9526 ( .A1(n7099), .A2(n8930), .ZN(n8417) );
  OAI22_X1 U9527 ( .A1(n8810), .A2(n8415), .B1(n8414), .B2(n10454), .ZN(n8416)
         );
  AOI211_X1 U9528 ( .C1(n9258), .C2(n8926), .A(n8417), .B(n8416), .ZN(n8422)
         );
  OAI21_X1 U9529 ( .B1(n8420), .B2(n8419), .A(n8418), .ZN(n9256) );
  NAND2_X1 U9530 ( .A1(n9256), .A2(n8933), .ZN(n8421) );
  OAI211_X1 U9531 ( .C1(n9260), .C2(n10466), .A(n8422), .B(n8421), .ZN(
        P2_U3281) );
  INV_X1 U9532 ( .A(n7105), .ZN(n8433) );
  OAI21_X1 U9533 ( .B1(n8425), .B2(n8424), .A(n8423), .ZN(n8426) );
  NAND2_X1 U9534 ( .A1(n8426), .A2(n8657), .ZN(n8432) );
  OAI22_X1 U9535 ( .A1(n8428), .A2(n8673), .B1(n8427), .B2(n8675), .ZN(n8936)
         );
  NOR2_X1 U9536 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6551), .ZN(n8704) );
  INV_X1 U9537 ( .A(n8944), .ZN(n8429) );
  NOR2_X1 U9538 ( .A1(n8678), .A2(n8429), .ZN(n8430) );
  AOI211_X1 U9539 ( .C1(n8680), .C2(n8936), .A(n8704), .B(n8430), .ZN(n8431)
         );
  OAI211_X1 U9540 ( .C1(n8433), .C2(n8683), .A(n8432), .B(n8431), .ZN(P2_U3228) );
  INV_X1 U9541 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n8436) );
  INV_X1 U9542 ( .A(n8434), .ZN(n8437) );
  OAI222_X1 U9543 ( .A1(n9300), .A2(n8436), .B1(n8219), .B2(n8437), .C1(
        P2_U3152), .C2(n8435), .ZN(P2_U3333) );
  INV_X1 U9544 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n8438) );
  OAI222_X1 U9545 ( .A1(n10119), .A2(n8438), .B1(n10113), .B2(n8437), .C1(
        P1_U3084), .C2(n6094), .ZN(P1_U3328) );
  INV_X1 U9546 ( .A(n8439), .ZN(n8441) );
  NAND2_X1 U9547 ( .A1(n8441), .A2(n8440), .ZN(n8442) );
  XNOR2_X1 U9548 ( .A(n8443), .B(n8442), .ZN(n8449) );
  NOR2_X1 U9549 ( .A1(n8678), .A2(n8454), .ZN(n8447) );
  INV_X1 U9550 ( .A(n8680), .ZN(n8445) );
  AOI22_X1 U9551 ( .A1(n8689), .A2(n8916), .B1(n8915), .B2(n8690), .ZN(n8460)
         );
  OAI22_X1 U9552 ( .A1(n8445), .A2(n8460), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8444), .ZN(n8446) );
  AOI211_X1 U9553 ( .C1(n9249), .C2(n8641), .A(n8447), .B(n8446), .ZN(n8448)
         );
  OAI21_X1 U9554 ( .B1(n8449), .B2(n8669), .A(n8448), .ZN(P2_U3230) );
  XNOR2_X1 U9555 ( .A(n8450), .B(n8459), .ZN(n9251) );
  INV_X1 U9556 ( .A(n8942), .ZN(n8452) );
  INV_X1 U9557 ( .A(n8923), .ZN(n8451) );
  AOI211_X1 U9558 ( .C1(n9249), .C2(n8452), .A(n10545), .B(n8451), .ZN(n9248)
         );
  NOR2_X1 U9559 ( .A1(n8453), .A2(n8930), .ZN(n8457) );
  INV_X1 U9560 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8455) );
  OAI22_X1 U9561 ( .A1(n8810), .A2(n8455), .B1(n8454), .B2(n10454), .ZN(n8456)
         );
  AOI211_X1 U9562 ( .C1(n9248), .C2(n8955), .A(n8457), .B(n8456), .ZN(n8464)
         );
  XNOR2_X1 U9563 ( .A(n8459), .B(n8458), .ZN(n8462) );
  OAI21_X1 U9564 ( .B1(n8462), .B2(n8461), .A(n8460), .ZN(n9247) );
  NAND2_X1 U9565 ( .A1(n9247), .A2(n8810), .ZN(n8463) );
  OAI211_X1 U9566 ( .C1(n9251), .C2(n8952), .A(n8464), .B(n8463), .ZN(P2_U3279) );
  INV_X1 U9567 ( .A(n8465), .ZN(n8497) );
  AOI22_X1 U9568 ( .A1(n6096), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n10107), .ZN(n8466) );
  OAI21_X1 U9569 ( .B1(n8497), .B2(n10113), .A(n8466), .ZN(P1_U3327) );
  NAND2_X1 U9570 ( .A1(n8467), .A2(n9670), .ZN(n8469) );
  NAND2_X1 U9571 ( .A1(n8469), .A2(n8468), .ZN(n8470) );
  NAND2_X1 U9572 ( .A1(n8470), .A2(n8472), .ZN(n8471) );
  NAND2_X1 U9573 ( .A1(n9963), .A2(n8471), .ZN(n10072) );
  INV_X1 U9574 ( .A(n10072), .ZN(n8485) );
  XNOR2_X1 U9575 ( .A(n8473), .B(n8472), .ZN(n8476) );
  NAND2_X1 U9576 ( .A1(n10072), .A2(n6266), .ZN(n8475) );
  AOI22_X1 U9577 ( .A1(n10391), .A2(n9707), .B1(n9709), .B2(n10393), .ZN(n8474) );
  OAI211_X1 U9578 ( .C1(n9972), .C2(n8476), .A(n8475), .B(n8474), .ZN(n10077)
         );
  NAND2_X1 U9579 ( .A1(n10077), .A2(n9940), .ZN(n8484) );
  NAND2_X1 U9580 ( .A1(n8477), .A2(n6157), .ZN(n8478) );
  INV_X1 U9581 ( .A(n6157), .ZN(n8481) );
  AOI22_X1 U9582 ( .A1(n10371), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n8479), .B2(
        n10409), .ZN(n8480) );
  OAI21_X1 U9583 ( .B1(n8481), .B2(n9969), .A(n8480), .ZN(n8482) );
  AOI21_X1 U9584 ( .B1(n10073), .B2(n10368), .A(n8482), .ZN(n8483) );
  OAI211_X1 U9585 ( .C1(n8485), .C2(n9779), .A(n8484), .B(n8483), .ZN(P1_U3278) );
  INV_X1 U9586 ( .A(n8486), .ZN(n8487) );
  NOR2_X1 U9587 ( .A1(n8488), .A2(n8487), .ZN(n8489) );
  XNOR2_X1 U9588 ( .A(n8490), .B(n8489), .ZN(n8495) );
  AOI22_X1 U9589 ( .A1(n8927), .A2(n8665), .B1(n8648), .B2(n8914), .ZN(n8491)
         );
  NAND2_X1 U9590 ( .A1(P2_U3152), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8739) );
  OAI211_X1 U9591 ( .C1(n8492), .C2(n8662), .A(n8491), .B(n8739), .ZN(n8493)
         );
  AOI21_X1 U9592 ( .B1(n9242), .B2(n8641), .A(n8493), .ZN(n8494) );
  OAI21_X1 U9593 ( .B1(n8495), .B2(n8669), .A(n8494), .ZN(P2_U3240) );
  INV_X1 U9594 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n8496) );
  OAI222_X1 U9595 ( .A1(P2_U3152), .A2(n8498), .B1(n8219), .B2(n8497), .C1(
        n8496), .C2(n9300), .ZN(P2_U3332) );
  INV_X1 U9596 ( .A(n8499), .ZN(n8513) );
  AOI21_X1 U9597 ( .B1(n10107), .B2(P2_DATAO_REG_27__SCAN_IN), .A(n8500), .ZN(
        n8501) );
  OAI21_X1 U9598 ( .B1(n8513), .B2(n10113), .A(n8501), .ZN(P1_U3326) );
  XNOR2_X1 U9599 ( .A(n8503), .B(n8502), .ZN(n8504) );
  XNOR2_X1 U9600 ( .A(n8505), .B(n8504), .ZN(n8511) );
  OR2_X1 U9601 ( .A1(n8687), .A2(n8673), .ZN(n8507) );
  NAND2_X1 U9602 ( .A1(n8689), .A2(n8915), .ZN(n8506) );
  NAND2_X1 U9603 ( .A1(n8507), .A2(n8506), .ZN(n8901) );
  NOR2_X1 U9604 ( .A1(n9118), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8764) );
  AOI21_X1 U9605 ( .B1(n8680), .B2(n8901), .A(n8764), .ZN(n8508) );
  OAI21_X1 U9606 ( .B1(n8678), .B2(n8906), .A(n8508), .ZN(n8509) );
  AOI21_X1 U9607 ( .B1(n9232), .B2(n8641), .A(n8509), .ZN(n8510) );
  OAI21_X1 U9608 ( .B1(n8511), .B2(n8669), .A(n8510), .ZN(P2_U3221) );
  INV_X1 U9609 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n8514) );
  OAI222_X1 U9610 ( .A1(n9300), .A2(n8514), .B1(n8219), .B2(n8513), .C1(n8512), 
        .C2(P2_U3152), .ZN(P2_U3331) );
  INV_X1 U9611 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n8517) );
  OAI222_X1 U9612 ( .A1(n10119), .A2(n8517), .B1(n10113), .B2(n8516), .C1(
        P1_U3084), .C2(n8515), .ZN(P1_U3331) );
  INV_X1 U9613 ( .A(n8518), .ZN(n10112) );
  OAI222_X1 U9614 ( .A1(P2_U3152), .A2(n8519), .B1(n8219), .B2(n10112), .C1(
        n9300), .C2(n6177), .ZN(P2_U3329) );
  NOR2_X1 U9615 ( .A1(n8617), .A2(n8542), .ZN(n8521) );
  XNOR2_X1 U9616 ( .A(n8999), .B(n8543), .ZN(n8522) );
  XOR2_X1 U9617 ( .A(n8521), .B(n8522), .Z(n8655) );
  NAND2_X1 U9618 ( .A1(n8654), .A2(n8523), .ZN(n8526) );
  XNOR2_X1 U9619 ( .A(n8993), .B(n8543), .ZN(n8524) );
  NOR2_X1 U9620 ( .A1(n8661), .A2(n8542), .ZN(n8615) );
  INV_X1 U9621 ( .A(n8524), .ZN(n8525) );
  OR2_X1 U9622 ( .A1(n8526), .A2(n8525), .ZN(n8527) );
  XNOR2_X1 U9623 ( .A(n8840), .B(n8543), .ZN(n8529) );
  NOR2_X1 U9624 ( .A1(n8629), .A2(n8542), .ZN(n8637) );
  XNOR2_X1 U9625 ( .A(n8982), .B(n8543), .ZN(n8531) );
  NOR2_X1 U9626 ( .A1(n8686), .A2(n8542), .ZN(n8530) );
  XNOR2_X1 U9627 ( .A(n8531), .B(n8530), .ZN(n8626) );
  XNOR2_X1 U9628 ( .A(n8801), .B(n8543), .ZN(n8534) );
  NOR2_X1 U9629 ( .A1(n8627), .A2(n8542), .ZN(n8533) );
  NAND2_X1 U9630 ( .A1(n8534), .A2(n8533), .ZN(n8536) );
  OAI21_X1 U9631 ( .B1(n8534), .B2(n8533), .A(n8536), .ZN(n8670) );
  INV_X1 U9632 ( .A(n8670), .ZN(n8535) );
  NAND2_X1 U9633 ( .A1(n8671), .A2(n8536), .ZN(n8607) );
  XNOR2_X1 U9634 ( .A(n8970), .B(n8537), .ZN(n8539) );
  OR2_X1 U9635 ( .A1(n8674), .A2(n8542), .ZN(n8538) );
  NOR2_X1 U9636 ( .A1(n8539), .A2(n8538), .ZN(n8540) );
  AOI21_X1 U9637 ( .B1(n8539), .B2(n8538), .A(n8540), .ZN(n8606) );
  NAND2_X1 U9638 ( .A1(n8607), .A2(n8606), .ZN(n8605) );
  INV_X1 U9639 ( .A(n8540), .ZN(n8541) );
  NAND2_X1 U9640 ( .A1(n8605), .A2(n8541), .ZN(n8547) );
  NOR2_X1 U9641 ( .A1(n8609), .A2(n8542), .ZN(n8544) );
  MUX2_X1 U9642 ( .A(n8544), .B(n8609), .S(n8543), .Z(n8545) );
  XNOR2_X1 U9643 ( .A(n8965), .B(n8545), .ZN(n8546) );
  XNOR2_X1 U9644 ( .A(n8547), .B(n8546), .ZN(n8554) );
  OAI22_X1 U9645 ( .A1(n8549), .A2(n8662), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8548), .ZN(n8552) );
  OAI22_X1 U9646 ( .A1(n8674), .A2(n8660), .B1(n8678), .B2(n8550), .ZN(n8551)
         );
  AOI211_X1 U9647 ( .C1(n8965), .C2(n8641), .A(n8552), .B(n8551), .ZN(n8553)
         );
  OAI21_X1 U9648 ( .B1(n8554), .B2(n8669), .A(n8553), .ZN(P2_U3222) );
  NAND2_X1 U9649 ( .A1(n9293), .A2(n8558), .ZN(n8557) );
  INV_X1 U9650 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n8555) );
  OR2_X1 U9651 ( .A1(n5528), .A2(n8555), .ZN(n8556) );
  NAND2_X1 U9652 ( .A1(n8602), .A2(n8558), .ZN(n8560) );
  OR2_X1 U9653 ( .A1(n5528), .A2(n8603), .ZN(n8559) );
  NAND2_X1 U9654 ( .A1(n9993), .A2(n9741), .ZN(n9989) );
  NAND2_X1 U9655 ( .A1(n4851), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n8564) );
  NAND2_X1 U9656 ( .A1(n4854), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n8563) );
  NAND2_X1 U9657 ( .A1(n8561), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n8562) );
  NAND3_X1 U9658 ( .A1(n8564), .A2(n8563), .A3(n8562), .ZN(n9702) );
  INV_X1 U9659 ( .A(n8565), .ZN(n8566) );
  NAND2_X1 U9660 ( .A1(n9702), .A2(n8566), .ZN(n9991) );
  NOR2_X1 U9661 ( .A1(n10371), .A2(n9991), .ZN(n9744) );
  INV_X1 U9662 ( .A(n9986), .ZN(n9440) );
  NOR2_X1 U9663 ( .A1(n9440), .A2(n9969), .ZN(n8567) );
  AOI211_X1 U9664 ( .C1(n10419), .C2(P1_REG2_REG_31__SCAN_IN), .A(n9744), .B(
        n8567), .ZN(n8568) );
  OAI21_X1 U9665 ( .B1(n9988), .B2(n9918), .A(n8568), .ZN(P1_U3261) );
  INV_X1 U9666 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n8570) );
  INV_X1 U9667 ( .A(n10115), .ZN(n8569) );
  OAI222_X1 U9668 ( .A1(n9300), .A2(n8570), .B1(n8219), .B2(n8569), .C1(n6741), 
        .C2(P2_U3152), .ZN(P2_U3330) );
  OAI21_X1 U9669 ( .B1(n8572), .B2(n8579), .A(n8571), .ZN(n10424) );
  INV_X1 U9670 ( .A(n10424), .ZN(n8586) );
  INV_X1 U9671 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n8573) );
  OAI22_X1 U9672 ( .A1(n9940), .A2(n8574), .B1(n8573), .B2(n10376), .ZN(n8578)
         );
  OR2_X1 U9673 ( .A1(n10420), .A2(n10388), .ZN(n8575) );
  NAND2_X1 U9674 ( .A1(n8576), .A2(n8575), .ZN(n10421) );
  NOR2_X1 U9675 ( .A1(n9918), .A2(n10421), .ZN(n8577) );
  AOI211_X1 U9676 ( .C1(n10367), .C2(n8590), .A(n8578), .B(n8577), .ZN(n8585)
         );
  XNOR2_X1 U9677 ( .A(n9588), .B(n8579), .ZN(n8583) );
  OAI22_X1 U9678 ( .A1(n9592), .A2(n9977), .B1(n8580), .B2(n9975), .ZN(n8581)
         );
  AOI21_X1 U9679 ( .B1(n10424), .B2(n6266), .A(n8581), .ZN(n8582) );
  OAI21_X1 U9680 ( .B1(n9972), .B2(n8583), .A(n8582), .ZN(n10422) );
  NAND2_X1 U9681 ( .A1(n10422), .A2(n9940), .ZN(n8584) );
  OAI211_X1 U9682 ( .C1(n8586), .C2(n9779), .A(n8585), .B(n8584), .ZN(P1_U3289) );
  XOR2_X1 U9683 ( .A(n8587), .B(n8588), .Z(n8593) );
  AOI22_X1 U9684 ( .A1(n9435), .A2(n8590), .B1(P1_REG3_REG_2__SCAN_IN), .B2(
        n8589), .ZN(n8592) );
  AOI22_X1 U9685 ( .A1(n9417), .A2(n9718), .B1(n9416), .B2(n9717), .ZN(n8591)
         );
  OAI211_X1 U9686 ( .C1(n8593), .C2(n9438), .A(n8592), .B(n8591), .ZN(P1_U3235) );
  AOI22_X1 U9687 ( .A1(n10371), .A2(P1_REG2_REG_28__SCAN_IN), .B1(n8594), .B2(
        n10409), .ZN(n8595) );
  OAI21_X1 U9688 ( .B1(n4982), .B2(n9969), .A(n8595), .ZN(n8598) );
  NOR2_X1 U9689 ( .A1(n8596), .A2(n9779), .ZN(n8597) );
  OAI21_X1 U9690 ( .B1(n8601), .B2(n10371), .A(n8600), .ZN(P1_U3263) );
  INV_X1 U9691 ( .A(n8602), .ZN(n9301) );
  OAI222_X1 U9692 ( .A1(P1_U3084), .A2(n8604), .B1(n10113), .B2(n9301), .C1(
        n8603), .C2(n10119), .ZN(P1_U3323) );
  OAI211_X1 U9693 ( .C1(n8607), .C2(n8606), .A(n8605), .B(n8657), .ZN(n8613)
         );
  NOR2_X1 U9694 ( .A1(n8627), .A2(n8660), .ZN(n8611) );
  OAI22_X1 U9695 ( .A1(n8609), .A2(n8662), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8608), .ZN(n8610) );
  AOI211_X1 U9696 ( .C1(n8665), .C2(n8787), .A(n8611), .B(n8610), .ZN(n8612)
         );
  OAI211_X1 U9697 ( .C1(n8790), .C2(n8683), .A(n8613), .B(n8612), .ZN(P2_U3216) );
  OAI211_X1 U9698 ( .C1(n8616), .C2(n8615), .A(n8614), .B(n8657), .ZN(n8621)
         );
  OAI22_X1 U9699 ( .A1(n8662), .A2(n8629), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9184), .ZN(n8619) );
  OAI22_X1 U9700 ( .A1(n8678), .A2(n8850), .B1(n8660), .B2(n8617), .ZN(n8618)
         );
  NAND2_X1 U9701 ( .A1(n8621), .A2(n8620), .ZN(P2_U3218) );
  INV_X1 U9703 ( .A(n8623), .ZN(n8625) );
  AOI21_X1 U9704 ( .B1(n8626), .B2(n8622), .A(n8625), .ZN(n8633) );
  OAI22_X1 U9705 ( .A1(n8627), .A2(n8662), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9197), .ZN(n8631) );
  INV_X1 U9706 ( .A(n8816), .ZN(n8628) );
  OAI22_X1 U9707 ( .A1(n8629), .A2(n8660), .B1(n8678), .B2(n8628), .ZN(n8630)
         );
  AOI211_X1 U9708 ( .C1(n8982), .C2(n8641), .A(n8631), .B(n8630), .ZN(n8632)
         );
  OAI21_X1 U9709 ( .B1(n8633), .B2(n8669), .A(n8632), .ZN(P2_U3227) );
  OAI211_X1 U9710 ( .C1(n8635), .C2(n8637), .A(n8636), .B(n8657), .ZN(n8643)
         );
  OAI22_X1 U9711 ( .A1(n8686), .A2(n8662), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8638), .ZN(n8640) );
  OAI22_X1 U9712 ( .A1(n8678), .A2(n8836), .B1(n8660), .B2(n8661), .ZN(n8639)
         );
  AOI211_X1 U9713 ( .C1(n8987), .C2(n8641), .A(n8640), .B(n8639), .ZN(n8642)
         );
  NAND2_X1 U9714 ( .A1(n8643), .A2(n8642), .ZN(P2_U3231) );
  AOI211_X1 U9715 ( .C1(n8646), .C2(n8645), .A(n8669), .B(n8644), .ZN(n8653)
         );
  AOI22_X1 U9716 ( .A1(n8647), .A2(n8887), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3152), .ZN(n8650) );
  AOI22_X1 U9717 ( .A1(n8892), .A2(n8665), .B1(n8648), .B2(n8917), .ZN(n8649)
         );
  OAI211_X1 U9718 ( .C1(n8651), .C2(n8683), .A(n8650), .B(n8649), .ZN(n8652)
         );
  OR2_X1 U9719 ( .A1(n8653), .A2(n8652), .ZN(P2_U3235) );
  INV_X1 U9720 ( .A(n8999), .ZN(n8861) );
  OAI21_X1 U9721 ( .B1(n8656), .B2(n8655), .A(n8654), .ZN(n8658) );
  NAND2_X1 U9722 ( .A1(n8658), .A2(n8657), .ZN(n8667) );
  NOR2_X1 U9723 ( .A1(n8660), .A2(n8659), .ZN(n8664) );
  OAI22_X1 U9724 ( .A1(n8662), .A2(n8661), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9209), .ZN(n8663) );
  AOI211_X1 U9725 ( .C1(n8665), .C2(n8859), .A(n8664), .B(n8663), .ZN(n8666)
         );
  OAI211_X1 U9726 ( .C1(n8861), .C2(n8683), .A(n8667), .B(n8666), .ZN(P2_U3237) );
  INV_X1 U9727 ( .A(n8801), .ZN(n8977) );
  AOI21_X1 U9728 ( .B1(n8668), .B2(n8670), .A(n8669), .ZN(n8672) );
  NAND2_X1 U9729 ( .A1(n8672), .A2(n8671), .ZN(n8682) );
  OR2_X1 U9730 ( .A1(n8674), .A2(n8673), .ZN(n8677) );
  OR2_X1 U9731 ( .A1(n8686), .A2(n8675), .ZN(n8676) );
  NAND2_X1 U9732 ( .A1(n8677), .A2(n8676), .ZN(n8805) );
  OAI22_X1 U9733 ( .A1(n8798), .A2(n8678), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9114), .ZN(n8679) );
  AOI21_X1 U9734 ( .B1(n8805), .B2(n8680), .A(n8679), .ZN(n8681) );
  OAI211_X1 U9735 ( .C1(n8977), .C2(n8683), .A(n8682), .B(n8681), .ZN(P2_U3242) );
  MUX2_X1 U9736 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n8684), .S(P2_U3966), .Z(
        P2_U3583) );
  MUX2_X1 U9737 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8685), .S(P2_U3966), .Z(
        P2_U3579) );
  MUX2_X1 U9738 ( .A(n8821), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8688), .Z(
        P2_U3578) );
  INV_X1 U9739 ( .A(n8686), .ZN(n8829) );
  MUX2_X1 U9740 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8829), .S(P2_U3966), .Z(
        P2_U3577) );
  MUX2_X1 U9741 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8871), .S(P2_U3966), .Z(
        P2_U3574) );
  MUX2_X1 U9742 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8887), .S(P2_U3966), .Z(
        P2_U3573) );
  INV_X1 U9743 ( .A(n8687), .ZN(n8870) );
  MUX2_X1 U9744 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8870), .S(P2_U3966), .Z(
        P2_U3572) );
  MUX2_X1 U9745 ( .A(n8917), .B(P2_DATAO_REG_19__SCAN_IN), .S(n8688), .Z(
        P2_U3571) );
  MUX2_X1 U9746 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n8689), .S(P2_U3966), .Z(
        P2_U3570) );
  MUX2_X1 U9747 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8914), .S(P2_U3966), .Z(
        P2_U3569) );
  MUX2_X1 U9748 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8690), .S(P2_U3966), .Z(
        P2_U3568) );
  MUX2_X1 U9749 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n8691), .S(P2_U3966), .Z(
        P2_U3565) );
  MUX2_X1 U9750 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n8692), .S(P2_U3966), .Z(
        P2_U3562) );
  MUX2_X1 U9751 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n8693), .S(P2_U3966), .Z(
        P2_U3561) );
  MUX2_X1 U9752 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n8694), .S(P2_U3966), .Z(
        P2_U3560) );
  MUX2_X1 U9753 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n8696), .S(P2_U3966), .Z(
        P2_U3559) );
  MUX2_X1 U9754 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(n8697), .S(P2_U3966), .Z(
        P2_U3557) );
  MUX2_X1 U9755 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n8698), .S(P2_U3966), .Z(
        P2_U3556) );
  MUX2_X1 U9756 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n8699), .S(P2_U3966), .Z(
        P2_U3553) );
  MUX2_X1 U9757 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n8700), .S(P2_U3966), .Z(
        P2_U3552) );
  NOR2_X1 U9758 ( .A1(n8701), .A2(n8708), .ZN(n8703) );
  XNOR2_X1 U9759 ( .A(n8723), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n8718) );
  XNOR2_X1 U9760 ( .A(n8717), .B(n8718), .ZN(n8716) );
  INV_X1 U9761 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n8706) );
  INV_X1 U9762 ( .A(n8704), .ZN(n8705) );
  OAI21_X1 U9763 ( .B1(n8741), .B2(n8706), .A(n8705), .ZN(n8714) );
  NAND2_X1 U9764 ( .A1(n8708), .A2(n8707), .ZN(n8710) );
  NAND2_X1 U9765 ( .A1(n8710), .A2(n8709), .ZN(n8712) );
  XNOR2_X1 U9766 ( .A(n8723), .B(P2_REG2_REG_16__SCAN_IN), .ZN(n8711) );
  NOR2_X1 U9767 ( .A1(n8712), .A2(n8711), .ZN(n8722) );
  AOI211_X1 U9768 ( .C1(n8712), .C2(n8711), .A(n10357), .B(n8722), .ZN(n8713)
         );
  AOI211_X1 U9769 ( .C1(n10364), .C2(n8723), .A(n8714), .B(n8713), .ZN(n8715)
         );
  OAI21_X1 U9770 ( .B1(n8716), .B2(n10353), .A(n8715), .ZN(P2_U3261) );
  XNOR2_X1 U9771 ( .A(n8738), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n8721) );
  INV_X1 U9772 ( .A(n8717), .ZN(n8719) );
  OAI22_X1 U9773 ( .A1(n8719), .A2(n8718), .B1(n8723), .B2(
        P2_REG1_REG_16__SCAN_IN), .ZN(n8720) );
  NOR2_X1 U9774 ( .A1(n8720), .A2(n8721), .ZN(n8737) );
  AOI211_X1 U9775 ( .C1(n8721), .C2(n8720), .A(n10353), .B(n8737), .ZN(n8732)
         );
  NAND2_X1 U9776 ( .A1(n8738), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n8724) );
  OAI21_X1 U9777 ( .B1(n8738), .B2(P2_REG2_REG_17__SCAN_IN), .A(n8724), .ZN(
        n8725) );
  NOR2_X1 U9778 ( .A1(n8726), .A2(n8725), .ZN(n8733) );
  AOI211_X1 U9779 ( .C1(n8726), .C2(n8725), .A(n10357), .B(n8733), .ZN(n8731)
         );
  INV_X1 U9780 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n8729) );
  NAND2_X1 U9781 ( .A1(n10364), .A2(n8738), .ZN(n8728) );
  NAND2_X1 U9782 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(P2_U3152), .ZN(n8727) );
  OAI211_X1 U9783 ( .C1(n8741), .C2(n8729), .A(n8728), .B(n8727), .ZN(n8730)
         );
  OR3_X1 U9784 ( .A1(n8732), .A2(n8731), .A3(n8730), .ZN(P2_U3262) );
  NOR2_X1 U9785 ( .A1(n8736), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n8748) );
  AND2_X1 U9786 ( .A1(n8736), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n8747) );
  NOR2_X1 U9787 ( .A1(n8748), .A2(n8747), .ZN(n8734) );
  XNOR2_X1 U9788 ( .A(n8746), .B(n8734), .ZN(n8735) );
  NAND2_X1 U9789 ( .A1(n8735), .A2(n10334), .ZN(n8745) );
  XNOR2_X1 U9790 ( .A(n8736), .B(n8752), .ZN(n8751) );
  XNOR2_X1 U9791 ( .A(n8751), .B(n8750), .ZN(n8743) );
  INV_X1 U9792 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n8740) );
  OAI21_X1 U9793 ( .B1(n8741), .B2(n8740), .A(n8739), .ZN(n8742) );
  AOI21_X1 U9794 ( .B1(n10333), .B2(n8743), .A(n8742), .ZN(n8744) );
  OAI211_X1 U9795 ( .C1(n10335), .C2(n8753), .A(n8745), .B(n8744), .ZN(
        P2_U3263) );
  INV_X1 U9796 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n8749) );
  XNOR2_X1 U9797 ( .A(n8759), .B(n8749), .ZN(n8757) );
  NAND2_X1 U9798 ( .A1(n8751), .A2(n8750), .ZN(n8755) );
  NAND2_X1 U9799 ( .A1(n8753), .A2(n8752), .ZN(n8754) );
  NAND2_X1 U9800 ( .A1(n8755), .A2(n8754), .ZN(n8758) );
  XNOR2_X1 U9801 ( .A(n8758), .B(n9238), .ZN(n8756) );
  OAI22_X1 U9802 ( .A1(n10357), .A2(n8757), .B1(n8756), .B2(n10353), .ZN(n8763) );
  XNOR2_X1 U9803 ( .A(n8758), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n8762) );
  XNOR2_X1 U9804 ( .A(n8759), .B(P2_REG2_REG_19__SCAN_IN), .ZN(n8760) );
  OR2_X1 U9805 ( .A1(n10357), .A2(n8760), .ZN(n8761) );
  XNOR2_X1 U9806 ( .A(n8957), .B(n8771), .ZN(n8959) );
  NOR2_X1 U9807 ( .A1(n8766), .A2(n8765), .ZN(n10548) );
  INV_X1 U9808 ( .A(n10548), .ZN(n8767) );
  NOR2_X1 U9809 ( .A1(n10466), .A2(n8767), .ZN(n8775) );
  NOR2_X1 U9810 ( .A1(n8768), .A2(n8930), .ZN(n8769) );
  AOI211_X1 U9811 ( .C1(n10466), .C2(P2_REG2_REG_31__SCAN_IN), .A(n8775), .B(
        n8769), .ZN(n8770) );
  OAI21_X1 U9812 ( .B1(n8959), .B2(n8777), .A(n8770), .ZN(P2_U3265) );
  NOR2_X1 U9813 ( .A1(n8773), .A2(n8930), .ZN(n8774) );
  AOI211_X1 U9814 ( .C1(n10466), .C2(P2_REG2_REG_30__SCAN_IN), .A(n8775), .B(
        n8774), .ZN(n8776) );
  OAI21_X1 U9815 ( .B1(n8777), .B2(n10546), .A(n8776), .ZN(P2_U3266) );
  NAND2_X1 U9816 ( .A1(n8779), .A2(n8778), .ZN(n8780) );
  XOR2_X1 U9817 ( .A(n8783), .B(n8780), .Z(n8782) );
  AOI222_X1 U9818 ( .A1(n8937), .A2(n8782), .B1(n8821), .B2(n8915), .C1(n8781), 
        .C2(n8916), .ZN(n8973) );
  XOR2_X1 U9819 ( .A(n8784), .B(n8783), .Z(n8974) );
  INV_X1 U9820 ( .A(n8974), .ZN(n8792) );
  AND2_X1 U9821 ( .A1(n8970), .A2(n8804), .ZN(n8785) );
  NOR2_X1 U9822 ( .A1(n8786), .A2(n8785), .ZN(n8971) );
  NAND2_X1 U9823 ( .A1(n8971), .A2(n8926), .ZN(n8789) );
  AOI22_X1 U9824 ( .A1(n8787), .A2(n8945), .B1(P2_REG2_REG_27__SCAN_IN), .B2(
        n10466), .ZN(n8788) );
  OAI211_X1 U9825 ( .C1(n8790), .C2(n8930), .A(n8789), .B(n8788), .ZN(n8791)
         );
  AOI21_X1 U9826 ( .B1(n8792), .B2(n8933), .A(n8791), .ZN(n8793) );
  OAI21_X1 U9827 ( .B1(n10466), .B2(n8973), .A(n8793), .ZN(P2_U3269) );
  XOR2_X1 U9828 ( .A(n8795), .B(n8794), .Z(n8980) );
  XNOR2_X1 U9829 ( .A(n8796), .B(n8795), .ZN(n8797) );
  NAND2_X1 U9830 ( .A1(n8797), .A2(n8937), .ZN(n8976) );
  INV_X1 U9831 ( .A(n8976), .ZN(n8811) );
  INV_X1 U9832 ( .A(n8798), .ZN(n8799) );
  AOI22_X1 U9833 ( .A1(n8799), .A2(n8945), .B1(P2_REG2_REG_26__SCAN_IN), .B2(
        n10466), .ZN(n8800) );
  OAI21_X1 U9834 ( .B1(n8977), .B2(n8930), .A(n8800), .ZN(n8809) );
  NAND2_X1 U9835 ( .A1(n8801), .A2(n8982), .ZN(n8803) );
  NAND2_X1 U9836 ( .A1(n8801), .A2(n8834), .ZN(n8802) );
  NAND4_X1 U9837 ( .A1(n8804), .A2(n10429), .A3(n8803), .A4(n8802), .ZN(n8807)
         );
  INV_X1 U9838 ( .A(n8805), .ZN(n8806) );
  AND2_X1 U9839 ( .A1(n8807), .A2(n8806), .ZN(n8975) );
  NOR2_X1 U9840 ( .A1(n8975), .A2(n8909), .ZN(n8808) );
  AOI211_X1 U9841 ( .C1(n8811), .C2(n8810), .A(n8809), .B(n8808), .ZN(n8812)
         );
  OAI21_X1 U9842 ( .B1(n8980), .B2(n8952), .A(n8812), .ZN(P2_U3270) );
  XNOR2_X1 U9843 ( .A(n8814), .B(n8813), .ZN(n8985) );
  XNOR2_X1 U9844 ( .A(n8982), .B(n8834), .ZN(n8815) );
  NOR2_X1 U9845 ( .A1(n8815), .A2(n10545), .ZN(n8981) );
  AOI22_X1 U9846 ( .A1(n10466), .A2(P2_REG2_REG_25__SCAN_IN), .B1(n8816), .B2(
        n8945), .ZN(n8817) );
  OAI21_X1 U9847 ( .B1(n8818), .B2(n8930), .A(n8817), .ZN(n8824) );
  XNOR2_X1 U9848 ( .A(n8820), .B(n8819), .ZN(n8822) );
  AOI222_X1 U9849 ( .A1(n8937), .A2(n8822), .B1(n8821), .B2(n8916), .C1(n8843), 
        .C2(n8915), .ZN(n8984) );
  NOR2_X1 U9850 ( .A1(n8984), .A2(n10466), .ZN(n8823) );
  AOI211_X1 U9851 ( .C1(n8955), .C2(n8981), .A(n8824), .B(n8823), .ZN(n8825)
         );
  OAI21_X1 U9852 ( .B1(n8985), .B2(n8952), .A(n8825), .ZN(P2_U3271) );
  NAND2_X1 U9853 ( .A1(n5367), .A2(n8826), .ZN(n8827) );
  XNOR2_X1 U9854 ( .A(n8828), .B(n8827), .ZN(n8830) );
  AOI222_X1 U9855 ( .A1(n8937), .A2(n8830), .B1(n8829), .B2(n8916), .C1(n8864), 
        .C2(n8915), .ZN(n8990) );
  OAI21_X1 U9856 ( .B1(n8833), .B2(n8832), .A(n8831), .ZN(n8986) );
  INV_X1 U9857 ( .A(n8849), .ZN(n8835) );
  AOI21_X1 U9858 ( .B1(n8987), .B2(n8835), .A(n5124), .ZN(n8988) );
  NAND2_X1 U9859 ( .A1(n8988), .A2(n8926), .ZN(n8839) );
  INV_X1 U9860 ( .A(n8836), .ZN(n8837) );
  AOI22_X1 U9861 ( .A1(n10466), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n8837), .B2(
        n8945), .ZN(n8838) );
  OAI211_X1 U9862 ( .C1(n8840), .C2(n8930), .A(n8839), .B(n8838), .ZN(n8841)
         );
  AOI21_X1 U9863 ( .B1(n8986), .B2(n8933), .A(n8841), .ZN(n8842) );
  OAI21_X1 U9864 ( .B1(n10466), .B2(n8990), .A(n8842), .ZN(P2_U3272) );
  OAI21_X1 U9865 ( .B1(n4880), .B2(n8845), .A(n5367), .ZN(n8844) );
  AOI222_X1 U9866 ( .A1(n8937), .A2(n8844), .B1(n8871), .B2(n8915), .C1(n8843), 
        .C2(n8916), .ZN(n8996) );
  INV_X1 U9867 ( .A(n8998), .ZN(n8847) );
  NAND2_X1 U9868 ( .A1(n8846), .A2(n8845), .ZN(n8992) );
  NAND3_X1 U9869 ( .A1(n8847), .A2(n8933), .A3(n8992), .ZN(n8856) );
  AND2_X1 U9870 ( .A1(n8993), .A2(n8858), .ZN(n8848) );
  NOR2_X1 U9871 ( .A1(n8849), .A2(n8848), .ZN(n8994) );
  INV_X1 U9872 ( .A(n8993), .ZN(n8853) );
  INV_X1 U9873 ( .A(n8850), .ZN(n8851) );
  AOI22_X1 U9874 ( .A1(n10466), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n8851), .B2(
        n8945), .ZN(n8852) );
  OAI21_X1 U9875 ( .B1(n8853), .B2(n8930), .A(n8852), .ZN(n8854) );
  AOI21_X1 U9876 ( .B1(n8994), .B2(n8926), .A(n8854), .ZN(n8855) );
  OAI211_X1 U9877 ( .C1(n10466), .C2(n8996), .A(n8856), .B(n8855), .ZN(
        P2_U3273) );
  XOR2_X1 U9878 ( .A(n8862), .B(n8857), .Z(n9003) );
  AOI21_X1 U9879 ( .B1(n8999), .B2(n8874), .A(n5125), .ZN(n9000) );
  AOI22_X1 U9880 ( .A1(n10466), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n8859), .B2(
        n8945), .ZN(n8860) );
  OAI21_X1 U9881 ( .B1(n8861), .B2(n8930), .A(n8860), .ZN(n8867) );
  XOR2_X1 U9882 ( .A(n8863), .B(n8862), .Z(n8865) );
  AOI222_X1 U9883 ( .A1(n8937), .A2(n8865), .B1(n8887), .B2(n8915), .C1(n8864), 
        .C2(n8916), .ZN(n9002) );
  NOR2_X1 U9884 ( .A1(n9002), .A2(n10466), .ZN(n8866) );
  AOI211_X1 U9885 ( .C1(n9000), .C2(n8926), .A(n8867), .B(n8866), .ZN(n8868)
         );
  OAI21_X1 U9886 ( .B1(n9003), .B2(n8952), .A(n8868), .ZN(P2_U3274) );
  XOR2_X1 U9887 ( .A(n8869), .B(n8882), .Z(n8872) );
  AOI222_X1 U9888 ( .A1(n8937), .A2(n8872), .B1(n8871), .B2(n8916), .C1(n8870), 
        .C2(n8915), .ZN(n9007) );
  INV_X1 U9889 ( .A(n8874), .ZN(n8875) );
  AOI21_X1 U9890 ( .B1(n9004), .B2(n8891), .A(n8875), .ZN(n9005) );
  INV_X1 U9891 ( .A(n8876), .ZN(n8877) );
  AOI22_X1 U9892 ( .A1(n10466), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n8877), .B2(
        n8945), .ZN(n8878) );
  OAI21_X1 U9893 ( .B1(n8879), .B2(n8930), .A(n8878), .ZN(n8884) );
  AOI21_X1 U9894 ( .B1(n8882), .B2(n8881), .A(n8880), .ZN(n9008) );
  NOR2_X1 U9895 ( .A1(n9008), .A2(n8952), .ZN(n8883) );
  AOI211_X1 U9896 ( .C1(n9005), .C2(n8926), .A(n8884), .B(n8883), .ZN(n8885)
         );
  OAI21_X1 U9897 ( .B1(n10466), .B2(n9007), .A(n8885), .ZN(P2_U3275) );
  XNOR2_X1 U9898 ( .A(n8896), .B(n8886), .ZN(n8888) );
  AOI222_X1 U9899 ( .A1(n8937), .A2(n8888), .B1(n8887), .B2(n8916), .C1(n8917), 
        .C2(n8915), .ZN(n9015) );
  NAND2_X1 U9900 ( .A1(n8889), .A2(n9011), .ZN(n8890) );
  AND2_X1 U9901 ( .A1(n8891), .A2(n8890), .ZN(n9012) );
  NAND2_X1 U9902 ( .A1(n9011), .A2(n8943), .ZN(n8894) );
  AOI22_X1 U9903 ( .A1(n10466), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n8892), .B2(
        n8945), .ZN(n8893) );
  NAND2_X1 U9904 ( .A1(n8894), .A2(n8893), .ZN(n8895) );
  AOI21_X1 U9905 ( .B1(n9012), .B2(n8926), .A(n8895), .ZN(n8899) );
  OR2_X1 U9906 ( .A1(n8897), .A2(n8896), .ZN(n9010) );
  NAND3_X1 U9907 ( .A1(n9010), .A2(n9009), .A3(n8933), .ZN(n8898) );
  OAI211_X1 U9908 ( .C1(n9015), .C2(n10466), .A(n8899), .B(n8898), .ZN(
        P2_U3276) );
  XNOR2_X1 U9909 ( .A(n8903), .B(n8900), .ZN(n8902) );
  AOI21_X1 U9910 ( .B1(n8902), .B2(n8937), .A(n8901), .ZN(n9235) );
  XNOR2_X1 U9911 ( .A(n8904), .B(n8903), .ZN(n9237) );
  NOR2_X1 U9912 ( .A1(n9242), .A2(n8923), .ZN(n8925) );
  XNOR2_X1 U9913 ( .A(n8925), .B(n9232), .ZN(n8905) );
  NAND2_X1 U9914 ( .A1(n8905), .A2(n10429), .ZN(n9233) );
  OAI22_X1 U9915 ( .A1(n8810), .A2(n8749), .B1(n8906), .B2(n10454), .ZN(n8907)
         );
  AOI21_X1 U9916 ( .B1(n9232), .B2(n8943), .A(n8907), .ZN(n8908) );
  OAI21_X1 U9917 ( .B1(n9233), .B2(n8909), .A(n8908), .ZN(n8910) );
  AOI21_X1 U9918 ( .B1(n9237), .B2(n8933), .A(n8910), .ZN(n8911) );
  OAI21_X1 U9919 ( .B1(n10466), .B2(n9235), .A(n8911), .ZN(P2_U3277) );
  OAI211_X1 U9920 ( .C1(n5302), .C2(n8913), .A(n8912), .B(n8937), .ZN(n8919)
         );
  AOI22_X1 U9921 ( .A1(n8917), .A2(n8916), .B1(n8915), .B2(n8914), .ZN(n8918)
         );
  OAI21_X1 U9922 ( .B1(n8922), .B2(n8921), .A(n8920), .ZN(n9241) );
  AND2_X1 U9923 ( .A1(n9242), .A2(n8923), .ZN(n8924) );
  NOR2_X1 U9924 ( .A1(n8925), .A2(n8924), .ZN(n9243) );
  NAND2_X1 U9925 ( .A1(n9243), .A2(n8926), .ZN(n8929) );
  AOI22_X1 U9926 ( .A1(n10466), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n8927), .B2(
        n8945), .ZN(n8928) );
  OAI211_X1 U9927 ( .C1(n8931), .C2(n8930), .A(n8929), .B(n8928), .ZN(n8932)
         );
  AOI21_X1 U9928 ( .B1(n9241), .B2(n8933), .A(n8932), .ZN(n8934) );
  OAI21_X1 U9929 ( .B1(n10466), .B2(n9245), .A(n8934), .ZN(P2_U3278) );
  XOR2_X1 U9930 ( .A(n8950), .B(n8935), .Z(n8938) );
  AOI21_X1 U9931 ( .B1(n8938), .B2(n8937), .A(n8936), .ZN(n9254) );
  NAND2_X1 U9932 ( .A1(n7105), .A2(n8939), .ZN(n8940) );
  NAND2_X1 U9933 ( .A1(n8940), .A2(n10429), .ZN(n8941) );
  NOR2_X1 U9934 ( .A1(n8942), .A2(n8941), .ZN(n9252) );
  INV_X1 U9935 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8948) );
  NAND2_X1 U9936 ( .A1(n7105), .A2(n8943), .ZN(n8947) );
  NAND2_X1 U9937 ( .A1(n8945), .A2(n8944), .ZN(n8946) );
  OAI211_X1 U9938 ( .C1(n8810), .C2(n8948), .A(n8947), .B(n8946), .ZN(n8954)
         );
  OAI21_X1 U9939 ( .B1(n8951), .B2(n8950), .A(n8949), .ZN(n9255) );
  NOR2_X1 U9940 ( .A1(n9255), .A2(n8952), .ZN(n8953) );
  AOI211_X1 U9941 ( .C1(n9252), .C2(n8955), .A(n8954), .B(n8953), .ZN(n8956)
         );
  OAI21_X1 U9942 ( .B1(n10466), .B2(n9254), .A(n8956), .ZN(P2_U3280) );
  AOI21_X1 U9943 ( .B1(n8957), .B2(n10550), .A(n10548), .ZN(n8958) );
  OAI21_X1 U9944 ( .B1(n8959), .B2(n10545), .A(n8958), .ZN(n9273) );
  MUX2_X1 U9945 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n9273), .S(n10553), .Z(
        P2_U3551) );
  AOI22_X1 U9946 ( .A1(n8961), .A2(n10429), .B1(n10550), .B2(n8960), .ZN(n8962) );
  OAI211_X1 U9947 ( .C1(n8964), .C2(n9271), .A(n8963), .B(n8962), .ZN(n9274)
         );
  MUX2_X1 U9948 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n9274), .S(n10553), .Z(
        P2_U3549) );
  AOI22_X1 U9949 ( .A1(n8966), .A2(n10429), .B1(n10550), .B2(n8965), .ZN(n8967) );
  OAI211_X1 U9950 ( .C1(n8969), .C2(n9271), .A(n8968), .B(n8967), .ZN(n9275)
         );
  MUX2_X1 U9951 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n9275), .S(n10553), .Z(
        P2_U3548) );
  AOI22_X1 U9952 ( .A1(n8971), .A2(n10429), .B1(n10550), .B2(n8970), .ZN(n8972) );
  OAI211_X1 U9953 ( .C1(n8974), .C2(n9271), .A(n8973), .B(n8972), .ZN(n9276)
         );
  MUX2_X1 U9954 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n9276), .S(n10553), .Z(
        P2_U3547) );
  OAI211_X1 U9955 ( .C1(n8977), .C2(n10536), .A(n8976), .B(n8975), .ZN(n8978)
         );
  INV_X1 U9956 ( .A(n8978), .ZN(n8979) );
  OAI21_X1 U9957 ( .B1(n8980), .B2(n9271), .A(n8979), .ZN(n9277) );
  MUX2_X1 U9958 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n9277), .S(n10553), .Z(
        P2_U3546) );
  AOI21_X1 U9959 ( .B1(n10550), .B2(n8982), .A(n8981), .ZN(n8983) );
  OAI211_X1 U9960 ( .C1(n8985), .C2(n9271), .A(n8984), .B(n8983), .ZN(n9278)
         );
  MUX2_X1 U9961 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n9278), .S(n10553), .Z(
        P2_U3545) );
  INV_X1 U9962 ( .A(n8986), .ZN(n8991) );
  AOI22_X1 U9963 ( .A1(n8988), .A2(n10429), .B1(n10550), .B2(n8987), .ZN(n8989) );
  OAI211_X1 U9964 ( .C1(n8991), .C2(n9271), .A(n8990), .B(n8989), .ZN(n9279)
         );
  MUX2_X1 U9965 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n9279), .S(n10553), .Z(
        P2_U3544) );
  NAND2_X1 U9966 ( .A1(n8992), .A2(n10541), .ZN(n8997) );
  AOI22_X1 U9967 ( .A1(n8994), .A2(n10429), .B1(n10550), .B2(n8993), .ZN(n8995) );
  OAI211_X1 U9968 ( .C1(n8998), .C2(n8997), .A(n8996), .B(n8995), .ZN(n9280)
         );
  MUX2_X1 U9969 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n9280), .S(n10553), .Z(
        P2_U3543) );
  AOI22_X1 U9970 ( .A1(n9000), .A2(n10429), .B1(n10550), .B2(n8999), .ZN(n9001) );
  OAI211_X1 U9971 ( .C1(n9003), .C2(n9271), .A(n9002), .B(n9001), .ZN(n9281)
         );
  MUX2_X1 U9972 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n9281), .S(n10553), .Z(
        P2_U3542) );
  AOI22_X1 U9973 ( .A1(n9005), .A2(n10429), .B1(n10550), .B2(n9004), .ZN(n9006) );
  OAI211_X1 U9974 ( .C1(n9008), .C2(n9271), .A(n9007), .B(n9006), .ZN(n9282)
         );
  MUX2_X1 U9975 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n9282), .S(n10553), .Z(
        P2_U3541) );
  NAND3_X1 U9976 ( .A1(n9010), .A2(n9009), .A3(n10541), .ZN(n9014) );
  AOI22_X1 U9977 ( .A1(n9012), .A2(n10429), .B1(n10550), .B2(n9011), .ZN(n9013) );
  NAND3_X1 U9978 ( .A1(n9015), .A2(n9014), .A3(n9013), .ZN(n9283) );
  MUX2_X1 U9979 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n9283), .S(n10553), .Z(
        P2_U3540) );
  XNOR2_X1 U9980 ( .A(n9222), .B(keyinput_125), .ZN(n9231) );
  INV_X1 U9981 ( .A(keyinput_124), .ZN(n9108) );
  INV_X1 U9982 ( .A(keyinput_123), .ZN(n9106) );
  INV_X1 U9983 ( .A(keyinput_122), .ZN(n9104) );
  INV_X1 U9984 ( .A(keyinput_118), .ZN(n9098) );
  OAI22_X1 U9985 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(keyinput_114), .B1(
        keyinput_115), .B2(P2_REG3_REG_24__SCAN_IN), .ZN(n9016) );
  AOI221_X1 U9986 ( .B1(P2_REG3_REG_17__SCAN_IN), .B2(keyinput_114), .C1(
        P2_REG3_REG_24__SCAN_IN), .C2(keyinput_115), .A(n9016), .ZN(n9096) );
  XOR2_X1 U9987 ( .A(P2_REG3_REG_7__SCAN_IN), .B(keyinput_99), .Z(n9077) );
  INV_X1 U9988 ( .A(keyinput_98), .ZN(n9071) );
  INV_X1 U9989 ( .A(keyinput_87), .ZN(n9053) );
  INV_X1 U9990 ( .A(SI_14_), .ZN(n9018) );
  OAI22_X1 U9991 ( .A1(n9121), .A2(keyinput_81), .B1(n9018), .B2(keyinput_82), 
        .ZN(n9017) );
  AOI221_X1 U9992 ( .B1(n9121), .B2(keyinput_81), .C1(keyinput_82), .C2(n9018), 
        .A(n9017), .ZN(n9051) );
  OAI22_X1 U9993 ( .A1(n9020), .A2(keyinput_76), .B1(keyinput_77), .B2(SI_19_), 
        .ZN(n9019) );
  AOI221_X1 U9994 ( .B1(n9020), .B2(keyinput_76), .C1(SI_19_), .C2(keyinput_77), .A(n9019), .ZN(n9041) );
  INV_X1 U9995 ( .A(keyinput_75), .ZN(n9039) );
  INV_X1 U9996 ( .A(SI_25_), .ZN(n9137) );
  INV_X1 U9997 ( .A(keyinput_71), .ZN(n9033) );
  INV_X1 U9998 ( .A(keyinput_70), .ZN(n9031) );
  INV_X1 U9999 ( .A(keyinput_69), .ZN(n9029) );
  AOI22_X1 U10000 ( .A1(P2_WR_REG_SCAN_IN), .A2(keyinput_64), .B1(SI_31_), 
        .B2(keyinput_65), .ZN(n9021) );
  OAI221_X1 U10001 ( .B1(P2_WR_REG_SCAN_IN), .B2(keyinput_64), .C1(SI_31_), 
        .C2(keyinput_65), .A(n9021), .ZN(n9025) );
  AOI22_X1 U10002 ( .A1(n9125), .A2(keyinput_67), .B1(n9023), .B2(keyinput_66), 
        .ZN(n9022) );
  OAI221_X1 U10003 ( .B1(n9125), .B2(keyinput_67), .C1(n9023), .C2(keyinput_66), .A(n9022), .ZN(n9024) );
  OAI22_X1 U10004 ( .A1(keyinput_68), .A2(n9027), .B1(n9025), .B2(n9024), .ZN(
        n9026) );
  AOI21_X1 U10005 ( .B1(keyinput_68), .B2(n9027), .A(n9026), .ZN(n9028) );
  AOI221_X1 U10006 ( .B1(SI_27_), .B2(keyinput_69), .C1(n9130), .C2(n9029), 
        .A(n9028), .ZN(n9030) );
  AOI221_X1 U10007 ( .B1(SI_26_), .B2(n9031), .C1(n9133), .C2(keyinput_70), 
        .A(n9030), .ZN(n9032) );
  AOI221_X1 U10008 ( .B1(SI_25_), .B2(keyinput_71), .C1(n9137), .C2(n9033), 
        .A(n9032), .ZN(n9036) );
  AOI22_X1 U10009 ( .A1(SI_23_), .A2(keyinput_73), .B1(SI_24_), .B2(
        keyinput_72), .ZN(n9034) );
  OAI221_X1 U10010 ( .B1(SI_23_), .B2(keyinput_73), .C1(SI_24_), .C2(
        keyinput_72), .A(n9034), .ZN(n9035) );
  AOI211_X1 U10011 ( .C1(SI_22_), .C2(keyinput_74), .A(n9036), .B(n9035), .ZN(
        n9037) );
  OAI21_X1 U10012 ( .B1(SI_22_), .B2(keyinput_74), .A(n9037), .ZN(n9038) );
  OAI221_X1 U10013 ( .B1(SI_21_), .B2(keyinput_75), .C1(n9144), .C2(n9039), 
        .A(n9038), .ZN(n9040) );
  INV_X1 U10014 ( .A(SI_18_), .ZN(n9149) );
  AOI22_X1 U10015 ( .A1(n9041), .A2(n9040), .B1(keyinput_78), .B2(n9149), .ZN(
        n9045) );
  INV_X1 U10016 ( .A(SI_16_), .ZN(n9043) );
  AOI22_X1 U10017 ( .A1(SI_17_), .A2(keyinput_79), .B1(n9043), .B2(keyinput_80), .ZN(n9042) );
  OAI221_X1 U10018 ( .B1(SI_17_), .B2(keyinput_79), .C1(n9043), .C2(
        keyinput_80), .A(n9042), .ZN(n9044) );
  AOI221_X1 U10019 ( .B1(keyinput_78), .B2(n9045), .C1(n9149), .C2(n9045), .A(
        n9044), .ZN(n9050) );
  INV_X1 U10020 ( .A(SI_13_), .ZN(n9152) );
  AOI22_X1 U10021 ( .A1(n9152), .A2(keyinput_83), .B1(keyinput_84), .B2(n9153), 
        .ZN(n9046) );
  OAI221_X1 U10022 ( .B1(n9152), .B2(keyinput_83), .C1(n9153), .C2(keyinput_84), .A(n9046), .ZN(n9049) );
  AOI22_X1 U10023 ( .A1(SI_10_), .A2(keyinput_86), .B1(SI_11_), .B2(
        keyinput_85), .ZN(n9047) );
  OAI221_X1 U10024 ( .B1(SI_10_), .B2(keyinput_86), .C1(SI_11_), .C2(
        keyinput_85), .A(n9047), .ZN(n9048) );
  AOI211_X1 U10025 ( .C1(n9051), .C2(n9050), .A(n9049), .B(n9048), .ZN(n9052)
         );
  AOI221_X1 U10026 ( .B1(SI_9_), .B2(n9053), .C1(n9161), .C2(keyinput_87), .A(
        n9052), .ZN(n9062) );
  AOI22_X1 U10027 ( .A1(SI_7_), .A2(keyinput_89), .B1(SI_8_), .B2(keyinput_88), 
        .ZN(n9054) );
  OAI221_X1 U10028 ( .B1(SI_7_), .B2(keyinput_89), .C1(SI_8_), .C2(keyinput_88), .A(n9054), .ZN(n9061) );
  OAI22_X1 U10029 ( .A1(SI_6_), .A2(keyinput_90), .B1(keyinput_91), .B2(SI_5_), 
        .ZN(n9055) );
  AOI221_X1 U10030 ( .B1(SI_6_), .B2(keyinput_90), .C1(SI_5_), .C2(keyinput_91), .A(n9055), .ZN(n9060) );
  XNOR2_X1 U10031 ( .A(n9056), .B(keyinput_93), .ZN(n9058) );
  XNOR2_X1 U10032 ( .A(SI_4_), .B(keyinput_92), .ZN(n9057) );
  NOR2_X1 U10033 ( .A1(n9058), .A2(n9057), .ZN(n9059) );
  OAI211_X1 U10034 ( .C1(n9062), .C2(n9061), .A(n9060), .B(n9059), .ZN(n9065)
         );
  INV_X1 U10035 ( .A(keyinput_94), .ZN(n9063) );
  MUX2_X1 U10036 ( .A(n9063), .B(keyinput_94), .S(SI_2_), .Z(n9064) );
  NAND2_X1 U10037 ( .A1(n9065), .A2(n9064), .ZN(n9068) );
  OAI22_X1 U10038 ( .A1(SI_0_), .A2(keyinput_96), .B1(keyinput_95), .B2(SI_1_), 
        .ZN(n9066) );
  AOI221_X1 U10039 ( .B1(SI_0_), .B2(keyinput_96), .C1(SI_1_), .C2(keyinput_95), .A(n9066), .ZN(n9067) );
  AOI22_X1 U10040 ( .A1(n9068), .A2(n9067), .B1(n5327), .B2(keyinput_97), .ZN(
        n9069) );
  OAI21_X1 U10041 ( .B1(n5327), .B2(keyinput_97), .A(n9069), .ZN(n9070) );
  OAI221_X1 U10042 ( .B1(P2_STATE_REG_SCAN_IN), .B2(n9071), .C1(P2_U3152), 
        .C2(keyinput_98), .A(n9070), .ZN(n9076) );
  AOI22_X1 U10043 ( .A1(n9184), .A2(keyinput_102), .B1(n6467), .B2(
        keyinput_103), .ZN(n9072) );
  OAI221_X1 U10044 ( .B1(n9184), .B2(keyinput_102), .C1(n6467), .C2(
        keyinput_103), .A(n9072), .ZN(n9075) );
  AOI22_X1 U10045 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(keyinput_100), .B1(
        P2_REG3_REG_14__SCAN_IN), .B2(keyinput_101), .ZN(n9073) );
  OAI221_X1 U10046 ( .B1(P2_REG3_REG_27__SCAN_IN), .B2(keyinput_100), .C1(
        P2_REG3_REG_14__SCAN_IN), .C2(keyinput_101), .A(n9073), .ZN(n9074) );
  AOI211_X1 U10047 ( .C1(n9077), .C2(n9076), .A(n9075), .B(n9074), .ZN(n9082)
         );
  INV_X1 U10048 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n9119) );
  AOI22_X1 U10049 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(keyinput_105), .B1(n9119), .B2(keyinput_104), .ZN(n9078) );
  OAI221_X1 U10050 ( .B1(P2_REG3_REG_19__SCAN_IN), .B2(keyinput_105), .C1(
        n9119), .C2(keyinput_104), .A(n9078), .ZN(n9081) );
  OAI22_X1 U10051 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(keyinput_107), .B1(
        keyinput_106), .B2(P2_REG3_REG_28__SCAN_IN), .ZN(n9079) );
  AOI221_X1 U10052 ( .B1(P2_REG3_REG_8__SCAN_IN), .B2(keyinput_107), .C1(
        P2_REG3_REG_28__SCAN_IN), .C2(keyinput_106), .A(n9079), .ZN(n9080) );
  OAI21_X1 U10053 ( .B1(n9082), .B2(n9081), .A(n9080), .ZN(n9087) );
  OAI22_X1 U10054 ( .A1(n9084), .A2(keyinput_109), .B1(keyinput_108), .B2(
        P2_REG3_REG_1__SCAN_IN), .ZN(n9083) );
  AOI221_X1 U10055 ( .B1(n9084), .B2(keyinput_109), .C1(P2_REG3_REG_1__SCAN_IN), .C2(keyinput_108), .A(n9083), .ZN(n9086) );
  NOR2_X1 U10056 ( .A1(n6495), .A2(keyinput_110), .ZN(n9085) );
  AOI221_X1 U10057 ( .B1(n9087), .B2(n9086), .C1(keyinput_110), .C2(n6495), 
        .A(n9085), .ZN(n9090) );
  AOI22_X1 U10058 ( .A1(P2_REG3_REG_25__SCAN_IN), .A2(keyinput_111), .B1(n6551), .B2(keyinput_112), .ZN(n9088) );
  OAI221_X1 U10059 ( .B1(P2_REG3_REG_25__SCAN_IN), .B2(keyinput_111), .C1(
        n6551), .C2(keyinput_112), .A(n9088), .ZN(n9089) );
  AOI211_X1 U10060 ( .C1(n9092), .C2(keyinput_113), .A(n9090), .B(n9089), .ZN(
        n9091) );
  OAI21_X1 U10061 ( .B1(n9092), .B2(keyinput_113), .A(n9091), .ZN(n9095) );
  AOI22_X1 U10062 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(keyinput_117), .B1(n9202), 
        .B2(keyinput_116), .ZN(n9093) );
  OAI221_X1 U10063 ( .B1(P2_REG3_REG_9__SCAN_IN), .B2(keyinput_117), .C1(n9202), .C2(keyinput_116), .A(n9093), .ZN(n9094) );
  AOI21_X1 U10064 ( .B1(n9096), .B2(n9095), .A(n9094), .ZN(n9097) );
  AOI221_X1 U10065 ( .B1(P2_REG3_REG_0__SCAN_IN), .B2(keyinput_118), .C1(n7294), .C2(n9098), .A(n9097), .ZN(n9101) );
  AOI22_X1 U10066 ( .A1(P2_REG3_REG_20__SCAN_IN), .A2(keyinput_119), .B1(n9210), .B2(keyinput_120), .ZN(n9099) );
  OAI221_X1 U10067 ( .B1(P2_REG3_REG_20__SCAN_IN), .B2(keyinput_119), .C1(
        n9210), .C2(keyinput_120), .A(n9099), .ZN(n9100) );
  AOI211_X1 U10068 ( .C1(n9209), .C2(keyinput_121), .A(n9101), .B(n9100), .ZN(
        n9102) );
  OAI21_X1 U10069 ( .B1(n9209), .B2(keyinput_121), .A(n9102), .ZN(n9103) );
  OAI221_X1 U10070 ( .B1(P2_REG3_REG_11__SCAN_IN), .B2(keyinput_122), .C1(
        n9215), .C2(n9104), .A(n9103), .ZN(n9105) );
  OAI221_X1 U10071 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(keyinput_123), .C1(n9219), .C2(n9106), .A(n9105), .ZN(n9107) );
  OAI221_X1 U10072 ( .B1(P2_REG3_REG_18__SCAN_IN), .B2(n9108), .C1(n6572), 
        .C2(keyinput_124), .A(n9107), .ZN(n9230) );
  INV_X1 U10073 ( .A(keyinput_127), .ZN(n9111) );
  OAI22_X1 U10074 ( .A1(n9112), .A2(keyinput_127), .B1(n9114), .B2(
        keyinput_126), .ZN(n9109) );
  AOI21_X1 U10075 ( .B1(n9114), .B2(keyinput_126), .A(n9109), .ZN(n9110) );
  OAI21_X1 U10076 ( .B1(P2_REG3_REG_15__SCAN_IN), .B2(n9111), .A(n9110), .ZN(
        n9229) );
  INV_X1 U10077 ( .A(keyinput_63), .ZN(n9227) );
  AOI22_X1 U10078 ( .A1(n9114), .A2(keyinput_62), .B1(n9112), .B2(keyinput_63), 
        .ZN(n9113) );
  OAI21_X1 U10079 ( .B1(n9114), .B2(keyinput_62), .A(n9113), .ZN(n9226) );
  INV_X1 U10080 ( .A(keyinput_60), .ZN(n9221) );
  INV_X1 U10081 ( .A(keyinput_59), .ZN(n9218) );
  INV_X1 U10082 ( .A(keyinput_58), .ZN(n9216) );
  INV_X1 U10083 ( .A(keyinput_54), .ZN(n9207) );
  OAI22_X1 U10084 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(keyinput_50), .B1(
        P2_REG3_REG_24__SCAN_IN), .B2(keyinput_51), .ZN(n9115) );
  AOI221_X1 U10085 ( .B1(P2_REG3_REG_17__SCAN_IN), .B2(keyinput_50), .C1(
        keyinput_51), .C2(P2_REG3_REG_24__SCAN_IN), .A(n9115), .ZN(n9205) );
  AOI22_X1 U10086 ( .A1(P2_REG3_REG_21__SCAN_IN), .A2(keyinput_45), .B1(n7653), 
        .B2(keyinput_44), .ZN(n9116) );
  OAI221_X1 U10087 ( .B1(P2_REG3_REG_21__SCAN_IN), .B2(keyinput_45), .C1(n7653), .C2(keyinput_44), .A(n9116), .ZN(n9194) );
  OAI22_X1 U10088 ( .A1(n9119), .A2(keyinput_40), .B1(n9118), .B2(keyinput_41), 
        .ZN(n9117) );
  AOI221_X1 U10089 ( .B1(n9119), .B2(keyinput_40), .C1(keyinput_41), .C2(n9118), .A(n9117), .ZN(n9192) );
  INV_X1 U10090 ( .A(keyinput_34), .ZN(n9181) );
  NOR2_X1 U10091 ( .A1(P2_RD_REG_SCAN_IN), .A2(keyinput_33), .ZN(n9179) );
  INV_X1 U10092 ( .A(keyinput_23), .ZN(n9162) );
  OAI22_X1 U10093 ( .A1(n9121), .A2(keyinput_17), .B1(keyinput_15), .B2(SI_17_), .ZN(n9120) );
  AOI221_X1 U10094 ( .B1(n9121), .B2(keyinput_17), .C1(SI_17_), .C2(
        keyinput_15), .A(n9120), .ZN(n9159) );
  OAI22_X1 U10095 ( .A1(SI_20_), .A2(keyinput_12), .B1(keyinput_13), .B2(
        SI_19_), .ZN(n9122) );
  AOI221_X1 U10096 ( .B1(SI_20_), .B2(keyinput_12), .C1(SI_19_), .C2(
        keyinput_13), .A(n9122), .ZN(n9146) );
  INV_X1 U10097 ( .A(keyinput_11), .ZN(n9143) );
  INV_X1 U10098 ( .A(keyinput_7), .ZN(n9136) );
  INV_X1 U10099 ( .A(keyinput_6), .ZN(n9134) );
  INV_X1 U10100 ( .A(keyinput_5), .ZN(n9131) );
  AOI22_X1 U10101 ( .A1(SI_31_), .A2(keyinput_1), .B1(SI_30_), .B2(keyinput_2), 
        .ZN(n9123) );
  OAI221_X1 U10102 ( .B1(SI_31_), .B2(keyinput_1), .C1(SI_30_), .C2(keyinput_2), .A(n9123), .ZN(n9127) );
  AOI22_X1 U10103 ( .A1(P2_WR_REG_SCAN_IN), .A2(keyinput_0), .B1(n9125), .B2(
        keyinput_3), .ZN(n9124) );
  OAI221_X1 U10104 ( .B1(P2_WR_REG_SCAN_IN), .B2(keyinput_0), .C1(n9125), .C2(
        keyinput_3), .A(n9124), .ZN(n9126) );
  OAI22_X1 U10105 ( .A1(n9127), .A2(n9126), .B1(keyinput_4), .B2(SI_28_), .ZN(
        n9128) );
  AOI21_X1 U10106 ( .B1(keyinput_4), .B2(SI_28_), .A(n9128), .ZN(n9129) );
  AOI221_X1 U10107 ( .B1(SI_27_), .B2(n9131), .C1(n9130), .C2(keyinput_5), .A(
        n9129), .ZN(n9132) );
  AOI221_X1 U10108 ( .B1(SI_26_), .B2(n9134), .C1(n9133), .C2(keyinput_6), .A(
        n9132), .ZN(n9135) );
  AOI221_X1 U10109 ( .B1(SI_25_), .B2(keyinput_7), .C1(n9137), .C2(n9136), .A(
        n9135), .ZN(n9140) );
  AOI22_X1 U10110 ( .A1(SI_22_), .A2(keyinput_10), .B1(SI_24_), .B2(keyinput_8), .ZN(n9138) );
  OAI221_X1 U10111 ( .B1(SI_22_), .B2(keyinput_10), .C1(SI_24_), .C2(
        keyinput_8), .A(n9138), .ZN(n9139) );
  AOI211_X1 U10112 ( .C1(SI_23_), .C2(keyinput_9), .A(n9140), .B(n9139), .ZN(
        n9141) );
  OAI21_X1 U10113 ( .B1(SI_23_), .B2(keyinput_9), .A(n9141), .ZN(n9142) );
  OAI221_X1 U10114 ( .B1(SI_21_), .B2(keyinput_11), .C1(n9144), .C2(n9143), 
        .A(n9142), .ZN(n9145) );
  AOI22_X1 U10115 ( .A1(n9146), .A2(n9145), .B1(keyinput_14), .B2(n9149), .ZN(
        n9150) );
  AOI22_X1 U10116 ( .A1(SI_14_), .A2(keyinput_18), .B1(SI_16_), .B2(
        keyinput_16), .ZN(n9147) );
  OAI221_X1 U10117 ( .B1(SI_14_), .B2(keyinput_18), .C1(SI_16_), .C2(
        keyinput_16), .A(n9147), .ZN(n9148) );
  AOI221_X1 U10118 ( .B1(keyinput_14), .B2(n9150), .C1(n9149), .C2(n9150), .A(
        n9148), .ZN(n9158) );
  AOI22_X1 U10119 ( .A1(n9153), .A2(keyinput_20), .B1(n9152), .B2(keyinput_19), 
        .ZN(n9151) );
  OAI221_X1 U10120 ( .B1(n9153), .B2(keyinput_20), .C1(n9152), .C2(keyinput_19), .A(n9151), .ZN(n9157) );
  AOI22_X1 U10121 ( .A1(SI_11_), .A2(keyinput_21), .B1(n9155), .B2(keyinput_22), .ZN(n9154) );
  OAI221_X1 U10122 ( .B1(SI_11_), .B2(keyinput_21), .C1(n9155), .C2(
        keyinput_22), .A(n9154), .ZN(n9156) );
  AOI211_X1 U10123 ( .C1(n9159), .C2(n9158), .A(n9157), .B(n9156), .ZN(n9160)
         );
  AOI221_X1 U10124 ( .B1(SI_9_), .B2(n9162), .C1(n9161), .C2(keyinput_23), .A(
        n9160), .ZN(n9170) );
  AOI22_X1 U10125 ( .A1(SI_7_), .A2(keyinput_25), .B1(SI_8_), .B2(keyinput_24), 
        .ZN(n9163) );
  OAI221_X1 U10126 ( .B1(SI_7_), .B2(keyinput_25), .C1(SI_8_), .C2(keyinput_24), .A(n9163), .ZN(n9169) );
  OAI22_X1 U10127 ( .A1(n9165), .A2(keyinput_27), .B1(keyinput_29), .B2(SI_3_), 
        .ZN(n9164) );
  AOI221_X1 U10128 ( .B1(n9165), .B2(keyinput_27), .C1(SI_3_), .C2(keyinput_29), .A(n9164), .ZN(n9168) );
  OAI22_X1 U10129 ( .A1(SI_6_), .A2(keyinput_26), .B1(SI_4_), .B2(keyinput_28), 
        .ZN(n9166) );
  AOI221_X1 U10130 ( .B1(SI_6_), .B2(keyinput_26), .C1(keyinput_28), .C2(SI_4_), .A(n9166), .ZN(n9167) );
  OAI211_X1 U10131 ( .C1(n9170), .C2(n9169), .A(n9168), .B(n9167), .ZN(n9177)
         );
  INV_X1 U10132 ( .A(keyinput_30), .ZN(n9171) );
  MUX2_X1 U10133 ( .A(n9171), .B(keyinput_30), .S(SI_2_), .Z(n9176) );
  XNOR2_X1 U10134 ( .A(n9172), .B(keyinput_31), .ZN(n9175) );
  INV_X1 U10135 ( .A(SI_0_), .ZN(n9173) );
  XNOR2_X1 U10136 ( .A(keyinput_32), .B(n9173), .ZN(n9174) );
  AOI211_X1 U10137 ( .C1(n9177), .C2(n9176), .A(n9175), .B(n9174), .ZN(n9178)
         );
  AOI211_X1 U10138 ( .C1(P2_RD_REG_SCAN_IN), .C2(keyinput_33), .A(n9179), .B(
        n9178), .ZN(n9180) );
  AOI221_X1 U10139 ( .B1(P2_STATE_REG_SCAN_IN), .B2(keyinput_34), .C1(P2_U3152), .C2(n9181), .A(n9180), .ZN(n9188) );
  XNOR2_X1 U10140 ( .A(P2_REG3_REG_7__SCAN_IN), .B(keyinput_35), .ZN(n9187) );
  OAI22_X1 U10141 ( .A1(n6467), .A2(keyinput_39), .B1(n6522), .B2(keyinput_37), 
        .ZN(n9182) );
  AOI221_X1 U10142 ( .B1(n6467), .B2(keyinput_39), .C1(keyinput_37), .C2(n6522), .A(n9182), .ZN(n9186) );
  OAI22_X1 U10143 ( .A1(n9184), .A2(keyinput_38), .B1(P2_REG3_REG_27__SCAN_IN), 
        .B2(keyinput_36), .ZN(n9183) );
  AOI221_X1 U10144 ( .B1(n9184), .B2(keyinput_38), .C1(keyinput_36), .C2(
        P2_REG3_REG_27__SCAN_IN), .A(n9183), .ZN(n9185) );
  OAI211_X1 U10145 ( .C1(n9188), .C2(n9187), .A(n9186), .B(n9185), .ZN(n9191)
         );
  AOI22_X1 U10146 ( .A1(n8548), .A2(keyinput_42), .B1(n6434), .B2(keyinput_43), 
        .ZN(n9189) );
  OAI221_X1 U10147 ( .B1(n8548), .B2(keyinput_42), .C1(n6434), .C2(keyinput_43), .A(n9189), .ZN(n9190) );
  AOI21_X1 U10148 ( .B1(n9192), .B2(n9191), .A(n9190), .ZN(n9193) );
  OAI22_X1 U10149 ( .A1(n9194), .A2(n9193), .B1(keyinput_46), .B2(
        P2_REG3_REG_12__SCAN_IN), .ZN(n9195) );
  AOI21_X1 U10150 ( .B1(keyinput_46), .B2(P2_REG3_REG_12__SCAN_IN), .A(n9195), 
        .ZN(n9199) );
  AOI22_X1 U10151 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(keyinput_48), .B1(n9197), 
        .B2(keyinput_47), .ZN(n9196) );
  OAI221_X1 U10152 ( .B1(P2_REG3_REG_16__SCAN_IN), .B2(keyinput_48), .C1(n9197), .C2(keyinput_47), .A(n9196), .ZN(n9198) );
  AOI211_X1 U10153 ( .C1(P2_REG3_REG_5__SCAN_IN), .C2(keyinput_49), .A(n9199), 
        .B(n9198), .ZN(n9200) );
  OAI21_X1 U10154 ( .B1(P2_REG3_REG_5__SCAN_IN), .B2(keyinput_49), .A(n9200), 
        .ZN(n9204) );
  AOI22_X1 U10155 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(keyinput_53), .B1(n9202), 
        .B2(keyinput_52), .ZN(n9201) );
  OAI221_X1 U10156 ( .B1(P2_REG3_REG_9__SCAN_IN), .B2(keyinput_53), .C1(n9202), 
        .C2(keyinput_52), .A(n9201), .ZN(n9203) );
  AOI21_X1 U10157 ( .B1(n9205), .B2(n9204), .A(n9203), .ZN(n9206) );
  AOI221_X1 U10158 ( .B1(P2_REG3_REG_0__SCAN_IN), .B2(keyinput_54), .C1(n7294), 
        .C2(n9207), .A(n9206), .ZN(n9213) );
  OAI22_X1 U10159 ( .A1(n9210), .A2(keyinput_56), .B1(n9209), .B2(keyinput_57), 
        .ZN(n9208) );
  AOI221_X1 U10160 ( .B1(n9210), .B2(keyinput_56), .C1(keyinput_57), .C2(n9209), .A(n9208), .ZN(n9211) );
  OAI21_X1 U10161 ( .B1(keyinput_55), .B2(P2_REG3_REG_20__SCAN_IN), .A(n9211), 
        .ZN(n9212) );
  AOI211_X1 U10162 ( .C1(keyinput_55), .C2(P2_REG3_REG_20__SCAN_IN), .A(n9213), 
        .B(n9212), .ZN(n9214) );
  AOI221_X1 U10163 ( .B1(P2_REG3_REG_11__SCAN_IN), .B2(n9216), .C1(n9215), 
        .C2(keyinput_58), .A(n9214), .ZN(n9217) );
  AOI221_X1 U10164 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(keyinput_59), .C1(n9219), 
        .C2(n9218), .A(n9217), .ZN(n9220) );
  AOI221_X1 U10165 ( .B1(P2_REG3_REG_18__SCAN_IN), .B2(keyinput_60), .C1(n6572), .C2(n9221), .A(n9220), .ZN(n9224) );
  XNOR2_X1 U10166 ( .A(n9222), .B(keyinput_61), .ZN(n9223) );
  NOR2_X1 U10167 ( .A1(n9224), .A2(n9223), .ZN(n9225) );
  AOI211_X1 U10168 ( .C1(P2_REG3_REG_15__SCAN_IN), .C2(n9227), .A(n9226), .B(
        n9225), .ZN(n9228) );
  AOI211_X1 U10169 ( .C1(n9231), .C2(n9230), .A(n9229), .B(n9228), .ZN(n9240)
         );
  NAND2_X1 U10170 ( .A1(n9232), .A2(n10550), .ZN(n9234) );
  NAND3_X1 U10171 ( .A1(n9235), .A2(n9234), .A3(n9233), .ZN(n9236) );
  AOI21_X1 U10172 ( .B1(n9237), .B2(n10541), .A(n9236), .ZN(n9284) );
  MUX2_X1 U10173 ( .A(n9238), .B(n9284), .S(n10553), .Z(n9239) );
  XNOR2_X1 U10174 ( .A(n9240), .B(n9239), .ZN(P2_U3539) );
  INV_X1 U10175 ( .A(n9241), .ZN(n9246) );
  AOI22_X1 U10176 ( .A1(n9243), .A2(n10429), .B1(n10550), .B2(n9242), .ZN(
        n9244) );
  OAI211_X1 U10177 ( .C1(n9246), .C2(n9271), .A(n9245), .B(n9244), .ZN(n9287)
         );
  MUX2_X1 U10178 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n9287), .S(n10553), .Z(
        P2_U3538) );
  AOI211_X1 U10179 ( .C1(n10550), .C2(n9249), .A(n9248), .B(n9247), .ZN(n9250)
         );
  OAI21_X1 U10180 ( .B1(n9271), .B2(n9251), .A(n9250), .ZN(n9288) );
  MUX2_X1 U10181 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n9288), .S(n10553), .Z(
        P2_U3537) );
  AOI21_X1 U10182 ( .B1(n10550), .B2(n7105), .A(n9252), .ZN(n9253) );
  OAI211_X1 U10183 ( .C1(n9255), .C2(n9271), .A(n9254), .B(n9253), .ZN(n9289)
         );
  MUX2_X1 U10184 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n9289), .S(n10553), .Z(
        P2_U3536) );
  INV_X1 U10185 ( .A(n9256), .ZN(n9261) );
  AOI22_X1 U10186 ( .A1(n9258), .A2(n10429), .B1(n10550), .B2(n9257), .ZN(
        n9259) );
  OAI211_X1 U10187 ( .C1(n9261), .C2(n9271), .A(n9260), .B(n9259), .ZN(n9290)
         );
  MUX2_X1 U10188 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n9290), .S(n10553), .Z(
        P2_U3535) );
  AOI22_X1 U10189 ( .A1(n9263), .A2(n10429), .B1(n10550), .B2(n9262), .ZN(
        n9264) );
  OAI211_X1 U10190 ( .C1(n9266), .C2(n9271), .A(n9265), .B(n9264), .ZN(n9291)
         );
  MUX2_X1 U10191 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n9291), .S(n10553), .Z(
        P2_U3534) );
  AOI22_X1 U10192 ( .A1(n9268), .A2(n10429), .B1(n10550), .B2(n9267), .ZN(
        n9269) );
  OAI211_X1 U10193 ( .C1(n9272), .C2(n9271), .A(n9270), .B(n9269), .ZN(n9292)
         );
  MUX2_X1 U10194 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n9292), .S(n10553), .Z(
        P2_U3533) );
  MUX2_X1 U10195 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n9273), .S(n10557), .Z(
        P2_U3519) );
  MUX2_X1 U10196 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n9274), .S(n10557), .Z(
        P2_U3517) );
  MUX2_X1 U10197 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n9275), .S(n10557), .Z(
        P2_U3516) );
  MUX2_X1 U10198 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n9276), .S(n10557), .Z(
        P2_U3515) );
  MUX2_X1 U10199 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n9277), .S(n10557), .Z(
        P2_U3514) );
  MUX2_X1 U10200 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n9278), .S(n10557), .Z(
        P2_U3513) );
  MUX2_X1 U10201 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n9279), .S(n10557), .Z(
        P2_U3512) );
  MUX2_X1 U10202 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n9280), .S(n10557), .Z(
        P2_U3511) );
  MUX2_X1 U10203 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n9281), .S(n10557), .Z(
        P2_U3510) );
  MUX2_X1 U10204 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n9282), .S(n10557), .Z(
        P2_U3509) );
  MUX2_X1 U10205 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n9283), .S(n10557), .Z(
        P2_U3508) );
  INV_X1 U10206 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n9285) );
  MUX2_X1 U10207 ( .A(n9285), .B(n9284), .S(n10557), .Z(n9286) );
  INV_X1 U10208 ( .A(n9286), .ZN(P2_U3507) );
  MUX2_X1 U10209 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n9287), .S(n10557), .Z(
        P2_U3505) );
  MUX2_X1 U10210 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n9288), .S(n10557), .Z(
        P2_U3502) );
  MUX2_X1 U10211 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n9289), .S(n10557), .Z(
        P2_U3499) );
  MUX2_X1 U10212 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n9290), .S(n10557), .Z(
        P2_U3496) );
  MUX2_X1 U10213 ( .A(P2_REG0_REG_14__SCAN_IN), .B(n9291), .S(n10557), .Z(
        P2_U3493) );
  MUX2_X1 U10214 ( .A(P2_REG0_REG_13__SCAN_IN), .B(n9292), .S(n10557), .Z(
        P2_U3490) );
  INV_X1 U10215 ( .A(n9293), .ZN(n10110) );
  NOR4_X1 U10216 ( .A1(n9295), .A2(P2_IR_REG_30__SCAN_IN), .A3(n9294), .A4(
        P2_U3152), .ZN(n9296) );
  AOI21_X1 U10217 ( .B1(P1_DATAO_REG_31__SCAN_IN), .B2(n9297), .A(n9296), .ZN(
        n9298) );
  OAI21_X1 U10218 ( .B1(n10110), .B2(n8219), .A(n9298), .ZN(P2_U3327) );
  OAI222_X1 U10219 ( .A1(P2_U3152), .A2(n9299), .B1(n8219), .B2(n9301), .C1(
        n9300), .C2(n6811), .ZN(P2_U3328) );
  INV_X1 U10220 ( .A(n9302), .ZN(n9303) );
  MUX2_X1 U10221 ( .A(P2_IR_REG_0__SCAN_IN), .B(n9303), .S(P2_U3152), .Z(
        P2_U3358) );
  NAND2_X1 U10222 ( .A1(n9305), .A2(n9304), .ZN(n9306) );
  XOR2_X1 U10223 ( .A(n9307), .B(n9306), .Z(n9312) );
  OAI22_X1 U10224 ( .A1(n9978), .A2(n9431), .B1(n9430), .B2(n9976), .ZN(n9308)
         );
  AOI211_X1 U10225 ( .C1(n9434), .C2(n9967), .A(n9309), .B(n9308), .ZN(n9311)
         );
  NAND2_X1 U10226 ( .A1(n10068), .A2(n9435), .ZN(n9310) );
  OAI211_X1 U10227 ( .C1(n9312), .C2(n9438), .A(n9311), .B(n9310), .ZN(
        P1_U3213) );
  NAND2_X1 U10228 ( .A1(n9313), .A2(n9370), .ZN(n9314) );
  XOR2_X1 U10229 ( .A(n9315), .B(n9314), .Z(n9322) );
  INV_X1 U10230 ( .A(n9820), .ZN(n10019) );
  INV_X1 U10231 ( .A(n9316), .ZN(n9817) );
  OAI22_X1 U10232 ( .A1(n9392), .A2(n9817), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9317), .ZN(n9320) );
  OAI22_X1 U10233 ( .A1(n9337), .A2(n9431), .B1(n9430), .B2(n9318), .ZN(n9319)
         );
  AOI211_X1 U10234 ( .C1(n10019), .C2(n9435), .A(n9320), .B(n9319), .ZN(n9321)
         );
  OAI21_X1 U10235 ( .B1(n9322), .B2(n9438), .A(n9321), .ZN(P1_U3214) );
  AOI21_X1 U10236 ( .B1(n9325), .B2(n9324), .A(n9323), .ZN(n9329) );
  AND2_X1 U10237 ( .A1(P1_U3084), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9738) );
  OAI22_X1 U10238 ( .A1(n9338), .A2(n9430), .B1(n9431), .B2(n9907), .ZN(n9326)
         );
  AOI211_X1 U10239 ( .C1(n9434), .C2(n9878), .A(n9738), .B(n9326), .ZN(n9328)
         );
  NAND2_X1 U10240 ( .A1(n10039), .A2(n9435), .ZN(n9327) );
  OAI211_X1 U10241 ( .C1(n9329), .C2(n9438), .A(n9328), .B(n9327), .ZN(
        P1_U3217) );
  INV_X1 U10242 ( .A(n9330), .ZN(n9332) );
  NAND2_X1 U10243 ( .A1(n9332), .A2(n9331), .ZN(n9333) );
  XNOR2_X1 U10244 ( .A(n9334), .B(n9333), .ZN(n9342) );
  INV_X1 U10245 ( .A(n9855), .ZN(n9336) );
  OAI22_X1 U10246 ( .A1(n9392), .A2(n9336), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9335), .ZN(n9340) );
  OAI22_X1 U10247 ( .A1(n9338), .A2(n9431), .B1(n9430), .B2(n9337), .ZN(n9339)
         );
  AOI211_X1 U10248 ( .C1(n10030), .C2(n9435), .A(n9340), .B(n9339), .ZN(n9341)
         );
  OAI21_X1 U10249 ( .B1(n9342), .B2(n9438), .A(n9341), .ZN(P1_U3221) );
  OAI21_X1 U10250 ( .B1(n9344), .B2(n9343), .A(n9411), .ZN(n9348) );
  AOI22_X1 U10251 ( .A1(n9434), .A2(n9790), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3084), .ZN(n9346) );
  AOI22_X1 U10252 ( .A1(n9417), .A2(n9824), .B1(n9416), .B2(n9785), .ZN(n9345)
         );
  OAI211_X1 U10253 ( .C1(n9792), .C2(n9409), .A(n9346), .B(n9345), .ZN(n9347)
         );
  AOI21_X1 U10254 ( .B1(n9348), .B2(n9413), .A(n9347), .ZN(n9349) );
  INV_X1 U10255 ( .A(n9349), .ZN(P1_U3223) );
  AOI21_X1 U10256 ( .B1(n9351), .B2(n9422), .A(n9350), .ZN(n9356) );
  AOI22_X1 U10257 ( .A1(n9416), .A2(n9899), .B1(n9417), .B2(n9706), .ZN(n9353)
         );
  OAI211_X1 U10258 ( .C1(n9392), .C2(n9932), .A(n9353), .B(n9352), .ZN(n9354)
         );
  AOI21_X1 U10259 ( .B1(n10058), .B2(n9435), .A(n9354), .ZN(n9355) );
  OAI21_X1 U10260 ( .B1(n9356), .B2(n9438), .A(n9355), .ZN(P1_U3224) );
  XNOR2_X1 U10261 ( .A(n9358), .B(n9357), .ZN(n9359) );
  XNOR2_X1 U10262 ( .A(n9360), .B(n9359), .ZN(n9366) );
  OAI21_X1 U10263 ( .B1(n9392), .B2(n9362), .A(n9361), .ZN(n9364) );
  OAI22_X1 U10264 ( .A1(n9947), .A2(n9431), .B1(n9430), .B2(n9907), .ZN(n9363)
         );
  AOI211_X1 U10265 ( .C1(n10049), .C2(n9435), .A(n9364), .B(n9363), .ZN(n9365)
         );
  OAI21_X1 U10266 ( .B1(n9366), .B2(n9438), .A(n9365), .ZN(P1_U3226) );
  INV_X1 U10267 ( .A(n9367), .ZN(n9372) );
  AOI21_X1 U10268 ( .B1(n9368), .B2(n9370), .A(n9369), .ZN(n9371) );
  OAI21_X1 U10269 ( .B1(n9372), .B2(n9371), .A(n9413), .ZN(n9376) );
  AOI22_X1 U10270 ( .A1(n9434), .A2(n9809), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3084), .ZN(n9375) );
  AOI22_X1 U10271 ( .A1(n9417), .A2(n9831), .B1(n9416), .B2(n9806), .ZN(n9374)
         );
  NAND2_X1 U10272 ( .A1(n10014), .A2(n9435), .ZN(n9373) );
  NAND4_X1 U10273 ( .A1(n9376), .A2(n9375), .A3(n9374), .A4(n9373), .ZN(
        P1_U3227) );
  INV_X1 U10274 ( .A(n9377), .ZN(n9379) );
  NOR2_X1 U10275 ( .A1(n9379), .A2(n9378), .ZN(n9380) );
  XNOR2_X1 U10276 ( .A(n9381), .B(n9380), .ZN(n9387) );
  INV_X1 U10277 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n9382) );
  OAI22_X1 U10278 ( .A1(n9392), .A2(n9383), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9382), .ZN(n9385) );
  OAI22_X1 U10279 ( .A1(n9405), .A2(n9431), .B1(n9430), .B2(n9393), .ZN(n9384)
         );
  AOI211_X1 U10280 ( .C1(n10035), .C2(n9435), .A(n9385), .B(n9384), .ZN(n9386)
         );
  OAI21_X1 U10281 ( .B1(n9387), .B2(n9438), .A(n9386), .ZN(P1_U3231) );
  XOR2_X1 U10282 ( .A(n9389), .B(n9388), .Z(n9398) );
  INV_X1 U10283 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n9390) );
  OAI22_X1 U10284 ( .A1(n9392), .A2(n9391), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9390), .ZN(n9396) );
  OAI22_X1 U10285 ( .A1(n9394), .A2(n9430), .B1(n9431), .B2(n9393), .ZN(n9395)
         );
  AOI211_X1 U10286 ( .C1(n9835), .C2(n9435), .A(n9396), .B(n9395), .ZN(n9397)
         );
  OAI21_X1 U10287 ( .B1(n9398), .B2(n9438), .A(n9397), .ZN(P1_U3233) );
  XNOR2_X1 U10288 ( .A(n9400), .B(n9399), .ZN(n9401) );
  XNOR2_X1 U10289 ( .A(n9402), .B(n9401), .ZN(n9403) );
  NAND2_X1 U10290 ( .A1(n9403), .A2(n9413), .ZN(n9408) );
  AND2_X1 U10291 ( .A1(P1_U3084), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n10303) );
  OAI22_X1 U10292 ( .A1(n9927), .A2(n9431), .B1(n9430), .B2(n9405), .ZN(n9406)
         );
  AOI211_X1 U10293 ( .C1(n9434), .C2(n9894), .A(n10303), .B(n9406), .ZN(n9407)
         );
  OAI211_X1 U10294 ( .C1(n9896), .C2(n9409), .A(n9408), .B(n9407), .ZN(
        P1_U3236) );
  OAI211_X1 U10295 ( .C1(n9415), .C2(n9414), .A(n9413), .B(n9412), .ZN(n9421)
         );
  AOI22_X1 U10296 ( .A1(n9434), .A2(n9776), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3084), .ZN(n9420) );
  AOI22_X1 U10297 ( .A1(n9417), .A2(n9806), .B1(n9416), .B2(n9704), .ZN(n9419)
         );
  NAND2_X1 U10298 ( .A1(n10003), .A2(n9435), .ZN(n9418) );
  NAND4_X1 U10299 ( .A1(n9421), .A2(n9420), .A3(n9419), .A4(n9418), .ZN(
        P1_U3238) );
  INV_X1 U10300 ( .A(n9422), .ZN(n9429) );
  INV_X1 U10301 ( .A(n9424), .ZN(n9426) );
  NAND2_X1 U10302 ( .A1(n9426), .A2(n9425), .ZN(n9428) );
  AOI22_X1 U10303 ( .A1(n9429), .A2(n9423), .B1(n9428), .B2(n9427), .ZN(n9439)
         );
  OAI22_X1 U10304 ( .A1(n9948), .A2(n9431), .B1(n9430), .B2(n9947), .ZN(n9432)
         );
  AOI211_X1 U10305 ( .C1(n9434), .C2(n9956), .A(n9433), .B(n9432), .ZN(n9437)
         );
  NAND2_X1 U10306 ( .A1(n10062), .A2(n9435), .ZN(n9436) );
  OAI211_X1 U10307 ( .C1(n9439), .C2(n9438), .A(n9437), .B(n9436), .ZN(
        P1_U3239) );
  NAND2_X1 U10308 ( .A1(n9622), .A2(n10411), .ZN(n9689) );
  NOR3_X1 U10309 ( .A1(n9647), .A2(n9441), .A3(n9442), .ZN(n9528) );
  INV_X1 U10310 ( .A(n9908), .ZN(n9673) );
  INV_X1 U10311 ( .A(n9449), .ZN(n9477) );
  MUX2_X1 U10312 ( .A(n9562), .B(n9564), .S(n9477), .Z(n9443) );
  INV_X1 U10313 ( .A(n9567), .ZN(n9445) );
  MUX2_X1 U10314 ( .A(n9445), .B(n9444), .S(n9449), .Z(n9491) );
  AND2_X1 U10315 ( .A1(n9530), .A2(n9477), .ZN(n9486) );
  INV_X1 U10316 ( .A(n9486), .ZN(n9489) );
  NAND2_X1 U10317 ( .A1(n9558), .A2(n9449), .ZN(n9480) );
  INV_X1 U10318 ( .A(n9480), .ZN(n9487) );
  MUX2_X1 U10319 ( .A(n9710), .B(n9446), .S(n9449), .Z(n9473) );
  INV_X1 U10320 ( .A(n9473), .ZN(n9476) );
  INV_X1 U10321 ( .A(n9547), .ZN(n9448) );
  MUX2_X1 U10322 ( .A(n9448), .B(n9447), .S(n9449), .Z(n9472) );
  OAI21_X1 U10323 ( .B1(n9477), .B2(n9624), .A(n9452), .ZN(n9453) );
  NAND2_X1 U10324 ( .A1(n9461), .A2(n9454), .ZN(n9542) );
  AOI21_X1 U10325 ( .B1(n9460), .B2(n9455), .A(n9542), .ZN(n9456) );
  NOR2_X1 U10326 ( .A1(n9456), .A2(n9459), .ZN(n9465) );
  INV_X1 U10327 ( .A(n9457), .ZN(n9458) );
  NOR3_X1 U10328 ( .A1(n9460), .A2(n9459), .A3(n9458), .ZN(n9463) );
  INV_X1 U10329 ( .A(n9461), .ZN(n9462) );
  NOR2_X1 U10330 ( .A1(n9463), .A2(n9462), .ZN(n9464) );
  MUX2_X1 U10331 ( .A(n9465), .B(n9464), .S(n9449), .Z(n9467) );
  MUX2_X1 U10332 ( .A(n9537), .B(n9546), .S(n9449), .Z(n9466) );
  INV_X1 U10333 ( .A(n9468), .ZN(n9531) );
  INV_X1 U10334 ( .A(n9545), .ZN(n9469) );
  MUX2_X1 U10335 ( .A(n9531), .B(n9469), .S(n9449), .Z(n9471) );
  INV_X1 U10336 ( .A(n9551), .ZN(n9478) );
  OAI21_X1 U10337 ( .B1(n9482), .B2(n9478), .A(n9477), .ZN(n9479) );
  MUX2_X1 U10338 ( .A(n9480), .B(n9479), .S(n9554), .Z(n9484) );
  INV_X1 U10339 ( .A(n9973), .ZN(n9964) );
  OAI211_X1 U10340 ( .C1(n9482), .C2(n9481), .A(n9556), .B(n9449), .ZN(n9483)
         );
  NAND3_X1 U10341 ( .A1(n9484), .A2(n9964), .A3(n9483), .ZN(n9485) );
  OAI21_X1 U10342 ( .B1(n9487), .B2(n9486), .A(n9485), .ZN(n9488) );
  MUX2_X1 U10343 ( .A(n9922), .B(n9559), .S(n9449), .Z(n9490) );
  MUX2_X1 U10344 ( .A(n9571), .B(n9569), .S(n9449), .Z(n9492) );
  MUX2_X1 U10345 ( .A(n9573), .B(n9572), .S(n9449), .Z(n9493) );
  AOI211_X1 U10346 ( .C1(n9494), .C2(n9493), .A(n5133), .B(n9846), .ZN(n9505)
         );
  NAND2_X1 U10347 ( .A1(n9498), .A2(n9495), .ZN(n9578) );
  NAND2_X1 U10348 ( .A1(n9578), .A2(n9499), .ZN(n9501) );
  INV_X1 U10349 ( .A(n9496), .ZN(n9497) );
  NAND2_X1 U10350 ( .A1(n9498), .A2(n9497), .ZN(n9500) );
  AND2_X1 U10351 ( .A1(n9500), .A2(n9499), .ZN(n9576) );
  MUX2_X1 U10352 ( .A(n9501), .B(n9576), .S(n9449), .Z(n9502) );
  NAND2_X1 U10353 ( .A1(n9502), .A2(n9841), .ZN(n9504) );
  MUX2_X1 U10354 ( .A(n9575), .B(n9579), .S(n9449), .Z(n9503) );
  MUX2_X1 U10355 ( .A(n9581), .B(n9633), .S(n9449), .Z(n9506) );
  MUX2_X1 U10356 ( .A(n9606), .B(n9631), .S(n9449), .Z(n9507) );
  MUX2_X1 U10357 ( .A(n9609), .B(n9607), .S(n9449), .Z(n9508) );
  MUX2_X1 U10358 ( .A(n9747), .B(n9610), .S(n9449), .Z(n9509) );
  NAND3_X1 U10359 ( .A1(n9510), .A2(n9748), .A3(n9509), .ZN(n9511) );
  OAI211_X1 U10360 ( .C1(n9636), .C2(n9449), .A(n9511), .B(n9678), .ZN(n9518)
         );
  INV_X1 U10361 ( .A(n9615), .ZN(n9512) );
  NOR2_X1 U10362 ( .A1(n9518), .A2(n9512), .ZN(n9514) );
  NAND2_X1 U10363 ( .A1(n9519), .A2(n9513), .ZN(n9646) );
  OAI211_X1 U10364 ( .C1(n9514), .C2(n9646), .A(n9643), .B(n9449), .ZN(n9517)
         );
  NOR2_X1 U10365 ( .A1(n9742), .A2(n9618), .ZN(n9529) );
  NAND2_X1 U10366 ( .A1(n9986), .A2(n9529), .ZN(n9516) );
  NAND2_X1 U10367 ( .A1(n9515), .A2(n9702), .ZN(n9523) );
  AND2_X1 U10368 ( .A1(n9742), .A2(n9523), .ZN(n9642) );
  AOI21_X1 U10369 ( .B1(n9517), .B2(n9516), .A(n9642), .ZN(n9527) );
  NAND3_X1 U10370 ( .A1(n9518), .A2(n9643), .A3(n9616), .ZN(n9520) );
  AOI21_X1 U10371 ( .B1(n9520), .B2(n9519), .A(n9642), .ZN(n9522) );
  INV_X1 U10372 ( .A(n9702), .ZN(n9521) );
  NAND2_X1 U10373 ( .A1(n9986), .A2(n9521), .ZN(n9683) );
  OAI21_X1 U10374 ( .B1(n9522), .B2(n9449), .A(n9683), .ZN(n9526) );
  INV_X1 U10375 ( .A(n9523), .ZN(n9525) );
  INV_X1 U10376 ( .A(n9683), .ZN(n9524) );
  AOI21_X1 U10377 ( .B1(n9993), .B2(n9525), .A(n9524), .ZN(n9649) );
  INV_X1 U10378 ( .A(n9529), .ZN(n9681) );
  NAND3_X1 U10379 ( .A1(n9576), .A2(n9575), .A3(n9572), .ZN(n9584) );
  AND2_X1 U10380 ( .A1(n9922), .A2(n9530), .ZN(n9543) );
  NAND2_X1 U10381 ( .A1(n9547), .A2(n9531), .ZN(n9532) );
  AND4_X1 U10382 ( .A1(n9553), .A2(n9534), .A3(n9533), .A4(n9532), .ZN(n9535)
         );
  NAND2_X1 U10383 ( .A1(n9554), .A2(n9535), .ZN(n9544) );
  NAND2_X1 U10384 ( .A1(n9537), .A2(n9536), .ZN(n9538) );
  NOR2_X1 U10385 ( .A1(n9544), .A2(n9538), .ZN(n9539) );
  AND4_X1 U10386 ( .A1(n9567), .A2(n9543), .A3(n9539), .A4(n9562), .ZN(n9540)
         );
  NAND2_X1 U10387 ( .A1(n9571), .A2(n9540), .ZN(n9541) );
  NOR2_X1 U10388 ( .A1(n9584), .A2(n9541), .ZN(n9628) );
  NAND2_X1 U10389 ( .A1(n9628), .A2(n9542), .ZN(n9587) );
  INV_X1 U10390 ( .A(n9543), .ZN(n9561) );
  INV_X1 U10391 ( .A(n9544), .ZN(n9549) );
  NAND3_X1 U10392 ( .A1(n9547), .A2(n9546), .A3(n9545), .ZN(n9548) );
  NAND2_X1 U10393 ( .A1(n9549), .A2(n9548), .ZN(n9557) );
  NAND2_X1 U10394 ( .A1(n9551), .A2(n9550), .ZN(n9552) );
  NAND3_X1 U10395 ( .A1(n9554), .A2(n9553), .A3(n9552), .ZN(n9555) );
  AND4_X1 U10396 ( .A1(n9558), .A2(n9557), .A3(n9556), .A4(n9555), .ZN(n9560)
         );
  OAI21_X1 U10397 ( .B1(n9561), .B2(n9560), .A(n9559), .ZN(n9563) );
  NAND2_X1 U10398 ( .A1(n9563), .A2(n9562), .ZN(n9565) );
  NAND2_X1 U10399 ( .A1(n9565), .A2(n9564), .ZN(n9566) );
  NAND3_X1 U10400 ( .A1(n9571), .A2(n9567), .A3(n9566), .ZN(n9583) );
  NAND2_X1 U10401 ( .A1(n9569), .A2(n9568), .ZN(n9570) );
  NAND3_X1 U10402 ( .A1(n9572), .A2(n9571), .A3(n9570), .ZN(n9574) );
  NAND2_X1 U10403 ( .A1(n9574), .A2(n9573), .ZN(n9577) );
  OAI211_X1 U10404 ( .C1(n9578), .C2(n9577), .A(n9576), .B(n9575), .ZN(n9580)
         );
  AND2_X1 U10405 ( .A1(n9580), .A2(n9579), .ZN(n9582) );
  OAI211_X1 U10406 ( .C1(n9584), .C2(n9583), .A(n9582), .B(n9581), .ZN(n9585)
         );
  INV_X1 U10407 ( .A(n9585), .ZN(n9586) );
  AND2_X1 U10408 ( .A1(n9587), .A2(n9586), .ZN(n9630) );
  INV_X1 U10409 ( .A(n9630), .ZN(n9605) );
  INV_X1 U10410 ( .A(n9588), .ZN(n9595) );
  INV_X1 U10411 ( .A(n9589), .ZN(n9590) );
  OAI211_X1 U10412 ( .C1(n9592), .C2(n10408), .A(n9591), .B(n9590), .ZN(n9593)
         );
  NAND4_X1 U10413 ( .A1(n9595), .A2(n9596), .A3(n9594), .A4(n9593), .ZN(n9599)
         );
  NAND3_X1 U10414 ( .A1(n9596), .A2(n10420), .A3(n10392), .ZN(n9597) );
  NAND4_X1 U10415 ( .A1(n9599), .A2(n9623), .A3(n9598), .A4(n9597), .ZN(n9600)
         );
  NAND3_X1 U10416 ( .A1(n9600), .A2(n9627), .A3(n5370), .ZN(n9602) );
  INV_X1 U10417 ( .A(n9628), .ZN(n9601) );
  AOI21_X1 U10418 ( .B1(n9603), .B2(n9602), .A(n9601), .ZN(n9604) );
  OAI21_X1 U10419 ( .B1(n9605), .B2(n9604), .A(n9633), .ZN(n9608) );
  NAND2_X1 U10420 ( .A1(n9607), .A2(n9606), .ZN(n9637) );
  AOI21_X1 U10421 ( .B1(n9608), .B2(n9631), .A(n9637), .ZN(n9612) );
  AND2_X1 U10422 ( .A1(n9610), .A2(n9609), .ZN(n9635) );
  INV_X1 U10423 ( .A(n9635), .ZN(n9611) );
  NOR3_X1 U10424 ( .A1(n9754), .A2(n9612), .A3(n9611), .ZN(n9617) );
  NAND2_X1 U10425 ( .A1(n9636), .A2(n9613), .ZN(n9614) );
  NAND3_X1 U10426 ( .A1(n9616), .A2(n9615), .A3(n9614), .ZN(n9641) );
  NOR2_X1 U10427 ( .A1(n9617), .A2(n9641), .ZN(n9619) );
  NAND2_X1 U10428 ( .A1(n9742), .A2(n9618), .ZN(n9680) );
  OAI211_X1 U10429 ( .C1(n9619), .C2(n9646), .A(n9643), .B(n9680), .ZN(n9620)
         );
  NAND3_X1 U10430 ( .A1(n9683), .A2(n9681), .A3(n9620), .ZN(n9621) );
  NAND2_X1 U10431 ( .A1(n9621), .A2(n9684), .ZN(n9694) );
  AOI21_X1 U10432 ( .B1(n9694), .B2(n10411), .A(n9622), .ZN(n9692) );
  NAND3_X1 U10433 ( .A1(n9625), .A2(n9624), .A3(n9623), .ZN(n9626) );
  NAND3_X1 U10434 ( .A1(n9628), .A2(n9627), .A3(n9626), .ZN(n9629) );
  NAND2_X1 U10435 ( .A1(n9630), .A2(n9629), .ZN(n9634) );
  INV_X1 U10436 ( .A(n9631), .ZN(n9632) );
  AOI21_X1 U10437 ( .B1(n9634), .B2(n9633), .A(n9632), .ZN(n9638) );
  OAI211_X1 U10438 ( .C1(n9638), .C2(n9637), .A(n9636), .B(n9635), .ZN(n9639)
         );
  INV_X1 U10439 ( .A(n9639), .ZN(n9640) );
  NOR2_X1 U10440 ( .A1(n9641), .A2(n9640), .ZN(n9645) );
  INV_X1 U10441 ( .A(n9642), .ZN(n9644) );
  OAI211_X1 U10442 ( .C1(n9646), .C2(n9645), .A(n9644), .B(n9643), .ZN(n9648)
         );
  AOI211_X1 U10443 ( .C1(n9649), .C2(n9648), .A(n9647), .B(n9685), .ZN(n9687)
         );
  INV_X1 U10444 ( .A(n9651), .ZN(n9654) );
  NAND4_X1 U10445 ( .A1(n9655), .A2(n9654), .A3(n9653), .A4(n9652), .ZN(n9657)
         );
  NOR2_X1 U10446 ( .A1(n9657), .A2(n9656), .ZN(n9663) );
  INV_X1 U10447 ( .A(n9658), .ZN(n9662) );
  AND2_X1 U10448 ( .A1(n9659), .A2(n10395), .ZN(n9660) );
  NAND4_X1 U10449 ( .A1(n9663), .A2(n9662), .A3(n9661), .A4(n9660), .ZN(n9665)
         );
  NOR2_X1 U10450 ( .A1(n9665), .A2(n9664), .ZN(n9666) );
  NAND3_X1 U10451 ( .A1(n9668), .A2(n9667), .A3(n9666), .ZN(n9669) );
  NOR4_X1 U10452 ( .A1(n9973), .A2(n9671), .A3(n9670), .A4(n9669), .ZN(n9672)
         );
  NAND4_X1 U10453 ( .A1(n9673), .A2(n5151), .A3(n9950), .A4(n9672), .ZN(n9674)
         );
  NOR2_X1 U10454 ( .A1(n9889), .A2(n9674), .ZN(n9675) );
  AND4_X1 U10455 ( .A1(n9850), .A2(n9882), .A3(n9869), .A4(n9675), .ZN(n9676)
         );
  AND4_X1 U10456 ( .A1(n9805), .A2(n9841), .A3(n9823), .A4(n9676), .ZN(n9677)
         );
  AND4_X1 U10457 ( .A1(n9678), .A2(n9796), .A3(n9770), .A4(n9677), .ZN(n9679)
         );
  AND4_X1 U10458 ( .A1(n6190), .A2(n9680), .A3(n9748), .A4(n9679), .ZN(n9682)
         );
  NAND4_X1 U10459 ( .A1(n9684), .A2(n9683), .A3(n9682), .A4(n9681), .ZN(n9686)
         );
  AND2_X1 U10460 ( .A1(n9686), .A2(n9685), .ZN(n9688) );
  INV_X1 U10461 ( .A(n9688), .ZN(n9690) );
  NOR2_X1 U10462 ( .A1(n9690), .A2(n9689), .ZN(n9691) );
  OAI21_X1 U10463 ( .B1(n9694), .B2(n9693), .A(n9697), .ZN(n9701) );
  NOR4_X1 U10464 ( .A1(n10242), .A2(n6130), .A3(n9696), .A4(n9695), .ZN(n9700)
         );
  INV_X1 U10465 ( .A(n9697), .ZN(n9698) );
  OAI21_X1 U10466 ( .B1(n9441), .B2(n9698), .A(P1_B_REG_SCAN_IN), .ZN(n9699)
         );
  MUX2_X1 U10467 ( .A(n9702), .B(P1_DATAO_REG_31__SCAN_IN), .S(n9719), .Z(
        P1_U3586) );
  INV_X1 U10468 ( .A(n9703), .ZN(n9750) );
  MUX2_X1 U10469 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9750), .S(P1_U4006), .Z(
        P1_U3583) );
  MUX2_X1 U10470 ( .A(n9704), .B(P1_DATAO_REG_27__SCAN_IN), .S(n9719), .Z(
        P1_U3582) );
  MUX2_X1 U10471 ( .A(n9785), .B(P1_DATAO_REG_26__SCAN_IN), .S(n9719), .Z(
        P1_U3581) );
  MUX2_X1 U10472 ( .A(n9806), .B(P1_DATAO_REG_25__SCAN_IN), .S(n9719), .Z(
        P1_U3580) );
  MUX2_X1 U10473 ( .A(n9824), .B(P1_DATAO_REG_24__SCAN_IN), .S(n9719), .Z(
        P1_U3579) );
  MUX2_X1 U10474 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9831), .S(P1_U4006), .Z(
        P1_U3578) );
  MUX2_X1 U10475 ( .A(n9851), .B(P1_DATAO_REG_22__SCAN_IN), .S(n9719), .Z(
        P1_U3577) );
  MUX2_X1 U10476 ( .A(n9870), .B(P1_DATAO_REG_21__SCAN_IN), .S(n9719), .Z(
        P1_U3576) );
  MUX2_X1 U10477 ( .A(n9883), .B(P1_DATAO_REG_20__SCAN_IN), .S(n9719), .Z(
        P1_U3575) );
  MUX2_X1 U10478 ( .A(n9900), .B(P1_DATAO_REG_19__SCAN_IN), .S(n9719), .Z(
        P1_U3574) );
  MUX2_X1 U10479 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9884), .S(P1_U4006), .Z(
        P1_U3573) );
  MUX2_X1 U10480 ( .A(n9899), .B(P1_DATAO_REG_17__SCAN_IN), .S(n9719), .Z(
        P1_U3572) );
  MUX2_X1 U10481 ( .A(n9705), .B(P1_DATAO_REG_16__SCAN_IN), .S(n9719), .Z(
        P1_U3571) );
  MUX2_X1 U10482 ( .A(n9706), .B(P1_DATAO_REG_15__SCAN_IN), .S(n9719), .Z(
        P1_U3570) );
  MUX2_X1 U10483 ( .A(n9707), .B(P1_DATAO_REG_14__SCAN_IN), .S(n9719), .Z(
        P1_U3569) );
  MUX2_X1 U10484 ( .A(n9708), .B(P1_DATAO_REG_13__SCAN_IN), .S(n9719), .Z(
        P1_U3568) );
  MUX2_X1 U10485 ( .A(n9709), .B(P1_DATAO_REG_12__SCAN_IN), .S(n9719), .Z(
        P1_U3567) );
  MUX2_X1 U10486 ( .A(n9710), .B(P1_DATAO_REG_11__SCAN_IN), .S(n9719), .Z(
        P1_U3566) );
  MUX2_X1 U10487 ( .A(n9711), .B(P1_DATAO_REG_10__SCAN_IN), .S(n9719), .Z(
        P1_U3565) );
  MUX2_X1 U10488 ( .A(n9712), .B(P1_DATAO_REG_9__SCAN_IN), .S(n9719), .Z(
        P1_U3564) );
  MUX2_X1 U10489 ( .A(n9713), .B(P1_DATAO_REG_7__SCAN_IN), .S(n9719), .Z(
        P1_U3562) );
  MUX2_X1 U10490 ( .A(n9714), .B(P1_DATAO_REG_6__SCAN_IN), .S(n9719), .Z(
        P1_U3561) );
  MUX2_X1 U10491 ( .A(n9715), .B(P1_DATAO_REG_5__SCAN_IN), .S(n9719), .Z(
        P1_U3560) );
  MUX2_X1 U10492 ( .A(n9716), .B(P1_DATAO_REG_4__SCAN_IN), .S(n9719), .Z(
        P1_U3559) );
  MUX2_X1 U10493 ( .A(n9717), .B(P1_DATAO_REG_3__SCAN_IN), .S(n9719), .Z(
        P1_U3558) );
  MUX2_X1 U10494 ( .A(n10392), .B(P1_DATAO_REG_2__SCAN_IN), .S(n9719), .Z(
        P1_U3557) );
  MUX2_X1 U10495 ( .A(n9718), .B(P1_DATAO_REG_1__SCAN_IN), .S(n9719), .Z(
        P1_U3556) );
  MUX2_X1 U10496 ( .A(n6205), .B(P1_DATAO_REG_0__SCAN_IN), .S(n9719), .Z(
        P1_U3555) );
  AOI21_X1 U10497 ( .B1(P1_REG1_REG_17__SCAN_IN), .B2(n9727), .A(n9720), .ZN(
        n10307) );
  INV_X1 U10498 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9722) );
  AOI22_X1 U10499 ( .A1(n10304), .A2(P1_REG1_REG_18__SCAN_IN), .B1(n9722), 
        .B2(n9721), .ZN(n10306) );
  NAND2_X1 U10500 ( .A1(n10307), .A2(n10306), .ZN(n10305) );
  OAI21_X1 U10501 ( .B1(P1_REG1_REG_18__SCAN_IN), .B2(n10304), .A(n10305), 
        .ZN(n9724) );
  XNOR2_X1 U10502 ( .A(n10411), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n9723) );
  XNOR2_X1 U10503 ( .A(n9724), .B(n9723), .ZN(n9740) );
  INV_X1 U10504 ( .A(n9725), .ZN(n9726) );
  AOI21_X1 U10505 ( .B1(n9727), .B2(P1_REG2_REG_17__SCAN_IN), .A(n9726), .ZN(
        n10301) );
  INV_X1 U10506 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9728) );
  OR2_X1 U10507 ( .A1(n10304), .A2(n9728), .ZN(n9730) );
  NAND2_X1 U10508 ( .A1(n10304), .A2(n9728), .ZN(n9729) );
  AND2_X1 U10509 ( .A1(n9730), .A2(n9729), .ZN(n10300) );
  NOR2_X1 U10510 ( .A1(n10301), .A2(n10300), .ZN(n10299) );
  AOI21_X1 U10511 ( .B1(n10304), .B2(P1_REG2_REG_18__SCAN_IN), .A(n10299), 
        .ZN(n9733) );
  INV_X1 U10512 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n9731) );
  MUX2_X1 U10513 ( .A(n9731), .B(P1_REG2_REG_19__SCAN_IN), .S(n10411), .Z(
        n9732) );
  XNOR2_X1 U10514 ( .A(n9733), .B(n9732), .ZN(n9734) );
  OAI22_X1 U10515 ( .A1(n9736), .A2(n9735), .B1(n10298), .B2(n9734), .ZN(n9737) );
  AOI211_X1 U10516 ( .C1(n10411), .C2(n10312), .A(n9738), .B(n9737), .ZN(n9739) );
  OAI21_X1 U10517 ( .B1(n9740), .B2(n10269), .A(n9739), .ZN(P1_U3260) );
  INV_X1 U10518 ( .A(n9741), .ZN(n9743) );
  NAND2_X1 U10519 ( .A1(n9743), .A2(n9742), .ZN(n9990) );
  NAND3_X1 U10520 ( .A1(n9990), .A2(n9989), .A3(n10368), .ZN(n9746) );
  AOI21_X1 U10521 ( .B1(n10419), .B2(P1_REG2_REG_30__SCAN_IN), .A(n9744), .ZN(
        n9745) );
  OAI211_X1 U10522 ( .C1(n9993), .C2(n9969), .A(n9746), .B(n9745), .ZN(
        P1_U3262) );
  NAND2_X1 U10523 ( .A1(n9766), .A2(n9747), .ZN(n9749) );
  XNOR2_X1 U10524 ( .A(n9755), .B(n9754), .ZN(n10002) );
  NAND2_X1 U10525 ( .A1(n10371), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n9756) );
  OAI21_X1 U10526 ( .B1(n10376), .B2(n9757), .A(n9756), .ZN(n9758) );
  AOI21_X1 U10527 ( .B1(n9998), .B2(n10367), .A(n9758), .ZN(n9763) );
  NAND2_X1 U10528 ( .A1(n9998), .A2(n9775), .ZN(n9760) );
  AND2_X1 U10529 ( .A1(n9761), .A2(n9760), .ZN(n9999) );
  NAND2_X1 U10530 ( .A1(n9999), .A2(n10368), .ZN(n9762) );
  OAI211_X1 U10531 ( .C1(n10002), .C2(n9985), .A(n9763), .B(n9762), .ZN(n9764)
         );
  INV_X1 U10532 ( .A(n9764), .ZN(n9765) );
  OAI21_X1 U10533 ( .B1(n10001), .B2(n10371), .A(n9765), .ZN(P1_U3264) );
  OAI21_X1 U10534 ( .B1(n9770), .B2(n9767), .A(n9766), .ZN(n9774) );
  OAI22_X1 U10535 ( .A1(n9769), .A2(n9977), .B1(n9768), .B2(n9975), .ZN(n9773)
         );
  XNOR2_X1 U10536 ( .A(n9771), .B(n9770), .ZN(n10007) );
  NOR2_X1 U10537 ( .A1(n10007), .A2(n10401), .ZN(n9772) );
  AOI21_X1 U10538 ( .B1(n10003), .B2(n9789), .A(n9759), .ZN(n10004) );
  INV_X1 U10539 ( .A(n10003), .ZN(n9778) );
  AOI22_X1 U10540 ( .A1(n10371), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n9776), 
        .B2(n10409), .ZN(n9777) );
  OAI21_X1 U10541 ( .B1(n9778), .B2(n9969), .A(n9777), .ZN(n9781) );
  NOR2_X1 U10542 ( .A1(n10007), .A2(n9779), .ZN(n9780) );
  AOI211_X1 U10543 ( .C1(n10004), .C2(n10368), .A(n9781), .B(n9780), .ZN(n9782) );
  OAI21_X1 U10544 ( .B1(n10006), .B2(n10419), .A(n9782), .ZN(P1_U3265) );
  OAI21_X1 U10545 ( .B1(n9796), .B2(n9784), .A(n9783), .ZN(n9786) );
  AOI222_X1 U10546 ( .A1(n10397), .A2(n9786), .B1(n9785), .B2(n10391), .C1(
        n9824), .C2(n10393), .ZN(n10011) );
  INV_X1 U10547 ( .A(n9808), .ZN(n9787) );
  NAND2_X1 U10548 ( .A1(n9787), .A2(n10008), .ZN(n9788) );
  AND2_X1 U10549 ( .A1(n9789), .A2(n9788), .ZN(n10009) );
  AOI22_X1 U10550 ( .A1(n10419), .A2(P1_REG2_REG_25__SCAN_IN), .B1(n9790), 
        .B2(n10409), .ZN(n9791) );
  OAI21_X1 U10551 ( .B1(n9792), .B2(n9969), .A(n9791), .ZN(n9798) );
  INV_X1 U10552 ( .A(n9793), .ZN(n9794) );
  AOI21_X1 U10553 ( .B1(n9796), .B2(n9795), .A(n9794), .ZN(n10012) );
  NOR2_X1 U10554 ( .A1(n10012), .A2(n9985), .ZN(n9797) );
  AOI211_X1 U10555 ( .C1(n10009), .C2(n10368), .A(n9798), .B(n9797), .ZN(n9799) );
  OAI21_X1 U10556 ( .B1(n10011), .B2(n10371), .A(n9799), .ZN(P1_U3266) );
  INV_X1 U10557 ( .A(n9805), .ZN(n9801) );
  OAI21_X1 U10558 ( .B1(n9802), .B2(n9801), .A(n9800), .ZN(n10017) );
  OAI21_X1 U10559 ( .B1(n9805), .B2(n9804), .A(n9803), .ZN(n9807) );
  AOI222_X1 U10560 ( .A1(n10397), .A2(n9807), .B1(n9806), .B2(n10391), .C1(
        n9831), .C2(n10393), .ZN(n10016) );
  AOI211_X1 U10561 ( .C1(n10014), .C2(n9816), .A(n10522), .B(n9808), .ZN(
        n10013) );
  AOI22_X1 U10562 ( .A1(n10013), .A2(n9856), .B1(n10409), .B2(n9809), .ZN(
        n9810) );
  AOI21_X1 U10563 ( .B1(n10016), .B2(n9810), .A(n10371), .ZN(n9811) );
  INV_X1 U10564 ( .A(n9811), .ZN(n9813) );
  AOI22_X1 U10565 ( .A1(n10014), .A2(n10367), .B1(n10419), .B2(
        P1_REG2_REG_24__SCAN_IN), .ZN(n9812) );
  OAI211_X1 U10566 ( .C1(n10017), .C2(n9985), .A(n9813), .B(n9812), .ZN(
        P1_U3267) );
  XNOR2_X1 U10567 ( .A(n9814), .B(n9823), .ZN(n10022) );
  OR2_X1 U10568 ( .A1(n9820), .A2(n9833), .ZN(n9815) );
  AND3_X1 U10569 ( .A1(n9816), .A2(n9815), .A3(n10386), .ZN(n10018) );
  NOR2_X1 U10570 ( .A1(n10376), .A2(n9817), .ZN(n9818) );
  AOI21_X1 U10571 ( .B1(n10419), .B2(P1_REG2_REG_23__SCAN_IN), .A(n9818), .ZN(
        n9819) );
  OAI21_X1 U10572 ( .B1(n9820), .B2(n9969), .A(n9819), .ZN(n9827) );
  OAI21_X1 U10573 ( .B1(n9823), .B2(n9822), .A(n9821), .ZN(n9825) );
  AOI222_X1 U10574 ( .A1(n10397), .A2(n9825), .B1(n9824), .B2(n10391), .C1(
        n9851), .C2(n10393), .ZN(n10021) );
  NOR2_X1 U10575 ( .A1(n10021), .A2(n10371), .ZN(n9826) );
  AOI211_X1 U10576 ( .C1(n10018), .C2(n9983), .A(n9827), .B(n9826), .ZN(n9828)
         );
  OAI21_X1 U10577 ( .B1(n10022), .B2(n9985), .A(n9828), .ZN(P1_U3268) );
  OAI21_X1 U10578 ( .B1(n9841), .B2(n9830), .A(n9829), .ZN(n9832) );
  AOI222_X1 U10579 ( .A1(n10397), .A2(n9832), .B1(n9870), .B2(n10393), .C1(
        n9831), .C2(n10391), .ZN(n10027) );
  AND2_X1 U10580 ( .A1(n9835), .A2(n9853), .ZN(n9834) );
  OR2_X1 U10581 ( .A1(n9834), .A2(n9833), .ZN(n10024) );
  INV_X1 U10582 ( .A(n10024), .ZN(n9844) );
  INV_X1 U10583 ( .A(n9835), .ZN(n10023) );
  AOI22_X1 U10584 ( .A1(n10371), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n9836), 
        .B2(n10409), .ZN(n9837) );
  OAI21_X1 U10585 ( .B1(n10023), .B2(n9969), .A(n9837), .ZN(n9843) );
  INV_X1 U10586 ( .A(n9838), .ZN(n9839) );
  AOI21_X1 U10587 ( .B1(n9841), .B2(n9840), .A(n9839), .ZN(n10028) );
  NOR2_X1 U10588 ( .A1(n10028), .A2(n9985), .ZN(n9842) );
  AOI211_X1 U10589 ( .C1(n9844), .C2(n10368), .A(n9843), .B(n9842), .ZN(n9845)
         );
  OAI21_X1 U10590 ( .B1(n10027), .B2(n10371), .A(n9845), .ZN(P1_U3269) );
  XNOR2_X1 U10591 ( .A(n9847), .B(n9846), .ZN(n10033) );
  OAI21_X1 U10592 ( .B1(n9850), .B2(n9849), .A(n9848), .ZN(n9852) );
  AOI222_X1 U10593 ( .A1(n10397), .A2(n9852), .B1(n9851), .B2(n10391), .C1(
        n9883), .C2(n10393), .ZN(n10032) );
  INV_X1 U10594 ( .A(n9853), .ZN(n9854) );
  AOI211_X1 U10595 ( .C1(n10030), .C2(n9862), .A(n10522), .B(n9854), .ZN(
        n10029) );
  AOI22_X1 U10596 ( .A1(n10029), .A2(n9856), .B1(n9855), .B2(n10409), .ZN(
        n9857) );
  AOI21_X1 U10597 ( .B1(n10032), .B2(n9857), .A(n10371), .ZN(n9858) );
  INV_X1 U10598 ( .A(n9858), .ZN(n9860) );
  AOI22_X1 U10599 ( .A1(n10030), .A2(n10367), .B1(n10419), .B2(
        P1_REG2_REG_21__SCAN_IN), .ZN(n9859) );
  OAI211_X1 U10600 ( .C1(n10033), .C2(n9985), .A(n9860), .B(n9859), .ZN(
        P1_U3270) );
  XNOR2_X1 U10601 ( .A(n9861), .B(n5133), .ZN(n10038) );
  INV_X1 U10602 ( .A(n9862), .ZN(n9863) );
  AOI211_X1 U10603 ( .C1(n10035), .C2(n4980), .A(n10522), .B(n9863), .ZN(
        n10034) );
  AOI22_X1 U10604 ( .A1(n10371), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9864), 
        .B2(n10409), .ZN(n9865) );
  OAI21_X1 U10605 ( .B1(n9866), .B2(n9969), .A(n9865), .ZN(n9873) );
  OAI21_X1 U10606 ( .B1(n9869), .B2(n9868), .A(n9867), .ZN(n9871) );
  AOI222_X1 U10607 ( .A1(n10397), .A2(n9871), .B1(n9870), .B2(n10391), .C1(
        n9900), .C2(n10393), .ZN(n10037) );
  NOR2_X1 U10608 ( .A1(n10037), .A2(n10371), .ZN(n9872) );
  AOI211_X1 U10609 ( .C1(n10034), .C2(n9983), .A(n9873), .B(n9872), .ZN(n9874)
         );
  OAI21_X1 U10610 ( .B1(n9985), .B2(n10038), .A(n9874), .ZN(P1_U3271) );
  XNOR2_X1 U10611 ( .A(n9876), .B(n9875), .ZN(n10043) );
  AOI21_X1 U10612 ( .B1(n10039), .B2(n9891), .A(n9877), .ZN(n10040) );
  AOI22_X1 U10613 ( .A1(n10371), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9878), 
        .B2(n10409), .ZN(n9879) );
  OAI21_X1 U10614 ( .B1(n4979), .B2(n9969), .A(n9879), .ZN(n9887) );
  OAI21_X1 U10615 ( .B1(n9882), .B2(n9881), .A(n4935), .ZN(n9885) );
  AOI222_X1 U10616 ( .A1(n10397), .A2(n9885), .B1(n9884), .B2(n10393), .C1(
        n9883), .C2(n10391), .ZN(n10042) );
  NOR2_X1 U10617 ( .A1(n10042), .A2(n10419), .ZN(n9886) );
  AOI211_X1 U10618 ( .C1(n10040), .C2(n10368), .A(n9887), .B(n9886), .ZN(n9888) );
  OAI21_X1 U10619 ( .B1(n9985), .B2(n10043), .A(n9888), .ZN(P1_U3272) );
  XNOR2_X1 U10620 ( .A(n9890), .B(n9889), .ZN(n10048) );
  INV_X1 U10621 ( .A(n9896), .ZN(n10044) );
  INV_X1 U10622 ( .A(n9914), .ZN(n9893) );
  INV_X1 U10623 ( .A(n9891), .ZN(n9892) );
  AOI21_X1 U10624 ( .B1(n10044), .B2(n9893), .A(n9892), .ZN(n10045) );
  AOI22_X1 U10625 ( .A1(n10371), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9894), 
        .B2(n10409), .ZN(n9895) );
  OAI21_X1 U10626 ( .B1(n9896), .B2(n9969), .A(n9895), .ZN(n9903) );
  OAI21_X1 U10627 ( .B1(n5238), .B2(n9898), .A(n9897), .ZN(n9901) );
  AOI222_X1 U10628 ( .A1(n10397), .A2(n9901), .B1(n9900), .B2(n10391), .C1(
        n9899), .C2(n10393), .ZN(n10047) );
  NOR2_X1 U10629 ( .A1(n10047), .A2(n10371), .ZN(n9902) );
  AOI211_X1 U10630 ( .C1(n10045), .C2(n10368), .A(n9903), .B(n9902), .ZN(n9904) );
  OAI21_X1 U10631 ( .B1(n9985), .B2(n10048), .A(n9904), .ZN(P1_U3273) );
  NOR2_X1 U10632 ( .A1(n9923), .A2(n9905), .ZN(n9906) );
  XNOR2_X1 U10633 ( .A(n9906), .B(n9908), .ZN(n9912) );
  OAI22_X1 U10634 ( .A1(n9947), .A2(n9977), .B1(n9907), .B2(n9975), .ZN(n9911)
         );
  XNOR2_X1 U10635 ( .A(n9909), .B(n9908), .ZN(n10055) );
  NOR2_X1 U10636 ( .A1(n10055), .A2(n10401), .ZN(n9910) );
  AOI211_X1 U10637 ( .C1(n9912), .C2(n10397), .A(n9911), .B(n9910), .ZN(n10054) );
  INV_X1 U10638 ( .A(n10055), .ZN(n9920) );
  AND2_X1 U10639 ( .A1(n10049), .A2(n9936), .ZN(n9913) );
  OR2_X1 U10640 ( .A1(n9914), .A2(n9913), .ZN(n10051) );
  AOI22_X1 U10641 ( .A1(n10371), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9915), 
        .B2(n10409), .ZN(n9917) );
  NAND2_X1 U10642 ( .A1(n10049), .A2(n10367), .ZN(n9916) );
  OAI211_X1 U10643 ( .C1(n10051), .C2(n9918), .A(n9917), .B(n9916), .ZN(n9919)
         );
  AOI21_X1 U10644 ( .B1(n9920), .B2(n10415), .A(n9919), .ZN(n9921) );
  OAI21_X1 U10645 ( .B1(n10054), .B2(n10419), .A(n9921), .ZN(P1_U3274) );
  NOR2_X1 U10646 ( .A1(n5151), .A2(n5148), .ZN(n9925) );
  AOI21_X1 U10647 ( .B1(n9925), .B2(n9924), .A(n9923), .ZN(n9926) );
  OAI222_X1 U10648 ( .A1(n9977), .A2(n9976), .B1(n9975), .B2(n9927), .C1(n9972), .C2(n9926), .ZN(n10056) );
  OAI21_X1 U10649 ( .B1(n9930), .B2(n9929), .A(n9928), .ZN(n10060) );
  NAND2_X1 U10650 ( .A1(n10419), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n9931) );
  OAI21_X1 U10651 ( .B1(n10376), .B2(n9932), .A(n9931), .ZN(n9933) );
  AOI21_X1 U10652 ( .B1(n10058), .B2(n10367), .A(n9933), .ZN(n9938) );
  OR2_X1 U10653 ( .A1(n9954), .A2(n9934), .ZN(n9935) );
  AND3_X1 U10654 ( .A1(n9936), .A2(n9935), .A3(n10386), .ZN(n10057) );
  NAND2_X1 U10655 ( .A1(n10057), .A2(n9983), .ZN(n9937) );
  OAI211_X1 U10656 ( .C1(n10060), .C2(n9985), .A(n9938), .B(n9937), .ZN(n9939)
         );
  AOI21_X1 U10657 ( .B1(n10056), .B2(n9940), .A(n9939), .ZN(n9941) );
  INV_X1 U10658 ( .A(n9941), .ZN(P1_U3275) );
  NAND2_X1 U10659 ( .A1(n9943), .A2(n9942), .ZN(n9946) );
  INV_X1 U10660 ( .A(n9944), .ZN(n9945) );
  AOI21_X1 U10661 ( .B1(n9950), .B2(n9946), .A(n9945), .ZN(n10061) );
  OAI22_X1 U10662 ( .A1(n9948), .A2(n9977), .B1(n9947), .B2(n9975), .ZN(n9953)
         );
  XOR2_X1 U10663 ( .A(n9950), .B(n9949), .Z(n9951) );
  NOR2_X1 U10664 ( .A1(n9951), .A2(n9972), .ZN(n9952) );
  AOI211_X1 U10665 ( .C1(n6266), .C2(n10061), .A(n9953), .B(n9952), .ZN(n10065) );
  INV_X1 U10666 ( .A(n9966), .ZN(n9955) );
  AOI21_X1 U10667 ( .B1(n10062), .B2(n9955), .A(n9954), .ZN(n10063) );
  NAND2_X1 U10668 ( .A1(n10063), .A2(n10368), .ZN(n9958) );
  AOI22_X1 U10669 ( .A1(n10419), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n9956), 
        .B2(n10409), .ZN(n9957) );
  OAI211_X1 U10670 ( .C1(n9959), .C2(n9969), .A(n9958), .B(n9957), .ZN(n9960)
         );
  AOI21_X1 U10671 ( .B1(n10061), .B2(n10415), .A(n9960), .ZN(n9961) );
  OAI21_X1 U10672 ( .B1(n10065), .B2(n10371), .A(n9961), .ZN(P1_U3276) );
  NAND2_X1 U10673 ( .A1(n9963), .A2(n9962), .ZN(n9965) );
  XNOR2_X1 U10674 ( .A(n9965), .B(n9964), .ZN(n10071) );
  AOI211_X1 U10675 ( .C1(n10068), .C2(n4913), .A(n10522), .B(n9966), .ZN(
        n10067) );
  INV_X1 U10676 ( .A(n10068), .ZN(n9970) );
  AOI22_X1 U10677 ( .A1(n10371), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n9967), 
        .B2(n10409), .ZN(n9968) );
  OAI21_X1 U10678 ( .B1(n9970), .B2(n9969), .A(n9968), .ZN(n9982) );
  AOI211_X1 U10679 ( .C1(n9974), .C2(n9973), .A(n9972), .B(n9971), .ZN(n9980)
         );
  OAI22_X1 U10680 ( .A1(n9978), .A2(n9977), .B1(n9976), .B2(n9975), .ZN(n9979)
         );
  NOR2_X1 U10681 ( .A1(n9980), .A2(n9979), .ZN(n10070) );
  NOR2_X1 U10682 ( .A1(n10070), .A2(n10371), .ZN(n9981) );
  AOI211_X1 U10683 ( .C1(n9983), .C2(n10067), .A(n9982), .B(n9981), .ZN(n9984)
         );
  OAI21_X1 U10684 ( .B1(n10071), .B2(n9985), .A(n9984), .ZN(P1_U3277) );
  NAND2_X1 U10685 ( .A1(n9986), .A2(n10502), .ZN(n9987) );
  OAI211_X1 U10686 ( .C1(n9988), .C2(n10522), .A(n9987), .B(n9991), .ZN(n10084) );
  MUX2_X1 U10687 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n10084), .S(n10531), .Z(
        P1_U3554) );
  NAND3_X1 U10688 ( .A1(n9990), .A2(n10386), .A3(n9989), .ZN(n9992) );
  OAI211_X1 U10689 ( .C1(n9993), .C2(n10520), .A(n9992), .B(n9991), .ZN(n10085) );
  MUX2_X1 U10690 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n10085), .S(n10531), .Z(
        P1_U3553) );
  MUX2_X1 U10691 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9997), .S(n10531), .Z(
        P1_U3551) );
  AOI22_X1 U10692 ( .A1(n9999), .A2(n10386), .B1(n10502), .B2(n9998), .ZN(
        n10000) );
  OAI211_X1 U10693 ( .C1(n10436), .C2(n10002), .A(n10001), .B(n10000), .ZN(
        n10087) );
  MUX2_X1 U10694 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n10087), .S(n10531), .Z(
        P1_U3550) );
  AOI22_X1 U10695 ( .A1(n10004), .A2(n10386), .B1(n10502), .B2(n10003), .ZN(
        n10005) );
  OAI211_X1 U10696 ( .C1(n10007), .C2(n10504), .A(n10006), .B(n10005), .ZN(
        n10088) );
  MUX2_X1 U10697 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n10088), .S(n10531), .Z(
        P1_U3549) );
  AOI22_X1 U10698 ( .A1(n10009), .A2(n10386), .B1(n10502), .B2(n10008), .ZN(
        n10010) );
  OAI211_X1 U10699 ( .C1(n10436), .C2(n10012), .A(n10011), .B(n10010), .ZN(
        n10089) );
  MUX2_X1 U10700 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n10089), .S(n10531), .Z(
        P1_U3548) );
  AOI21_X1 U10701 ( .B1(n10502), .B2(n10014), .A(n10013), .ZN(n10015) );
  OAI211_X1 U10702 ( .C1(n10436), .C2(n10017), .A(n10016), .B(n10015), .ZN(
        n10090) );
  MUX2_X1 U10703 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n10090), .S(n10531), .Z(
        P1_U3547) );
  AOI21_X1 U10704 ( .B1(n10502), .B2(n10019), .A(n10018), .ZN(n10020) );
  OAI211_X1 U10705 ( .C1(n10436), .C2(n10022), .A(n10021), .B(n10020), .ZN(
        n10091) );
  MUX2_X1 U10706 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n10091), .S(n10531), .Z(
        P1_U3546) );
  OAI22_X1 U10707 ( .A1(n10024), .A2(n10522), .B1(n10023), .B2(n10520), .ZN(
        n10025) );
  INV_X1 U10708 ( .A(n10025), .ZN(n10026) );
  OAI211_X1 U10709 ( .C1(n10436), .C2(n10028), .A(n10027), .B(n10026), .ZN(
        n10092) );
  MUX2_X1 U10710 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n10092), .S(n10531), .Z(
        P1_U3545) );
  AOI21_X1 U10711 ( .B1(n10502), .B2(n10030), .A(n10029), .ZN(n10031) );
  OAI211_X1 U10712 ( .C1(n10436), .C2(n10033), .A(n10032), .B(n10031), .ZN(
        n10093) );
  MUX2_X1 U10713 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n10093), .S(n10531), .Z(
        P1_U3544) );
  AOI21_X1 U10714 ( .B1(n10502), .B2(n10035), .A(n10034), .ZN(n10036) );
  OAI211_X1 U10715 ( .C1(n10436), .C2(n10038), .A(n10037), .B(n10036), .ZN(
        n10094) );
  MUX2_X1 U10716 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n10094), .S(n10531), .Z(
        P1_U3543) );
  AOI22_X1 U10717 ( .A1(n10040), .A2(n10386), .B1(n10502), .B2(n10039), .ZN(
        n10041) );
  OAI211_X1 U10718 ( .C1(n10436), .C2(n10043), .A(n10042), .B(n10041), .ZN(
        n10095) );
  MUX2_X1 U10719 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n10095), .S(n10531), .Z(
        P1_U3542) );
  AOI22_X1 U10720 ( .A1(n10045), .A2(n10386), .B1(n10502), .B2(n10044), .ZN(
        n10046) );
  OAI211_X1 U10721 ( .C1(n10436), .C2(n10048), .A(n10047), .B(n10046), .ZN(
        n10096) );
  MUX2_X1 U10722 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n10096), .S(n10531), .Z(
        P1_U3541) );
  INV_X1 U10723 ( .A(n10049), .ZN(n10050) );
  OAI22_X1 U10724 ( .A1(n10051), .A2(n10522), .B1(n10050), .B2(n10520), .ZN(
        n10052) );
  INV_X1 U10725 ( .A(n10052), .ZN(n10053) );
  OAI211_X1 U10726 ( .C1(n10504), .C2(n10055), .A(n10054), .B(n10053), .ZN(
        n10097) );
  MUX2_X1 U10727 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n10097), .S(n10531), .Z(
        P1_U3540) );
  AOI211_X1 U10728 ( .C1(n10502), .C2(n10058), .A(n10057), .B(n10056), .ZN(
        n10059) );
  OAI21_X1 U10729 ( .B1(n10436), .B2(n10060), .A(n10059), .ZN(n10098) );
  MUX2_X1 U10730 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n10098), .S(n10531), .Z(
        P1_U3539) );
  INV_X1 U10731 ( .A(n10061), .ZN(n10066) );
  AOI22_X1 U10732 ( .A1(n10063), .A2(n10386), .B1(n10502), .B2(n10062), .ZN(
        n10064) );
  OAI211_X1 U10733 ( .C1(n10504), .C2(n10066), .A(n10065), .B(n10064), .ZN(
        n10099) );
  MUX2_X1 U10734 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n10099), .S(n10531), .Z(
        P1_U3538) );
  AOI21_X1 U10735 ( .B1(n10502), .B2(n10068), .A(n10067), .ZN(n10069) );
  OAI211_X1 U10736 ( .C1(n10436), .C2(n10071), .A(n10070), .B(n10069), .ZN(
        n10100) );
  MUX2_X1 U10737 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n10100), .S(n10531), .Z(
        P1_U3537) );
  INV_X1 U10738 ( .A(n10504), .ZN(n10525) );
  NAND2_X1 U10739 ( .A1(n10072), .A2(n10525), .ZN(n10075) );
  AOI22_X1 U10740 ( .A1(n10073), .A2(n10386), .B1(n10502), .B2(n6157), .ZN(
        n10074) );
  NAND2_X1 U10741 ( .A1(n10075), .A2(n10074), .ZN(n10076) );
  MUX2_X1 U10742 ( .A(n10101), .B(P1_REG1_REG_13__SCAN_IN), .S(n10529), .Z(
        P1_U3536) );
  AOI211_X1 U10743 ( .C1(n10502), .C2(n10080), .A(n10079), .B(n10078), .ZN(
        n10081) );
  OAI21_X1 U10744 ( .B1(n10436), .B2(n10082), .A(n10081), .ZN(n10102) );
  MUX2_X1 U10745 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n10102), .S(n10531), .Z(
        P1_U3535) );
  MUX2_X1 U10746 ( .A(n10083), .B(P1_REG1_REG_0__SCAN_IN), .S(n10529), .Z(
        P1_U3523) );
  MUX2_X1 U10747 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n10084), .S(n10535), .Z(
        P1_U3522) );
  MUX2_X1 U10748 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n10085), .S(n10535), .Z(
        P1_U3521) );
  MUX2_X1 U10749 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n10086), .S(n10535), .Z(
        P1_U3520) );
  MUX2_X1 U10750 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n10087), .S(n10535), .Z(
        P1_U3518) );
  MUX2_X1 U10751 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n10088), .S(n10535), .Z(
        P1_U3517) );
  MUX2_X1 U10752 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n10089), .S(n10535), .Z(
        P1_U3516) );
  MUX2_X1 U10753 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n10090), .S(n10535), .Z(
        P1_U3515) );
  MUX2_X1 U10754 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n10091), .S(n10535), .Z(
        P1_U3514) );
  MUX2_X1 U10755 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n10092), .S(n10535), .Z(
        P1_U3513) );
  MUX2_X1 U10756 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n10093), .S(n10535), .Z(
        P1_U3512) );
  MUX2_X1 U10757 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n10094), .S(n10535), .Z(
        P1_U3511) );
  MUX2_X1 U10758 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n10095), .S(n10535), .Z(
        P1_U3510) );
  MUX2_X1 U10759 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n10096), .S(n10535), .Z(
        P1_U3508) );
  MUX2_X1 U10760 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n10097), .S(n10535), .Z(
        P1_U3505) );
  MUX2_X1 U10761 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n10098), .S(n10535), .Z(
        P1_U3502) );
  MUX2_X1 U10762 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n10099), .S(n10535), .Z(
        P1_U3499) );
  MUX2_X1 U10763 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n10100), .S(n10535), .Z(
        P1_U3496) );
  MUX2_X1 U10764 ( .A(n10101), .B(P1_REG0_REG_13__SCAN_IN), .S(n10532), .Z(
        P1_U3493) );
  MUX2_X1 U10765 ( .A(P1_REG0_REG_12__SCAN_IN), .B(n10102), .S(n10535), .Z(
        P1_U3490) );
  MUX2_X1 U10766 ( .A(n10103), .B(P1_D_REG_0__SCAN_IN), .S(n10242), .Z(
        P1_U3440) );
  INV_X1 U10767 ( .A(n10104), .ZN(n10106) );
  NAND4_X1 U10768 ( .A1(n10106), .A2(P1_IR_REG_31__SCAN_IN), .A3(
        P1_STATE_REG_SCAN_IN), .A4(n10105), .ZN(n10109) );
  NAND2_X1 U10769 ( .A1(n10107), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n10108) );
  OAI211_X1 U10770 ( .C1(n10110), .C2(n10113), .A(n10109), .B(n10108), .ZN(
        P1_U3322) );
  OAI222_X1 U10771 ( .A1(n10113), .A2(n10112), .B1(P1_U3084), .B2(n10111), 
        .C1(n10119), .C2(n6184), .ZN(P1_U3324) );
  NAND2_X1 U10772 ( .A1(n10115), .A2(n10114), .ZN(n10117) );
  OAI211_X1 U10773 ( .C1(n10119), .C2(n10118), .A(n10117), .B(n10116), .ZN(
        P1_U3325) );
  MUX2_X1 U10774 ( .A(n10120), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3353) );
  NOR2_X4 U10775 ( .A1(n10121), .A2(n10242), .ZN(n10146) );
  INV_X1 U10776 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n10122) );
  NOR2_X1 U10777 ( .A1(n10146), .A2(n10122), .ZN(P1_U3321) );
  INV_X1 U10778 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n10123) );
  NOR2_X1 U10779 ( .A1(n10146), .A2(n10123), .ZN(P1_U3320) );
  INV_X1 U10780 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n10124) );
  NOR2_X1 U10781 ( .A1(n10146), .A2(n10124), .ZN(P1_U3319) );
  INV_X1 U10782 ( .A(P1_D_REG_5__SCAN_IN), .ZN(n10125) );
  NOR2_X1 U10783 ( .A1(n10146), .A2(n10125), .ZN(P1_U3318) );
  INV_X1 U10784 ( .A(P1_D_REG_6__SCAN_IN), .ZN(n10126) );
  NOR2_X1 U10785 ( .A1(n10146), .A2(n10126), .ZN(P1_U3317) );
  INV_X1 U10786 ( .A(P1_D_REG_7__SCAN_IN), .ZN(n10127) );
  NOR2_X1 U10787 ( .A1(n10146), .A2(n10127), .ZN(P1_U3316) );
  INV_X1 U10788 ( .A(P1_D_REG_8__SCAN_IN), .ZN(n10128) );
  NOR2_X1 U10789 ( .A1(n10146), .A2(n10128), .ZN(P1_U3315) );
  INV_X1 U10790 ( .A(P1_D_REG_9__SCAN_IN), .ZN(n10129) );
  NOR2_X1 U10791 ( .A1(n10146), .A2(n10129), .ZN(P1_U3314) );
  INV_X1 U10792 ( .A(P1_D_REG_10__SCAN_IN), .ZN(n10130) );
  NOR2_X1 U10793 ( .A1(n10146), .A2(n10130), .ZN(P1_U3313) );
  INV_X1 U10794 ( .A(P1_D_REG_11__SCAN_IN), .ZN(n10131) );
  NOR2_X1 U10795 ( .A1(n10146), .A2(n10131), .ZN(P1_U3312) );
  INV_X1 U10796 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n10132) );
  NOR2_X1 U10797 ( .A1(n10146), .A2(n10132), .ZN(P1_U3311) );
  INV_X1 U10798 ( .A(P1_D_REG_13__SCAN_IN), .ZN(n10133) );
  NOR2_X1 U10799 ( .A1(n10146), .A2(n10133), .ZN(P1_U3310) );
  INV_X1 U10800 ( .A(P1_D_REG_14__SCAN_IN), .ZN(n10134) );
  NOR2_X1 U10801 ( .A1(n10146), .A2(n10134), .ZN(P1_U3309) );
  INV_X1 U10802 ( .A(P1_D_REG_15__SCAN_IN), .ZN(n10135) );
  NOR2_X1 U10803 ( .A1(n10146), .A2(n10135), .ZN(P1_U3308) );
  INV_X1 U10804 ( .A(P1_D_REG_16__SCAN_IN), .ZN(n10136) );
  NOR2_X1 U10805 ( .A1(n10146), .A2(n10136), .ZN(P1_U3307) );
  INV_X1 U10806 ( .A(P1_D_REG_17__SCAN_IN), .ZN(n10137) );
  NOR2_X1 U10807 ( .A1(n10146), .A2(n10137), .ZN(P1_U3306) );
  INV_X1 U10808 ( .A(P1_D_REG_18__SCAN_IN), .ZN(n10138) );
  NOR2_X1 U10809 ( .A1(n10146), .A2(n10138), .ZN(P1_U3305) );
  INV_X1 U10810 ( .A(P1_D_REG_19__SCAN_IN), .ZN(n10139) );
  NOR2_X1 U10811 ( .A1(n10146), .A2(n10139), .ZN(P1_U3304) );
  INV_X1 U10812 ( .A(P1_D_REG_20__SCAN_IN), .ZN(n10140) );
  NOR2_X1 U10813 ( .A1(n10146), .A2(n10140), .ZN(P1_U3303) );
  INV_X1 U10814 ( .A(P1_D_REG_21__SCAN_IN), .ZN(n10141) );
  NOR2_X1 U10815 ( .A1(n10146), .A2(n10141), .ZN(P1_U3302) );
  INV_X1 U10816 ( .A(P1_D_REG_22__SCAN_IN), .ZN(n10142) );
  NOR2_X1 U10817 ( .A1(n10146), .A2(n10142), .ZN(P1_U3301) );
  INV_X1 U10818 ( .A(P1_D_REG_23__SCAN_IN), .ZN(n10143) );
  NOR2_X1 U10819 ( .A1(n10146), .A2(n10143), .ZN(P1_U3300) );
  INV_X1 U10820 ( .A(P1_D_REG_24__SCAN_IN), .ZN(n10144) );
  NOR2_X1 U10821 ( .A1(n10146), .A2(n10144), .ZN(P1_U3299) );
  INV_X1 U10822 ( .A(P1_D_REG_25__SCAN_IN), .ZN(n10145) );
  NOR2_X1 U10823 ( .A1(n10146), .A2(n10145), .ZN(P1_U3298) );
  INV_X1 U10824 ( .A(P1_D_REG_26__SCAN_IN), .ZN(n10147) );
  NOR2_X1 U10825 ( .A1(n10146), .A2(n10147), .ZN(P1_U3297) );
  INV_X1 U10826 ( .A(P1_D_REG_27__SCAN_IN), .ZN(n10148) );
  NOR2_X1 U10827 ( .A1(n10146), .A2(n10148), .ZN(P1_U3296) );
  INV_X1 U10828 ( .A(P1_D_REG_28__SCAN_IN), .ZN(n10149) );
  NOR2_X1 U10829 ( .A1(n10146), .A2(n10149), .ZN(P1_U3295) );
  INV_X1 U10830 ( .A(P1_D_REG_29__SCAN_IN), .ZN(n10150) );
  NOR2_X1 U10831 ( .A1(n10146), .A2(n10150), .ZN(P1_U3294) );
  INV_X1 U10832 ( .A(P1_D_REG_30__SCAN_IN), .ZN(n10151) );
  NOR2_X1 U10833 ( .A1(n10146), .A2(n10151), .ZN(P1_U3293) );
  INV_X1 U10834 ( .A(P1_D_REG_31__SCAN_IN), .ZN(n10152) );
  NOR2_X1 U10835 ( .A1(n10146), .A2(n10152), .ZN(P1_U3292) );
  INV_X1 U10836 ( .A(n10153), .ZN(n10157) );
  INV_X1 U10837 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n10156) );
  AOI22_X1 U10838 ( .A1(n10157), .A2(n10331), .B1(n10156), .B2(n10329), .ZN(
        P2_U3438) );
  AND2_X1 U10839 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n10329), .ZN(P2_U3326) );
  AND2_X1 U10840 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n10329), .ZN(P2_U3325) );
  AND2_X1 U10841 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n10329), .ZN(P2_U3324) );
  AND2_X1 U10842 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n10329), .ZN(P2_U3323) );
  AND2_X1 U10843 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n10329), .ZN(P2_U3322) );
  AND2_X1 U10844 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n10329), .ZN(P2_U3321) );
  AND2_X1 U10845 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n10329), .ZN(P2_U3320) );
  AND2_X1 U10846 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n10329), .ZN(P2_U3319) );
  AND2_X1 U10847 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n10329), .ZN(P2_U3318) );
  AND2_X1 U10848 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n10329), .ZN(P2_U3317) );
  AND2_X1 U10849 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n10329), .ZN(P2_U3316) );
  AND2_X1 U10850 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n10329), .ZN(P2_U3315) );
  AND2_X1 U10851 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n10329), .ZN(P2_U3314) );
  AND2_X1 U10852 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n10329), .ZN(P2_U3313) );
  AND2_X1 U10853 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n10329), .ZN(P2_U3312) );
  AND2_X1 U10854 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n10329), .ZN(P2_U3311) );
  AND2_X1 U10855 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n10329), .ZN(P2_U3310) );
  AND2_X1 U10856 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n10329), .ZN(P2_U3309) );
  AND2_X1 U10857 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n10329), .ZN(P2_U3308) );
  AND2_X1 U10858 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n10329), .ZN(P2_U3307) );
  AND2_X1 U10859 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n10329), .ZN(P2_U3306) );
  AND2_X1 U10860 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n10329), .ZN(P2_U3305) );
  AND2_X1 U10861 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n10329), .ZN(P2_U3304) );
  AND2_X1 U10862 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n10329), .ZN(P2_U3303) );
  AND2_X1 U10863 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n10329), .ZN(P2_U3302) );
  AND2_X1 U10864 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n10329), .ZN(P2_U3301) );
  AND2_X1 U10865 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n10329), .ZN(P2_U3300) );
  AND2_X1 U10866 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n10329), .ZN(P2_U3299) );
  AND2_X1 U10867 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n10329), .ZN(P2_U3298) );
  AND2_X1 U10868 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n10329), .ZN(P2_U3297) );
  XOR2_X1 U10869 ( .A(P2_ADDR_REG_0__SCAN_IN), .B(P1_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1071_U46) );
  NAND3_X1 U10870 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_0__SCAN_IN), .ZN(n10160) );
  AOI21_X1 U10871 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10162) );
  INV_X1 U10872 ( .A(n10162), .ZN(n10158) );
  NAND2_X1 U10873 ( .A1(n10160), .A2(n10158), .ZN(n10159) );
  XNOR2_X1 U10874 ( .A(P2_ADDR_REG_1__SCAN_IN), .B(n10159), .ZN(ADD_1071_U5)
         );
  XOR2_X1 U10875 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(P2_ADDR_REG_2__SCAN_IN), .Z(
        n10164) );
  INV_X1 U10876 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10161) );
  OAI21_X1 U10877 ( .B1(n10162), .B2(n10161), .A(n10160), .ZN(n10163) );
  XOR2_X1 U10878 ( .A(n10164), .B(n10163), .Z(ADD_1071_U54) );
  XOR2_X1 U10879 ( .A(P2_ADDR_REG_3__SCAN_IN), .B(P1_ADDR_REG_3__SCAN_IN), .Z(
        n10168) );
  NAND2_X1 U10880 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n10166) );
  NAND2_X1 U10881 ( .A1(n10164), .A2(n10163), .ZN(n10165) );
  NAND2_X1 U10882 ( .A1(n10166), .A2(n10165), .ZN(n10167) );
  XOR2_X1 U10883 ( .A(n10168), .B(n10167), .Z(ADD_1071_U53) );
  XNOR2_X1 U10884 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10172) );
  NAND2_X1 U10885 ( .A1(P2_ADDR_REG_3__SCAN_IN), .A2(P1_ADDR_REG_3__SCAN_IN), 
        .ZN(n10170) );
  NAND2_X1 U10886 ( .A1(n10168), .A2(n10167), .ZN(n10169) );
  NAND2_X1 U10887 ( .A1(n10170), .A2(n10169), .ZN(n10171) );
  XNOR2_X1 U10888 ( .A(n10172), .B(n10171), .ZN(ADD_1071_U52) );
  NOR2_X1 U10889 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10174) );
  NOR2_X1 U10890 ( .A1(n10172), .A2(n10171), .ZN(n10173) );
  NOR2_X1 U10891 ( .A1(n10174), .A2(n10173), .ZN(n10175) );
  AND2_X1 U10892 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n10175), .ZN(n10178) );
  NOR2_X1 U10893 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n10175), .ZN(n10180) );
  NOR2_X1 U10894 ( .A1(n10178), .A2(n10180), .ZN(n10177) );
  XNOR2_X1 U10895 ( .A(n10177), .B(n10176), .ZN(ADD_1071_U51) );
  NOR2_X1 U10896 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n10178), .ZN(n10179) );
  NOR2_X1 U10897 ( .A1(n10180), .A2(n10179), .ZN(n10182) );
  XOR2_X1 U10898 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(n10182), .Z(n10183) );
  XNOR2_X1 U10899 ( .A(n10183), .B(n10181), .ZN(ADD_1071_U50) );
  NAND2_X1 U10900 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(n10182), .ZN(n10185) );
  NAND2_X1 U10901 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(n10183), .ZN(n10184) );
  NAND2_X1 U10902 ( .A1(n10185), .A2(n10184), .ZN(n10187) );
  XOR2_X1 U10903 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n10187), .Z(n10188) );
  XNOR2_X1 U10904 ( .A(n10188), .B(n10186), .ZN(ADD_1071_U49) );
  NAND2_X1 U10905 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n10187), .ZN(n10190) );
  NAND2_X1 U10906 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n10188), .ZN(n10189) );
  NAND2_X1 U10907 ( .A1(n10190), .A2(n10189), .ZN(n10192) );
  XOR2_X1 U10908 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(n10192), .Z(n10193) );
  XNOR2_X1 U10909 ( .A(n10193), .B(n10191), .ZN(ADD_1071_U48) );
  NAND2_X1 U10910 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n10192), .ZN(n10195) );
  NAND2_X1 U10911 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n10193), .ZN(n10194) );
  NAND2_X1 U10912 ( .A1(n10195), .A2(n10194), .ZN(n10197) );
  XOR2_X1 U10913 ( .A(P1_ADDR_REG_9__SCAN_IN), .B(n10197), .Z(n10198) );
  XNOR2_X1 U10914 ( .A(n10198), .B(n10196), .ZN(ADD_1071_U47) );
  XOR2_X1 U10915 ( .A(P2_ADDR_REG_10__SCAN_IN), .B(P1_ADDR_REG_10__SCAN_IN), 
        .Z(n10202) );
  NAND2_X1 U10916 ( .A1(P1_ADDR_REG_9__SCAN_IN), .A2(n10197), .ZN(n10200) );
  NAND2_X1 U10917 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n10198), .ZN(n10199) );
  NAND2_X1 U10918 ( .A1(n10200), .A2(n10199), .ZN(n10201) );
  XOR2_X1 U10919 ( .A(n10202), .B(n10201), .Z(ADD_1071_U63) );
  XOR2_X1 U10920 ( .A(P2_ADDR_REG_11__SCAN_IN), .B(P1_ADDR_REG_11__SCAN_IN), 
        .Z(n10206) );
  NAND2_X1 U10921 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n10204) );
  NAND2_X1 U10922 ( .A1(n10202), .A2(n10201), .ZN(n10203) );
  NAND2_X1 U10923 ( .A1(n10204), .A2(n10203), .ZN(n10205) );
  XOR2_X1 U10924 ( .A(n10206), .B(n10205), .Z(ADD_1071_U62) );
  NAND2_X1 U10925 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n10208) );
  NAND2_X1 U10926 ( .A1(n10206), .A2(n10205), .ZN(n10207) );
  NAND2_X1 U10927 ( .A1(n10208), .A2(n10207), .ZN(n10210) );
  XNOR2_X1 U10928 ( .A(P2_ADDR_REG_12__SCAN_IN), .B(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n10209) );
  XNOR2_X1 U10929 ( .A(n10210), .B(n10209), .ZN(ADD_1071_U61) );
  NOR2_X1 U10930 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n10212) );
  NOR2_X1 U10931 ( .A1(n10210), .A2(n10209), .ZN(n10211) );
  XNOR2_X1 U10932 ( .A(P2_ADDR_REG_13__SCAN_IN), .B(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n10213) );
  XNOR2_X1 U10933 ( .A(n10214), .B(n10213), .ZN(ADD_1071_U60) );
  NOR2_X1 U10934 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n10216) );
  NOR2_X1 U10935 ( .A1(n10214), .A2(n10213), .ZN(n10215) );
  XNOR2_X1 U10936 ( .A(P2_ADDR_REG_14__SCAN_IN), .B(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n10217) );
  XNOR2_X1 U10937 ( .A(n10218), .B(n10217), .ZN(ADD_1071_U59) );
  NOR2_X1 U10938 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n10220) );
  NOR2_X1 U10939 ( .A1(n10218), .A2(n10217), .ZN(n10219) );
  NOR2_X1 U10940 ( .A1(n10220), .A2(n10219), .ZN(n10222) );
  XNOR2_X1 U10941 ( .A(P2_ADDR_REG_15__SCAN_IN), .B(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n10221) );
  XNOR2_X1 U10942 ( .A(n10222), .B(n10221), .ZN(ADD_1071_U58) );
  NOR2_X1 U10943 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n10224) );
  NOR2_X1 U10944 ( .A1(n10222), .A2(n10221), .ZN(n10223) );
  NOR2_X1 U10945 ( .A1(n10224), .A2(n10223), .ZN(n10226) );
  XNOR2_X1 U10946 ( .A(P2_ADDR_REG_16__SCAN_IN), .B(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n10225) );
  XNOR2_X1 U10947 ( .A(n10226), .B(n10225), .ZN(ADD_1071_U57) );
  NOR2_X1 U10948 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n10228) );
  NOR2_X1 U10949 ( .A1(n10226), .A2(n10225), .ZN(n10227) );
  NOR2_X1 U10950 ( .A1(n10228), .A2(n10227), .ZN(n10230) );
  XNOR2_X1 U10951 ( .A(P2_ADDR_REG_17__SCAN_IN), .B(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n10229) );
  XNOR2_X1 U10952 ( .A(n10230), .B(n10229), .ZN(ADD_1071_U56) );
  NOR2_X1 U10953 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n10232) );
  NOR2_X1 U10954 ( .A1(n10230), .A2(n10229), .ZN(n10231) );
  NOR2_X1 U10955 ( .A1(n10232), .A2(n10231), .ZN(n10233) );
  NOR2_X1 U10956 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(n10233), .ZN(n10236) );
  AND2_X1 U10957 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(n10233), .ZN(n10235) );
  NOR2_X1 U10958 ( .A1(n10236), .A2(n10235), .ZN(n10234) );
  XOR2_X1 U10959 ( .A(P1_ADDR_REG_18__SCAN_IN), .B(n10234), .Z(ADD_1071_U55)
         );
  NOR2_X1 U10960 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n10235), .ZN(n10237) );
  NOR2_X1 U10961 ( .A1(n10237), .A2(n10236), .ZN(n10239) );
  XNOR2_X1 U10962 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(P1_ADDR_REG_19__SCAN_IN), 
        .ZN(n10238) );
  XNOR2_X1 U10963 ( .A(n10239), .B(n10238), .ZN(ADD_1071_U4) );
  AOI21_X1 U10964 ( .B1(n10242), .B2(n10241), .A(n10240), .ZN(P1_U3441) );
  INV_X1 U10965 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n10375) );
  INV_X1 U10966 ( .A(n10243), .ZN(n10244) );
  OAI21_X1 U10967 ( .B1(n10245), .B2(P1_REG1_REG_0__SCAN_IN), .A(n10244), .ZN(
        n10252) );
  NOR4_X1 U10968 ( .A1(n10248), .A2(n10247), .A3(n10246), .A4(P1_U3084), .ZN(
        n10249) );
  AOI21_X1 U10969 ( .B1(n10320), .B2(n10250), .A(n10249), .ZN(n10251) );
  AOI21_X1 U10970 ( .B1(n10253), .B2(n10252), .A(n10251), .ZN(n10254) );
  AOI21_X1 U10971 ( .B1(n10313), .B2(P1_ADDR_REG_0__SCAN_IN), .A(n10254), .ZN(
        n10255) );
  OAI21_X1 U10972 ( .B1(P1_STATE_REG_SCAN_IN), .B2(n10375), .A(n10255), .ZN(
        P1_U3241) );
  AOI22_X1 U10973 ( .A1(n10313), .A2(P1_ADDR_REG_6__SCAN_IN), .B1(n10312), 
        .B2(n10256), .ZN(n10267) );
  AOI21_X1 U10974 ( .B1(n10259), .B2(n10258), .A(n10257), .ZN(n10260) );
  NAND2_X1 U10975 ( .A1(n10318), .A2(n10260), .ZN(n10265) );
  OAI211_X1 U10976 ( .C1(n10263), .C2(n10262), .A(n10320), .B(n10261), .ZN(
        n10264) );
  NAND4_X1 U10977 ( .A1(n10267), .A2(n10266), .A3(n10265), .A4(n10264), .ZN(
        P1_U3247) );
  AOI22_X1 U10978 ( .A1(n10313), .A2(P1_ADDR_REG_11__SCAN_IN), .B1(n10312), 
        .B2(n10268), .ZN(n10285) );
  NOR3_X1 U10979 ( .A1(n10269), .A2(n10530), .A3(n10278), .ZN(n10276) );
  AOI211_X1 U10980 ( .C1(n10271), .C2(n10273), .A(n10270), .B(n10298), .ZN(
        n10275) );
  AOI211_X1 U10981 ( .C1(n10277), .C2(n10276), .A(n10275), .B(n4916), .ZN(
        n10284) );
  NAND3_X1 U10982 ( .A1(n10279), .A2(n10530), .A3(n10278), .ZN(n10280) );
  NAND3_X1 U10983 ( .A1(n10320), .A2(n10281), .A3(n10280), .ZN(n10282) );
  NAND4_X1 U10984 ( .A1(n10285), .A2(n10284), .A3(n10283), .A4(n10282), .ZN(
        P1_U3252) );
  OAI21_X1 U10985 ( .B1(n10288), .B2(n10287), .A(n10286), .ZN(n10289) );
  AOI22_X1 U10986 ( .A1(n10289), .A2(n10320), .B1(n10313), .B2(
        P1_ADDR_REG_13__SCAN_IN), .ZN(n10297) );
  OAI211_X1 U10987 ( .C1(n10292), .C2(n10291), .A(n10318), .B(n10290), .ZN(
        n10295) );
  NAND2_X1 U10988 ( .A1(n10312), .A2(n10293), .ZN(n10294) );
  NAND4_X1 U10989 ( .A1(n10297), .A2(n10296), .A3(n10295), .A4(n10294), .ZN(
        P1_U3254) );
  AOI211_X1 U10990 ( .C1(n10301), .C2(n10300), .A(n10299), .B(n10298), .ZN(
        n10302) );
  AOI211_X1 U10991 ( .C1(n10304), .C2(n10312), .A(n10303), .B(n10302), .ZN(
        n10310) );
  OAI21_X1 U10992 ( .B1(n10307), .B2(n10306), .A(n10305), .ZN(n10308) );
  AOI22_X1 U10993 ( .A1(n10308), .A2(n10320), .B1(n10313), .B2(
        P1_ADDR_REG_18__SCAN_IN), .ZN(n10309) );
  NAND2_X1 U10994 ( .A1(n10310), .A2(n10309), .ZN(P1_U3259) );
  AOI22_X1 U10995 ( .A1(n10313), .A2(P1_ADDR_REG_5__SCAN_IN), .B1(n10312), 
        .B2(n10311), .ZN(n10326) );
  OAI21_X1 U10996 ( .B1(n10316), .B2(n10315), .A(n10314), .ZN(n10317) );
  NAND2_X1 U10997 ( .A1(n10318), .A2(n10317), .ZN(n10324) );
  OAI211_X1 U10998 ( .C1(n10322), .C2(n10321), .A(n10320), .B(n10319), .ZN(
        n10323) );
  NAND4_X1 U10999 ( .A1(n10326), .A2(n10325), .A3(n10324), .A4(n10323), .ZN(
        P1_U3246) );
  NOR2_X1 U11000 ( .A1(n10328), .A2(n10327), .ZN(n10332) );
  INV_X1 U11001 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n10330) );
  AOI22_X1 U11002 ( .A1(n10332), .A2(n10331), .B1(n10330), .B2(n10329), .ZN(
        P2_U3437) );
  AOI22_X1 U11003 ( .A1(n10334), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n10333), .ZN(n10340) );
  AOI22_X1 U11004 ( .A1(n10352), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3152), .ZN(n10339) );
  OAI21_X1 U11005 ( .B1(P2_REG1_REG_0__SCAN_IN), .B2(n10353), .A(n10335), .ZN(
        n10337) );
  NOR2_X1 U11006 ( .A1(n10357), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n10336) );
  OAI21_X1 U11007 ( .B1(n10337), .B2(n10336), .A(P2_IR_REG_0__SCAN_IN), .ZN(
        n10338) );
  OAI211_X1 U11008 ( .C1(P2_IR_REG_0__SCAN_IN), .C2(n10340), .A(n10339), .B(
        n10338), .ZN(P2_U3245) );
  AOI22_X1 U11009 ( .A1(n10352), .A2(P2_ADDR_REG_1__SCAN_IN), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(P2_U3152), .ZN(n10351) );
  AOI211_X1 U11010 ( .C1(n10343), .C2(n10342), .A(n10341), .B(n10353), .ZN(
        n10348) );
  AOI211_X1 U11011 ( .C1(n10346), .C2(n10345), .A(n10344), .B(n10357), .ZN(
        n10347) );
  AOI211_X1 U11012 ( .C1(n10364), .C2(n10349), .A(n10348), .B(n10347), .ZN(
        n10350) );
  NAND2_X1 U11013 ( .A1(n10351), .A2(n10350), .ZN(P2_U3246) );
  AOI22_X1 U11014 ( .A1(n10352), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3152), .ZN(n10366) );
  AOI211_X1 U11015 ( .C1(n10356), .C2(n10355), .A(n10354), .B(n10353), .ZN(
        n10362) );
  AOI211_X1 U11016 ( .C1(n10360), .C2(n10359), .A(n10358), .B(n10357), .ZN(
        n10361) );
  AOI211_X1 U11017 ( .C1(n10364), .C2(n10363), .A(n10362), .B(n10361), .ZN(
        n10365) );
  NAND2_X1 U11018 ( .A1(n10366), .A2(n10365), .ZN(P2_U3247) );
  XNOR2_X1 U11019 ( .A(P2_RD_REG_SCAN_IN), .B(P1_RD_REG_SCAN_IN), .ZN(U126) );
  NAND2_X1 U11020 ( .A1(n10419), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n10370) );
  OAI21_X1 U11021 ( .B1(n10368), .B2(n10367), .A(n10385), .ZN(n10369) );
  OAI211_X1 U11022 ( .C1(n10372), .C2(n10371), .A(n10370), .B(n10369), .ZN(
        n10373) );
  INV_X1 U11023 ( .A(n10373), .ZN(n10374) );
  OAI21_X1 U11024 ( .B1(n10376), .B2(n10375), .A(n10374), .ZN(P1_U3291) );
  AOI22_X1 U11025 ( .A1(n10541), .A2(n10379), .B1(n10378), .B2(n10377), .ZN(
        n10380) );
  AND2_X1 U11026 ( .A1(n10381), .A2(n10380), .ZN(n10383) );
  AOI22_X1 U11027 ( .A1(n10553), .A2(n10383), .B1(n6342), .B2(n10551), .ZN(
        P2_U3520) );
  INV_X1 U11028 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n10382) );
  AOI22_X1 U11029 ( .A1(n10557), .A2(n10383), .B1(n10382), .B2(n10554), .ZN(
        P2_U3451) );
  XOR2_X1 U11030 ( .A(n10384), .B(n10395), .Z(n10402) );
  INV_X1 U11031 ( .A(n10402), .ZN(n10416) );
  INV_X1 U11032 ( .A(n10408), .ZN(n10390) );
  NAND2_X1 U11033 ( .A1(n10408), .A2(n10385), .ZN(n10387) );
  NAND2_X1 U11034 ( .A1(n10387), .A2(n10386), .ZN(n10389) );
  OR2_X1 U11035 ( .A1(n10389), .A2(n10388), .ZN(n10412) );
  OAI21_X1 U11036 ( .B1(n10390), .B2(n10520), .A(n10412), .ZN(n10403) );
  AOI22_X1 U11037 ( .A1(n10393), .A2(n6205), .B1(n10392), .B2(n10391), .ZN(
        n10400) );
  OAI21_X1 U11038 ( .B1(n10396), .B2(n10395), .A(n10394), .ZN(n10398) );
  NAND2_X1 U11039 ( .A1(n10398), .A2(n10397), .ZN(n10399) );
  OAI211_X1 U11040 ( .C1(n10402), .C2(n10401), .A(n10400), .B(n10399), .ZN(
        n10414) );
  AOI211_X1 U11041 ( .C1(n10525), .C2(n10416), .A(n10403), .B(n10414), .ZN(
        n10405) );
  AOI22_X1 U11042 ( .A1(n10531), .A2(n10405), .B1(n7185), .B2(n10529), .ZN(
        P1_U3524) );
  INV_X1 U11043 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n10404) );
  AOI22_X1 U11044 ( .A1(n10535), .A2(n10405), .B1(n10404), .B2(n10532), .ZN(
        P1_U3457) );
  INV_X1 U11045 ( .A(n10406), .ZN(n10407) );
  AOI22_X1 U11046 ( .A1(n10409), .A2(P1_REG3_REG_1__SCAN_IN), .B1(n10408), 
        .B2(n10407), .ZN(n10410) );
  OAI21_X1 U11047 ( .B1(n10412), .B2(n10411), .A(n10410), .ZN(n10413) );
  NOR2_X1 U11048 ( .A1(n10414), .A2(n10413), .ZN(n10418) );
  AOI22_X1 U11049 ( .A1(n10416), .A2(n10415), .B1(P1_REG2_REG_1__SCAN_IN), 
        .B2(n10419), .ZN(n10417) );
  OAI21_X1 U11050 ( .B1(n10419), .B2(n10418), .A(n10417), .ZN(P1_U3290) );
  OAI22_X1 U11051 ( .A1(n10421), .A2(n10522), .B1(n10420), .B2(n10520), .ZN(
        n10423) );
  AOI211_X1 U11052 ( .C1(n10525), .C2(n10424), .A(n10423), .B(n10422), .ZN(
        n10427) );
  INV_X1 U11053 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n10425) );
  AOI22_X1 U11054 ( .A1(n10531), .A2(n10427), .B1(n10425), .B2(n10529), .ZN(
        P1_U3525) );
  INV_X1 U11055 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n10426) );
  AOI22_X1 U11056 ( .A1(n10535), .A2(n10427), .B1(n10426), .B2(n10532), .ZN(
        P1_U3460) );
  INV_X1 U11057 ( .A(n10428), .ZN(n10433) );
  AOI22_X1 U11058 ( .A1(n10430), .A2(n10429), .B1(n10550), .B2(n7054), .ZN(
        n10431) );
  OAI211_X1 U11059 ( .C1(n10433), .C2(n10510), .A(n10432), .B(n10431), .ZN(
        n10434) );
  INV_X1 U11060 ( .A(n10434), .ZN(n10435) );
  AOI22_X1 U11061 ( .A1(n10553), .A2(n10435), .B1(n7379), .B2(n10551), .ZN(
        P2_U3522) );
  AOI22_X1 U11062 ( .A1(n10557), .A2(n10435), .B1(n6351), .B2(n10554), .ZN(
        P2_U3457) );
  INV_X1 U11063 ( .A(n10436), .ZN(n10441) );
  OAI22_X1 U11064 ( .A1(n10437), .A2(n10522), .B1(n4989), .B2(n10520), .ZN(
        n10439) );
  AOI211_X1 U11065 ( .C1(n10441), .C2(n10440), .A(n10439), .B(n10438), .ZN(
        n10444) );
  AOI22_X1 U11066 ( .A1(n10531), .A2(n10444), .B1(n10442), .B2(n10529), .ZN(
        P1_U3527) );
  INV_X1 U11067 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n10443) );
  AOI22_X1 U11068 ( .A1(n10535), .A2(n10444), .B1(n10443), .B2(n10532), .ZN(
        P1_U3466) );
  OAI22_X1 U11069 ( .A1(n10446), .A2(n10545), .B1(n10445), .B2(n10536), .ZN(
        n10447) );
  AOI211_X1 U11070 ( .C1(n10449), .C2(n10541), .A(n10448), .B(n10447), .ZN(
        n10451) );
  AOI22_X1 U11071 ( .A1(n10553), .A2(n10451), .B1(n6385), .B2(n10551), .ZN(
        P2_U3524) );
  INV_X1 U11072 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n10450) );
  AOI22_X1 U11073 ( .A1(n10557), .A2(n10451), .B1(n10450), .B2(n10554), .ZN(
        P2_U3463) );
  INV_X1 U11074 ( .A(n10452), .ZN(n10455) );
  OAI22_X1 U11075 ( .A1(n10456), .A2(n10455), .B1(n10454), .B2(n10453), .ZN(
        n10457) );
  INV_X1 U11076 ( .A(n10457), .ZN(n10458) );
  OAI211_X1 U11077 ( .C1(n10461), .C2(n10460), .A(n10459), .B(n10458), .ZN(
        n10462) );
  AOI21_X1 U11078 ( .B1(n10464), .B2(n10463), .A(n10462), .ZN(n10465) );
  AOI22_X1 U11079 ( .A1(n10466), .A2(n6396), .B1(n10465), .B2(n8810), .ZN(
        P2_U3291) );
  OAI22_X1 U11080 ( .A1(n10468), .A2(n10522), .B1(n10467), .B2(n10520), .ZN(
        n10470) );
  AOI211_X1 U11081 ( .C1(n10525), .C2(n10471), .A(n10470), .B(n10469), .ZN(
        n10473) );
  AOI22_X1 U11082 ( .A1(n10531), .A2(n10473), .B1(n7184), .B2(n10529), .ZN(
        P1_U3529) );
  INV_X1 U11083 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n10472) );
  AOI22_X1 U11084 ( .A1(n10535), .A2(n10473), .B1(n10472), .B2(n10532), .ZN(
        P1_U3472) );
  OAI22_X1 U11085 ( .A1(n10475), .A2(n10545), .B1(n10474), .B2(n10536), .ZN(
        n10477) );
  AOI211_X1 U11086 ( .C1(n10541), .C2(n10478), .A(n10477), .B(n10476), .ZN(
        n10480) );
  AOI22_X1 U11087 ( .A1(n10553), .A2(n10480), .B1(n6412), .B2(n10551), .ZN(
        P2_U3526) );
  INV_X1 U11088 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10479) );
  AOI22_X1 U11089 ( .A1(n10557), .A2(n10480), .B1(n10479), .B2(n10554), .ZN(
        P2_U3469) );
  OAI22_X1 U11090 ( .A1(n10482), .A2(n10522), .B1(n10481), .B2(n10520), .ZN(
        n10484) );
  AOI211_X1 U11091 ( .C1(n10525), .C2(n10485), .A(n10484), .B(n10483), .ZN(
        n10488) );
  AOI22_X1 U11092 ( .A1(n10531), .A2(n10488), .B1(n10486), .B2(n10529), .ZN(
        P1_U3531) );
  INV_X1 U11093 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n10487) );
  AOI22_X1 U11094 ( .A1(n10535), .A2(n10488), .B1(n10487), .B2(n10532), .ZN(
        P1_U3478) );
  INV_X1 U11095 ( .A(n10489), .ZN(n10495) );
  INV_X1 U11096 ( .A(n10490), .ZN(n10491) );
  OAI22_X1 U11097 ( .A1(n10492), .A2(n10522), .B1(n10491), .B2(n10520), .ZN(
        n10494) );
  AOI211_X1 U11098 ( .C1(n10525), .C2(n10495), .A(n10494), .B(n10493), .ZN(
        n10498) );
  AOI22_X1 U11099 ( .A1(n10531), .A2(n10498), .B1(n10496), .B2(n10529), .ZN(
        P1_U3532) );
  INV_X1 U11100 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n10497) );
  AOI22_X1 U11101 ( .A1(n10535), .A2(n10498), .B1(n10497), .B2(n10532), .ZN(
        P1_U3481) );
  INV_X1 U11102 ( .A(n10505), .ZN(n10507) );
  AOI211_X1 U11103 ( .C1(n10502), .C2(n10501), .A(n10500), .B(n10499), .ZN(
        n10503) );
  OAI21_X1 U11104 ( .B1(n10505), .B2(n10504), .A(n10503), .ZN(n10506) );
  AOI21_X1 U11105 ( .B1(n6266), .B2(n10507), .A(n10506), .ZN(n10509) );
  AOI22_X1 U11106 ( .A1(n10531), .A2(n10509), .B1(n7498), .B2(n10529), .ZN(
        P1_U3533) );
  INV_X1 U11107 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n10508) );
  AOI22_X1 U11108 ( .A1(n10535), .A2(n10509), .B1(n10508), .B2(n10532), .ZN(
        P1_U3484) );
  INV_X1 U11109 ( .A(n10510), .ZN(n10518) );
  INV_X1 U11110 ( .A(n10511), .ZN(n10517) );
  INV_X1 U11111 ( .A(n10512), .ZN(n10513) );
  OAI22_X1 U11112 ( .A1(n10514), .A2(n10545), .B1(n10513), .B2(n10536), .ZN(
        n10516) );
  AOI211_X1 U11113 ( .C1(n10518), .C2(n10517), .A(n10516), .B(n10515), .ZN(
        n10519) );
  AOI22_X1 U11114 ( .A1(n10553), .A2(n10519), .B1(n7524), .B2(n10551), .ZN(
        P2_U3530) );
  AOI22_X1 U11115 ( .A1(n10557), .A2(n10519), .B1(n6470), .B2(n10554), .ZN(
        P2_U3481) );
  OAI22_X1 U11116 ( .A1(n10523), .A2(n10522), .B1(n10521), .B2(n10520), .ZN(
        n10524) );
  AOI21_X1 U11117 ( .B1(n10526), .B2(n10525), .A(n10524), .ZN(n10527) );
  AND2_X1 U11118 ( .A1(n10528), .A2(n10527), .ZN(n10534) );
  AOI22_X1 U11119 ( .A1(n10531), .A2(n10534), .B1(n10530), .B2(n10529), .ZN(
        P1_U3534) );
  INV_X1 U11120 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n10533) );
  AOI22_X1 U11121 ( .A1(n10535), .A2(n10534), .B1(n10533), .B2(n10532), .ZN(
        P1_U3487) );
  OAI22_X1 U11122 ( .A1(n10538), .A2(n10545), .B1(n10537), .B2(n10536), .ZN(
        n10540) );
  AOI211_X1 U11123 ( .C1(n10542), .C2(n10541), .A(n10540), .B(n10539), .ZN(
        n10544) );
  AOI22_X1 U11124 ( .A1(n10553), .A2(n10544), .B1(n7884), .B2(n10551), .ZN(
        P2_U3532) );
  INV_X1 U11125 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n10543) );
  AOI22_X1 U11126 ( .A1(n10557), .A2(n10544), .B1(n10543), .B2(n10554), .ZN(
        P2_U3487) );
  NOR2_X1 U11127 ( .A1(n10546), .A2(n10545), .ZN(n10547) );
  INV_X1 U11128 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n10552) );
  AOI22_X1 U11129 ( .A1(n10553), .A2(n10556), .B1(n10552), .B2(n10551), .ZN(
        P2_U3550) );
  INV_X1 U11130 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n10555) );
  AOI22_X1 U11131 ( .A1(n10557), .A2(n10556), .B1(n10555), .B2(n10554), .ZN(
        P2_U3518) );
  XNOR2_X1 U11132 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  NAND2_X1 U6093 ( .A1(n6318), .A2(n6314), .ZN(n8512) );
  CLKBUF_X3 U5018 ( .A(n5519), .Z(n4854) );
  NAND2_X1 U6003 ( .A1(n4928), .A2(n10377), .ZN(n7286) );
  NAND2_X1 U7238 ( .A1(n6157), .A2(n9978), .ZN(n9554) );
  NAND3_X1 U6009 ( .A1(n5325), .A2(n6300), .A3(n5324), .ZN(n6314) );
  CLKBUF_X1 U4947 ( .A(n6865), .Z(n7001) );
  CLKBUF_X1 U5022 ( .A(n6307), .Z(n6305) );
  NAND2_X2 U5113 ( .A1(n6741), .A2(n8512), .ZN(n6348) );
  CLKBUF_X3 U6235 ( .A(n5548), .Z(n4855) );
  CLKBUF_X1 U6283 ( .A(n6703), .Z(n10461) );
endmodule

