

module b20_C_2inp_gates_syn ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, ADD_1068_U4, 
        ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58, ADD_1068_U59, 
        ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63, ADD_1068_U47, 
        ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51, ADD_1068_U52, 
        ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46, U126, U123, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439, P1_U3440, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462, P1_U3465, P1_U3468, 
        P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, 
        P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3509, 
        P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, 
        P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, 
        P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, 
        P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, 
        P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, 
        P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, 
        P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3554, P1_U3555, 
        P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, 
        P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, 
        P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, 
        P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, 
        P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U3973, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376, P2_U3377, P2_U3263, 
        P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, 
        P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, 
        P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, 
        P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, 
        P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399, P2_U3402, P2_U3405, 
        P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420, P2_U3423, P2_U3426, 
        P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441, P2_U3444, P2_U3446, 
        P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451, P2_U3452, P2_U3453, 
        P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458, P2_U3459, P2_U3460, 
        P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465, P2_U3466, P2_U3467, 
        P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472, P2_U3473, P2_U3474, 
        P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479, P2_U3480, P2_U3481, 
        P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486, P2_U3487, P2_U3488, 
        P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, 
        P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, 
        P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, 
        P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3491, P2_U3492, 
        P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, 
        P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, 
        P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, 
        P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, 
        P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180, P2_U3179, P2_U3178, 
        P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, P2_U3171, 
        P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, P2_U3164, 
        P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, P2_U3157, 
        P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151, P2_U3150, P2_U3893, 
        keyinput127, keyinput126, keyinput125, keyinput124, keyinput123, 
        keyinput122, keyinput121, keyinput120, keyinput119, keyinput118, 
        keyinput117, keyinput116, keyinput115, keyinput114, keyinput113, 
        keyinput112, keyinput111, keyinput110, keyinput109, keyinput108, 
        keyinput107, keyinput106, keyinput105, keyinput104, keyinput103, 
        keyinput102, keyinput101, keyinput100, keyinput99, keyinput98, 
        keyinput97, keyinput96, keyinput95, keyinput94, keyinput93, keyinput92, 
        keyinput91, keyinput90, keyinput89, keyinput88, keyinput87, keyinput86, 
        keyinput85, keyinput84, keyinput83, keyinput82, keyinput81, keyinput80, 
        keyinput79, keyinput78, keyinput77, keyinput76, keyinput75, keyinput74, 
        keyinput73, keyinput72, keyinput71, keyinput70, keyinput69, keyinput68, 
        keyinput67, keyinput66, keyinput65, keyinput64, keyinput63, keyinput62, 
        keyinput61, keyinput60, keyinput59, keyinput58, keyinput57, keyinput56, 
        keyinput55, keyinput54, keyinput53, keyinput52, keyinput51, keyinput50, 
        keyinput49, keyinput48, keyinput47, keyinput46, keyinput45, keyinput44, 
        keyinput43, keyinput42, keyinput41, keyinput40, keyinput39, keyinput38, 
        keyinput37, keyinput36, keyinput35, keyinput34, keyinput33, keyinput32, 
        keyinput31, keyinput30, keyinput29, keyinput28, keyinput27, keyinput26, 
        keyinput25, keyinput24, keyinput23, keyinput22, keyinput21, keyinput20, 
        keyinput19, keyinput18, keyinput17, keyinput16, keyinput15, keyinput14, 
        keyinput13, keyinput12, keyinput11, keyinput10, keyinput9, keyinput8, 
        keyinput7, keyinput6, keyinput5, keyinput4, keyinput3, keyinput2, 
        keyinput1, keyinput0 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, keyinput127, keyinput126, keyinput125,
         keyinput124, keyinput123, keyinput122, keyinput121, keyinput120,
         keyinput119, keyinput118, keyinput117, keyinput116, keyinput115,
         keyinput114, keyinput113, keyinput112, keyinput111, keyinput110,
         keyinput109, keyinput108, keyinput107, keyinput106, keyinput105,
         keyinput104, keyinput103, keyinput102, keyinput101, keyinput100,
         keyinput99, keyinput98, keyinput97, keyinput96, keyinput95,
         keyinput94, keyinput93, keyinput92, keyinput91, keyinput90,
         keyinput89, keyinput88, keyinput87, keyinput86, keyinput85,
         keyinput84, keyinput83, keyinput82, keyinput81, keyinput80,
         keyinput79, keyinput78, keyinput77, keyinput76, keyinput75,
         keyinput74, keyinput73, keyinput72, keyinput71, keyinput70,
         keyinput69, keyinput68, keyinput67, keyinput66, keyinput65,
         keyinput64, keyinput63, keyinput62, keyinput61, keyinput60,
         keyinput59, keyinput58, keyinput57, keyinput56, keyinput55,
         keyinput54, keyinput53, keyinput52, keyinput51, keyinput50,
         keyinput49, keyinput48, keyinput47, keyinput46, keyinput45,
         keyinput44, keyinput43, keyinput42, keyinput41, keyinput40,
         keyinput39, keyinput38, keyinput37, keyinput36, keyinput35,
         keyinput34, keyinput33, keyinput32, keyinput31, keyinput30,
         keyinput29, keyinput28, keyinput27, keyinput26, keyinput25,
         keyinput24, keyinput23, keyinput22, keyinput21, keyinput20,
         keyinput19, keyinput18, keyinput17, keyinput16, keyinput15,
         keyinput14, keyinput13, keyinput12, keyinput11, keyinput10, keyinput9,
         keyinput8, keyinput7, keyinput6, keyinput5, keyinput4, keyinput3,
         keyinput2, keyinput1, keyinput0;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420,
         n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430,
         n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440,
         n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450,
         n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460,
         n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470,
         n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480,
         n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490,
         n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500,
         n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510,
         n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520,
         n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530,
         n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540,
         n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550,
         n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560,
         n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570,
         n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580,
         n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590,
         n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600,
         n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610,
         n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620,
         n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630,
         n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640,
         n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650,
         n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660,
         n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670,
         n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680,
         n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690,
         n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700,
         n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710,
         n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720,
         n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730,
         n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740,
         n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750,
         n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760,
         n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770,
         n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780,
         n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790,
         n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800,
         n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810,
         n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820,
         n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830,
         n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840,
         n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850,
         n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860,
         n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870,
         n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880,
         n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890,
         n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900,
         n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910,
         n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920,
         n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930,
         n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940,
         n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950,
         n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960,
         n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970,
         n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980,
         n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990,
         n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000,
         n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010,
         n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020,
         n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030,
         n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040,
         n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050,
         n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060,
         n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070,
         n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080,
         n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090,
         n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100,
         n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110,
         n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120,
         n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130,
         n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140,
         n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150,
         n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160,
         n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170,
         n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180,
         n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190,
         n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200,
         n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210,
         n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220,
         n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230,
         n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240,
         n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250,
         n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260,
         n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270,
         n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280,
         n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290,
         n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300,
         n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310,
         n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320,
         n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330,
         n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340,
         n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350,
         n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360,
         n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370,
         n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380,
         n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390,
         n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400,
         n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410,
         n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420,
         n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430,
         n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440,
         n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450,
         n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460,
         n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470,
         n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480,
         n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490,
         n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500,
         n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510,
         n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520,
         n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530,
         n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540,
         n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550,
         n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560,
         n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570,
         n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580,
         n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590,
         n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600,
         n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610,
         n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620,
         n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630,
         n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640,
         n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650,
         n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660,
         n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670,
         n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680,
         n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690,
         n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700,
         n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710,
         n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720,
         n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730,
         n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740,
         n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750,
         n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760,
         n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770,
         n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780,
         n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790,
         n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800,
         n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810,
         n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820,
         n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830,
         n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840,
         n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850,
         n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860,
         n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870,
         n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880,
         n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890,
         n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900,
         n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910,
         n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920,
         n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930,
         n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940,
         n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950,
         n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960,
         n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970,
         n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980,
         n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990,
         n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000,
         n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010,
         n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020,
         n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030,
         n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040,
         n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050,
         n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060,
         n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070,
         n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080,
         n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090,
         n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100,
         n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110,
         n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120,
         n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130,
         n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140,
         n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150,
         n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160,
         n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170,
         n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180,
         n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190,
         n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200,
         n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210,
         n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220,
         n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230,
         n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240,
         n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250,
         n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260,
         n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270,
         n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280,
         n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290,
         n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300,
         n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310,
         n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320,
         n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330,
         n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340,
         n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350,
         n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360,
         n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370,
         n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380,
         n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390,
         n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400,
         n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410,
         n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420,
         n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430,
         n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440,
         n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450,
         n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460,
         n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470,
         n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480,
         n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490,
         n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500,
         n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510,
         n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520,
         n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530,
         n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540,
         n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550,
         n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560,
         n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570,
         n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580,
         n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590,
         n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600,
         n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610,
         n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620,
         n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630,
         n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640,
         n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650,
         n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660,
         n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670,
         n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680,
         n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690,
         n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700,
         n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710,
         n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720,
         n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730,
         n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740,
         n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750,
         n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760,
         n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770,
         n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780,
         n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790,
         n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800,
         n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810,
         n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820,
         n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830,
         n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840,
         n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850,
         n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860,
         n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870,
         n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880,
         n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890,
         n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900,
         n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910,
         n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920,
         n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930,
         n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940,
         n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950,
         n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960,
         n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970,
         n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980,
         n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990,
         n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000,
         n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010,
         n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020,
         n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030,
         n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040,
         n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050,
         n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060,
         n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070,
         n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080,
         n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090,
         n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100,
         n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110,
         n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120,
         n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130,
         n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140,
         n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150,
         n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160,
         n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170,
         n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180,
         n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190,
         n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200,
         n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210,
         n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220,
         n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230,
         n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240,
         n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250,
         n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260,
         n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270,
         n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280,
         n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290,
         n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300,
         n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310,
         n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320,
         n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330,
         n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340,
         n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350,
         n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360,
         n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370,
         n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380,
         n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390,
         n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400,
         n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410,
         n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420,
         n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430,
         n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440,
         n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450,
         n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460,
         n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470,
         n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480,
         n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490,
         n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500,
         n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510,
         n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520,
         n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530,
         n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540,
         n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550,
         n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560,
         n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570,
         n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580,
         n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590,
         n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600,
         n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610,
         n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620,
         n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630,
         n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640,
         n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650,
         n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660,
         n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670,
         n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680,
         n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690,
         n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700,
         n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710,
         n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720,
         n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730,
         n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740,
         n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750,
         n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760,
         n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770,
         n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780,
         n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790,
         n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800,
         n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810,
         n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820,
         n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830,
         n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840,
         n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850,
         n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860,
         n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870,
         n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880,
         n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890,
         n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900,
         n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910,
         n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920,
         n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930,
         n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940,
         n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950,
         n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960,
         n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970,
         n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980,
         n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990,
         n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000,
         n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010,
         n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020,
         n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030,
         n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040,
         n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050,
         n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060,
         n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070,
         n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080,
         n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090,
         n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100,
         n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110,
         n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120,
         n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130,
         n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140,
         n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150,
         n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160,
         n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170,
         n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180,
         n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190,
         n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200,
         n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210,
         n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220,
         n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230,
         n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240,
         n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250,
         n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260,
         n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270,
         n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280,
         n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290,
         n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300,
         n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310,
         n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320,
         n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330,
         n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340,
         n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350,
         n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360,
         n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370,
         n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380,
         n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390,
         n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400,
         n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410,
         n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420,
         n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430,
         n8431, n8432, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441,
         n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451,
         n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461,
         n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471,
         n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481,
         n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491,
         n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501,
         n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511,
         n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521,
         n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531,
         n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541,
         n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551,
         n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561,
         n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571,
         n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581,
         n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591,
         n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601,
         n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611,
         n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621,
         n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631,
         n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641,
         n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651,
         n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661,
         n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671,
         n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681,
         n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691,
         n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701,
         n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711,
         n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721,
         n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731,
         n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741,
         n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751,
         n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761,
         n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771,
         n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781,
         n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791,
         n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801,
         n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811,
         n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821,
         n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831,
         n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841,
         n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851,
         n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861,
         n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871,
         n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881,
         n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891,
         n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901,
         n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911,
         n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921,
         n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931,
         n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941,
         n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951,
         n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961,
         n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971,
         n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981,
         n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991,
         n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001,
         n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011,
         n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021,
         n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031,
         n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041,
         n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051,
         n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061,
         n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071,
         n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081,
         n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091,
         n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101,
         n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111,
         n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121,
         n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131,
         n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141,
         n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151,
         n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161,
         n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171,
         n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181,
         n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191,
         n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201,
         n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211,
         n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221,
         n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231,
         n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241,
         n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251,
         n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261,
         n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271,
         n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281,
         n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291,
         n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301,
         n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311,
         n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321,
         n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331,
         n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341,
         n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351,
         n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361,
         n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371,
         n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381,
         n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391,
         n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401,
         n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411,
         n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421,
         n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431,
         n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441,
         n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451,
         n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461,
         n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471,
         n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481,
         n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491,
         n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501,
         n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511,
         n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521,
         n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531,
         n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541,
         n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551,
         n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561,
         n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571,
         n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581,
         n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591,
         n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601,
         n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611,
         n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621,
         n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631,
         n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641,
         n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651,
         n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661,
         n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671,
         n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681,
         n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691,
         n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701,
         n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711,
         n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721,
         n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731,
         n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741,
         n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751,
         n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761,
         n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771,
         n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781,
         n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791,
         n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801,
         n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811,
         n9812, n9813, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
         n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
         n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
         n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
         n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
         n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
         n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
         n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
         n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
         n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
         n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
         n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
         n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
         n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
         n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
         n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
         n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
         n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
         n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
         n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
         n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193,
         n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
         n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209,
         n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217,
         n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
         n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233,
         n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
         n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
         n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
         n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265,
         n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273,
         n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281,
         n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289,
         n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297,
         n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305,
         n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313,
         n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321,
         n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329,
         n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337,
         n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345,
         n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353,
         n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361,
         n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369,
         n10370, n10371, n10372;

  NAND2_X1 U4917 ( .A1(n8254), .A2(n8256), .ZN(n7531) );
  INV_X1 U4918 ( .A(n5308), .ZN(n6639) );
  NAND4_X2 U4919 ( .A1(n5134), .A2(n5133), .A3(n5132), .A4(n5131), .ZN(n6427)
         );
  INV_X2 U4920 ( .A(n5763), .ZN(n8202) );
  BUF_X2 U4921 ( .A(n7197), .Z(n4412) );
  CLKBUF_X2 U4922 ( .A(n5757), .Z(n8208) );
  BUF_X1 U4923 ( .A(n6428), .Z(n9087) );
  AOI21_X1 U4924 ( .B1(n8035), .B2(n4647), .A(n4645), .ZN(n8879) );
  INV_X1 U4925 ( .A(n6424), .ZN(n9085) );
  INV_X2 U4926 ( .A(n5797), .ZN(n6061) );
  OR2_X1 U4927 ( .A1(n6125), .A2(n5715), .ZN(n5717) );
  INV_X1 U4929 ( .A(n5154), .ZN(n6635) );
  INV_X1 U4930 ( .A(n7191), .ZN(n6440) );
  XNOR2_X1 U4931 ( .A(n8170), .B(n8169), .ZN(n8460) );
  INV_X1 U4932 ( .A(n8443), .ZN(n8580) );
  INV_X1 U4933 ( .A(n4412), .ZN(n6195) );
  XOR2_X1 U4934 ( .A(n6453), .B(n6574), .Z(n4411) );
  CLKBUF_X3 U4935 ( .A(n9103), .Z(n4417) );
  OAI21_X2 U4936 ( .B1(n8536), .B2(n8532), .A(n8533), .ZN(n8170) );
  INV_X2 U4937 ( .A(n7175), .ZN(n6411) );
  XNOR2_X2 U4938 ( .A(n5717), .B(n5716), .ZN(n6106) );
  NOR3_X2 U4939 ( .A1(n5378), .A2(n4755), .A3(n5580), .ZN(n5610) );
  NAND2_X2 U4940 ( .A1(n5330), .A2(n4921), .ZN(n5378) );
  XNOR2_X2 U4941 ( .A(n5421), .B(n5114), .ZN(n7648) );
  INV_X2 U4942 ( .A(n5882), .ZN(n7880) );
  OAI22_X2 U4943 ( .A1(n7880), .A2(n5894), .B1(n8585), .B2(n10014), .ZN(n8035)
         );
  OR2_X1 U4944 ( .A1(n6395), .A2(n8190), .ZN(n8397) );
  NAND2_X1 U4945 ( .A1(n7953), .A2(n5327), .ZN(n8099) );
  NAND2_X1 U4946 ( .A1(n6514), .A2(n6517), .ZN(n9050) );
  INV_X2 U4947 ( .A(n8182), .ZN(n8186) );
  INV_X1 U4948 ( .A(n8278), .ZN(n9990) );
  NAND2_X1 U4949 ( .A1(n6420), .A2(n6424), .ZN(n6428) );
  INV_X1 U4950 ( .A(n9264), .ZN(n7406) );
  CLKBUF_X1 U4952 ( .A(n5665), .Z(n4418) );
  NAND2_X2 U4953 ( .A1(n5737), .A2(n6915), .ZN(n5764) );
  BUF_X4 U4954 ( .A(n5144), .Z(n4413) );
  XNOR2_X1 U4955 ( .A(n5586), .B(n10290), .ZN(n8128) );
  AND2_X1 U4956 ( .A1(n5688), .A2(n4989), .ZN(n5689) );
  AND2_X1 U4957 ( .A1(n5659), .A2(n5658), .ZN(n5660) );
  NOR2_X1 U4958 ( .A1(n9653), .A2(n9652), .ZN(n9654) );
  AND2_X1 U4959 ( .A1(n5677), .A2(n5674), .ZN(n5685) );
  XNOR2_X1 U4960 ( .A(n8203), .B(n4568), .ZN(n8755) );
  NAND2_X1 U4961 ( .A1(n9221), .A2(n6583), .ZN(n9222) );
  NAND2_X1 U4962 ( .A1(n5571), .A2(n5570), .ZN(n6821) );
  NAND2_X1 U4963 ( .A1(n9445), .A2(n5525), .ZN(n4903) );
  NAND2_X1 U4964 ( .A1(n5569), .A2(n6625), .ZN(n9821) );
  OR2_X1 U4965 ( .A1(n5568), .A2(SI_29_), .ZN(n5569) );
  OR2_X1 U4966 ( .A1(n4443), .A2(n4781), .ZN(n4780) );
  XNOR2_X1 U4967 ( .A(n6623), .B(n6621), .ZN(n5568) );
  NAND2_X1 U4968 ( .A1(n9516), .A2(n9517), .ZN(n9515) );
  NOR2_X1 U4969 ( .A1(n8721), .A2(n8720), .ZN(n8719) );
  INV_X1 U4970 ( .A(n4722), .ZN(n9516) );
  NAND2_X1 U4971 ( .A1(n9235), .A2(n9234), .ZN(n9233) );
  OAI21_X1 U4972 ( .B1(n9544), .B2(n6707), .A(n6667), .ZN(n4722) );
  AND2_X1 U4973 ( .A1(n4754), .A2(n6521), .ZN(n9235) );
  OR2_X1 U4974 ( .A1(n6520), .A2(n6519), .ZN(n4754) );
  OAI21_X1 U4975 ( .B1(n8099), .B2(n4907), .A(n4905), .ZN(n4904) );
  NAND2_X1 U4976 ( .A1(n4708), .A2(n4463), .ZN(n9590) );
  NAND2_X1 U4977 ( .A1(n7855), .A2(n7856), .ZN(n7957) );
  NOR2_X1 U4978 ( .A1(n8621), .A2(n6336), .ZN(n6337) );
  OAI21_X1 U4979 ( .B1(n7684), .B2(n6163), .A(n8303), .ZN(n7805) );
  NAND2_X1 U4980 ( .A1(n9105), .A2(n4975), .ZN(n7174) );
  OAI21_X1 U4981 ( .B1(n7431), .B2(n6157), .A(n6158), .ZN(n7515) );
  AOI21_X1 U4982 ( .B1(n7311), .B2(n8606), .A(n8607), .ZN(n8610) );
  OR2_X1 U4983 ( .A1(n8588), .A2(n9994), .ZN(n8303) );
  AND2_X2 U4984 ( .A1(n6361), .A2(n9943), .ZN(n9960) );
  AND2_X1 U4985 ( .A1(n5835), .A2(n5834), .ZN(n9994) );
  NAND2_X2 U4986 ( .A1(n5673), .A2(n9886), .ZN(n9560) );
  NAND2_X1 U4987 ( .A1(n4562), .A2(n4559), .ZN(n5068) );
  BUF_X2 U4988 ( .A(n6508), .Z(n6587) );
  OR2_X1 U4989 ( .A1(n5772), .A2(n9972), .ZN(n8261) );
  NAND3_X1 U4990 ( .A1(n6408), .A2(n6404), .A3(n6403), .ZN(n6420) );
  NAND2_X2 U4991 ( .A1(n8250), .A2(n8425), .ZN(n8402) );
  NAND4_X1 U4992 ( .A1(n5731), .A2(n5730), .A3(n5729), .A4(n5728), .ZN(n7537)
         );
  INV_X1 U4993 ( .A(n5740), .ZN(n9961) );
  NAND4_X1 U4994 ( .A1(n5171), .A2(n5170), .A3(n5169), .A4(n5168), .ZN(n9263)
         );
  NAND4_X1 U4995 ( .A1(n5150), .A2(n5149), .A3(n5148), .A4(n5147), .ZN(n9264)
         );
  NAND4_X1 U4996 ( .A1(n5762), .A2(n5761), .A3(n5760), .A4(n5759), .ZN(n5772)
         );
  INV_X1 U4997 ( .A(n5369), .ZN(n5146) );
  INV_X2 U4998 ( .A(n5155), .ZN(n5535) );
  INV_X1 U4999 ( .A(n5764), .ZN(n8201) );
  NAND2_X1 U5000 ( .A1(n5021), .A2(n9820), .ZN(n5308) );
  XNOR2_X1 U5001 ( .A(n5593), .B(P1_IR_REG_21__SCAN_IN), .ZN(n5665) );
  NAND2_X1 U5002 ( .A1(n5597), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5593) );
  NAND2_X1 U5003 ( .A1(n9048), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5702) );
  NAND2_X1 U5004 ( .A1(n5597), .A2(n5596), .ZN(n7667) );
  NAND2_X2 U5005 ( .A1(n6106), .A2(n6290), .ZN(n5737) );
  INV_X1 U5006 ( .A(n9820), .ZN(n5023) );
  XNOR2_X1 U5007 ( .A(n5720), .B(n5719), .ZN(n6290) );
  XNOR2_X1 U5008 ( .A(n5121), .B(P1_IR_REG_27__SCAN_IN), .ZN(n5650) );
  OAI21_X1 U5009 ( .B1(n5121), .B2(n5118), .A(n5117), .ZN(n5120) );
  XNOR2_X1 U5010 ( .A(n5020), .B(n5019), .ZN(n9820) );
  XNOR2_X1 U5011 ( .A(n5594), .B(P1_IR_REG_22__SCAN_IN), .ZN(n6843) );
  NAND2_X1 U5012 ( .A1(n5749), .A2(n5748), .ZN(n7021) );
  NAND2_X1 U5013 ( .A1(n5806), .A2(n5807), .ZN(n5820) );
  NOR2_X1 U5014 ( .A1(n5013), .A2(n4688), .ZN(n4920) );
  AND3_X1 U5015 ( .A1(n5722), .A2(n4674), .A3(n4673), .ZN(n5806) );
  NAND2_X2 U5016 ( .A1(n4850), .A2(n4848), .ZN(n5122) );
  AND2_X1 U5017 ( .A1(n5008), .A2(n5009), .ZN(n4921) );
  NAND2_X1 U5018 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(n5015), .ZN(n5117) );
  NAND2_X1 U5019 ( .A1(n4994), .A2(P1_IR_REG_28__SCAN_IN), .ZN(n5118) );
  AND2_X1 U5020 ( .A1(n5692), .A2(n4937), .ZN(n4673) );
  AND2_X1 U5021 ( .A1(n5691), .A2(n5693), .ZN(n4674) );
  INV_X1 U5022 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n5612) );
  NOR2_X2 U5023 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n5173) );
  INV_X1 U5024 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n5393) );
  INV_X1 U5025 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5392) );
  INV_X4 U5026 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  NOR2_X1 U5027 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n5007) );
  INV_X1 U5028 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n5265) );
  INV_X1 U5029 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5579) );
  INV_X1 U5030 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n4852) );
  INV_X1 U5031 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4851) );
  INV_X1 U5032 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n5264) );
  INV_X1 U5033 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5977) );
  NOR2_X2 U5034 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5722) );
  INV_X4 U5035 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  NAND2_X1 U5036 ( .A1(n6873), .A2(n5732), .ZN(n4414) );
  NAND2_X1 U5037 ( .A1(n6873), .A2(n5732), .ZN(n5155) );
  OAI21_X2 U5038 ( .B1(n6186), .B2(n8386), .A(n8388), .ZN(n6380) );
  NAND2_X1 U5039 ( .A1(n6873), .A2(n6915), .ZN(n4415) );
  NAND2_X1 U5040 ( .A1(n6873), .A2(n6915), .ZN(n5154) );
  AOI22_X2 U5041 ( .A1(n9508), .A2(n5636), .B1(n9499), .B2(n9689), .ZN(n9493)
         );
  OAI22_X2 U5042 ( .A1(n9522), .A2(n5434), .B1(n9545), .B2(n9696), .ZN(n9508)
         );
  NAND2_X1 U5043 ( .A1(n6420), .A2(n6424), .ZN(n4416) );
  OAI21_X2 U5044 ( .B1(n9515), .B2(n6797), .A(n4718), .ZN(n9461) );
  OAI211_X1 U5045 ( .C1(n6873), .C2(n6916), .A(n5129), .B(n5128), .ZN(n9103)
         );
  AOI21_X2 U5046 ( .B1(n7624), .B2(n7620), .A(n7622), .ZN(n7836) );
  NAND2_X1 U5047 ( .A1(n5021), .A2(n5023), .ZN(n5144) );
  OAI22_X2 U5048 ( .A1(n4742), .A2(n7363), .B1(n4411), .B2(n7524), .ZN(n7609)
         );
  NOR2_X2 U5049 ( .A1(n7364), .A2(n7365), .ZN(n7363) );
  OAI22_X2 U5050 ( .A1(n7253), .A2(n7252), .B1(n6446), .B2(n6445), .ZN(n7364)
         );
  AOI21_X2 U5051 ( .B1(n7836), .B2(n6483), .A(n6482), .ZN(n7909) );
  XNOR2_X1 U5052 ( .A(n6447), .B(n6574), .ZN(n6449) );
  INV_X4 U5053 ( .A(n9085), .ZN(n6574) );
  NAND2_X2 U5054 ( .A1(n6408), .A2(n5667), .ZN(n6418) );
  NAND2_X2 U5055 ( .A1(n5608), .A2(n4723), .ZN(n6408) );
  NAND2_X1 U5056 ( .A1(n8364), .A2(n8362), .ZN(n4549) );
  NOR2_X1 U5057 ( .A1(P2_IR_REG_14__SCAN_IN), .A2(P2_IR_REG_9__SCAN_IN), .ZN(
        n5695) );
  OAI21_X1 U5058 ( .B1(n4880), .B2(n4424), .A(n5077), .ZN(n4877) );
  OR2_X1 U5059 ( .A1(n9031), .A2(n8565), .ZN(n8350) );
  INV_X1 U5060 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n5692) );
  OR2_X1 U5061 ( .A1(n6842), .A2(n6843), .ZN(n6404) );
  OAI21_X1 U5062 ( .B1(n5122), .B2(P1_DATAO_REG_4__SCAN_IN), .A(n4565), .ZN(
        n5047) );
  NAND2_X1 U5063 ( .A1(n5122), .A2(n6932), .ZN(n4565) );
  NAND2_X1 U5064 ( .A1(n8311), .A2(n8402), .ZN(n4571) );
  NAND2_X1 U5065 ( .A1(n8310), .A2(n8406), .ZN(n4572) );
  OAI22_X1 U5066 ( .A1(n4638), .A2(n6825), .B1(n4634), .B2(n6837), .ZN(n4631)
         );
  OR2_X1 U5067 ( .A1(n6737), .A2(n6738), .ZN(n4638) );
  NAND2_X1 U5068 ( .A1(n4636), .A2(n4635), .ZN(n4634) );
  NAND2_X1 U5069 ( .A1(n6733), .A2(n4627), .ZN(n4629) );
  NAND2_X1 U5070 ( .A1(n4633), .A2(n4632), .ZN(n4627) );
  NAND2_X1 U5071 ( .A1(n4471), .A2(n6837), .ZN(n4633) );
  NAND2_X1 U5072 ( .A1(n4540), .A2(n4451), .ZN(n4539) );
  NAND2_X1 U5073 ( .A1(n4542), .A2(n4541), .ZN(n4540) );
  NAND2_X1 U5074 ( .A1(n4573), .A2(n8345), .ZN(n8353) );
  NAND2_X1 U5075 ( .A1(n4575), .A2(n4574), .ZN(n4573) );
  AOI21_X1 U5076 ( .B1(n4548), .B2(n4550), .A(n8369), .ZN(n4547) );
  INV_X1 U5077 ( .A(n8364), .ZN(n4550) );
  NAND2_X1 U5078 ( .A1(n4569), .A2(n8390), .ZN(n8393) );
  OR4_X1 U5079 ( .A1(n6810), .A2(n6848), .A3(n6809), .A4(n6825), .ZN(n6815) );
  NOR2_X1 U5080 ( .A1(n5094), .A2(n4886), .ZN(n4885) );
  INV_X1 U5081 ( .A(n5092), .ZN(n4886) );
  INV_X1 U5082 ( .A(n5349), .ZN(n5091) );
  INV_X1 U5083 ( .A(SI_15_), .ZN(n5090) );
  NOR2_X1 U5084 ( .A1(n4971), .A2(n7282), .ZN(n4968) );
  NOR2_X1 U5085 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .ZN(
        n5697) );
  NOR2_X1 U5086 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), .ZN(
        n5696) );
  NOR2_X1 U5087 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n5694) );
  XNOR2_X1 U5088 ( .A(n5706), .B(P2_IR_REG_29__SCAN_IN), .ZN(n5708) );
  NAND2_X1 U5089 ( .A1(n4532), .A2(n4531), .ZN(n4530) );
  NOR2_X1 U5090 ( .A1(n6216), .A2(n6218), .ZN(n4531) );
  NOR2_X1 U5091 ( .A1(n7769), .A2(n6331), .ZN(n6332) );
  AND2_X1 U5092 ( .A1(n6943), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n6331) );
  OR2_X1 U5093 ( .A1(n8183), .A2(n8561), .ZN(n8388) );
  XNOR2_X1 U5094 ( .A(n8192), .B(n8580), .ZN(n8235) );
  OR2_X1 U5095 ( .A1(n4431), .A2(n4487), .ZN(n4670) );
  AND2_X1 U5096 ( .A1(n6172), .A2(n8819), .ZN(n8784) );
  AND2_X1 U5097 ( .A1(n4788), .A2(n8355), .ZN(n4783) );
  OR2_X1 U5098 ( .A1(n8956), .A2(n8509), .ZN(n8354) );
  INV_X1 U5099 ( .A(n5908), .ZN(n4657) );
  AND2_X1 U5100 ( .A1(n6115), .A2(n4979), .ZN(n5718) );
  OR2_X1 U5101 ( .A1(P2_IR_REG_27__SCAN_IN), .A2(P2_IR_REG_26__SCAN_IN), .ZN(
        n5701) );
  INV_X1 U5102 ( .A(n5713), .ZN(n5714) );
  INV_X1 U5103 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n6093) );
  INV_X1 U5104 ( .A(n6092), .ZN(n6096) );
  INV_X1 U5105 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n4937) );
  INV_X1 U5106 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n5691) );
  NOR2_X1 U5107 ( .A1(n9565), .A2(n9703), .ZN(n9550) );
  NAND2_X1 U5108 ( .A1(n5567), .A2(n5566), .ZN(n6623) );
  INV_X1 U5109 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5004) );
  INV_X1 U5110 ( .A(n4921), .ZN(n4688) );
  NAND2_X1 U5111 ( .A1(n4756), .A2(n5581), .ZN(n4755) );
  INV_X1 U5112 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5581) );
  INV_X1 U5113 ( .A(n4757), .ZN(n4756) );
  AOI21_X1 U5114 ( .B1(n4868), .B2(n4865), .A(n4508), .ZN(n4864) );
  OAI21_X1 U5115 ( .B1(n5391), .B2(n5106), .A(n5105), .ZN(n5403) );
  NAND2_X1 U5116 ( .A1(n5088), .A2(n5087), .ZN(n5348) );
  NAND2_X1 U5117 ( .A1(n4875), .A2(n4873), .ZN(n5315) );
  AOI21_X1 U5118 ( .B1(n4876), .B2(n4874), .A(n4477), .ZN(n4873) );
  NOR2_X1 U5119 ( .A1(n4877), .A2(n5080), .ZN(n4871) );
  INV_X1 U5120 ( .A(n4560), .ZN(n4559) );
  OAI21_X1 U5121 ( .B1(n4563), .B2(n4561), .A(n4995), .ZN(n4560) );
  INV_X1 U5122 ( .A(n5062), .ZN(n4561) );
  NAND3_X1 U5123 ( .A1(n4849), .A2(P1_ADDR_REG_19__SCAN_IN), .A3(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n4848) );
  NAND3_X1 U5124 ( .A1(n5032), .A2(n4852), .A3(n4851), .ZN(n4850) );
  INV_X1 U5125 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4849) );
  OAI21_X1 U5126 ( .B1(n4440), .B2(n4952), .A(n4951), .ZN(n4950) );
  AND2_X1 U5127 ( .A1(n8439), .A2(n8185), .ZN(n4952) );
  NAND2_X1 U5128 ( .A1(n4440), .A2(n8185), .ZN(n4951) );
  INV_X1 U5129 ( .A(n5756), .ZN(n6101) );
  AND4_X1 U5130 ( .A1(n5946), .A2(n5945), .A3(n5944), .A4(n5943), .ZN(n8565)
         );
  XNOR2_X1 U5131 ( .A(n6219), .B(n6320), .ZN(n7128) );
  NAND2_X1 U5132 ( .A1(n4530), .A2(n4527), .ZN(n6219) );
  INV_X1 U5133 ( .A(n4529), .ZN(n4527) );
  AND2_X1 U5134 ( .A1(n4530), .A2(n4528), .ZN(n6220) );
  NOR2_X1 U5135 ( .A1(n4529), .A2(n6320), .ZN(n4528) );
  NAND2_X1 U5136 ( .A1(n4835), .A2(n4833), .ZN(n4523) );
  AND2_X1 U5137 ( .A1(n4834), .A2(n4510), .ZN(n4833) );
  NAND2_X1 U5138 ( .A1(n4664), .A2(n4661), .ZN(n6187) );
  AOI21_X1 U5139 ( .B1(n4663), .B2(n4666), .A(n4662), .ZN(n4661) );
  NOR2_X1 U5140 ( .A1(n8178), .A2(n6067), .ZN(n4662) );
  OR2_X1 U5141 ( .A1(n8952), .A2(n8868), .ZN(n8358) );
  INV_X1 U5142 ( .A(n8585), .ZN(n8087) );
  INV_X1 U5144 ( .A(n8907), .ZN(n9951) );
  OR2_X1 U5145 ( .A1(n10014), .A2(n8087), .ZN(n8323) );
  NAND2_X1 U5146 ( .A1(n5737), .A2(n5732), .ZN(n5763) );
  XNOR2_X1 U5147 ( .A(n5780), .B(P2_IR_REG_4__SCAN_IN), .ZN(n6316) );
  AOI22_X1 U5148 ( .A1(n4416), .A2(n7191), .B1(n6508), .B2(n9263), .ZN(n6443)
         );
  NOR2_X1 U5149 ( .A1(n9752), .A2(n9394), .ZN(n6857) );
  AND2_X1 U5150 ( .A1(n9752), .A2(n9394), .ZN(n6839) );
  NOR2_X1 U5151 ( .A1(n5607), .A2(n8128), .ZN(n4723) );
  NAND2_X1 U5152 ( .A1(n4903), .A2(n4901), .ZN(n4899) );
  AND2_X1 U5153 ( .A1(n4902), .A2(n5526), .ZN(n4901) );
  OR2_X1 U5154 ( .A1(n9509), .A2(n9499), .ZN(n6659) );
  OR2_X1 U5155 ( .A1(n9210), .A2(n9255), .ZN(n5294) );
  NAND2_X1 U5156 ( .A1(n4890), .A2(n4888), .ZN(n7590) );
  AND2_X1 U5157 ( .A1(n4889), .A2(n7591), .ZN(n4888) );
  NAND2_X1 U5158 ( .A1(n4891), .A2(n4893), .ZN(n4889) );
  OR2_X1 U5159 ( .A1(n9263), .A2(n7191), .ZN(n5172) );
  INV_X1 U5160 ( .A(n6427), .ZN(n7087) );
  INV_X1 U5161 ( .A(n4904), .ZN(n9599) );
  AOI21_X1 U5162 ( .B1(n9618), .B2(n4906), .A(n5374), .ZN(n4905) );
  NAND2_X1 U5163 ( .A1(n9618), .A2(n4911), .ZN(n4907) );
  INV_X1 U5164 ( .A(n5737), .ZN(n6209) );
  INV_X1 U5165 ( .A(n8806), .ZN(n8777) );
  OR2_X1 U5166 ( .A1(n9821), .A2(n5154), .ZN(n5571) );
  NAND2_X1 U5167 ( .A1(n8321), .A2(n8406), .ZN(n4542) );
  NAND2_X1 U5168 ( .A1(n8316), .A2(n8315), .ZN(n8320) );
  NOR2_X1 U5169 ( .A1(n4631), .A2(n6740), .ZN(n4628) );
  NAND2_X1 U5170 ( .A1(n4600), .A2(n4599), .ZN(n4598) );
  NOR2_X1 U5171 ( .A1(n8102), .A2(n6746), .ZN(n4599) );
  NAND2_X1 U5172 ( .A1(n4601), .A2(n8100), .ZN(n4600) );
  NAND2_X1 U5173 ( .A1(n4547), .A2(n4434), .ZN(n4544) );
  OAI21_X1 U5174 ( .B1(n6803), .B2(n6802), .A(n4613), .ZN(n4612) );
  AND2_X1 U5175 ( .A1(n9476), .A2(n6801), .ZN(n4613) );
  NAND2_X1 U5176 ( .A1(n6807), .A2(n4610), .ZN(n4609) );
  AND2_X1 U5177 ( .A1(n6806), .A2(n6819), .ZN(n4610) );
  NAND2_X1 U5178 ( .A1(n4679), .A2(n9658), .ZN(n4678) );
  NAND2_X1 U5179 ( .A1(n4709), .A2(n4713), .ZN(n4708) );
  INV_X1 U5180 ( .A(n4711), .ZN(n4710) );
  OAI21_X1 U5181 ( .B1(n9623), .B2(n4712), .A(n6655), .ZN(n4711) );
  NOR2_X1 U5182 ( .A1(n9739), .A2(n9059), .ZN(n4692) );
  INV_X1 U5183 ( .A(n5361), .ZN(n5093) );
  NOR2_X1 U5184 ( .A1(n4412), .A2(n7199), .ZN(n7200) );
  INV_X1 U5185 ( .A(n8405), .ZN(n4795) );
  NOR2_X1 U5186 ( .A1(n4796), .A2(n4792), .ZN(n4791) );
  INV_X1 U5187 ( .A(n6381), .ZN(n4792) );
  INV_X1 U5188 ( .A(n8397), .ZN(n4796) );
  NAND2_X1 U5189 ( .A1(n4526), .A2(n4459), .ZN(n4824) );
  NAND2_X1 U5190 ( .A1(n4824), .A2(n7054), .ZN(n4825) );
  NAND2_X1 U5191 ( .A1(n6315), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n4816) );
  NAND3_X1 U5192 ( .A1(n4811), .A2(n4809), .A3(n4455), .ZN(n6323) );
  INV_X1 U5193 ( .A(n8383), .ZN(n4779) );
  INV_X1 U5194 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n8018) );
  NAND2_X1 U5195 ( .A1(n5813), .A2(n5812), .ZN(n5827) );
  INV_X1 U5196 ( .A(n5814), .ZN(n5813) );
  INV_X1 U5197 ( .A(n8284), .ZN(n4770) );
  AND2_X1 U5198 ( .A1(n8285), .A2(n8248), .ZN(n6161) );
  NAND2_X1 U5199 ( .A1(n7269), .A2(n5753), .ZN(n8260) );
  NAND2_X1 U5200 ( .A1(n8254), .A2(n7532), .ZN(n8251) );
  AND2_X1 U5201 ( .A1(n8406), .A2(n7198), .ZN(n7100) );
  INV_X1 U5202 ( .A(n8340), .ZN(n4786) );
  NAND2_X1 U5203 ( .A1(n5949), .A2(n4650), .ZN(n4646) );
  INV_X1 U5204 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5719) );
  NOR2_X1 U5205 ( .A1(n6123), .A2(P2_IR_REG_26__SCAN_IN), .ZN(n6125) );
  INV_X1 U5206 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n5963) );
  AOI21_X1 U5207 ( .B1(n6556), .B2(n4731), .A(n9177), .ZN(n4729) );
  INV_X1 U5208 ( .A(n9062), .ZN(n4747) );
  OR2_X1 U5209 ( .A1(n9809), .A2(n5606), .ZN(n6598) );
  MUX2_X1 U5210 ( .A(n6828), .B(n6837), .S(n9401), .Z(n6829) );
  OR2_X1 U5211 ( .A1(n4425), .A2(n4625), .ZN(n4620) );
  OAI21_X1 U5212 ( .B1(n6817), .B2(n4619), .A(n4618), .ZN(n6827) );
  INV_X1 U5213 ( .A(n4621), .ZN(n4619) );
  AOI21_X1 U5214 ( .B1(n4624), .B2(n4621), .A(n4432), .ZN(n4618) );
  NOR2_X1 U5215 ( .A1(n4425), .A2(n4622), .ZN(n4621) );
  INV_X1 U5216 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n10082) );
  OR2_X1 U5217 ( .A1(n9323), .A2(n4594), .ZN(n4593) );
  AND2_X1 U5218 ( .A1(n9324), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n4594) );
  NOR2_X1 U5219 ( .A1(n6821), .A2(n4678), .ZN(n4677) );
  OR2_X1 U5220 ( .A1(n9649), .A2(n9432), .ZN(n6818) );
  NAND2_X1 U5221 ( .A1(n9658), .A2(n9441), .ZN(n4902) );
  NOR2_X1 U5222 ( .A1(n9450), .A2(n9764), .ZN(n9423) );
  OR2_X1 U5223 ( .A1(n9465), .A2(n9478), .ZN(n9437) );
  NOR2_X1 U5224 ( .A1(n9496), .A2(n4721), .ZN(n4720) );
  INV_X1 U5225 ( .A(n6659), .ZN(n4721) );
  NOR2_X1 U5226 ( .A1(n9801), .A2(n4691), .ZN(n4690) );
  INV_X1 U5227 ( .A(n4692), .ZN(n4691) );
  OR2_X1 U5228 ( .A1(n9210), .A2(n7981), .ZN(n6741) );
  OR2_X1 U5229 ( .A1(n9173), .A2(n7439), .ZN(n6739) );
  OR2_X1 U5230 ( .A1(n9424), .A2(n9441), .ZN(n6819) );
  AND2_X1 U5231 ( .A1(n9801), .A2(n9722), .ZN(n5374) );
  OR2_X1 U5232 ( .A1(n9801), .A2(n9607), .ZN(n6767) );
  AND2_X1 U5233 ( .A1(n5589), .A2(n9810), .ZN(n6599) );
  INV_X1 U5234 ( .A(n7667), .ZN(n6678) );
  AND2_X1 U5235 ( .A1(n5508), .A2(n5494), .ZN(n5506) );
  AND2_X1 U5236 ( .A1(n5489), .A2(n5476), .ZN(n5487) );
  NAND2_X1 U5237 ( .A1(n4478), .A2(n4990), .ZN(n5580) );
  AOI21_X1 U5238 ( .B1(n4509), .B2(n5419), .A(n4869), .ZN(n4868) );
  NOR2_X1 U5239 ( .A1(n5112), .A2(SI_20_), .ZN(n4869) );
  INV_X1 U5240 ( .A(n5375), .ZN(n4882) );
  INV_X1 U5241 ( .A(n5071), .ZN(n4878) );
  INV_X1 U5242 ( .A(n4877), .ZN(n4876) );
  NOR2_X1 U5243 ( .A1(n5263), .A2(n4881), .ZN(n4558) );
  INV_X1 U5244 ( .A(n4558), .ZN(n4556) );
  NAND2_X1 U5245 ( .A1(n5058), .A2(n5057), .ZN(n5235) );
  INV_X1 U5246 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n4591) );
  INV_X1 U5247 ( .A(n8481), .ZN(n4934) );
  OR2_X1 U5248 ( .A1(n4442), .A2(n8505), .ZN(n4964) );
  OR2_X1 U5249 ( .A1(n5827), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5839) );
  NAND2_X1 U5250 ( .A1(n7789), .A2(n4940), .ZN(n4939) );
  INV_X1 U5251 ( .A(n7778), .ZN(n4940) );
  AND2_X1 U5252 ( .A1(n4942), .A2(n7671), .ZN(n4941) );
  INV_X1 U5253 ( .A(n7669), .ZN(n4942) );
  NOR2_X1 U5254 ( .A1(n4934), .A2(n4930), .ZN(n4929) );
  INV_X1 U5255 ( .A(n8523), .ZN(n4930) );
  AOI21_X1 U5256 ( .B1(n4974), .B2(n4981), .A(n4426), .ZN(n4966) );
  NOR2_X1 U5257 ( .A1(n7573), .A2(n7574), .ZN(n7670) );
  OR2_X1 U5258 ( .A1(n8515), .A2(n4927), .ZN(n4926) );
  INV_X1 U5259 ( .A(n8175), .ZN(n4927) );
  NAND2_X1 U5260 ( .A1(n4978), .A2(n4959), .ZN(n4958) );
  NOR2_X1 U5261 ( .A1(n5700), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n4959) );
  AND2_X1 U5262 ( .A1(n8212), .A2(n6105), .ZN(n8190) );
  NAND2_X1 U5263 ( .A1(n5796), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n5745) );
  OR2_X1 U5264 ( .A1(n5774), .A2(n6257), .ZN(n5711) );
  NAND2_X1 U5265 ( .A1(n6151), .A2(n6150), .ZN(n7098) );
  AND2_X1 U5266 ( .A1(n6149), .A2(n6148), .ZN(n6150) );
  NAND2_X1 U5267 ( .A1(n7021), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6312) );
  OR2_X1 U5268 ( .A1(n7027), .A2(n7026), .ZN(n4526) );
  NAND2_X1 U5269 ( .A1(n4825), .A2(n4823), .ZN(n7058) );
  NAND2_X1 U5270 ( .A1(n6215), .A2(n6313), .ZN(n4823) );
  INV_X1 U5271 ( .A(n4824), .ZN(n6215) );
  INV_X1 U5272 ( .A(n4825), .ZN(n6216) );
  INV_X1 U5273 ( .A(n9923), .ZN(n4533) );
  NOR2_X1 U5274 ( .A1(n7058), .A2(n5758), .ZN(n7057) );
  OAI21_X1 U5275 ( .B1(n7128), .B2(n4839), .A(n4838), .ZN(n7238) );
  NAND2_X1 U5276 ( .A1(n4842), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n4839) );
  INV_X1 U5277 ( .A(n7239), .ZN(n4842) );
  OR2_X1 U5278 ( .A1(n7128), .A2(n5787), .ZN(n4841) );
  NAND2_X1 U5279 ( .A1(n6321), .A2(n4810), .ZN(n4809) );
  INV_X1 U5280 ( .A(n7244), .ZN(n4810) );
  OR2_X1 U5281 ( .A1(n7130), .A2(n4812), .ZN(n4811) );
  OR2_X1 U5282 ( .A1(n7244), .A2(n7517), .ZN(n4812) );
  OR2_X1 U5283 ( .A1(n7130), .A2(n7517), .ZN(n4814) );
  OR2_X1 U5284 ( .A1(n8604), .A2(n6227), .ZN(n6228) );
  XNOR2_X1 U5285 ( .A(n6228), .B(n6939), .ZN(n7658) );
  NAND2_X1 U5286 ( .A1(n4819), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n4818) );
  NAND2_X1 U5287 ( .A1(n6329), .A2(n4819), .ZN(n4817) );
  INV_X1 U5288 ( .A(n7770), .ZN(n4819) );
  AOI21_X1 U5289 ( .B1(P2_REG1_REG_12__SCAN_IN), .B2(n6953), .A(n8615), .ZN(
        n6233) );
  NAND2_X1 U5290 ( .A1(n4828), .A2(n4827), .ZN(n4525) );
  NAND2_X1 U5291 ( .A1(n6237), .A2(n4832), .ZN(n4827) );
  OR2_X1 U5292 ( .A1(n8667), .A2(n4829), .ZN(n4828) );
  NAND2_X1 U5293 ( .A1(n4832), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n4829) );
  NOR2_X1 U5294 ( .A1(n4525), .A2(n4524), .ZN(n6238) );
  NOR2_X1 U5295 ( .A1(n8688), .A2(n8962), .ZN(n4524) );
  AOI21_X1 U5296 ( .B1(P2_REG2_REG_16__SCAN_IN), .B2(n7164), .A(n8683), .ZN(
        n6343) );
  NOR2_X1 U5297 ( .A1(n8443), .A2(n9953), .ZN(n6189) );
  NAND2_X1 U5298 ( .A1(n8388), .A2(n8389), .ZN(n8386) );
  OR2_X1 U5299 ( .A1(n6023), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6036) );
  OR2_X1 U5300 ( .A1(n6014), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6023) );
  NAND2_X1 U5301 ( .A1(n8852), .A2(n4460), .ZN(n8837) );
  INV_X1 U5302 ( .A(n8842), .ZN(n6000) );
  AND2_X1 U5303 ( .A1(n8365), .A2(n8828), .ZN(n8842) );
  AND3_X1 U5304 ( .A1(n5999), .A2(n5998), .A3(n5997), .ZN(n8856) );
  NAND2_X1 U5305 ( .A1(n4659), .A2(n8853), .ZN(n8852) );
  OR2_X1 U5306 ( .A1(n5918), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5931) );
  AOI21_X1 U5307 ( .B1(n4421), .B2(n4774), .A(n4773), .ZN(n4772) );
  AND2_X1 U5308 ( .A1(n8323), .A2(n8324), .ZN(n7879) );
  OR2_X1 U5309 ( .A1(n5868), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5887) );
  OR2_X1 U5310 ( .A1(n5853), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5868) );
  NAND2_X1 U5311 ( .A1(n4776), .A2(n8225), .ZN(n4775) );
  INV_X1 U5312 ( .A(n7805), .ZN(n4776) );
  AND2_X1 U5313 ( .A1(n8315), .A2(n8307), .ZN(n8224) );
  AND2_X1 U5314 ( .A1(n8299), .A2(n8306), .ZN(n8225) );
  OR2_X1 U5315 ( .A1(n5799), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5814) );
  OAI21_X1 U5316 ( .B1(n7515), .B2(n7512), .A(n7511), .ZN(n7565) );
  NAND2_X1 U5317 ( .A1(n7428), .A2(n8284), .ZN(n7514) );
  NAND2_X1 U5318 ( .A1(n5727), .A2(n5726), .ZN(n5740) );
  AND2_X1 U5319 ( .A1(n4492), .A2(n5725), .ZN(n5727) );
  OR2_X1 U5320 ( .A1(n7537), .A2(n7206), .ZN(n7532) );
  AOI22_X1 U5321 ( .A1(n6187), .A2(n8386), .B1(n8768), .B2(n8183), .ZN(n6373)
         );
  OR2_X1 U5322 ( .A1(n8383), .A2(n8384), .ZN(n8766) );
  AOI21_X1 U5323 ( .B1(n4669), .B2(n6044), .A(n4436), .ZN(n4666) );
  NOR2_X1 U5324 ( .A1(n6175), .A2(n8243), .ZN(n4781) );
  INV_X1 U5325 ( .A(n8766), .ZN(n8764) );
  OR2_X1 U5326 ( .A1(n8991), .A2(n8777), .ZN(n8786) );
  NAND2_X1 U5327 ( .A1(n6171), .A2(n8242), .ZN(n8783) );
  AOI21_X1 U5328 ( .B1(n4799), .B2(n8853), .A(n4798), .ZN(n4797) );
  INV_X1 U5329 ( .A(n8363), .ZN(n4798) );
  NAND2_X1 U5330 ( .A1(n6003), .A2(n6002), .ZN(n8478) );
  NAND2_X1 U5331 ( .A1(n5992), .A2(n5991), .ZN(n8521) );
  NAND2_X1 U5332 ( .A1(n8858), .A2(n8857), .ZN(n8860) );
  NOR2_X1 U5333 ( .A1(n6167), .A2(n4789), .ZN(n4788) );
  INV_X1 U5334 ( .A(n8338), .ZN(n4789) );
  INV_X1 U5335 ( .A(n8341), .ZN(n8880) );
  NAND2_X1 U5336 ( .A1(n8406), .A2(n7212), .ZN(n9953) );
  OR2_X1 U5337 ( .A1(n8904), .A2(n8216), .ZN(n6166) );
  INV_X1 U5338 ( .A(n4653), .ZN(n4652) );
  OAI21_X1 U5339 ( .B1(n5924), .B2(n4654), .A(n4658), .ZN(n4653) );
  NAND2_X1 U5340 ( .A1(n5909), .A2(n5908), .ZN(n4654) );
  NAND2_X1 U5341 ( .A1(n8035), .A2(n4655), .ZN(n4651) );
  NAND2_X1 U5342 ( .A1(n4758), .A2(n4760), .ZN(n8904) );
  AOI21_X1 U5343 ( .B1(n8334), .B2(n8329), .A(n4761), .ZN(n4760) );
  NAND2_X1 U5344 ( .A1(n6165), .A2(n4759), .ZN(n4758) );
  INV_X1 U5345 ( .A(n8335), .ZN(n4761) );
  INV_X1 U5346 ( .A(n8330), .ZN(n4765) );
  AND2_X1 U5347 ( .A1(n6109), .A2(n8406), .ZN(n8907) );
  AND3_X1 U5348 ( .A1(n5770), .A2(n5769), .A3(n5768), .ZN(n9972) );
  AND3_X1 U5349 ( .A1(n5752), .A2(n5751), .A3(n5750), .ZN(n9966) );
  NAND2_X1 U5350 ( .A1(n6099), .A2(n6194), .ZN(n8912) );
  NAND2_X1 U5351 ( .A1(n6128), .A2(n6148), .ZN(n6132) );
  NAND2_X1 U5352 ( .A1(n5718), .A2(n5719), .ZN(n5704) );
  NAND2_X1 U5353 ( .A1(n5704), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5706) );
  INV_X1 U5354 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n10121) );
  NAND2_X1 U5355 ( .A1(n6117), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6119) );
  INV_X1 U5356 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n6118) );
  NOR2_X1 U5357 ( .A1(n5975), .A2(P2_IR_REG_18__SCAN_IN), .ZN(n6091) );
  AND2_X1 U5358 ( .A1(n5925), .A2(n5915), .ZN(n8656) );
  NOR2_X1 U5359 ( .A1(n5849), .A2(P2_IR_REG_9__SCAN_IN), .ZN(n5861) );
  INV_X1 U5360 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5860) );
  XNOR2_X1 U5361 ( .A(n5793), .B(P2_IR_REG_5__SCAN_IN), .ZN(n6320) );
  NOR2_X1 U5362 ( .A1(n5748), .A2(n4936), .ZN(n5792) );
  NAND2_X1 U5363 ( .A1(n4937), .A2(n5692), .ZN(n4936) );
  INV_X1 U5364 ( .A(n5748), .ZN(n4935) );
  NAND2_X1 U5365 ( .A1(n5722), .A2(n5691), .ZN(n5748) );
  NAND2_X1 U5366 ( .A1(n4750), .A2(n9187), .ZN(n4749) );
  INV_X1 U5367 ( .A(n6562), .ZN(n4750) );
  NAND2_X1 U5368 ( .A1(n6562), .A2(n4753), .ZN(n4752) );
  INV_X1 U5369 ( .A(n9187), .ZN(n4753) );
  INV_X1 U5370 ( .A(n7363), .ZN(n4740) );
  NOR2_X1 U5371 ( .A1(n4992), .A2(n4411), .ZN(n4739) );
  AND3_X1 U5372 ( .A1(n6600), .A2(n6599), .A3(n6598), .ZN(n6617) );
  AOI21_X1 U5373 ( .B1(n9756), .B2(n9249), .A(n6857), .ZN(n6684) );
  XNOR2_X1 U5374 ( .A(n4593), .B(n9338), .ZN(n9325) );
  OAI21_X1 U5375 ( .B1(n9861), .B2(n4596), .A(n9867), .ZN(n9367) );
  OR2_X1 U5376 ( .A1(n9370), .A2(n9369), .ZN(n4577) );
  NAND2_X1 U5377 ( .A1(n4457), .A2(n4902), .ZN(n4900) );
  INV_X1 U5378 ( .A(n9532), .ZN(n9499) );
  AND2_X1 U5379 ( .A1(n9515), .A2(n4720), .ZN(n9494) );
  NAND2_X1 U5380 ( .A1(n8050), .A2(n6766), .ZN(n9622) );
  NAND2_X1 U5381 ( .A1(n9622), .A2(n9623), .ZN(n9621) );
  NAND2_X1 U5382 ( .A1(n4703), .A2(n4701), .ZN(n8050) );
  NOR2_X1 U5383 ( .A1(n4702), .A2(n8053), .ZN(n4701) );
  INV_X1 U5384 ( .A(n4705), .ZN(n4702) );
  NAND2_X1 U5385 ( .A1(n4704), .A2(n6764), .ZN(n4703) );
  INV_X1 U5386 ( .A(n7957), .ZN(n4704) );
  AOI21_X1 U5387 ( .B1(n6764), .B2(n4707), .A(n4706), .ZN(n4705) );
  INV_X1 U5388 ( .A(n6761), .ZN(n4706) );
  INV_X1 U5389 ( .A(n5635), .ZN(n4707) );
  OR2_X1 U5390 ( .A1(n7821), .A2(n9210), .ZN(n7858) );
  OR2_X1 U5391 ( .A1(n7756), .A2(n9256), .ZN(n5279) );
  INV_X1 U5392 ( .A(n7442), .ZN(n4893) );
  AOI21_X1 U5393 ( .B1(n7442), .B2(n4892), .A(n4465), .ZN(n4891) );
  INV_X1 U5394 ( .A(n5233), .ZN(n4892) );
  NAND3_X1 U5395 ( .A1(n4895), .A2(n4894), .A3(n5219), .ZN(n7414) );
  NAND2_X1 U5396 ( .A1(n4896), .A2(n4898), .ZN(n4894) );
  NAND2_X1 U5397 ( .A1(n6721), .A2(n6713), .ZN(n7180) );
  OR2_X1 U5398 ( .A1(n9876), .A2(n6899), .ZN(n9591) );
  INV_X1 U5399 ( .A(n9893), .ZN(n9498) );
  OR2_X1 U5400 ( .A1(n9567), .A2(n4519), .ZN(n6605) );
  AND2_X1 U5401 ( .A1(n5616), .A2(n9811), .ZN(n6600) );
  OR2_X1 U5402 ( .A1(n9809), .A2(P1_D_REG_0__SCAN_IN), .ZN(n5616) );
  NAND2_X1 U5403 ( .A1(n9764), .A2(n5524), .ZN(n5525) );
  INV_X1 U5404 ( .A(n9469), .ZN(n9668) );
  INV_X1 U5405 ( .A(n5636), .ZN(n9517) );
  NAND2_X1 U5406 ( .A1(n5401), .A2(n4917), .ZN(n4916) );
  NOR2_X1 U5407 ( .A1(n4470), .A2(n4918), .ZN(n4917) );
  INV_X1 U5408 ( .A(n4984), .ZN(n4918) );
  INV_X1 U5409 ( .A(n9526), .ZN(n9543) );
  AOI21_X1 U5410 ( .B1(n4911), .B2(n4909), .A(n4466), .ZN(n4908) );
  INV_X1 U5411 ( .A(n5347), .ZN(n4909) );
  OR2_X1 U5412 ( .A1(n9744), .A2(n9253), .ZN(n5327) );
  INV_X1 U5413 ( .A(n6873), .ZN(n5406) );
  INV_X1 U5414 ( .A(n4897), .ZN(n4896) );
  OAI21_X1 U5415 ( .B1(n7488), .B2(n4898), .A(n7334), .ZN(n4897) );
  INV_X1 U5416 ( .A(n5002), .ZN(n4898) );
  NAND2_X1 U5417 ( .A1(n7489), .A2(n7488), .ZN(n7487) );
  INV_X1 U5418 ( .A(n9899), .ZN(n9745) );
  INV_X1 U5419 ( .A(n9723), .ZN(n9705) );
  NAND2_X1 U5420 ( .A1(n6408), .A2(n5664), .ZN(n9807) );
  NAND2_X1 U5421 ( .A1(n6625), .A2(n6624), .ZN(n6630) );
  INV_X1 U5422 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n5019) );
  NAND2_X1 U5423 ( .A1(n5568), .A2(SI_29_), .ZN(n6625) );
  AND2_X1 U5424 ( .A1(n5297), .A2(n4614), .ZN(n4616) );
  NOR2_X1 U5425 ( .A1(n5016), .A2(n4615), .ZN(n4614) );
  INV_X1 U5426 ( .A(n5007), .ZN(n4615) );
  NAND2_X1 U5427 ( .A1(n4726), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4725) );
  NAND2_X1 U5428 ( .A1(n4883), .A2(n4884), .ZN(n5376) );
  NAND2_X1 U5429 ( .A1(n4887), .A2(n5092), .ZN(n5363) );
  NAND2_X1 U5430 ( .A1(n4879), .A2(n5071), .ZN(n5281) );
  AND2_X1 U5431 ( .A1(n5176), .A2(n5163), .ZN(n4855) );
  NAND2_X1 U5432 ( .A1(n4564), .A2(n4467), .ZN(n4698) );
  NAND2_X1 U5433 ( .A1(n4857), .A2(n5176), .ZN(n4564) );
  XNOR2_X1 U5434 ( .A(n5047), .B(SI_4_), .ZN(n5176) );
  NOR2_X1 U5435 ( .A1(n4947), .A2(n8571), .ZN(n4945) );
  AND2_X1 U5436 ( .A1(n4950), .A2(n4490), .ZN(n4947) );
  INV_X1 U5437 ( .A(n8185), .ZN(n4949) );
  NAND2_X1 U5438 ( .A1(n4950), .A2(n4953), .ZN(n4948) );
  NAND2_X1 U5439 ( .A1(n4440), .A2(n4954), .ZN(n4953) );
  INV_X1 U5440 ( .A(n8439), .ZN(n4954) );
  AND4_X1 U5441 ( .A1(n5845), .A2(n5844), .A3(n5843), .A4(n5842), .ZN(n7991)
         );
  AND4_X1 U5442 ( .A1(n5989), .A2(n5988), .A3(n5987), .A4(n5986), .ZN(n8868)
         );
  AND2_X1 U5443 ( .A1(n6079), .A2(n6078), .ZN(n8561) );
  NAND2_X1 U5444 ( .A1(n7120), .A2(n9943), .ZN(n8576) );
  INV_X1 U5445 ( .A(n7545), .ZN(n8420) );
  INV_X1 U5446 ( .A(n8561), .ZN(n8768) );
  NAND2_X1 U5447 ( .A1(n6043), .A2(n6042), .ZN(n8806) );
  INV_X1 U5448 ( .A(n8827), .ZN(n8807) );
  INV_X1 U5449 ( .A(n8565), .ZN(n8910) );
  NAND2_X1 U5450 ( .A1(n4520), .A2(n7933), .ZN(n4521) );
  OR2_X1 U5451 ( .A1(n8634), .A2(n5898), .ZN(n4846) );
  OR2_X1 U5452 ( .A1(n8667), .A2(n8965), .ZN(n4831) );
  INV_X1 U5453 ( .A(n4807), .ZN(n8671) );
  NAND2_X1 U5454 ( .A1(n4804), .A2(n4803), .ZN(n8683) );
  NAND2_X1 U5455 ( .A1(n6341), .A2(n4808), .ZN(n4803) );
  OR2_X1 U5456 ( .A1(n8672), .A2(n4805), .ZN(n4804) );
  NAND2_X1 U5457 ( .A1(n4808), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n4805) );
  INV_X1 U5458 ( .A(n7248), .ZN(n9918) );
  NAND2_X1 U5459 ( .A1(n5885), .A2(n5884), .ZN(n10014) );
  NAND2_X1 U5460 ( .A1(n6356), .A2(n7109), .ZN(n9943) );
  INV_X2 U5461 ( .A(n9960), .ZN(n8913) );
  INV_X1 U5462 ( .A(n8950), .ZN(n8966) );
  NOR2_X1 U5463 ( .A1(n8749), .A2(n6394), .ZN(n6402) );
  AND2_X1 U5464 ( .A1(n6393), .A2(n6392), .ZN(n6394) );
  NAND2_X1 U5465 ( .A1(n5897), .A2(n5896), .ZN(n8096) );
  XNOR2_X1 U5466 ( .A(n5911), .B(P2_IR_REG_13__SCAN_IN), .ZN(n8643) );
  NAND2_X1 U5467 ( .A1(n4738), .A2(n4498), .ZN(n9102) );
  NAND2_X1 U5468 ( .A1(n6494), .A2(n4977), .ZN(n6495) );
  NAND2_X1 U5469 ( .A1(n5124), .A2(n5123), .ZN(n9703) );
  NAND2_X1 U5470 ( .A1(n5444), .A2(n5443), .ZN(n9509) );
  INV_X1 U5471 ( .A(n9247), .ZN(n9209) );
  OR2_X1 U5472 ( .A1(n5308), .A2(n5130), .ZN(n5132) );
  OR2_X1 U5473 ( .A1(n5446), .A2(n7394), .ZN(n5133) );
  NAND2_X1 U5474 ( .A1(n9828), .A2(n9827), .ZN(n9826) );
  OR2_X1 U5475 ( .A1(n6992), .A2(n6993), .ZN(n4588) );
  NAND2_X1 U5476 ( .A1(n4588), .A2(n4587), .ZN(n4586) );
  NAND2_X1 U5477 ( .A1(n7068), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n4587) );
  AND2_X1 U5478 ( .A1(n4586), .A2(n4585), .ZN(n7289) );
  INV_X1 U5479 ( .A(n7069), .ZN(n4585) );
  INV_X1 U5480 ( .A(n9722), .ZN(n9607) );
  AND2_X1 U5481 ( .A1(n9560), .A2(n5669), .ZN(n9446) );
  AND2_X1 U5482 ( .A1(n9560), .A2(n5670), .ZN(n9620) );
  OR2_X1 U5483 ( .A1(n6605), .A2(n9807), .ZN(n9886) );
  AND2_X1 U5484 ( .A1(n6638), .A2(n6637), .ZN(n9752) );
  XNOR2_X1 U5485 ( .A(n5577), .B(n6824), .ZN(n5684) );
  INV_X1 U5486 ( .A(n6734), .ZN(n4636) );
  INV_X1 U5487 ( .A(n7585), .ZN(n4635) );
  NAND2_X1 U5488 ( .A1(n4637), .A2(n6825), .ZN(n4632) );
  NOR2_X1 U5489 ( .A1(n6734), .A2(n7413), .ZN(n4637) );
  AOI21_X1 U5490 ( .B1(n8322), .B2(n8402), .A(n8327), .ZN(n4541) );
  INV_X1 U5491 ( .A(n4631), .ZN(n4630) );
  AND2_X1 U5492 ( .A1(n8880), .A2(n4485), .ZN(n4574) );
  NAND2_X1 U5493 ( .A1(n4602), .A2(n7956), .ZN(n4601) );
  NAND2_X1 U5494 ( .A1(n4639), .A2(n7812), .ZN(n6742) );
  NAND2_X1 U5495 ( .A1(n4538), .A2(n8336), .ZN(n8337) );
  NAND2_X1 U5496 ( .A1(n4539), .A2(n8333), .ZN(n4538) );
  INV_X1 U5497 ( .A(n8359), .ZN(n4552) );
  NOR2_X1 U5498 ( .A1(n4606), .A2(n6837), .ZN(n4605) );
  INV_X1 U5499 ( .A(n6782), .ZN(n4606) );
  OAI211_X1 U5500 ( .C1(n6773), .C2(n6825), .A(n9608), .B(n4607), .ZN(n6785)
         );
  OR2_X1 U5501 ( .A1(n6772), .A2(n6837), .ZN(n4607) );
  AOI21_X1 U5502 ( .B1(n4598), .B2(n6749), .A(n6748), .ZN(n6750) );
  AOI21_X1 U5503 ( .B1(n4547), .B2(n4546), .A(n4473), .ZN(n4545) );
  INV_X1 U5504 ( .A(n4548), .ZN(n4546) );
  NAND2_X1 U5505 ( .A1(n8382), .A2(n8764), .ZN(n4570) );
  OAI21_X1 U5506 ( .B1(n6805), .B2(n6825), .A(n4608), .ZN(n6816) );
  AOI21_X1 U5507 ( .B1(n4612), .B2(n4611), .A(n4609), .ZN(n4608) );
  NOR2_X1 U5508 ( .A1(n6837), .A2(n6661), .ZN(n4611) );
  NOR2_X1 U5509 ( .A1(n8393), .A2(n4566), .ZN(n8407) );
  NAND2_X1 U5510 ( .A1(n4568), .A2(n4567), .ZN(n4566) );
  OR2_X1 U5511 ( .A1(n6132), .A2(n6147), .ZN(n7094) );
  INV_X1 U5512 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n6114) );
  NAND2_X1 U5513 ( .A1(n4626), .A2(n9401), .ZN(n4622) );
  NAND2_X1 U5514 ( .A1(n5272), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5305) );
  NAND2_X1 U5515 ( .A1(n7583), .A2(n6739), .ZN(n6734) );
  AND2_X1 U5516 ( .A1(n4868), .A2(n4867), .ZN(n4862) );
  INV_X1 U5517 ( .A(n5437), .ZN(n4867) );
  NOR2_X1 U5518 ( .A1(n4866), .A2(n5437), .ZN(n4865) );
  INV_X1 U5519 ( .A(n4870), .ZN(n4866) );
  INV_X1 U5520 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n5102) );
  INV_X1 U5521 ( .A(SI_17_), .ZN(n5096) );
  INV_X1 U5522 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n5009) );
  AND2_X1 U5523 ( .A1(n4424), .A2(n5295), .ZN(n4874) );
  INV_X1 U5524 ( .A(n7571), .ZN(n4973) );
  INV_X1 U5525 ( .A(n7572), .ZN(n4974) );
  NOR2_X1 U5526 ( .A1(n4533), .A2(n6218), .ZN(n4529) );
  NOR2_X1 U5527 ( .A1(n8627), .A2(n6335), .ZN(n6336) );
  INV_X1 U5528 ( .A(n8692), .ZN(n4832) );
  INV_X1 U5529 ( .A(n6068), .ZN(n4665) );
  NOR2_X1 U5530 ( .A1(n4669), .A2(n6068), .ZN(n4663) );
  INV_X1 U5531 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n10087) );
  OR2_X1 U5532 ( .A1(n5941), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5955) );
  INV_X1 U5533 ( .A(n8313), .ZN(n4773) );
  INV_X1 U5534 ( .A(n8225), .ZN(n4774) );
  INV_X1 U5535 ( .A(n9966), .ZN(n5753) );
  OR2_X1 U5536 ( .A1(n8985), .A2(n8176), .ZN(n8379) );
  NOR2_X1 U5537 ( .A1(n4764), .A2(n4762), .ZN(n4759) );
  INV_X1 U5538 ( .A(n8334), .ZN(n4762) );
  NAND2_X1 U5539 ( .A1(n7094), .A2(n7109), .ZN(n6200) );
  INV_X1 U5540 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n10253) );
  NAND2_X1 U5541 ( .A1(n4978), .A2(n4957), .ZN(n4956) );
  OR2_X1 U5542 ( .A1(n5863), .A2(P2_IR_REG_11__SCAN_IN), .ZN(n5895) );
  OAI21_X1 U5543 ( .B1(n7885), .B2(n4737), .A(n4736), .ZN(n6513) );
  AOI21_X1 U5544 ( .B1(n6500), .B2(n7971), .A(n4472), .ZN(n4736) );
  INV_X1 U5545 ( .A(n7971), .ZN(n4737) );
  AND2_X1 U5546 ( .A1(P1_REG3_REG_19__SCAN_IN), .A2(n5024), .ZN(n5025) );
  NAND2_X1 U5547 ( .A1(n9127), .A2(n4445), .ZN(n4730) );
  NOR2_X1 U5548 ( .A1(n5340), .A2(n5339), .ZN(n5338) );
  NAND2_X1 U5549 ( .A1(n6673), .A2(n9405), .ZN(n6848) );
  INV_X1 U5550 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n10209) );
  INV_X1 U5551 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5008) );
  INV_X1 U5552 ( .A(n4678), .ZN(n4676) );
  NOR2_X1 U5553 ( .A1(n9685), .A2(n4685), .ZN(n4684) );
  INV_X1 U5554 ( .A(n4686), .ZN(n4685) );
  NOR2_X1 U5555 ( .A1(n9696), .A2(n9509), .ZN(n4686) );
  NOR2_X1 U5556 ( .A1(n9143), .A2(n9141), .ZN(n5397) );
  OR2_X1 U5557 ( .A1(n5305), .A2(n5304), .ZN(n5321) );
  NOR2_X1 U5558 ( .A1(n7858), .A2(n7889), .ZN(n7859) );
  NOR2_X1 U5559 ( .A1(n5255), .A2(n10209), .ZN(n5254) );
  OAI21_X1 U5560 ( .B1(n6734), .B2(n7585), .A(n6751), .ZN(n5629) );
  OR2_X1 U5561 ( .A1(n4716), .A2(n6734), .ZN(n6692) );
  NAND2_X1 U5562 ( .A1(n6720), .A2(n6735), .ZN(n4716) );
  INV_X1 U5563 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n5240) );
  OR2_X1 U5564 ( .A1(n5241), .A2(n5240), .ZN(n5255) );
  NAND2_X1 U5565 ( .A1(n7362), .A2(n9262), .ZN(n6722) );
  NAND2_X1 U5566 ( .A1(n4708), .A2(n4710), .ZN(n9588) );
  INV_X1 U5567 ( .A(n9587), .ZN(n4715) );
  INV_X1 U5568 ( .A(n4908), .ZN(n4906) );
  NAND2_X1 U5569 ( .A1(n8106), .A2(n4692), .ZN(n9627) );
  NOR2_X1 U5570 ( .A1(n7593), .A2(n9173), .ZN(n7744) );
  NOR2_X1 U5571 ( .A1(n7221), .A2(n7322), .ZN(n7490) );
  NAND2_X1 U5572 ( .A1(n4675), .A2(n6440), .ZN(n7221) );
  NAND2_X1 U5573 ( .A1(n4991), .A2(n5015), .ZN(n5016) );
  AND2_X1 U5574 ( .A1(n5547), .A2(n5534), .ZN(n5545) );
  AND2_X1 U5575 ( .A1(n5529), .A2(n5513), .ZN(n5527) );
  NAND2_X1 U5576 ( .A1(n5377), .A2(n5392), .ZN(n4757) );
  AOI21_X1 U5577 ( .B1(n4885), .B2(n5089), .A(n4479), .ZN(n4884) );
  NOR2_X1 U5578 ( .A1(n5072), .A2(n4881), .ZN(n4880) );
  INV_X1 U5579 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5003) );
  INV_X1 U5580 ( .A(n5046), .ZN(n4857) );
  OAI21_X1 U5581 ( .B1(n5122), .B2(P1_DATAO_REG_2__SCAN_IN), .A(n5039), .ZN(
        n5040) );
  NAND2_X1 U5582 ( .A1(n5122), .A2(n6924), .ZN(n5039) );
  NAND2_X1 U5583 ( .A1(n4694), .A2(n4693), .ZN(n5035) );
  NAND2_X1 U5584 ( .A1(n5122), .A2(n6918), .ZN(n4693) );
  NAND2_X1 U5585 ( .A1(n4696), .A2(n4695), .ZN(n4694) );
  OR2_X1 U5586 ( .A1(n8010), .A2(n8064), .ZN(n8013) );
  NAND2_X1 U5587 ( .A1(n7278), .A2(n5772), .ZN(n7279) );
  NAND2_X1 U5588 ( .A1(n5982), .A2(n5981), .ZN(n5995) );
  INV_X1 U5589 ( .A(n5983), .ZN(n5982) );
  AOI21_X1 U5590 ( .B1(n4419), .B2(n4427), .A(n4963), .ZN(n4962) );
  NAND2_X1 U5591 ( .A1(n5954), .A2(n5953), .ZN(n5968) );
  INV_X1 U5592 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n5953) );
  INV_X1 U5593 ( .A(n5955), .ZN(n5954) );
  NAND2_X1 U5594 ( .A1(n5930), .A2(n5929), .ZN(n5941) );
  INV_X1 U5595 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n5929) );
  INV_X1 U5596 ( .A(n5931), .ZN(n5930) );
  INV_X1 U5597 ( .A(n4794), .ZN(n4793) );
  OAI211_X1 U5598 ( .C1(n8748), .C2(n8923), .A(n8415), .B(n4795), .ZN(n4794)
         );
  NAND2_X1 U5599 ( .A1(n4480), .A2(n5723), .ZN(n4802) );
  OAI21_X1 U5600 ( .B1(n6977), .B2(n6211), .A(n6212), .ZN(n6974) );
  INV_X1 U5601 ( .A(n4816), .ZN(n4815) );
  AND2_X1 U5602 ( .A1(n4422), .A2(n4816), .ZN(n9927) );
  INV_X1 U5603 ( .A(n4841), .ZN(n7127) );
  INV_X1 U5604 ( .A(n6323), .ZN(n6325) );
  NAND2_X1 U5605 ( .A1(n6222), .A2(n4505), .ZN(n6223) );
  INV_X1 U5606 ( .A(n7238), .ZN(n6222) );
  NAND2_X1 U5607 ( .A1(n6323), .A2(n7310), .ZN(n8606) );
  AOI21_X1 U5608 ( .B1(P2_REG2_REG_8__SCAN_IN), .B2(n8598), .A(n8610), .ZN(
        n6328) );
  NAND2_X1 U5609 ( .A1(n4836), .A2(n4439), .ZN(n4835) );
  INV_X1 U5610 ( .A(n7658), .ZN(n4836) );
  AND2_X1 U5611 ( .A1(n6333), .A2(n6948), .ZN(n6334) );
  NOR2_X1 U5612 ( .A1(n8639), .A2(n5903), .ZN(n8638) );
  OAI21_X1 U5613 ( .B1(n8639), .B2(n4821), .A(n4820), .ZN(n8658) );
  NAND2_X1 U5614 ( .A1(n4822), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n4821) );
  NAND2_X1 U5615 ( .A1(n6338), .A2(n4822), .ZN(n4820) );
  INV_X1 U5616 ( .A(n8659), .ZN(n4822) );
  INV_X1 U5617 ( .A(n8684), .ZN(n4808) );
  INV_X1 U5618 ( .A(n9938), .ZN(n8709) );
  AND2_X1 U5619 ( .A1(n8705), .A2(n8883), .ZN(n8706) );
  INV_X1 U5620 ( .A(n6100), .ZN(n8743) );
  NAND2_X1 U5621 ( .A1(n8401), .A2(n8443), .ZN(n6374) );
  AND2_X1 U5622 ( .A1(n4780), .A2(n4779), .ZN(n4778) );
  OR2_X1 U5623 ( .A1(n6171), .A2(n4443), .ZN(n4777) );
  OR2_X1 U5624 ( .A1(n6058), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n6073) );
  NAND2_X1 U5625 ( .A1(n6035), .A2(n6034), .ZN(n6049) );
  INV_X1 U5626 ( .A(n6036), .ZN(n6035) );
  NAND2_X1 U5627 ( .A1(n6004), .A2(n10087), .ZN(n6014) );
  INV_X1 U5628 ( .A(n6005), .ZN(n6004) );
  INV_X1 U5629 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n5899) );
  INV_X1 U5630 ( .A(n5901), .ZN(n5900) );
  NAND2_X1 U5631 ( .A1(n5886), .A2(n8018), .ZN(n5901) );
  INV_X1 U5632 ( .A(n5887), .ZN(n5886) );
  INV_X1 U5633 ( .A(n5839), .ZN(n5838) );
  AOI21_X1 U5634 ( .B1(n4642), .B2(n4644), .A(n4448), .ZN(n4640) );
  INV_X1 U5635 ( .A(n4643), .ZN(n4642) );
  OAI21_X1 U5636 ( .B1(n7553), .B2(n4644), .A(n8221), .ZN(n4643) );
  INV_X1 U5637 ( .A(n5825), .ZN(n4644) );
  NAND2_X1 U5638 ( .A1(n7549), .A2(n5825), .ZN(n7686) );
  NAND2_X1 U5639 ( .A1(n7550), .A2(n7553), .ZN(n7549) );
  NAND2_X1 U5640 ( .A1(n4770), .A2(n8287), .ZN(n4769) );
  INV_X1 U5641 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5783) );
  NAND2_X1 U5642 ( .A1(n7375), .A2(n5773), .ZN(n7431) );
  AND2_X1 U5643 ( .A1(n8251), .A2(n8256), .ZN(n9941) );
  NOR2_X1 U5644 ( .A1(n6200), .A2(n7100), .ZN(n6355) );
  OR2_X1 U5645 ( .A1(n6199), .A2(n6137), .ZN(n6354) );
  AND2_X1 U5646 ( .A1(n8742), .A2(n8741), .ZN(n8970) );
  INV_X1 U5647 ( .A(n8235), .ZN(n6090) );
  NAND2_X1 U5648 ( .A1(n6070), .A2(n6069), .ZN(n8183) );
  OR2_X1 U5649 ( .A1(n5764), .A2(n8197), .ZN(n6069) );
  AND2_X1 U5650 ( .A1(n8379), .A2(n8380), .ZN(n8774) );
  AOI21_X1 U5651 ( .B1(n4786), .B2(n8355), .A(n4785), .ZN(n4784) );
  INV_X1 U5652 ( .A(n8342), .ZN(n4785) );
  NOR2_X1 U5653 ( .A1(n4648), .A2(n4656), .ZN(n4647) );
  NAND2_X1 U5654 ( .A1(n4481), .A2(n4646), .ZN(n4645) );
  INV_X1 U5655 ( .A(n5949), .ZN(n4648) );
  NAND2_X1 U5656 ( .A1(n4651), .A2(n4649), .ZN(n8891) );
  OAI21_X1 U5657 ( .B1(n8035), .B2(n5909), .A(n5908), .ZN(n8026) );
  OR2_X1 U5658 ( .A1(n6201), .A2(n8425), .ZN(n10000) );
  INV_X1 U5659 ( .A(n10005), .ZN(n10015) );
  INV_X1 U5660 ( .A(n9970), .ZN(n10010) );
  NOR2_X1 U5661 ( .A1(n7104), .A2(n6200), .ZN(n7119) );
  AND2_X1 U5662 ( .A1(n7114), .A2(n9944), .ZN(n7101) );
  OR2_X1 U5663 ( .A1(n7095), .A2(n6200), .ZN(n7121) );
  INV_X1 U5664 ( .A(n7535), .ZN(n7206) );
  AND2_X1 U5665 ( .A1(n7098), .A2(n8135), .ZN(n7109) );
  INV_X1 U5666 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5716) );
  AND2_X1 U5667 ( .A1(n6127), .A2(n6126), .ZN(n6148) );
  NAND2_X1 U5668 ( .A1(n6094), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6095) );
  INV_X1 U5669 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5693) );
  MUX2_X1 U5670 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5721), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n5724) );
  NAND2_X1 U5671 ( .A1(n9911), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5721) );
  NAND2_X1 U5672 ( .A1(n6425), .A2(n9085), .ZN(n6426) );
  INV_X1 U5673 ( .A(n4729), .ZN(n4727) );
  INV_X1 U5674 ( .A(n9127), .ZN(n4728) );
  INV_X1 U5675 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n9141) );
  AOI21_X1 U5676 ( .B1(n4430), .B2(n4751), .A(n4747), .ZN(n4746) );
  INV_X1 U5677 ( .A(n4752), .ZN(n4751) );
  NAND2_X1 U5678 ( .A1(n5445), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n5462) );
  AND2_X1 U5679 ( .A1(n5425), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n5445) );
  NAND2_X1 U5680 ( .A1(n6448), .A2(n6427), .ZN(n6432) );
  OR2_X1 U5681 ( .A1(n7158), .A2(n6418), .ZN(n6433) );
  XNOR2_X1 U5682 ( .A(n6431), .B(n9085), .ZN(n6434) );
  AOI22_X1 U5683 ( .A1(n6428), .A2(n7175), .B1(n6508), .B2(n9264), .ZN(n6410)
         );
  INV_X1 U5684 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n5211) );
  NAND2_X1 U5685 ( .A1(n4744), .A2(n4743), .ZN(n4742) );
  NAND2_X1 U5686 ( .A1(n4411), .A2(n7524), .ZN(n4743) );
  INV_X1 U5687 ( .A(n4992), .ZN(n4744) );
  NAND3_X1 U5688 ( .A1(n6831), .A2(n6832), .A3(n6830), .ZN(n6836) );
  NOR4_X1 U5689 ( .A1(n6706), .A2(n6839), .A3(n6705), .A4(n6704), .ZN(n6861)
         );
  INV_X1 U5690 ( .A(n5664), .ZN(n6871) );
  NOR2_X1 U5691 ( .A1(n6986), .A2(n4582), .ZN(n7042) );
  NOR2_X1 U5692 ( .A1(n6922), .A2(n4583), .ZN(n4582) );
  INV_X1 U5693 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n4583) );
  NOR2_X1 U5694 ( .A1(n7042), .A2(n7041), .ZN(n9841) );
  NOR2_X1 U5695 ( .A1(n7289), .A2(n4584), .ZN(n7347) );
  AND2_X1 U5696 ( .A1(n7296), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n4584) );
  INV_X1 U5697 ( .A(n4593), .ZN(n9344) );
  AND2_X1 U5698 ( .A1(n9423), .A2(n4493), .ZN(n9399) );
  NAND2_X1 U5699 ( .A1(n5537), .A2(n5536), .ZN(n9424) );
  NAND2_X1 U5700 ( .A1(n5496), .A2(n5495), .ZN(n9465) );
  INV_X1 U5701 ( .A(n4719), .ZN(n4718) );
  OAI21_X1 U5702 ( .B1(n6797), .B2(n4720), .A(n6795), .ZN(n4719) );
  AND2_X1 U5703 ( .A1(n9437), .A2(n6668), .ZN(n9460) );
  NAND2_X1 U5704 ( .A1(n9461), .A2(n9460), .ZN(n9459) );
  AND2_X1 U5705 ( .A1(n9550), .A2(n4682), .ZN(n9483) );
  AND2_X1 U5706 ( .A1(n4684), .A2(n4683), .ZN(n4682) );
  NAND2_X1 U5707 ( .A1(n9550), .A2(n4684), .ZN(n9501) );
  AND4_X1 U5708 ( .A1(n5503), .A2(n5502), .A3(n5501), .A4(n5500), .ZN(n9478)
         );
  INV_X1 U5709 ( .A(n9675), .ZN(n9519) );
  NAND2_X1 U5710 ( .A1(n9550), .A2(n9536), .ZN(n9535) );
  AND2_X1 U5711 ( .A1(n9572), .A2(n6777), .ZN(n9544) );
  NAND2_X1 U5712 ( .A1(n9573), .A2(n9574), .ZN(n9572) );
  AND2_X1 U5713 ( .A1(n8106), .A2(n4689), .ZN(n9601) );
  AND2_X1 U5714 ( .A1(n9600), .A2(n4690), .ZN(n4689) );
  AND2_X1 U5715 ( .A1(n7859), .A2(n7979), .ZN(n8106) );
  NAND2_X1 U5716 ( .A1(n8106), .A2(n8115), .ZN(n8105) );
  NAND2_X1 U5717 ( .A1(n7957), .A2(n5635), .ZN(n8101) );
  NAND2_X1 U5718 ( .A1(n7744), .A2(n7915), .ZN(n7821) );
  NAND2_X1 U5719 ( .A1(n4717), .A2(n6692), .ZN(n7738) );
  INV_X1 U5720 ( .A(n5629), .ZN(n4717) );
  AND4_X1 U5721 ( .A1(n5246), .A2(n5245), .A3(n5244), .A4(n5243), .ZN(n7588)
         );
  NAND2_X1 U5722 ( .A1(n4681), .A2(n4680), .ZN(n7593) );
  AND2_X1 U5723 ( .A1(n7490), .A2(n9900), .ZN(n7491) );
  AND2_X1 U5724 ( .A1(n6712), .A2(n5627), .ZN(n7183) );
  INV_X1 U5725 ( .A(n9263), .ZN(n7086) );
  BUF_X1 U5726 ( .A(n5623), .Z(n7152) );
  INV_X1 U5727 ( .A(n9647), .ZN(n9653) );
  INV_X1 U5728 ( .A(n6800), .ZN(n9476) );
  AND2_X1 U5729 ( .A1(n4919), .A2(n4433), .ZN(n4915) );
  OR2_X1 U5730 ( .A1(n9703), .A2(n9695), .ZN(n4919) );
  NAND2_X1 U5731 ( .A1(n9621), .A2(n6770), .ZN(n9609) );
  NAND2_X1 U5732 ( .A1(n5353), .A2(n5352), .ZN(n9739) );
  NAND2_X1 U5733 ( .A1(n5319), .A2(n5318), .ZN(n9744) );
  INV_X1 U5734 ( .A(n9255), .ZN(n7981) );
  AND4_X1 U5735 ( .A1(n5278), .A2(n5277), .A3(n5276), .A4(n5275), .ZN(n7830)
         );
  NAND2_X1 U5736 ( .A1(n7087), .A2(n7158), .ZN(n5141) );
  INV_X1 U5737 ( .A(n6600), .ZN(n5663) );
  AND2_X1 U5738 ( .A1(n5615), .A2(n5662), .ZN(n5683) );
  NAND2_X1 U5739 ( .A1(n5642), .A2(n5641), .ZN(n9893) );
  XNOR2_X1 U5740 ( .A(n6630), .B(n6629), .ZN(n8429) );
  NAND2_X1 U5741 ( .A1(n5586), .A2(n5116), .ZN(n5121) );
  AND2_X1 U5742 ( .A1(n5566), .A2(n5552), .ZN(n5564) );
  XNOR2_X1 U5743 ( .A(n5546), .B(n5545), .ZN(n8194) );
  INV_X1 U5744 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n10290) );
  NAND2_X1 U5745 ( .A1(n5582), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5584) );
  INV_X1 U5746 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5583) );
  NAND2_X1 U5747 ( .A1(n5584), .A2(n5583), .ZN(n4726) );
  AND2_X1 U5748 ( .A1(n5471), .A2(n5458), .ZN(n5469) );
  XNOR2_X1 U5749 ( .A(n5613), .B(n5612), .ZN(n6679) );
  NAND2_X1 U5750 ( .A1(n4863), .A2(n4868), .ZN(n5438) );
  OR2_X1 U5751 ( .A1(n5113), .A2(n4870), .ZN(n4863) );
  NAND2_X1 U5752 ( .A1(n5592), .A2(n5010), .ZN(n5597) );
  NAND2_X1 U5753 ( .A1(n5404), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5405) );
  AND2_X1 U5754 ( .A1(n5301), .A2(n5316), .ZN(n7293) );
  NAND2_X1 U5755 ( .A1(n4872), .A2(n4876), .ZN(n5296) );
  OR2_X1 U5756 ( .A1(n5068), .A2(n4424), .ZN(n4872) );
  NAND3_X1 U5757 ( .A1(n4557), .A2(n4553), .A3(n4555), .ZN(n6942) );
  OR2_X1 U5758 ( .A1(n4559), .A2(n4556), .ZN(n4555) );
  XNOR2_X1 U5759 ( .A(n5247), .B(n4995), .ZN(n6937) );
  OAI21_X1 U5760 ( .B1(n5235), .B2(n5234), .A(n5062), .ZN(n5247) );
  AOI21_X1 U5761 ( .B1(n5190), .B2(n4698), .A(n4476), .ZN(n4697) );
  CLKBUF_X1 U5762 ( .A(n5203), .Z(n5204) );
  XNOR2_X1 U5763 ( .A(n5035), .B(SI_1_), .ZN(n5127) );
  AND3_X1 U5764 ( .A1(n5125), .A2(n4590), .A3(n4589), .ZN(n6905) );
  NAND2_X1 U5765 ( .A1(n4483), .A2(P1_IR_REG_1__SCAN_IN), .ZN(n4589) );
  NAND2_X1 U5766 ( .A1(n4591), .A2(n9815), .ZN(n4590) );
  NAND2_X1 U5767 ( .A1(n4943), .A2(n4941), .ZN(n7779) );
  INV_X1 U5768 ( .A(n7670), .ZN(n4943) );
  NAND2_X1 U5769 ( .A1(n7779), .A2(n7778), .ZN(n7790) );
  AND3_X1 U5770 ( .A1(n6018), .A2(n6017), .A3(n6016), .ZN(n8827) );
  NAND2_X1 U5771 ( .A1(n8514), .A2(n8515), .ZN(n4925) );
  OR2_X1 U5772 ( .A1(n8572), .A2(n4427), .ZN(n4961) );
  INV_X1 U5773 ( .A(n4938), .ZN(n7792) );
  INV_X1 U5774 ( .A(n8568), .ZN(n8550) );
  NAND2_X1 U5775 ( .A1(n4928), .A2(n4932), .ZN(n8536) );
  AOI21_X1 U5776 ( .B1(n8481), .B2(n4933), .A(n4435), .ZN(n4932) );
  NAND2_X1 U5777 ( .A1(n7113), .A2(n7112), .ZN(n8558) );
  AOI21_X1 U5778 ( .B1(n4429), .B2(n4927), .A(n4502), .ZN(n4923) );
  NAND2_X1 U5779 ( .A1(n6029), .A2(n6028), .ZN(n8819) );
  AND4_X1 U5780 ( .A1(n5874), .A2(n5873), .A3(n5872), .A4(n5871), .ZN(n8063)
         );
  INV_X1 U5781 ( .A(n7991), .ZN(n8587) );
  NAND4_X1 U5782 ( .A1(n5779), .A2(n5778), .A3(n5777), .A4(n5776), .ZN(n8592)
         );
  OR2_X1 U5783 ( .A1(n5797), .A2(n5741), .ZN(n5744) );
  OR2_X1 U5784 ( .A1(n5757), .A2(n6256), .ZN(n5709) );
  OR2_X1 U5785 ( .A1(n7098), .A2(n6207), .ZN(n8727) );
  OR2_X1 U5786 ( .A1(n5774), .A2(n7360), .ZN(n5728) );
  INV_X1 U5787 ( .A(n4526), .ZN(n7025) );
  NAND2_X1 U5788 ( .A1(n4422), .A2(n6315), .ZN(n7055) );
  INV_X1 U5789 ( .A(n4534), .ZN(n9924) );
  OR2_X1 U5790 ( .A1(n7057), .A2(n6216), .ZN(n4534) );
  INV_X1 U5791 ( .A(n6220), .ZN(n4840) );
  NAND2_X1 U5792 ( .A1(n4811), .A2(n4809), .ZN(n7243) );
  NOR2_X1 U5793 ( .A1(n7651), .A2(n5836), .ZN(n7650) );
  OR2_X1 U5794 ( .A1(P2_U3150), .A2(n6298), .ZN(n8735) );
  NOR2_X1 U5795 ( .A1(n7658), .A2(n5841), .ZN(n7657) );
  AND2_X1 U5796 ( .A1(n4522), .A2(n6232), .ZN(n8617) );
  INV_X1 U5797 ( .A(n6234), .ZN(n4845) );
  NAND2_X1 U5798 ( .A1(n4847), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n4844) );
  NAND2_X1 U5799 ( .A1(n6234), .A2(n4847), .ZN(n4843) );
  INV_X1 U5800 ( .A(n8651), .ZN(n4847) );
  OR2_X1 U5801 ( .A1(n8672), .A2(n8914), .ZN(n4807) );
  INV_X1 U5802 ( .A(n6341), .ZN(n4806) );
  AOI21_X1 U5803 ( .B1(n4446), .B2(n8692), .A(n4525), .ZN(n8693) );
  INV_X1 U5804 ( .A(n6237), .ZN(n4830) );
  NAND2_X1 U5805 ( .A1(n4536), .A2(n4535), .ZN(n8724) );
  AOI21_X1 U5806 ( .B1(n4423), .B2(n8959), .A(n8722), .ZN(n4536) );
  INV_X1 U5807 ( .A(n8608), .ZN(n9929) );
  NOR2_X1 U5808 ( .A1(n6344), .A2(n8707), .ZN(n8721) );
  AND2_X1 U5809 ( .A1(n9914), .A2(n6107), .ZN(n8737) );
  OAI21_X1 U5810 ( .B1(n6191), .B2(n9949), .A(n6190), .ZN(n8756) );
  NOR2_X1 U5811 ( .A1(n6189), .A2(n6188), .ZN(n6190) );
  NOR2_X1 U5812 ( .A1(n8178), .A2(n9951), .ZN(n6188) );
  AND2_X1 U5813 ( .A1(n8810), .A2(n8917), .ZN(n4853) );
  NAND2_X1 U5814 ( .A1(n8860), .A2(n4799), .ZN(n8829) );
  NAND2_X1 U5815 ( .A1(n8852), .A2(n5990), .ZN(n8839) );
  NAND2_X1 U5816 ( .A1(n8860), .A2(n8358), .ZN(n8843) );
  NAND2_X1 U5817 ( .A1(n5980), .A2(n5979), .ZN(n8952) );
  NAND2_X1 U5818 ( .A1(n5967), .A2(n5966), .ZN(n8956) );
  NAND2_X1 U5819 ( .A1(n4775), .A2(n4421), .ZN(n7868) );
  AND2_X1 U5820 ( .A1(n4775), .A2(n8299), .ZN(n7898) );
  NAND2_X1 U5821 ( .A1(n7514), .A2(n8287), .ZN(n7560) );
  INV_X1 U5822 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n7380) );
  NAND2_X1 U5823 ( .A1(n6182), .A2(n7355), .ZN(n9939) );
  NAND2_X1 U5824 ( .A1(n7199), .A2(n7848), .ZN(n10005) );
  INV_X1 U5825 ( .A(n8846), .ZN(n8918) );
  INV_X1 U5826 ( .A(n8183), .ZN(n8759) );
  NAND2_X1 U5827 ( .A1(n6057), .A2(n6056), .ZN(n8979) );
  OR2_X1 U5828 ( .A1(n5764), .A2(n10143), .ZN(n6056) );
  NAND2_X1 U5829 ( .A1(n4660), .A2(n4666), .ZN(n8767) );
  AOI21_X1 U5830 ( .B1(n6171), .B2(n4781), .A(n4443), .ZN(n8765) );
  NAND2_X1 U5831 ( .A1(n6033), .A2(n6032), .ZN(n8991) );
  NAND2_X1 U5832 ( .A1(n6013), .A2(n6012), .ZN(n9002) );
  INV_X1 U5833 ( .A(n8521), .ZN(n9014) );
  NAND2_X1 U5834 ( .A1(n5952), .A2(n5951), .ZN(n9025) );
  NAND2_X1 U5835 ( .A1(n4787), .A2(n8340), .ZN(n8878) );
  NAND2_X1 U5836 ( .A1(n6166), .A2(n4788), .ZN(n4787) );
  NAND2_X1 U5837 ( .A1(n5940), .A2(n5939), .ZN(n9031) );
  NAND2_X1 U5838 ( .A1(n6166), .A2(n8338), .ZN(n8889) );
  NAND2_X1 U5839 ( .A1(n5928), .A2(n5927), .ZN(n9037) );
  NAND2_X1 U5840 ( .A1(n4651), .A2(n4652), .ZN(n8906) );
  NAND2_X1 U5841 ( .A1(n4766), .A2(n8328), .ZN(n8025) );
  NAND2_X1 U5842 ( .A1(n6165), .A2(n4763), .ZN(n4766) );
  NAND2_X1 U5843 ( .A1(n6165), .A2(n8323), .ZN(n8034) );
  AND3_X1 U5844 ( .A1(n5824), .A2(n5823), .A3(n5822), .ZN(n8304) );
  INV_X1 U5845 ( .A(n6958), .ZN(n8139) );
  INV_X1 U5846 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n9042) );
  INV_X1 U5847 ( .A(n5704), .ZN(n5703) );
  XNOR2_X1 U5848 ( .A(n5706), .B(n5705), .ZN(n8431) );
  INV_X1 U5849 ( .A(n6148), .ZN(n8136) );
  NAND2_X1 U5850 ( .A1(n6120), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6121) );
  INV_X1 U5851 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n10235) );
  INV_X1 U5852 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n7946) );
  INV_X1 U5853 ( .A(n8425), .ZN(n7848) );
  INV_X1 U5854 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n10344) );
  INV_X1 U5855 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7694) );
  INV_X1 U5856 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7546) );
  XNOR2_X1 U5857 ( .A(n5978), .B(n5977), .ZN(n7545) );
  INV_X1 U5858 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n10055) );
  INV_X1 U5859 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n10164) );
  INV_X1 U5860 ( .A(n8656), .ZN(n7016) );
  INV_X1 U5861 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n10300) );
  XNOR2_X1 U5862 ( .A(n5850), .B(n5860), .ZN(n6943) );
  INV_X1 U5863 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n10277) );
  INV_X1 U5864 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n10343) );
  NAND2_X1 U5865 ( .A1(n5748), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5765) );
  NAND2_X1 U5866 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n5746) );
  NAND2_X1 U5867 ( .A1(n5724), .A2(n5723), .ZN(n6977) );
  CLKBUF_X2 U5868 ( .A(P2_IR_REG_0__SCAN_IN), .Z(n9911) );
  INV_X1 U5869 ( .A(n9424), .ZN(n9658) );
  NAND2_X1 U5870 ( .A1(n4748), .A2(n4752), .ZN(n9064) );
  NAND2_X1 U5871 ( .A1(n6563), .A2(n4749), .ZN(n4748) );
  OAI21_X1 U5872 ( .B1(n7363), .B2(n4992), .A(n4411), .ZN(n4741) );
  NAND2_X1 U5873 ( .A1(n9127), .A2(n9129), .ZN(n4735) );
  NAND2_X1 U5874 ( .A1(n7970), .A2(n7971), .ZN(n7969) );
  NAND2_X1 U5875 ( .A1(n7885), .A2(n6501), .ZN(n7970) );
  NOR2_X1 U5876 ( .A1(n6563), .A2(n6562), .ZN(n9186) );
  AND4_X1 U5877 ( .A1(n5232), .A2(n5231), .A3(n5230), .A4(n5229), .ZN(n7841)
         );
  OR2_X1 U5878 ( .A1(n6611), .A2(n9591), .ZN(n9227) );
  AND2_X1 U5879 ( .A1(n9223), .A2(n9220), .ZN(n6583) );
  INV_X1 U5880 ( .A(n9229), .ZN(n9239) );
  AND2_X1 U5881 ( .A1(n6618), .A2(n9886), .ZN(n9247) );
  AND2_X1 U5882 ( .A1(n6617), .A2(n6602), .ZN(n9236) );
  INV_X1 U5883 ( .A(n9227), .ZN(n9244) );
  NAND2_X1 U5884 ( .A1(n6836), .A2(n4603), .ZN(n6841) );
  NAND2_X1 U5885 ( .A1(n6857), .A2(n6837), .ZN(n4603) );
  INV_X1 U5886 ( .A(n8114), .ZN(n9253) );
  XNOR2_X1 U5887 ( .A(n6905), .B(P1_REG2_REG_1__SCAN_IN), .ZN(n6875) );
  OAI21_X1 U5888 ( .B1(n7042), .B2(n4579), .A(n4578), .ZN(n9843) );
  NAND2_X1 U5889 ( .A1(n9840), .A2(n4581), .ZN(n4578) );
  NAND2_X1 U5890 ( .A1(n9840), .A2(n4580), .ZN(n4579) );
  INV_X1 U5891 ( .A(n7041), .ZN(n4580) );
  NAND2_X1 U5892 ( .A1(n9314), .A2(n9313), .ZN(n9312) );
  AND2_X1 U5893 ( .A1(n9312), .A2(n4592), .ZN(n9828) );
  NAND2_X1 U5894 ( .A1(n7002), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n4592) );
  NOR2_X1 U5895 ( .A1(n7473), .A2(n4595), .ZN(n7477) );
  AND2_X1 U5896 ( .A1(n7474), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n4595) );
  NOR2_X1 U5897 ( .A1(n7477), .A2(n7476), .ZN(n9323) );
  NOR2_X1 U5898 ( .A1(n9364), .A2(n4597), .ZN(n9861) );
  AND2_X1 U5899 ( .A1(n9365), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n4597) );
  INV_X1 U5900 ( .A(n4577), .ZN(n9378) );
  XNOR2_X1 U5901 ( .A(n4576), .B(P1_REG2_REG_19__SCAN_IN), .ZN(n9384) );
  NAND2_X1 U5902 ( .A1(n4577), .A2(n9377), .ZN(n4576) );
  INV_X1 U5903 ( .A(n9384), .ZN(n9387) );
  AND2_X1 U5904 ( .A1(n6965), .A2(n8195), .ZN(n9386) );
  INV_X1 U5905 ( .A(n9648), .ZN(n9441) );
  NAND2_X1 U5906 ( .A1(n4899), .A2(n4900), .ZN(n9412) );
  NAND2_X1 U5907 ( .A1(n4899), .A2(n4461), .ZN(n9645) );
  INV_X1 U5908 ( .A(n9465), .ZN(n9669) );
  NAND2_X1 U5909 ( .A1(n9515), .A2(n6659), .ZN(n9495) );
  INV_X1 U5910 ( .A(n9545), .ZN(n9688) );
  INV_X1 U5911 ( .A(n9695), .ZN(n9524) );
  NAND2_X1 U5912 ( .A1(n4703), .A2(n4705), .ZN(n8052) );
  AND2_X1 U5913 ( .A1(n4912), .A2(n4913), .ZN(n8049) );
  NAND2_X1 U5914 ( .A1(n8099), .A2(n5347), .ZN(n4912) );
  NAND2_X1 U5915 ( .A1(n5337), .A2(n5336), .ZN(n9059) );
  OAI21_X1 U5916 ( .B1(n7412), .B2(n4893), .A(n4891), .ZN(n7592) );
  NAND2_X1 U5917 ( .A1(n7443), .A2(n7442), .ZN(n7441) );
  NAND2_X1 U5918 ( .A1(n7412), .A2(n5233), .ZN(n7443) );
  INV_X1 U5919 ( .A(n9620), .ZN(n9585) );
  OR2_X1 U5920 ( .A1(n5673), .A2(n5666), .ZN(n9489) );
  NAND2_X1 U5921 ( .A1(n7732), .A2(n7849), .ZN(n9877) );
  NAND2_X1 U5922 ( .A1(n4418), .A2(n6843), .ZN(n9876) );
  OR2_X1 U5923 ( .A1(n5155), .A2(n6921), .ZN(n5165) );
  INV_X1 U5924 ( .A(n9644), .ZN(n9734) );
  AND2_X2 U5925 ( .A1(n5683), .A2(n6600), .ZN(n9910) );
  NAND2_X1 U5926 ( .A1(n4903), .A2(n5526), .ZN(n9422) );
  OR3_X1 U5927 ( .A1(n9709), .A2(n9708), .A3(n9707), .ZN(n9784) );
  AND2_X1 U5928 ( .A1(n4916), .A2(n4433), .ZN(n9541) );
  NAND2_X1 U5929 ( .A1(n5396), .A2(n5395), .ZN(n9792) );
  NAND2_X1 U5930 ( .A1(n5366), .A2(n5365), .ZN(n9801) );
  OAI21_X1 U5931 ( .B1(n8099), .B2(n4910), .A(n4908), .ZN(n9619) );
  NAND2_X1 U5932 ( .A1(n5285), .A2(n5284), .ZN(n9210) );
  INV_X1 U5933 ( .A(n9786), .ZN(n9803) );
  NAND2_X1 U5934 ( .A1(n7487), .A2(n5002), .ZN(n7335) );
  XNOR2_X1 U5935 ( .A(n6634), .B(n6633), .ZN(n9812) );
  OAI22_X1 U5936 ( .A1(n6630), .A2(n6629), .B1(SI_30_), .B2(n6628), .ZN(n6634)
         );
  INV_X1 U5937 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n5017) );
  NAND2_X1 U5938 ( .A1(n9813), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5018) );
  NAND2_X1 U5939 ( .A1(n4617), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5020) );
  CLKBUF_X1 U5940 ( .A(n5650), .Z(n8195) );
  INV_X1 U5941 ( .A(n5608), .ZN(n8082) );
  INV_X1 U5942 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n10271) );
  INV_X1 U5943 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7851) );
  INV_X1 U5944 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7734) );
  INV_X1 U5945 ( .A(n4418), .ZN(n7732) );
  INV_X1 U5946 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7548) );
  CLKBUF_X1 U5947 ( .A(n5617), .Z(n4519) );
  NOR2_X1 U5948 ( .A1(n6915), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9817) );
  INV_X1 U5949 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n7169) );
  INV_X1 U5950 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n10285) );
  INV_X1 U5951 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n6941) );
  NAND2_X1 U5952 ( .A1(n4700), .A2(n4856), .ZN(n5189) );
  INV_X1 U5953 ( .A(n4698), .ZN(n4856) );
  NAND2_X1 U5954 ( .A1(n4855), .A2(n5164), .ZN(n4700) );
  NAND2_X1 U5955 ( .A1(n4858), .A2(n5046), .ZN(n5177) );
  INV_X1 U5956 ( .A(n6905), .ZN(n6916) );
  NAND2_X1 U5957 ( .A1(n4948), .A2(n8545), .ZN(n4946) );
  NAND2_X1 U5958 ( .A1(n4521), .A2(n6232), .ZN(n7925) );
  INV_X1 U5959 ( .A(n4846), .ZN(n8633) );
  INV_X1 U5960 ( .A(n4831), .ZN(n8666) );
  INV_X1 U5961 ( .A(n4826), .ZN(n8699) );
  OAI21_X1 U5962 ( .B1(n6363), .B2(n8922), .A(n6362), .ZN(n6364) );
  INV_X1 U5963 ( .A(n6400), .ZN(n6401) );
  OAI22_X1 U5964 ( .A1(n6399), .A2(n8950), .B1(n10029), .B2(n10302), .ZN(n6400) );
  NOR2_X1 U5965 ( .A1(n5000), .A2(n6183), .ZN(n6184) );
  NOR2_X1 U5966 ( .A1(n8401), .A2(n8950), .ZN(n6183) );
  AOI21_X1 U5967 ( .B1(n8997), .B2(n8967), .A(n4501), .ZN(n8938) );
  NAND2_X1 U5968 ( .A1(n6395), .A2(n6396), .ZN(n6398) );
  AND2_X1 U5969 ( .A1(n6370), .A2(n4499), .ZN(n6371) );
  AOI21_X1 U5970 ( .B1(n8997), .B2(n9038), .A(n4500), .ZN(n8998) );
  INV_X1 U5971 ( .A(n4588), .ZN(n7067) );
  INV_X1 U5972 ( .A(n4586), .ZN(n7070) );
  AND2_X1 U5973 ( .A1(n5680), .A2(n5679), .ZN(n5681) );
  OAI211_X1 U5974 ( .C1(n6873), .C2(n7048), .A(n5166), .B(n5165), .ZN(n7191)
         );
  AND2_X1 U5975 ( .A1(n4964), .A2(n8504), .ZN(n4419) );
  OR2_X1 U5976 ( .A1(n9139), .A2(n6533), .ZN(n4420) );
  AND2_X1 U5977 ( .A1(n8299), .A2(n8315), .ZN(n4421) );
  NAND2_X2 U5978 ( .A1(n5022), .A2(n9820), .ZN(n5369) );
  OR2_X1 U5979 ( .A1(n6314), .A2(n6313), .ZN(n4422) );
  OR2_X1 U5980 ( .A1(n8708), .A2(n6238), .ZN(n4423) );
  XNOR2_X1 U5981 ( .A(n6096), .B(P2_IR_REG_20__SCAN_IN), .ZN(n7197) );
  OR2_X1 U5982 ( .A1(n4878), .A2(n5280), .ZN(n4424) );
  AND2_X1 U5983 ( .A1(n6824), .A2(n4453), .ZN(n4425) );
  AND2_X1 U5984 ( .A1(n4973), .A2(n4972), .ZN(n4426) );
  INV_X1 U5985 ( .A(n8176), .ZN(n8793) );
  OR2_X1 U5986 ( .A1(n8505), .A2(n8573), .ZN(n4427) );
  AND2_X1 U5987 ( .A1(n6556), .A2(n4733), .ZN(n4428) );
  AND2_X1 U5988 ( .A1(n4926), .A2(n8488), .ZN(n4429) );
  AND2_X1 U5989 ( .A1(n4504), .A2(n4749), .ZN(n4430) );
  NAND2_X1 U5990 ( .A1(n5303), .A2(n5302), .ZN(n7889) );
  AND2_X1 U5991 ( .A1(n4854), .A2(n8819), .ZN(n4431) );
  AND2_X1 U5992 ( .A1(n9756), .A2(n6825), .ZN(n4432) );
  OR2_X1 U5993 ( .A1(n9714), .A2(n9554), .ZN(n4433) );
  INV_X1 U5994 ( .A(n8392), .ZN(n4567) );
  AND3_X1 U5995 ( .A1(n4543), .A2(n8357), .A3(n4551), .ZN(n4434) );
  AND2_X1 U5996 ( .A1(n8167), .A2(n8841), .ZN(n4435) );
  AND2_X1 U5997 ( .A1(n8358), .A2(n8359), .ZN(n8857) );
  OAI21_X1 U5998 ( .B1(n6785), .B2(n6784), .A(n4475), .ZN(n4604) );
  AND2_X1 U5999 ( .A1(n8176), .A2(n4671), .ZN(n4436) );
  AND2_X1 U6000 ( .A1(n4735), .A2(n4734), .ZN(n4437) );
  AND2_X1 U6001 ( .A1(n4939), .A2(n4458), .ZN(n4438) );
  AND4_X1 U6002 ( .A1(n5523), .A2(n5522), .A3(n5521), .A4(n5520), .ZN(n9657)
         );
  AND2_X1 U6003 ( .A1(n4837), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n4439) );
  INV_X1 U6004 ( .A(n4741), .ZN(n7523) );
  XOR2_X1 U6005 ( .A(n8235), .B(n8186), .Z(n4440) );
  NAND2_X1 U6006 ( .A1(n6408), .A2(n6407), .ZN(n6424) );
  NOR2_X1 U6007 ( .A1(n7563), .A2(n7562), .ZN(n4441) );
  XNOR2_X1 U6008 ( .A(n6119), .B(n6118), .ZN(n6129) );
  AND2_X1 U6009 ( .A1(n8495), .A2(n8496), .ZN(n4442) );
  NAND2_X1 U6010 ( .A1(n4730), .A2(n4733), .ZN(n9070) );
  OAI21_X1 U6011 ( .B1(n7204), .B2(n7203), .A(n7202), .ZN(n7209) );
  NAND2_X1 U6012 ( .A1(n4935), .A2(n5692), .ZN(n5766) );
  XNOR2_X1 U6013 ( .A(n5018), .B(n5017), .ZN(n5021) );
  NOR2_X1 U6014 ( .A1(n6179), .A2(n6178), .ZN(n4443) );
  AND2_X1 U6015 ( .A1(n9423), .A2(n9658), .ZN(n4444) );
  AND2_X1 U6016 ( .A1(n4420), .A2(n9129), .ZN(n4445) );
  INV_X1 U6017 ( .A(n4981), .ZN(n4969) );
  AND2_X1 U6018 ( .A1(n4831), .A2(n4830), .ZN(n4446) );
  INV_X1 U6019 ( .A(n8401), .ZN(n8192) );
  AND2_X1 U6020 ( .A1(n6082), .A2(n6081), .ZN(n8401) );
  OR2_X1 U6021 ( .A1(n5820), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n4447) );
  INV_X1 U6022 ( .A(n6770), .ZN(n4714) );
  NAND2_X1 U6023 ( .A1(n4924), .A2(n4923), .ZN(n8556) );
  NAND2_X1 U6024 ( .A1(n4925), .A2(n8175), .ZN(n8487) );
  NAND2_X1 U6025 ( .A1(n4523), .A2(n6948), .ZN(n6232) );
  OR2_X1 U6026 ( .A1(n7991), .A2(n7950), .ZN(n8299) );
  NAND4_X1 U6027 ( .A1(n5745), .A2(n5744), .A3(n5743), .A4(n5742), .ZN(n5755)
         );
  AND2_X1 U6028 ( .A1(n8588), .A2(n7785), .ZN(n4448) );
  AND2_X1 U6029 ( .A1(n9139), .A2(n6533), .ZN(n4449) );
  AND2_X1 U6030 ( .A1(n6563), .A2(n6562), .ZN(n4450) );
  NAND2_X1 U6031 ( .A1(n5424), .A2(n5423), .ZN(n9696) );
  AND2_X1 U6032 ( .A1(n8325), .A2(n8326), .ZN(n4451) );
  OR2_X1 U6033 ( .A1(n9037), .A2(n8894), .ZN(n4452) );
  INV_X1 U6034 ( .A(n9252), .ZN(n9240) );
  INV_X1 U6035 ( .A(n6044), .ZN(n4672) );
  AND2_X1 U6036 ( .A1(n6820), .A2(n6837), .ZN(n4453) );
  INV_X1 U6037 ( .A(n5067), .ZN(n4881) );
  NAND2_X1 U6038 ( .A1(n5460), .A2(n5459), .ZN(n9685) );
  OR2_X1 U6039 ( .A1(n9002), .A2(n8827), .ZN(n8242) );
  NAND2_X1 U6040 ( .A1(n6022), .A2(n6021), .ZN(n4854) );
  INV_X1 U6041 ( .A(n4911), .ZN(n4910) );
  NOR2_X1 U6042 ( .A1(n4454), .A2(n5346), .ZN(n4911) );
  INV_X1 U6043 ( .A(n4669), .ZN(n4667) );
  AOI21_X1 U6044 ( .B1(n4670), .B2(n4672), .A(n8774), .ZN(n4669) );
  NOR2_X1 U6045 ( .A1(n9739), .A2(n9624), .ZN(n4454) );
  NAND2_X1 U6046 ( .A1(n7237), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n4455) );
  OAI21_X1 U6047 ( .B1(n4445), .B2(n4732), .A(n6546), .ZN(n4731) );
  NAND2_X1 U6048 ( .A1(n5381), .A2(n5380), .ZN(n9724) );
  AND2_X1 U6049 ( .A1(n5263), .A2(n4881), .ZN(n4456) );
  INV_X1 U6050 ( .A(n6821), .ZN(n5687) );
  INV_X1 U6051 ( .A(n9059), .ZN(n8115) );
  NAND2_X1 U6052 ( .A1(n5115), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5586) );
  AND2_X1 U6053 ( .A1(n6819), .A2(n9405), .ZN(n4457) );
  NAND2_X1 U6054 ( .A1(n7788), .A2(n7804), .ZN(n4458) );
  NAND2_X1 U6055 ( .A1(n7021), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n4459) );
  AND2_X1 U6056 ( .A1(n6000), .A2(n5990), .ZN(n4460) );
  AND2_X1 U6057 ( .A1(n4900), .A2(n6703), .ZN(n4461) );
  INV_X1 U6058 ( .A(n4713), .ZN(n4712) );
  NOR2_X1 U6059 ( .A1(n6774), .A2(n4714), .ZN(n4713) );
  AND2_X1 U6060 ( .A1(n4807), .A2(n4806), .ZN(n4462) );
  AND2_X1 U6061 ( .A1(n4710), .A2(n4715), .ZN(n4463) );
  NAND2_X1 U6062 ( .A1(n4826), .A2(n4423), .ZN(n4464) );
  NAND2_X1 U6063 ( .A1(n4616), .A2(n4920), .ZN(n4617) );
  INV_X1 U6064 ( .A(n4733), .ZN(n4732) );
  NAND2_X1 U6065 ( .A1(n4482), .A2(n4420), .ZN(n4733) );
  INV_X1 U6066 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n9815) );
  NOR2_X1 U6067 ( .A1(n9258), .A2(n7839), .ZN(n4465) );
  NOR2_X1 U6068 ( .A1(n9248), .A2(n9134), .ZN(n4466) );
  NAND2_X1 U6069 ( .A1(n5048), .A2(SI_4_), .ZN(n4467) );
  INV_X1 U6070 ( .A(n4650), .ZN(n4649) );
  NAND2_X1 U6071 ( .A1(n4652), .A2(n4452), .ZN(n4650) );
  OR2_X1 U6072 ( .A1(n5308), .A2(n5136), .ZN(n4468) );
  INV_X1 U6073 ( .A(n4764), .ZN(n4763) );
  NAND2_X1 U6074 ( .A1(n8323), .A2(n4765), .ZN(n4764) );
  AND2_X1 U6075 ( .A1(n4974), .A2(n4968), .ZN(n4469) );
  AND2_X1 U6076 ( .A1(n9714), .A2(n9554), .ZN(n4470) );
  INV_X1 U6077 ( .A(n9756), .ZN(n9401) );
  AND2_X1 U6078 ( .A1(n6627), .A2(n6626), .ZN(n9756) );
  NOR2_X1 U6079 ( .A1(n6737), .A2(n7413), .ZN(n4471) );
  NOR2_X1 U6080 ( .A1(n6507), .A2(n6506), .ZN(n4472) );
  INV_X1 U6081 ( .A(n5234), .ZN(n4563) );
  NOR2_X2 U6082 ( .A1(n5820), .A2(n4958), .ZN(n6115) );
  OR2_X1 U6083 ( .A1(n8817), .A2(n8368), .ZN(n4473) );
  XNOR2_X1 U6084 ( .A(n5405), .B(n5579), .ZN(n5617) );
  NAND2_X1 U6085 ( .A1(n8397), .A2(n8204), .ZN(n8394) );
  INV_X1 U6086 ( .A(n8394), .ZN(n4568) );
  AND2_X1 U6087 ( .A1(n4629), .A2(n4630), .ZN(n4474) );
  AND2_X1 U6088 ( .A1(n6783), .A2(n4605), .ZN(n4475) );
  AND2_X1 U6089 ( .A1(n5050), .A2(SI_5_), .ZN(n4476) );
  AND2_X1 U6090 ( .A1(n5079), .A2(SI_12_), .ZN(n4477) );
  INV_X1 U6091 ( .A(n4656), .ZN(n4655) );
  OR2_X1 U6092 ( .A1(n5924), .A2(n4657), .ZN(n4656) );
  AND2_X1 U6093 ( .A1(n5010), .A2(n5393), .ZN(n4478) );
  AND2_X1 U6094 ( .A1(n5093), .A2(SI_16_), .ZN(n4479) );
  OR2_X1 U6095 ( .A1(n7360), .A2(n9911), .ZN(n4480) );
  OR2_X1 U6096 ( .A1(n5948), .A2(n8888), .ZN(n4481) );
  OR2_X1 U6097 ( .A1(n9128), .A2(n4449), .ZN(n4482) );
  INV_X1 U6098 ( .A(n4624), .ZN(n4623) );
  NAND2_X1 U6099 ( .A1(n6824), .A2(n6818), .ZN(n4624) );
  AND2_X1 U6100 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n4483) );
  OR2_X1 U6101 ( .A1(n8521), .A2(n8856), .ZN(n8365) );
  INV_X1 U6102 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n5377) );
  INV_X1 U6103 ( .A(n4626), .ZN(n4625) );
  NAND2_X1 U6104 ( .A1(n6822), .A2(n6823), .ZN(n4626) );
  NOR2_X1 U6105 ( .A1(n6031), .A2(n4431), .ZN(n4484) );
  NAND2_X1 U6106 ( .A1(n5408), .A2(n5407), .ZN(n9714) );
  OR2_X1 U6107 ( .A1(n8340), .A2(n8406), .ZN(n4485) );
  OR3_X1 U6108 ( .A1(n5378), .A2(n4757), .A3(n5580), .ZN(n4486) );
  AND2_X1 U6109 ( .A1(n8991), .A2(n8806), .ZN(n4487) );
  NAND2_X1 U6110 ( .A1(n5478), .A2(n5477), .ZN(n9676) );
  INV_X1 U6111 ( .A(n9676), .ZN(n4683) );
  AND2_X1 U6112 ( .A1(n4668), .A2(n4672), .ZN(n4488) );
  AND2_X1 U6113 ( .A1(n4884), .A2(n4882), .ZN(n4489) );
  OR2_X1 U6114 ( .A1(n4440), .A2(n4949), .ZN(n4490) );
  AND2_X1 U6115 ( .A1(n6148), .A2(n4922), .ZN(n4491) );
  OR2_X1 U6116 ( .A1(n5737), .A2(n6977), .ZN(n4492) );
  AND2_X1 U6117 ( .A1(n9756), .A2(n4677), .ZN(n4493) );
  AOI21_X1 U6118 ( .B1(n8347), .B2(n8402), .A(n4552), .ZN(n4551) );
  OR2_X1 U6119 ( .A1(n8478), .A2(n8841), .ZN(n8366) );
  NAND2_X1 U6120 ( .A1(n4941), .A2(n7789), .ZN(n4494) );
  INV_X1 U6121 ( .A(n4800), .ZN(n4799) );
  NAND2_X1 U6122 ( .A1(n8365), .A2(n8358), .ZN(n4800) );
  INV_X1 U6123 ( .A(n5617), .ZN(n5666) );
  INV_X2 U6124 ( .A(n6420), .ZN(n6448) );
  INV_X1 U6125 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n4695) );
  AND2_X1 U6126 ( .A1(n4965), .A2(n4442), .ZN(n4495) );
  AND2_X1 U6127 ( .A1(n4961), .A2(n4419), .ZN(n4496) );
  AND2_X1 U6128 ( .A1(n8106), .A2(n4690), .ZN(n4497) );
  NAND2_X1 U6129 ( .A1(n8166), .A2(n8523), .ZN(n8479) );
  INV_X1 U6130 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5010) );
  AND2_X1 U6131 ( .A1(n5330), .A2(n5008), .ZN(n5333) );
  XNOR2_X1 U6132 ( .A(n4725), .B(P1_IR_REG_25__SCAN_IN), .ZN(n5608) );
  NAND2_X1 U6133 ( .A1(n5401), .A2(n4984), .ZN(n9563) );
  INV_X1 U6134 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n4957) );
  NAND2_X1 U6135 ( .A1(n6377), .A2(n6376), .ZN(n6395) );
  INV_X1 U6136 ( .A(n8480), .ZN(n4933) );
  NAND2_X1 U6137 ( .A1(n4726), .A2(n4724), .ZN(n5607) );
  AND3_X1 U6138 ( .A1(n9092), .A2(n9236), .A3(n9091), .ZN(n4498) );
  NAND2_X1 U6139 ( .A1(n6046), .A2(n6045), .ZN(n8985) );
  INV_X1 U6140 ( .A(n8985), .ZN(n4671) );
  OR2_X1 U6141 ( .A1(n8401), .A2(n9013), .ZN(n4499) );
  AND2_X1 U6142 ( .A1(n4854), .A2(n6396), .ZN(n4500) );
  AND2_X1 U6143 ( .A1(n4854), .A2(n8966), .ZN(n4501) );
  OR2_X1 U6144 ( .A1(n8572), .A2(n8573), .ZN(n4965) );
  AND2_X1 U6145 ( .A1(n8177), .A2(n8176), .ZN(n4502) );
  NAND2_X1 U6146 ( .A1(n5554), .A2(n5553), .ZN(n9649) );
  INV_X1 U6147 ( .A(n9649), .ZN(n4679) );
  NOR2_X1 U6148 ( .A1(n8638), .A2(n6338), .ZN(n4503) );
  OR2_X1 U6149 ( .A1(n6566), .A2(n6565), .ZN(n4504) );
  INV_X1 U6150 ( .A(n8841), .ZN(n8818) );
  AND3_X1 U6151 ( .A1(n6009), .A2(n6008), .A3(n6007), .ZN(n8841) );
  INV_X1 U6152 ( .A(n7933), .ZN(n6948) );
  AND2_X1 U6153 ( .A1(n5864), .A2(n5895), .ZN(n7933) );
  NAND2_X1 U6154 ( .A1(n9550), .A2(n4686), .ZN(n4687) );
  NAND2_X1 U6155 ( .A1(n7237), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n4505) );
  AND2_X1 U6156 ( .A1(n4846), .A2(n4845), .ZN(n4506) );
  OR2_X1 U6157 ( .A1(n5378), .A2(P1_IR_REG_16__SCAN_IN), .ZN(n4507) );
  INV_X1 U6158 ( .A(n9764), .ZN(n9452) );
  NAND2_X1 U6159 ( .A1(n5515), .A2(n5514), .ZN(n9764) );
  AOI21_X1 U6160 ( .B1(n8479), .B2(n8480), .A(n4934), .ZN(n4931) );
  AND2_X1 U6161 ( .A1(n5436), .A2(SI_21_), .ZN(n4508) );
  NAND2_X1 U6162 ( .A1(n5112), .A2(SI_20_), .ZN(n4509) );
  NAND2_X1 U6163 ( .A1(n6943), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n4510) );
  XNOR2_X1 U6164 ( .A(n6095), .B(P2_IR_REG_21__SCAN_IN), .ZN(n7196) );
  INV_X2 U6165 ( .A(n10017), .ZN(n10016) );
  OR2_X1 U6166 ( .A1(n6843), .A2(n4519), .ZN(n6825) );
  INV_X1 U6167 ( .A(n6825), .ZN(n6837) );
  XNOR2_X1 U6168 ( .A(n6121), .B(n10121), .ZN(n6133) );
  AND2_X1 U6169 ( .A1(n4970), .A2(n4969), .ZN(n4511) );
  INV_X1 U6170 ( .A(n8543), .ZN(n4963) );
  NOR2_X1 U6171 ( .A1(n7657), .A2(n6230), .ZN(n4512) );
  INV_X1 U6172 ( .A(n9128), .ZN(n4734) );
  AND2_X1 U6173 ( .A1(n4740), .A2(n4739), .ZN(n4513) );
  INV_X1 U6174 ( .A(n4681), .ZN(n7444) );
  NOR2_X1 U6175 ( .A1(n7331), .A2(n7457), .ZN(n4681) );
  NOR2_X1 U6176 ( .A1(n7650), .A2(n6329), .ZN(n4514) );
  INV_X1 U6177 ( .A(SI_20_), .ZN(n5420) );
  INV_X1 U6178 ( .A(n5346), .ZN(n4913) );
  INV_X1 U6179 ( .A(n8591), .ZN(n4972) );
  NAND2_X1 U6180 ( .A1(n5120), .A2(n4617), .ZN(n5643) );
  AND3_X2 U6181 ( .A1(n6153), .A2(n6355), .A3(n7104), .ZN(n10029) );
  INV_X1 U6182 ( .A(n7839), .ZN(n4680) );
  NAND2_X1 U6183 ( .A1(n7531), .A2(n5738), .ZN(n7534) );
  OR2_X1 U6184 ( .A1(n7312), .A2(n5811), .ZN(n7311) );
  INV_X1 U6185 ( .A(n8722), .ZN(n4537) );
  INV_X1 U6186 ( .A(n8688), .ZN(n7164) );
  NAND2_X1 U6187 ( .A1(n7088), .A2(n6411), .ZN(n7187) );
  INV_X1 U6188 ( .A(n7187), .ZN(n4675) );
  AND2_X1 U6189 ( .A1(n4814), .A2(n4813), .ZN(n4515) );
  AND2_X1 U6190 ( .A1(n4841), .A2(n4840), .ZN(n4516) );
  AND2_X1 U6191 ( .A1(n4422), .A2(n4815), .ZN(n4517) );
  OR2_X1 U6192 ( .A1(n5623), .A2(n7148), .ZN(n7146) );
  AND2_X1 U6193 ( .A1(n4534), .A2(n4533), .ZN(n4518) );
  INV_X1 U6194 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n5304) );
  AND4_X1 U6195 ( .A1(n4468), .A2(n5140), .A3(n5139), .A4(n5138), .ZN(n6419)
         );
  INV_X1 U6196 ( .A(n9839), .ZN(n4581) );
  INV_X1 U6197 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n4596) );
  XNOR2_X1 U6198 ( .A(n6337), .B(n8643), .ZN(n8639) );
  XNOR2_X1 U6199 ( .A(n6233), .B(n8643), .ZN(n8634) );
  NAND2_X1 U6200 ( .A1(n9120), .A2(n9121), .ZN(n9221) );
  INV_X1 U6201 ( .A(n9093), .ZN(n4738) );
  INV_X1 U6202 ( .A(n6513), .ZN(n6511) );
  OAI21_X2 U6203 ( .B1(n6560), .B2(n6559), .A(n9111), .ZN(n6563) );
  AOI21_X1 U6204 ( .B1(n7173), .B2(n7174), .A(n4996), .ZN(n7253) );
  OAI21_X2 U6205 ( .B1(n5378), .B2(n4757), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n5591) );
  NAND2_X1 U6206 ( .A1(n4570), .A2(n8387), .ZN(n4569) );
  OAI211_X1 U6207 ( .C1(n8378), .C2(n8402), .A(n4860), .B(n8774), .ZN(n4859)
         );
  NAND2_X1 U6208 ( .A1(n4859), .A2(n8381), .ZN(n8382) );
  INV_X1 U6209 ( .A(n4523), .ZN(n4520) );
  NAND3_X1 U6210 ( .A1(n4521), .A2(P2_REG1_REG_11__SCAN_IN), .A3(n6232), .ZN(
        n4522) );
  INV_X1 U6211 ( .A(n4522), .ZN(n7924) );
  NOR2_X1 U6212 ( .A1(n6973), .A2(n6213), .ZN(n7027) );
  INV_X1 U6213 ( .A(n7057), .ZN(n4532) );
  NAND2_X1 U6214 ( .A1(n8700), .A2(n4423), .ZN(n4535) );
  OR2_X1 U6215 ( .A1(n8700), .A2(n8959), .ZN(n4826) );
  INV_X1 U6216 ( .A(n8724), .ZN(n8723) );
  NAND2_X1 U6217 ( .A1(n8346), .A2(n8406), .ZN(n4543) );
  NAND2_X1 U6218 ( .A1(n4544), .A2(n4545), .ZN(n8370) );
  AND2_X1 U6219 ( .A1(n4549), .A2(n8366), .ZN(n4548) );
  NAND2_X1 U6220 ( .A1(n5235), .A2(n5062), .ZN(n4562) );
  INV_X1 U6221 ( .A(n4562), .ZN(n4554) );
  AOI21_X1 U6222 ( .B1(n4554), .B2(n4558), .A(n4456), .ZN(n4553) );
  NAND3_X1 U6223 ( .A1(n4562), .A2(n4559), .A3(n5263), .ZN(n4557) );
  NAND3_X1 U6224 ( .A1(n8312), .A2(n4572), .A3(n4571), .ZN(n8316) );
  NAND3_X1 U6225 ( .A1(n8339), .A2(n8340), .A3(n8406), .ZN(n4575) );
  NAND3_X1 U6226 ( .A1(n6744), .A2(n6743), .A3(n6756), .ZN(n4602) );
  NAND2_X1 U6227 ( .A1(n5330), .A2(n4920), .ZN(n5115) );
  AND2_X2 U6228 ( .A1(n5297), .A2(n5007), .ZN(n5330) );
  INV_X1 U6229 ( .A(n4617), .ZN(n5119) );
  AOI21_X1 U6230 ( .B1(n6817), .B2(n4623), .A(n4620), .ZN(n6828) );
  NAND2_X1 U6231 ( .A1(n4629), .A2(n4628), .ZN(n4639) );
  NAND2_X1 U6232 ( .A1(n5739), .A2(n9961), .ZN(n8256) );
  OR2_X1 U6233 ( .A1(n9961), .A2(n5739), .ZN(n8254) );
  NAND2_X1 U6234 ( .A1(n8432), .A2(n8431), .ZN(n5797) );
  NAND3_X1 U6235 ( .A1(n8432), .A2(n8431), .A3(P2_REG0_REG_1__SCAN_IN), .ZN(
        n5710) );
  XNOR2_X2 U6236 ( .A(n5702), .B(n9042), .ZN(n8432) );
  OAI21_X1 U6237 ( .B1(n7550), .B2(n4644), .A(n4642), .ZN(n7685) );
  NAND2_X1 U6238 ( .A1(n4641), .A2(n4640), .ZN(n7801) );
  NAND2_X1 U6239 ( .A1(n7550), .A2(n4642), .ZN(n4641) );
  OR2_X1 U6240 ( .A1(n8145), .A2(n8908), .ZN(n4658) );
  INV_X1 U6241 ( .A(n8851), .ZN(n4659) );
  OR2_X1 U6242 ( .A1(n6031), .A2(n4667), .ZN(n4660) );
  OR2_X1 U6243 ( .A1(n6031), .A2(n4670), .ZN(n4668) );
  NAND3_X1 U6244 ( .A1(n6031), .A2(n4666), .A3(n4665), .ZN(n4664) );
  AND2_X1 U6245 ( .A1(n9423), .A2(n4676), .ZN(n9416) );
  NAND2_X1 U6246 ( .A1(n9423), .A2(n4677), .ZN(n9400) );
  INV_X1 U6247 ( .A(n4687), .ZN(n9500) );
  INV_X1 U6248 ( .A(n5122), .ZN(n4696) );
  NAND2_X1 U6249 ( .A1(n5127), .A2(n5126), .ZN(n5038) );
  NAND2_X1 U6250 ( .A1(n4699), .A2(n4697), .ZN(n5207) );
  NAND3_X1 U6251 ( .A1(n4855), .A2(n5190), .A3(n5164), .ZN(n4699) );
  INV_X1 U6252 ( .A(n9622), .ZN(n4709) );
  OR2_X1 U6253 ( .A1(n5584), .A2(n5583), .ZN(n4724) );
  AOI21_X2 U6254 ( .B1(n4728), .B2(n4428), .A(n4727), .ZN(n9112) );
  AND2_X2 U6255 ( .A1(n9222), .A2(n6597), .ZN(n9093) );
  NAND2_X1 U6256 ( .A1(n6563), .A2(n4430), .ZN(n4745) );
  NAND2_X1 U6257 ( .A1(n4745), .A2(n4746), .ZN(n9153) );
  NAND2_X1 U6258 ( .A1(n9051), .A2(n6517), .ZN(n6520) );
  NAND2_X1 U6259 ( .A1(n6516), .A2(n6515), .ZN(n9051) );
  NAND2_X1 U6260 ( .A1(n6430), .A2(n6429), .ZN(n6431) );
  NAND2_X1 U6261 ( .A1(n6413), .A2(n6412), .ZN(n6437) );
  NAND3_X1 U6262 ( .A1(n4768), .A2(n8246), .A3(n4767), .ZN(n7554) );
  NAND3_X1 U6263 ( .A1(n6161), .A2(n4769), .A3(n8282), .ZN(n4767) );
  NAND3_X1 U6264 ( .A1(n7428), .A2(n4769), .A3(n6161), .ZN(n4768) );
  NAND2_X1 U6265 ( .A1(n7805), .A2(n4421), .ZN(n4771) );
  NAND2_X1 U6266 ( .A1(n4771), .A2(n4772), .ZN(n6164) );
  NAND2_X1 U6267 ( .A1(n4777), .A2(n4778), .ZN(n6180) );
  NAND2_X1 U6268 ( .A1(n6166), .A2(n4783), .ZN(n4782) );
  NAND2_X1 U6269 ( .A1(n4782), .A2(n4784), .ZN(n8869) );
  NAND2_X1 U6270 ( .A1(n6382), .A2(n4791), .ZN(n4790) );
  NAND2_X1 U6271 ( .A1(n6382), .A2(n6381), .ZN(n8203) );
  NAND2_X1 U6272 ( .A1(n4790), .A2(n4793), .ZN(n8239) );
  OAI21_X1 U6273 ( .B1(n8858), .B2(n4800), .A(n4797), .ZN(n6170) );
  INV_X1 U6274 ( .A(n5724), .ZN(n4801) );
  OAI21_X1 U6275 ( .B1(n4802), .B2(n4801), .A(n6310), .ZN(n6972) );
  XNOR2_X1 U6276 ( .A(n6340), .B(n8674), .ZN(n8672) );
  INV_X1 U6277 ( .A(n4814), .ZN(n7129) );
  INV_X1 U6278 ( .A(n6321), .ZN(n4813) );
  OAI21_X1 U6279 ( .B1(n7651), .B2(n4818), .A(n4817), .ZN(n7769) );
  XNOR2_X1 U6280 ( .A(n6236), .B(n8674), .ZN(n8667) );
  NAND2_X1 U6281 ( .A1(n6230), .A2(n4837), .ZN(n4834) );
  NAND2_X1 U6282 ( .A1(n4835), .A2(n4834), .ZN(n7760) );
  INV_X1 U6283 ( .A(n7761), .ZN(n4837) );
  NAND2_X1 U6284 ( .A1(n6220), .A2(n4842), .ZN(n4838) );
  OAI21_X1 U6285 ( .B1(n8634), .B2(n4844), .A(n4843), .ZN(n8650) );
  INV_X1 U6286 ( .A(n4854), .ZN(n6172) );
  NAND2_X1 U6287 ( .A1(n4854), .A2(n8539), .ZN(n8798) );
  NOR2_X1 U6288 ( .A1(n4854), .A2(n8819), .ZN(n6030) );
  AOI21_X1 U6289 ( .B1(n4854), .B2(n8918), .A(n4853), .ZN(n8811) );
  AOI21_X1 U6290 ( .B1(n4854), .B2(n8576), .A(n8463), .ZN(n8464) );
  XNOR2_X1 U6291 ( .A(n4854), .B(n8186), .ZN(n8169) );
  NAND2_X1 U6292 ( .A1(n5164), .A2(n5163), .ZN(n4858) );
  NAND3_X1 U6293 ( .A1(n8377), .A2(n8402), .A3(n8376), .ZN(n4860) );
  NAND2_X1 U6294 ( .A1(n5113), .A2(n4862), .ZN(n4861) );
  NAND2_X1 U6295 ( .A1(n4861), .A2(n4864), .ZN(n5453) );
  NAND2_X1 U6296 ( .A1(n5113), .A2(n5112), .ZN(n5421) );
  NOR2_X1 U6297 ( .A1(n5419), .A2(n5420), .ZN(n4870) );
  NAND2_X1 U6298 ( .A1(n5068), .A2(n4871), .ZN(n4875) );
  NAND2_X1 U6299 ( .A1(n5068), .A2(n4880), .ZN(n4879) );
  NAND2_X1 U6300 ( .A1(n5348), .A2(n4885), .ZN(n4883) );
  NAND2_X1 U6301 ( .A1(n4883), .A2(n4489), .ZN(n5101) );
  OR2_X1 U6302 ( .A1(n5348), .A2(n5089), .ZN(n4887) );
  NAND2_X1 U6303 ( .A1(n7412), .A2(n4891), .ZN(n4890) );
  OAI21_X1 U6304 ( .B1(n7489), .B2(n4898), .A(n4896), .ZN(n7333) );
  NAND2_X1 U6305 ( .A1(n4896), .A2(n7489), .ZN(n4895) );
  NOR2_X4 U6306 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n5151) );
  NAND3_X1 U6307 ( .A1(n5151), .A2(n5173), .A3(n4914), .ZN(n5201) );
  NAND4_X1 U6308 ( .A1(n5151), .A2(n5173), .A3(n4914), .A4(n5003), .ZN(n5203)
         );
  NOR2_X2 U6309 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_4__SCAN_IN), .ZN(
        n4914) );
  NAND2_X1 U6310 ( .A1(n4916), .A2(n4915), .ZN(n5417) );
  NAND2_X1 U6311 ( .A1(n6128), .A2(n4491), .ZN(n6130) );
  INV_X1 U6312 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n4922) );
  NAND2_X1 U6313 ( .A1(n8514), .A2(n4429), .ZN(n4924) );
  NAND2_X1 U6314 ( .A1(n8166), .A2(n4929), .ZN(n4928) );
  OAI21_X1 U6315 ( .B1(n7670), .B2(n4494), .A(n4438), .ZN(n4938) );
  NOR2_X1 U6316 ( .A1(n7670), .A2(n7669), .ZN(n7672) );
  NAND2_X1 U6317 ( .A1(n8438), .A2(n4945), .ZN(n4944) );
  OAI211_X1 U6318 ( .C1(n8438), .C2(n4946), .A(n4944), .B(n8193), .ZN(P2_U3160) );
  OR2_X1 U6319 ( .A1(n8438), .A2(n8439), .ZN(n8440) );
  NOR2_X1 U6320 ( .A1(n5820), .A2(n4956), .ZN(n4955) );
  INV_X1 U6321 ( .A(n4955), .ZN(n5937) );
  NAND2_X1 U6322 ( .A1(n8572), .A2(n4419), .ZN(n4960) );
  NAND2_X1 U6323 ( .A1(n4960), .A2(n4962), .ZN(n8158) );
  INV_X1 U6324 ( .A(n4965), .ZN(n8494) );
  NAND2_X1 U6325 ( .A1(n4469), .A2(n7280), .ZN(n4967) );
  NAND2_X1 U6326 ( .A1(n7280), .A2(n4968), .ZN(n4970) );
  NAND2_X1 U6327 ( .A1(n4967), .A2(n4966), .ZN(n7573) );
  NAND2_X1 U6328 ( .A1(n7280), .A2(n7279), .ZN(n7281) );
  INV_X1 U6329 ( .A(n4970), .ZN(n7465) );
  INV_X1 U6330 ( .A(n7279), .ZN(n4971) );
  NAND2_X1 U6331 ( .A1(n5490), .A2(n5489), .ZN(n5507) );
  NOR2_X1 U6332 ( .A1(n7150), .A2(n6419), .ZN(n7148) );
  NAND2_X1 U6333 ( .A1(n6391), .A2(n6390), .ZN(n8749) );
  NOR2_X1 U6334 ( .A1(n8707), .A2(n8706), .ZN(n8713) );
  NAND2_X1 U6335 ( .A1(n6314), .A2(n6313), .ZN(n6315) );
  XNOR2_X1 U6336 ( .A(n5528), .B(n5527), .ZN(n8125) );
  NAND2_X1 U6337 ( .A1(n6673), .A2(n6818), .ZN(n9411) );
  AOI21_X1 U6338 ( .B1(n8182), .B2(n7206), .A(n7205), .ZN(n7268) );
  NAND2_X1 U6339 ( .A1(n7146), .A2(n5141), .ZN(n7089) );
  OAI21_X2 U6340 ( .B1(n8391), .B2(n4567), .A(n4568), .ZN(n8409) );
  OR2_X1 U6341 ( .A1(n5718), .A2(n5715), .ZN(n5720) );
  NAND2_X1 U6342 ( .A1(n9646), .A2(n9903), .ZN(n9655) );
  NAND2_X1 U6343 ( .A1(n6427), .A2(n6508), .ZN(n6430) );
  NAND2_X2 U6344 ( .A1(n5707), .A2(n8431), .ZN(n5774) );
  INV_X1 U6345 ( .A(n5021), .ZN(n5022) );
  NAND2_X1 U6346 ( .A1(n5548), .A2(n5547), .ZN(n5565) );
  INV_X1 U6347 ( .A(n5677), .ZN(n5678) );
  NAND2_X1 U6348 ( .A1(n8260), .A2(n8262), .ZN(n8268) );
  AND2_X1 U6349 ( .A1(n8416), .A2(n8415), .ZN(n8417) );
  XNOR2_X1 U6350 ( .A(n7209), .B(n9961), .ZN(n7207) );
  NAND2_X1 U6351 ( .A1(n8432), .A2(n5708), .ZN(n5757) );
  INV_X1 U6352 ( .A(n8432), .ZN(n5707) );
  AOI21_X2 U6353 ( .B1(n9599), .B2(n5389), .A(n5388), .ZN(n9580) );
  OR2_X1 U6354 ( .A1(n6436), .A2(n6435), .ZN(n4975) );
  AND2_X1 U6355 ( .A1(n8013), .A2(n8012), .ZN(n4976) );
  OR2_X1 U6356 ( .A1(n6493), .A2(n9201), .ZN(n4977) );
  INV_X1 U6357 ( .A(n6316), .ZN(n9937) );
  INV_X1 U6358 ( .A(n6107), .ZN(n6243) );
  INV_X1 U6359 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n6317) );
  AND4_X1 U6360 ( .A1(n5697), .A2(n5696), .A3(n5695), .A4(n5694), .ZN(n4978)
         );
  NOR2_X1 U6361 ( .A1(n5713), .A2(n5701), .ZN(n4979) );
  AND3_X1 U6362 ( .A1(n5387), .A2(n5386), .A3(n5385), .ZN(n9592) );
  INV_X1 U6363 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6217) );
  AND2_X1 U6364 ( .A1(n7016), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n4980) );
  AND2_X1 U6365 ( .A1(n7464), .A2(n7468), .ZN(n4981) );
  NAND2_X1 U6366 ( .A1(n10016), .A2(n10015), .ZN(n9013) );
  INV_X1 U6367 ( .A(n9013), .ZN(n6396) );
  AND2_X1 U6368 ( .A1(n6398), .A2(n6397), .ZN(n4982) );
  OR2_X1 U6369 ( .A1(n8759), .A2(n8950), .ZN(n4983) );
  OR2_X1 U6370 ( .A1(n9586), .A2(n10056), .ZN(n4984) );
  AND2_X1 U6371 ( .A1(n8142), .A2(n8584), .ZN(n4985) );
  AND2_X1 U6372 ( .A1(n7208), .A2(n7269), .ZN(n4986) );
  OR2_X1 U6373 ( .A1(n8759), .A2(n9013), .ZN(n4987) );
  OR2_X1 U6374 ( .A1(n9658), .A2(n9247), .ZN(n4988) );
  OR2_X1 U6375 ( .A1(n5687), .A2(n9644), .ZN(n4989) );
  AND2_X1 U6376 ( .A1(n5579), .A2(n5578), .ZN(n4990) );
  AND2_X1 U6377 ( .A1(n10290), .A2(n5014), .ZN(n4991) );
  AND2_X1 U6378 ( .A1(n6452), .A2(n6451), .ZN(n4992) );
  AND4_X1 U6379 ( .A1(n5578), .A2(n5392), .A3(n5377), .A4(n5612), .ZN(n4993)
         );
  INV_X1 U6380 ( .A(n9755), .ZN(n5657) );
  INV_X1 U6381 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n5032) );
  NAND2_X1 U6382 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), 
        .ZN(n4994) );
  AND2_X1 U6383 ( .A1(n5067), .A2(n5066), .ZN(n4995) );
  INV_X1 U6384 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5705) );
  AND2_X1 U6385 ( .A1(n6439), .A2(n6438), .ZN(n4996) );
  OR2_X1 U6386 ( .A1(n8401), .A2(n8443), .ZN(n4997) );
  AND2_X1 U6387 ( .A1(n6089), .A2(n6088), .ZN(n8443) );
  INV_X1 U6388 ( .A(n4413), .ZN(n5257) );
  OR2_X1 U6389 ( .A1(n9792), .A2(n9610), .ZN(n4998) );
  AND2_X1 U6390 ( .A1(n6890), .A2(n6426), .ZN(n4999) );
  AND2_X1 U6391 ( .A1(n6369), .A2(n8967), .ZN(n5000) );
  OR2_X1 U6392 ( .A1(n9262), .A2(n7322), .ZN(n5001) );
  OR2_X1 U6393 ( .A1(n9261), .A2(n7493), .ZN(n5002) );
  OAI21_X1 U6394 ( .B1(n6791), .B2(n6790), .A(n6789), .ZN(n6792) );
  INV_X1 U6395 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5578) );
  INV_X1 U6396 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n6335) );
  INV_X1 U6397 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n6226) );
  INV_X1 U6398 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5014) );
  NOR2_X1 U6399 ( .A1(n6316), .A2(n6217), .ZN(n6218) );
  OR2_X1 U6400 ( .A1(n5764), .A2(n4695), .ZN(n5725) );
  NAND2_X1 U6401 ( .A1(n6428), .A2(n4417), .ZN(n6429) );
  NAND2_X1 U6402 ( .A1(n6508), .A2(n6414), .ZN(n6415) );
  INV_X1 U6403 ( .A(n9685), .ZN(n5655) );
  INV_X1 U6404 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n5095) );
  NAND2_X1 U6405 ( .A1(n7992), .A2(n8587), .ZN(n7993) );
  INV_X1 U6406 ( .A(n8908), .ZN(n8147) );
  INV_X1 U6407 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n5812) );
  OAI22_X1 U6408 ( .A1(n8866), .A2(n5974), .B1(n8881), .B2(n8956), .ZN(n8851)
         );
  INV_X1 U6409 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5837) );
  INV_X1 U6410 ( .A(n8775), .ZN(n8178) );
  NOR2_X1 U6411 ( .A1(n6545), .A2(n6544), .ZN(n6546) );
  AND2_X1 U6412 ( .A1(n5025), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n5425) );
  INV_X1 U6413 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n5339) );
  AND2_X1 U6414 ( .A1(n5254), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n5272) );
  INV_X1 U6415 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5015) );
  INV_X1 U6416 ( .A(n5435), .ZN(n5436) );
  INV_X1 U6417 ( .A(SI_8_), .ZN(n10062) );
  AND2_X1 U6418 ( .A1(n7668), .A2(n8590), .ZN(n7669) );
  INV_X1 U6419 ( .A(n7277), .ZN(n7278) );
  OR2_X1 U6420 ( .A1(n6083), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n6100) );
  INV_X1 U6421 ( .A(n8208), .ZN(n6060) );
  INV_X1 U6422 ( .A(n6228), .ZN(n6229) );
  AOI21_X1 U6423 ( .B1(P2_REG2_REG_14__SCAN_IN), .B2(n7016), .A(n8658), .ZN(
        n6340) );
  INV_X1 U6424 ( .A(n6049), .ZN(n6048) );
  NAND2_X1 U6425 ( .A1(n5900), .A2(n5899), .ZN(n5918) );
  NAND2_X1 U6426 ( .A1(n5838), .A2(n5837), .ZN(n5853) );
  OR2_X1 U6427 ( .A1(n6132), .A2(P2_D_REG_1__SCAN_IN), .ZN(n6135) );
  OAI21_X1 U6428 ( .B1(n8755), .B2(n9939), .A(n6388), .ZN(n6389) );
  OR2_X1 U6429 ( .A1(n9037), .A2(n8454), .ZN(n8338) );
  OR2_X1 U6430 ( .A1(n8402), .A2(n7198), .ZN(n7355) );
  OR2_X1 U6431 ( .A1(n5321), .A2(n10341), .ZN(n5340) );
  AND2_X1 U6432 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n5180) );
  OR2_X1 U6433 ( .A1(n5539), .A2(n5538), .ZN(n5556) );
  OR2_X1 U6434 ( .A1(n5367), .A2(n9131), .ZN(n9143) );
  INV_X1 U6435 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n10341) );
  INV_X1 U6436 ( .A(n5462), .ZN(n5479) );
  NAND2_X1 U6437 ( .A1(n7989), .A2(n7962), .ZN(n5313) );
  OR2_X1 U6438 ( .A1(n9173), .A2(n9257), .ZN(n5262) );
  INV_X1 U6439 ( .A(n9567), .ZN(n9628) );
  OR2_X1 U6440 ( .A1(n6623), .A2(n6622), .ZN(n6624) );
  NAND2_X1 U6441 ( .A1(n5530), .A2(n5529), .ZN(n5546) );
  INV_X1 U6442 ( .A(SI_12_), .ZN(n5078) );
  OR2_X1 U6443 ( .A1(n5267), .A2(n5266), .ZN(n5282) );
  INV_X1 U6444 ( .A(n8881), .ZN(n8509) );
  OR2_X1 U6445 ( .A1(n5968), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5983) );
  NAND2_X1 U6446 ( .A1(n7122), .A2(n7212), .ZN(n8566) );
  OR2_X1 U6447 ( .A1(n5757), .A2(n6214), .ZN(n5742) );
  AND2_X1 U6448 ( .A1(n8711), .A2(n8710), .ZN(n8712) );
  NAND2_X1 U6449 ( .A1(n6048), .A2(n6047), .ZN(n6058) );
  OR2_X1 U6450 ( .A1(n8071), .A2(n8063), .ZN(n8317) );
  NAND2_X1 U6451 ( .A1(n6159), .A2(n6158), .ZN(n8270) );
  NAND2_X1 U6452 ( .A1(n6135), .A2(n6134), .ZN(n6199) );
  NAND2_X1 U6453 ( .A1(n6111), .A2(n6110), .ZN(n6112) );
  OR2_X1 U6454 ( .A1(n8784), .A2(n8374), .ZN(n8804) );
  AND2_X1 U6455 ( .A1(n8348), .A2(n8338), .ZN(n8905) );
  INV_X1 U6456 ( .A(n9953), .ZN(n8909) );
  INV_X1 U6457 ( .A(n8586), .ZN(n8006) );
  INV_X1 U6458 ( .A(n8912), .ZN(n9949) );
  AND2_X1 U6459 ( .A1(n6543), .A2(n6542), .ZN(n9214) );
  INV_X1 U6460 ( .A(n9225), .ZN(n9241) );
  AND2_X1 U6461 ( .A1(n6679), .A2(P1_STATE_REG_SCAN_IN), .ZN(n5664) );
  INV_X1 U6462 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n9131) );
  AND2_X1 U6463 ( .A1(n6779), .A2(n6777), .ZN(n9574) );
  NOR2_X1 U6464 ( .A1(n9059), .A2(n9252), .ZN(n5346) );
  NAND2_X1 U6465 ( .A1(n9651), .A2(n9650), .ZN(n9652) );
  INV_X1 U6466 ( .A(n9703), .ZN(n9558) );
  NOR2_X1 U6467 ( .A1(n9625), .A2(n9724), .ZN(n5388) );
  OR2_X1 U6468 ( .A1(n9877), .A2(n6680), .ZN(n9899) );
  OR2_X1 U6469 ( .A1(n9877), .A2(n6678), .ZN(n9567) );
  AND2_X1 U6470 ( .A1(n6598), .A2(n5614), .ZN(n5662) );
  INV_X1 U6471 ( .A(n8571), .ZN(n8545) );
  AND2_X1 U6472 ( .A1(n6055), .A2(n6054), .ZN(n8176) );
  AND4_X1 U6473 ( .A1(n5960), .A2(n5959), .A3(n5958), .A4(n5957), .ZN(n8896)
         );
  OR2_X1 U6474 ( .A1(n10005), .A2(n6358), .ZN(n9944) );
  INV_X1 U6475 ( .A(n9994), .ZN(n7785) );
  INV_X1 U6476 ( .A(n9943), .ZN(n8917) );
  INV_X1 U6477 ( .A(n8922), .ZN(n8848) );
  AND2_X1 U6478 ( .A1(n10029), .A2(n9970), .ZN(n8967) );
  OR2_X1 U6479 ( .A1(n7204), .A2(n6199), .ZN(n7104) );
  NOR2_X1 U6480 ( .A1(n10017), .A2(n10010), .ZN(n9038) );
  NAND2_X1 U6481 ( .A1(n9939), .A2(n10000), .ZN(n9970) );
  XNOR2_X1 U6482 ( .A(n6152), .B(n10253), .ZN(n7097) );
  XNOR2_X1 U6483 ( .A(n6098), .B(P2_IR_REG_22__SCAN_IN), .ZN(n8425) );
  INV_X1 U6484 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5807) );
  AND2_X1 U6485 ( .A1(n6915), .A2(P2_U3151), .ZN(n9044) );
  AND2_X1 U6486 ( .A1(n6612), .A2(n9723), .ZN(n9225) );
  AND2_X1 U6487 ( .A1(n9142), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9229) );
  AOI21_X1 U6488 ( .B1(n6839), .B2(n5666), .A(n6838), .ZN(n6840) );
  AND4_X1 U6489 ( .A1(n5562), .A2(n5561), .A3(n5560), .A4(n5559), .ZN(n9432)
         );
  AND4_X1 U6490 ( .A1(n5416), .A2(n5415), .A3(n5414), .A4(n5413), .ZN(n9706)
         );
  AND4_X1 U6491 ( .A1(n5326), .A2(n5325), .A3(n5324), .A4(n5323), .ZN(n8114)
         );
  OR3_X1 U6492 ( .A1(n6881), .A2(n8195), .A3(n5643), .ZN(n9844) );
  INV_X1 U6493 ( .A(n9844), .ZN(n9872) );
  NAND2_X1 U6494 ( .A1(n5678), .A2(n9560), .ZN(n5679) );
  INV_X1 U6495 ( .A(n9574), .ZN(n9564) );
  AND2_X1 U6496 ( .A1(n5644), .A2(n6899), .ZN(n9723) );
  INV_X1 U6497 ( .A(n9489), .ZN(n9578) );
  INV_X1 U6498 ( .A(n9591), .ZN(n9881) );
  AND2_X1 U6499 ( .A1(n9910), .A2(n9903), .ZN(n9711) );
  NAND2_X1 U6500 ( .A1(n6821), .A2(n5657), .ZN(n5658) );
  INV_X1 U6501 ( .A(n9460), .ZN(n9457) );
  AND2_X1 U6502 ( .A1(n6787), .A2(n6788), .ZN(n9528) );
  AND2_X1 U6503 ( .A1(n9906), .A2(n9903), .ZN(n9786) );
  NAND2_X1 U6504 ( .A1(n5668), .A2(n5620), .ZN(n9903) );
  NAND2_X1 U6505 ( .A1(n5588), .A2(n5587), .ZN(n9809) );
  AND2_X1 U6506 ( .A1(n5335), .A2(n5334), .ZN(n9324) );
  INV_X1 U6507 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n10126) );
  INV_X1 U6508 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n10339) );
  INV_X1 U6509 ( .A(n8576), .ZN(n8554) );
  AND2_X1 U6510 ( .A1(n7118), .A2(n7117), .ZN(n8571) );
  NAND2_X1 U6511 ( .A1(n6066), .A2(n6065), .ZN(n8775) );
  AND2_X1 U6512 ( .A1(n6297), .A2(n6296), .ZN(n9938) );
  INV_X1 U6513 ( .A(n8737), .ZN(n9930) );
  OR2_X1 U6514 ( .A1(n6361), .A2(n9944), .ZN(n8846) );
  OR2_X1 U6515 ( .A1(n6361), .A2(n6359), .ZN(n9956) );
  AND2_X1 U6516 ( .A1(n6360), .A2(n9956), .ZN(n8922) );
  NAND2_X1 U6517 ( .A1(n10029), .A2(n10015), .ZN(n8950) );
  INV_X1 U6518 ( .A(n10029), .ZN(n10027) );
  INV_X1 U6519 ( .A(n8478), .ZN(n9009) );
  INV_X1 U6520 ( .A(n9038), .ZN(n9022) );
  AND2_X1 U6521 ( .A1(n6203), .A2(n6202), .ZN(n10017) );
  AND2_X1 U6522 ( .A1(n7109), .A2(n6132), .ZN(n6958) );
  AND2_X1 U6523 ( .A1(n7097), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8135) );
  INV_X1 U6524 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n10301) );
  INV_X1 U6525 ( .A(n9875), .ZN(n9352) );
  INV_X1 U6526 ( .A(n9696), .ZN(n9536) );
  INV_X1 U6527 ( .A(n9236), .ZN(n9205) );
  INV_X1 U6528 ( .A(n9792), .ZN(n9586) );
  NAND2_X1 U6529 ( .A1(n6841), .A2(n6840), .ZN(n6868) );
  NAND4_X1 U6530 ( .A1(n5031), .A2(n5030), .A3(n5029), .A4(n5028), .ZN(n9695)
         );
  INV_X1 U6531 ( .A(n9592), .ZN(n9625) );
  INV_X1 U6532 ( .A(n7588), .ZN(n9258) );
  INV_X1 U6533 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n9858) );
  INV_X1 U6534 ( .A(n9386), .ZN(n9869) );
  OR2_X1 U6535 ( .A1(n6881), .A2(n6899), .ZN(n9866) );
  INV_X1 U6536 ( .A(n9446), .ZN(n9637) );
  INV_X2 U6537 ( .A(n9560), .ZN(n9889) );
  NAND2_X1 U6538 ( .A1(n9910), .A2(n9745), .ZN(n9644) );
  INV_X1 U6539 ( .A(n9910), .ZN(n9908) );
  NAND2_X1 U6540 ( .A1(n9906), .A2(n9745), .ZN(n9755) );
  INV_X1 U6541 ( .A(n9906), .ZN(n9905) );
  AND2_X2 U6542 ( .A1(n5683), .A2(n5663), .ZN(n9906) );
  INV_X1 U6543 ( .A(n9891), .ZN(n9890) );
  AND2_X1 U6544 ( .A1(n9809), .A2(n9808), .ZN(n9891) );
  INV_X1 U6545 ( .A(n6843), .ZN(n7849) );
  INV_X1 U6546 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n7266) );
  INV_X1 U6547 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6950) );
  INV_X1 U6548 ( .A(n8727), .ZN(P2_U3893) );
  INV_X1 U6549 ( .A(n10054), .ZN(P1_U3973) );
  NOR2_X1 U6550 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n5005) );
  NAND4_X1 U6551 ( .A1(n5005), .A2(n5004), .A3(n5265), .A4(n5264), .ZN(n5006)
         );
  NOR2_X2 U6552 ( .A1(n5203), .A2(n5006), .ZN(n5297) );
  NOR2_X1 U6553 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_24__SCAN_IN), .ZN(
        n5012) );
  NOR2_X1 U6554 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_25__SCAN_IN), .ZN(
        n5011) );
  NAND4_X1 U6555 ( .A1(n4993), .A2(n4478), .A3(n5012), .A4(n5011), .ZN(n5013)
         );
  NAND2_X1 U6556 ( .A1(n5119), .A2(n5019), .ZN(n9813) );
  NAND2_X1 U6557 ( .A1(n5257), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n5031) );
  INV_X1 U6558 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n10333) );
  OR2_X1 U6559 ( .A1(n5308), .A2(n10333), .ZN(n5030) );
  INV_X1 U6560 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n9552) );
  OR2_X1 U6561 ( .A1(n5649), .A2(n9552), .ZN(n5029) );
  NAND2_X2 U6562 ( .A1(n5023), .A2(n5022), .ZN(n5446) );
  NAND2_X1 U6563 ( .A1(n5180), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n5212) );
  NOR2_X1 U6564 ( .A1(n5212), .A2(n5211), .ZN(n5210) );
  NAND2_X1 U6565 ( .A1(n5210), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5241) );
  NAND2_X1 U6566 ( .A1(n5338), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n5367) );
  NAND2_X1 U6567 ( .A1(n5397), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n5409) );
  INV_X1 U6568 ( .A(n5409), .ZN(n5024) );
  INV_X1 U6569 ( .A(n5425), .ZN(n5427) );
  INV_X1 U6570 ( .A(n5025), .ZN(n5412) );
  INV_X1 U6571 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n5026) );
  NAND2_X1 U6572 ( .A1(n5412), .A2(n5026), .ZN(n5027) );
  NAND2_X1 U6573 ( .A1(n5427), .A2(n5027), .ZN(n9551) );
  OR2_X1 U6574 ( .A1(n5572), .A2(n9551), .ZN(n5028) );
  INV_X1 U6575 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6918) );
  NAND3_X1 U6576 ( .A1(n5122), .A2(SI_0_), .A3(P2_DATAO_REG_0__SCAN_IN), .ZN(
        n5034) );
  INV_X1 U6577 ( .A(n5122), .ZN(n5732) );
  AND2_X1 U6578 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n5033) );
  NAND2_X1 U6579 ( .A1(n5732), .A2(n5033), .ZN(n5735) );
  NAND2_X1 U6580 ( .A1(n5034), .A2(n5735), .ZN(n5126) );
  INV_X1 U6581 ( .A(n5035), .ZN(n5036) );
  NAND2_X1 U6582 ( .A1(n5036), .A2(SI_1_), .ZN(n5037) );
  NAND2_X1 U6583 ( .A1(n5038), .A2(n5037), .ZN(n5153) );
  INV_X1 U6584 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6913) );
  INV_X1 U6585 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6924) );
  XNOR2_X1 U6586 ( .A(n5040), .B(SI_2_), .ZN(n5152) );
  NAND2_X1 U6587 ( .A1(n5153), .A2(n5152), .ZN(n5043) );
  INV_X1 U6588 ( .A(n5040), .ZN(n5041) );
  NAND2_X1 U6589 ( .A1(n5041), .A2(SI_2_), .ZN(n5042) );
  NAND2_X1 U6590 ( .A1(n5043), .A2(n5042), .ZN(n5164) );
  INV_X1 U6591 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n10272) );
  INV_X1 U6592 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6921) );
  MUX2_X1 U6593 ( .A(n10272), .B(n6921), .S(n5122), .Z(n5044) );
  XNOR2_X1 U6594 ( .A(n5044), .B(SI_3_), .ZN(n5163) );
  INV_X1 U6595 ( .A(n5044), .ZN(n5045) );
  NAND2_X1 U6596 ( .A1(n5045), .A2(SI_3_), .ZN(n5046) );
  INV_X1 U6597 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n10270) );
  INV_X1 U6598 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6932) );
  INV_X1 U6599 ( .A(n5047), .ZN(n5048) );
  MUX2_X1 U6600 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n5122), .Z(n5050) );
  INV_X1 U6601 ( .A(SI_5_), .ZN(n5049) );
  XNOR2_X1 U6602 ( .A(n5050), .B(n5049), .ZN(n5190) );
  INV_X1 U6603 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6928) );
  BUF_X4 U6604 ( .A(n5122), .Z(n6915) );
  MUX2_X1 U6605 ( .A(n10343), .B(n6928), .S(n6915), .Z(n5051) );
  XNOR2_X1 U6606 ( .A(n5051), .B(SI_6_), .ZN(n5206) );
  NAND2_X1 U6607 ( .A1(n5207), .A2(n5206), .ZN(n5054) );
  INV_X1 U6608 ( .A(n5051), .ZN(n5052) );
  NAND2_X1 U6609 ( .A1(n5052), .A2(SI_6_), .ZN(n5053) );
  NAND2_X1 U6610 ( .A1(n5054), .A2(n5053), .ZN(n5221) );
  INV_X1 U6611 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6919) );
  INV_X1 U6612 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6926) );
  MUX2_X1 U6613 ( .A(n6919), .B(n6926), .S(n6915), .Z(n5055) );
  XNOR2_X1 U6614 ( .A(n5055), .B(SI_7_), .ZN(n5220) );
  NAND2_X1 U6615 ( .A1(n5221), .A2(n5220), .ZN(n5058) );
  INV_X1 U6616 ( .A(n5055), .ZN(n5056) );
  NAND2_X1 U6617 ( .A1(n5056), .A2(SI_7_), .ZN(n5057) );
  INV_X1 U6618 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6936) );
  INV_X1 U6619 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n6934) );
  MUX2_X1 U6620 ( .A(n6936), .B(n6934), .S(n6915), .Z(n5059) );
  NAND2_X1 U6621 ( .A1(n5059), .A2(n10062), .ZN(n5062) );
  INV_X1 U6622 ( .A(n5059), .ZN(n5060) );
  NAND2_X1 U6623 ( .A1(n5060), .A2(SI_8_), .ZN(n5061) );
  NAND2_X1 U6624 ( .A1(n5062), .A2(n5061), .ZN(n5234) );
  INV_X1 U6625 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6938) );
  MUX2_X1 U6626 ( .A(n6938), .B(n6941), .S(n6915), .Z(n5064) );
  INV_X1 U6627 ( .A(SI_9_), .ZN(n5063) );
  NAND2_X1 U6628 ( .A1(n5064), .A2(n5063), .ZN(n5067) );
  INV_X1 U6629 ( .A(n5064), .ZN(n5065) );
  NAND2_X1 U6630 ( .A1(n5065), .A2(SI_9_), .ZN(n5066) );
  MUX2_X1 U6631 ( .A(n10277), .B(n10285), .S(n6915), .Z(n5069) );
  XNOR2_X1 U6632 ( .A(n5069), .B(SI_10_), .ZN(n5263) );
  INV_X1 U6633 ( .A(n5263), .ZN(n5072) );
  INV_X1 U6634 ( .A(n5069), .ZN(n5070) );
  NAND2_X1 U6635 ( .A1(n5070), .A2(SI_10_), .ZN(n5071) );
  MUX2_X1 U6636 ( .A(n10300), .B(n6950), .S(n6915), .Z(n5074) );
  INV_X1 U6637 ( .A(SI_11_), .ZN(n5073) );
  NAND2_X1 U6638 ( .A1(n5074), .A2(n5073), .ZN(n5077) );
  INV_X1 U6639 ( .A(n5074), .ZN(n5075) );
  NAND2_X1 U6640 ( .A1(n5075), .A2(SI_11_), .ZN(n5076) );
  NAND2_X1 U6641 ( .A1(n5077), .A2(n5076), .ZN(n5280) );
  MUX2_X1 U6642 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .S(n6915), .Z(n5079) );
  XNOR2_X1 U6643 ( .A(n5079), .B(n5078), .ZN(n5295) );
  INV_X1 U6644 ( .A(n5295), .ZN(n5080) );
  MUX2_X1 U6645 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n6915), .Z(n5082) );
  XNOR2_X1 U6646 ( .A(n5082), .B(SI_13_), .ZN(n5314) );
  INV_X1 U6647 ( .A(n5314), .ZN(n5081) );
  NAND2_X1 U6648 ( .A1(n5315), .A2(n5081), .ZN(n5084) );
  NAND2_X1 U6649 ( .A1(n5082), .A2(SI_13_), .ZN(n5083) );
  NAND2_X1 U6650 ( .A1(n5084), .A2(n5083), .ZN(n5328) );
  MUX2_X1 U6651 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n6915), .Z(n5086) );
  XNOR2_X1 U6652 ( .A(n5086), .B(SI_14_), .ZN(n5329) );
  INV_X1 U6653 ( .A(n5329), .ZN(n5085) );
  NAND2_X1 U6654 ( .A1(n5328), .A2(n5085), .ZN(n5088) );
  NAND2_X1 U6655 ( .A1(n5086), .A2(SI_14_), .ZN(n5087) );
  MUX2_X1 U6656 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .S(n6915), .Z(n5349) );
  NOR2_X1 U6657 ( .A1(n5091), .A2(n5090), .ZN(n5089) );
  NAND2_X1 U6658 ( .A1(n5091), .A2(n5090), .ZN(n5092) );
  MUX2_X1 U6659 ( .A(n10164), .B(n7169), .S(n6915), .Z(n5361) );
  NOR2_X1 U6660 ( .A1(n5093), .A2(SI_16_), .ZN(n5094) );
  MUX2_X1 U6661 ( .A(n5095), .B(n7266), .S(n6915), .Z(n5097) );
  NAND2_X1 U6662 ( .A1(n5097), .A2(n5096), .ZN(n5100) );
  INV_X1 U6663 ( .A(n5097), .ZN(n5098) );
  NAND2_X1 U6664 ( .A1(n5098), .A2(SI_17_), .ZN(n5099) );
  NAND2_X1 U6665 ( .A1(n5100), .A2(n5099), .ZN(n5375) );
  NAND2_X1 U6666 ( .A1(n5101), .A2(n5100), .ZN(n5391) );
  MUX2_X1 U6667 ( .A(n10055), .B(n5102), .S(n6915), .Z(n5103) );
  XNOR2_X1 U6668 ( .A(n5103), .B(SI_18_), .ZN(n5390) );
  INV_X1 U6669 ( .A(n5390), .ZN(n5106) );
  INV_X1 U6670 ( .A(n5103), .ZN(n5104) );
  NAND2_X1 U6671 ( .A1(n5104), .A2(SI_18_), .ZN(n5105) );
  INV_X1 U6672 ( .A(n5403), .ZN(n5111) );
  MUX2_X1 U6673 ( .A(n7546), .B(n7548), .S(n6915), .Z(n5107) );
  NAND2_X1 U6674 ( .A1(n5107), .A2(n10094), .ZN(n5112) );
  INV_X1 U6675 ( .A(n5107), .ZN(n5108) );
  NAND2_X1 U6676 ( .A1(n5108), .A2(SI_19_), .ZN(n5109) );
  NAND2_X1 U6677 ( .A1(n5112), .A2(n5109), .ZN(n5402) );
  INV_X1 U6678 ( .A(n5402), .ZN(n5110) );
  NAND2_X1 U6679 ( .A1(n5111), .A2(n5110), .ZN(n5113) );
  MUX2_X1 U6680 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(P2_DATAO_REG_20__SCAN_IN), 
        .S(n6915), .Z(n5418) );
  XNOR2_X1 U6681 ( .A(n5418), .B(n5420), .ZN(n5114) );
  NAND2_X1 U6682 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_26__SCAN_IN), 
        .ZN(n5116) );
  NAND2_X4 U6683 ( .A1(n5643), .A2(n5650), .ZN(n6873) );
  NAND2_X1 U6684 ( .A1(n7648), .A2(n6635), .ZN(n5124) );
  NAND2_X1 U6685 ( .A1(n5535), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n5123) );
  INV_X1 U6686 ( .A(n5151), .ZN(n5125) );
  OR2_X1 U6687 ( .A1(n4414), .A2(n6918), .ZN(n5129) );
  XNOR2_X1 U6688 ( .A(n5127), .B(n5126), .ZN(n6917) );
  OR2_X1 U6689 ( .A1(n4415), .A2(n6917), .ZN(n5128) );
  NAND2_X1 U6690 ( .A1(n5146), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5134) );
  INV_X1 U6691 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n7394) );
  INV_X1 U6692 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n5130) );
  INV_X1 U6693 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n6878) );
  OR2_X1 U6694 ( .A1(n5144), .A2(n6878), .ZN(n5131) );
  XNOR2_X1 U6695 ( .A(n9103), .B(n6427), .ZN(n5623) );
  NAND2_X1 U6696 ( .A1(n6915), .A2(SI_0_), .ZN(n5135) );
  XNOR2_X1 U6697 ( .A(n5135), .B(P2_DATAO_REG_0__SCAN_IN), .ZN(n9825) );
  MUX2_X1 U6698 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9825), .S(n6873), .Z(n9879) );
  INV_X1 U6699 ( .A(n9879), .ZN(n7150) );
  INV_X1 U6700 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n5136) );
  INV_X1 U6701 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n7144) );
  OR2_X1 U6702 ( .A1(n5446), .A2(n7144), .ZN(n5140) );
  INV_X1 U6703 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n5137) );
  OR2_X1 U6704 ( .A1(n5369), .A2(n5137), .ZN(n5139) );
  INV_X1 U6705 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n6876) );
  OR2_X1 U6706 ( .A1(n4413), .A2(n6876), .ZN(n5138) );
  INV_X1 U6707 ( .A(n4417), .ZN(n7158) );
  INV_X1 U6708 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n5142) );
  OR2_X1 U6709 ( .A1(n5446), .A2(n5142), .ZN(n5150) );
  INV_X1 U6710 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n5143) );
  OR2_X1 U6711 ( .A1(n4413), .A2(n5143), .ZN(n5149) );
  INV_X1 U6712 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n5145) );
  OR2_X1 U6713 ( .A1(n5308), .A2(n5145), .ZN(n5148) );
  NAND2_X1 U6714 ( .A1(n5146), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5147) );
  OR2_X1 U6715 ( .A1(n5151), .A2(n9815), .ZN(n5175) );
  INV_X1 U6716 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n10275) );
  XNOR2_X1 U6717 ( .A(n5175), .B(n10275), .ZN(n6922) );
  XNOR2_X1 U6718 ( .A(n5153), .B(n5152), .ZN(n6923) );
  OR2_X1 U6719 ( .A1(n5154), .A2(n6923), .ZN(n5157) );
  OR2_X1 U6720 ( .A1(n4414), .A2(n6924), .ZN(n5156) );
  OAI211_X1 U6721 ( .C1(n6873), .C2(n6922), .A(n5157), .B(n5156), .ZN(n7175)
         );
  NAND2_X1 U6722 ( .A1(n7406), .A2(n7175), .ZN(n5626) );
  NAND2_X1 U6723 ( .A1(n6411), .A2(n9264), .ZN(n5627) );
  NAND2_X1 U6724 ( .A1(n5626), .A2(n5627), .ZN(n6687) );
  NAND2_X1 U6725 ( .A1(n7089), .A2(n6687), .ZN(n5159) );
  OR2_X1 U6726 ( .A1(n9264), .A2(n7175), .ZN(n5158) );
  NAND2_X1 U6727 ( .A1(n5159), .A2(n5158), .ZN(n7181) );
  NAND2_X1 U6728 ( .A1(n5175), .A2(n10275), .ZN(n5160) );
  NAND2_X1 U6729 ( .A1(n5160), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5162) );
  INV_X1 U6730 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n5161) );
  XNOR2_X1 U6731 ( .A(n5162), .B(n5161), .ZN(n7048) );
  XNOR2_X1 U6732 ( .A(n5164), .B(n5163), .ZN(n6920) );
  OR2_X1 U6733 ( .A1(n4415), .A2(n6920), .ZN(n5166) );
  NAND2_X1 U6734 ( .A1(n5146), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5171) );
  OR2_X1 U6735 ( .A1(n5446), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n5170) );
  INV_X1 U6736 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6995) );
  OR2_X1 U6737 ( .A1(n4413), .A2(n6995), .ZN(n5169) );
  INV_X1 U6738 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n5167) );
  OR2_X1 U6739 ( .A1(n5308), .A2(n5167), .ZN(n5168) );
  NAND2_X1 U6740 ( .A1(n6440), .A2(n9263), .ZN(n6721) );
  NAND2_X1 U6741 ( .A1(n7086), .A2(n7191), .ZN(n6713) );
  NAND2_X1 U6742 ( .A1(n7181), .A2(n7180), .ZN(n7179) );
  NAND2_X1 U6743 ( .A1(n7179), .A2(n5172), .ZN(n7220) );
  OR2_X1 U6744 ( .A1(n5173), .A2(n9815), .ZN(n5174) );
  NAND2_X1 U6745 ( .A1(n5175), .A2(n5174), .ZN(n5186) );
  XNOR2_X1 U6746 ( .A(n5186), .B(P1_IR_REG_4__SCAN_IN), .ZN(n9845) );
  XNOR2_X1 U6747 ( .A(n5177), .B(n5176), .ZN(n6931) );
  OR2_X1 U6748 ( .A1(n5154), .A2(n6931), .ZN(n5179) );
  OR2_X1 U6749 ( .A1(n5155), .A2(n6932), .ZN(n5178) );
  OAI211_X1 U6750 ( .C1(n9845), .C2(n6873), .A(n5179), .B(n5178), .ZN(n7322)
         );
  INV_X1 U6751 ( .A(n7322), .ZN(n7362) );
  NAND2_X1 U6752 ( .A1(n6639), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5184) );
  INV_X1 U6753 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6989) );
  OR2_X1 U6754 ( .A1(n5369), .A2(n6989), .ZN(n5183) );
  INV_X1 U6755 ( .A(n5180), .ZN(n5194) );
  OAI21_X1 U6756 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(n5194), .ZN(n7320) );
  OR2_X1 U6757 ( .A1(n5446), .A2(n7320), .ZN(n5182) );
  INV_X1 U6758 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n6996) );
  OR2_X1 U6759 ( .A1(n4413), .A2(n6996), .ZN(n5181) );
  NAND4_X1 U6760 ( .A1(n5184), .A2(n5183), .A3(n5182), .A4(n5181), .ZN(n9262)
         );
  INV_X1 U6761 ( .A(n9262), .ZN(n5185) );
  NAND2_X1 U6762 ( .A1(n5185), .A2(n7322), .ZN(n6714) );
  NAND2_X1 U6763 ( .A1(n6722), .A2(n6714), .ZN(n7219) );
  NAND2_X1 U6764 ( .A1(n7220), .A2(n7219), .ZN(n7218) );
  NAND2_X1 U6765 ( .A1(n7218), .A2(n5001), .ZN(n7489) );
  OAI21_X1 U6766 ( .B1(n5186), .B2(P1_IR_REG_4__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5188) );
  INV_X1 U6767 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n5187) );
  XNOR2_X1 U6768 ( .A(n5188), .B(n5187), .ZN(n9266) );
  XNOR2_X1 U6769 ( .A(n5189), .B(n5190), .ZN(n6929) );
  OR2_X1 U6770 ( .A1(n4415), .A2(n6929), .ZN(n5192) );
  INV_X1 U6771 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6930) );
  OR2_X1 U6772 ( .A1(n5155), .A2(n6930), .ZN(n5191) );
  OAI211_X1 U6773 ( .C1(n6873), .C2(n9266), .A(n5192), .B(n5191), .ZN(n7493)
         );
  INV_X1 U6774 ( .A(n7493), .ZN(n9900) );
  NAND2_X1 U6775 ( .A1(n6639), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n5200) );
  INV_X1 U6777 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n6990) );
  OR2_X1 U6778 ( .A1(n5649), .A2(n6990), .ZN(n5199) );
  INV_X1 U6779 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n5193) );
  NAND2_X1 U6780 ( .A1(n5194), .A2(n5193), .ZN(n5195) );
  NAND2_X1 U6781 ( .A1(n5212), .A2(n5195), .ZN(n7494) );
  OR2_X1 U6782 ( .A1(n5572), .A2(n7494), .ZN(n5198) );
  INV_X1 U6783 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n5196) );
  OR2_X1 U6784 ( .A1(n4413), .A2(n5196), .ZN(n5197) );
  NAND4_X1 U6785 ( .A1(n5200), .A2(n5199), .A3(n5198), .A4(n5197), .ZN(n9261)
         );
  NAND2_X1 U6786 ( .A1(n9900), .A2(n9261), .ZN(n6719) );
  INV_X1 U6787 ( .A(n9261), .ZN(n7614) );
  NAND2_X1 U6788 ( .A1(n7614), .A2(n7493), .ZN(n6717) );
  NAND2_X1 U6789 ( .A1(n6719), .A2(n6717), .ZN(n7488) );
  NAND2_X1 U6790 ( .A1(n5201), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5202) );
  MUX2_X1 U6791 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5202), .S(
        P1_IR_REG_6__SCAN_IN), .Z(n5205) );
  NAND2_X1 U6792 ( .A1(n5205), .A2(n5204), .ZN(n9285) );
  XNOR2_X1 U6793 ( .A(n5207), .B(n5206), .ZN(n6927) );
  OR2_X1 U6794 ( .A1(n6927), .A2(n5154), .ZN(n5209) );
  NAND2_X1 U6795 ( .A1(n5535), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n5208) );
  OAI211_X1 U6796 ( .C1(n6873), .C2(n9285), .A(n5209), .B(n5208), .ZN(n7616)
         );
  INV_X1 U6797 ( .A(n7616), .ZN(n7387) );
  NAND2_X1 U6798 ( .A1(n5146), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n5218) );
  INV_X1 U6799 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n6998) );
  OR2_X1 U6800 ( .A1(n4413), .A2(n6998), .ZN(n5217) );
  INV_X1 U6801 ( .A(n5210), .ZN(n5226) );
  NAND2_X1 U6802 ( .A1(n5212), .A2(n5211), .ZN(n5213) );
  NAND2_X1 U6803 ( .A1(n5226), .A2(n5213), .ZN(n7619) );
  OR2_X1 U6804 ( .A1(n5446), .A2(n7619), .ZN(n5216) );
  INV_X1 U6805 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n5214) );
  OR2_X1 U6806 ( .A1(n5308), .A2(n5214), .ZN(n5215) );
  NAND4_X1 U6807 ( .A1(n5218), .A2(n5217), .A3(n5216), .A4(n5215), .ZN(n9260)
         );
  NAND2_X1 U6808 ( .A1(n7387), .A2(n9260), .ZN(n6720) );
  INV_X1 U6809 ( .A(n9260), .ZN(n7454) );
  NAND2_X1 U6810 ( .A1(n7616), .A2(n7454), .ZN(n7418) );
  NAND2_X1 U6811 ( .A1(n6720), .A2(n7418), .ZN(n7334) );
  OR2_X1 U6812 ( .A1(n9260), .A2(n7616), .ZN(n5219) );
  XNOR2_X1 U6813 ( .A(n5221), .B(n5220), .ZN(n6925) );
  OR2_X1 U6814 ( .A1(n6925), .A2(n4415), .ZN(n5224) );
  NAND2_X1 U6815 ( .A1(n5204), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5222) );
  XNOR2_X1 U6816 ( .A(n5222), .B(P1_IR_REG_7__SCAN_IN), .ZN(n7001) );
  AOI22_X1 U6817 ( .A1(n5535), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n5406), .B2(
        n7001), .ZN(n5223) );
  NAND2_X1 U6818 ( .A1(n5224), .A2(n5223), .ZN(n7457) );
  NAND2_X1 U6819 ( .A1(n6639), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5232) );
  INV_X1 U6820 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n7424) );
  OR2_X1 U6821 ( .A1(n5369), .A2(n7424), .ZN(n5231) );
  INV_X1 U6822 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n5225) );
  NAND2_X1 U6823 ( .A1(n5226), .A2(n5225), .ZN(n5227) );
  NAND2_X1 U6824 ( .A1(n5241), .A2(n5227), .ZN(n7625) );
  OR2_X1 U6825 ( .A1(n5446), .A2(n7625), .ZN(n5230) );
  INV_X1 U6826 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n5228) );
  OR2_X1 U6827 ( .A1(n4413), .A2(n5228), .ZN(n5229) );
  OR2_X1 U6828 ( .A1(n7457), .A2(n7841), .ZN(n6735) );
  NAND2_X1 U6829 ( .A1(n7457), .A2(n7841), .ZN(n7437) );
  NAND2_X1 U6830 ( .A1(n6735), .A2(n7437), .ZN(n7413) );
  NAND2_X1 U6831 ( .A1(n7414), .A2(n7413), .ZN(n7412) );
  INV_X1 U6832 ( .A(n7841), .ZN(n9259) );
  OR2_X1 U6833 ( .A1(n9259), .A2(n7457), .ZN(n5233) );
  XNOR2_X1 U6834 ( .A(n5235), .B(n5234), .ZN(n6933) );
  NAND2_X1 U6835 ( .A1(n6933), .A2(n6635), .ZN(n5239) );
  INV_X1 U6836 ( .A(n5204), .ZN(n5237) );
  INV_X1 U6837 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n5236) );
  NAND2_X1 U6838 ( .A1(n5237), .A2(n5236), .ZN(n5267) );
  NAND2_X1 U6839 ( .A1(n5267), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5248) );
  XNOR2_X1 U6840 ( .A(n5248), .B(P1_IR_REG_8__SCAN_IN), .ZN(n7002) );
  AOI22_X1 U6841 ( .A1(n5535), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n5406), .B2(
        n7002), .ZN(n5238) );
  NAND2_X1 U6842 ( .A1(n5239), .A2(n5238), .ZN(n7839) );
  NAND2_X1 U6843 ( .A1(n5146), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n5246) );
  INV_X1 U6844 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n10312) );
  OR2_X1 U6845 ( .A1(n5308), .A2(n10312), .ZN(n5245) );
  NAND2_X1 U6846 ( .A1(n5241), .A2(n5240), .ZN(n5242) );
  NAND2_X1 U6847 ( .A1(n5255), .A2(n5242), .ZN(n7840) );
  OR2_X1 U6848 ( .A1(n5572), .A2(n7840), .ZN(n5244) );
  INV_X1 U6849 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n7003) );
  OR2_X1 U6850 ( .A1(n4413), .A2(n7003), .ZN(n5243) );
  OR2_X1 U6851 ( .A1(n7839), .A2(n7588), .ZN(n7583) );
  NAND2_X1 U6852 ( .A1(n7839), .A2(n7588), .ZN(n6736) );
  NAND2_X1 U6853 ( .A1(n7583), .A2(n6736), .ZN(n7442) );
  NAND2_X1 U6854 ( .A1(n6937), .A2(n6635), .ZN(n5252) );
  NAND2_X1 U6855 ( .A1(n5248), .A2(n5265), .ZN(n5249) );
  NAND2_X1 U6856 ( .A1(n5249), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5250) );
  XNOR2_X1 U6857 ( .A(n5250), .B(P1_IR_REG_9__SCAN_IN), .ZN(n7005) );
  AOI22_X1 U6858 ( .A1(n5535), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n5406), .B2(
        n7005), .ZN(n5251) );
  NAND2_X1 U6859 ( .A1(n5252), .A2(n5251), .ZN(n9173) );
  NAND2_X1 U6860 ( .A1(n6639), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5261) );
  INV_X1 U6861 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n5253) );
  OR2_X1 U6862 ( .A1(n5649), .A2(n5253), .ZN(n5260) );
  INV_X1 U6863 ( .A(n5254), .ZN(n5273) );
  NAND2_X1 U6864 ( .A1(n5255), .A2(n10209), .ZN(n5256) );
  NAND2_X1 U6865 ( .A1(n5273), .A2(n5256), .ZN(n7596) );
  OR2_X1 U6866 ( .A1(n5572), .A2(n7596), .ZN(n5259) );
  INV_X1 U6867 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n7004) );
  OR2_X1 U6868 ( .A1(n4413), .A2(n7004), .ZN(n5258) );
  NAND4_X1 U6869 ( .A1(n5261), .A2(n5260), .A3(n5259), .A4(n5258), .ZN(n9257)
         );
  INV_X1 U6870 ( .A(n9257), .ZN(n7439) );
  NAND2_X1 U6871 ( .A1(n9173), .A2(n7439), .ZN(n6751) );
  NAND2_X1 U6872 ( .A1(n6739), .A2(n6751), .ZN(n7591) );
  NAND2_X1 U6873 ( .A1(n7590), .A2(n5262), .ZN(n7737) );
  NAND2_X1 U6874 ( .A1(n6942), .A2(n6635), .ZN(n5270) );
  NAND2_X1 U6875 ( .A1(n5265), .A2(n5264), .ZN(n5266) );
  NAND2_X1 U6876 ( .A1(n5282), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5268) );
  XNOR2_X1 U6877 ( .A(n5268), .B(P1_IR_REG_10__SCAN_IN), .ZN(n7068) );
  AOI22_X1 U6878 ( .A1(n5535), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n5406), .B2(
        n7068), .ZN(n5269) );
  NAND2_X1 U6879 ( .A1(n5270), .A2(n5269), .ZN(n7756) );
  NAND2_X1 U6880 ( .A1(n6639), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5278) );
  INV_X1 U6881 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n5271) );
  OR2_X1 U6882 ( .A1(n5649), .A2(n5271), .ZN(n5277) );
  INV_X1 U6883 ( .A(n5272), .ZN(n5288) );
  NAND2_X1 U6884 ( .A1(n5273), .A2(n10192), .ZN(n5274) );
  NAND2_X1 U6885 ( .A1(n5288), .A2(n5274), .ZN(n7914) );
  OR2_X1 U6886 ( .A1(n5446), .A2(n7914), .ZN(n5276) );
  INV_X1 U6887 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n7007) );
  OR2_X1 U6888 ( .A1(n4413), .A2(n7007), .ZN(n5275) );
  OR2_X1 U6889 ( .A1(n7756), .A2(n7830), .ZN(n6754) );
  NAND2_X1 U6890 ( .A1(n7756), .A2(n7830), .ZN(n7812) );
  NAND2_X1 U6891 ( .A1(n6754), .A2(n7812), .ZN(n7736) );
  NAND2_X1 U6892 ( .A1(n7737), .A2(n7736), .ZN(n7735) );
  INV_X1 U6893 ( .A(n7830), .ZN(n9256) );
  NAND2_X1 U6894 ( .A1(n7735), .A2(n5279), .ZN(n7818) );
  XNOR2_X1 U6895 ( .A(n5281), .B(n5280), .ZN(n6947) );
  NAND2_X1 U6896 ( .A1(n6947), .A2(n6635), .ZN(n5285) );
  OAI21_X1 U6897 ( .B1(n5282), .B2(P1_IR_REG_10__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5283) );
  XNOR2_X1 U6898 ( .A(n5283), .B(P1_IR_REG_11__SCAN_IN), .ZN(n7296) );
  AOI22_X1 U6899 ( .A1(n5535), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n5406), .B2(
        n7296), .ZN(n5284) );
  NAND2_X1 U6900 ( .A1(n6639), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5293) );
  INV_X1 U6901 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n5286) );
  OR2_X1 U6902 ( .A1(n5369), .A2(n5286), .ZN(n5292) );
  INV_X1 U6903 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n5287) );
  NAND2_X1 U6904 ( .A1(n5288), .A2(n5287), .ZN(n5289) );
  NAND2_X1 U6905 ( .A1(n5305), .A2(n5289), .ZN(n7819) );
  OR2_X1 U6906 ( .A1(n5572), .A2(n7819), .ZN(n5291) );
  INV_X1 U6907 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n7073) );
  OR2_X1 U6908 ( .A1(n4413), .A2(n7073), .ZN(n5290) );
  NAND4_X1 U6909 ( .A1(n5293), .A2(n5292), .A3(n5291), .A4(n5290), .ZN(n9255)
         );
  NAND2_X1 U6910 ( .A1(n9210), .A2(n7981), .ZN(n6743) );
  NAND2_X1 U6911 ( .A1(n6741), .A2(n6743), .ZN(n7817) );
  NAND2_X1 U6912 ( .A1(n7818), .A2(n7817), .ZN(n7816) );
  NAND2_X1 U6913 ( .A1(n7816), .A2(n5294), .ZN(n7854) );
  XNOR2_X1 U6914 ( .A(n5296), .B(n5295), .ZN(n6952) );
  NAND2_X1 U6915 ( .A1(n6952), .A2(n6635), .ZN(n5303) );
  OR2_X1 U6916 ( .A1(n5297), .A2(n9815), .ZN(n5300) );
  INV_X1 U6917 ( .A(n5300), .ZN(n5298) );
  NAND2_X1 U6918 ( .A1(n5298), .A2(P1_IR_REG_12__SCAN_IN), .ZN(n5301) );
  INV_X1 U6919 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n5299) );
  NAND2_X1 U6920 ( .A1(n5300), .A2(n5299), .ZN(n5316) );
  AOI22_X1 U6921 ( .A1(n5535), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n5406), .B2(
        n7293), .ZN(n5302) );
  NAND2_X1 U6922 ( .A1(n5257), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n5312) );
  INV_X1 U6923 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n7290) );
  OR2_X1 U6924 ( .A1(n5369), .A2(n7290), .ZN(n5311) );
  NAND2_X1 U6925 ( .A1(n5305), .A2(n5304), .ZN(n5306) );
  NAND2_X1 U6926 ( .A1(n5321), .A2(n5306), .ZN(n7861) );
  OR2_X1 U6927 ( .A1(n5572), .A2(n7861), .ZN(n5310) );
  INV_X1 U6928 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n5307) );
  OR2_X1 U6929 ( .A1(n5308), .A2(n5307), .ZN(n5309) );
  NAND4_X1 U6930 ( .A1(n5312), .A2(n5311), .A3(n5310), .A4(n5309), .ZN(n9254)
         );
  INV_X1 U6931 ( .A(n9254), .ZN(n7962) );
  OR2_X1 U6932 ( .A1(n7889), .A2(n7962), .ZN(n7956) );
  NAND2_X1 U6933 ( .A1(n7889), .A2(n7962), .ZN(n6756) );
  NAND2_X1 U6934 ( .A1(n7956), .A2(n6756), .ZN(n7853) );
  NAND2_X1 U6935 ( .A1(n7854), .A2(n7853), .ZN(n7852) );
  NAND2_X1 U6936 ( .A1(n7852), .A2(n5313), .ZN(n7954) );
  XNOR2_X1 U6937 ( .A(n5315), .B(n5314), .ZN(n6956) );
  NAND2_X1 U6938 ( .A1(n6956), .A2(n6635), .ZN(n5319) );
  NAND2_X1 U6939 ( .A1(n5316), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5317) );
  XNOR2_X1 U6940 ( .A(n5317), .B(P1_IR_REG_13__SCAN_IN), .ZN(n7474) );
  AOI22_X1 U6941 ( .A1(n5535), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n5406), .B2(
        n7474), .ZN(n5318) );
  NAND2_X1 U6942 ( .A1(n6639), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n5326) );
  INV_X1 U6943 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n5320) );
  OR2_X1 U6944 ( .A1(n5369), .A2(n5320), .ZN(n5325) );
  NAND2_X1 U6945 ( .A1(n5321), .A2(n10341), .ZN(n5322) );
  NAND2_X1 U6946 ( .A1(n5340), .A2(n5322), .ZN(n7964) );
  OR2_X1 U6947 ( .A1(n5446), .A2(n7964), .ZN(n5324) );
  INV_X1 U6948 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n7479) );
  OR2_X1 U6949 ( .A1(n4413), .A2(n7479), .ZN(n5323) );
  OR2_X1 U6950 ( .A1(n9744), .A2(n8114), .ZN(n6759) );
  NAND2_X1 U6951 ( .A1(n9744), .A2(n8114), .ZN(n8100) );
  NAND2_X1 U6952 ( .A1(n6759), .A2(n8100), .ZN(n7960) );
  NAND2_X1 U6953 ( .A1(n7954), .A2(n7960), .ZN(n7953) );
  XNOR2_X1 U6954 ( .A(n5328), .B(n5329), .ZN(n7014) );
  NAND2_X1 U6955 ( .A1(n7014), .A2(n6635), .ZN(n5337) );
  NOR2_X1 U6956 ( .A1(n5330), .A2(n9815), .ZN(n5331) );
  MUX2_X1 U6957 ( .A(n9815), .B(n5331), .S(P1_IR_REG_14__SCAN_IN), .Z(n5332)
         );
  INV_X1 U6958 ( .A(n5332), .ZN(n5335) );
  INV_X1 U6959 ( .A(n5333), .ZN(n5334) );
  AOI22_X1 U6960 ( .A1(n5535), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n5406), .B2(
        n9324), .ZN(n5336) );
  NAND2_X1 U6961 ( .A1(n6639), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5345) );
  INV_X1 U6962 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n8107) );
  OR2_X1 U6963 ( .A1(n5649), .A2(n8107), .ZN(n5344) );
  INV_X1 U6964 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n9332) );
  OR2_X1 U6965 ( .A1(n4413), .A2(n9332), .ZN(n5343) );
  INV_X1 U6966 ( .A(n5338), .ZN(n5354) );
  NAND2_X1 U6967 ( .A1(n5340), .A2(n5339), .ZN(n5341) );
  NAND2_X1 U6968 ( .A1(n5354), .A2(n5341), .ZN(n9057) );
  OR2_X1 U6969 ( .A1(n5572), .A2(n9057), .ZN(n5342) );
  NAND4_X1 U6970 ( .A1(n5345), .A2(n5344), .A3(n5343), .A4(n5342), .ZN(n9252)
         );
  NAND2_X1 U6971 ( .A1(n9059), .A2(n9252), .ZN(n5347) );
  XNOR2_X1 U6972 ( .A(n5349), .B(SI_15_), .ZN(n5350) );
  XNOR2_X1 U6973 ( .A(n5348), .B(n5350), .ZN(n7019) );
  NAND2_X1 U6974 ( .A1(n7019), .A2(n6635), .ZN(n5353) );
  OR2_X1 U6975 ( .A1(n5333), .A2(n9815), .ZN(n5351) );
  XNOR2_X1 U6976 ( .A(n5351), .B(P1_IR_REG_15__SCAN_IN), .ZN(n9338) );
  AOI22_X1 U6977 ( .A1(n5535), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n5406), .B2(
        n9338), .ZN(n5352) );
  NAND2_X1 U6978 ( .A1(n5146), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n5360) );
  INV_X1 U6979 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n10076) );
  OR2_X1 U6980 ( .A1(n5308), .A2(n10076), .ZN(n5359) );
  INV_X1 U6981 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n10340) );
  NAND2_X1 U6982 ( .A1(n5354), .A2(n10340), .ZN(n5355) );
  NAND2_X1 U6983 ( .A1(n5367), .A2(n5355), .ZN(n9238) );
  OR2_X1 U6984 ( .A1(n5446), .A2(n9238), .ZN(n5358) );
  INV_X1 U6985 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n5356) );
  OR2_X1 U6986 ( .A1(n4413), .A2(n5356), .ZN(n5357) );
  NAND4_X1 U6987 ( .A1(n5360), .A2(n5359), .A3(n5358), .A4(n5357), .ZN(n9624)
         );
  INV_X1 U6988 ( .A(n9739), .ZN(n9248) );
  INV_X1 U6989 ( .A(n9624), .ZN(n9134) );
  XNOR2_X1 U6990 ( .A(n5361), .B(SI_16_), .ZN(n5362) );
  XNOR2_X1 U6991 ( .A(n5363), .B(n5362), .ZN(n7163) );
  NAND2_X1 U6992 ( .A1(n7163), .A2(n6635), .ZN(n5366) );
  NAND2_X1 U6993 ( .A1(n5378), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5364) );
  XNOR2_X1 U6994 ( .A(n5364), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9365) );
  AOI22_X1 U6995 ( .A1(n5535), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n5406), .B2(
        n9365), .ZN(n5365) );
  NAND2_X1 U6996 ( .A1(n5367), .A2(n9131), .ZN(n5368) );
  AND2_X1 U6997 ( .A1(n9143), .A2(n5368), .ZN(n9631) );
  INV_X1 U6998 ( .A(n5572), .ZN(n5384) );
  NAND2_X1 U6999 ( .A1(n9631), .A2(n5384), .ZN(n5373) );
  NAND2_X1 U7000 ( .A1(n6639), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n5372) );
  INV_X1 U7001 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n10147) );
  OR2_X1 U7002 ( .A1(n5369), .A2(n10147), .ZN(n5371) );
  INV_X1 U7003 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9357) );
  OR2_X1 U7004 ( .A1(n4413), .A2(n9357), .ZN(n5370) );
  NAND4_X1 U7005 ( .A1(n5373), .A2(n5372), .A3(n5371), .A4(n5370), .ZN(n9722)
         );
  NAND2_X1 U7006 ( .A1(n9801), .A2(n9607), .ZN(n6770) );
  NAND2_X1 U7007 ( .A1(n6767), .A2(n6770), .ZN(n9618) );
  XNOR2_X1 U7008 ( .A(n5376), .B(n5375), .ZN(n7250) );
  NAND2_X1 U7009 ( .A1(n7250), .A2(n6635), .ZN(n5381) );
  NAND2_X1 U7010 ( .A1(n4507), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5379) );
  XNOR2_X1 U7011 ( .A(n5379), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9859) );
  AOI22_X1 U7012 ( .A1(n5535), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n5406), .B2(
        n9859), .ZN(n5380) );
  NAND2_X1 U7013 ( .A1(n6639), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n5383) );
  NAND2_X1 U7014 ( .A1(n5146), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n5382) );
  AND2_X1 U7015 ( .A1(n5383), .A2(n5382), .ZN(n5387) );
  XNOR2_X1 U7016 ( .A(n9143), .B(P1_REG3_REG_17__SCAN_IN), .ZN(n9603) );
  NAND2_X1 U7017 ( .A1(n9603), .A2(n5384), .ZN(n5386) );
  INV_X1 U7018 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9728) );
  OR2_X1 U7019 ( .A1(n4413), .A2(n9728), .ZN(n5385) );
  NAND2_X1 U7020 ( .A1(n9724), .A2(n9625), .ZN(n5389) );
  INV_X1 U7021 ( .A(n9724), .ZN(n9600) );
  XNOR2_X1 U7022 ( .A(n5391), .B(n5390), .ZN(n7275) );
  NAND2_X1 U7023 ( .A1(n7275), .A2(n6635), .ZN(n5396) );
  NAND2_X1 U7024 ( .A1(n5591), .A2(n5393), .ZN(n5404) );
  OR2_X1 U7025 ( .A1(n5591), .A2(n5393), .ZN(n5394) );
  AND2_X1 U7026 ( .A1(n5404), .A2(n5394), .ZN(n9381) );
  AOI22_X1 U7027 ( .A1(n5535), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n5406), .B2(
        n9381), .ZN(n5395) );
  OR2_X1 U7028 ( .A1(n5397), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n5398) );
  NAND2_X1 U7029 ( .A1(n5398), .A2(n5409), .ZN(n9582) );
  AOI22_X1 U7030 ( .A1(n5146), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n6639), .B2(
        P1_REG0_REG_18__SCAN_IN), .ZN(n5400) );
  NAND2_X1 U7031 ( .A1(n5257), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n5399) );
  OAI211_X1 U7032 ( .C1(n9582), .C2(n5572), .A(n5400), .B(n5399), .ZN(n9610)
         );
  NAND2_X1 U7033 ( .A1(n9580), .A2(n4998), .ZN(n5401) );
  INV_X1 U7034 ( .A(n9610), .ZN(n10056) );
  XNOR2_X1 U7035 ( .A(n5403), .B(n5402), .ZN(n7544) );
  NAND2_X1 U7036 ( .A1(n7544), .A2(n6635), .ZN(n5408) );
  AOI22_X1 U7037 ( .A1(n5535), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n5666), .B2(
        n5406), .ZN(n5407) );
  NAND2_X1 U7038 ( .A1(n6639), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n5416) );
  INV_X1 U7039 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n9379) );
  OR2_X1 U7040 ( .A1(n5649), .A2(n9379), .ZN(n5415) );
  INV_X1 U7041 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n10297) );
  OR2_X1 U7042 ( .A1(n4413), .A2(n10297), .ZN(n5414) );
  INV_X1 U7043 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n5410) );
  NAND2_X1 U7044 ( .A1(n5410), .A2(n5409), .ZN(n5411) );
  NAND2_X1 U7045 ( .A1(n5412), .A2(n5411), .ZN(n9568) );
  OR2_X1 U7046 ( .A1(n5572), .A2(n9568), .ZN(n5413) );
  INV_X1 U7047 ( .A(n9706), .ZN(n9554) );
  INV_X1 U7048 ( .A(n9714), .ZN(n9571) );
  OAI21_X1 U7049 ( .B1(n9524), .B2(n9558), .A(n5417), .ZN(n9522) );
  INV_X1 U7050 ( .A(n5418), .ZN(n5419) );
  MUX2_X1 U7051 ( .A(n7694), .B(n7734), .S(n6915), .Z(n5435) );
  XNOR2_X1 U7052 ( .A(n5435), .B(SI_21_), .ZN(n5422) );
  XNOR2_X1 U7053 ( .A(n5438), .B(n5422), .ZN(n7693) );
  NAND2_X1 U7054 ( .A1(n7693), .A2(n6635), .ZN(n5424) );
  NAND2_X1 U7055 ( .A1(n5535), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n5423) );
  NAND2_X1 U7056 ( .A1(n6639), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n5433) );
  INV_X1 U7057 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n9523) );
  OR2_X1 U7058 ( .A1(n5649), .A2(n9523), .ZN(n5432) );
  INV_X1 U7059 ( .A(n5445), .ZN(n5429) );
  INV_X1 U7060 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n5426) );
  NAND2_X1 U7061 ( .A1(n5427), .A2(n5426), .ZN(n5428) );
  NAND2_X1 U7062 ( .A1(n5429), .A2(n5428), .ZN(n9537) );
  OR2_X1 U7063 ( .A1(n5572), .A2(n9537), .ZN(n5431) );
  INV_X1 U7064 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n9701) );
  OR2_X1 U7065 ( .A1(n4413), .A2(n9701), .ZN(n5430) );
  NAND4_X1 U7066 ( .A1(n5433), .A2(n5432), .A3(n5431), .A4(n5430), .ZN(n9545)
         );
  NOR2_X1 U7067 ( .A1(n9536), .A2(n9688), .ZN(n5434) );
  NOR2_X1 U7068 ( .A1(n5436), .A2(SI_21_), .ZN(n5437) );
  MUX2_X1 U7069 ( .A(n10344), .B(n7851), .S(n6915), .Z(n5440) );
  INV_X1 U7070 ( .A(SI_22_), .ZN(n5439) );
  NAND2_X1 U7071 ( .A1(n5440), .A2(n5439), .ZN(n5451) );
  INV_X1 U7072 ( .A(n5440), .ZN(n5441) );
  NAND2_X1 U7073 ( .A1(n5441), .A2(SI_22_), .ZN(n5442) );
  NAND2_X1 U7074 ( .A1(n5451), .A2(n5442), .ZN(n5452) );
  XNOR2_X1 U7075 ( .A(n5453), .B(n5452), .ZN(n7847) );
  NAND2_X1 U7076 ( .A1(n7847), .A2(n6635), .ZN(n5444) );
  NAND2_X1 U7077 ( .A1(n5535), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n5443) );
  NAND2_X1 U7078 ( .A1(n5257), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n5450) );
  INV_X1 U7079 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n10334) );
  OR2_X1 U7080 ( .A1(n5649), .A2(n10334), .ZN(n5449) );
  OAI21_X1 U7081 ( .B1(n5445), .B2(P1_REG3_REG_22__SCAN_IN), .A(n5462), .ZN(
        n9510) );
  OR2_X1 U7082 ( .A1(n5446), .A2(n9510), .ZN(n5448) );
  INV_X1 U7083 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n9777) );
  OR2_X1 U7084 ( .A1(n5308), .A2(n9777), .ZN(n5447) );
  NAND4_X1 U7085 ( .A1(n5450), .A2(n5449), .A3(n5448), .A4(n5447), .ZN(n9532)
         );
  NAND2_X1 U7086 ( .A1(n9509), .A2(n9499), .ZN(n6665) );
  NAND2_X1 U7087 ( .A1(n6659), .A2(n6665), .ZN(n5636) );
  INV_X1 U7088 ( .A(n9509), .ZN(n9689) );
  OAI21_X1 U7089 ( .B1(n5453), .B2(n5452), .A(n5451), .ZN(n5470) );
  INV_X1 U7090 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n5454) );
  MUX2_X1 U7091 ( .A(n7946), .B(n5454), .S(n6915), .Z(n5456) );
  INV_X1 U7092 ( .A(SI_23_), .ZN(n5455) );
  NAND2_X1 U7093 ( .A1(n5456), .A2(n5455), .ZN(n5471) );
  INV_X1 U7094 ( .A(n5456), .ZN(n5457) );
  NAND2_X1 U7095 ( .A1(n5457), .A2(SI_23_), .ZN(n5458) );
  XNOR2_X1 U7096 ( .A(n5470), .B(n5469), .ZN(n7943) );
  NAND2_X1 U7097 ( .A1(n7943), .A2(n6635), .ZN(n5460) );
  NAND2_X1 U7098 ( .A1(n5535), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n5459) );
  NAND2_X1 U7099 ( .A1(n6639), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n5467) );
  INV_X1 U7100 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n5461) );
  OR2_X1 U7101 ( .A1(n5649), .A2(n5461), .ZN(n5466) );
  XNOR2_X1 U7102 ( .A(P1_REG3_REG_23__SCAN_IN), .B(n5479), .ZN(n9503) );
  OR2_X1 U7103 ( .A1(n5572), .A2(n9503), .ZN(n5465) );
  INV_X1 U7104 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n5463) );
  OR2_X1 U7105 ( .A1(n4413), .A2(n5463), .ZN(n5464) );
  NAND4_X1 U7106 ( .A1(n5467), .A2(n5466), .A3(n5465), .A4(n5464), .ZN(n9675)
         );
  NAND2_X1 U7107 ( .A1(n5655), .A2(n9519), .ZN(n5468) );
  AOI22_X1 U7108 ( .A1(n9493), .A2(n5468), .B1(n9685), .B2(n9675), .ZN(n9474)
         );
  NAND2_X1 U7109 ( .A1(n5470), .A2(n5469), .ZN(n5472) );
  NAND2_X1 U7110 ( .A1(n5472), .A2(n5471), .ZN(n5488) );
  MUX2_X1 U7111 ( .A(n10235), .B(n10271), .S(n6915), .Z(n5474) );
  INV_X1 U7112 ( .A(SI_24_), .ZN(n5473) );
  NAND2_X1 U7113 ( .A1(n5474), .A2(n5473), .ZN(n5489) );
  INV_X1 U7114 ( .A(n5474), .ZN(n5475) );
  NAND2_X1 U7115 ( .A1(n5475), .A2(SI_24_), .ZN(n5476) );
  XNOR2_X1 U7116 ( .A(n5488), .B(n5487), .ZN(n8005) );
  NAND2_X1 U7117 ( .A1(n8005), .A2(n6635), .ZN(n5478) );
  OR2_X1 U7118 ( .A1(n5155), .A2(n10271), .ZN(n5477) );
  NAND2_X1 U7119 ( .A1(n6639), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n5485) );
  INV_X1 U7120 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n9485) );
  OR2_X1 U7121 ( .A1(n5649), .A2(n9485), .ZN(n5484) );
  NAND3_X1 U7122 ( .A1(P1_REG3_REG_23__SCAN_IN), .A2(P1_REG3_REG_24__SCAN_IN), 
        .A3(n5479), .ZN(n5498) );
  INV_X1 U7123 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n10098) );
  NAND2_X1 U7124 ( .A1(P1_REG3_REG_23__SCAN_IN), .A2(n5479), .ZN(n5480) );
  NAND2_X1 U7125 ( .A1(n10098), .A2(n5480), .ZN(n5481) );
  NAND2_X1 U7126 ( .A1(n5498), .A2(n5481), .ZN(n9484) );
  OR2_X1 U7127 ( .A1(n5572), .A2(n9484), .ZN(n5483) );
  INV_X1 U7128 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n9681) );
  OR2_X1 U7129 ( .A1(n4413), .A2(n9681), .ZN(n5482) );
  NAND4_X1 U7130 ( .A1(n5485), .A2(n5484), .A3(n5483), .A4(n5482), .ZN(n9469)
         );
  NAND2_X1 U7131 ( .A1(n9676), .A2(n9469), .ZN(n5486) );
  AOI22_X1 U7132 ( .A1(n9474), .A2(n5486), .B1(n4683), .B2(n9668), .ZN(n9458)
         );
  NAND2_X1 U7133 ( .A1(n5488), .A2(n5487), .ZN(n5490) );
  INV_X1 U7134 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n8133) );
  INV_X1 U7135 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n8081) );
  MUX2_X1 U7136 ( .A(n8133), .B(n8081), .S(n6915), .Z(n5492) );
  INV_X1 U7137 ( .A(SI_25_), .ZN(n5491) );
  NAND2_X1 U7138 ( .A1(n5492), .A2(n5491), .ZN(n5508) );
  INV_X1 U7139 ( .A(n5492), .ZN(n5493) );
  NAND2_X1 U7140 ( .A1(n5493), .A2(SI_25_), .ZN(n5494) );
  XNOR2_X1 U7141 ( .A(n5507), .B(n5506), .ZN(n8080) );
  NAND2_X1 U7142 ( .A1(n8080), .A2(n6635), .ZN(n5496) );
  NAND2_X1 U7143 ( .A1(n5535), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n5495) );
  NAND2_X1 U7144 ( .A1(n6639), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n5503) );
  INV_X1 U7145 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n9467) );
  OR2_X1 U7146 ( .A1(n5649), .A2(n9467), .ZN(n5502) );
  INV_X1 U7147 ( .A(n5498), .ZN(n5497) );
  NAND2_X1 U7148 ( .A1(n5497), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n5518) );
  INV_X1 U7149 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n10058) );
  NAND2_X1 U7150 ( .A1(n5498), .A2(n10058), .ZN(n5499) );
  NAND2_X1 U7151 ( .A1(n5518), .A2(n5499), .ZN(n9466) );
  OR2_X1 U7152 ( .A1(n5572), .A2(n9466), .ZN(n5501) );
  INV_X1 U7153 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n9673) );
  OR2_X1 U7154 ( .A1(n4413), .A2(n9673), .ZN(n5500) );
  NAND2_X1 U7155 ( .A1(n9669), .A2(n9478), .ZN(n5505) );
  NOR2_X1 U7156 ( .A1(n9669), .A2(n9478), .ZN(n5504) );
  AOI21_X1 U7157 ( .B1(n9458), .B2(n5505), .A(n5504), .ZN(n9445) );
  NAND2_X1 U7158 ( .A1(n5507), .A2(n5506), .ZN(n5509) );
  NAND2_X1 U7159 ( .A1(n5509), .A2(n5508), .ZN(n5528) );
  INV_X1 U7160 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n10143) );
  INV_X1 U7161 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n8126) );
  MUX2_X1 U7162 ( .A(n10143), .B(n8126), .S(n6915), .Z(n5511) );
  INV_X1 U7163 ( .A(SI_26_), .ZN(n5510) );
  NAND2_X1 U7164 ( .A1(n5511), .A2(n5510), .ZN(n5529) );
  INV_X1 U7165 ( .A(n5511), .ZN(n5512) );
  NAND2_X1 U7166 ( .A1(n5512), .A2(SI_26_), .ZN(n5513) );
  NAND2_X1 U7167 ( .A1(n8125), .A2(n6635), .ZN(n5515) );
  NAND2_X1 U7168 ( .A1(n5535), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n5514) );
  NAND2_X1 U7169 ( .A1(n6639), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n5523) );
  INV_X1 U7170 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n9449) );
  OR2_X1 U7171 ( .A1(n5649), .A2(n9449), .ZN(n5522) );
  INV_X1 U7172 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n10284) );
  OR2_X1 U7173 ( .A1(n4413), .A2(n10284), .ZN(n5521) );
  INV_X1 U7174 ( .A(n5518), .ZN(n5516) );
  NAND2_X1 U7175 ( .A1(n5516), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n5539) );
  INV_X1 U7176 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n5517) );
  NAND2_X1 U7177 ( .A1(n5518), .A2(n5517), .ZN(n5519) );
  NAND2_X1 U7178 ( .A1(n5539), .A2(n5519), .ZN(n9448) );
  OR2_X1 U7179 ( .A1(n5572), .A2(n9448), .ZN(n5520) );
  INV_X1 U7180 ( .A(n9657), .ZN(n5524) );
  NAND2_X1 U7181 ( .A1(n9452), .A2(n9657), .ZN(n5526) );
  NAND2_X1 U7182 ( .A1(n5528), .A2(n5527), .ZN(n5530) );
  INV_X1 U7183 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n8197) );
  INV_X1 U7184 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n8196) );
  MUX2_X1 U7185 ( .A(n8197), .B(n8196), .S(n6915), .Z(n5532) );
  INV_X1 U7186 ( .A(SI_27_), .ZN(n5531) );
  NAND2_X1 U7187 ( .A1(n5532), .A2(n5531), .ZN(n5547) );
  INV_X1 U7188 ( .A(n5532), .ZN(n5533) );
  NAND2_X1 U7189 ( .A1(n5533), .A2(SI_27_), .ZN(n5534) );
  NAND2_X1 U7190 ( .A1(n8194), .A2(n6635), .ZN(n5537) );
  NAND2_X1 U7191 ( .A1(n5535), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n5536) );
  NAND2_X1 U7192 ( .A1(n5146), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n5544) );
  INV_X1 U7193 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n9759) );
  OR2_X1 U7194 ( .A1(n5308), .A2(n9759), .ZN(n5543) );
  INV_X1 U7195 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n5538) );
  NAND2_X1 U7196 ( .A1(n5539), .A2(n5538), .ZN(n5540) );
  NAND2_X1 U7197 ( .A1(n5556), .A2(n5540), .ZN(n6604) );
  OR2_X1 U7198 ( .A1(n5572), .A2(n6604), .ZN(n5542) );
  INV_X1 U7199 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n9662) );
  OR2_X1 U7200 ( .A1(n4413), .A2(n9662), .ZN(n5541) );
  NAND4_X1 U7201 ( .A1(n5544), .A2(n5543), .A3(n5542), .A4(n5541), .ZN(n9648)
         );
  NAND2_X1 U7202 ( .A1(n9424), .A2(n9441), .ZN(n9405) );
  NAND2_X1 U7203 ( .A1(n5546), .A2(n5545), .ZN(n5548) );
  INV_X1 U7204 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n8132) );
  MUX2_X1 U7205 ( .A(n10301), .B(n8132), .S(n6915), .Z(n5550) );
  INV_X1 U7206 ( .A(SI_28_), .ZN(n5549) );
  NAND2_X1 U7207 ( .A1(n5550), .A2(n5549), .ZN(n5566) );
  INV_X1 U7208 ( .A(n5550), .ZN(n5551) );
  NAND2_X1 U7209 ( .A1(n5551), .A2(SI_28_), .ZN(n5552) );
  XNOR2_X1 U7210 ( .A(n5565), .B(n5564), .ZN(n6080) );
  NAND2_X1 U7211 ( .A1(n6080), .A2(n6635), .ZN(n5554) );
  OR2_X1 U7212 ( .A1(n5155), .A2(n8132), .ZN(n5553) );
  NAND2_X1 U7213 ( .A1(n5146), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n5562) );
  INV_X1 U7214 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n10281) );
  OR2_X1 U7215 ( .A1(n5308), .A2(n10281), .ZN(n5561) );
  INV_X1 U7216 ( .A(n5556), .ZN(n5555) );
  NAND2_X1 U7217 ( .A1(n5555), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n5671) );
  INV_X1 U7218 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n10280) );
  NAND2_X1 U7219 ( .A1(n5556), .A2(n10280), .ZN(n5557) );
  NAND2_X1 U7220 ( .A1(n5671), .A2(n5557), .ZN(n9413) );
  OR2_X1 U7221 ( .A1(n5572), .A2(n9413), .ZN(n5560) );
  INV_X1 U7222 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n5558) );
  OR2_X1 U7223 ( .A1(n4413), .A2(n5558), .ZN(n5559) );
  NAND2_X1 U7224 ( .A1(n9649), .A2(n9432), .ZN(n6673) );
  NAND2_X1 U7225 ( .A1(n9412), .A2(n9411), .ZN(n9646) );
  INV_X1 U7226 ( .A(n9432), .ZN(n9250) );
  NAND2_X1 U7227 ( .A1(n9649), .A2(n9250), .ZN(n5563) );
  NAND2_X1 U7228 ( .A1(n9646), .A2(n5563), .ZN(n5577) );
  NAND2_X1 U7229 ( .A1(n5565), .A2(n5564), .ZN(n5567) );
  MUX2_X1 U7230 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .S(n6915), .Z(n6621) );
  INV_X1 U7231 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n9823) );
  OR2_X1 U7232 ( .A1(n5155), .A2(n9823), .ZN(n5570) );
  NAND2_X1 U7233 ( .A1(n6639), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n5576) );
  INV_X1 U7234 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n5672) );
  OR2_X1 U7235 ( .A1(n5649), .A2(n5672), .ZN(n5575) );
  INV_X1 U7236 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n5686) );
  OR2_X1 U7237 ( .A1(n4413), .A2(n5686), .ZN(n5574) );
  OR2_X1 U7238 ( .A1(n5572), .A2(n5671), .ZN(n5573) );
  NAND4_X1 U7239 ( .A1(n5576), .A2(n5575), .A3(n5574), .A4(n5573), .ZN(n9410)
         );
  XNOR2_X1 U7240 ( .A(n6821), .B(n9410), .ZN(n6824) );
  NAND2_X1 U7241 ( .A1(n5610), .A2(n5612), .ZN(n5582) );
  NAND2_X1 U7242 ( .A1(n8082), .A2(P1_B_REG_SCAN_IN), .ZN(n5585) );
  MUX2_X1 U7243 ( .A(P1_B_REG_SCAN_IN), .B(n5585), .S(n5607), .Z(n5588) );
  INV_X1 U7244 ( .A(n8128), .ZN(n5587) );
  OR2_X1 U7245 ( .A1(n9809), .A2(P1_D_REG_1__SCAN_IN), .ZN(n5589) );
  NAND2_X1 U7246 ( .A1(n8082), .A2(n8128), .ZN(n9810) );
  OAI21_X1 U7247 ( .B1(P1_IR_REG_18__SCAN_IN), .B2(P1_IR_REG_19__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5590) );
  NAND2_X1 U7248 ( .A1(n5591), .A2(n5590), .ZN(n5595) );
  INV_X1 U7249 ( .A(n5595), .ZN(n5592) );
  NAND2_X1 U7250 ( .A1(n4486), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5594) );
  NAND2_X1 U7251 ( .A1(n5595), .A2(P1_IR_REG_20__SCAN_IN), .ZN(n5596) );
  INV_X1 U7252 ( .A(n6605), .ZN(n5598) );
  NOR2_X1 U7253 ( .A1(n6599), .A2(n5598), .ZN(n5615) );
  NOR2_X1 U7254 ( .A1(P1_D_REG_12__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .ZN(
        n10322) );
  NOR2_X1 U7255 ( .A1(P1_D_REG_31__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .ZN(
        n10319) );
  NOR4_X1 U7256 ( .A1(P1_D_REG_30__SCAN_IN), .A2(P1_D_REG_20__SCAN_IN), .A3(
        P1_D_REG_2__SCAN_IN), .A4(P1_D_REG_29__SCAN_IN), .ZN(n5605) );
  INV_X1 U7257 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n10064) );
  INV_X1 U7258 ( .A(P1_D_REG_26__SCAN_IN), .ZN(n10159) );
  INV_X1 U7259 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n10238) );
  INV_X1 U7260 ( .A(P1_D_REG_18__SCAN_IN), .ZN(n10237) );
  NAND4_X1 U7261 ( .A1(n10064), .A2(n10159), .A3(n10238), .A4(n10237), .ZN(
        n10296) );
  NOR4_X1 U7262 ( .A1(P1_D_REG_11__SCAN_IN), .A2(P1_D_REG_9__SCAN_IN), .A3(
        P1_D_REG_10__SCAN_IN), .A4(P1_D_REG_28__SCAN_IN), .ZN(n5602) );
  NOR4_X1 U7263 ( .A1(P1_D_REG_8__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_5__SCAN_IN), .A4(P1_D_REG_6__SCAN_IN), .ZN(n5601) );
  NOR4_X1 U7264 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_16__SCAN_IN), .A3(
        P1_D_REG_17__SCAN_IN), .A4(P1_D_REG_22__SCAN_IN), .ZN(n5600) );
  NOR4_X1 U7265 ( .A1(P1_D_REG_27__SCAN_IN), .A2(P1_D_REG_24__SCAN_IN), .A3(
        P1_D_REG_25__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n5599) );
  NAND4_X1 U7266 ( .A1(n5602), .A2(n5601), .A3(n5600), .A4(n5599), .ZN(n5603)
         );
  NOR4_X1 U7267 ( .A1(P1_D_REG_21__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        n10296), .A4(n5603), .ZN(n5604) );
  AND4_X1 U7268 ( .A1(n10322), .A2(n10319), .A3(n5605), .A4(n5604), .ZN(n5606)
         );
  NAND2_X1 U7269 ( .A1(n5617), .A2(n7667), .ZN(n6842) );
  INV_X1 U7270 ( .A(n6842), .ZN(n6680) );
  OR2_X1 U7271 ( .A1(n9876), .A2(n6680), .ZN(n5609) );
  NAND2_X1 U7272 ( .A1(n6408), .A2(n5609), .ZN(n6607) );
  INV_X1 U7273 ( .A(n5610), .ZN(n5611) );
  NAND2_X1 U7274 ( .A1(n5611), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5613) );
  NOR2_X1 U7275 ( .A1(n6607), .A2(n6871), .ZN(n5614) );
  NAND2_X1 U7276 ( .A1(n5607), .A2(n8128), .ZN(n9811) );
  NAND2_X1 U7277 ( .A1(n5617), .A2(n6843), .ZN(n6406) );
  NAND2_X1 U7278 ( .A1(n6842), .A2(n6406), .ZN(n5618) );
  AND2_X1 U7279 ( .A1(n9877), .A2(n5618), .ZN(n5619) );
  NAND2_X1 U7280 ( .A1(n5619), .A2(n9876), .ZN(n5668) );
  NAND2_X1 U7281 ( .A1(n6837), .A2(n7667), .ZN(n5620) );
  NAND2_X1 U7282 ( .A1(n5684), .A2(n9786), .ZN(n5661) );
  INV_X1 U7283 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n5656) );
  INV_X1 U7284 ( .A(n6824), .ZN(n5640) );
  INV_X1 U7285 ( .A(n9405), .ZN(n5621) );
  NOR2_X1 U7286 ( .A1(n9411), .A2(n5621), .ZN(n5638) );
  OR2_X1 U7287 ( .A1(n9764), .A2(n9657), .ZN(n6811) );
  NAND2_X1 U7288 ( .A1(n9764), .A2(n9657), .ZN(n6669) );
  NAND2_X1 U7289 ( .A1(n6811), .A2(n6669), .ZN(n9444) );
  INV_X1 U7290 ( .A(n9437), .ZN(n5622) );
  NOR2_X1 U7291 ( .A1(n9444), .A2(n5622), .ZN(n5637) );
  OR2_X1 U7292 ( .A1(n9059), .A2(n9240), .ZN(n6761) );
  NAND2_X1 U7293 ( .A1(n9059), .A2(n9240), .ZN(n6653) );
  NAND2_X1 U7294 ( .A1(n6761), .A2(n6653), .ZN(n8102) );
  INV_X1 U7295 ( .A(n8100), .ZN(n6745) );
  NOR2_X1 U7296 ( .A1(n8102), .A2(n6745), .ZN(n6764) );
  AND2_X1 U7297 ( .A1(n6419), .A2(n9879), .ZN(n7151) );
  NAND2_X1 U7298 ( .A1(n7152), .A2(n7151), .ZN(n5625) );
  NAND2_X1 U7299 ( .A1(n7087), .A2(n4417), .ZN(n5624) );
  NAND2_X1 U7300 ( .A1(n5625), .A2(n5624), .ZN(n7084) );
  INV_X1 U7301 ( .A(n5626), .ZN(n6709) );
  OR2_X1 U7302 ( .A1(n7084), .A2(n6709), .ZN(n6712) );
  INV_X1 U7303 ( .A(n7180), .ZN(n7184) );
  NAND2_X1 U7304 ( .A1(n7183), .A2(n7184), .ZN(n7182) );
  AND2_X1 U7305 ( .A1(n7182), .A2(n6713), .ZN(n7225) );
  NAND2_X1 U7306 ( .A1(n7225), .A2(n6714), .ZN(n7223) );
  NAND2_X1 U7307 ( .A1(n7223), .A2(n6722), .ZN(n7497) );
  INV_X1 U7308 ( .A(n7488), .ZN(n7498) );
  NAND2_X1 U7309 ( .A1(n7497), .A2(n7498), .ZN(n7496) );
  NAND2_X1 U7310 ( .A1(n7496), .A2(n6719), .ZN(n7329) );
  AND2_X1 U7311 ( .A1(n6736), .A2(n7437), .ZN(n7585) );
  INV_X1 U7312 ( .A(n7418), .ZN(n5628) );
  NOR2_X1 U7313 ( .A1(n5629), .A2(n5628), .ZN(n6694) );
  NAND2_X1 U7314 ( .A1(n7329), .A2(n6694), .ZN(n7739) );
  INV_X1 U7315 ( .A(n7736), .ZN(n7741) );
  AND2_X1 U7316 ( .A1(n7738), .A2(n7741), .ZN(n5630) );
  NAND2_X1 U7317 ( .A1(n7739), .A2(n5630), .ZN(n7740) );
  INV_X1 U7318 ( .A(n7812), .ZN(n5631) );
  NOR2_X1 U7319 ( .A1(n7817), .A2(n5631), .ZN(n5632) );
  NAND2_X1 U7320 ( .A1(n7740), .A2(n5632), .ZN(n5633) );
  NAND2_X1 U7321 ( .A1(n5633), .A2(n6741), .ZN(n7855) );
  INV_X1 U7322 ( .A(n7853), .ZN(n7856) );
  INV_X1 U7323 ( .A(n7956), .ZN(n5634) );
  NOR2_X1 U7324 ( .A1(n7960), .A2(n5634), .ZN(n5635) );
  OR2_X1 U7325 ( .A1(n9739), .A2(n9134), .ZN(n6762) );
  NAND2_X1 U7326 ( .A1(n9739), .A2(n9134), .ZN(n6766) );
  NAND2_X1 U7327 ( .A1(n6762), .A2(n6766), .ZN(n8053) );
  INV_X1 U7328 ( .A(n9618), .ZN(n9623) );
  XNOR2_X1 U7329 ( .A(n9724), .B(n9592), .ZN(n6774) );
  OR2_X1 U7330 ( .A1(n9724), .A2(n9592), .ZN(n6655) );
  OR2_X1 U7331 ( .A1(n9792), .A2(n10056), .ZN(n6656) );
  NAND2_X1 U7332 ( .A1(n9792), .A2(n10056), .ZN(n6776) );
  NAND2_X1 U7333 ( .A1(n6656), .A2(n6776), .ZN(n9587) );
  NAND2_X1 U7334 ( .A1(n9590), .A2(n6776), .ZN(n9573) );
  OR2_X1 U7335 ( .A1(n9714), .A2(n9706), .ZN(n6779) );
  NAND2_X1 U7336 ( .A1(n9714), .A2(n9706), .ZN(n6777) );
  OR2_X1 U7337 ( .A1(n9696), .A2(n9688), .ZN(n6787) );
  OR2_X1 U7338 ( .A1(n9703), .A2(n9524), .ZN(n9527) );
  NAND2_X1 U7339 ( .A1(n6787), .A2(n9527), .ZN(n6707) );
  NAND2_X1 U7340 ( .A1(n9696), .A2(n9688), .ZN(n6788) );
  NAND2_X1 U7341 ( .A1(n9703), .A2(n9524), .ZN(n6782) );
  NAND2_X1 U7342 ( .A1(n6788), .A2(n6782), .ZN(n6708) );
  NAND2_X1 U7343 ( .A1(n6708), .A2(n6787), .ZN(n6667) );
  OR2_X1 U7344 ( .A1(n9685), .A2(n9519), .ZN(n6801) );
  NAND2_X1 U7345 ( .A1(n9685), .A2(n9519), .ZN(n6666) );
  NAND2_X1 U7346 ( .A1(n6801), .A2(n6666), .ZN(n9496) );
  OR2_X1 U7347 ( .A1(n9676), .A2(n9668), .ZN(n6795) );
  NAND2_X1 U7348 ( .A1(n9676), .A2(n9668), .ZN(n6804) );
  NAND2_X1 U7349 ( .A1(n6795), .A2(n6804), .ZN(n6800) );
  INV_X1 U7350 ( .A(n6666), .ZN(n9475) );
  OR2_X1 U7351 ( .A1(n6800), .A2(n9475), .ZN(n6797) );
  NAND2_X1 U7352 ( .A1(n9465), .A2(n9478), .ZN(n6668) );
  NAND2_X1 U7353 ( .A1(n5637), .A2(n9459), .ZN(n9439) );
  NAND2_X1 U7354 ( .A1(n9439), .A2(n6669), .ZN(n9430) );
  NAND2_X1 U7355 ( .A1(n9430), .A2(n4457), .ZN(n9429) );
  NAND2_X1 U7356 ( .A1(n5638), .A2(n9429), .ZN(n9406) );
  NAND2_X1 U7357 ( .A1(n9406), .A2(n6818), .ZN(n5639) );
  XNOR2_X1 U7358 ( .A(n5640), .B(n5639), .ZN(n5654) );
  NAND2_X1 U7359 ( .A1(n4418), .A2(n6678), .ZN(n5642) );
  OR2_X1 U7360 ( .A1(n7849), .A2(n4519), .ZN(n5641) );
  INV_X1 U7361 ( .A(n9876), .ZN(n5644) );
  INV_X1 U7362 ( .A(n5643), .ZN(n6899) );
  INV_X1 U7363 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n5648) );
  INV_X1 U7364 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n5645) );
  OR2_X1 U7365 ( .A1(n4413), .A2(n5645), .ZN(n5647) );
  NAND2_X1 U7366 ( .A1(n6639), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n5646) );
  OAI211_X1 U7367 ( .C1(n5649), .C2(n5648), .A(n5647), .B(n5646), .ZN(n9249)
         );
  INV_X1 U7368 ( .A(P1_B_REG_SCAN_IN), .ZN(n5651) );
  OR2_X1 U7369 ( .A1(n8195), .A2(n5651), .ZN(n9393) );
  NAND3_X1 U7370 ( .A1(n9881), .A2(n9249), .A3(n9393), .ZN(n5652) );
  OAI21_X1 U7371 ( .B1(n9705), .B2(n9432), .A(n5652), .ZN(n5653) );
  AOI21_X1 U7372 ( .B1(n5654), .B2(n9893), .A(n5653), .ZN(n5677) );
  NOR2_X1 U7373 ( .A1(n4417), .A2(n9879), .ZN(n7088) );
  NAND2_X1 U7374 ( .A1(n7491), .A2(n7387), .ZN(n7331) );
  INV_X1 U7375 ( .A(n7756), .ZN(n7915) );
  INV_X1 U7376 ( .A(n9744), .ZN(n7979) );
  NAND2_X1 U7377 ( .A1(n9601), .A2(n9586), .ZN(n9581) );
  OR2_X1 U7378 ( .A1(n9581), .A2(n9714), .ZN(n9565) );
  NAND2_X1 U7379 ( .A1(n9483), .A2(n9669), .ZN(n9450) );
  OAI211_X1 U7380 ( .C1(n5687), .C2(n9416), .A(n9628), .B(n9400), .ZN(n5674)
         );
  MUX2_X1 U7381 ( .A(n5656), .B(n5685), .S(n9906), .Z(n5659) );
  NAND2_X1 U7382 ( .A1(n5661), .A2(n5660), .ZN(P1_U3519) );
  NAND3_X1 U7383 ( .A1(n5663), .A2(n5662), .A3(n6599), .ZN(n5673) );
  NAND2_X1 U7384 ( .A1(n5665), .A2(n7667), .ZN(n6405) );
  INV_X1 U7385 ( .A(n6405), .ZN(n5667) );
  NAND2_X1 U7386 ( .A1(n5667), .A2(n5666), .ZN(n6403) );
  NAND2_X1 U7387 ( .A1(n5668), .A2(n6403), .ZN(n5669) );
  NAND2_X1 U7388 ( .A1(n5684), .A2(n9446), .ZN(n5682) );
  OR2_X1 U7389 ( .A1(n9877), .A2(n7667), .ZN(n6615) );
  INV_X1 U7390 ( .A(n6615), .ZN(n5670) );
  OAI22_X1 U7391 ( .A1(n9560), .A2(n5672), .B1(n5671), .B2(n9886), .ZN(n5676)
         );
  NOR2_X1 U7392 ( .A1(n5674), .A2(n9489), .ZN(n5675) );
  AOI211_X1 U7393 ( .C1(n9620), .C2(n6821), .A(n5676), .B(n5675), .ZN(n5680)
         );
  NAND2_X1 U7394 ( .A1(n5682), .A2(n5681), .ZN(P1_U3356) );
  NAND2_X1 U7395 ( .A1(n5684), .A2(n9711), .ZN(n5690) );
  MUX2_X1 U7396 ( .A(n5686), .B(n5685), .S(n9910), .Z(n5688) );
  NAND2_X1 U7397 ( .A1(n5690), .A2(n5689), .ZN(P1_U3551) );
  NOR2_X1 U7398 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), .ZN(
        n5699) );
  NOR2_X1 U7399 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n5698) );
  NAND4_X1 U7400 ( .A1(n5699), .A2(n5698), .A3(n6093), .A4(n5977), .ZN(n5700)
         );
  NAND4_X1 U7401 ( .A1(n10121), .A2(n10253), .A3(n6114), .A4(n6118), .ZN(n5713) );
  NAND2_X1 U7402 ( .A1(n5703), .A2(n5705), .ZN(n9048) );
  NAND2_X2 U7403 ( .A1(n5707), .A2(n5708), .ZN(n5756) );
  INV_X1 U7404 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n7533) );
  OR2_X1 U7405 ( .A1(n5756), .A2(n7533), .ZN(n5712) );
  INV_X1 U7406 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n6257) );
  INV_X1 U7407 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n6256) );
  NAND4_X2 U7408 ( .A1(n5712), .A2(n5711), .A3(n5710), .A4(n5709), .ZN(n5739)
         );
  NAND2_X1 U7409 ( .A1(n6115), .A2(n5714), .ZN(n6123) );
  INV_X1 U7410 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n5715) );
  INV_X1 U7411 ( .A(n5722), .ZN(n5723) );
  OR2_X1 U7412 ( .A1(n5763), .A2(n6917), .ZN(n5726) );
  NAND2_X1 U7413 ( .A1(n6061), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5731) );
  INV_X1 U7414 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n7125) );
  OR2_X1 U7415 ( .A1(n5756), .A2(n7125), .ZN(n5730) );
  INV_X1 U7416 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n6210) );
  OR2_X1 U7417 ( .A1(n5757), .A2(n6210), .ZN(n5729) );
  INV_X1 U7418 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n7360) );
  NAND2_X1 U7419 ( .A1(n5732), .A2(SI_0_), .ZN(n5734) );
  INV_X1 U7420 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5733) );
  NAND2_X1 U7421 ( .A1(n5734), .A2(n5733), .ZN(n5736) );
  AND2_X1 U7422 ( .A1(n5736), .A2(n5735), .ZN(n9049) );
  MUX2_X1 U7423 ( .A(n9911), .B(n9049), .S(n5737), .Z(n7535) );
  NAND2_X1 U7424 ( .A1(n7537), .A2(n7535), .ZN(n5738) );
  OR2_X1 U7425 ( .A1(n5739), .A2(n5740), .ZN(n9945) );
  NAND2_X1 U7426 ( .A1(n7534), .A2(n9945), .ZN(n5754) );
  INV_X2 U7427 ( .A(n5774), .ZN(n5796) );
  INV_X1 U7428 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n5741) );
  INV_X1 U7429 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n9942) );
  OR2_X1 U7430 ( .A1(n5756), .A2(n9942), .ZN(n5743) );
  INV_X1 U7431 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n6214) );
  OAI22_X1 U7432 ( .A1(n5722), .A2(n5746), .B1(P2_IR_REG_2__SCAN_IN), .B2(
        P2_IR_REG_31__SCAN_IN), .ZN(n5747) );
  INV_X1 U7433 ( .A(n5747), .ZN(n5749) );
  OR2_X1 U7434 ( .A1(n5737), .A2(n7021), .ZN(n5752) );
  OR2_X1 U7435 ( .A1(n5764), .A2(n6913), .ZN(n5751) );
  OR2_X1 U7436 ( .A1(n5763), .A2(n6923), .ZN(n5750) );
  NAND2_X1 U7437 ( .A1(n5755), .A2(n9966), .ZN(n8262) );
  NAND2_X1 U7438 ( .A1(n5754), .A2(n8268), .ZN(n7376) );
  OR2_X1 U7439 ( .A1(n5755), .A2(n5753), .ZN(n7377) );
  NAND2_X1 U7440 ( .A1(n7376), .A2(n7377), .ZN(n5771) );
  NAND2_X1 U7441 ( .A1(n6061), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5762) );
  OR2_X1 U7442 ( .A1(n5774), .A2(n7056), .ZN(n5761) );
  OR2_X1 U7443 ( .A1(n5756), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n5760) );
  INV_X1 U7444 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n5758) );
  OR2_X1 U7445 ( .A1(n8208), .A2(n5758), .ZN(n5759) );
  OR2_X1 U7446 ( .A1(n5763), .A2(n6920), .ZN(n5770) );
  OR2_X1 U7447 ( .A1(n5764), .A2(n10272), .ZN(n5769) );
  MUX2_X1 U7448 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5765), .S(
        P2_IR_REG_3__SCAN_IN), .Z(n5767) );
  NAND2_X1 U7449 ( .A1(n5767), .A2(n5766), .ZN(n7054) );
  OR2_X1 U7450 ( .A1(n5737), .A2(n7054), .ZN(n5768) );
  NAND2_X1 U7451 ( .A1(n5772), .A2(n9972), .ZN(n8263) );
  NAND2_X1 U7452 ( .A1(n8261), .A2(n8263), .ZN(n7373) );
  NAND2_X1 U7453 ( .A1(n5771), .A2(n7373), .ZN(n7375) );
  INV_X1 U7454 ( .A(n5772), .ZN(n9952) );
  INV_X1 U7455 ( .A(n9972), .ZN(n7381) );
  OR2_X1 U7456 ( .A1(n5772), .A2(n7381), .ZN(n5773) );
  NAND2_X1 U7457 ( .A1(n6061), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n5779) );
  OR2_X1 U7458 ( .A1(n5774), .A2(n6317), .ZN(n5778) );
  NAND2_X1 U7459 ( .A1(n10082), .A2(n7380), .ZN(n5785) );
  NAND2_X1 U7460 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n5775) );
  AND2_X1 U7461 ( .A1(n5785), .A2(n5775), .ZN(n7285) );
  OR2_X1 U7462 ( .A1(n5756), .A2(n7285), .ZN(n5777) );
  OR2_X1 U7463 ( .A1(n8208), .A2(n6217), .ZN(n5776) );
  NAND2_X1 U7464 ( .A1(n5766), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5780) );
  OR2_X1 U7465 ( .A1(n5763), .A2(n6931), .ZN(n5782) );
  OR2_X1 U7466 ( .A1(n5764), .A2(n10270), .ZN(n5781) );
  OAI211_X1 U7467 ( .C1(n5737), .C2(n9937), .A(n5782), .B(n5781), .ZN(n7434)
         );
  NOR2_X1 U7468 ( .A1(n8592), .A2(n7434), .ZN(n6157) );
  NAND2_X1 U7469 ( .A1(n8592), .A2(n7434), .ZN(n6158) );
  NAND2_X1 U7470 ( .A1(n6061), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5791) );
  INV_X1 U7471 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n7517) );
  OR2_X1 U7472 ( .A1(n5774), .A2(n7517), .ZN(n5790) );
  INV_X1 U7473 ( .A(n5785), .ZN(n5784) );
  NAND2_X1 U7474 ( .A1(n5784), .A2(n5783), .ZN(n5799) );
  NAND2_X1 U7475 ( .A1(n5785), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5786) );
  AND2_X1 U7476 ( .A1(n5799), .A2(n5786), .ZN(n7518) );
  OR2_X1 U7477 ( .A1(n5756), .A2(n7518), .ZN(n5789) );
  INV_X1 U7478 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n5787) );
  OR2_X1 U7479 ( .A1(n8208), .A2(n5787), .ZN(n5788) );
  NAND4_X1 U7480 ( .A1(n5791), .A2(n5790), .A3(n5789), .A4(n5788), .ZN(n8591)
         );
  OR2_X1 U7481 ( .A1(n5792), .A2(n5715), .ZN(n5793) );
  INV_X1 U7482 ( .A(n6320), .ZN(n7126) );
  OR2_X1 U7483 ( .A1(n5763), .A2(n6929), .ZN(n5795) );
  INV_X1 U7484 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6914) );
  OR2_X1 U7485 ( .A1(n5764), .A2(n6914), .ZN(n5794) );
  OAI211_X1 U7486 ( .C1(n5737), .C2(n7126), .A(n5795), .B(n5794), .ZN(n7520)
         );
  AND2_X1 U7487 ( .A1(n8591), .A2(n7520), .ZN(n7512) );
  OR2_X1 U7488 ( .A1(n8591), .A2(n7520), .ZN(n7511) );
  NAND2_X1 U7489 ( .A1(n5796), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n5805) );
  INV_X1 U7490 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n5798) );
  OR2_X1 U7491 ( .A1(n5797), .A2(n5798), .ZN(n5804) );
  NAND2_X1 U7492 ( .A1(n5799), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5800) );
  AND2_X1 U7493 ( .A1(n5814), .A2(n5800), .ZN(n7582) );
  OR2_X1 U7494 ( .A1(n5756), .A2(n7582), .ZN(n5803) );
  INV_X1 U7495 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n5801) );
  OR2_X1 U7496 ( .A1(n8208), .A2(n5801), .ZN(n5802) );
  NAND4_X1 U7497 ( .A1(n5805), .A2(n5804), .A3(n5803), .A4(n5802), .ZN(n8590)
         );
  OR2_X1 U7498 ( .A1(n5806), .A2(n5715), .ZN(n5808) );
  XNOR2_X1 U7499 ( .A(n5808), .B(n5807), .ZN(n7237) );
  OR2_X1 U7500 ( .A1(n5763), .A2(n6927), .ZN(n5810) );
  OR2_X1 U7501 ( .A1(n5764), .A2(n10343), .ZN(n5809) );
  OAI211_X1 U7502 ( .C1(n5737), .C2(n7237), .A(n5810), .B(n5809), .ZN(n8278)
         );
  NOR2_X1 U7503 ( .A1(n8590), .A2(n8278), .ZN(n7563) );
  NAND2_X1 U7504 ( .A1(n8590), .A2(n8278), .ZN(n7561) );
  OAI21_X2 U7505 ( .B1(n7565), .B2(n7563), .A(n7561), .ZN(n7550) );
  NAND2_X1 U7506 ( .A1(n6061), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5819) );
  INV_X1 U7507 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n5811) );
  OR2_X1 U7508 ( .A1(n5774), .A2(n5811), .ZN(n5818) );
  NAND2_X1 U7509 ( .A1(n5814), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5815) );
  AND2_X1 U7510 ( .A1(n5827), .A2(n5815), .ZN(n7555) );
  OR2_X1 U7511 ( .A1(n5756), .A2(n7555), .ZN(n5817) );
  OR2_X1 U7512 ( .A1(n8208), .A2(n7306), .ZN(n5816) );
  NAND4_X1 U7513 ( .A1(n5819), .A2(n5818), .A3(n5817), .A4(n5816), .ZN(n8589)
         );
  OR2_X1 U7514 ( .A1(n5763), .A2(n6925), .ZN(n5824) );
  OR2_X1 U7515 ( .A1(n5764), .A2(n6919), .ZN(n5823) );
  NAND2_X1 U7516 ( .A1(n5820), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5821) );
  XNOR2_X1 U7517 ( .A(n5821), .B(n4957), .ZN(n7310) );
  OR2_X1 U7518 ( .A1(n5737), .A2(n7310), .ZN(n5822) );
  XNOR2_X1 U7519 ( .A(n8589), .B(n8304), .ZN(n7553) );
  INV_X1 U7520 ( .A(n8304), .ZN(n7676) );
  NAND2_X1 U7521 ( .A1(n8589), .A2(n7676), .ZN(n5825) );
  NAND2_X1 U7522 ( .A1(n5796), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n5832) );
  INV_X1 U7523 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n5826) );
  OR2_X1 U7524 ( .A1(n5797), .A2(n5826), .ZN(n5831) );
  NAND2_X1 U7525 ( .A1(n5827), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5828) );
  AND2_X1 U7526 ( .A1(n5839), .A2(n5828), .ZN(n7690) );
  OR2_X1 U7527 ( .A1(n5756), .A2(n7690), .ZN(n5830) );
  OR2_X1 U7528 ( .A1(n8208), .A2(n6226), .ZN(n5829) );
  NAND4_X1 U7529 ( .A1(n5832), .A2(n5831), .A3(n5830), .A4(n5829), .ZN(n8588)
         );
  NAND2_X1 U7530 ( .A1(n6933), .A2(n8202), .ZN(n5835) );
  NAND2_X1 U7531 ( .A1(n4447), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5833) );
  XNOR2_X1 U7532 ( .A(n5833), .B(P2_IR_REG_8__SCAN_IN), .ZN(n6327) );
  AOI22_X1 U7533 ( .A1(n8201), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n6209), .B2(
        n6327), .ZN(n5834) );
  NAND2_X1 U7534 ( .A1(n8588), .A2(n9994), .ZN(n8298) );
  NAND2_X1 U7535 ( .A1(n8303), .A2(n8298), .ZN(n8221) );
  NAND2_X1 U7536 ( .A1(n6061), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5845) );
  INV_X1 U7537 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n5836) );
  OR2_X1 U7538 ( .A1(n5774), .A2(n5836), .ZN(n5844) );
  NAND2_X1 U7539 ( .A1(n5839), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n5840) );
  AND2_X1 U7540 ( .A1(n5853), .A2(n5840), .ZN(n7807) );
  OR2_X1 U7541 ( .A1(n5756), .A2(n7807), .ZN(n5843) );
  INV_X1 U7542 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n5841) );
  OR2_X1 U7543 ( .A1(n8208), .A2(n5841), .ZN(n5842) );
  NAND2_X1 U7544 ( .A1(n6937), .A2(n8202), .ZN(n5848) );
  OR2_X1 U7545 ( .A1(n4447), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n5849) );
  NAND2_X1 U7546 ( .A1(n5849), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5846) );
  XNOR2_X1 U7547 ( .A(n5846), .B(P2_IR_REG_9__SCAN_IN), .ZN(n7655) );
  AOI22_X1 U7548 ( .A1(n8201), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6209), .B2(
        n7655), .ZN(n5847) );
  NAND2_X1 U7549 ( .A1(n5848), .A2(n5847), .ZN(n7950) );
  NAND2_X1 U7550 ( .A1(n7991), .A2(n7950), .ZN(n8306) );
  NAND2_X1 U7551 ( .A1(n6942), .A2(n8202), .ZN(n5852) );
  OR2_X1 U7552 ( .A1(n5861), .A2(n5715), .ZN(n5850) );
  INV_X1 U7553 ( .A(n6943), .ZN(n7766) );
  AOI22_X1 U7554 ( .A1(n8201), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6209), .B2(
        n7766), .ZN(n5851) );
  NAND2_X1 U7555 ( .A1(n5852), .A2(n5851), .ZN(n7996) );
  NAND2_X1 U7556 ( .A1(n6061), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5859) );
  INV_X1 U7557 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7905) );
  OR2_X1 U7558 ( .A1(n5774), .A2(n7905), .ZN(n5858) );
  NAND2_X1 U7559 ( .A1(n5853), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5854) );
  AND2_X1 U7560 ( .A1(n5868), .A2(n5854), .ZN(n7995) );
  OR2_X1 U7561 ( .A1(n5756), .A2(n7995), .ZN(n5857) );
  INV_X1 U7562 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n5855) );
  OR2_X1 U7563 ( .A1(n8208), .A2(n5855), .ZN(n5856) );
  NAND4_X1 U7564 ( .A1(n5859), .A2(n5858), .A3(n5857), .A4(n5856), .ZN(n8586)
         );
  AND2_X1 U7565 ( .A1(n7996), .A2(n8586), .ZN(n5878) );
  OR2_X1 U7566 ( .A1(n8225), .A2(n5878), .ZN(n7870) );
  NAND2_X1 U7567 ( .A1(n6947), .A2(n8202), .ZN(n5866) );
  NAND2_X1 U7568 ( .A1(n5861), .A2(n5860), .ZN(n5863) );
  NAND2_X1 U7569 ( .A1(n5863), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5862) );
  MUX2_X1 U7570 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5862), .S(
        P2_IR_REG_11__SCAN_IN), .Z(n5864) );
  AOI22_X1 U7571 ( .A1(n8201), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n6209), .B2(
        n7933), .ZN(n5865) );
  NAND2_X1 U7572 ( .A1(n5866), .A2(n5865), .ZN(n8071) );
  NAND2_X1 U7573 ( .A1(n6061), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5874) );
  INV_X1 U7574 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n5867) );
  OR2_X1 U7575 ( .A1(n5774), .A2(n5867), .ZN(n5873) );
  NAND2_X1 U7576 ( .A1(n5868), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5869) );
  AND2_X1 U7577 ( .A1(n5887), .A2(n5869), .ZN(n8067) );
  OR2_X1 U7578 ( .A1(n5756), .A2(n8067), .ZN(n5872) );
  INV_X1 U7579 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n5870) );
  OR2_X1 U7580 ( .A1(n8208), .A2(n5870), .ZN(n5871) );
  INV_X1 U7581 ( .A(n8063), .ZN(n8011) );
  AND2_X1 U7582 ( .A1(n8071), .A2(n8011), .ZN(n5880) );
  OR2_X1 U7583 ( .A1(n7870), .A2(n5880), .ZN(n5875) );
  NAND2_X1 U7584 ( .A1(n8071), .A2(n8063), .ZN(n8319) );
  NAND2_X1 U7585 ( .A1(n8317), .A2(n8319), .ZN(n8228) );
  OR2_X1 U7586 ( .A1(n7996), .A2(n8586), .ZN(n5876) );
  OR2_X1 U7587 ( .A1(n7950), .A2(n8587), .ZN(n7899) );
  AND2_X1 U7588 ( .A1(n5876), .A2(n7899), .ZN(n5877) );
  OR2_X1 U7589 ( .A1(n5878), .A2(n5877), .ZN(n7871) );
  AND2_X1 U7590 ( .A1(n8228), .A2(n7871), .ZN(n5879) );
  OR2_X1 U7591 ( .A1(n5880), .A2(n5879), .ZN(n5881) );
  OAI21_X1 U7592 ( .B1(n7801), .B2(n5875), .A(n5881), .ZN(n5882) );
  NAND2_X1 U7593 ( .A1(n6952), .A2(n8202), .ZN(n5885) );
  NAND2_X1 U7594 ( .A1(n5895), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5883) );
  XNOR2_X1 U7595 ( .A(n5883), .B(P2_IR_REG_12__SCAN_IN), .ZN(n8627) );
  AOI22_X1 U7596 ( .A1(n8201), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6209), .B2(
        n8627), .ZN(n5884) );
  NAND2_X1 U7597 ( .A1(n6061), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5893) );
  OR2_X1 U7598 ( .A1(n5774), .A2(n6335), .ZN(n5892) );
  NAND2_X1 U7599 ( .A1(n5887), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5888) );
  AND2_X1 U7600 ( .A1(n5901), .A2(n5888), .ZN(n8017) );
  OR2_X1 U7601 ( .A1(n5756), .A2(n8017), .ZN(n5891) );
  INV_X1 U7602 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n5889) );
  OR2_X1 U7603 ( .A1(n8208), .A2(n5889), .ZN(n5890) );
  NAND4_X1 U7604 ( .A1(n5893), .A2(n5892), .A3(n5891), .A4(n5890), .ZN(n8585)
         );
  AND2_X1 U7605 ( .A1(n10014), .A2(n8585), .ZN(n5894) );
  NAND2_X1 U7606 ( .A1(n6956), .A2(n8202), .ZN(n5897) );
  OAI21_X1 U7607 ( .B1(n5895), .B2(P2_IR_REG_12__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5911) );
  AOI22_X1 U7608 ( .A1(n8201), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6209), .B2(
        n8643), .ZN(n5896) );
  NAND2_X1 U7609 ( .A1(n6061), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5907) );
  INV_X1 U7610 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n5898) );
  OR2_X1 U7611 ( .A1(n8208), .A2(n5898), .ZN(n5906) );
  NAND2_X1 U7612 ( .A1(n5901), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n5902) );
  AND2_X1 U7613 ( .A1(n5918), .A2(n5902), .ZN(n8094) );
  OR2_X1 U7614 ( .A1(n5756), .A2(n8094), .ZN(n5905) );
  INV_X1 U7615 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n5903) );
  OR2_X1 U7616 ( .A1(n5774), .A2(n5903), .ZN(n5904) );
  NAND4_X1 U7617 ( .A1(n5907), .A2(n5906), .A3(n5905), .A4(n5904), .ZN(n8584)
         );
  NOR2_X1 U7618 ( .A1(n8096), .A2(n8584), .ZN(n5909) );
  NAND2_X1 U7619 ( .A1(n8096), .A2(n8584), .ZN(n5908) );
  NAND2_X1 U7620 ( .A1(n7014), .A2(n8202), .ZN(n5917) );
  INV_X1 U7621 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5910) );
  NAND2_X1 U7622 ( .A1(n5911), .A2(n5910), .ZN(n5912) );
  NAND2_X1 U7623 ( .A1(n5912), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5914) );
  INV_X1 U7624 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5913) );
  NAND2_X1 U7625 ( .A1(n5914), .A2(n5913), .ZN(n5925) );
  OR2_X1 U7626 ( .A1(n5914), .A2(n5913), .ZN(n5915) );
  AOI22_X1 U7627 ( .A1(n8201), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n6209), .B2(
        n8656), .ZN(n5916) );
  NAND2_X1 U7628 ( .A1(n5917), .A2(n5916), .ZN(n8145) );
  NAND2_X1 U7629 ( .A1(n6061), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5923) );
  INV_X1 U7630 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n6339) );
  OR2_X1 U7631 ( .A1(n5774), .A2(n6339), .ZN(n5922) );
  NAND2_X1 U7632 ( .A1(n5918), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5919) );
  AND2_X1 U7633 ( .A1(n5931), .A2(n5919), .ZN(n8451) );
  OR2_X1 U7634 ( .A1(n5756), .A2(n8451), .ZN(n5921) );
  INV_X1 U7635 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n6235) );
  OR2_X1 U7636 ( .A1(n8208), .A2(n6235), .ZN(n5920) );
  NAND4_X1 U7637 ( .A1(n5923), .A2(n5922), .A3(n5921), .A4(n5920), .ZN(n8908)
         );
  AND2_X1 U7638 ( .A1(n8145), .A2(n8908), .ZN(n5924) );
  NAND2_X1 U7639 ( .A1(n7019), .A2(n8202), .ZN(n5928) );
  NAND2_X1 U7640 ( .A1(n5925), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5926) );
  XNOR2_X1 U7641 ( .A(n5926), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8674) );
  AOI22_X1 U7642 ( .A1(n8674), .A2(n6209), .B1(n8201), .B2(
        P1_DATAO_REG_15__SCAN_IN), .ZN(n5927) );
  NAND2_X1 U7643 ( .A1(n6061), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n5936) );
  INV_X1 U7644 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n8965) );
  OR2_X1 U7645 ( .A1(n8208), .A2(n8965), .ZN(n5935) );
  NAND2_X1 U7646 ( .A1(n5931), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5932) );
  AND2_X1 U7647 ( .A1(n5941), .A2(n5932), .ZN(n8915) );
  OR2_X1 U7648 ( .A1(n5756), .A2(n8915), .ZN(n5934) );
  INV_X1 U7649 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n8914) );
  OR2_X1 U7650 ( .A1(n5774), .A2(n8914), .ZN(n5933) );
  NAND4_X1 U7651 ( .A1(n5936), .A2(n5935), .A3(n5934), .A4(n5933), .ZN(n8894)
         );
  NAND2_X1 U7652 ( .A1(n9037), .A2(n8894), .ZN(n8890) );
  NAND2_X1 U7653 ( .A1(n7163), .A2(n8202), .ZN(n5940) );
  NAND2_X1 U7654 ( .A1(n5937), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5938) );
  XNOR2_X1 U7655 ( .A(n5938), .B(P2_IR_REG_16__SCAN_IN), .ZN(n8688) );
  AOI22_X1 U7656 ( .A1(n8201), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n6209), .B2(
        n8688), .ZN(n5939) );
  NAND2_X1 U7657 ( .A1(n6061), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n5946) );
  INV_X1 U7658 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8899) );
  OR2_X1 U7659 ( .A1(n5774), .A2(n8899), .ZN(n5945) );
  NAND2_X1 U7660 ( .A1(n5941), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5942) );
  AND2_X1 U7661 ( .A1(n5955), .A2(n5942), .ZN(n8498) );
  OR2_X1 U7662 ( .A1(n5756), .A2(n8498), .ZN(n5944) );
  INV_X1 U7663 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8962) );
  OR2_X1 U7664 ( .A1(n8208), .A2(n8962), .ZN(n5943) );
  NAND2_X1 U7665 ( .A1(n9031), .A2(n8910), .ZN(n5947) );
  AND2_X1 U7666 ( .A1(n8890), .A2(n5947), .ZN(n5949) );
  INV_X1 U7667 ( .A(n5947), .ZN(n5948) );
  NAND2_X1 U7668 ( .A1(n9031), .A2(n8565), .ZN(n8340) );
  NAND2_X1 U7669 ( .A1(n8350), .A2(n8340), .ZN(n8888) );
  NAND2_X1 U7670 ( .A1(n7250), .A2(n8202), .ZN(n5952) );
  NOR2_X1 U7671 ( .A1(n5937), .A2(P2_IR_REG_16__SCAN_IN), .ZN(n5964) );
  OR2_X1 U7672 ( .A1(n5964), .A2(n5715), .ZN(n5950) );
  XNOR2_X1 U7673 ( .A(n5950), .B(P2_IR_REG_17__SCAN_IN), .ZN(n8708) );
  AOI22_X1 U7674 ( .A1(n8201), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n6209), .B2(
        n8708), .ZN(n5951) );
  INV_X1 U7675 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8883) );
  OR2_X1 U7676 ( .A1(n5774), .A2(n8883), .ZN(n5960) );
  INV_X1 U7677 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n10086) );
  OR2_X1 U7678 ( .A1(n5797), .A2(n10086), .ZN(n5959) );
  NAND2_X1 U7679 ( .A1(n5955), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n5956) );
  AND2_X1 U7680 ( .A1(n5968), .A2(n5956), .ZN(n8507) );
  OR2_X1 U7681 ( .A1(n5756), .A2(n8507), .ZN(n5958) );
  INV_X1 U7682 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n8959) );
  OR2_X1 U7683 ( .A1(n8208), .A2(n8959), .ZN(n5957) );
  OR2_X1 U7684 ( .A1(n9025), .A2(n8896), .ZN(n8355) );
  NAND2_X1 U7685 ( .A1(n9025), .A2(n8896), .ZN(n8342) );
  NAND2_X1 U7686 ( .A1(n8355), .A2(n8342), .ZN(n8341) );
  NAND2_X1 U7687 ( .A1(n8879), .A2(n8341), .ZN(n5962) );
  INV_X1 U7688 ( .A(n8896), .ZN(n8583) );
  NAND2_X1 U7689 ( .A1(n9025), .A2(n8583), .ZN(n5961) );
  NAND2_X1 U7690 ( .A1(n5962), .A2(n5961), .ZN(n8866) );
  NAND2_X1 U7691 ( .A1(n7275), .A2(n8202), .ZN(n5967) );
  NAND2_X1 U7692 ( .A1(n5964), .A2(n5963), .ZN(n5975) );
  NAND2_X1 U7693 ( .A1(n5975), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5965) );
  XNOR2_X1 U7694 ( .A(n5965), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8730) );
  AOI22_X1 U7695 ( .A1(n8201), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6209), .B2(
        n8730), .ZN(n5966) );
  NAND2_X1 U7696 ( .A1(n5968), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5969) );
  NAND2_X1 U7697 ( .A1(n5983), .A2(n5969), .ZN(n8873) );
  NAND2_X1 U7698 ( .A1(n6101), .A2(n8873), .ZN(n5973) );
  INV_X1 U7699 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n6345) );
  OR2_X1 U7700 ( .A1(n5774), .A2(n6345), .ZN(n5972) );
  INV_X1 U7701 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n9020) );
  OR2_X1 U7702 ( .A1(n5797), .A2(n9020), .ZN(n5971) );
  INV_X1 U7703 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n10276) );
  OR2_X1 U7704 ( .A1(n8208), .A2(n10276), .ZN(n5970) );
  NAND4_X1 U7705 ( .A1(n5973), .A2(n5972), .A3(n5971), .A4(n5970), .ZN(n8881)
         );
  AND2_X1 U7706 ( .A1(n8956), .A2(n8881), .ZN(n5974) );
  NAND2_X1 U7707 ( .A1(n7544), .A2(n8202), .ZN(n5980) );
  INV_X1 U7708 ( .A(n6091), .ZN(n5976) );
  NAND2_X1 U7709 ( .A1(n5976), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5978) );
  AOI22_X1 U7710 ( .A1(n8201), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n8420), .B2(
        n6209), .ZN(n5979) );
  INV_X1 U7711 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n5981) );
  NAND2_X1 U7712 ( .A1(n5983), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n5984) );
  NAND2_X1 U7713 ( .A1(n5995), .A2(n5984), .ZN(n8861) );
  NAND2_X1 U7714 ( .A1(n6101), .A2(n8861), .ZN(n5989) );
  INV_X1 U7715 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n5985) );
  OR2_X1 U7716 ( .A1(n5774), .A2(n5985), .ZN(n5988) );
  INV_X1 U7717 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n9016) );
  OR2_X1 U7718 ( .A1(n5797), .A2(n9016), .ZN(n5987) );
  INV_X1 U7719 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n8953) );
  OR2_X1 U7720 ( .A1(n8208), .A2(n8953), .ZN(n5986) );
  NAND2_X1 U7721 ( .A1(n8952), .A2(n8868), .ZN(n8359) );
  INV_X1 U7722 ( .A(n8868), .ZN(n8582) );
  NAND2_X1 U7723 ( .A1(n8952), .A2(n8582), .ZN(n5990) );
  NAND2_X1 U7724 ( .A1(n7648), .A2(n8202), .ZN(n5992) );
  INV_X1 U7725 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7649) );
  OR2_X1 U7726 ( .A1(n5764), .A2(n7649), .ZN(n5991) );
  INV_X1 U7727 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n10314) );
  OR2_X1 U7728 ( .A1(n5774), .A2(n10314), .ZN(n5994) );
  INV_X1 U7729 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n9011) );
  OR2_X1 U7730 ( .A1(n5797), .A2(n9011), .ZN(n5993) );
  AND2_X1 U7731 ( .A1(n5994), .A2(n5993), .ZN(n5999) );
  OR2_X2 U7732 ( .A1(n5995), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n6005) );
  NAND2_X1 U7733 ( .A1(n5995), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n5996) );
  NAND2_X1 U7734 ( .A1(n6005), .A2(n5996), .ZN(n8844) );
  NAND2_X1 U7735 ( .A1(n8844), .A2(n6101), .ZN(n5998) );
  INV_X1 U7736 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n10195) );
  OR2_X1 U7737 ( .A1(n8208), .A2(n10195), .ZN(n5997) );
  NAND2_X1 U7738 ( .A1(n8521), .A2(n8856), .ZN(n8828) );
  INV_X1 U7739 ( .A(n8856), .ZN(n8581) );
  OR2_X1 U7740 ( .A1(n8521), .A2(n8581), .ZN(n6001) );
  NAND2_X1 U7741 ( .A1(n8837), .A2(n6001), .ZN(n8825) );
  NAND2_X1 U7742 ( .A1(n7693), .A2(n8202), .ZN(n6003) );
  OR2_X1 U7743 ( .A1(n5764), .A2(n7694), .ZN(n6002) );
  NAND2_X1 U7744 ( .A1(n6005), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n6006) );
  NAND2_X1 U7745 ( .A1(n6014), .A2(n6006), .ZN(n8832) );
  NAND2_X1 U7746 ( .A1(n8832), .A2(n6101), .ZN(n6009) );
  AOI22_X1 U7747 ( .A1(n5796), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n6061), .B2(
        P2_REG0_REG_21__SCAN_IN), .ZN(n6008) );
  NAND2_X1 U7748 ( .A1(n6060), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n6007) );
  NAND2_X1 U7749 ( .A1(n8478), .A2(n8841), .ZN(n8367) );
  NAND2_X1 U7750 ( .A1(n8366), .A2(n8367), .ZN(n8215) );
  NAND2_X1 U7751 ( .A1(n8825), .A2(n8215), .ZN(n6011) );
  OR2_X1 U7752 ( .A1(n8478), .A2(n8818), .ZN(n6010) );
  NAND2_X1 U7753 ( .A1(n6011), .A2(n6010), .ZN(n8816) );
  NAND2_X1 U7754 ( .A1(n7847), .A2(n8202), .ZN(n6013) );
  OR2_X1 U7755 ( .A1(n5764), .A2(n10344), .ZN(n6012) );
  NAND2_X1 U7756 ( .A1(n6014), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6015) );
  NAND2_X1 U7757 ( .A1(n6023), .A2(n6015), .ZN(n8822) );
  NAND2_X1 U7758 ( .A1(n8822), .A2(n6101), .ZN(n6018) );
  AOI22_X1 U7759 ( .A1(n5796), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n6061), .B2(
        P2_REG0_REG_22__SCAN_IN), .ZN(n6017) );
  NAND2_X1 U7760 ( .A1(n6060), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n6016) );
  NAND2_X1 U7761 ( .A1(n9002), .A2(n8827), .ZN(n8245) );
  NAND2_X1 U7762 ( .A1(n8242), .A2(n8245), .ZN(n8817) );
  NAND2_X1 U7763 ( .A1(n8816), .A2(n8817), .ZN(n6020) );
  OR2_X1 U7764 ( .A1(n9002), .A2(n8807), .ZN(n6019) );
  NAND2_X1 U7765 ( .A1(n6020), .A2(n6019), .ZN(n8805) );
  NAND2_X1 U7766 ( .A1(n7943), .A2(n8202), .ZN(n6022) );
  OR2_X1 U7767 ( .A1(n5764), .A2(n7946), .ZN(n6021) );
  NAND2_X1 U7768 ( .A1(n6023), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6024) );
  NAND2_X1 U7769 ( .A1(n6036), .A2(n6024), .ZN(n8810) );
  NAND2_X1 U7770 ( .A1(n8810), .A2(n6101), .ZN(n6029) );
  INV_X1 U7771 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n8937) );
  NAND2_X1 U7772 ( .A1(n5796), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n6026) );
  NAND2_X1 U7773 ( .A1(n6061), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n6025) );
  OAI211_X1 U7774 ( .C1(n8937), .C2(n8208), .A(n6026), .B(n6025), .ZN(n6027)
         );
  INV_X1 U7775 ( .A(n6027), .ZN(n6028) );
  NOR2_X1 U7776 ( .A1(n8805), .A2(n6030), .ZN(n6031) );
  NAND2_X1 U7777 ( .A1(n8005), .A2(n8202), .ZN(n6033) );
  OR2_X1 U7778 ( .A1(n5764), .A2(n10235), .ZN(n6032) );
  INV_X1 U7779 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n6034) );
  NAND2_X1 U7780 ( .A1(n6036), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n6037) );
  NAND2_X1 U7781 ( .A1(n6049), .A2(n6037), .ZN(n8797) );
  NAND2_X1 U7782 ( .A1(n8797), .A2(n6101), .ZN(n6043) );
  INV_X1 U7783 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n6040) );
  NAND2_X1 U7784 ( .A1(n6061), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n6039) );
  NAND2_X1 U7785 ( .A1(n6060), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n6038) );
  OAI211_X1 U7786 ( .C1(n5774), .C2(n6040), .A(n6039), .B(n6038), .ZN(n6041)
         );
  INV_X1 U7787 ( .A(n6041), .ZN(n6042) );
  NOR2_X1 U7788 ( .A1(n8991), .A2(n8806), .ZN(n6044) );
  NAND2_X1 U7789 ( .A1(n8080), .A2(n8202), .ZN(n6046) );
  OR2_X1 U7790 ( .A1(n5764), .A2(n8133), .ZN(n6045) );
  INV_X1 U7791 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n6047) );
  NAND2_X1 U7792 ( .A1(n6049), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n6050) );
  NAND2_X1 U7793 ( .A1(n6058), .A2(n6050), .ZN(n8782) );
  NAND2_X1 U7794 ( .A1(n8782), .A2(n6101), .ZN(n6055) );
  INV_X1 U7795 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n8931) );
  NAND2_X1 U7796 ( .A1(n5796), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n6052) );
  NAND2_X1 U7797 ( .A1(n6061), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n6051) );
  OAI211_X1 U7798 ( .C1(n8931), .C2(n8208), .A(n6052), .B(n6051), .ZN(n6053)
         );
  INV_X1 U7799 ( .A(n6053), .ZN(n6054) );
  NAND2_X1 U7800 ( .A1(n8985), .A2(n8176), .ZN(n8380) );
  NAND2_X1 U7801 ( .A1(n8125), .A2(n8202), .ZN(n6057) );
  NAND2_X1 U7802 ( .A1(n6058), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n6059) );
  NAND2_X1 U7803 ( .A1(n6073), .A2(n6059), .ZN(n8771) );
  NAND2_X1 U7804 ( .A1(n8771), .A2(n6101), .ZN(n6066) );
  INV_X1 U7805 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n8770) );
  NAND2_X1 U7806 ( .A1(n6060), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n6063) );
  NAND2_X1 U7807 ( .A1(n6061), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n6062) );
  OAI211_X1 U7808 ( .C1(n5774), .C2(n8770), .A(n6063), .B(n6062), .ZN(n6064)
         );
  INV_X1 U7809 ( .A(n6064), .ZN(n6065) );
  NOR2_X1 U7810 ( .A1(n8979), .A2(n8775), .ZN(n6068) );
  INV_X1 U7811 ( .A(n8979), .ZN(n6067) );
  NAND2_X1 U7812 ( .A1(n8194), .A2(n8202), .ZN(n6070) );
  INV_X1 U7813 ( .A(n6073), .ZN(n6072) );
  INV_X1 U7814 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n6071) );
  NAND2_X1 U7815 ( .A1(n6072), .A2(n6071), .ZN(n6083) );
  NAND2_X1 U7816 ( .A1(n6073), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n6074) );
  NAND2_X1 U7817 ( .A1(n6083), .A2(n6074), .ZN(n8757) );
  NAND2_X1 U7818 ( .A1(n8757), .A2(n6101), .ZN(n6079) );
  INV_X1 U7819 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n6192) );
  NAND2_X1 U7820 ( .A1(n5796), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n6076) );
  NAND2_X1 U7821 ( .A1(n6061), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n6075) );
  OAI211_X1 U7822 ( .C1(n6192), .C2(n8208), .A(n6076), .B(n6075), .ZN(n6077)
         );
  INV_X1 U7823 ( .A(n6077), .ZN(n6078) );
  NAND2_X1 U7824 ( .A1(n8183), .A2(n8561), .ZN(n8389) );
  NAND2_X1 U7825 ( .A1(n6080), .A2(n8202), .ZN(n6082) );
  OR2_X1 U7826 ( .A1(n5764), .A2(n10301), .ZN(n6081) );
  NAND2_X1 U7827 ( .A1(n6083), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n6084) );
  NAND2_X1 U7828 ( .A1(n6100), .A2(n6084), .ZN(n8187) );
  NAND2_X1 U7829 ( .A1(n8187), .A2(n6101), .ZN(n6089) );
  INV_X1 U7830 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n6154) );
  NAND2_X1 U7831 ( .A1(n5796), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n6086) );
  NAND2_X1 U7832 ( .A1(n6061), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n6085) );
  OAI211_X1 U7833 ( .C1(n6154), .C2(n8208), .A(n6086), .B(n6085), .ZN(n6087)
         );
  INV_X1 U7834 ( .A(n6087), .ZN(n6088) );
  XNOR2_X1 U7835 ( .A(n6373), .B(n6090), .ZN(n6113) );
  AOI21_X1 U7836 ( .B1(n6091), .B2(n5977), .A(n5715), .ZN(n6092) );
  NAND2_X1 U7837 ( .A1(n6096), .A2(n6093), .ZN(n6094) );
  NAND2_X1 U7838 ( .A1(n8250), .A2(n4412), .ZN(n6099) );
  INV_X1 U7839 ( .A(n6115), .ZN(n6097) );
  NAND2_X1 U7840 ( .A1(n6097), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6098) );
  NAND2_X1 U7841 ( .A1(n8420), .A2(n8425), .ZN(n6194) );
  NAND2_X1 U7842 ( .A1(n8743), .A2(n6101), .ZN(n8212) );
  INV_X1 U7843 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n10302) );
  NAND2_X1 U7844 ( .A1(n6061), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n6103) );
  NAND2_X1 U7845 ( .A1(n5796), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n6102) );
  OAI211_X1 U7846 ( .C1(n8208), .C2(n10302), .A(n6103), .B(n6102), .ZN(n6104)
         );
  INV_X1 U7847 ( .A(n6104), .ZN(n6105) );
  INV_X1 U7848 ( .A(n8190), .ZN(n8579) );
  INV_X4 U7849 ( .A(n8402), .ZN(n8406) );
  INV_X1 U7850 ( .A(n6290), .ZN(n8422) );
  BUF_X4 U7851 ( .A(n6106), .Z(n6107) );
  NAND2_X1 U7852 ( .A1(n8422), .A2(n6243), .ZN(n6108) );
  NAND2_X1 U7853 ( .A1(n5737), .A2(n6108), .ZN(n7212) );
  NAND2_X1 U7854 ( .A1(n8579), .A2(n8909), .ZN(n6111) );
  INV_X1 U7855 ( .A(n7212), .ZN(n6109) );
  NAND2_X1 U7856 ( .A1(n8768), .A2(n8907), .ZN(n6110) );
  AOI21_X1 U7857 ( .B1(n6113), .B2(n8912), .A(n6112), .ZN(n6367) );
  NAND2_X1 U7858 ( .A1(n6115), .A2(n6114), .ZN(n6116) );
  NAND2_X1 U7859 ( .A1(n6116), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6152) );
  NAND2_X1 U7860 ( .A1(n6152), .A2(n10253), .ZN(n6117) );
  XNOR2_X1 U7861 ( .A(n6129), .B(P2_B_REG_SCAN_IN), .ZN(n6122) );
  NAND2_X1 U7862 ( .A1(n6119), .A2(n6118), .ZN(n6120) );
  NAND2_X1 U7863 ( .A1(n6122), .A2(n6133), .ZN(n6128) );
  NAND2_X1 U7864 ( .A1(n6123), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6124) );
  MUX2_X1 U7865 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6124), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n6127) );
  INV_X1 U7866 ( .A(n6125), .ZN(n6126) );
  NAND2_X1 U7867 ( .A1(n6129), .A2(n8136), .ZN(n6959) );
  NAND2_X1 U7868 ( .A1(n6130), .A2(n6959), .ZN(n7204) );
  NAND3_X1 U7869 ( .A1(n4412), .A2(n8425), .A3(n7545), .ZN(n6131) );
  NAND2_X1 U7870 ( .A1(n8402), .A2(n6131), .ZN(n6136) );
  OR2_X1 U7871 ( .A1(n7204), .A2(n6136), .ZN(n6353) );
  NAND2_X1 U7872 ( .A1(n6195), .A2(n8420), .ZN(n6201) );
  NOR2_X1 U7873 ( .A1(n10000), .A2(n8250), .ZN(n6356) );
  NAND2_X1 U7874 ( .A1(n6133), .A2(n8136), .ZN(n6134) );
  INV_X1 U7875 ( .A(n6136), .ZN(n6137) );
  OAI21_X1 U7876 ( .B1(n6353), .B2(n6356), .A(n6354), .ZN(n6153) );
  INV_X1 U7877 ( .A(P2_D_REG_12__SCAN_IN), .ZN(n10060) );
  INV_X1 U7878 ( .A(P2_D_REG_18__SCAN_IN), .ZN(n10132) );
  INV_X1 U7879 ( .A(P2_D_REG_23__SCAN_IN), .ZN(n10145) );
  INV_X1 U7880 ( .A(P2_D_REG_17__SCAN_IN), .ZN(n10229) );
  NAND4_X1 U7881 ( .A1(n10060), .A2(n10132), .A3(n10145), .A4(n10229), .ZN(
        n10287) );
  INV_X1 U7882 ( .A(n10287), .ZN(n6140) );
  NOR2_X1 U7883 ( .A1(P2_D_REG_25__SCAN_IN), .A2(P2_D_REG_24__SCAN_IN), .ZN(
        n6139) );
  NOR4_X1 U7884 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_9__SCAN_IN), .A3(
        P2_D_REG_10__SCAN_IN), .A4(P2_D_REG_3__SCAN_IN), .ZN(n10353) );
  NOR4_X1 U7885 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_15__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n6138) );
  NAND4_X1 U7886 ( .A1(n6140), .A2(n6139), .A3(n10353), .A4(n6138), .ZN(n6146)
         );
  NOR4_X1 U7887 ( .A1(P2_D_REG_19__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_30__SCAN_IN), .ZN(n6144) );
  NOR4_X1 U7888 ( .A1(P2_D_REG_5__SCAN_IN), .A2(P2_D_REG_8__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_21__SCAN_IN), .ZN(n6143) );
  NOR4_X1 U7889 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_28__SCAN_IN), .A3(
        P2_D_REG_27__SCAN_IN), .A4(P2_D_REG_14__SCAN_IN), .ZN(n6142) );
  NOR4_X1 U7890 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_16__SCAN_IN), .A3(
        P2_D_REG_22__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n6141) );
  NAND4_X1 U7891 ( .A1(n6144), .A2(n6143), .A3(n6142), .A4(n6141), .ZN(n6145)
         );
  NOR2_X1 U7892 ( .A1(n6146), .A2(n6145), .ZN(n6147) );
  INV_X1 U7893 ( .A(n6133), .ZN(n6151) );
  INV_X1 U7894 ( .A(n6129), .ZN(n6149) );
  NAND2_X1 U7895 ( .A1(n6195), .A2(n7545), .ZN(n7198) );
  NAND2_X1 U7896 ( .A1(n6367), .A2(n10029), .ZN(n6156) );
  NAND2_X1 U7897 ( .A1(n10027), .A2(n6154), .ZN(n6155) );
  NAND2_X1 U7898 ( .A1(n6156), .A2(n6155), .ZN(n6185) );
  INV_X1 U7899 ( .A(n8268), .ZN(n9946) );
  NAND2_X1 U7900 ( .A1(n9941), .A2(n9946), .ZN(n9940) );
  NAND2_X1 U7901 ( .A1(n9940), .A2(n8260), .ZN(n7370) );
  INV_X1 U7902 ( .A(n7373), .ZN(n8219) );
  NAND2_X1 U7903 ( .A1(n7370), .A2(n8219), .ZN(n7371) );
  NAND2_X1 U7904 ( .A1(n7371), .A2(n8261), .ZN(n6160) );
  INV_X1 U7905 ( .A(n6157), .ZN(n6159) );
  NAND2_X1 U7906 ( .A1(n6160), .A2(n8270), .ZN(n7428) );
  INV_X1 U7907 ( .A(n7434), .ZN(n9978) );
  OR2_X1 U7908 ( .A1(n8592), .A2(n9978), .ZN(n8284) );
  INV_X1 U7909 ( .A(n7520), .ZN(n9984) );
  NAND2_X1 U7910 ( .A1(n8591), .A2(n9984), .ZN(n8287) );
  OR2_X1 U7911 ( .A1(n8591), .A2(n9984), .ZN(n8285) );
  OR2_X1 U7912 ( .A1(n8590), .A2(n9990), .ZN(n8248) );
  NAND2_X1 U7913 ( .A1(n8590), .A2(n9990), .ZN(n8246) );
  INV_X1 U7914 ( .A(n7553), .ZN(n8294) );
  NAND2_X1 U7915 ( .A1(n7554), .A2(n8294), .ZN(n6162) );
  NAND2_X1 U7916 ( .A1(n8589), .A2(n8304), .ZN(n8297) );
  NAND2_X1 U7917 ( .A1(n6162), .A2(n8297), .ZN(n7684) );
  INV_X1 U7918 ( .A(n8298), .ZN(n6163) );
  OR2_X1 U7919 ( .A1(n7996), .A2(n8006), .ZN(n8315) );
  NAND2_X1 U7920 ( .A1(n7996), .A2(n8006), .ZN(n8307) );
  AND2_X1 U7921 ( .A1(n8319), .A2(n8307), .ZN(n8313) );
  NAND2_X1 U7922 ( .A1(n6164), .A2(n8317), .ZN(n7878) );
  NAND2_X1 U7923 ( .A1(n10014), .A2(n8087), .ZN(n8324) );
  NAND2_X1 U7924 ( .A1(n7878), .A2(n7879), .ZN(n6165) );
  INV_X1 U7925 ( .A(n8584), .ZN(n8140) );
  NOR2_X1 U7926 ( .A1(n8096), .A2(n8140), .ZN(n8330) );
  NAND2_X1 U7927 ( .A1(n8096), .A2(n8140), .ZN(n8328) );
  OR2_X1 U7928 ( .A1(n8145), .A2(n8147), .ZN(n8334) );
  NAND2_X1 U7929 ( .A1(n8145), .A2(n8147), .ZN(n8335) );
  INV_X1 U7930 ( .A(n8894), .ZN(n8454) );
  AND2_X1 U7931 ( .A1(n9037), .A2(n8454), .ZN(n8216) );
  INV_X1 U7932 ( .A(n8350), .ZN(n6167) );
  INV_X1 U7933 ( .A(n8869), .ZN(n6169) );
  NAND2_X1 U7934 ( .A1(n8956), .A2(n8509), .ZN(n8343) );
  NAND2_X1 U7935 ( .A1(n8354), .A2(n8343), .ZN(n8870) );
  INV_X1 U7936 ( .A(n8870), .ZN(n6168) );
  NAND2_X1 U7937 ( .A1(n6169), .A2(n6168), .ZN(n8872) );
  NAND2_X1 U7938 ( .A1(n8872), .A2(n8354), .ZN(n8858) );
  AND2_X1 U7939 ( .A1(n8828), .A2(n8367), .ZN(n8363) );
  NAND2_X1 U7940 ( .A1(n6170), .A2(n8366), .ZN(n8815) );
  NAND2_X1 U7941 ( .A1(n8815), .A2(n8245), .ZN(n6171) );
  INV_X1 U7942 ( .A(n8380), .ZN(n6173) );
  NOR2_X1 U7943 ( .A1(n6173), .A2(n8786), .ZN(n6177) );
  OR2_X1 U7944 ( .A1(n8784), .A2(n6177), .ZN(n6174) );
  INV_X1 U7945 ( .A(n8379), .ZN(n6179) );
  OR2_X1 U7946 ( .A1(n6174), .A2(n6179), .ZN(n6175) );
  NAND2_X1 U7947 ( .A1(n8991), .A2(n8777), .ZN(n8376) );
  INV_X1 U7948 ( .A(n8819), .ZN(n8539) );
  AND2_X1 U7949 ( .A1(n8376), .A2(n8798), .ZN(n8785) );
  AND2_X1 U7950 ( .A1(n8785), .A2(n8380), .ZN(n6176) );
  OR2_X1 U7951 ( .A1(n6177), .A2(n6176), .ZN(n6178) );
  NOR2_X1 U7952 ( .A1(n8979), .A2(n8178), .ZN(n8383) );
  NAND2_X1 U7953 ( .A1(n8979), .A2(n8178), .ZN(n8214) );
  NAND2_X1 U7954 ( .A1(n6180), .A2(n8214), .ZN(n6186) );
  XOR2_X1 U7955 ( .A(n8235), .B(n6380), .Z(n6369) );
  AOI21_X1 U7956 ( .B1(n4412), .B2(n7848), .A(n8420), .ZN(n6181) );
  AND2_X1 U7957 ( .A1(n10005), .A2(n6181), .ZN(n6182) );
  NAND2_X1 U7958 ( .A1(n6185), .A2(n6184), .ZN(P2_U3487) );
  XOR2_X1 U7959 ( .A(n6186), .B(n8386), .Z(n8761) );
  XNOR2_X1 U7960 ( .A(n6187), .B(n8386), .ZN(n6191) );
  AOI21_X1 U7961 ( .B1(n8761), .B2(n9970), .A(n8756), .ZN(n6204) );
  MUX2_X1 U7962 ( .A(n6192), .B(n6204), .S(n10029), .Z(n6193) );
  NAND2_X1 U7963 ( .A1(n6193), .A2(n4983), .ZN(P2_U3486) );
  INV_X1 U7964 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n6205) );
  INV_X1 U7965 ( .A(n6194), .ZN(n6196) );
  NAND2_X1 U7966 ( .A1(n6196), .A2(n4412), .ZN(n6197) );
  OR2_X1 U7967 ( .A1(n8250), .A2(n6197), .ZN(n7116) );
  NAND2_X1 U7968 ( .A1(n7355), .A2(n7116), .ZN(n6198) );
  NAND2_X1 U7969 ( .A1(n7119), .A2(n6198), .ZN(n6203) );
  NAND2_X1 U7970 ( .A1(n7204), .A2(n6199), .ZN(n7095) );
  NAND3_X1 U7971 ( .A1(n7116), .A2(n8402), .A3(n10005), .ZN(n7114) );
  INV_X1 U7972 ( .A(n6201), .ZN(n6358) );
  OR2_X1 U7973 ( .A1(n7121), .A2(n7101), .ZN(n6202) );
  MUX2_X1 U7974 ( .A(n6205), .B(n6204), .S(n10016), .Z(n6206) );
  NAND2_X1 U7975 ( .A1(n6206), .A2(n4987), .ZN(P2_U3454) );
  INV_X1 U7976 ( .A(n8135), .ZN(n6207) );
  INV_X1 U7977 ( .A(n7097), .ZN(n7944) );
  OR2_X1 U7978 ( .A1(n8402), .A2(n7944), .ZN(n6208) );
  OR2_X1 U7979 ( .A1(n7098), .A2(n7944), .ZN(n6294) );
  NAND2_X1 U7980 ( .A1(n6208), .A2(n6294), .ZN(n6289) );
  OAI21_X1 U7981 ( .B1(n6289), .B2(n6209), .A(P2_STATE_REG_SCAN_IN), .ZN(
        P2_U3150) );
  XNOR2_X1 U7982 ( .A(n7545), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n6244) );
  INV_X1 U7983 ( .A(n8627), .ZN(n6953) );
  NOR2_X1 U7984 ( .A1(n6210), .A2(n9911), .ZN(n6211) );
  NAND2_X1 U7985 ( .A1(n5722), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6212) );
  NOR2_X1 U7986 ( .A1(n6974), .A2(n6256), .ZN(n6973) );
  INV_X1 U7987 ( .A(n6212), .ZN(n6213) );
  MUX2_X1 U7988 ( .A(n6214), .B(P2_REG1_REG_2__SCAN_IN), .S(n7021), .Z(n7026)
         );
  INV_X1 U7989 ( .A(n7054), .ZN(n6313) );
  AOI22_X1 U7990 ( .A1(P2_REG1_REG_4__SCAN_IN), .A2(n6316), .B1(n9937), .B2(
        n6217), .ZN(n9923) );
  NAND2_X1 U7991 ( .A1(P2_REG1_REG_6__SCAN_IN), .A2(n7237), .ZN(n6221) );
  OAI21_X1 U7992 ( .B1(P2_REG1_REG_6__SCAN_IN), .B2(n7237), .A(n6221), .ZN(
        n7239) );
  NAND2_X1 U7993 ( .A1(n6223), .A2(n7310), .ZN(n8600) );
  OAI21_X1 U7994 ( .B1(n6223), .B2(n7310), .A(n8600), .ZN(n7305) );
  INV_X1 U7995 ( .A(n7305), .ZN(n6224) );
  INV_X1 U7996 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n7306) );
  NAND2_X1 U7997 ( .A1(n6224), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n7304) );
  XNOR2_X1 U7998 ( .A(n6327), .B(P2_REG1_REG_8__SCAN_IN), .ZN(n8601) );
  INV_X1 U7999 ( .A(n8601), .ZN(n6225) );
  AOI21_X1 U8000 ( .B1(n7304), .B2(n8600), .A(n6225), .ZN(n8604) );
  INV_X1 U8001 ( .A(n6327), .ZN(n8598) );
  NOR2_X1 U8002 ( .A1(n6327), .A2(n6226), .ZN(n6227) );
  INV_X1 U8003 ( .A(n7655), .ZN(n6939) );
  NOR2_X1 U8004 ( .A1(n7655), .A2(n6229), .ZN(n6230) );
  NAND2_X1 U8005 ( .A1(P2_REG1_REG_10__SCAN_IN), .A2(n6943), .ZN(n6231) );
  OAI21_X1 U8006 ( .B1(P2_REG1_REG_10__SCAN_IN), .B2(n6943), .A(n6231), .ZN(
        n7761) );
  AOI22_X1 U8007 ( .A1(n8627), .A2(P2_REG1_REG_12__SCAN_IN), .B1(n5889), .B2(
        n6953), .ZN(n8616) );
  NOR2_X1 U8008 ( .A1(n8617), .A2(n8616), .ZN(n8615) );
  NOR2_X1 U8009 ( .A1(n8643), .A2(n6233), .ZN(n6234) );
  AOI22_X1 U8010 ( .A1(P2_REG1_REG_14__SCAN_IN), .A2(n8656), .B1(n7016), .B2(
        n6235), .ZN(n8651) );
  NOR2_X1 U8011 ( .A1(n8650), .A2(n4980), .ZN(n6236) );
  NOR2_X1 U8012 ( .A1(n8674), .A2(n6236), .ZN(n6237) );
  AOI22_X1 U8013 ( .A1(P2_REG1_REG_16__SCAN_IN), .A2(n8688), .B1(n7164), .B2(
        n8962), .ZN(n8692) );
  XNOR2_X1 U8014 ( .A(n6238), .B(n8708), .ZN(n8700) );
  INV_X1 U8015 ( .A(n8730), .ZN(n8731) );
  AOI22_X1 U8016 ( .A1(P2_REG1_REG_18__SCAN_IN), .A2(n8730), .B1(n8731), .B2(
        n10276), .ZN(n8722) );
  NOR2_X1 U8017 ( .A1(n8730), .A2(n10276), .ZN(n6239) );
  OAI21_X1 U8018 ( .B1(n8723), .B2(n6239), .A(n6244), .ZN(n6240) );
  OR2_X1 U8019 ( .A1(n6290), .A2(P2_U3151), .ZN(n8129) );
  NOR2_X1 U8020 ( .A1(n6289), .A2(n8129), .ZN(n9914) );
  OAI211_X1 U8021 ( .C1(n6244), .C2(n8723), .A(n6240), .B(n8737), .ZN(n6352)
         );
  AND2_X1 U8022 ( .A1(n9914), .A2(n6243), .ZN(n8608) );
  MUX2_X1 U8023 ( .A(n5985), .B(P2_REG2_REG_19__SCAN_IN), .S(n7545), .Z(n6349)
         );
  INV_X1 U8024 ( .A(n6349), .ZN(n6241) );
  NAND2_X1 U8025 ( .A1(n6241), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n6288) );
  INV_X1 U8026 ( .A(n6244), .ZN(n6242) );
  NAND3_X1 U8027 ( .A1(n8737), .A2(P2_REG1_REG_18__SCAN_IN), .A3(n6242), .ZN(
        n6287) );
  MUX2_X1 U8028 ( .A(n6244), .B(n6349), .S(n6243), .Z(n6306) );
  NAND2_X1 U8029 ( .A1(P2_U3893), .A2(n6290), .ZN(n7248) );
  MUX2_X1 U8030 ( .A(n8883), .B(n8959), .S(n6107), .Z(n6245) );
  NAND2_X1 U8031 ( .A1(n6245), .A2(n8708), .ZN(n6285) );
  XOR2_X1 U8032 ( .A(n8708), .B(n6245), .Z(n8703) );
  MUX2_X1 U8033 ( .A(P2_REG2_REG_16__SCAN_IN), .B(P2_REG1_REG_16__SCAN_IN), 
        .S(n6107), .Z(n6246) );
  OR2_X1 U8034 ( .A1(n6246), .A2(n7164), .ZN(n6284) );
  XNOR2_X1 U8035 ( .A(n6246), .B(n8688), .ZN(n8687) );
  MUX2_X1 U8036 ( .A(P2_REG2_REG_15__SCAN_IN), .B(P2_REG1_REG_15__SCAN_IN), 
        .S(n6107), .Z(n6248) );
  INV_X1 U8037 ( .A(n6248), .ZN(n6247) );
  NAND2_X1 U8038 ( .A1(n8674), .A2(n6247), .ZN(n6283) );
  XNOR2_X1 U8039 ( .A(n8674), .B(n6248), .ZN(n8670) );
  MUX2_X1 U8040 ( .A(P2_REG2_REG_14__SCAN_IN), .B(P2_REG1_REG_14__SCAN_IN), 
        .S(n6107), .Z(n6249) );
  OR2_X1 U8041 ( .A1(n6249), .A2(n7016), .ZN(n6282) );
  XNOR2_X1 U8042 ( .A(n8656), .B(n6249), .ZN(n8654) );
  MUX2_X1 U8043 ( .A(P2_REG2_REG_13__SCAN_IN), .B(P2_REG1_REG_13__SCAN_IN), 
        .S(n6107), .Z(n6251) );
  INV_X1 U8044 ( .A(n6251), .ZN(n6250) );
  NAND2_X1 U8045 ( .A1(n8643), .A2(n6250), .ZN(n6281) );
  XNOR2_X1 U8046 ( .A(n6251), .B(n8643), .ZN(n8637) );
  MUX2_X1 U8047 ( .A(P2_REG2_REG_12__SCAN_IN), .B(P2_REG1_REG_12__SCAN_IN), 
        .S(n6107), .Z(n6252) );
  OR2_X1 U8048 ( .A1(n6252), .A2(n6953), .ZN(n6280) );
  XNOR2_X1 U8049 ( .A(n6252), .B(n8627), .ZN(n8620) );
  MUX2_X1 U8050 ( .A(P2_REG2_REG_11__SCAN_IN), .B(P2_REG1_REG_11__SCAN_IN), 
        .S(n6107), .Z(n6253) );
  OR2_X1 U8051 ( .A1(n6253), .A2(n6948), .ZN(n6279) );
  XNOR2_X1 U8052 ( .A(n6253), .B(n7933), .ZN(n7928) );
  MUX2_X1 U8053 ( .A(P2_REG2_REG_10__SCAN_IN), .B(P2_REG1_REG_10__SCAN_IN), 
        .S(n6107), .Z(n6254) );
  OR2_X1 U8054 ( .A1(n6254), .A2(n6943), .ZN(n6278) );
  XNOR2_X1 U8055 ( .A(n6254), .B(n7766), .ZN(n7764) );
  MUX2_X1 U8056 ( .A(P2_REG2_REG_9__SCAN_IN), .B(P2_REG1_REG_9__SCAN_IN), .S(
        n6107), .Z(n6255) );
  OR2_X1 U8057 ( .A1(n6255), .A2(n6939), .ZN(n6277) );
  XNOR2_X1 U8058 ( .A(n6255), .B(n7655), .ZN(n7654) );
  MUX2_X1 U8059 ( .A(P2_REG2_REG_8__SCAN_IN), .B(P2_REG1_REG_8__SCAN_IN), .S(
        n6107), .Z(n6275) );
  OR2_X1 U8060 ( .A1(n6275), .A2(n8598), .ZN(n6276) );
  INV_X1 U8061 ( .A(n7237), .ZN(n6273) );
  MUX2_X1 U8062 ( .A(P2_REG2_REG_6__SCAN_IN), .B(P2_REG1_REG_6__SCAN_IN), .S(
        n6107), .Z(n6271) );
  INV_X1 U8063 ( .A(n6271), .ZN(n6272) );
  MUX2_X1 U8064 ( .A(P2_REG2_REG_5__SCAN_IN), .B(P2_REG1_REG_5__SCAN_IN), .S(
        n6107), .Z(n6269) );
  INV_X1 U8065 ( .A(n6269), .ZN(n6270) );
  MUX2_X1 U8066 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n6107), .Z(n6267) );
  INV_X1 U8067 ( .A(n6267), .ZN(n6268) );
  MUX2_X1 U8068 ( .A(n6257), .B(n6256), .S(n6107), .Z(n6258) );
  XNOR2_X1 U8069 ( .A(n6258), .B(n6977), .ZN(n6982) );
  MUX2_X1 U8070 ( .A(n7360), .B(n6210), .S(n6107), .Z(n9912) );
  NAND2_X1 U8071 ( .A1(n9912), .A2(n9911), .ZN(n6981) );
  NAND2_X1 U8072 ( .A1(n6982), .A2(n6981), .ZN(n6980) );
  INV_X1 U8073 ( .A(n6258), .ZN(n6259) );
  NAND2_X1 U8074 ( .A1(n6259), .A2(n6977), .ZN(n6260) );
  NAND2_X1 U8075 ( .A1(n6980), .A2(n6260), .ZN(n7034) );
  MUX2_X1 U8076 ( .A(P2_REG2_REG_2__SCAN_IN), .B(P2_REG1_REG_2__SCAN_IN), .S(
        n6107), .Z(n6262) );
  INV_X1 U8077 ( .A(n7021), .ZN(n6261) );
  XNOR2_X1 U8078 ( .A(n6262), .B(n6261), .ZN(n7033) );
  NAND2_X1 U8079 ( .A1(n7034), .A2(n7033), .ZN(n7032) );
  NAND2_X1 U8080 ( .A1(n6262), .A2(n7021), .ZN(n6263) );
  NAND2_X1 U8081 ( .A1(n7032), .A2(n6263), .ZN(n7051) );
  MUX2_X1 U8082 ( .A(P2_REG2_REG_3__SCAN_IN), .B(P2_REG1_REG_3__SCAN_IN), .S(
        n6107), .Z(n6264) );
  XNOR2_X1 U8083 ( .A(n6264), .B(n7054), .ZN(n7052) );
  OR2_X1 U8084 ( .A1(n7051), .A2(n7052), .ZN(n7049) );
  INV_X1 U8085 ( .A(n6264), .ZN(n6265) );
  NAND2_X1 U8086 ( .A1(n6265), .A2(n6313), .ZN(n6266) );
  AND2_X1 U8087 ( .A1(n7049), .A2(n6266), .ZN(n9921) );
  XNOR2_X1 U8088 ( .A(n6267), .B(n6316), .ZN(n9920) );
  NAND2_X1 U8089 ( .A1(n9921), .A2(n9920), .ZN(n9919) );
  OAI21_X1 U8090 ( .B1(n6316), .B2(n6268), .A(n9919), .ZN(n7137) );
  XNOR2_X1 U8091 ( .A(n6269), .B(n6320), .ZN(n7136) );
  NAND2_X1 U8092 ( .A1(n7137), .A2(n7136), .ZN(n7135) );
  OAI21_X1 U8093 ( .B1(n6320), .B2(n6270), .A(n7135), .ZN(n7235) );
  XNOR2_X1 U8094 ( .A(n6271), .B(n7237), .ZN(n7236) );
  NOR2_X1 U8095 ( .A1(n7235), .A2(n7236), .ZN(n7234) );
  AOI21_X1 U8096 ( .B1(n6273), .B2(n6272), .A(n7234), .ZN(n7308) );
  MUX2_X1 U8097 ( .A(P2_REG2_REG_7__SCAN_IN), .B(P2_REG1_REG_7__SCAN_IN), .S(
        n6107), .Z(n6274) );
  XNOR2_X1 U8098 ( .A(n6274), .B(n7310), .ZN(n7307) );
  OAI22_X1 U8099 ( .A1(n7308), .A2(n7307), .B1(n6274), .B2(n7310), .ZN(n8595)
         );
  XNOR2_X1 U8100 ( .A(n6275), .B(n6327), .ZN(n8594) );
  NAND2_X1 U8101 ( .A1(n8595), .A2(n8594), .ZN(n8593) );
  NAND2_X1 U8102 ( .A1(n6276), .A2(n8593), .ZN(n7653) );
  NAND2_X1 U8103 ( .A1(n7654), .A2(n7653), .ZN(n7652) );
  NAND2_X1 U8104 ( .A1(n6277), .A2(n7652), .ZN(n7763) );
  NAND2_X1 U8105 ( .A1(n7764), .A2(n7763), .ZN(n7762) );
  NAND2_X1 U8106 ( .A1(n6278), .A2(n7762), .ZN(n7927) );
  NAND2_X1 U8107 ( .A1(n7928), .A2(n7927), .ZN(n7926) );
  NAND2_X1 U8108 ( .A1(n6279), .A2(n7926), .ZN(n8619) );
  NAND2_X1 U8109 ( .A1(n8620), .A2(n8619), .ZN(n8618) );
  NAND2_X1 U8110 ( .A1(n6280), .A2(n8618), .ZN(n8636) );
  NAND2_X1 U8111 ( .A1(n8637), .A2(n8636), .ZN(n8635) );
  NAND2_X1 U8112 ( .A1(n6281), .A2(n8635), .ZN(n8653) );
  NAND2_X1 U8113 ( .A1(n8654), .A2(n8653), .ZN(n8652) );
  NAND2_X1 U8114 ( .A1(n6282), .A2(n8652), .ZN(n8669) );
  NAND2_X1 U8115 ( .A1(n8670), .A2(n8669), .ZN(n8668) );
  NAND2_X1 U8116 ( .A1(n6283), .A2(n8668), .ZN(n8686) );
  NAND2_X1 U8117 ( .A1(n8687), .A2(n8686), .ZN(n8685) );
  NAND2_X1 U8118 ( .A1(n6284), .A2(n8685), .ZN(n8702) );
  NAND2_X1 U8119 ( .A1(n8703), .A2(n8702), .ZN(n8701) );
  NAND2_X1 U8120 ( .A1(n6285), .A2(n8701), .ZN(n6300) );
  MUX2_X1 U8121 ( .A(n6345), .B(n10276), .S(n6107), .Z(n6301) );
  NAND2_X1 U8122 ( .A1(n6300), .A2(n6301), .ZN(n8725) );
  NAND3_X1 U8123 ( .A1(n6306), .A2(n9918), .A3(n8725), .ZN(n6286) );
  OAI211_X1 U8124 ( .C1(n9929), .C2(n6288), .A(n6287), .B(n6286), .ZN(n6309)
         );
  INV_X1 U8125 ( .A(n6289), .ZN(n6293) );
  NOR2_X1 U8126 ( .A1(n6107), .A2(P2_U3151), .ZN(n6291) );
  AND2_X1 U8127 ( .A1(n6291), .A2(n6290), .ZN(n6292) );
  NAND2_X1 U8128 ( .A1(n6293), .A2(n6292), .ZN(n6297) );
  INV_X1 U8129 ( .A(n6294), .ZN(n6298) );
  INV_X1 U8130 ( .A(n8129), .ZN(n6295) );
  NAND2_X1 U8131 ( .A1(n6298), .A2(n6295), .ZN(n6296) );
  INV_X1 U8132 ( .A(n8735), .ZN(n9934) );
  NAND2_X1 U8133 ( .A1(n9934), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n6299) );
  NAND2_X1 U8134 ( .A1(P2_U3151), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8472) );
  OAI211_X1 U8135 ( .C1(n9938), .C2(n7545), .A(n6299), .B(n8472), .ZN(n6308)
         );
  INV_X1 U8136 ( .A(n6300), .ZN(n6303) );
  INV_X1 U8137 ( .A(n6301), .ZN(n6302) );
  NAND2_X1 U8138 ( .A1(n6303), .A2(n6302), .ZN(n8726) );
  NAND2_X1 U8139 ( .A1(n8725), .A2(n8731), .ZN(n6304) );
  AOI21_X1 U8140 ( .B1(n6304), .B2(n8726), .A(n6306), .ZN(n6305) );
  AOI211_X1 U8141 ( .C1(n6306), .C2(n8726), .A(n7248), .B(n6305), .ZN(n6307)
         );
  AOI211_X1 U8142 ( .C1(n8731), .C2(n6309), .A(n6308), .B(n6307), .ZN(n6351)
         );
  NAND2_X1 U8143 ( .A1(n5722), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6310) );
  NOR2_X1 U8144 ( .A1(n6972), .A2(n6257), .ZN(n6971) );
  INV_X1 U8145 ( .A(n6310), .ZN(n6311) );
  NOR2_X1 U8146 ( .A1(n6971), .A2(n6311), .ZN(n7024) );
  OAI21_X1 U8147 ( .B1(n7021), .B2(P2_REG2_REG_2__SCAN_IN), .A(n6312), .ZN(
        n7023) );
  NOR2_X1 U8148 ( .A1(n7024), .A2(n7023), .ZN(n7022) );
  AOI21_X1 U8149 ( .B1(P2_REG2_REG_2__SCAN_IN), .B2(n7021), .A(n7022), .ZN(
        n6314) );
  INV_X1 U8150 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n7056) );
  AOI22_X1 U8151 ( .A1(P2_REG2_REG_4__SCAN_IN), .A2(n6316), .B1(n9937), .B2(
        n6317), .ZN(n9926) );
  NOR2_X1 U8152 ( .A1(n9927), .A2(n9926), .ZN(n9925) );
  NOR2_X1 U8153 ( .A1(n6316), .A2(n6317), .ZN(n6318) );
  NOR2_X1 U8154 ( .A1(n9925), .A2(n6318), .ZN(n6319) );
  XNOR2_X1 U8155 ( .A(n6319), .B(n6320), .ZN(n7130) );
  NOR2_X1 U8156 ( .A1(n6320), .A2(n6319), .ZN(n6321) );
  NAND2_X1 U8157 ( .A1(P2_REG2_REG_6__SCAN_IN), .A2(n7237), .ZN(n6322) );
  OAI21_X1 U8158 ( .B1(P2_REG2_REG_6__SCAN_IN), .B2(n7237), .A(n6322), .ZN(
        n7244) );
  INV_X1 U8159 ( .A(n7310), .ZN(n6324) );
  NAND2_X1 U8160 ( .A1(n6325), .A2(n6324), .ZN(n6326) );
  NAND2_X1 U8161 ( .A1(n8606), .A2(n6326), .ZN(n7312) );
  INV_X1 U8162 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7689) );
  XNOR2_X1 U8163 ( .A(n6327), .B(n7689), .ZN(n8607) );
  XNOR2_X1 U8164 ( .A(n6328), .B(n7655), .ZN(n7651) );
  NOR2_X1 U8165 ( .A1(n7655), .A2(n6328), .ZN(n6329) );
  NAND2_X1 U8166 ( .A1(P2_REG2_REG_10__SCAN_IN), .A2(n6943), .ZN(n6330) );
  OAI21_X1 U8167 ( .B1(n6943), .B2(P2_REG2_REG_10__SCAN_IN), .A(n6330), .ZN(
        n7770) );
  XNOR2_X1 U8168 ( .A(n6332), .B(n7933), .ZN(n7930) );
  NOR2_X1 U8169 ( .A1(n7930), .A2(n5867), .ZN(n7929) );
  INV_X1 U8170 ( .A(n6332), .ZN(n6333) );
  NOR2_X1 U8171 ( .A1(n7929), .A2(n6334), .ZN(n8623) );
  MUX2_X1 U8172 ( .A(P2_REG2_REG_12__SCAN_IN), .B(n6335), .S(n8627), .Z(n8622)
         );
  NOR2_X1 U8173 ( .A1(n8623), .A2(n8622), .ZN(n8621) );
  NOR2_X1 U8174 ( .A1(n8643), .A2(n6337), .ZN(n6338) );
  MUX2_X1 U8175 ( .A(P2_REG2_REG_14__SCAN_IN), .B(n6339), .S(n8656), .Z(n8659)
         );
  NOR2_X1 U8176 ( .A1(n8674), .A2(n6340), .ZN(n6341) );
  NAND2_X1 U8177 ( .A1(P2_REG2_REG_16__SCAN_IN), .A2(n7164), .ZN(n6342) );
  OAI21_X1 U8178 ( .B1(n7164), .B2(P2_REG2_REG_16__SCAN_IN), .A(n6342), .ZN(
        n8684) );
  NOR2_X1 U8179 ( .A1(n8708), .A2(n6343), .ZN(n6344) );
  XNOR2_X1 U8180 ( .A(n8708), .B(n6343), .ZN(n8705) );
  NOR2_X1 U8181 ( .A1(n8883), .A2(n8705), .ZN(n8707) );
  NOR2_X1 U8182 ( .A1(n8730), .A2(n6345), .ZN(n6347) );
  INV_X1 U8183 ( .A(n6347), .ZN(n6346) );
  OAI21_X1 U8184 ( .B1(P2_REG2_REG_18__SCAN_IN), .B2(n8731), .A(n6346), .ZN(
        n8720) );
  OAI21_X1 U8185 ( .B1(n8719), .B2(n6347), .A(n6349), .ZN(n6348) );
  OAI211_X1 U8186 ( .C1(n6349), .C2(n8719), .A(n6348), .B(n8608), .ZN(n6350)
         );
  NAND3_X1 U8187 ( .A1(n6352), .A2(n6351), .A3(n6350), .ZN(P2_U3201) );
  INV_X1 U8188 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n6357) );
  NAND4_X1 U8189 ( .A1(n6355), .A2(n7095), .A3(n6354), .A4(n6353), .ZN(n6361)
         );
  MUX2_X1 U8190 ( .A(n6357), .B(n6367), .S(n8913), .Z(n6366) );
  INV_X1 U8191 ( .A(n6369), .ZN(n6363) );
  OR2_X1 U8192 ( .A1(n9960), .A2(n9939), .ZN(n6360) );
  NAND2_X1 U8193 ( .A1(n6358), .A2(n8250), .ZN(n6359) );
  AOI22_X1 U8194 ( .A1(n8192), .A2(n8918), .B1(n8917), .B2(n8187), .ZN(n6362)
         );
  INV_X1 U8195 ( .A(n6364), .ZN(n6365) );
  NAND2_X1 U8196 ( .A1(n6366), .A2(n6365), .ZN(P2_U3205) );
  INV_X1 U8197 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n6368) );
  MUX2_X1 U8198 ( .A(n6368), .B(n6367), .S(n10016), .Z(n6372) );
  NAND2_X1 U8199 ( .A1(n6369), .A2(n9038), .ZN(n6370) );
  NAND2_X1 U8200 ( .A1(n6372), .A2(n6371), .ZN(P2_U3455) );
  NAND2_X1 U8201 ( .A1(n6373), .A2(n4997), .ZN(n6375) );
  NAND2_X1 U8202 ( .A1(n6375), .A2(n6374), .ZN(n6378) );
  OR2_X1 U8203 ( .A1(n9821), .A2(n5763), .ZN(n6377) );
  INV_X1 U8204 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n8430) );
  OR2_X1 U8205 ( .A1(n5764), .A2(n8430), .ZN(n6376) );
  NAND2_X1 U8206 ( .A1(n6395), .A2(n8190), .ZN(n8204) );
  XNOR2_X1 U8207 ( .A(n6378), .B(n8394), .ZN(n6379) );
  NAND2_X1 U8208 ( .A1(n6379), .A2(n8912), .ZN(n6391) );
  NAND2_X1 U8209 ( .A1(n6380), .A2(n8235), .ZN(n6382) );
  OR2_X1 U8210 ( .A1(n8192), .A2(n8443), .ZN(n6381) );
  INV_X1 U8211 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n8927) );
  NAND2_X1 U8212 ( .A1(n5796), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n6384) );
  NAND2_X1 U8213 ( .A1(n6061), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n6383) );
  OAI211_X1 U8214 ( .C1(n8927), .C2(n8208), .A(n6384), .B(n6383), .ZN(n6385)
         );
  INV_X1 U8215 ( .A(n6385), .ZN(n6386) );
  NAND2_X1 U8216 ( .A1(n8212), .A2(n6386), .ZN(n8578) );
  AND2_X1 U8217 ( .A1(n5737), .A2(P2_B_REG_SCAN_IN), .ZN(n6387) );
  NOR2_X1 U8218 ( .A1(n9953), .A2(n6387), .ZN(n8741) );
  AOI22_X1 U8219 ( .A1(n8907), .A2(n8580), .B1(n8578), .B2(n8741), .ZN(n6388)
         );
  INV_X1 U8220 ( .A(n6389), .ZN(n6390) );
  INV_X1 U8221 ( .A(n8755), .ZN(n6393) );
  INV_X1 U8222 ( .A(n10000), .ZN(n6392) );
  INV_X1 U8223 ( .A(n6395), .ZN(n6399) );
  NAND2_X1 U8224 ( .A1(n10017), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n6397) );
  OAI21_X1 U8225 ( .B1(n6402), .B2(n10017), .A(n4982), .ZN(P2_U3456) );
  OAI21_X1 U8226 ( .B1(n6402), .B2(n10027), .A(n6401), .ZN(P2_U3488) );
  INV_X2 U8227 ( .A(n6418), .ZN(n6508) );
  INV_X2 U8228 ( .A(n6448), .ZN(n6589) );
  AOI22_X1 U8229 ( .A1(n9696), .A2(n6587), .B1(n6448), .B2(n9545), .ZN(n6558)
         );
  INV_X1 U8230 ( .A(n6558), .ZN(n6560) );
  AND2_X1 U8231 ( .A1(n6406), .A2(n6405), .ZN(n6407) );
  AOI22_X1 U8232 ( .A1(n9696), .A2(n4416), .B1(n6508), .B2(n9545), .ZN(n6409)
         );
  XNOR2_X1 U8233 ( .A(n6409), .B(n6574), .ZN(n6557) );
  INV_X1 U8234 ( .A(n6557), .ZN(n6559) );
  XNOR2_X1 U8235 ( .A(n6410), .B(n6574), .ZN(n6438) );
  OR2_X1 U8236 ( .A1(n6411), .A2(n6590), .ZN(n6413) );
  OR2_X1 U8237 ( .A1(n6589), .A2(n7406), .ZN(n6412) );
  XNOR2_X1 U8238 ( .A(n6438), .B(n6437), .ZN(n7173) );
  NAND2_X1 U8239 ( .A1(n6428), .A2(n9879), .ZN(n6416) );
  INV_X1 U8240 ( .A(n6419), .ZN(n6414) );
  NAND2_X1 U8241 ( .A1(n6416), .A2(n6415), .ZN(n6423) );
  NOR2_X1 U8242 ( .A1(n6408), .A2(n6876), .ZN(n6417) );
  OR2_X1 U8243 ( .A1(n6423), .A2(n6417), .ZN(n6891) );
  INV_X1 U8244 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n6961) );
  OR2_X1 U8245 ( .A1(n6418), .A2(n7150), .ZN(n6422) );
  OR2_X1 U8246 ( .A1(n6420), .A2(n6419), .ZN(n6421) );
  OAI211_X1 U8247 ( .C1(n6408), .C2(n6961), .A(n6422), .B(n6421), .ZN(n6892)
         );
  NAND2_X1 U8248 ( .A1(n6891), .A2(n6892), .ZN(n6890) );
  INV_X1 U8249 ( .A(n6423), .ZN(n6425) );
  NAND2_X1 U8250 ( .A1(n6433), .A2(n6432), .ZN(n6435) );
  XNOR2_X1 U8251 ( .A(n6434), .B(n6435), .ZN(n9106) );
  NAND2_X1 U8252 ( .A1(n4999), .A2(n9106), .ZN(n9105) );
  INV_X1 U8253 ( .A(n6434), .ZN(n6436) );
  INV_X1 U8254 ( .A(n6437), .ZN(n6439) );
  OR2_X1 U8255 ( .A1(n6440), .A2(n6418), .ZN(n6442) );
  OR2_X1 U8256 ( .A1(n6589), .A2(n7086), .ZN(n6441) );
  NAND2_X1 U8257 ( .A1(n6442), .A2(n6441), .ZN(n6445) );
  XNOR2_X1 U8258 ( .A(n6443), .B(n6574), .ZN(n6444) );
  XOR2_X1 U8259 ( .A(n6445), .B(n6444), .Z(n7252) );
  INV_X1 U8260 ( .A(n6444), .ZN(n6446) );
  AOI22_X1 U8261 ( .A1(n9087), .A2(n7322), .B1(n6587), .B2(n9262), .ZN(n6447)
         );
  AOI22_X1 U8262 ( .A1(n6587), .A2(n7322), .B1(n6448), .B2(n9262), .ZN(n6450)
         );
  XNOR2_X1 U8263 ( .A(n6449), .B(n6450), .ZN(n7365) );
  INV_X1 U8264 ( .A(n6449), .ZN(n6452) );
  INV_X1 U8265 ( .A(n6450), .ZN(n6451) );
  AOI22_X1 U8266 ( .A1(n9087), .A2(n7493), .B1(n6587), .B2(n9261), .ZN(n6453)
         );
  OR2_X1 U8267 ( .A1(n9900), .A2(n6590), .ZN(n6455) );
  OR2_X1 U8268 ( .A1(n6589), .A2(n7614), .ZN(n6454) );
  NAND2_X1 U8269 ( .A1(n6455), .A2(n6454), .ZN(n7524) );
  AOI22_X1 U8270 ( .A1(n9087), .A2(n7616), .B1(n6508), .B2(n9260), .ZN(n6456)
         );
  XOR2_X1 U8271 ( .A(n6574), .B(n6456), .Z(n7611) );
  OR2_X1 U8272 ( .A1(n7387), .A2(n6590), .ZN(n6458) );
  OR2_X1 U8273 ( .A1(n6589), .A2(n7454), .ZN(n6457) );
  NAND2_X1 U8274 ( .A1(n6458), .A2(n6457), .ZN(n6459) );
  NOR2_X1 U8275 ( .A1(n7611), .A2(n6459), .ZN(n6461) );
  INV_X1 U8276 ( .A(n7611), .ZN(n6460) );
  INV_X1 U8277 ( .A(n6459), .ZN(n7610) );
  OAI22_X2 U8278 ( .A1(n7609), .A2(n6461), .B1(n6460), .B2(n7610), .ZN(n7624)
         );
  NAND2_X1 U8279 ( .A1(n9087), .A2(n7457), .ZN(n6463) );
  OR2_X1 U8280 ( .A1(n6590), .A2(n7841), .ZN(n6462) );
  NAND2_X1 U8281 ( .A1(n6463), .A2(n6462), .ZN(n6464) );
  XNOR2_X1 U8282 ( .A(n6464), .B(n9085), .ZN(n6468) );
  NAND2_X1 U8283 ( .A1(n6587), .A2(n7457), .ZN(n6466) );
  OR2_X1 U8284 ( .A1(n6589), .A2(n7841), .ZN(n6465) );
  AND2_X1 U8285 ( .A1(n6466), .A2(n6465), .ZN(n6467) );
  NAND2_X1 U8286 ( .A1(n6468), .A2(n6467), .ZN(n7620) );
  NOR2_X1 U8287 ( .A1(n6468), .A2(n6467), .ZN(n7622) );
  AOI22_X1 U8288 ( .A1(n9173), .A2(n9087), .B1(n6587), .B2(n9257), .ZN(n6469)
         );
  XOR2_X1 U8289 ( .A(n6574), .B(n6469), .Z(n9167) );
  NAND2_X1 U8290 ( .A1(n9173), .A2(n6587), .ZN(n6471) );
  OR2_X1 U8291 ( .A1(n6589), .A2(n7439), .ZN(n6470) );
  NAND2_X1 U8292 ( .A1(n6471), .A2(n6470), .ZN(n6477) );
  NAND2_X1 U8293 ( .A1(n7839), .A2(n6587), .ZN(n6473) );
  OR2_X1 U8294 ( .A1(n6589), .A2(n7588), .ZN(n6472) );
  NAND2_X1 U8295 ( .A1(n6473), .A2(n6472), .ZN(n7838) );
  NAND2_X1 U8296 ( .A1(n7839), .A2(n9087), .ZN(n6475) );
  OR2_X1 U8297 ( .A1(n6590), .A2(n7588), .ZN(n6474) );
  NAND2_X1 U8298 ( .A1(n6475), .A2(n6474), .ZN(n6476) );
  XNOR2_X1 U8299 ( .A(n6476), .B(n6574), .ZN(n6480) );
  AOI22_X1 U8300 ( .A1(n9167), .A2(n6477), .B1(n7838), .B2(n6480), .ZN(n6483)
         );
  INV_X1 U8301 ( .A(n6480), .ZN(n9165) );
  INV_X1 U8302 ( .A(n7838), .ZN(n6478) );
  INV_X1 U8303 ( .A(n6477), .ZN(n9166) );
  AOI21_X1 U8304 ( .B1(n9165), .B2(n6478), .A(n9166), .ZN(n6481) );
  NAND2_X1 U8305 ( .A1(n9166), .A2(n6478), .ZN(n6479) );
  OAI22_X1 U8306 ( .A1(n9167), .A2(n6481), .B1(n6480), .B2(n6479), .ZN(n6482)
         );
  AOI22_X1 U8307 ( .A1(n9210), .A2(n9087), .B1(n6508), .B2(n9255), .ZN(n6484)
         );
  XNOR2_X1 U8308 ( .A(n6484), .B(n6574), .ZN(n9202) );
  NOR2_X1 U8309 ( .A1(n6589), .A2(n7981), .ZN(n6485) );
  AOI21_X1 U8310 ( .B1(n9210), .B2(n6587), .A(n6485), .ZN(n9201) );
  NAND2_X1 U8311 ( .A1(n7756), .A2(n6587), .ZN(n6487) );
  OR2_X1 U8312 ( .A1(n6589), .A2(n7830), .ZN(n6486) );
  NAND2_X1 U8313 ( .A1(n6487), .A2(n6486), .ZN(n6491) );
  INV_X1 U8314 ( .A(n6491), .ZN(n7912) );
  NAND2_X1 U8315 ( .A1(n7756), .A2(n9087), .ZN(n6489) );
  OR2_X1 U8316 ( .A1(n6418), .A2(n7830), .ZN(n6488) );
  NAND2_X1 U8317 ( .A1(n6489), .A2(n6488), .ZN(n6490) );
  XNOR2_X1 U8318 ( .A(n6490), .B(n6574), .ZN(n9200) );
  INV_X1 U8319 ( .A(n9200), .ZN(n7910) );
  AOI22_X1 U8320 ( .A1(n9202), .A2(n9201), .B1(n7912), .B2(n7910), .ZN(n6496)
         );
  NAND2_X1 U8321 ( .A1(n9200), .A2(n6491), .ZN(n6493) );
  AOI21_X1 U8322 ( .B1(n9201), .B2(n6493), .A(n9202), .ZN(n6492) );
  INV_X1 U8323 ( .A(n6492), .ZN(n6494) );
  AOI21_X2 U8324 ( .B1(n7909), .B2(n6496), .A(n6495), .ZN(n7887) );
  AOI22_X1 U8325 ( .A1(n7889), .A2(n9087), .B1(n6508), .B2(n9254), .ZN(n6497)
         );
  XOR2_X1 U8326 ( .A(n6574), .B(n6497), .Z(n6499) );
  INV_X1 U8327 ( .A(n7889), .ZN(n7989) );
  OAI22_X1 U8328 ( .A1(n7989), .A2(n6418), .B1(n7962), .B2(n6589), .ZN(n6498)
         );
  NOR2_X1 U8329 ( .A1(n6499), .A2(n6498), .ZN(n6500) );
  AOI21_X1 U8330 ( .B1(n6499), .B2(n6498), .A(n6500), .ZN(n7886) );
  NAND2_X1 U8331 ( .A1(n7887), .A2(n7886), .ZN(n7885) );
  INV_X1 U8332 ( .A(n6500), .ZN(n6501) );
  NAND2_X1 U8333 ( .A1(n9744), .A2(n9087), .ZN(n6503) );
  OR2_X1 U8334 ( .A1(n6590), .A2(n8114), .ZN(n6502) );
  NAND2_X1 U8335 ( .A1(n6503), .A2(n6502), .ZN(n6504) );
  XNOR2_X1 U8336 ( .A(n6504), .B(n6574), .ZN(n6507) );
  AOI22_X1 U8337 ( .A1(n9744), .A2(n6587), .B1(n6448), .B2(n9253), .ZN(n6505)
         );
  XNOR2_X1 U8338 ( .A(n6507), .B(n6505), .ZN(n7971) );
  INV_X1 U8339 ( .A(n6505), .ZN(n6506) );
  AOI22_X1 U8340 ( .A1(n9059), .A2(n4416), .B1(n6508), .B2(n9252), .ZN(n6509)
         );
  XNOR2_X1 U8341 ( .A(n6509), .B(n6574), .ZN(n6512) );
  INV_X1 U8342 ( .A(n6512), .ZN(n6510) );
  NAND2_X1 U8343 ( .A1(n6511), .A2(n6510), .ZN(n6514) );
  NAND2_X1 U8344 ( .A1(n6513), .A2(n6512), .ZN(n6517) );
  INV_X1 U8345 ( .A(n9050), .ZN(n6516) );
  OAI22_X1 U8346 ( .A1(n8115), .A2(n6590), .B1(n9240), .B2(n6589), .ZN(n9053)
         );
  INV_X1 U8347 ( .A(n9053), .ZN(n6515) );
  AOI22_X1 U8348 ( .A1(n9739), .A2(n9087), .B1(n6587), .B2(n9624), .ZN(n6518)
         );
  XNOR2_X1 U8349 ( .A(n6518), .B(n6574), .ZN(n6519) );
  NAND2_X1 U8350 ( .A1(n6520), .A2(n6519), .ZN(n6521) );
  AOI22_X1 U8351 ( .A1(n9739), .A2(n6587), .B1(n6448), .B2(n9624), .ZN(n9234)
         );
  NAND2_X1 U8352 ( .A1(n9233), .A2(n6521), .ZN(n9127) );
  NOR2_X1 U8353 ( .A1(n6418), .A2(n9607), .ZN(n6522) );
  AOI21_X1 U8354 ( .B1(n9801), .B2(n9087), .A(n6522), .ZN(n6523) );
  XNOR2_X1 U8355 ( .A(n6523), .B(n6574), .ZN(n6528) );
  INV_X1 U8356 ( .A(n6528), .ZN(n6526) );
  NOR2_X1 U8357 ( .A1(n6589), .A2(n9607), .ZN(n6524) );
  AOI21_X1 U8358 ( .B1(n9801), .B2(n6587), .A(n6524), .ZN(n6527) );
  INV_X1 U8359 ( .A(n6527), .ZN(n6525) );
  NAND2_X1 U8360 ( .A1(n6526), .A2(n6525), .ZN(n9129) );
  AND2_X1 U8361 ( .A1(n6528), .A2(n6527), .ZN(n9128) );
  NAND2_X1 U8362 ( .A1(n9724), .A2(n4416), .ZN(n6530) );
  OR2_X1 U8363 ( .A1(n6590), .A2(n9592), .ZN(n6529) );
  NAND2_X1 U8364 ( .A1(n6530), .A2(n6529), .ZN(n6531) );
  XNOR2_X1 U8365 ( .A(n6531), .B(n9085), .ZN(n9139) );
  NOR2_X1 U8366 ( .A1(n6589), .A2(n9592), .ZN(n6532) );
  AOI21_X1 U8367 ( .B1(n9724), .B2(n6587), .A(n6532), .ZN(n6533) );
  INV_X1 U8368 ( .A(n6533), .ZN(n9138) );
  NAND2_X1 U8369 ( .A1(n9714), .A2(n9087), .ZN(n6535) );
  OR2_X1 U8370 ( .A1(n6418), .A2(n9706), .ZN(n6534) );
  NAND2_X1 U8371 ( .A1(n6535), .A2(n6534), .ZN(n6536) );
  XNOR2_X1 U8372 ( .A(n6536), .B(n6574), .ZN(n9075) );
  NAND2_X1 U8373 ( .A1(n9714), .A2(n6587), .ZN(n6538) );
  OR2_X1 U8374 ( .A1(n6589), .A2(n9706), .ZN(n6537) );
  NAND2_X1 U8375 ( .A1(n6538), .A2(n6537), .ZN(n9073) );
  NAND2_X1 U8376 ( .A1(n9075), .A2(n9073), .ZN(n9175) );
  INV_X1 U8377 ( .A(n9175), .ZN(n6545) );
  NAND2_X1 U8378 ( .A1(n9792), .A2(n4416), .ZN(n6540) );
  NAND2_X1 U8379 ( .A1(n6587), .A2(n9610), .ZN(n6539) );
  NAND2_X1 U8380 ( .A1(n6540), .A2(n6539), .ZN(n6541) );
  XNOR2_X1 U8381 ( .A(n6541), .B(n9085), .ZN(n9072) );
  NAND2_X1 U8382 ( .A1(n9792), .A2(n6587), .ZN(n6543) );
  NAND2_X1 U8383 ( .A1(n6448), .A2(n9610), .ZN(n6542) );
  NOR2_X1 U8384 ( .A1(n9072), .A2(n9214), .ZN(n6544) );
  INV_X1 U8385 ( .A(n9075), .ZN(n6551) );
  INV_X1 U8386 ( .A(n9072), .ZN(n9071) );
  INV_X1 U8387 ( .A(n9214), .ZN(n6547) );
  OAI21_X1 U8388 ( .B1(n9071), .B2(n6547), .A(n9073), .ZN(n6550) );
  NOR3_X1 U8389 ( .A1(n9071), .A2(n9073), .A3(n6547), .ZN(n6549) );
  AOI22_X1 U8390 ( .A1(n9703), .A2(n9087), .B1(n6587), .B2(n9695), .ZN(n6548)
         );
  XOR2_X1 U8391 ( .A(n6574), .B(n6548), .Z(n6552) );
  OAI22_X1 U8392 ( .A1(n9558), .A2(n6590), .B1(n9524), .B2(n6589), .ZN(n6553)
         );
  NOR2_X1 U8393 ( .A1(n6552), .A2(n6553), .ZN(n9178) );
  AOI211_X1 U8394 ( .C1(n6551), .C2(n6550), .A(n6549), .B(n9178), .ZN(n6556)
         );
  INV_X1 U8395 ( .A(n6552), .ZN(n6555) );
  INV_X1 U8396 ( .A(n6553), .ZN(n6554) );
  NOR2_X1 U8397 ( .A1(n6555), .A2(n6554), .ZN(n9177) );
  XOR2_X1 U8398 ( .A(n6558), .B(n6557), .Z(n9113) );
  NAND2_X1 U8399 ( .A1(n9112), .A2(n9113), .ZN(n9111) );
  AOI22_X1 U8400 ( .A1(n9509), .A2(n9087), .B1(n6587), .B2(n9532), .ZN(n6561)
         );
  XNOR2_X1 U8401 ( .A(n6561), .B(n6574), .ZN(n6562) );
  OAI22_X1 U8402 ( .A1(n9689), .A2(n6418), .B1(n9499), .B2(n6589), .ZN(n9187)
         );
  AOI22_X1 U8403 ( .A1(n9685), .A2(n9087), .B1(n6587), .B2(n9675), .ZN(n6564)
         );
  XNOR2_X1 U8404 ( .A(n6564), .B(n6574), .ZN(n6566) );
  AOI22_X1 U8405 ( .A1(n9685), .A2(n6587), .B1(n6448), .B2(n9675), .ZN(n6565)
         );
  NAND2_X1 U8406 ( .A1(n6566), .A2(n6565), .ZN(n9062) );
  AOI22_X1 U8407 ( .A1(n9676), .A2(n4416), .B1(n6587), .B2(n9469), .ZN(n6567)
         );
  XOR2_X1 U8408 ( .A(n6574), .B(n6567), .Z(n6569) );
  OAI22_X1 U8409 ( .A1(n4683), .A2(n6418), .B1(n9668), .B2(n6589), .ZN(n6568)
         );
  NOR2_X1 U8410 ( .A1(n6569), .A2(n6568), .ZN(n6570) );
  AOI21_X1 U8411 ( .B1(n6569), .B2(n6568), .A(n6570), .ZN(n9154) );
  NAND2_X1 U8412 ( .A1(n9153), .A2(n9154), .ZN(n9152) );
  INV_X1 U8413 ( .A(n6570), .ZN(n6571) );
  NAND2_X1 U8414 ( .A1(n9152), .A2(n6571), .ZN(n9120) );
  NAND2_X1 U8415 ( .A1(n9465), .A2(n4416), .ZN(n6573) );
  OR2_X1 U8416 ( .A1(n6590), .A2(n9478), .ZN(n6572) );
  NAND2_X1 U8417 ( .A1(n6573), .A2(n6572), .ZN(n6575) );
  XNOR2_X1 U8418 ( .A(n6575), .B(n6574), .ZN(n6580) );
  INV_X1 U8419 ( .A(n9478), .ZN(n9251) );
  AOI22_X1 U8420 ( .A1(n9465), .A2(n6587), .B1(n6448), .B2(n9251), .ZN(n6581)
         );
  XNOR2_X1 U8421 ( .A(n6580), .B(n6581), .ZN(n9121) );
  NAND2_X1 U8422 ( .A1(n9764), .A2(n4416), .ZN(n6577) );
  OR2_X1 U8423 ( .A1(n6590), .A2(n9657), .ZN(n6576) );
  NAND2_X1 U8424 ( .A1(n6577), .A2(n6576), .ZN(n6578) );
  XNOR2_X1 U8425 ( .A(n6578), .B(n6574), .ZN(n6586) );
  NOR2_X1 U8426 ( .A1(n6589), .A2(n9657), .ZN(n6579) );
  AOI21_X1 U8427 ( .B1(n9764), .B2(n6587), .A(n6579), .ZN(n6584) );
  XNOR2_X1 U8428 ( .A(n6586), .B(n6584), .ZN(n9223) );
  INV_X1 U8429 ( .A(n6580), .ZN(n6582) );
  NAND2_X1 U8430 ( .A1(n6582), .A2(n6581), .ZN(n9220) );
  INV_X1 U8431 ( .A(n6584), .ZN(n6585) );
  NAND2_X1 U8432 ( .A1(n6586), .A2(n6585), .ZN(n6594) );
  AOI22_X1 U8433 ( .A1(n9424), .A2(n9087), .B1(n6587), .B2(n9648), .ZN(n6588)
         );
  XOR2_X1 U8434 ( .A(n6574), .B(n6588), .Z(n6592) );
  OAI22_X1 U8435 ( .A1(n9658), .A2(n6590), .B1(n9441), .B2(n6589), .ZN(n6591)
         );
  NOR2_X1 U8436 ( .A1(n6592), .A2(n6591), .ZN(n9098) );
  AOI21_X1 U8437 ( .B1(n6592), .B2(n6591), .A(n9098), .ZN(n6593) );
  AOI21_X1 U8438 ( .B1(n9222), .B2(n6594), .A(n6593), .ZN(n6603) );
  INV_X1 U8439 ( .A(n6593), .ZN(n6596) );
  INV_X1 U8440 ( .A(n6594), .ZN(n6595) );
  NOR2_X1 U8441 ( .A1(n6596), .A2(n6595), .ZN(n6597) );
  NAND2_X1 U8442 ( .A1(n9899), .A2(n9876), .ZN(n6601) );
  NOR2_X1 U8443 ( .A1(n9807), .A2(n6601), .ZN(n6602) );
  OAI21_X1 U8444 ( .B1(n6603), .B2(n9093), .A(n9236), .ZN(n6620) );
  INV_X1 U8445 ( .A(n6604), .ZN(n9425) );
  INV_X1 U8446 ( .A(n6617), .ZN(n6606) );
  NAND2_X1 U8447 ( .A1(n6606), .A2(n6605), .ZN(n6609) );
  INV_X1 U8448 ( .A(n6679), .ZN(n6872) );
  NOR2_X1 U8449 ( .A1(n6607), .A2(n6872), .ZN(n6608) );
  NAND2_X1 U8450 ( .A1(n6609), .A2(n6608), .ZN(n9142) );
  NOR2_X1 U8451 ( .A1(n9807), .A2(n6842), .ZN(n6610) );
  AND2_X1 U8452 ( .A1(n6617), .A2(n6610), .ZN(n6612) );
  INV_X1 U8453 ( .A(n6612), .ZN(n6611) );
  AOI22_X1 U8454 ( .A1(n9225), .A2(n5524), .B1(P1_REG3_REG_27__SCAN_IN), .B2(
        P1_U3086), .ZN(n6613) );
  OAI21_X1 U8455 ( .B1(n9432), .B2(n9227), .A(n6613), .ZN(n6614) );
  AOI21_X1 U8456 ( .B1(n9425), .B2(n9229), .A(n6614), .ZN(n6619) );
  NOR2_X1 U8457 ( .A1(n9807), .A2(n6615), .ZN(n6616) );
  NAND2_X1 U8458 ( .A1(n6617), .A2(n6616), .ZN(n6618) );
  NAND3_X1 U8459 ( .A1(n6620), .A2(n6619), .A3(n4988), .ZN(P1_U3214) );
  INV_X1 U8460 ( .A(n6621), .ZN(n6622) );
  MUX2_X1 U8461 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(P2_DATAO_REG_30__SCAN_IN), 
        .S(n6915), .Z(n6628) );
  XNOR2_X1 U8462 ( .A(n6628), .B(SI_30_), .ZN(n6629) );
  NAND2_X1 U8463 ( .A1(n8429), .A2(n6635), .ZN(n6627) );
  INV_X1 U8464 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n10303) );
  OR2_X1 U8465 ( .A1(n5155), .A2(n10303), .ZN(n6626) );
  INV_X1 U8466 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n6631) );
  INV_X1 U8467 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n6636) );
  MUX2_X1 U8468 ( .A(n6631), .B(n6636), .S(n6915), .Z(n6632) );
  XNOR2_X1 U8469 ( .A(n6632), .B(SI_31_), .ZN(n6633) );
  NAND2_X1 U8470 ( .A1(n9812), .A2(n6635), .ZN(n6638) );
  OR2_X1 U8471 ( .A1(n5155), .A2(n6636), .ZN(n6637) );
  INV_X1 U8472 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n6642) );
  INV_X1 U8473 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n9639) );
  OR2_X1 U8474 ( .A1(n4413), .A2(n9639), .ZN(n6641) );
  NAND2_X1 U8475 ( .A1(n6639), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n6640) );
  OAI211_X1 U8476 ( .C1(n5649), .C2(n6642), .A(n6641), .B(n6640), .ZN(n9394)
         );
  AND2_X1 U8477 ( .A1(n6743), .A2(n7812), .ZN(n6752) );
  OR2_X1 U8478 ( .A1(n9879), .A2(n6419), .ZN(n6688) );
  OAI211_X1 U8479 ( .C1(n7087), .C2(n4417), .A(n6688), .B(n4418), .ZN(n6643)
         );
  INV_X1 U8480 ( .A(n6643), .ZN(n6644) );
  OAI211_X1 U8481 ( .C1(n6712), .C2(n6644), .A(n5627), .B(n6721), .ZN(n6645)
         );
  INV_X1 U8482 ( .A(n6722), .ZN(n7222) );
  AOI21_X1 U8483 ( .B1(n6645), .B2(n6713), .A(n7222), .ZN(n6646) );
  NAND2_X1 U8484 ( .A1(n6714), .A2(n6717), .ZN(n6724) );
  OAI21_X1 U8485 ( .B1(n6646), .B2(n6724), .A(n6719), .ZN(n6647) );
  NAND2_X1 U8486 ( .A1(n6694), .A2(n6647), .ZN(n6648) );
  NAND3_X1 U8487 ( .A1(n6648), .A2(n6754), .A3(n7738), .ZN(n6649) );
  NAND2_X1 U8488 ( .A1(n7956), .A2(n6741), .ZN(n6757) );
  AOI21_X1 U8489 ( .B1(n6752), .B2(n6649), .A(n6757), .ZN(n6651) );
  NAND2_X1 U8490 ( .A1(n8100), .A2(n6756), .ZN(n6650) );
  OAI211_X1 U8491 ( .C1(n6651), .C2(n6650), .A(n6761), .B(n6759), .ZN(n6652)
         );
  INV_X1 U8492 ( .A(n6652), .ZN(n6654) );
  NAND2_X1 U8493 ( .A1(n6766), .A2(n6653), .ZN(n6747) );
  OAI211_X1 U8494 ( .C1(n6654), .C2(n6747), .A(n6767), .B(n6762), .ZN(n6657)
         );
  NAND2_X1 U8495 ( .A1(n6656), .A2(n6655), .ZN(n6686) );
  NAND2_X1 U8496 ( .A1(n6779), .A2(n6656), .ZN(n6784) );
  AOI211_X1 U8497 ( .C1(n6770), .C2(n6657), .A(n6686), .B(n6784), .ZN(n6663)
         );
  NAND2_X1 U8498 ( .A1(n9724), .A2(n9592), .ZN(n6658) );
  AND2_X1 U8499 ( .A1(n6776), .A2(n6658), .ZN(n6685) );
  OAI21_X1 U8500 ( .B1(n6784), .B2(n6685), .A(n6777), .ZN(n6781) );
  NAND2_X1 U8501 ( .A1(n6801), .A2(n6659), .ZN(n6793) );
  INV_X1 U8502 ( .A(n6795), .ZN(n6660) );
  AOI21_X1 U8503 ( .B1(n6666), .B2(n6793), .A(n6660), .ZN(n6662) );
  INV_X1 U8504 ( .A(n6804), .ZN(n6661) );
  OAI21_X1 U8505 ( .B1(n6662), .B2(n6661), .A(n9437), .ZN(n6664) );
  NOR2_X1 U8506 ( .A1(n6664), .A2(n6707), .ZN(n6844) );
  OAI21_X1 U8507 ( .B1(n6663), .B2(n6781), .A(n6844), .ZN(n6672) );
  INV_X1 U8508 ( .A(n6664), .ZN(n6671) );
  AND2_X1 U8509 ( .A1(n6666), .A2(n6665), .ZN(n6799) );
  NAND3_X1 U8510 ( .A1(n6804), .A2(n6799), .A3(n6667), .ZN(n6670) );
  NAND2_X1 U8511 ( .A1(n6669), .A2(n6668), .ZN(n6812) );
  AOI21_X1 U8512 ( .B1(n6671), .B2(n6670), .A(n6812), .ZN(n6845) );
  NAND2_X1 U8513 ( .A1(n6819), .A2(n6811), .ZN(n6847) );
  AOI21_X1 U8514 ( .B1(n6672), .B2(n6845), .A(n6847), .ZN(n6674) );
  NOR2_X1 U8515 ( .A1(n6674), .A2(n6848), .ZN(n6676) );
  INV_X1 U8516 ( .A(n9410), .ZN(n6675) );
  OAI21_X1 U8517 ( .B1(n6821), .B2(n6675), .A(n6818), .ZN(n6852) );
  NOR2_X1 U8518 ( .A1(n9756), .A2(n9249), .ZN(n6705) );
  AOI21_X1 U8519 ( .B1(n6675), .B2(n6821), .A(n6705), .ZN(n6853) );
  OAI21_X1 U8520 ( .B1(n6676), .B2(n6852), .A(n6853), .ZN(n6677) );
  AOI21_X1 U8521 ( .B1(n6684), .B2(n6677), .A(n6839), .ZN(n6682) );
  OR2_X1 U8522 ( .A1(n6678), .A2(n4519), .ZN(n9880) );
  OR2_X1 U8523 ( .A1(n6679), .A2(P1_U3086), .ZN(n7941) );
  NOR2_X1 U8524 ( .A1(n6682), .A2(n6680), .ZN(n6681) );
  AOI211_X1 U8525 ( .C1(n6682), .C2(n9880), .A(n7941), .B(n6681), .ZN(n6683)
         );
  INV_X1 U8526 ( .A(n6683), .ZN(n6870) );
  INV_X1 U8527 ( .A(n6684), .ZN(n6706) );
  INV_X1 U8528 ( .A(n9411), .ZN(n6703) );
  INV_X1 U8529 ( .A(n9496), .ZN(n6700) );
  XNOR2_X1 U8530 ( .A(n9703), .B(n9524), .ZN(n9526) );
  INV_X1 U8531 ( .A(n6685), .ZN(n6698) );
  INV_X1 U8532 ( .A(n6686), .ZN(n6775) );
  INV_X1 U8533 ( .A(n7817), .ZN(n7813) );
  INV_X1 U8534 ( .A(n6687), .ZN(n7090) );
  INV_X1 U8535 ( .A(n6688), .ZN(n6689) );
  OR2_X1 U8536 ( .A1(n7151), .A2(n6689), .ZN(n9892) );
  NOR4_X1 U8537 ( .A1(n6687), .A2(n9892), .A3(n7180), .A4(n4418), .ZN(n6690)
         );
  INV_X1 U8538 ( .A(n7219), .ZN(n7224) );
  NAND4_X1 U8539 ( .A1(n6690), .A2(n7498), .A3(n7224), .A4(n7152), .ZN(n6691)
         );
  NOR3_X1 U8540 ( .A1(n7736), .A2(n6692), .A3(n6691), .ZN(n6693) );
  NAND4_X1 U8541 ( .A1(n7856), .A2(n7813), .A3(n6694), .A4(n6693), .ZN(n6695)
         );
  NOR4_X1 U8542 ( .A1(n8053), .A2(n8102), .A3(n7960), .A4(n6695), .ZN(n6696)
         );
  NAND3_X1 U8543 ( .A1(n6775), .A2(n9623), .A3(n6696), .ZN(n6697) );
  NOR4_X1 U8544 ( .A1(n9526), .A2(n9564), .A3(n6698), .A4(n6697), .ZN(n6699)
         );
  NAND4_X1 U8545 ( .A1(n6700), .A2(n9517), .A3(n9528), .A4(n6699), .ZN(n6701)
         );
  NOR4_X1 U8546 ( .A1(n9444), .A2(n9457), .A3(n6800), .A4(n6701), .ZN(n6702)
         );
  NAND4_X1 U8547 ( .A1(n6824), .A2(n6703), .A3(n4457), .A4(n6702), .ZN(n6704)
         );
  INV_X1 U8548 ( .A(n6861), .ZN(n6835) );
  INV_X1 U8549 ( .A(n6848), .ZN(n6807) );
  NAND2_X1 U8550 ( .A1(n6811), .A2(n9437), .ZN(n6808) );
  NOR2_X1 U8551 ( .A1(n6808), .A2(n6812), .ZN(n6806) );
  MUX2_X1 U8552 ( .A(n6708), .B(n6707), .S(n6825), .Z(n6791) );
  AOI21_X1 U8553 ( .B1(n7084), .B2(n5627), .A(n6709), .ZN(n6710) );
  MUX2_X1 U8554 ( .A(n5627), .B(n6710), .S(n6825), .Z(n6711) );
  NAND2_X1 U8555 ( .A1(n6711), .A2(n7184), .ZN(n6730) );
  INV_X1 U8556 ( .A(n6712), .ZN(n6715) );
  OAI211_X1 U8557 ( .C1(n6730), .C2(n6715), .A(n6714), .B(n6713), .ZN(n6716)
         );
  NAND2_X1 U8558 ( .A1(n6716), .A2(n6722), .ZN(n6718) );
  NAND4_X1 U8559 ( .A1(n6718), .A2(n6837), .A3(n7418), .A4(n6717), .ZN(n6732)
         );
  NAND2_X1 U8560 ( .A1(n6720), .A2(n6719), .ZN(n7419) );
  NAND3_X1 U8561 ( .A1(n6722), .A2(n6721), .A3(n6825), .ZN(n6723) );
  NOR2_X1 U8562 ( .A1(n7419), .A2(n6723), .ZN(n6729) );
  NAND2_X1 U8563 ( .A1(n6724), .A2(n6825), .ZN(n6727) );
  NAND3_X1 U8564 ( .A1(n7419), .A2(n6837), .A3(n7418), .ZN(n6726) );
  OR2_X1 U8565 ( .A1(n7418), .A2(n6837), .ZN(n6725) );
  OAI211_X1 U8566 ( .C1(n7419), .C2(n6727), .A(n6726), .B(n6725), .ZN(n6728)
         );
  AOI21_X1 U8567 ( .B1(n6730), .B2(n6729), .A(n6728), .ZN(n6731) );
  NAND2_X1 U8568 ( .A1(n6732), .A2(n6731), .ZN(n6733) );
  INV_X1 U8569 ( .A(n7413), .ZN(n7422) );
  AND2_X1 U8570 ( .A1(n7583), .A2(n6735), .ZN(n6738) );
  NAND2_X1 U8571 ( .A1(n6751), .A2(n6736), .ZN(n6737) );
  INV_X1 U8572 ( .A(n6739), .ZN(n6740) );
  NAND3_X1 U8573 ( .A1(n6742), .A2(n6754), .A3(n6741), .ZN(n6744) );
  INV_X1 U8574 ( .A(n6759), .ZN(n6746) );
  INV_X1 U8575 ( .A(n6747), .ZN(n6749) );
  INV_X1 U8576 ( .A(n6762), .ZN(n6748) );
  OAI21_X1 U8577 ( .B1(n6750), .B2(n4714), .A(n6767), .ZN(n6773) );
  NAND2_X1 U8578 ( .A1(n4474), .A2(n6751), .ZN(n6755) );
  INV_X1 U8579 ( .A(n6752), .ZN(n6753) );
  AOI21_X1 U8580 ( .B1(n6755), .B2(n6754), .A(n6753), .ZN(n6758) );
  OAI21_X1 U8581 ( .B1(n6758), .B2(n6757), .A(n6756), .ZN(n6760) );
  NAND2_X1 U8582 ( .A1(n6760), .A2(n6759), .ZN(n6765) );
  NAND2_X1 U8583 ( .A1(n6762), .A2(n6761), .ZN(n6763) );
  AOI21_X1 U8584 ( .B1(n6765), .B2(n6764), .A(n6763), .ZN(n6769) );
  INV_X1 U8585 ( .A(n6766), .ZN(n6768) );
  OAI21_X1 U8586 ( .B1(n6769), .B2(n6768), .A(n6767), .ZN(n6771) );
  NAND2_X1 U8587 ( .A1(n6771), .A2(n6770), .ZN(n6772) );
  INV_X1 U8588 ( .A(n6774), .ZN(n9608) );
  NAND2_X1 U8589 ( .A1(n6785), .A2(n6775), .ZN(n6778) );
  NAND3_X1 U8590 ( .A1(n6778), .A2(n6777), .A3(n6776), .ZN(n6780) );
  NAND3_X1 U8591 ( .A1(n6780), .A2(n9527), .A3(n6779), .ZN(n6786) );
  INV_X1 U8592 ( .A(n6781), .ZN(n6783) );
  OAI21_X1 U8593 ( .B1(n6786), .B2(n6825), .A(n4604), .ZN(n6790) );
  MUX2_X1 U8594 ( .A(n6788), .B(n6787), .S(n6837), .Z(n6789) );
  NAND2_X1 U8595 ( .A1(n6792), .A2(n9517), .ZN(n6798) );
  INV_X1 U8596 ( .A(n6793), .ZN(n6794) );
  AND2_X1 U8597 ( .A1(n6798), .A2(n6794), .ZN(n6796) );
  OAI21_X1 U8598 ( .B1(n6797), .B2(n6796), .A(n6795), .ZN(n6805) );
  INV_X1 U8599 ( .A(n6798), .ZN(n6803) );
  INV_X1 U8600 ( .A(n6799), .ZN(n6802) );
  AND2_X1 U8601 ( .A1(n6812), .A2(n6811), .ZN(n6810) );
  INV_X1 U8602 ( .A(n6808), .ZN(n6809) );
  NAND2_X1 U8603 ( .A1(n6848), .A2(n6825), .ZN(n6814) );
  NAND4_X1 U8604 ( .A1(n6819), .A2(n6825), .A3(n6812), .A4(n6811), .ZN(n6813)
         );
  NAND4_X1 U8605 ( .A1(n6816), .A2(n6815), .A3(n6814), .A4(n6813), .ZN(n6817)
         );
  OAI21_X1 U8606 ( .B1(n6848), .B2(n6819), .A(n6818), .ZN(n6820) );
  NAND2_X1 U8607 ( .A1(n6821), .A2(n9410), .ZN(n6823) );
  MUX2_X1 U8608 ( .A(n9410), .B(n6821), .S(n6825), .Z(n6822) );
  INV_X1 U8609 ( .A(n9752), .ZN(n6826) );
  NAND3_X1 U8610 ( .A1(n6827), .A2(n9249), .A3(n6826), .ZN(n6832) );
  NAND2_X1 U8611 ( .A1(n9249), .A2(n9394), .ZN(n6854) );
  INV_X1 U8612 ( .A(n6839), .ZN(n6859) );
  NAND3_X1 U8613 ( .A1(n6829), .A2(n6854), .A3(n6859), .ZN(n6831) );
  INV_X1 U8614 ( .A(n6857), .ZN(n6830) );
  AOI21_X1 U8615 ( .B1(n6836), .B2(n6843), .A(n7732), .ZN(n6833) );
  INV_X1 U8616 ( .A(n6833), .ZN(n6834) );
  NOR2_X1 U8617 ( .A1(n7941), .A2(n7667), .ZN(n6860) );
  NAND4_X1 U8618 ( .A1(n6835), .A2(n6834), .A3(n5666), .A4(n6860), .ZN(n6869)
         );
  NAND3_X1 U8619 ( .A1(n6860), .A2(n4418), .A3(n7849), .ZN(n6838) );
  NOR4_X1 U8620 ( .A1(n9807), .A2(n9705), .A3(n8195), .A4(n6842), .ZN(n6865)
         );
  OAI21_X1 U8621 ( .B1(n7941), .B2(n6843), .A(P1_B_REG_SCAN_IN), .ZN(n6864) );
  INV_X1 U8622 ( .A(n6844), .ZN(n6846) );
  OAI21_X1 U8623 ( .B1(n9544), .B2(n6846), .A(n6845), .ZN(n6850) );
  INV_X1 U8624 ( .A(n6847), .ZN(n6849) );
  AOI21_X1 U8625 ( .B1(n6850), .B2(n6849), .A(n6848), .ZN(n6851) );
  OAI22_X1 U8626 ( .A1(n9756), .A2(n9394), .B1(n6852), .B2(n6851), .ZN(n6856)
         );
  INV_X1 U8627 ( .A(n6853), .ZN(n6855) );
  OAI22_X1 U8628 ( .A1(n6856), .A2(n6855), .B1(n9401), .B2(n6854), .ZN(n6858)
         );
  AOI211_X1 U8629 ( .C1(n6859), .C2(n6858), .A(n9876), .B(n6857), .ZN(n6862)
         );
  OAI211_X1 U8630 ( .C1(n6862), .C2(n6861), .A(n6860), .B(n4519), .ZN(n6863)
         );
  OAI21_X1 U8631 ( .B1(n6865), .B2(n6864), .A(n6863), .ZN(n6866) );
  INV_X1 U8632 ( .A(n6866), .ZN(n6867) );
  NAND4_X1 U8633 ( .A1(n6870), .A2(n6869), .A3(n6868), .A4(n6867), .ZN(
        P1_U3242) );
  OR2_X2 U8634 ( .A1(n6408), .A2(n6871), .ZN(n10054) );
  NAND2_X1 U8635 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n6893) );
  NOR2_X1 U8636 ( .A1(n6875), .A2(n6893), .ZN(n6901) );
  NAND2_X1 U8637 ( .A1(n9807), .A2(n7941), .ZN(n6884) );
  OR2_X1 U8638 ( .A1(n9876), .A2(n6872), .ZN(n6874) );
  AND2_X1 U8639 ( .A1(n6874), .A2(n6873), .ZN(n6882) );
  NAND2_X1 U8640 ( .A1(n6884), .A2(n6882), .ZN(n6881) );
  AOI211_X1 U8641 ( .C1(n6893), .C2(n6875), .A(n6901), .B(n9844), .ZN(n6889)
         );
  INV_X1 U8642 ( .A(n6881), .ZN(n6965) );
  MUX2_X1 U8643 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n6878), .S(n6916), .Z(n6877)
         );
  NOR3_X1 U8644 ( .A1(n6877), .A2(n6876), .A3(n6961), .ZN(n6904) );
  MUX2_X1 U8645 ( .A(n6878), .B(P1_REG1_REG_1__SCAN_IN), .S(n6916), .Z(n6879)
         );
  AOI21_X1 U8646 ( .B1(P1_IR_REG_0__SCAN_IN), .B2(P1_REG1_REG_0__SCAN_IN), .A(
        n6879), .ZN(n6880) );
  NOR3_X1 U8647 ( .A1(n9869), .A2(n6904), .A3(n6880), .ZN(n6888) );
  NOR2_X1 U8648 ( .A1(n9866), .A2(n6916), .ZN(n6887) );
  INV_X1 U8649 ( .A(n6882), .ZN(n6883) );
  NAND2_X1 U8650 ( .A1(n6884), .A2(n6883), .ZN(n9875) );
  INV_X1 U8651 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n6885) );
  OAI22_X1 U8652 ( .A1(n9875), .A2(n6885), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n7394), .ZN(n6886) );
  OR4_X1 U8653 ( .A1(n6889), .A2(n6888), .A3(n6887), .A4(n6886), .ZN(P1_U3244)
         );
  OAI21_X1 U8654 ( .B1(n6892), .B2(n6891), .A(n6890), .ZN(n7141) );
  INV_X1 U8655 ( .A(n6893), .ZN(n6895) );
  INV_X1 U8656 ( .A(n8195), .ZN(n6894) );
  MUX2_X1 U8657 ( .A(n7141), .B(n6895), .S(n6894), .Z(n6900) );
  OR2_X1 U8658 ( .A1(n8195), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n6896) );
  NAND2_X1 U8659 ( .A1(n6899), .A2(n6896), .ZN(n6963) );
  AND2_X1 U8660 ( .A1(n6963), .A2(n6961), .ZN(n6897) );
  OR2_X1 U8661 ( .A1(n10054), .A2(n6897), .ZN(n6898) );
  AOI21_X1 U8662 ( .B1(n6900), .B2(n6899), .A(n6898), .ZN(n9855) );
  AOI21_X1 U8663 ( .B1(P1_REG2_REG_1__SCAN_IN), .B2(n6905), .A(n6901), .ZN(
        n6903) );
  INV_X1 U8664 ( .A(n6922), .ZN(n6994) );
  XNOR2_X1 U8665 ( .A(n6994), .B(P1_REG2_REG_2__SCAN_IN), .ZN(n6902) );
  NOR2_X1 U8666 ( .A1(n6903), .A2(n6902), .ZN(n6986) );
  AOI211_X1 U8667 ( .C1(n6903), .C2(n6902), .A(n6986), .B(n9844), .ZN(n6912)
         );
  AOI21_X1 U8668 ( .B1(P1_REG1_REG_1__SCAN_IN), .B2(n6905), .A(n6904), .ZN(
        n6908) );
  MUX2_X1 U8669 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n5143), .S(n6922), .Z(n6907)
         );
  OR2_X1 U8670 ( .A1(n6908), .A2(n6907), .ZN(n7039) );
  INV_X1 U8671 ( .A(n7039), .ZN(n6906) );
  AOI211_X1 U8672 ( .C1(n6908), .C2(n6907), .A(n6906), .B(n9869), .ZN(n6911)
         );
  AOI22_X1 U8673 ( .A1(n9352), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n6909) );
  OAI21_X1 U8674 ( .B1(n6922), .B2(n9866), .A(n6909), .ZN(n6910) );
  OR4_X1 U8675 ( .A1(n9855), .A2(n6912), .A3(n6911), .A4(n6910), .ZN(P1_U3245)
         );
  INV_X2 U8676 ( .A(n9044), .ZN(n8437) );
  NOR2_X1 U8677 ( .A1(n6915), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9043) );
  INV_X2 U8678 ( .A(n9043), .ZN(n8435) );
  OAI222_X1 U8679 ( .A1(n8437), .A2(n4695), .B1(n8435), .B2(n6917), .C1(
        P2_U3151), .C2(n6977), .ZN(P2_U3294) );
  OAI222_X1 U8680 ( .A1(n8437), .A2(n6913), .B1(n8435), .B2(n6923), .C1(
        P2_U3151), .C2(n7021), .ZN(P2_U3293) );
  OAI222_X1 U8681 ( .A1(n8437), .A2(n10270), .B1(n8435), .B2(n6931), .C1(
        P2_U3151), .C2(n9937), .ZN(P2_U3291) );
  OAI222_X1 U8682 ( .A1(n8437), .A2(n10272), .B1(n8435), .B2(n6920), .C1(
        P2_U3151), .C2(n7054), .ZN(P2_U3292) );
  OAI222_X1 U8683 ( .A1(n8437), .A2(n6914), .B1(n8435), .B2(n6929), .C1(
        P2_U3151), .C2(n7126), .ZN(P2_U3290) );
  INV_X2 U8684 ( .A(n9817), .ZN(n9824) );
  NAND2_X2 U8685 ( .A1(n6915), .A2(P1_U3086), .ZN(n9822) );
  OAI222_X1 U8686 ( .A1(n9824), .A2(n6918), .B1(n9822), .B2(n6917), .C1(
        P1_U3086), .C2(n6916), .ZN(P1_U3354) );
  OAI222_X1 U8687 ( .A1(n8437), .A2(n10343), .B1(n8435), .B2(n6927), .C1(
        P2_U3151), .C2(n7237), .ZN(P2_U3289) );
  OAI222_X1 U8688 ( .A1(n8437), .A2(n6919), .B1(n8435), .B2(n6925), .C1(
        P2_U3151), .C2(n7310), .ZN(P2_U3288) );
  OAI222_X1 U8689 ( .A1(n9824), .A2(n6921), .B1(n9822), .B2(n6920), .C1(
        P1_U3086), .C2(n7048), .ZN(P1_U3352) );
  OAI222_X1 U8690 ( .A1(n9824), .A2(n6924), .B1(n9822), .B2(n6923), .C1(
        P1_U3086), .C2(n6922), .ZN(P1_U3353) );
  INV_X1 U8691 ( .A(n7001), .ZN(n9294) );
  OAI222_X1 U8692 ( .A1(n9824), .A2(n6926), .B1(n9822), .B2(n6925), .C1(
        P1_U3086), .C2(n9294), .ZN(P1_U3348) );
  OAI222_X1 U8693 ( .A1(n9824), .A2(n6928), .B1(n9822), .B2(n6927), .C1(
        P1_U3086), .C2(n9285), .ZN(P1_U3349) );
  OAI222_X1 U8694 ( .A1(n9824), .A2(n6930), .B1(n9822), .B2(n6929), .C1(
        P1_U3086), .C2(n9266), .ZN(P1_U3350) );
  OAI222_X1 U8695 ( .A1(n6932), .A2(n9824), .B1(P1_U3086), .B2(n9845), .C1(
        n9822), .C2(n6931), .ZN(P1_U3351) );
  INV_X1 U8696 ( .A(n6933), .ZN(n6935) );
  INV_X1 U8697 ( .A(n7002), .ZN(n9309) );
  OAI222_X1 U8698 ( .A1(n9824), .A2(n6934), .B1(n9822), .B2(n6935), .C1(
        P1_U3086), .C2(n9309), .ZN(P1_U3347) );
  OAI222_X1 U8699 ( .A1(n8437), .A2(n6936), .B1(n8435), .B2(n6935), .C1(
        P2_U3151), .C2(n8598), .ZN(P2_U3287) );
  INV_X1 U8700 ( .A(n6937), .ZN(n6940) );
  OAI222_X1 U8701 ( .A1(n8435), .A2(n6940), .B1(n6939), .B2(P2_U3151), .C1(
        n6938), .C2(n8437), .ZN(P2_U3286) );
  INV_X1 U8702 ( .A(n7005), .ZN(n9832) );
  OAI222_X1 U8703 ( .A1(n9824), .A2(n6941), .B1(n9822), .B2(n6940), .C1(n9832), 
        .C2(P1_U3086), .ZN(P1_U3346) );
  INV_X1 U8704 ( .A(n6942), .ZN(n6944) );
  OAI222_X1 U8705 ( .A1(n8435), .A2(n6944), .B1(n6943), .B2(P2_U3151), .C1(
        n10277), .C2(n8437), .ZN(P2_U3285) );
  INV_X1 U8706 ( .A(n7068), .ZN(n7072) );
  OAI222_X1 U8707 ( .A1(n9824), .A2(n10285), .B1(n9822), .B2(n6944), .C1(n7072), .C2(P1_U3086), .ZN(P1_U3345) );
  NOR2_X1 U8708 ( .A1(n6958), .A2(n10145), .ZN(P2_U3242) );
  INV_X1 U8709 ( .A(P2_D_REG_15__SCAN_IN), .ZN(n10248) );
  NOR2_X1 U8710 ( .A1(n6958), .A2(n10248), .ZN(P2_U3250) );
  NOR2_X1 U8711 ( .A1(n6958), .A2(n10060), .ZN(P2_U3253) );
  NOR2_X1 U8712 ( .A1(n6958), .A2(n10132), .ZN(P2_U3247) );
  INV_X1 U8713 ( .A(P2_D_REG_9__SCAN_IN), .ZN(n10133) );
  NOR2_X1 U8714 ( .A1(n6958), .A2(n10133), .ZN(P2_U3256) );
  NOR2_X1 U8715 ( .A1(n6958), .A2(n10229), .ZN(P2_U3248) );
  INV_X1 U8716 ( .A(P2_D_REG_10__SCAN_IN), .ZN(n10173) );
  NOR2_X1 U8717 ( .A1(n6958), .A2(n10173), .ZN(P2_U3255) );
  INV_X1 U8718 ( .A(P2_D_REG_3__SCAN_IN), .ZN(n10200) );
  NOR2_X1 U8719 ( .A1(n6958), .A2(n10200), .ZN(P2_U3262) );
  INV_X1 U8720 ( .A(P2_D_REG_7__SCAN_IN), .ZN(n10093) );
  NOR2_X1 U8721 ( .A1(n6958), .A2(n10093), .ZN(P2_U3258) );
  INV_X1 U8722 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n6946) );
  NAND2_X1 U8723 ( .A1(n7537), .A2(P2_U3893), .ZN(n6945) );
  OAI21_X1 U8724 ( .B1(P2_U3893), .B2(n6946), .A(n6945), .ZN(P2_U3491) );
  INV_X1 U8725 ( .A(n6947), .ZN(n6949) );
  OAI222_X1 U8726 ( .A1(n8437), .A2(n10300), .B1(n8435), .B2(n6949), .C1(
        P2_U3151), .C2(n6948), .ZN(P2_U3284) );
  INV_X1 U8727 ( .A(n7296), .ZN(n7079) );
  OAI222_X1 U8728 ( .A1(n9824), .A2(n6950), .B1(n9822), .B2(n6949), .C1(
        P1_U3086), .C2(n7079), .ZN(P1_U3344) );
  NOR2_X1 U8729 ( .A1(n9352), .A2(P1_U3973), .ZN(P1_U3085) );
  MUX2_X1 U8730 ( .A(n6950), .B(n8063), .S(P2_U3893), .Z(n6951) );
  INV_X1 U8731 ( .A(n6951), .ZN(P2_U3502) );
  INV_X1 U8732 ( .A(n6952), .ZN(n6954) );
  INV_X1 U8733 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n10298) );
  OAI222_X1 U8734 ( .A1(n8435), .A2(n6954), .B1(n6953), .B2(P2_U3151), .C1(
        n10298), .C2(n8437), .ZN(P2_U3283) );
  INV_X1 U8735 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n6955) );
  INV_X1 U8736 ( .A(n7293), .ZN(n7354) );
  OAI222_X1 U8737 ( .A1(n9824), .A2(n6955), .B1(n9822), .B2(n6954), .C1(n7354), 
        .C2(P1_U3086), .ZN(P1_U3343) );
  INV_X1 U8738 ( .A(n6956), .ZN(n6969) );
  AOI22_X1 U8739 ( .A1(n8643), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_13__SCAN_IN), .B2(n9044), .ZN(n6957) );
  OAI21_X1 U8740 ( .B1(n6969), .B2(n8435), .A(n6957), .ZN(P2_U3282) );
  AND2_X1 U8741 ( .A1(n8139), .A2(P2_D_REG_14__SCAN_IN), .ZN(P2_U3251) );
  AND2_X1 U8742 ( .A1(n8139), .A2(P2_D_REG_29__SCAN_IN), .ZN(P2_U3236) );
  AND2_X1 U8743 ( .A1(n8139), .A2(P2_D_REG_11__SCAN_IN), .ZN(P2_U3254) );
  AND2_X1 U8744 ( .A1(n8139), .A2(P2_D_REG_31__SCAN_IN), .ZN(P2_U3234) );
  AND2_X1 U8745 ( .A1(n8139), .A2(P2_D_REG_13__SCAN_IN), .ZN(P2_U3252) );
  AND2_X1 U8746 ( .A1(n8139), .A2(P2_D_REG_5__SCAN_IN), .ZN(P2_U3260) );
  AND2_X1 U8747 ( .A1(n8139), .A2(P2_D_REG_6__SCAN_IN), .ZN(P2_U3259) );
  AND2_X1 U8748 ( .A1(n8139), .A2(P2_D_REG_24__SCAN_IN), .ZN(P2_U3241) );
  AND2_X1 U8749 ( .A1(n8139), .A2(P2_D_REG_26__SCAN_IN), .ZN(P2_U3239) );
  AND2_X1 U8750 ( .A1(n8139), .A2(P2_D_REG_27__SCAN_IN), .ZN(P2_U3238) );
  AND2_X1 U8751 ( .A1(n8139), .A2(P2_D_REG_4__SCAN_IN), .ZN(P2_U3261) );
  AND2_X1 U8752 ( .A1(n8139), .A2(P2_D_REG_2__SCAN_IN), .ZN(P2_U3263) );
  AND2_X1 U8753 ( .A1(n8139), .A2(P2_D_REG_8__SCAN_IN), .ZN(P2_U3257) );
  AND2_X1 U8754 ( .A1(n8139), .A2(P2_D_REG_30__SCAN_IN), .ZN(P2_U3235) );
  AND2_X1 U8755 ( .A1(n8139), .A2(P2_D_REG_25__SCAN_IN), .ZN(P2_U3240) );
  AND2_X1 U8756 ( .A1(n8139), .A2(P2_D_REG_21__SCAN_IN), .ZN(P2_U3244) );
  AND2_X1 U8757 ( .A1(n8139), .A2(P2_D_REG_20__SCAN_IN), .ZN(P2_U3245) );
  AND2_X1 U8758 ( .A1(n8139), .A2(P2_D_REG_28__SCAN_IN), .ZN(P2_U3237) );
  AND2_X1 U8759 ( .A1(n8139), .A2(P2_D_REG_16__SCAN_IN), .ZN(P2_U3249) );
  AND2_X1 U8760 ( .A1(n8139), .A2(P2_D_REG_19__SCAN_IN), .ZN(P2_U3246) );
  AND2_X1 U8761 ( .A1(n8139), .A2(P2_D_REG_22__SCAN_IN), .ZN(P2_U3243) );
  INV_X1 U8762 ( .A(n6959), .ZN(n6960) );
  AOI22_X1 U8763 ( .A1(n8139), .A2(n4922), .B1(n8135), .B2(n6960), .ZN(
        P2_U3376) );
  INV_X1 U8764 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n6968) );
  NAND3_X1 U8765 ( .A1(n9386), .A2(P1_IR_REG_0__SCAN_IN), .A3(n6876), .ZN(
        n6967) );
  AOI21_X1 U8766 ( .B1(n8195), .B2(n6876), .A(n6963), .ZN(n6962) );
  MUX2_X1 U8767 ( .A(n6963), .B(n6962), .S(n6961), .Z(n6964) );
  AOI22_X1 U8768 ( .A1(n6965), .A2(n6964), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        P1_U3086), .ZN(n6966) );
  OAI211_X1 U8769 ( .C1(n9875), .C2(n6968), .A(n6967), .B(n6966), .ZN(P1_U3243) );
  INV_X1 U8770 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n6970) );
  INV_X1 U8771 ( .A(n7474), .ZN(n7480) );
  OAI222_X1 U8772 ( .A1(n9824), .A2(n6970), .B1(n9822), .B2(n6969), .C1(
        P1_U3086), .C2(n7480), .ZN(P1_U3342) );
  INV_X1 U8773 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n6985) );
  AOI21_X1 U8774 ( .B1(n6257), .B2(n6972), .A(n6971), .ZN(n6976) );
  AOI21_X1 U8775 ( .B1(n6256), .B2(n6974), .A(n6973), .ZN(n6975) );
  OAI22_X1 U8776 ( .A1(n6976), .A2(n9929), .B1(n9930), .B2(n6975), .ZN(n6979)
         );
  OAI22_X1 U8777 ( .A1(n9938), .A2(n6977), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7533), .ZN(n6978) );
  NOR2_X1 U8778 ( .A1(n6979), .A2(n6978), .ZN(n6984) );
  OAI211_X1 U8779 ( .C1(n6982), .C2(n6981), .A(n9918), .B(n6980), .ZN(n6983)
         );
  OAI211_X1 U8780 ( .C1(n6985), .C2(n8735), .A(n6984), .B(n6983), .ZN(P2_U3183) );
  AOI22_X1 U8781 ( .A1(n7068), .A2(n5271), .B1(P1_REG2_REG_10__SCAN_IN), .B2(
        n7072), .ZN(n6993) );
  INV_X1 U8782 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n7386) );
  INV_X1 U8783 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n7405) );
  OR2_X1 U8784 ( .A1(n7048), .A2(n7405), .ZN(n9839) );
  NAND2_X1 U8785 ( .A1(n7048), .A2(n7405), .ZN(n6987) );
  NAND2_X1 U8786 ( .A1(n9839), .A2(n6987), .ZN(n7041) );
  MUX2_X1 U8787 ( .A(n6989), .B(P1_REG2_REG_4__SCAN_IN), .S(n9845), .Z(n9840)
         );
  INV_X1 U8788 ( .A(n9843), .ZN(n6988) );
  OAI21_X1 U8789 ( .B1(n9845), .B2(n6989), .A(n6988), .ZN(n9270) );
  MUX2_X1 U8790 ( .A(n6990), .B(P1_REG2_REG_5__SCAN_IN), .S(n9266), .Z(n9271)
         );
  NAND2_X1 U8791 ( .A1(n9270), .A2(n9271), .ZN(n9269) );
  OAI21_X1 U8792 ( .B1(n6990), .B2(n9266), .A(n9269), .ZN(n9282) );
  XNOR2_X1 U8793 ( .A(n9285), .B(P1_REG2_REG_6__SCAN_IN), .ZN(n9283) );
  NAND2_X1 U8794 ( .A1(n9282), .A2(n9283), .ZN(n9281) );
  OAI21_X1 U8795 ( .B1(n7386), .B2(n9285), .A(n9281), .ZN(n9299) );
  MUX2_X1 U8796 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n7424), .S(n7001), .Z(n9298)
         );
  NAND2_X1 U8797 ( .A1(n9299), .A2(n9298), .ZN(n9297) );
  OAI21_X1 U8798 ( .B1(n9294), .B2(n7424), .A(n9297), .ZN(n9314) );
  INV_X1 U8799 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n7445) );
  MUX2_X1 U8800 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n7445), .S(n7002), .Z(n9313)
         );
  NOR2_X1 U8801 ( .A1(n7005), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6991) );
  AOI21_X1 U8802 ( .B1(n7005), .B2(P1_REG2_REG_9__SCAN_IN), .A(n6991), .ZN(
        n9827) );
  OAI21_X1 U8803 ( .B1(n7005), .B2(P1_REG2_REG_9__SCAN_IN), .A(n9826), .ZN(
        n6992) );
  AOI211_X1 U8804 ( .C1(n6993), .C2(n6992), .A(n7067), .B(n9844), .ZN(n7013)
         );
  NAND2_X1 U8805 ( .A1(n6994), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n7038) );
  MUX2_X1 U8806 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n6995), .S(n7048), .Z(n7037)
         );
  AOI21_X1 U8807 ( .B1(n7039), .B2(n7038), .A(n7037), .ZN(n9849) );
  NOR2_X1 U8808 ( .A1(n7048), .A2(n6995), .ZN(n9848) );
  MUX2_X1 U8809 ( .A(n6996), .B(P1_REG1_REG_4__SCAN_IN), .S(n9845), .Z(n9847)
         );
  OAI21_X1 U8810 ( .B1(n9849), .B2(n9848), .A(n9847), .ZN(n9846) );
  INV_X1 U8811 ( .A(n9845), .ZN(n6997) );
  NAND2_X1 U8812 ( .A1(n6997), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n9274) );
  MUX2_X1 U8813 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n5196), .S(n9266), .Z(n9273)
         );
  AOI21_X1 U8814 ( .B1(n9846), .B2(n9274), .A(n9273), .ZN(n9272) );
  NOR2_X1 U8815 ( .A1(n9266), .A2(n5196), .ZN(n9284) );
  MUX2_X1 U8816 ( .A(n6998), .B(P1_REG1_REG_6__SCAN_IN), .S(n9285), .Z(n6999)
         );
  OAI21_X1 U8817 ( .B1(n9272), .B2(n9284), .A(n6999), .ZN(n9302) );
  INV_X1 U8818 ( .A(n9285), .ZN(n7000) );
  NAND2_X1 U8819 ( .A1(n7000), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n9301) );
  MUX2_X1 U8820 ( .A(n5228), .B(P1_REG1_REG_7__SCAN_IN), .S(n7001), .Z(n9300)
         );
  AOI21_X1 U8821 ( .B1(n9302), .B2(n9301), .A(n9300), .ZN(n9317) );
  NOR2_X1 U8822 ( .A1(n9294), .A2(n5228), .ZN(n9316) );
  MUX2_X1 U8823 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n7003), .S(n7002), .Z(n9315)
         );
  OAI21_X1 U8824 ( .B1(n9317), .B2(n9316), .A(n9315), .ZN(n9319) );
  OAI21_X1 U8825 ( .B1(n7003), .B2(n9309), .A(n9319), .ZN(n9830) );
  MUX2_X1 U8826 ( .A(n7004), .B(P1_REG1_REG_9__SCAN_IN), .S(n7005), .Z(n9831)
         );
  NOR2_X1 U8827 ( .A1(n9830), .A2(n9831), .ZN(n9829) );
  NOR2_X1 U8828 ( .A1(n7005), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n7006) );
  NOR2_X1 U8829 ( .A1(n9829), .A2(n7006), .ZN(n7009) );
  MUX2_X1 U8830 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n7007), .S(n7068), .Z(n7008)
         );
  NAND2_X1 U8831 ( .A1(n7008), .A2(n7009), .ZN(n7071) );
  OAI211_X1 U8832 ( .C1(n7009), .C2(n7008), .A(n9386), .B(n7071), .ZN(n7011)
         );
  INV_X1 U8833 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n10192) );
  NOR2_X1 U8834 ( .A1(n10192), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7916) );
  AOI21_X1 U8835 ( .B1(n9352), .B2(P1_ADDR_REG_10__SCAN_IN), .A(n7916), .ZN(
        n7010) );
  OAI211_X1 U8836 ( .C1(n9866), .C2(n7072), .A(n7011), .B(n7010), .ZN(n7012)
         );
  OR2_X1 U8837 ( .A1(n7013), .A2(n7012), .ZN(P1_U3253) );
  INV_X1 U8838 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n7015) );
  INV_X1 U8839 ( .A(n7014), .ZN(n7017) );
  INV_X1 U8840 ( .A(n9324), .ZN(n9331) );
  OAI222_X1 U8841 ( .A1(n9824), .A2(n7015), .B1(n9822), .B2(n7017), .C1(
        P1_U3086), .C2(n9331), .ZN(P1_U3341) );
  INV_X1 U8842 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n7018) );
  OAI222_X1 U8843 ( .A1(n8437), .A2(n7018), .B1(n8435), .B2(n7017), .C1(
        P2_U3151), .C2(n7016), .ZN(P2_U3281) );
  INV_X1 U8844 ( .A(n7019), .ZN(n7065) );
  AOI22_X1 U8845 ( .A1(n8674), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_15__SCAN_IN), .B2(n9044), .ZN(n7020) );
  OAI21_X1 U8846 ( .B1(n7065), .B2(n8435), .A(n7020), .ZN(P2_U3280) );
  OAI22_X1 U8847 ( .A1(n9938), .A2(n7021), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9942), .ZN(n7031) );
  AOI21_X1 U8848 ( .B1(n7024), .B2(n7023), .A(n7022), .ZN(n7029) );
  AOI21_X1 U8849 ( .B1(n7027), .B2(n7026), .A(n7025), .ZN(n7028) );
  OAI22_X1 U8850 ( .A1(n7029), .A2(n9929), .B1(n9930), .B2(n7028), .ZN(n7030)
         );
  AOI211_X1 U8851 ( .C1(n9934), .C2(P2_ADDR_REG_2__SCAN_IN), .A(n7031), .B(
        n7030), .ZN(n7036) );
  OAI211_X1 U8852 ( .C1(n7034), .C2(n7033), .A(n7032), .B(n9918), .ZN(n7035)
         );
  NAND2_X1 U8853 ( .A1(n7036), .A2(n7035), .ZN(P2_U3184) );
  AND3_X1 U8854 ( .A1(n7039), .A2(n7038), .A3(n7037), .ZN(n7040) );
  NOR3_X1 U8855 ( .A1(n9869), .A2(n9849), .A3(n7040), .ZN(n7044) );
  AOI211_X1 U8856 ( .C1(n7042), .C2(n7041), .A(n9841), .B(n9844), .ZN(n7043)
         );
  NOR2_X1 U8857 ( .A1(n7044), .A2(n7043), .ZN(n7047) );
  NAND2_X1 U8858 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_U3086), .ZN(n7254) );
  INV_X1 U8859 ( .A(n7254), .ZN(n7045) );
  AOI21_X1 U8860 ( .B1(n9352), .B2(P1_ADDR_REG_3__SCAN_IN), .A(n7045), .ZN(
        n7046) );
  OAI211_X1 U8861 ( .C1(n7048), .C2(n9866), .A(n7047), .B(n7046), .ZN(P1_U3246) );
  INV_X1 U8862 ( .A(n7049), .ZN(n7050) );
  AOI21_X1 U8863 ( .B1(n7052), .B2(n7051), .A(n7050), .ZN(n7064) );
  NOR2_X1 U8864 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7380), .ZN(n7215) );
  INV_X1 U8865 ( .A(n7215), .ZN(n7053) );
  OAI21_X1 U8866 ( .B1(n9938), .B2(n7054), .A(n7053), .ZN(n7062) );
  AOI21_X1 U8867 ( .B1(n7055), .B2(n7056), .A(n4517), .ZN(n7060) );
  AOI21_X1 U8868 ( .B1(n7058), .B2(n5758), .A(n7057), .ZN(n7059) );
  OAI22_X1 U8869 ( .A1(n7060), .A2(n9929), .B1(n9930), .B2(n7059), .ZN(n7061)
         );
  AOI211_X1 U8870 ( .C1(n9934), .C2(P2_ADDR_REG_3__SCAN_IN), .A(n7062), .B(
        n7061), .ZN(n7063) );
  OAI21_X1 U8871 ( .B1(n7064), .B2(n7248), .A(n7063), .ZN(P2_U3185) );
  INV_X1 U8872 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n7066) );
  INV_X1 U8873 ( .A(n9338), .ZN(n9343) );
  OAI222_X1 U8874 ( .A1(n9824), .A2(n7066), .B1(n9822), .B2(n7065), .C1(
        P1_U3086), .C2(n9343), .ZN(P1_U3340) );
  AOI22_X1 U8875 ( .A1(P1_REG2_REG_11__SCAN_IN), .A2(n7079), .B1(n7296), .B2(
        n5286), .ZN(n7069) );
  AOI211_X1 U8876 ( .C1(n7070), .C2(n7069), .A(n7289), .B(n9844), .ZN(n7081)
         );
  OAI21_X1 U8877 ( .B1(n7072), .B2(n7007), .A(n7071), .ZN(n7075) );
  MUX2_X1 U8878 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n7073), .S(n7296), .Z(n7074)
         );
  NAND2_X1 U8879 ( .A1(n7074), .A2(n7075), .ZN(n7294) );
  OAI211_X1 U8880 ( .C1(n7075), .C2(n7074), .A(n9386), .B(n7294), .ZN(n7078)
         );
  NAND2_X1 U8881 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n9196) );
  INV_X1 U8882 ( .A(n9196), .ZN(n7076) );
  AOI21_X1 U8883 ( .B1(n9352), .B2(P1_ADDR_REG_11__SCAN_IN), .A(n7076), .ZN(
        n7077) );
  OAI211_X1 U8884 ( .C1(n9866), .C2(n7079), .A(n7078), .B(n7077), .ZN(n7080)
         );
  OR2_X1 U8885 ( .A1(n7081), .A2(n7080), .ZN(P1_U3254) );
  NAND2_X1 U8886 ( .A1(n7537), .A2(n7206), .ZN(n8253) );
  NAND2_X1 U8887 ( .A1(n7532), .A2(n8253), .ZN(n8217) );
  OAI21_X1 U8888 ( .B1(n8912), .B2(n9970), .A(n8217), .ZN(n7082) );
  NAND2_X1 U8889 ( .A1(n5739), .A2(n8909), .ZN(n7356) );
  OAI211_X1 U8890 ( .C1(n7206), .C2(n10005), .A(n7082), .B(n7356), .ZN(n7170)
         );
  NAND2_X1 U8891 ( .A1(n7170), .A2(n10029), .ZN(n7083) );
  OAI21_X1 U8892 ( .B1(n10029), .B2(n6210), .A(n7083), .ZN(P2_U3459) );
  XNOR2_X1 U8893 ( .A(n7084), .B(n6687), .ZN(n7085) );
  OAI222_X1 U8894 ( .A1(n9705), .A2(n7087), .B1(n9591), .B2(n7086), .C1(n7085), 
        .C2(n9498), .ZN(n7504) );
  INV_X1 U8895 ( .A(n7088), .ZN(n7149) );
  AOI211_X1 U8896 ( .C1(n7175), .C2(n7149), .A(n9567), .B(n4675), .ZN(n7505)
         );
  NOR2_X1 U8897 ( .A1(n7504), .A2(n7505), .ZN(n7167) );
  INV_X1 U8898 ( .A(n7089), .ZN(n7091) );
  XNOR2_X1 U8899 ( .A(n7091), .B(n7090), .ZN(n7508) );
  OAI22_X1 U8900 ( .A1(n9644), .A2(n6411), .B1(n9910), .B2(n5143), .ZN(n7092)
         );
  AOI21_X1 U8901 ( .B1(n9711), .B2(n7508), .A(n7092), .ZN(n7093) );
  OAI21_X1 U8902 ( .B1(n7167), .B2(n9908), .A(n7093), .ZN(P1_U3524) );
  INV_X1 U8903 ( .A(n7094), .ZN(n7103) );
  OR2_X1 U8904 ( .A1(n7095), .A2(n7103), .ZN(n7111) );
  INV_X1 U8905 ( .A(n7116), .ZN(n7096) );
  NAND2_X1 U8906 ( .A1(n7111), .A2(n7096), .ZN(n7107) );
  NAND2_X1 U8907 ( .A1(n7098), .A2(n7097), .ZN(n7099) );
  NOR2_X1 U8908 ( .A1(n7100), .A2(n7099), .ZN(n7106) );
  INV_X1 U8909 ( .A(n7101), .ZN(n7102) );
  OAI21_X1 U8910 ( .B1(n7104), .B2(n7103), .A(n7102), .ZN(n7105) );
  NAND3_X1 U8911 ( .A1(n7107), .A2(n7106), .A3(n7105), .ZN(n7108) );
  NAND2_X1 U8912 ( .A1(n7108), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7113) );
  INV_X1 U8913 ( .A(n7109), .ZN(n7110) );
  NOR2_X1 U8914 ( .A1(n7110), .A2(n7355), .ZN(n8423) );
  NAND2_X1 U8915 ( .A1(n7111), .A2(n8423), .ZN(n7112) );
  NOR2_X1 U8916 ( .A1(n8558), .A2(P2_U3151), .ZN(n7270) );
  INV_X1 U8917 ( .A(n7114), .ZN(n7115) );
  NAND2_X1 U8918 ( .A1(n7119), .A2(n7115), .ZN(n7118) );
  OR2_X1 U8919 ( .A1(n7121), .A2(n7116), .ZN(n7117) );
  NAND2_X1 U8920 ( .A1(n7119), .A2(n10015), .ZN(n7120) );
  AOI22_X1 U8921 ( .A1(n8545), .A2(n8217), .B1(n7535), .B2(n8576), .ZN(n7124)
         );
  OR2_X1 U8922 ( .A1(n7121), .A2(n7355), .ZN(n7213) );
  INV_X1 U8923 ( .A(n7213), .ZN(n7122) );
  INV_X1 U8924 ( .A(n8566), .ZN(n8548) );
  NAND2_X1 U8925 ( .A1(n8548), .A2(n5739), .ZN(n7123) );
  OAI211_X1 U8926 ( .C1(n7270), .C2(n7125), .A(n7124), .B(n7123), .ZN(P2_U3172) );
  NAND2_X1 U8927 ( .A1(P2_U3151), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n7467) );
  OAI21_X1 U8928 ( .B1(n9938), .B2(n7126), .A(n7467), .ZN(n7134) );
  AOI21_X1 U8929 ( .B1(n5787), .B2(n7128), .A(n7127), .ZN(n7132) );
  AOI21_X1 U8930 ( .B1(n7517), .B2(n7130), .A(n7129), .ZN(n7131) );
  OAI22_X1 U8931 ( .A1(n7132), .A2(n9930), .B1(n9929), .B2(n7131), .ZN(n7133)
         );
  AOI211_X1 U8932 ( .C1(n9934), .C2(P2_ADDR_REG_5__SCAN_IN), .A(n7134), .B(
        n7133), .ZN(n7139) );
  OAI211_X1 U8933 ( .C1(n7137), .C2(n7136), .A(n7135), .B(n9918), .ZN(n7138)
         );
  NAND2_X1 U8934 ( .A1(n7139), .A2(n7138), .ZN(P2_U3187) );
  INV_X1 U8935 ( .A(n9142), .ZN(n7140) );
  NAND2_X1 U8936 ( .A1(n7140), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9104) );
  INV_X1 U8937 ( .A(n9104), .ZN(n7145) );
  OAI22_X1 U8938 ( .A1(n9205), .A2(n7141), .B1(n9247), .B2(n7150), .ZN(n7142)
         );
  AOI21_X1 U8939 ( .B1(n9244), .B2(n6427), .A(n7142), .ZN(n7143) );
  OAI21_X1 U8940 ( .B1(n7145), .B2(n7144), .A(n7143), .ZN(P1_U3232) );
  INV_X1 U8941 ( .A(n7146), .ZN(n7147) );
  AOI21_X1 U8942 ( .B1(n7148), .B2(n7152), .A(n7147), .ZN(n7401) );
  INV_X1 U8943 ( .A(n7401), .ZN(n7157) );
  OAI211_X1 U8944 ( .C1(n7158), .C2(n7150), .A(n7149), .B(n9628), .ZN(n7395)
         );
  OAI21_X1 U8945 ( .B1(n6419), .B2(n9705), .A(n7395), .ZN(n7156) );
  XNOR2_X1 U8946 ( .A(n7152), .B(n7151), .ZN(n7154) );
  AND2_X1 U8947 ( .A1(n9881), .A2(n9264), .ZN(n7153) );
  AOI21_X1 U8948 ( .B1(n7154), .B2(n9893), .A(n7153), .ZN(n7396) );
  INV_X1 U8949 ( .A(n7396), .ZN(n7155) );
  AOI211_X1 U8950 ( .C1(n9903), .C2(n7157), .A(n7156), .B(n7155), .ZN(n7162)
         );
  OAI22_X1 U8951 ( .A1(n9755), .A2(n7158), .B1(n9906), .B2(n5130), .ZN(n7159)
         );
  INV_X1 U8952 ( .A(n7159), .ZN(n7160) );
  OAI21_X1 U8953 ( .B1(n7162), .B2(n9905), .A(n7160), .ZN(P1_U3456) );
  AOI22_X1 U8954 ( .A1(n9734), .A2(n4417), .B1(n9908), .B2(
        P1_REG1_REG_1__SCAN_IN), .ZN(n7161) );
  OAI21_X1 U8955 ( .B1(n7162), .B2(n9908), .A(n7161), .ZN(P1_U3523) );
  INV_X1 U8956 ( .A(n7163), .ZN(n7168) );
  OAI222_X1 U8957 ( .A1(n8435), .A2(n7168), .B1(n7164), .B2(P2_U3151), .C1(
        n10164), .C2(n8437), .ZN(P2_U3279) );
  OAI22_X1 U8958 ( .A1(n9755), .A2(n6411), .B1(n9906), .B2(n5145), .ZN(n7165)
         );
  AOI21_X1 U8959 ( .B1(n9786), .B2(n7508), .A(n7165), .ZN(n7166) );
  OAI21_X1 U8960 ( .B1(n7167), .B2(n9905), .A(n7166), .ZN(P1_U3459) );
  INV_X1 U8961 ( .A(n9365), .ZN(n9358) );
  OAI222_X1 U8962 ( .A1(n9824), .A2(n7169), .B1(n9822), .B2(n7168), .C1(n9358), 
        .C2(P1_U3086), .ZN(P1_U3339) );
  INV_X1 U8963 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n7172) );
  NAND2_X1 U8964 ( .A1(n7170), .A2(n10016), .ZN(n7171) );
  OAI21_X1 U8965 ( .B1(n10016), .B2(n7172), .A(n7171), .ZN(P2_U3390) );
  XOR2_X1 U8966 ( .A(n7174), .B(n7173), .Z(n7178) );
  AOI22_X1 U8967 ( .A1(n7175), .A2(n9209), .B1(n9244), .B2(n9263), .ZN(n7177)
         );
  AOI22_X1 U8968 ( .A1(n9225), .A2(n6427), .B1(n9104), .B2(
        P1_REG3_REG_2__SCAN_IN), .ZN(n7176) );
  OAI211_X1 U8969 ( .C1(n7178), .C2(n9205), .A(n7177), .B(n7176), .ZN(P1_U3237) );
  OAI21_X1 U8970 ( .B1(n7181), .B2(n7180), .A(n7179), .ZN(n7409) );
  OAI21_X1 U8971 ( .B1(n7184), .B2(n7183), .A(n7182), .ZN(n7185) );
  AOI22_X1 U8972 ( .A1(n7185), .A2(n9893), .B1(n9881), .B2(n9262), .ZN(n7411)
         );
  INV_X1 U8973 ( .A(n7411), .ZN(n7190) );
  INV_X1 U8974 ( .A(n7221), .ZN(n7186) );
  AOI211_X1 U8975 ( .C1(n7191), .C2(n7187), .A(n9567), .B(n7186), .ZN(n7403)
         );
  INV_X1 U8976 ( .A(n7403), .ZN(n7188) );
  OAI21_X1 U8977 ( .B1(n7406), .B2(n9705), .A(n7188), .ZN(n7189) );
  AOI211_X1 U8978 ( .C1(n9903), .C2(n7409), .A(n7190), .B(n7189), .ZN(n7195)
         );
  AOI22_X1 U8979 ( .A1(n9734), .A2(n7191), .B1(n9908), .B2(
        P1_REG1_REG_3__SCAN_IN), .ZN(n7192) );
  OAI21_X1 U8980 ( .B1(n7195), .B2(n9908), .A(n7192), .ZN(P1_U3525) );
  OAI22_X1 U8981 ( .A1(n9755), .A2(n6440), .B1(n9906), .B2(n5167), .ZN(n7193)
         );
  INV_X1 U8982 ( .A(n7193), .ZN(n7194) );
  OAI21_X1 U8983 ( .B1(n7195), .B2(n9905), .A(n7194), .ZN(P1_U3462) );
  INV_X1 U8984 ( .A(n8558), .ZN(n8570) );
  INV_X1 U8985 ( .A(n7196), .ZN(n7199) );
  NAND2_X1 U8986 ( .A1(n7199), .A2(n4412), .ZN(n7203) );
  INV_X1 U8987 ( .A(n7198), .ZN(n7201) );
  NOR2_X1 U8988 ( .A1(n7201), .A2(n7200), .ZN(n7202) );
  XNOR2_X1 U8989 ( .A(n7207), .B(n5739), .ZN(n7267) );
  INV_X1 U8990 ( .A(n7209), .ZN(n8182) );
  INV_X1 U8991 ( .A(n7532), .ZN(n7205) );
  OAI22_X1 U8992 ( .A1(n7267), .A2(n7268), .B1(n7207), .B2(n5739), .ZN(n7260)
         );
  XNOR2_X1 U8993 ( .A(n7209), .B(n5753), .ZN(n7208) );
  XNOR2_X1 U8994 ( .A(n7208), .B(n5755), .ZN(n7259) );
  INV_X1 U8995 ( .A(n5755), .ZN(n7269) );
  AOI21_X1 U8996 ( .B1(n7260), .B2(n7259), .A(n4986), .ZN(n7211) );
  XNOR2_X1 U8997 ( .A(n7209), .B(n7381), .ZN(n7277) );
  XNOR2_X1 U8998 ( .A(n7277), .B(n5772), .ZN(n7210) );
  NAND2_X1 U8999 ( .A1(n7211), .A2(n7210), .ZN(n7280) );
  OAI211_X1 U9000 ( .C1(n7211), .C2(n7210), .A(n7280), .B(n8545), .ZN(n7217)
         );
  NOR2_X2 U9001 ( .A1(n7213), .A2(n7212), .ZN(n8568) );
  INV_X1 U9002 ( .A(n8592), .ZN(n7468) );
  OAI22_X1 U9003 ( .A1(n8550), .A2(n7269), .B1(n7468), .B2(n8566), .ZN(n7214)
         );
  AOI211_X1 U9004 ( .C1(n7381), .C2(n8576), .A(n7215), .B(n7214), .ZN(n7216)
         );
  OAI211_X1 U9005 ( .C1(P2_REG3_REG_3__SCAN_IN), .C2(n8570), .A(n7217), .B(
        n7216), .ZN(P2_U3158) );
  OAI21_X1 U9006 ( .B1(n7220), .B2(n7219), .A(n7218), .ZN(n7326) );
  AOI211_X1 U9007 ( .C1(n7322), .C2(n7221), .A(n9567), .B(n7490), .ZN(n7321)
         );
  NOR2_X1 U9008 ( .A1(n7223), .A2(n7222), .ZN(n7228) );
  OAI21_X1 U9009 ( .B1(n7225), .B2(n7224), .A(n9893), .ZN(n7227) );
  AOI22_X1 U9010 ( .A1(n9881), .A2(n9261), .B1(n9723), .B2(n9263), .ZN(n7226)
         );
  OAI21_X1 U9011 ( .B1(n7228), .B2(n7227), .A(n7226), .ZN(n7319) );
  AOI211_X1 U9012 ( .C1(n9903), .C2(n7326), .A(n7321), .B(n7319), .ZN(n7233)
         );
  INV_X1 U9013 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n7229) );
  OAI22_X1 U9014 ( .A1(n9755), .A2(n7362), .B1(n9906), .B2(n7229), .ZN(n7230)
         );
  INV_X1 U9015 ( .A(n7230), .ZN(n7231) );
  OAI21_X1 U9016 ( .B1(n7233), .B2(n9905), .A(n7231), .ZN(P1_U3465) );
  AOI22_X1 U9017 ( .A1(n9734), .A2(n7322), .B1(n9908), .B2(
        P1_REG1_REG_4__SCAN_IN), .ZN(n7232) );
  OAI21_X1 U9018 ( .B1(n7233), .B2(n9908), .A(n7232), .ZN(P1_U3526) );
  AOI21_X1 U9019 ( .B1(n7236), .B2(n7235), .A(n7234), .ZN(n7249) );
  NAND2_X1 U9020 ( .A1(P2_U3151), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n7576) );
  OAI21_X1 U9021 ( .B1(n9938), .B2(n7237), .A(n7576), .ZN(n7242) );
  AOI21_X1 U9022 ( .B1(n4516), .B2(n7239), .A(n7238), .ZN(n7240) );
  NOR2_X1 U9023 ( .A1(n7240), .A2(n9930), .ZN(n7241) );
  AOI211_X1 U9024 ( .C1(n9934), .C2(P2_ADDR_REG_6__SCAN_IN), .A(n7242), .B(
        n7241), .ZN(n7247) );
  AOI21_X1 U9025 ( .B1(n4515), .B2(n7244), .A(n7243), .ZN(n7245) );
  OR2_X1 U9026 ( .A1(n7245), .A2(n9929), .ZN(n7246) );
  OAI211_X1 U9027 ( .C1(n7249), .C2(n7248), .A(n7247), .B(n7246), .ZN(P2_U3188) );
  INV_X1 U9028 ( .A(n7250), .ZN(n7265) );
  AOI22_X1 U9029 ( .A1(n8708), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_17__SCAN_IN), .B2(n9044), .ZN(n7251) );
  OAI21_X1 U9030 ( .B1(n7265), .B2(n8435), .A(n7251), .ZN(P2_U3278) );
  XOR2_X1 U9031 ( .A(n7253), .B(n7252), .Z(n7258) );
  INV_X1 U9032 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n7402) );
  AOI22_X1 U9033 ( .A1(n9244), .A2(n9262), .B1(n9225), .B2(n9264), .ZN(n7255)
         );
  OAI211_X1 U9034 ( .C1(n6440), .C2(n9247), .A(n7255), .B(n7254), .ZN(n7256)
         );
  AOI21_X1 U9035 ( .B1(n9229), .B2(n7402), .A(n7256), .ZN(n7257) );
  OAI21_X1 U9036 ( .B1(n7258), .B2(n9205), .A(n7257), .ZN(P1_U3218) );
  XOR2_X1 U9037 ( .A(n7260), .B(n7259), .Z(n7264) );
  OAI22_X1 U9038 ( .A1(n8554), .A2(n9966), .B1(n8566), .B2(n9952), .ZN(n7262)
         );
  NOR2_X1 U9039 ( .A1(n7270), .A2(n9942), .ZN(n7261) );
  AOI211_X1 U9040 ( .C1(n8568), .C2(n5739), .A(n7262), .B(n7261), .ZN(n7263)
         );
  OAI21_X1 U9041 ( .B1(n7264), .B2(n8571), .A(n7263), .ZN(P2_U3177) );
  INV_X1 U9042 ( .A(n9859), .ZN(n9867) );
  OAI222_X1 U9043 ( .A1(n9824), .A2(n7266), .B1(n9822), .B2(n7265), .C1(
        P1_U3086), .C2(n9867), .ZN(P1_U3338) );
  XOR2_X1 U9044 ( .A(n7267), .B(n7268), .Z(n7274) );
  OAI22_X1 U9045 ( .A1(n8554), .A2(n9961), .B1(n8566), .B2(n7269), .ZN(n7272)
         );
  NOR2_X1 U9046 ( .A1(n7270), .A2(n7533), .ZN(n7271) );
  AOI211_X1 U9047 ( .C1(n8568), .C2(n7537), .A(n7272), .B(n7271), .ZN(n7273)
         );
  OAI21_X1 U9048 ( .B1(n8571), .B2(n7274), .A(n7273), .ZN(P2_U3162) );
  INV_X1 U9049 ( .A(n7275), .ZN(n7303) );
  AOI22_X1 U9050 ( .A1(n9381), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n9817), .ZN(n7276) );
  OAI21_X1 U9051 ( .B1(n7303), .B2(n9822), .A(n7276), .ZN(P1_U3337) );
  XNOR2_X1 U9052 ( .A(n7209), .B(n9978), .ZN(n7463) );
  XNOR2_X1 U9053 ( .A(n7463), .B(n8592), .ZN(n7282) );
  AOI21_X1 U9054 ( .B1(n7282), .B2(n7281), .A(n7465), .ZN(n7288) );
  NAND2_X1 U9055 ( .A1(P2_U3151), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n9935) );
  INV_X1 U9056 ( .A(n9935), .ZN(n7284) );
  OAI22_X1 U9057 ( .A1(n8550), .A2(n9952), .B1(n4972), .B2(n8566), .ZN(n7283)
         );
  AOI211_X1 U9058 ( .C1(n7434), .C2(n8576), .A(n7284), .B(n7283), .ZN(n7287)
         );
  INV_X1 U9059 ( .A(n7285), .ZN(n7433) );
  NAND2_X1 U9060 ( .A1(n8558), .A2(n7433), .ZN(n7286) );
  OAI211_X1 U9061 ( .C1(n7288), .C2(n8571), .A(n7287), .B(n7286), .ZN(P2_U3170) );
  AOI22_X1 U9062 ( .A1(n7474), .A2(n5320), .B1(P1_REG2_REG_13__SCAN_IN), .B2(
        n7480), .ZN(n7292) );
  XNOR2_X1 U9063 ( .A(n7293), .B(n7290), .ZN(n7345) );
  NAND2_X1 U9064 ( .A1(n7347), .A2(n7345), .ZN(n7346) );
  OAI21_X1 U9065 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(n7293), .A(n7346), .ZN(
        n7291) );
  NOR2_X1 U9066 ( .A1(n7292), .A2(n7291), .ZN(n7473) );
  AOI211_X1 U9067 ( .C1(n7292), .C2(n7291), .A(n7473), .B(n9844), .ZN(n7302)
         );
  XNOR2_X1 U9068 ( .A(n7480), .B(P1_REG1_REG_13__SCAN_IN), .ZN(n7298) );
  INV_X1 U9069 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n7987) );
  MUX2_X1 U9070 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n7987), .S(n7293), .Z(n7343)
         );
  INV_X1 U9071 ( .A(n7294), .ZN(n7295) );
  AOI21_X1 U9072 ( .B1(n7296), .B2(P1_REG1_REG_11__SCAN_IN), .A(n7295), .ZN(
        n7344) );
  AND2_X1 U9073 ( .A1(n7343), .A2(n7344), .ZN(n7341) );
  AOI21_X1 U9074 ( .B1(n7987), .B2(n7354), .A(n7341), .ZN(n7297) );
  NAND2_X1 U9075 ( .A1(n7297), .A2(n7298), .ZN(n7478) );
  OAI211_X1 U9076 ( .C1(n7298), .C2(n7297), .A(n9386), .B(n7478), .ZN(n7300)
         );
  NOR2_X1 U9077 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n10341), .ZN(n7973) );
  AOI21_X1 U9078 ( .B1(n9352), .B2(P1_ADDR_REG_13__SCAN_IN), .A(n7973), .ZN(
        n7299) );
  OAI211_X1 U9079 ( .C1(n9866), .C2(n7480), .A(n7300), .B(n7299), .ZN(n7301)
         );
  OR2_X1 U9080 ( .A1(n7302), .A2(n7301), .ZN(P1_U3256) );
  OAI222_X1 U9081 ( .A1(n8435), .A2(n7303), .B1(n8731), .B2(P2_U3151), .C1(
        n10055), .C2(n8437), .ZN(P2_U3277) );
  INV_X1 U9082 ( .A(n7304), .ZN(n8603) );
  AOI21_X1 U9083 ( .B1(n7306), .B2(n7305), .A(n8603), .ZN(n7318) );
  XNOR2_X1 U9084 ( .A(n7308), .B(n7307), .ZN(n7309) );
  NAND2_X1 U9085 ( .A1(n7309), .A2(n9918), .ZN(n7317) );
  NAND2_X1 U9086 ( .A1(P2_U3151), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n7673) );
  OAI21_X1 U9087 ( .B1(n9938), .B2(n7310), .A(n7673), .ZN(n7315) );
  NAND2_X1 U9088 ( .A1(n7312), .A2(n5811), .ZN(n7313) );
  AOI21_X1 U9089 ( .B1(n7311), .B2(n7313), .A(n9929), .ZN(n7314) );
  AOI211_X1 U9090 ( .C1(n9934), .C2(P2_ADDR_REG_7__SCAN_IN), .A(n7315), .B(
        n7314), .ZN(n7316) );
  OAI211_X1 U9091 ( .C1(n7318), .C2(n9930), .A(n7317), .B(n7316), .ZN(P2_U3189) );
  INV_X1 U9092 ( .A(n7319), .ZN(n7328) );
  INV_X1 U9093 ( .A(n7320), .ZN(n7368) );
  INV_X1 U9094 ( .A(n9886), .ZN(n9632) );
  AOI22_X1 U9095 ( .A1(n7321), .A2(n9578), .B1(n7368), .B2(n9632), .ZN(n7324)
         );
  NAND2_X1 U9096 ( .A1(n9620), .A2(n7322), .ZN(n7323) );
  OAI211_X1 U9097 ( .C1(n6989), .C2(n9560), .A(n7324), .B(n7323), .ZN(n7325)
         );
  AOI21_X1 U9098 ( .B1(n9446), .B2(n7326), .A(n7325), .ZN(n7327) );
  OAI21_X1 U9099 ( .B1(n9889), .B2(n7328), .A(n7327), .ZN(P1_U3289) );
  XOR2_X1 U9100 ( .A(n7334), .B(n7329), .Z(n7330) );
  OAI222_X1 U9101 ( .A1(n9591), .A2(n7841), .B1(n9705), .B2(n7614), .C1(n9498), 
        .C2(n7330), .ZN(n7385) );
  INV_X1 U9102 ( .A(n7491), .ZN(n7332) );
  INV_X1 U9103 ( .A(n7331), .ZN(n7415) );
  AOI211_X1 U9104 ( .C1(n7616), .C2(n7332), .A(n9567), .B(n7415), .ZN(n7390)
         );
  NOR2_X1 U9105 ( .A1(n7385), .A2(n7390), .ZN(n7340) );
  OAI21_X1 U9106 ( .B1(n7335), .B2(n7334), .A(n7333), .ZN(n7384) );
  OAI22_X1 U9107 ( .A1(n9644), .A2(n7387), .B1(n9910), .B2(n6998), .ZN(n7336)
         );
  AOI21_X1 U9108 ( .B1(n7384), .B2(n9711), .A(n7336), .ZN(n7337) );
  OAI21_X1 U9109 ( .B1(n7340), .B2(n9908), .A(n7337), .ZN(P1_U3528) );
  OAI22_X1 U9110 ( .A1(n9755), .A2(n7387), .B1(n9906), .B2(n5214), .ZN(n7338)
         );
  AOI21_X1 U9111 ( .B1(n7384), .B2(n9786), .A(n7338), .ZN(n7339) );
  OAI21_X1 U9112 ( .B1(n7340), .B2(n9905), .A(n7339), .ZN(P1_U3471) );
  INV_X1 U9113 ( .A(n7341), .ZN(n7342) );
  OAI21_X1 U9114 ( .B1(n7344), .B2(n7343), .A(n7342), .ZN(n7352) );
  INV_X1 U9115 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n7350) );
  NOR2_X1 U9116 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n5304), .ZN(n7888) );
  AOI221_X1 U9117 ( .B1(n7347), .B2(n7346), .C1(n7345), .C2(n7346), .A(n9844), 
        .ZN(n7348) );
  NOR2_X1 U9118 ( .A1(n7888), .A2(n7348), .ZN(n7349) );
  OAI21_X1 U9119 ( .B1(n9875), .B2(n7350), .A(n7349), .ZN(n7351) );
  AOI21_X1 U9120 ( .B1(n9386), .B2(n7352), .A(n7351), .ZN(n7353) );
  OAI21_X1 U9121 ( .B1(n7354), .B2(n9866), .A(n7353), .ZN(P1_U3255) );
  NAND3_X1 U9122 ( .A1(n8217), .A2(n10005), .A3(n7355), .ZN(n7357) );
  OAI211_X1 U9123 ( .C1(n7125), .C2(n9943), .A(n7357), .B(n7356), .ZN(n7358)
         );
  AOI22_X1 U9124 ( .A1(n7358), .A2(n8913), .B1(n8918), .B2(n7535), .ZN(n7359)
         );
  OAI21_X1 U9125 ( .B1(n7360), .B2(n8913), .A(n7359), .ZN(P2_U3233) );
  AOI22_X1 U9126 ( .A1(n9244), .A2(n9261), .B1(n9225), .B2(n9263), .ZN(n7361)
         );
  NAND2_X1 U9127 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_U3086), .ZN(n9856) );
  OAI211_X1 U9128 ( .C1(n7362), .C2(n9247), .A(n7361), .B(n9856), .ZN(n7367)
         );
  AOI211_X1 U9129 ( .C1(n7365), .C2(n7364), .A(n9205), .B(n7363), .ZN(n7366)
         );
  AOI211_X1 U9130 ( .C1(n9229), .C2(n7368), .A(n7367), .B(n7366), .ZN(n7369)
         );
  INV_X1 U9131 ( .A(n7369), .ZN(P1_U3230) );
  INV_X1 U9132 ( .A(n7370), .ZN(n7374) );
  INV_X1 U9133 ( .A(n7371), .ZN(n7372) );
  AOI21_X1 U9134 ( .B1(n7374), .B2(n7373), .A(n7372), .ZN(n9973) );
  NAND3_X1 U9135 ( .A1(n7376), .A2(n8219), .A3(n7377), .ZN(n7378) );
  NAND2_X1 U9136 ( .A1(n7375), .A2(n7378), .ZN(n7379) );
  AOI222_X1 U9137 ( .A1(n8912), .A2(n7379), .B1(n8592), .B2(n8909), .C1(n5755), 
        .C2(n8907), .ZN(n9971) );
  MUX2_X1 U9138 ( .A(n7056), .B(n9971), .S(n8913), .Z(n7383) );
  AOI22_X1 U9139 ( .A1(n8918), .A2(n7381), .B1(n8917), .B2(n7380), .ZN(n7382)
         );
  OAI211_X1 U9140 ( .C1(n8922), .C2(n9973), .A(n7383), .B(n7382), .ZN(P2_U3230) );
  INV_X1 U9141 ( .A(n7384), .ZN(n7393) );
  NAND2_X1 U9142 ( .A1(n7385), .A2(n9560), .ZN(n7392) );
  OAI22_X1 U9143 ( .A1(n9560), .A2(n7386), .B1(n7619), .B2(n9886), .ZN(n7389)
         );
  NOR2_X1 U9144 ( .A1(n9585), .A2(n7387), .ZN(n7388) );
  AOI211_X1 U9145 ( .C1(n7390), .C2(n9578), .A(n7389), .B(n7388), .ZN(n7391)
         );
  OAI211_X1 U9146 ( .C1(n7393), .C2(n9637), .A(n7392), .B(n7391), .ZN(P1_U3287) );
  OAI22_X1 U9147 ( .A1(n9489), .A2(n7395), .B1(n7394), .B2(n9886), .ZN(n7398)
         );
  NOR2_X1 U9148 ( .A1(n9889), .A2(n7396), .ZN(n7397) );
  AOI211_X1 U9149 ( .C1(n9889), .C2(P1_REG2_REG_1__SCAN_IN), .A(n7398), .B(
        n7397), .ZN(n7400) );
  NAND2_X1 U9150 ( .A1(n9560), .A2(n9723), .ZN(n9606) );
  INV_X1 U9151 ( .A(n9606), .ZN(n9555) );
  AOI22_X1 U9152 ( .A1(n9555), .A2(n6414), .B1(n9620), .B2(n4417), .ZN(n7399)
         );
  OAI211_X1 U9153 ( .C1(n7401), .C2(n9637), .A(n7400), .B(n7399), .ZN(P1_U3292) );
  AOI22_X1 U9154 ( .A1(n7403), .A2(n9578), .B1(n9632), .B2(n7402), .ZN(n7404)
         );
  OAI21_X1 U9155 ( .B1(n7405), .B2(n9560), .A(n7404), .ZN(n7408) );
  OAI22_X1 U9156 ( .A1(n9585), .A2(n6440), .B1(n7406), .B2(n9606), .ZN(n7407)
         );
  AOI211_X1 U9157 ( .C1(n9446), .C2(n7409), .A(n7408), .B(n7407), .ZN(n7410)
         );
  OAI21_X1 U9158 ( .B1(n9889), .B2(n7411), .A(n7410), .ZN(P1_U3290) );
  OAI21_X1 U9159 ( .B1(n7414), .B2(n7413), .A(n7412), .ZN(n7456) );
  INV_X1 U9160 ( .A(n7456), .ZN(n7427) );
  INV_X1 U9161 ( .A(n7457), .ZN(n7627) );
  OAI22_X1 U9162 ( .A1(n9585), .A2(n7627), .B1(n7625), .B2(n9886), .ZN(n7417)
         );
  OAI211_X1 U9163 ( .C1(n7415), .C2(n7627), .A(n9628), .B(n7444), .ZN(n7452)
         );
  NOR2_X1 U9164 ( .A1(n7452), .A2(n9489), .ZN(n7416) );
  AOI211_X1 U9165 ( .C1(n9555), .C2(n9260), .A(n7417), .B(n7416), .ZN(n7426)
         );
  INV_X1 U9166 ( .A(n7496), .ZN(n7420) );
  OAI21_X1 U9167 ( .B1(n7420), .B2(n7419), .A(n7418), .ZN(n7421) );
  NAND2_X1 U9168 ( .A1(n7421), .A2(n7422), .ZN(n7586) );
  OAI21_X1 U9169 ( .B1(n7422), .B2(n7421), .A(n7586), .ZN(n7423) );
  AOI22_X1 U9170 ( .A1(n7423), .A2(n9893), .B1(n9881), .B2(n9258), .ZN(n7453)
         );
  MUX2_X1 U9171 ( .A(n7424), .B(n7453), .S(n9560), .Z(n7425) );
  OAI211_X1 U9172 ( .C1(n7427), .C2(n9637), .A(n7426), .B(n7425), .ZN(P1_U3286) );
  INV_X1 U9173 ( .A(n8261), .ZN(n8249) );
  NOR2_X1 U9174 ( .A1(n8270), .A2(n8249), .ZN(n7430) );
  INV_X1 U9175 ( .A(n7428), .ZN(n7429) );
  AOI21_X1 U9176 ( .B1(n7430), .B2(n7371), .A(n7429), .ZN(n9979) );
  XOR2_X1 U9177 ( .A(n7431), .B(n8270), .Z(n7432) );
  AOI222_X1 U9178 ( .A1(n8912), .A2(n7432), .B1(n5772), .B2(n8907), .C1(n8591), 
        .C2(n8909), .ZN(n9977) );
  MUX2_X1 U9179 ( .A(n6317), .B(n9977), .S(n8913), .Z(n7436) );
  AOI22_X1 U9180 ( .A1(n8918), .A2(n7434), .B1(n8917), .B2(n7433), .ZN(n7435)
         );
  OAI211_X1 U9181 ( .C1(n8922), .C2(n9979), .A(n7436), .B(n7435), .ZN(P2_U3229) );
  NAND2_X1 U9182 ( .A1(n7586), .A2(n7437), .ZN(n7438) );
  XNOR2_X1 U9183 ( .A(n7438), .B(n7442), .ZN(n7440) );
  OAI22_X1 U9184 ( .A1(n7440), .A2(n9498), .B1(n7439), .B2(n9591), .ZN(n7604)
         );
  INV_X1 U9185 ( .A(n7604), .ZN(n7451) );
  OAI21_X1 U9186 ( .B1(n7443), .B2(n7442), .A(n7441), .ZN(n7605) );
  OAI211_X1 U9187 ( .C1(n4680), .C2(n4681), .A(n7593), .B(n9628), .ZN(n7602)
         );
  OAI22_X1 U9188 ( .A1(n9560), .A2(n7445), .B1(n7840), .B2(n9886), .ZN(n7447)
         );
  NOR2_X1 U9189 ( .A1(n9606), .A2(n7841), .ZN(n7446) );
  AOI211_X1 U9190 ( .C1(n9620), .C2(n7839), .A(n7447), .B(n7446), .ZN(n7448)
         );
  OAI21_X1 U9191 ( .B1(n9489), .B2(n7602), .A(n7448), .ZN(n7449) );
  AOI21_X1 U9192 ( .B1(n7605), .B2(n9446), .A(n7449), .ZN(n7450) );
  OAI21_X1 U9193 ( .B1(n9889), .B2(n7451), .A(n7450), .ZN(P1_U3285) );
  OAI211_X1 U9194 ( .C1(n7454), .C2(n9705), .A(n7453), .B(n7452), .ZN(n7455)
         );
  AOI21_X1 U9195 ( .B1(n9903), .B2(n7456), .A(n7455), .ZN(n7462) );
  AOI22_X1 U9196 ( .A1(n9734), .A2(n7457), .B1(n9908), .B2(
        P1_REG1_REG_7__SCAN_IN), .ZN(n7458) );
  OAI21_X1 U9197 ( .B1(n7462), .B2(n9908), .A(n7458), .ZN(P1_U3529) );
  INV_X1 U9198 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n7459) );
  OAI22_X1 U9199 ( .A1(n9755), .A2(n7627), .B1(n9906), .B2(n7459), .ZN(n7460)
         );
  INV_X1 U9200 ( .A(n7460), .ZN(n7461) );
  OAI21_X1 U9201 ( .B1(n7462), .B2(n9905), .A(n7461), .ZN(P1_U3474) );
  INV_X1 U9202 ( .A(n7463), .ZN(n7464) );
  XNOR2_X1 U9203 ( .A(n7209), .B(n9984), .ZN(n7571) );
  XNOR2_X1 U9204 ( .A(n7571), .B(n8591), .ZN(n7572) );
  XNOR2_X1 U9205 ( .A(n4511), .B(n7572), .ZN(n7466) );
  NAND2_X1 U9206 ( .A1(n7466), .A2(n8545), .ZN(n7472) );
  INV_X1 U9207 ( .A(n7467), .ZN(n7470) );
  INV_X1 U9208 ( .A(n8590), .ZN(n8277) );
  OAI22_X1 U9209 ( .A1(n8550), .A2(n7468), .B1(n8277), .B2(n8566), .ZN(n7469)
         );
  AOI211_X1 U9210 ( .C1(n7520), .C2(n8576), .A(n7470), .B(n7469), .ZN(n7471)
         );
  OAI211_X1 U9211 ( .C1(n7518), .C2(n8570), .A(n7472), .B(n7471), .ZN(P2_U3167) );
  NAND2_X1 U9212 ( .A1(n9324), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n7475) );
  OAI21_X1 U9213 ( .B1(n9324), .B2(P1_REG2_REG_14__SCAN_IN), .A(n7475), .ZN(
        n7476) );
  AOI211_X1 U9214 ( .C1(n7477), .C2(n7476), .A(n9323), .B(n9844), .ZN(n7486)
         );
  XNOR2_X1 U9215 ( .A(n9331), .B(P1_REG1_REG_14__SCAN_IN), .ZN(n7482) );
  OAI21_X1 U9216 ( .B1(n7480), .B2(n7479), .A(n7478), .ZN(n7481) );
  NAND2_X1 U9217 ( .A1(n7482), .A2(n7481), .ZN(n9330) );
  OAI211_X1 U9218 ( .C1(n7482), .C2(n7481), .A(n9386), .B(n9330), .ZN(n7484)
         );
  AND2_X1 U9219 ( .A1(P1_U3086), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n9055) );
  AOI21_X1 U9220 ( .B1(n9352), .B2(P1_ADDR_REG_14__SCAN_IN), .A(n9055), .ZN(
        n7483) );
  OAI211_X1 U9221 ( .C1(n9866), .C2(n9331), .A(n7484), .B(n7483), .ZN(n7485)
         );
  OR2_X1 U9222 ( .A1(n7486), .A2(n7485), .ZN(P1_U3257) );
  OAI21_X1 U9223 ( .B1(n7489), .B2(n7488), .A(n7487), .ZN(n9904) );
  INV_X1 U9224 ( .A(n7490), .ZN(n7492) );
  AOI211_X1 U9225 ( .C1(n7493), .C2(n7492), .A(n9567), .B(n7491), .ZN(n9897)
         );
  INV_X1 U9226 ( .A(n7494), .ZN(n7528) );
  AOI22_X1 U9227 ( .A1(n9897), .A2(n9578), .B1(n7528), .B2(n9632), .ZN(n7495)
         );
  OAI21_X1 U9228 ( .B1(n9900), .B2(n9585), .A(n7495), .ZN(n7502) );
  OAI211_X1 U9229 ( .C1(n7498), .C2(n7497), .A(n7496), .B(n9893), .ZN(n7500)
         );
  AOI22_X1 U9230 ( .A1(n9881), .A2(n9260), .B1(n9723), .B2(n9262), .ZN(n7499)
         );
  NAND2_X1 U9231 ( .A1(n7500), .A2(n7499), .ZN(n9902) );
  MUX2_X1 U9232 ( .A(n9902), .B(P1_REG2_REG_5__SCAN_IN), .S(n9889), .Z(n7501)
         );
  AOI211_X1 U9233 ( .C1(n9446), .C2(n9904), .A(n7502), .B(n7501), .ZN(n7503)
         );
  INV_X1 U9234 ( .A(n7503), .ZN(P1_U3288) );
  AOI21_X1 U9235 ( .B1(P1_REG3_REG_2__SCAN_IN), .B2(n9632), .A(n7504), .ZN(
        n7510) );
  AOI22_X1 U9236 ( .A1(P1_REG2_REG_2__SCAN_IN), .A2(n9889), .B1(n9578), .B2(
        n7505), .ZN(n7506) );
  OAI21_X1 U9237 ( .B1(n9585), .B2(n6411), .A(n7506), .ZN(n7507) );
  AOI21_X1 U9238 ( .B1(n9446), .B2(n7508), .A(n7507), .ZN(n7509) );
  OAI21_X1 U9239 ( .B1(n9889), .B2(n7510), .A(n7509), .ZN(P1_U3291) );
  INV_X1 U9240 ( .A(n7511), .ZN(n7513) );
  NOR2_X1 U9241 ( .A1(n7513), .A2(n7512), .ZN(n8222) );
  XNOR2_X1 U9242 ( .A(n7514), .B(n8222), .ZN(n9985) );
  XOR2_X1 U9243 ( .A(n8222), .B(n7515), .Z(n7516) );
  AOI222_X1 U9244 ( .A1(n8912), .A2(n7516), .B1(n8590), .B2(n8909), .C1(n8592), 
        .C2(n8907), .ZN(n9983) );
  MUX2_X1 U9245 ( .A(n7517), .B(n9983), .S(n8913), .Z(n7522) );
  INV_X1 U9246 ( .A(n7518), .ZN(n7519) );
  AOI22_X1 U9247 ( .A1(n8918), .A2(n7520), .B1(n8917), .B2(n7519), .ZN(n7521)
         );
  OAI211_X1 U9248 ( .C1(n8922), .C2(n9985), .A(n7522), .B(n7521), .ZN(P2_U3228) );
  NOR2_X1 U9249 ( .A1(n7523), .A2(n4513), .ZN(n7525) );
  XNOR2_X1 U9250 ( .A(n7525), .B(n7524), .ZN(n7530) );
  AOI22_X1 U9251 ( .A1(n9244), .A2(n9260), .B1(n9225), .B2(n9262), .ZN(n7526)
         );
  NAND2_X1 U9252 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n9265) );
  OAI211_X1 U9253 ( .C1(n9900), .C2(n9247), .A(n7526), .B(n9265), .ZN(n7527)
         );
  AOI21_X1 U9254 ( .B1(n7528), .B2(n9229), .A(n7527), .ZN(n7529) );
  OAI21_X1 U9255 ( .B1(n7530), .B2(n9205), .A(n7529), .ZN(P1_U3227) );
  XNOR2_X1 U9256 ( .A(n7531), .B(n7532), .ZN(n9964) );
  OAI22_X1 U9257 ( .A1(n8846), .A2(n9961), .B1(n7533), .B2(n9943), .ZN(n7542)
         );
  NAND2_X1 U9258 ( .A1(n7535), .A2(n8912), .ZN(n7536) );
  OAI21_X1 U9259 ( .B1(n7531), .B2(n7536), .A(n9951), .ZN(n7538) );
  NAND2_X1 U9260 ( .A1(n7538), .A2(n7537), .ZN(n7540) );
  NAND2_X1 U9261 ( .A1(n5755), .A2(n8909), .ZN(n7539) );
  OAI211_X1 U9262 ( .C1(n7534), .C2(n9949), .A(n7540), .B(n7539), .ZN(n9962)
         );
  MUX2_X1 U9263 ( .A(n9962), .B(P2_REG2_REG_1__SCAN_IN), .S(n9960), .Z(n7541)
         );
  AOI211_X1 U9264 ( .C1(n8848), .C2(n9964), .A(n7542), .B(n7541), .ZN(n7543)
         );
  INV_X1 U9265 ( .A(n7543), .ZN(P2_U3232) );
  INV_X1 U9266 ( .A(n7544), .ZN(n7547) );
  OAI222_X1 U9267 ( .A1(n8437), .A2(n7546), .B1(n8435), .B2(n7547), .C1(n7545), 
        .C2(P2_U3151), .ZN(P2_U3276) );
  OAI222_X1 U9268 ( .A1(n9824), .A2(n7548), .B1(n9822), .B2(n7547), .C1(
        P1_U3086), .C2(n4519), .ZN(P1_U3336) );
  OAI211_X1 U9269 ( .C1(n7550), .C2(n7553), .A(n7549), .B(n8912), .ZN(n7552)
         );
  AOI22_X1 U9270 ( .A1(n8909), .A2(n8588), .B1(n8590), .B2(n8907), .ZN(n7551)
         );
  NAND2_X1 U9271 ( .A1(n7552), .A2(n7551), .ZN(n7641) );
  INV_X1 U9272 ( .A(n7641), .ZN(n7559) );
  XNOR2_X1 U9273 ( .A(n7554), .B(n7553), .ZN(n7642) );
  INV_X1 U9274 ( .A(n7555), .ZN(n7675) );
  AOI22_X1 U9275 ( .A1(n9960), .A2(P2_REG2_REG_7__SCAN_IN), .B1(n8917), .B2(
        n7675), .ZN(n7556) );
  OAI21_X1 U9276 ( .B1(n8304), .B2(n8846), .A(n7556), .ZN(n7557) );
  AOI21_X1 U9277 ( .B1(n7642), .B2(n8848), .A(n7557), .ZN(n7558) );
  OAI21_X1 U9278 ( .B1(n7559), .B2(n9960), .A(n7558), .ZN(P2_U3226) );
  NAND2_X1 U9279 ( .A1(n7560), .A2(n8285), .ZN(n7564) );
  INV_X1 U9280 ( .A(n7561), .ZN(n7562) );
  XNOR2_X1 U9281 ( .A(n7564), .B(n4441), .ZN(n9991) );
  INV_X1 U9282 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n7567) );
  XNOR2_X1 U9283 ( .A(n7565), .B(n4441), .ZN(n7566) );
  AOI222_X1 U9284 ( .A1(n8912), .A2(n7566), .B1(n8589), .B2(n8909), .C1(n8591), 
        .C2(n8907), .ZN(n9989) );
  MUX2_X1 U9285 ( .A(n7567), .B(n9989), .S(n8913), .Z(n7570) );
  INV_X1 U9286 ( .A(n7582), .ZN(n7568) );
  AOI22_X1 U9287 ( .A1(n8918), .A2(n8278), .B1(n8917), .B2(n7568), .ZN(n7569)
         );
  OAI211_X1 U9288 ( .C1(n8922), .C2(n9991), .A(n7570), .B(n7569), .ZN(P2_U3227) );
  XNOR2_X1 U9289 ( .A(n8186), .B(n9990), .ZN(n7668) );
  XNOR2_X1 U9290 ( .A(n7668), .B(n8590), .ZN(n7574) );
  AOI211_X1 U9291 ( .C1(n7574), .C2(n7573), .A(n8571), .B(n7670), .ZN(n7575)
         );
  INV_X1 U9292 ( .A(n7575), .ZN(n7581) );
  INV_X1 U9293 ( .A(n7576), .ZN(n7579) );
  INV_X1 U9294 ( .A(n8589), .ZN(n7577) );
  OAI22_X1 U9295 ( .A1(n8550), .A2(n4972), .B1(n7577), .B2(n8566), .ZN(n7578)
         );
  AOI211_X1 U9296 ( .C1(n8278), .C2(n8576), .A(n7579), .B(n7578), .ZN(n7580)
         );
  OAI211_X1 U9297 ( .C1(n7582), .C2(n8570), .A(n7581), .B(n7580), .ZN(P2_U3179) );
  INV_X1 U9298 ( .A(n7583), .ZN(n7584) );
  AOI21_X1 U9299 ( .B1(n7586), .B2(n7585), .A(n7584), .ZN(n7587) );
  XNOR2_X1 U9300 ( .A(n7587), .B(n7591), .ZN(n7589) );
  OAI22_X1 U9301 ( .A1(n7589), .A2(n9498), .B1(n7588), .B2(n9705), .ZN(n7633)
         );
  INV_X1 U9302 ( .A(n7633), .ZN(n7601) );
  OAI21_X1 U9303 ( .B1(n7592), .B2(n7591), .A(n7590), .ZN(n7634) );
  INV_X1 U9304 ( .A(n9173), .ZN(n7636) );
  INV_X1 U9305 ( .A(n7593), .ZN(n7594) );
  OAI21_X1 U9306 ( .B1(n7594), .B2(n7636), .A(n9628), .ZN(n7595) );
  OAI22_X1 U9307 ( .A1(n7595), .A2(n7744), .B1(n7830), .B2(n9591), .ZN(n7632)
         );
  AND2_X1 U9308 ( .A1(n9560), .A2(n4519), .ZN(n9615) );
  NAND2_X1 U9309 ( .A1(n7632), .A2(n9615), .ZN(n7598) );
  INV_X1 U9310 ( .A(n7596), .ZN(n9160) );
  AOI22_X1 U9311 ( .A1(n9889), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n9160), .B2(
        n9632), .ZN(n7597) );
  OAI211_X1 U9312 ( .C1(n7636), .C2(n9585), .A(n7598), .B(n7597), .ZN(n7599)
         );
  AOI21_X1 U9313 ( .B1(n7634), .B2(n9446), .A(n7599), .ZN(n7600) );
  OAI21_X1 U9314 ( .B1(n9889), .B2(n7601), .A(n7600), .ZN(P1_U3284) );
  OAI21_X1 U9315 ( .B1(n7841), .B2(n9705), .A(n7602), .ZN(n7603) );
  AOI211_X1 U9316 ( .C1(n7605), .C2(n9903), .A(n7604), .B(n7603), .ZN(n7608)
         );
  AOI22_X1 U9317 ( .A1(n9734), .A2(n7839), .B1(n9908), .B2(
        P1_REG1_REG_8__SCAN_IN), .ZN(n7606) );
  OAI21_X1 U9318 ( .B1(n7608), .B2(n9908), .A(n7606), .ZN(P1_U3530) );
  AOI22_X1 U9319 ( .A1(n5657), .A2(n7839), .B1(n9905), .B2(
        P1_REG0_REG_8__SCAN_IN), .ZN(n7607) );
  OAI21_X1 U9320 ( .B1(n7608), .B2(n9905), .A(n7607), .ZN(P1_U3477) );
  XNOR2_X1 U9321 ( .A(n7611), .B(n7610), .ZN(n7612) );
  XNOR2_X1 U9322 ( .A(n7609), .B(n7612), .ZN(n7613) );
  NAND2_X1 U9323 ( .A1(n7613), .A2(n9236), .ZN(n7618) );
  AND2_X1 U9324 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n9280) );
  OAI22_X1 U9325 ( .A1(n9241), .A2(n7614), .B1(n7841), .B2(n9227), .ZN(n7615)
         );
  AOI211_X1 U9326 ( .C1(n7616), .C2(n9209), .A(n9280), .B(n7615), .ZN(n7617)
         );
  OAI211_X1 U9327 ( .C1(n9239), .C2(n7619), .A(n7618), .B(n7617), .ZN(P1_U3239) );
  INV_X1 U9328 ( .A(n7620), .ZN(n7621) );
  NOR2_X1 U9329 ( .A1(n7622), .A2(n7621), .ZN(n7623) );
  XNOR2_X1 U9330 ( .A(n7624), .B(n7623), .ZN(n7631) );
  INV_X1 U9331 ( .A(n7625), .ZN(n7629) );
  AOI22_X1 U9332 ( .A1(n9244), .A2(n9258), .B1(n9225), .B2(n9260), .ZN(n7626)
         );
  NAND2_X1 U9333 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3086), .ZN(n9293) );
  OAI211_X1 U9334 ( .C1(n7627), .C2(n9247), .A(n7626), .B(n9293), .ZN(n7628)
         );
  AOI21_X1 U9335 ( .B1(n7629), .B2(n9229), .A(n7628), .ZN(n7630) );
  OAI21_X1 U9336 ( .B1(n7631), .B2(n9205), .A(n7630), .ZN(P1_U3213) );
  AOI211_X1 U9337 ( .C1(n7634), .C2(n9903), .A(n7633), .B(n7632), .ZN(n7640)
         );
  INV_X1 U9338 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n7635) );
  OAI22_X1 U9339 ( .A1(n9755), .A2(n7636), .B1(n9906), .B2(n7635), .ZN(n7637)
         );
  INV_X1 U9340 ( .A(n7637), .ZN(n7638) );
  OAI21_X1 U9341 ( .B1(n7640), .B2(n9905), .A(n7638), .ZN(P1_U3480) );
  AOI22_X1 U9342 ( .A1(n9734), .A2(n9173), .B1(n9908), .B2(
        P1_REG1_REG_9__SCAN_IN), .ZN(n7639) );
  OAI21_X1 U9343 ( .B1(n7640), .B2(n9908), .A(n7639), .ZN(P1_U3531) );
  AOI21_X1 U9344 ( .B1(n7642), .B2(n9970), .A(n7641), .ZN(n7647) );
  INV_X1 U9345 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n7643) );
  OAI22_X1 U9346 ( .A1(n9013), .A2(n8304), .B1(n7643), .B2(n10016), .ZN(n7644)
         );
  INV_X1 U9347 ( .A(n7644), .ZN(n7645) );
  OAI21_X1 U9348 ( .B1(n7647), .B2(n10017), .A(n7645), .ZN(P2_U3411) );
  AOI22_X1 U9349 ( .A1(n8966), .A2(n7676), .B1(n10027), .B2(
        P2_REG1_REG_7__SCAN_IN), .ZN(n7646) );
  OAI21_X1 U9350 ( .B1(n7647), .B2(n10027), .A(n7646), .ZN(P2_U3466) );
  INV_X1 U9351 ( .A(n7648), .ZN(n7666) );
  OAI222_X1 U9352 ( .A1(n8435), .A2(n7666), .B1(P2_U3151), .B2(n6195), .C1(
        n7649), .C2(n8437), .ZN(P2_U3275) );
  AOI21_X1 U9353 ( .B1(n7651), .B2(n5836), .A(n7650), .ZN(n7664) );
  OAI21_X1 U9354 ( .B1(n7654), .B2(n7653), .A(n7652), .ZN(n7662) );
  INV_X1 U9355 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n10317) );
  AND2_X1 U9356 ( .A1(P2_U3151), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n7793) );
  AOI21_X1 U9357 ( .B1(n8709), .B2(n7655), .A(n7793), .ZN(n7656) );
  OAI21_X1 U9358 ( .B1(n10317), .B2(n8735), .A(n7656), .ZN(n7661) );
  AOI21_X1 U9359 ( .B1(n5841), .B2(n7658), .A(n7657), .ZN(n7659) );
  NOR2_X1 U9360 ( .A1(n7659), .A2(n9930), .ZN(n7660) );
  AOI211_X1 U9361 ( .C1(n9918), .C2(n7662), .A(n7661), .B(n7660), .ZN(n7663)
         );
  OAI21_X1 U9362 ( .B1(n7664), .B2(n9929), .A(n7663), .ZN(P2_U3191) );
  INV_X1 U9363 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7665) );
  OAI222_X1 U9364 ( .A1(P1_U3086), .A2(n7667), .B1(n9822), .B2(n7666), .C1(
        n7665), .C2(n9824), .ZN(P1_U3335) );
  XNOR2_X1 U9365 ( .A(n8186), .B(n7676), .ZN(n7777) );
  XNOR2_X1 U9366 ( .A(n7777), .B(n8589), .ZN(n7671) );
  OAI21_X1 U9367 ( .B1(n7672), .B2(n7671), .A(n7779), .ZN(n7682) );
  INV_X1 U9368 ( .A(n7673), .ZN(n7674) );
  AOI21_X1 U9369 ( .B1(n8568), .B2(n8590), .A(n7674), .ZN(n7680) );
  NAND2_X1 U9370 ( .A1(n8558), .A2(n7675), .ZN(n7679) );
  NAND2_X1 U9371 ( .A1(n8576), .A2(n7676), .ZN(n7678) );
  INV_X1 U9372 ( .A(n8588), .ZN(n7804) );
  OR2_X1 U9373 ( .A1(n8566), .A2(n7804), .ZN(n7677) );
  NAND4_X1 U9374 ( .A1(n7680), .A2(n7679), .A3(n7678), .A4(n7677), .ZN(n7681)
         );
  AOI21_X1 U9375 ( .B1(n7682), .B2(n8545), .A(n7681), .ZN(n7683) );
  INV_X1 U9376 ( .A(n7683), .ZN(P2_U3153) );
  XOR2_X1 U9377 ( .A(n8221), .B(n7684), .Z(n9995) );
  OAI211_X1 U9378 ( .C1(n7686), .C2(n8221), .A(n7685), .B(n8912), .ZN(n7688)
         );
  AOI22_X1 U9379 ( .A1(n8587), .A2(n8909), .B1(n8907), .B2(n8589), .ZN(n7687)
         );
  AND2_X1 U9380 ( .A1(n7688), .A2(n7687), .ZN(n9996) );
  MUX2_X1 U9381 ( .A(n9996), .B(n7689), .S(n9960), .Z(n7692) );
  INV_X1 U9382 ( .A(n7690), .ZN(n7781) );
  AOI22_X1 U9383 ( .A1(n8918), .A2(n7785), .B1(n8917), .B2(n7781), .ZN(n7691)
         );
  OAI211_X1 U9384 ( .C1(n8922), .C2(n9995), .A(n7692), .B(n7691), .ZN(P2_U3225) );
  INV_X1 U9385 ( .A(n7693), .ZN(n7733) );
  OAI222_X1 U9386 ( .A1(n8435), .A2(n7733), .B1(P2_U3151), .B2(n7199), .C1(
        n7694), .C2(n8437), .ZN(P2_U3274) );
  INV_X1 U9387 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n10099) );
  INV_X1 U9388 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n8704) );
  INV_X1 U9389 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n10181) );
  NOR2_X1 U9390 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n7727) );
  NOR2_X1 U9391 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n7724) );
  NOR2_X1 U9392 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n7721) );
  NOR2_X1 U9393 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n7718) );
  NOR2_X1 U9394 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n10318) );
  INV_X1 U9395 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n7935) );
  NOR2_X1 U9396 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n7713) );
  NOR2_X1 U9397 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n7710) );
  NOR2_X1 U9398 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n7708) );
  NOR2_X1 U9399 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n7706) );
  NOR2_X1 U9400 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n7704) );
  NOR2_X1 U9401 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n10278) );
  NOR2_X1 U9402 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n7701) );
  NAND2_X1 U9403 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n7699) );
  XOR2_X1 U9404 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(P2_ADDR_REG_3__SCAN_IN), .Z(
        n10370) );
  NAND2_X1 U9405 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n7697) );
  AOI21_X1 U9406 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(P2_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10030) );
  INV_X1 U9407 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n10034) );
  NOR2_X1 U9408 ( .A1(n6968), .A2(n10034), .ZN(n10033) );
  AND2_X1 U9409 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(n10033), .ZN(n10031) );
  NOR2_X1 U9410 ( .A1(P2_ADDR_REG_1__SCAN_IN), .A2(n10031), .ZN(n7695) );
  NOR2_X1 U9411 ( .A1(n10030), .A2(n7695), .ZN(n10368) );
  XOR2_X1 U9412 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(P2_ADDR_REG_2__SCAN_IN), .Z(
        n10367) );
  NAND2_X1 U9413 ( .A1(n10368), .A2(n10367), .ZN(n7696) );
  NAND2_X1 U9414 ( .A1(n7697), .A2(n7696), .ZN(n10369) );
  NAND2_X1 U9415 ( .A1(n10370), .A2(n10369), .ZN(n7698) );
  NAND2_X1 U9416 ( .A1(n7699), .A2(n7698), .ZN(n10372) );
  XOR2_X1 U9417 ( .A(n9858), .B(P2_ADDR_REG_4__SCAN_IN), .Z(n10371) );
  NOR2_X1 U9418 ( .A1(n10372), .A2(n10371), .ZN(n7700) );
  NOR2_X1 U9419 ( .A1(n7701), .A2(n7700), .ZN(n10360) );
  XOR2_X1 U9420 ( .A(n10126), .B(P1_ADDR_REG_5__SCAN_IN), .Z(n10359) );
  NOR2_X1 U9421 ( .A1(n10360), .A2(n10359), .ZN(n7702) );
  NOR2_X1 U9422 ( .A1(n10278), .A2(n7702), .ZN(n10358) );
  INV_X1 U9423 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n10065) );
  XOR2_X1 U9424 ( .A(n10065), .B(P1_ADDR_REG_6__SCAN_IN), .Z(n10357) );
  NOR2_X1 U9425 ( .A1(n10358), .A2(n10357), .ZN(n7703) );
  NOR2_X1 U9426 ( .A1(n7704), .A2(n7703), .ZN(n10364) );
  XNOR2_X1 U9427 ( .A(P2_ADDR_REG_7__SCAN_IN), .B(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n10363) );
  NOR2_X1 U9428 ( .A1(n10364), .A2(n10363), .ZN(n7705) );
  NOR2_X1 U9429 ( .A1(n7706), .A2(n7705), .ZN(n10366) );
  XNOR2_X1 U9430 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n10365) );
  NOR2_X1 U9431 ( .A1(n10366), .A2(n10365), .ZN(n7707) );
  NOR2_X1 U9432 ( .A1(n7708), .A2(n7707), .ZN(n10362) );
  INV_X1 U9433 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n9838) );
  AOI22_X1 U9434 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n9838), .B1(
        P1_ADDR_REG_9__SCAN_IN), .B2(n10317), .ZN(n10361) );
  NOR2_X1 U9435 ( .A1(n10362), .A2(n10361), .ZN(n7709) );
  NOR2_X1 U9436 ( .A1(n7710), .A2(n7709), .ZN(n10053) );
  INV_X1 U9437 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n7711) );
  INV_X1 U9438 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n7768) );
  AOI22_X1 U9439 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(n7711), .B1(
        P1_ADDR_REG_10__SCAN_IN), .B2(n7768), .ZN(n10052) );
  NOR2_X1 U9440 ( .A1(n10053), .A2(n10052), .ZN(n7712) );
  NOR2_X1 U9441 ( .A1(n7713), .A2(n7712), .ZN(n10051) );
  AOI22_X1 U9442 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(n10339), .B1(
        P1_ADDR_REG_11__SCAN_IN), .B2(n7935), .ZN(n10050) );
  NOR2_X1 U9443 ( .A1(n10051), .A2(n10050), .ZN(n7714) );
  AOI21_X1 U9444 ( .B1(n7935), .B2(n10339), .A(n7714), .ZN(n10049) );
  INV_X1 U9445 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n10071) );
  AOI22_X1 U9446 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(n7350), .B1(
        P1_ADDR_REG_12__SCAN_IN), .B2(n10071), .ZN(n10048) );
  NOR2_X1 U9447 ( .A1(n10049), .A2(n10048), .ZN(n7715) );
  NOR2_X1 U9448 ( .A1(n10318), .A2(n7715), .ZN(n10047) );
  INV_X1 U9449 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n7716) );
  INV_X1 U9450 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n8645) );
  AOI22_X1 U9451 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(n7716), .B1(
        P1_ADDR_REG_13__SCAN_IN), .B2(n8645), .ZN(n10046) );
  NOR2_X1 U9452 ( .A1(n10047), .A2(n10046), .ZN(n7717) );
  NOR2_X1 U9453 ( .A1(n7718), .A2(n7717), .ZN(n10045) );
  INV_X1 U9454 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n7719) );
  INV_X1 U9455 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n10342) );
  AOI22_X1 U9456 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(n7719), .B1(
        P1_ADDR_REG_14__SCAN_IN), .B2(n10342), .ZN(n10044) );
  NOR2_X1 U9457 ( .A1(n10045), .A2(n10044), .ZN(n7720) );
  NOR2_X1 U9458 ( .A1(n7721), .A2(n7720), .ZN(n10043) );
  INV_X1 U9459 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n7722) );
  INV_X1 U9460 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n8677) );
  AOI22_X1 U9461 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(n7722), .B1(
        P1_ADDR_REG_15__SCAN_IN), .B2(n8677), .ZN(n10042) );
  NOR2_X1 U9462 ( .A1(n10043), .A2(n10042), .ZN(n7723) );
  NOR2_X1 U9463 ( .A1(n7724), .A2(n7723), .ZN(n10041) );
  INV_X1 U9464 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n7725) );
  INV_X1 U9465 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n8691) );
  AOI22_X1 U9466 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(n7725), .B1(
        P1_ADDR_REG_16__SCAN_IN), .B2(n8691), .ZN(n10040) );
  NOR2_X1 U9467 ( .A1(n10041), .A2(n10040), .ZN(n7726) );
  NOR2_X1 U9468 ( .A1(n7727), .A2(n7726), .ZN(n10039) );
  AOI22_X1 U9469 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(n10181), .B1(
        P1_ADDR_REG_17__SCAN_IN), .B2(n8704), .ZN(n10038) );
  NOR2_X1 U9470 ( .A1(n10039), .A2(n10038), .ZN(n7728) );
  AOI21_X1 U9471 ( .B1(n8704), .B2(n10181), .A(n7728), .ZN(n10036) );
  NOR2_X1 U9472 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n10036), .ZN(n7729) );
  NAND2_X1 U9473 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n10036), .ZN(n10035) );
  OAI21_X1 U9474 ( .B1(n10099), .B2(n7729), .A(n10035), .ZN(n7731) );
  XNOR2_X1 U9475 ( .A(P1_ADDR_REG_19__SCAN_IN), .B(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n7730) );
  XNOR2_X1 U9476 ( .A(n7731), .B(n7730), .ZN(ADD_1068_U4) );
  OAI222_X1 U9477 ( .A1(n9824), .A2(n7734), .B1(n9822), .B2(n7733), .C1(n7732), 
        .C2(P1_U3086), .ZN(P1_U3334) );
  OAI21_X1 U9478 ( .B1(n7737), .B2(n7736), .A(n7735), .ZN(n7752) );
  INV_X1 U9479 ( .A(n7752), .ZN(n7751) );
  INV_X1 U9480 ( .A(n9711), .ZN(n9736) );
  AND2_X1 U9481 ( .A1(n7739), .A2(n7738), .ZN(n7742) );
  OAI21_X1 U9482 ( .B1(n7742), .B2(n7741), .A(n7740), .ZN(n7743) );
  AOI222_X1 U9483 ( .A1(n9893), .A2(n7743), .B1(n9257), .B2(n9723), .C1(n9255), 
        .C2(n9881), .ZN(n7759) );
  OAI211_X1 U9484 ( .C1(n7744), .C2(n7915), .A(n9628), .B(n7821), .ZN(n7753)
         );
  NAND2_X1 U9485 ( .A1(n7759), .A2(n7753), .ZN(n7749) );
  OAI22_X1 U9486 ( .A1(n9644), .A2(n7915), .B1(n9910), .B2(n7007), .ZN(n7745)
         );
  AOI21_X1 U9487 ( .B1(n7749), .B2(n9910), .A(n7745), .ZN(n7746) );
  OAI21_X1 U9488 ( .B1(n7751), .B2(n9736), .A(n7746), .ZN(P1_U3532) );
  INV_X1 U9489 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n7747) );
  OAI22_X1 U9490 ( .A1(n9755), .A2(n7915), .B1(n9906), .B2(n7747), .ZN(n7748)
         );
  AOI21_X1 U9491 ( .B1(n7749), .B2(n9906), .A(n7748), .ZN(n7750) );
  OAI21_X1 U9492 ( .B1(n7751), .B2(n9803), .A(n7750), .ZN(P1_U3483) );
  NAND2_X1 U9493 ( .A1(n7752), .A2(n9446), .ZN(n7758) );
  OAI22_X1 U9494 ( .A1(n9560), .A2(n5271), .B1(n7914), .B2(n9886), .ZN(n7755)
         );
  NOR2_X1 U9495 ( .A1(n7753), .A2(n9489), .ZN(n7754) );
  AOI211_X1 U9496 ( .C1(n9620), .C2(n7756), .A(n7755), .B(n7754), .ZN(n7757)
         );
  OAI211_X1 U9497 ( .C1(n9889), .C2(n7759), .A(n7758), .B(n7757), .ZN(P1_U3283) );
  AOI21_X1 U9498 ( .B1(n4512), .B2(n7761), .A(n7760), .ZN(n7776) );
  OAI21_X1 U9499 ( .B1(n7764), .B2(n7763), .A(n7762), .ZN(n7774) );
  INV_X1 U9500 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n7765) );
  NOR2_X1 U9501 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7765), .ZN(n7997) );
  AOI21_X1 U9502 ( .B1(n8709), .B2(n7766), .A(n7997), .ZN(n7767) );
  OAI21_X1 U9503 ( .B1(n7768), .B2(n8735), .A(n7767), .ZN(n7773) );
  AOI21_X1 U9504 ( .B1(n4514), .B2(n7770), .A(n7769), .ZN(n7771) );
  NOR2_X1 U9505 ( .A1(n7771), .A2(n9929), .ZN(n7772) );
  AOI211_X1 U9506 ( .C1(n9918), .C2(n7774), .A(n7773), .B(n7772), .ZN(n7775)
         );
  OAI21_X1 U9507 ( .B1(n7776), .B2(n9930), .A(n7775), .ZN(P2_U3192) );
  NAND2_X1 U9508 ( .A1(n7777), .A2(n7577), .ZN(n7778) );
  XNOR2_X1 U9509 ( .A(n8186), .B(n7785), .ZN(n7788) );
  XNOR2_X1 U9510 ( .A(n7788), .B(n8588), .ZN(n7789) );
  XOR2_X1 U9511 ( .A(n7790), .B(n7789), .Z(n7787) );
  NAND2_X1 U9512 ( .A1(P2_U3151), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n8597) );
  INV_X1 U9513 ( .A(n8597), .ZN(n7780) );
  AOI21_X1 U9514 ( .B1(n8568), .B2(n8589), .A(n7780), .ZN(n7783) );
  NAND2_X1 U9515 ( .A1(n8558), .A2(n7781), .ZN(n7782) );
  OAI211_X1 U9516 ( .C1(n7991), .C2(n8566), .A(n7783), .B(n7782), .ZN(n7784)
         );
  AOI21_X1 U9517 ( .B1(n7785), .B2(n8576), .A(n7784), .ZN(n7786) );
  OAI21_X1 U9518 ( .B1(n7787), .B2(n8571), .A(n7786), .ZN(P2_U3161) );
  XNOR2_X1 U9519 ( .A(n8186), .B(n7950), .ZN(n7990) );
  XNOR2_X1 U9520 ( .A(n7990), .B(n8587), .ZN(n7791) );
  NAND2_X1 U9521 ( .A1(n7792), .A2(n7791), .ZN(n7994) );
  OAI211_X1 U9522 ( .C1(n7792), .C2(n7791), .A(n7994), .B(n8545), .ZN(n7800)
         );
  INV_X1 U9523 ( .A(n7807), .ZN(n7798) );
  INV_X1 U9524 ( .A(n7950), .ZN(n7806) );
  NOR2_X1 U9525 ( .A1(n8554), .A2(n7806), .ZN(n7797) );
  NAND2_X1 U9526 ( .A1(n8568), .A2(n8588), .ZN(n7795) );
  INV_X1 U9527 ( .A(n7793), .ZN(n7794) );
  OAI211_X1 U9528 ( .C1(n8566), .C2(n8006), .A(n7795), .B(n7794), .ZN(n7796)
         );
  AOI211_X1 U9529 ( .C1(n7798), .C2(n8558), .A(n7797), .B(n7796), .ZN(n7799)
         );
  NAND2_X1 U9530 ( .A1(n7800), .A2(n7799), .ZN(P2_U3171) );
  OR2_X1 U9531 ( .A1(n7801), .A2(n8225), .ZN(n7900) );
  INV_X1 U9532 ( .A(n7900), .ZN(n7802) );
  AOI21_X1 U9533 ( .B1(n8225), .B2(n7801), .A(n7802), .ZN(n7803) );
  OAI222_X1 U9534 ( .A1(n9951), .A2(n7804), .B1(n9953), .B2(n8006), .C1(n9949), 
        .C2(n7803), .ZN(n7947) );
  INV_X1 U9535 ( .A(n7947), .ZN(n7811) );
  XNOR2_X1 U9536 ( .A(n7805), .B(n8225), .ZN(n7948) );
  NOR2_X1 U9537 ( .A1(n8846), .A2(n7806), .ZN(n7809) );
  OAI22_X1 U9538 ( .A1(n8913), .A2(n5836), .B1(n7807), .B2(n9943), .ZN(n7808)
         );
  AOI211_X1 U9539 ( .C1(n7948), .C2(n8848), .A(n7809), .B(n7808), .ZN(n7810)
         );
  OAI21_X1 U9540 ( .B1(n7811), .B2(n9960), .A(n7810), .ZN(P2_U3224) );
  NAND2_X1 U9541 ( .A1(n7740), .A2(n7812), .ZN(n7814) );
  XNOR2_X1 U9542 ( .A(n7814), .B(n7813), .ZN(n7815) );
  AOI22_X1 U9543 ( .A1(n7815), .A2(n9893), .B1(n9881), .B2(n9254), .ZN(n7829)
         );
  OAI21_X1 U9544 ( .B1(n7818), .B2(n7817), .A(n7816), .ZN(n7832) );
  NAND2_X1 U9545 ( .A1(n7832), .A2(n9446), .ZN(n7827) );
  INV_X1 U9546 ( .A(n7819), .ZN(n9194) );
  AOI22_X1 U9547 ( .A1(n9889), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n9194), .B2(
        n9632), .ZN(n7820) );
  OAI21_X1 U9548 ( .B1(n7830), .B2(n9606), .A(n7820), .ZN(n7825) );
  INV_X1 U9549 ( .A(n7821), .ZN(n7823) );
  INV_X1 U9550 ( .A(n9210), .ZN(n7822) );
  OAI211_X1 U9551 ( .C1(n7823), .C2(n7822), .A(n9628), .B(n7858), .ZN(n7828)
         );
  NOR2_X1 U9552 ( .A1(n7828), .A2(n9489), .ZN(n7824) );
  AOI211_X1 U9553 ( .C1(n9620), .C2(n9210), .A(n7825), .B(n7824), .ZN(n7826)
         );
  OAI211_X1 U9554 ( .C1(n9889), .C2(n7829), .A(n7827), .B(n7826), .ZN(P1_U3282) );
  OAI211_X1 U9555 ( .C1(n7830), .C2(n9705), .A(n7829), .B(n7828), .ZN(n7831)
         );
  AOI21_X1 U9556 ( .B1(n7832), .B2(n9903), .A(n7831), .ZN(n7835) );
  AOI22_X1 U9557 ( .A1(n5657), .A2(n9210), .B1(n9905), .B2(
        P1_REG0_REG_11__SCAN_IN), .ZN(n7833) );
  OAI21_X1 U9558 ( .B1(n7835), .B2(n9905), .A(n7833), .ZN(P1_U3486) );
  AOI22_X1 U9559 ( .A1(n9734), .A2(n9210), .B1(n9908), .B2(
        P1_REG1_REG_11__SCAN_IN), .ZN(n7834) );
  OAI21_X1 U9560 ( .B1(n7835), .B2(n9908), .A(n7834), .ZN(P1_U3533) );
  XNOR2_X1 U9561 ( .A(n7836), .B(n9165), .ZN(n7837) );
  NOR2_X1 U9562 ( .A1(n7837), .A2(n7838), .ZN(n9164) );
  AOI21_X1 U9563 ( .B1(n7838), .B2(n7837), .A(n9164), .ZN(n7846) );
  AOI22_X1 U9564 ( .A1(n7839), .A2(n9209), .B1(n9244), .B2(n9257), .ZN(n7845)
         );
  INV_X1 U9565 ( .A(n7840), .ZN(n7843) );
  NAND2_X1 U9566 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_U3086), .ZN(n9308) );
  OAI21_X1 U9567 ( .B1(n9241), .B2(n7841), .A(n9308), .ZN(n7842) );
  AOI21_X1 U9568 ( .B1(n7843), .B2(n9229), .A(n7842), .ZN(n7844) );
  OAI211_X1 U9569 ( .C1(n7846), .C2(n9205), .A(n7845), .B(n7844), .ZN(P1_U3221) );
  INV_X1 U9570 ( .A(n7847), .ZN(n7850) );
  OAI222_X1 U9571 ( .A1(n8437), .A2(n10344), .B1(n8435), .B2(n7850), .C1(n7848), .C2(P2_U3151), .ZN(P2_U3273) );
  OAI222_X1 U9572 ( .A1(n9824), .A2(n7851), .B1(n9822), .B2(n7850), .C1(
        P1_U3086), .C2(n7849), .ZN(P1_U3333) );
  OAI21_X1 U9573 ( .B1(n7854), .B2(n7853), .A(n7852), .ZN(n7984) );
  INV_X1 U9574 ( .A(n7984), .ZN(n7867) );
  OAI211_X1 U9575 ( .C1(n7856), .C2(n7855), .A(n7957), .B(n9893), .ZN(n7857)
         );
  OAI21_X1 U9576 ( .B1(n8114), .B2(n9591), .A(n7857), .ZN(n7983) );
  INV_X1 U9577 ( .A(n7858), .ZN(n7860) );
  INV_X1 U9578 ( .A(n7859), .ZN(n7963) );
  OAI211_X1 U9579 ( .C1(n7989), .C2(n7860), .A(n7963), .B(n9628), .ZN(n7980)
         );
  INV_X1 U9580 ( .A(n7861), .ZN(n7890) );
  AOI22_X1 U9581 ( .A1(n9889), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n7890), .B2(
        n9632), .ZN(n7862) );
  OAI21_X1 U9582 ( .B1(n7981), .B2(n9606), .A(n7862), .ZN(n7863) );
  AOI21_X1 U9583 ( .B1(n9620), .B2(n7889), .A(n7863), .ZN(n7864) );
  OAI21_X1 U9584 ( .B1(n7980), .B2(n9489), .A(n7864), .ZN(n7865) );
  AOI21_X1 U9585 ( .B1(n9560), .B2(n7983), .A(n7865), .ZN(n7866) );
  OAI21_X1 U9586 ( .B1(n7867), .B2(n9637), .A(n7866), .ZN(P1_U3281) );
  NAND2_X1 U9587 ( .A1(n7868), .A2(n8307), .ZN(n7869) );
  XNOR2_X1 U9588 ( .A(n7869), .B(n8228), .ZN(n10007) );
  OR2_X1 U9589 ( .A1(n7801), .A2(n7870), .ZN(n7872) );
  AND2_X1 U9590 ( .A1(n7872), .A2(n7871), .ZN(n7873) );
  XNOR2_X1 U9591 ( .A(n7873), .B(n8228), .ZN(n7874) );
  OAI222_X1 U9592 ( .A1(n9951), .A2(n8006), .B1(n9953), .B2(n8087), .C1(n7874), 
        .C2(n9949), .ZN(n10009) );
  NAND2_X1 U9593 ( .A1(n10009), .A2(n8913), .ZN(n7877) );
  OAI22_X1 U9594 ( .A1(n8913), .A2(n5867), .B1(n8067), .B2(n9943), .ZN(n7875)
         );
  AOI21_X1 U9595 ( .B1(n8918), .B2(n8071), .A(n7875), .ZN(n7876) );
  OAI211_X1 U9596 ( .C1(n8922), .C2(n10007), .A(n7877), .B(n7876), .ZN(
        P2_U3222) );
  XNOR2_X1 U9597 ( .A(n7878), .B(n7879), .ZN(n10011) );
  INV_X1 U9598 ( .A(n7879), .ZN(n8327) );
  XNOR2_X1 U9599 ( .A(n7880), .B(n8327), .ZN(n7881) );
  OAI222_X1 U9600 ( .A1(n9951), .A2(n8063), .B1(n9953), .B2(n8140), .C1(n7881), 
        .C2(n9949), .ZN(n10012) );
  NAND2_X1 U9601 ( .A1(n10012), .A2(n8913), .ZN(n7884) );
  OAI22_X1 U9602 ( .A1(n8913), .A2(n6335), .B1(n8017), .B2(n9943), .ZN(n7882)
         );
  AOI21_X1 U9603 ( .B1(n8918), .B2(n10014), .A(n7882), .ZN(n7883) );
  OAI211_X1 U9604 ( .C1(n8922), .C2(n10011), .A(n7884), .B(n7883), .ZN(
        P2_U3221) );
  OAI21_X1 U9605 ( .B1(n7887), .B2(n7886), .A(n7885), .ZN(n7896) );
  AOI21_X1 U9606 ( .B1(n9244), .B2(n9253), .A(n7888), .ZN(n7894) );
  NAND2_X1 U9607 ( .A1(n9209), .A2(n7889), .ZN(n7893) );
  NAND2_X1 U9608 ( .A1(n9229), .A2(n7890), .ZN(n7892) );
  NAND2_X1 U9609 ( .A1(n9225), .A2(n9255), .ZN(n7891) );
  NAND4_X1 U9610 ( .A1(n7894), .A2(n7893), .A3(n7892), .A4(n7891), .ZN(n7895)
         );
  AOI21_X1 U9611 ( .B1(n7896), .B2(n9236), .A(n7895), .ZN(n7897) );
  INV_X1 U9612 ( .A(n7897), .ZN(P1_U3224) );
  XOR2_X1 U9613 ( .A(n7898), .B(n8224), .Z(n10001) );
  AOI22_X1 U9614 ( .A1(n8909), .A2(n8011), .B1(n8587), .B2(n8907), .ZN(n7904)
         );
  NAND2_X1 U9615 ( .A1(n7900), .A2(n7899), .ZN(n7901) );
  XOR2_X1 U9616 ( .A(n8224), .B(n7901), .Z(n7902) );
  NAND2_X1 U9617 ( .A1(n7902), .A2(n8912), .ZN(n7903) );
  OAI211_X1 U9618 ( .C1(n10001), .C2(n9939), .A(n7904), .B(n7903), .ZN(n10003)
         );
  NAND2_X1 U9619 ( .A1(n10003), .A2(n8913), .ZN(n7908) );
  OAI22_X1 U9620 ( .A1(n8913), .A2(n7905), .B1(n7995), .B2(n9943), .ZN(n7906)
         );
  AOI21_X1 U9621 ( .B1(n8918), .B2(n7996), .A(n7906), .ZN(n7907) );
  OAI211_X1 U9622 ( .C1(n10001), .C2(n9956), .A(n7908), .B(n7907), .ZN(
        P2_U3223) );
  XNOR2_X1 U9623 ( .A(n7909), .B(n7910), .ZN(n7911) );
  NAND2_X1 U9624 ( .A1(n7911), .A2(n7912), .ZN(n9199) );
  OAI21_X1 U9625 ( .B1(n7912), .B2(n7911), .A(n9199), .ZN(n7913) );
  NAND2_X1 U9626 ( .A1(n7913), .A2(n9236), .ZN(n7923) );
  INV_X1 U9627 ( .A(n7914), .ZN(n7921) );
  NOR2_X1 U9628 ( .A1(n9247), .A2(n7915), .ZN(n7920) );
  NAND2_X1 U9629 ( .A1(n9225), .A2(n9257), .ZN(n7918) );
  INV_X1 U9630 ( .A(n7916), .ZN(n7917) );
  OAI211_X1 U9631 ( .C1(n7981), .C2(n9227), .A(n7918), .B(n7917), .ZN(n7919)
         );
  AOI211_X1 U9632 ( .C1(n9229), .C2(n7921), .A(n7920), .B(n7919), .ZN(n7922)
         );
  NAND2_X1 U9633 ( .A1(n7923), .A2(n7922), .ZN(P1_U3217) );
  AOI21_X1 U9634 ( .B1(n7925), .B2(n5870), .A(n7924), .ZN(n7939) );
  OAI21_X1 U9635 ( .B1(n7928), .B2(n7927), .A(n7926), .ZN(n7937) );
  AND2_X1 U9636 ( .A1(P2_U3151), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n8068) );
  AOI21_X1 U9637 ( .B1(n5867), .B2(n7930), .A(n7929), .ZN(n7931) );
  NOR2_X1 U9638 ( .A1(n9929), .A2(n7931), .ZN(n7932) );
  AOI211_X1 U9639 ( .C1(n7933), .C2(n8709), .A(n8068), .B(n7932), .ZN(n7934)
         );
  OAI21_X1 U9640 ( .B1(n7935), .B2(n8735), .A(n7934), .ZN(n7936) );
  AOI21_X1 U9641 ( .B1(n9918), .B2(n7937), .A(n7936), .ZN(n7938) );
  OAI21_X1 U9642 ( .B1(n7939), .B2(n9930), .A(n7938), .ZN(P2_U3193) );
  INV_X1 U9643 ( .A(n7943), .ZN(n7942) );
  NAND2_X1 U9644 ( .A1(n9817), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n7940) );
  OAI211_X1 U9645 ( .C1(n7942), .C2(n9822), .A(n7941), .B(n7940), .ZN(P1_U3332) );
  NAND2_X1 U9646 ( .A1(n7943), .A2(n9043), .ZN(n7945) );
  NAND2_X1 U9647 ( .A1(n7944), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8427) );
  OAI211_X1 U9648 ( .C1(n7946), .C2(n8437), .A(n7945), .B(n8427), .ZN(P2_U3272) );
  AOI21_X1 U9649 ( .B1(n7948), .B2(n9970), .A(n7947), .ZN(n7952) );
  AOI22_X1 U9650 ( .A1(n8966), .A2(n7950), .B1(n10027), .B2(
        P2_REG1_REG_9__SCAN_IN), .ZN(n7949) );
  OAI21_X1 U9651 ( .B1(n7952), .B2(n10027), .A(n7949), .ZN(P2_U3468) );
  AOI22_X1 U9652 ( .A1(n6396), .A2(n7950), .B1(n10017), .B2(
        P2_REG0_REG_9__SCAN_IN), .ZN(n7951) );
  OAI21_X1 U9653 ( .B1(n7952), .B2(n10017), .A(n7951), .ZN(P2_U3417) );
  OAI21_X1 U9654 ( .B1(n7954), .B2(n7960), .A(n7953), .ZN(n7955) );
  INV_X1 U9655 ( .A(n7955), .ZN(n9748) );
  NAND2_X1 U9656 ( .A1(n7957), .A2(n7956), .ZN(n7959) );
  INV_X1 U9657 ( .A(n8101), .ZN(n7958) );
  AOI21_X1 U9658 ( .B1(n7960), .B2(n7959), .A(n7958), .ZN(n7961) );
  OAI222_X1 U9659 ( .A1(n9591), .A2(n9240), .B1(n9705), .B2(n7962), .C1(n9498), 
        .C2(n7961), .ZN(n9742) );
  AOI211_X1 U9660 ( .C1(n9744), .C2(n7963), .A(n9567), .B(n8106), .ZN(n9743)
         );
  NAND2_X1 U9661 ( .A1(n9743), .A2(n9578), .ZN(n7966) );
  INV_X1 U9662 ( .A(n7964), .ZN(n7976) );
  AOI22_X1 U9663 ( .A1(n9889), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n7976), .B2(
        n9632), .ZN(n7965) );
  OAI211_X1 U9664 ( .C1(n7979), .C2(n9585), .A(n7966), .B(n7965), .ZN(n7967)
         );
  AOI21_X1 U9665 ( .B1(n9560), .B2(n9742), .A(n7967), .ZN(n7968) );
  OAI21_X1 U9666 ( .B1(n9748), .B2(n9637), .A(n7968), .ZN(P1_U3280) );
  OAI21_X1 U9667 ( .B1(n7971), .B2(n7970), .A(n7969), .ZN(n7972) );
  NAND2_X1 U9668 ( .A1(n7972), .A2(n9236), .ZN(n7978) );
  AOI21_X1 U9669 ( .B1(n9225), .B2(n9254), .A(n7973), .ZN(n7974) );
  OAI21_X1 U9670 ( .B1(n9240), .B2(n9227), .A(n7974), .ZN(n7975) );
  AOI21_X1 U9671 ( .B1(n7976), .B2(n9229), .A(n7975), .ZN(n7977) );
  OAI211_X1 U9672 ( .C1(n7979), .C2(n9247), .A(n7978), .B(n7977), .ZN(P1_U3234) );
  OAI21_X1 U9673 ( .B1(n7981), .B2(n9705), .A(n7980), .ZN(n7982) );
  AOI211_X1 U9674 ( .C1(n7984), .C2(n9903), .A(n7983), .B(n7982), .ZN(n7986)
         );
  MUX2_X1 U9675 ( .A(n5307), .B(n7986), .S(n9906), .Z(n7985) );
  OAI21_X1 U9676 ( .B1(n7989), .B2(n9755), .A(n7985), .ZN(P1_U3489) );
  MUX2_X1 U9677 ( .A(n7987), .B(n7986), .S(n9910), .Z(n7988) );
  OAI21_X1 U9678 ( .B1(n7989), .B2(n9644), .A(n7988), .ZN(P1_U3534) );
  INV_X1 U9679 ( .A(n7990), .ZN(n7992) );
  NAND2_X1 U9680 ( .A1(n7994), .A2(n7993), .ZN(n8008) );
  XNOR2_X1 U9681 ( .A(n8008), .B(n8586), .ZN(n8062) );
  XNOR2_X1 U9682 ( .A(n7996), .B(n8186), .ZN(n8009) );
  XNOR2_X1 U9683 ( .A(n8062), .B(n8009), .ZN(n8004) );
  INV_X1 U9684 ( .A(n7995), .ZN(n8002) );
  INV_X1 U9685 ( .A(n7996), .ZN(n9999) );
  NOR2_X1 U9686 ( .A1(n8554), .A2(n9999), .ZN(n8001) );
  NAND2_X1 U9687 ( .A1(n8568), .A2(n8587), .ZN(n7999) );
  INV_X1 U9688 ( .A(n7997), .ZN(n7998) );
  OAI211_X1 U9689 ( .C1(n8566), .C2(n8063), .A(n7999), .B(n7998), .ZN(n8000)
         );
  AOI211_X1 U9690 ( .C1(n8002), .C2(n8558), .A(n8001), .B(n8000), .ZN(n8003)
         );
  OAI21_X1 U9691 ( .B1(n8004), .B2(n8571), .A(n8003), .ZN(P2_U3157) );
  INV_X1 U9692 ( .A(n8005), .ZN(n8077) );
  OAI222_X1 U9693 ( .A1(n5607), .A2(P1_U3086), .B1(n9822), .B2(n8077), .C1(
        n10271), .C2(n9824), .ZN(P1_U3331) );
  INV_X1 U9694 ( .A(n10014), .ZN(n8024) );
  XNOR2_X1 U9695 ( .A(n8071), .B(n8186), .ZN(n8064) );
  AOI22_X1 U9696 ( .A1(n8064), .A2(n8063), .B1(n8006), .B2(n8009), .ZN(n8007)
         );
  NAND2_X1 U9697 ( .A1(n8008), .A2(n8007), .ZN(n8014) );
  INV_X1 U9698 ( .A(n8009), .ZN(n8061) );
  AOI21_X1 U9699 ( .B1(n8061), .B2(n8586), .A(n8011), .ZN(n8010) );
  NAND3_X1 U9700 ( .A1(n8061), .A2(n8011), .A3(n8586), .ZN(n8012) );
  NAND2_X1 U9701 ( .A1(n8014), .A2(n4976), .ZN(n8016) );
  XNOR2_X1 U9702 ( .A(n10014), .B(n8186), .ZN(n8088) );
  XNOR2_X1 U9703 ( .A(n8088), .B(n8585), .ZN(n8015) );
  NAND2_X1 U9704 ( .A1(n8016), .A2(n8015), .ZN(n8090) );
  OAI211_X1 U9705 ( .C1(n8016), .C2(n8015), .A(n8090), .B(n8545), .ZN(n8023)
         );
  INV_X1 U9706 ( .A(n8017), .ZN(n8021) );
  NOR2_X1 U9707 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8018), .ZN(n8626) );
  AOI21_X1 U9708 ( .B1(n8548), .B2(n8584), .A(n8626), .ZN(n8019) );
  OAI21_X1 U9709 ( .B1(n8063), .B2(n8550), .A(n8019), .ZN(n8020) );
  AOI21_X1 U9710 ( .B1(n8021), .B2(n8558), .A(n8020), .ZN(n8022) );
  OAI211_X1 U9711 ( .C1(n8024), .C2(n8554), .A(n8023), .B(n8022), .ZN(P2_U3164) );
  NAND2_X1 U9712 ( .A1(n8334), .A2(n8335), .ZN(n8332) );
  XNOR2_X1 U9713 ( .A(n8025), .B(n8332), .ZN(n8084) );
  INV_X1 U9714 ( .A(n8332), .ZN(n8027) );
  XNOR2_X1 U9715 ( .A(n8026), .B(n8027), .ZN(n8028) );
  NAND2_X1 U9716 ( .A1(n8028), .A2(n8912), .ZN(n8030) );
  AOI22_X1 U9717 ( .A1(n8907), .A2(n8584), .B1(n8894), .B2(n8909), .ZN(n8029)
         );
  NAND2_X1 U9718 ( .A1(n8030), .A2(n8029), .ZN(n8083) );
  INV_X1 U9719 ( .A(n8145), .ZN(n8459) );
  OAI22_X1 U9720 ( .A1(n8459), .A2(n9944), .B1(n8451), .B2(n9943), .ZN(n8031)
         );
  OAI21_X1 U9721 ( .B1(n8083), .B2(n8031), .A(n8913), .ZN(n8033) );
  NAND2_X1 U9722 ( .A1(n9960), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n8032) );
  OAI211_X1 U9723 ( .C1(n8922), .C2(n8084), .A(n8033), .B(n8032), .ZN(P2_U3219) );
  XNOR2_X1 U9724 ( .A(n8096), .B(n8584), .ZN(n8326) );
  XNOR2_X1 U9725 ( .A(n8034), .B(n8326), .ZN(n8048) );
  INV_X1 U9726 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n8037) );
  XOR2_X1 U9727 ( .A(n8035), .B(n8326), .Z(n8036) );
  AOI222_X1 U9728 ( .A1(n8912), .A2(n8036), .B1(n8908), .B2(n8909), .C1(n8585), 
        .C2(n8907), .ZN(n8042) );
  MUX2_X1 U9729 ( .A(n8037), .B(n8042), .S(n10016), .Z(n8039) );
  NAND2_X1 U9730 ( .A1(n8096), .A2(n6396), .ZN(n8038) );
  OAI211_X1 U9731 ( .C1(n9022), .C2(n8048), .A(n8039), .B(n8038), .ZN(P2_U3429) );
  INV_X1 U9732 ( .A(n8967), .ZN(n8958) );
  MUX2_X1 U9733 ( .A(n5898), .B(n8042), .S(n10029), .Z(n8041) );
  NAND2_X1 U9734 ( .A1(n8096), .A2(n8966), .ZN(n8040) );
  OAI211_X1 U9735 ( .C1(n8048), .C2(n8958), .A(n8041), .B(n8040), .ZN(P2_U3472) );
  INV_X1 U9736 ( .A(n8042), .ZN(n8045) );
  INV_X1 U9737 ( .A(n8096), .ZN(n8043) );
  OAI22_X1 U9738 ( .A1(n8043), .A2(n9944), .B1(n8094), .B2(n9943), .ZN(n8044)
         );
  OAI21_X1 U9739 ( .B1(n8045), .B2(n8044), .A(n8913), .ZN(n8047) );
  NAND2_X1 U9740 ( .A1(n9960), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n8046) );
  OAI211_X1 U9741 ( .C1(n8922), .C2(n8048), .A(n8047), .B(n8046), .ZN(P2_U3220) );
  XNOR2_X1 U9742 ( .A(n8049), .B(n8053), .ZN(n9741) );
  INV_X1 U9743 ( .A(n8050), .ZN(n8051) );
  AOI21_X1 U9744 ( .B1(n8053), .B2(n8052), .A(n8051), .ZN(n8054) );
  OAI222_X1 U9745 ( .A1(n9591), .A2(n9607), .B1(n9705), .B2(n9240), .C1(n9498), 
        .C2(n8054), .ZN(n9737) );
  INV_X1 U9746 ( .A(n9627), .ZN(n8055) );
  AOI211_X1 U9747 ( .C1(n9739), .C2(n8105), .A(n9567), .B(n8055), .ZN(n9738)
         );
  NAND2_X1 U9748 ( .A1(n9738), .A2(n9578), .ZN(n8058) );
  INV_X1 U9749 ( .A(n9238), .ZN(n8056) );
  AOI22_X1 U9750 ( .A1(n9889), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n8056), .B2(
        n9632), .ZN(n8057) );
  OAI211_X1 U9751 ( .C1(n9248), .C2(n9585), .A(n8058), .B(n8057), .ZN(n8059)
         );
  AOI21_X1 U9752 ( .B1(n9560), .B2(n9737), .A(n8059), .ZN(n8060) );
  OAI21_X1 U9753 ( .B1(n9741), .B2(n9637), .A(n8060), .ZN(P1_U3278) );
  OAI22_X1 U9754 ( .A1(n8062), .A2(n8061), .B1(n8008), .B2(n8586), .ZN(n8066)
         );
  XNOR2_X1 U9755 ( .A(n8064), .B(n8063), .ZN(n8065) );
  XNOR2_X1 U9756 ( .A(n8066), .B(n8065), .ZN(n8076) );
  INV_X1 U9757 ( .A(n8067), .ZN(n8074) );
  NAND2_X1 U9758 ( .A1(n8568), .A2(n8586), .ZN(n8070) );
  INV_X1 U9759 ( .A(n8068), .ZN(n8069) );
  OAI211_X1 U9760 ( .C1(n8566), .C2(n8087), .A(n8070), .B(n8069), .ZN(n8073)
         );
  INV_X1 U9761 ( .A(n8071), .ZN(n10006) );
  NOR2_X1 U9762 ( .A1(n10006), .A2(n8554), .ZN(n8072) );
  AOI211_X1 U9763 ( .C1(n8074), .C2(n8558), .A(n8073), .B(n8072), .ZN(n8075)
         );
  OAI21_X1 U9764 ( .B1(n8076), .B2(n8571), .A(n8075), .ZN(P2_U3176) );
  OAI222_X1 U9765 ( .A1(n8435), .A2(n8077), .B1(P2_U3151), .B2(n6129), .C1(
        n10235), .C2(n8437), .ZN(P2_U3271) );
  MUX2_X1 U9766 ( .A(n8083), .B(P2_REG0_REG_14__SCAN_IN), .S(n10017), .Z(n8079) );
  OAI22_X1 U9767 ( .A1(n8084), .A2(n9022), .B1(n8459), .B2(n9013), .ZN(n8078)
         );
  OR2_X1 U9768 ( .A1(n8079), .A2(n8078), .ZN(P2_U3432) );
  INV_X1 U9769 ( .A(n8080), .ZN(n8134) );
  OAI222_X1 U9770 ( .A1(n8082), .A2(P1_U3086), .B1(n9822), .B2(n8134), .C1(
        n8081), .C2(n9824), .ZN(P1_U3330) );
  MUX2_X1 U9771 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n8083), .S(n10029), .Z(n8086) );
  OAI22_X1 U9772 ( .A1(n8084), .A2(n8958), .B1(n8459), .B2(n8950), .ZN(n8085)
         );
  OR2_X1 U9773 ( .A1(n8086), .A2(n8085), .ZN(P2_U3473) );
  OR2_X1 U9774 ( .A1(n8088), .A2(n8087), .ZN(n8089) );
  NAND2_X1 U9775 ( .A1(n8090), .A2(n8089), .ZN(n8144) );
  XNOR2_X1 U9776 ( .A(n8096), .B(n8186), .ZN(n8141) );
  XNOR2_X1 U9777 ( .A(n8141), .B(n8584), .ZN(n8091) );
  XNOR2_X1 U9778 ( .A(n8144), .B(n8091), .ZN(n8098) );
  AND2_X1 U9779 ( .A1(P2_U3151), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n8642) );
  NOR2_X1 U9780 ( .A1(n8566), .A2(n8147), .ZN(n8092) );
  AOI211_X1 U9781 ( .C1(n8568), .C2(n8585), .A(n8642), .B(n8092), .ZN(n8093)
         );
  OAI21_X1 U9782 ( .B1(n8094), .B2(n8570), .A(n8093), .ZN(n8095) );
  AOI21_X1 U9783 ( .B1(n8096), .B2(n8576), .A(n8095), .ZN(n8097) );
  OAI21_X1 U9784 ( .B1(n8098), .B2(n8571), .A(n8097), .ZN(P2_U3174) );
  XOR2_X1 U9785 ( .A(n8099), .B(n8102), .Z(n8124) );
  NAND2_X1 U9786 ( .A1(n8101), .A2(n8100), .ZN(n8103) );
  XNOR2_X1 U9787 ( .A(n8103), .B(n8102), .ZN(n8104) );
  OAI22_X1 U9788 ( .A1(n8104), .A2(n9498), .B1(n9134), .B2(n9591), .ZN(n8118)
         );
  OAI211_X1 U9789 ( .C1(n8106), .C2(n8115), .A(n9628), .B(n8105), .ZN(n8113)
         );
  NOR2_X1 U9790 ( .A1(n9606), .A2(n8114), .ZN(n8109) );
  OAI22_X1 U9791 ( .A1(n9560), .A2(n8107), .B1(n9057), .B2(n9886), .ZN(n8108)
         );
  AOI211_X1 U9792 ( .C1(n9059), .C2(n9620), .A(n8109), .B(n8108), .ZN(n8110)
         );
  OAI21_X1 U9793 ( .B1(n8113), .B2(n9489), .A(n8110), .ZN(n8111) );
  AOI21_X1 U9794 ( .B1(n8118), .B2(n9560), .A(n8111), .ZN(n8112) );
  OAI21_X1 U9795 ( .B1(n8124), .B2(n9637), .A(n8112), .ZN(P1_U3279) );
  INV_X1 U9796 ( .A(n8113), .ZN(n8117) );
  OAI22_X1 U9797 ( .A1(n8115), .A2(n9899), .B1(n8114), .B2(n9705), .ZN(n8116)
         );
  NOR3_X1 U9798 ( .A1(n8118), .A2(n8117), .A3(n8116), .ZN(n8121) );
  NOR2_X1 U9799 ( .A1(n8121), .A2(n9905), .ZN(n8119) );
  AOI21_X1 U9800 ( .B1(P1_REG0_REG_14__SCAN_IN), .B2(n9905), .A(n8119), .ZN(
        n8120) );
  OAI21_X1 U9801 ( .B1(n8124), .B2(n9803), .A(n8120), .ZN(P1_U3495) );
  NOR2_X1 U9802 ( .A1(n8121), .A2(n9908), .ZN(n8122) );
  AOI21_X1 U9803 ( .B1(P1_REG1_REG_14__SCAN_IN), .B2(n9908), .A(n8122), .ZN(
        n8123) );
  OAI21_X1 U9804 ( .B1(n8124), .B2(n9736), .A(n8123), .ZN(P1_U3536) );
  INV_X1 U9805 ( .A(n8125), .ZN(n8127) );
  OAI222_X1 U9806 ( .A1(n8435), .A2(n8127), .B1(P2_U3151), .B2(n8136), .C1(
        n10143), .C2(n8437), .ZN(P2_U3269) );
  OAI222_X1 U9807 ( .A1(n8128), .A2(P1_U3086), .B1(n9822), .B2(n8127), .C1(
        n8126), .C2(n9824), .ZN(P1_U3329) );
  NAND2_X1 U9808 ( .A1(n6080), .A2(n9043), .ZN(n8130) );
  OAI211_X1 U9809 ( .C1(n8437), .C2(n10301), .A(n8130), .B(n8129), .ZN(
        P2_U3267) );
  INV_X1 U9810 ( .A(n6080), .ZN(n8131) );
  OAI222_X1 U9811 ( .A1(n9824), .A2(n8132), .B1(n9822), .B2(n8131), .C1(n5643), 
        .C2(P1_U3086), .ZN(P1_U3327) );
  OAI222_X1 U9812 ( .A1(n8435), .A2(n8134), .B1(P2_U3151), .B2(n6133), .C1(
        n8133), .C2(n8437), .ZN(P2_U3270) );
  INV_X1 U9813 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n8138) );
  AND2_X1 U9814 ( .A1(n8136), .A2(n8135), .ZN(n8137) );
  AOI22_X1 U9815 ( .A1(n8139), .A2(n8138), .B1(n8137), .B2(n6133), .ZN(
        P2_U3377) );
  NAND2_X1 U9816 ( .A1(n8141), .A2(n8140), .ZN(n8143) );
  INV_X1 U9817 ( .A(n8141), .ZN(n8142) );
  AOI21_X1 U9818 ( .B1(n8144), .B2(n8143), .A(n4985), .ZN(n8449) );
  XNOR2_X1 U9819 ( .A(n8145), .B(n8186), .ZN(n8146) );
  XNOR2_X1 U9820 ( .A(n8146), .B(n8908), .ZN(n8448) );
  NAND2_X1 U9821 ( .A1(n8449), .A2(n8448), .ZN(n8447) );
  NAND2_X1 U9822 ( .A1(n8146), .A2(n8147), .ZN(n8148) );
  NAND2_X1 U9823 ( .A1(n8447), .A2(n8148), .ZN(n8572) );
  XNOR2_X1 U9824 ( .A(n9037), .B(n8186), .ZN(n8150) );
  XNOR2_X1 U9825 ( .A(n8150), .B(n8454), .ZN(n8573) );
  XNOR2_X1 U9826 ( .A(n9031), .B(n8182), .ZN(n8149) );
  NOR2_X1 U9827 ( .A1(n8149), .A2(n8910), .ZN(n8505) );
  AOI21_X1 U9828 ( .B1(n8149), .B2(n8910), .A(n8505), .ZN(n8495) );
  INV_X1 U9829 ( .A(n8150), .ZN(n8151) );
  NAND2_X1 U9830 ( .A1(n8151), .A2(n8894), .ZN(n8496) );
  XNOR2_X1 U9831 ( .A(n9025), .B(n8186), .ZN(n8152) );
  NAND2_X1 U9832 ( .A1(n8152), .A2(n8896), .ZN(n8543) );
  INV_X1 U9833 ( .A(n8152), .ZN(n8153) );
  NAND2_X1 U9834 ( .A1(n8153), .A2(n8583), .ZN(n8154) );
  AND2_X1 U9835 ( .A1(n8543), .A2(n8154), .ZN(n8504) );
  XNOR2_X1 U9836 ( .A(n8956), .B(n8186), .ZN(n8155) );
  NAND2_X1 U9837 ( .A1(n8155), .A2(n8509), .ZN(n8467) );
  INV_X1 U9838 ( .A(n8155), .ZN(n8156) );
  NAND2_X1 U9839 ( .A1(n8156), .A2(n8881), .ZN(n8157) );
  AND2_X1 U9840 ( .A1(n8467), .A2(n8157), .ZN(n8544) );
  NAND2_X1 U9841 ( .A1(n8158), .A2(n8544), .ZN(n8466) );
  NAND2_X1 U9842 ( .A1(n8466), .A2(n8467), .ZN(n8162) );
  XNOR2_X1 U9843 ( .A(n8952), .B(n8186), .ZN(n8159) );
  NAND2_X1 U9844 ( .A1(n8159), .A2(n8868), .ZN(n8522) );
  INV_X1 U9845 ( .A(n8159), .ZN(n8160) );
  NAND2_X1 U9846 ( .A1(n8160), .A2(n8582), .ZN(n8161) );
  AND2_X1 U9847 ( .A1(n8522), .A2(n8161), .ZN(n8468) );
  NAND2_X1 U9848 ( .A1(n8162), .A2(n8468), .ZN(n8470) );
  NAND2_X1 U9849 ( .A1(n8470), .A2(n8522), .ZN(n8166) );
  XNOR2_X1 U9850 ( .A(n8521), .B(n8186), .ZN(n8163) );
  NAND2_X1 U9851 ( .A1(n8163), .A2(n8856), .ZN(n8480) );
  INV_X1 U9852 ( .A(n8163), .ZN(n8164) );
  NAND2_X1 U9853 ( .A1(n8164), .A2(n8581), .ZN(n8165) );
  AND2_X1 U9854 ( .A1(n8480), .A2(n8165), .ZN(n8523) );
  XNOR2_X1 U9855 ( .A(n8478), .B(n8186), .ZN(n8167) );
  XNOR2_X1 U9856 ( .A(n8167), .B(n8818), .ZN(n8481) );
  XNOR2_X1 U9857 ( .A(n9002), .B(n8182), .ZN(n8168) );
  NOR2_X1 U9858 ( .A1(n8168), .A2(n8807), .ZN(n8532) );
  NAND2_X1 U9859 ( .A1(n8168), .A2(n8807), .ZN(n8533) );
  NAND2_X1 U9860 ( .A1(n8460), .A2(n8539), .ZN(n8173) );
  INV_X1 U9861 ( .A(n8169), .ZN(n8171) );
  OR2_X1 U9862 ( .A1(n8171), .A2(n8170), .ZN(n8172) );
  NAND2_X1 U9863 ( .A1(n8173), .A2(n8172), .ZN(n8514) );
  XNOR2_X1 U9864 ( .A(n8991), .B(n8186), .ZN(n8174) );
  XNOR2_X1 U9865 ( .A(n8174), .B(n8806), .ZN(n8515) );
  NAND2_X1 U9866 ( .A1(n8174), .A2(n8777), .ZN(n8175) );
  XNOR2_X1 U9867 ( .A(n8985), .B(n8186), .ZN(n8177) );
  XNOR2_X1 U9868 ( .A(n8177), .B(n8793), .ZN(n8488) );
  XNOR2_X1 U9869 ( .A(n8979), .B(n8186), .ZN(n8179) );
  XNOR2_X1 U9870 ( .A(n8179), .B(n8775), .ZN(n8557) );
  NAND2_X1 U9871 ( .A1(n8556), .A2(n8557), .ZN(n8181) );
  NAND2_X1 U9872 ( .A1(n8179), .A2(n8178), .ZN(n8180) );
  NAND2_X1 U9873 ( .A1(n8181), .A2(n8180), .ZN(n8438) );
  XNOR2_X1 U9874 ( .A(n8183), .B(n8182), .ZN(n8184) );
  NAND2_X1 U9875 ( .A1(n8184), .A2(n8768), .ZN(n8185) );
  OAI21_X1 U9876 ( .B1(n8184), .B2(n8768), .A(n8185), .ZN(n8439) );
  AOI22_X1 U9877 ( .A1(n8768), .A2(n8568), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3151), .ZN(n8189) );
  NAND2_X1 U9878 ( .A1(n8187), .A2(n8558), .ZN(n8188) );
  OAI211_X1 U9879 ( .C1(n8190), .C2(n8566), .A(n8189), .B(n8188), .ZN(n8191)
         );
  AOI21_X1 U9880 ( .B1(n8192), .B2(n8576), .A(n8191), .ZN(n8193) );
  INV_X1 U9881 ( .A(n8194), .ZN(n8198) );
  OAI222_X1 U9882 ( .A1(n9824), .A2(n8196), .B1(P1_U3086), .B2(n8195), .C1(
        n8198), .C2(n9822), .ZN(P1_U3328) );
  OAI222_X1 U9883 ( .A1(n8435), .A2(n8198), .B1(n6107), .B2(P2_U3151), .C1(
        n8197), .C2(n8437), .ZN(P2_U3268) );
  NAND2_X1 U9884 ( .A1(n8429), .A2(n8202), .ZN(n8200) );
  INV_X1 U9885 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n8436) );
  OR2_X1 U9886 ( .A1(n5764), .A2(n8436), .ZN(n8199) );
  NAND2_X1 U9887 ( .A1(n8200), .A2(n8199), .ZN(n8973) );
  INV_X1 U9888 ( .A(n8973), .ZN(n8748) );
  AOI22_X1 U9889 ( .A1(n9812), .A2(n8202), .B1(n8201), .B2(
        P1_DATAO_REG_31__SCAN_IN), .ZN(n8972) );
  INV_X1 U9890 ( .A(n8972), .ZN(n8923) );
  INV_X1 U9891 ( .A(n8578), .ZN(n8403) );
  NAND2_X1 U9892 ( .A1(n8973), .A2(n8403), .ZN(n8213) );
  NAND2_X1 U9893 ( .A1(n8213), .A2(n8204), .ZN(n8405) );
  INV_X1 U9894 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n8209) );
  NAND2_X1 U9895 ( .A1(n6061), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n8207) );
  INV_X1 U9896 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n8205) );
  OR2_X1 U9897 ( .A1(n5774), .A2(n8205), .ZN(n8206) );
  OAI211_X1 U9898 ( .C1(n8209), .C2(n8208), .A(n8207), .B(n8206), .ZN(n8210)
         );
  INV_X1 U9899 ( .A(n8210), .ZN(n8211) );
  NAND2_X1 U9900 ( .A1(n8212), .A2(n8211), .ZN(n8742) );
  NAND2_X1 U9901 ( .A1(n8972), .A2(n8742), .ZN(n8415) );
  INV_X1 U9902 ( .A(n8213), .ZN(n8237) );
  AND2_X1 U9903 ( .A1(n8748), .A2(n8578), .ZN(n8395) );
  INV_X1 U9904 ( .A(n8214), .ZN(n8384) );
  INV_X1 U9905 ( .A(n8386), .ZN(n8234) );
  INV_X1 U9906 ( .A(n8774), .ZN(n8788) );
  NAND2_X1 U9907 ( .A1(n8786), .A2(n8376), .ZN(n8801) );
  INV_X1 U9908 ( .A(n8798), .ZN(n8374) );
  INV_X1 U9909 ( .A(n8817), .ZN(n8814) );
  INV_X1 U9910 ( .A(n8215), .ZN(n8830) );
  INV_X1 U9911 ( .A(n8857), .ZN(n8853) );
  INV_X1 U9912 ( .A(n8888), .ZN(n8892) );
  INV_X1 U9913 ( .A(n8216), .ZN(n8348) );
  NOR3_X1 U9914 ( .A1(n8217), .A2(n8268), .A3(n8250), .ZN(n8220) );
  INV_X1 U9915 ( .A(n7531), .ZN(n8218) );
  NAND4_X1 U9916 ( .A1(n8220), .A2(n8219), .A3(n8218), .A4(n8270), .ZN(n8223)
         );
  NOR4_X1 U9917 ( .A1(n8223), .A2(n8222), .A3(n4441), .A4(n8221), .ZN(n8226)
         );
  NAND4_X1 U9918 ( .A1(n8226), .A2(n8225), .A3(n8224), .A4(n8294), .ZN(n8227)
         );
  NOR4_X1 U9919 ( .A1(n8332), .A2(n8327), .A3(n8228), .A4(n8227), .ZN(n8229)
         );
  NAND4_X1 U9920 ( .A1(n8892), .A2(n8905), .A3(n8229), .A4(n8326), .ZN(n8230)
         );
  NOR4_X1 U9921 ( .A1(n8853), .A2(n8341), .A3(n8870), .A4(n8230), .ZN(n8231)
         );
  NAND4_X1 U9922 ( .A1(n8814), .A2(n8842), .A3(n8830), .A4(n8231), .ZN(n8232)
         );
  NOR4_X1 U9923 ( .A1(n8788), .A2(n8801), .A3(n8804), .A4(n8232), .ZN(n8233)
         );
  NAND4_X1 U9924 ( .A1(n8235), .A2(n8764), .A3(n8234), .A4(n8233), .ZN(n8236)
         );
  NOR4_X1 U9925 ( .A1(n8237), .A2(n8395), .A3(n8394), .A4(n8236), .ZN(n8238)
         );
  AOI22_X1 U9926 ( .A1(n8239), .A2(n8250), .B1(n8238), .B2(n8415), .ZN(n8419)
         );
  NOR2_X1 U9927 ( .A1(n8972), .A2(n8742), .ZN(n8410) );
  NOR2_X1 U9928 ( .A1(n8410), .A2(n6195), .ZN(n8241) );
  NAND2_X1 U9929 ( .A1(n8923), .A2(n8395), .ZN(n8240) );
  NAND2_X1 U9930 ( .A1(n8241), .A2(n8240), .ZN(n8418) );
  INV_X1 U9931 ( .A(n8242), .ZN(n8243) );
  NOR2_X1 U9932 ( .A1(n8784), .A2(n8243), .ZN(n8244) );
  MUX2_X1 U9933 ( .A(n8245), .B(n8244), .S(n8406), .Z(n8371) );
  INV_X1 U9934 ( .A(n8343), .ZN(n8347) );
  NAND2_X1 U9935 ( .A1(n8246), .A2(n8402), .ZN(n8283) );
  NAND2_X1 U9936 ( .A1(n8287), .A2(n8263), .ZN(n8247) );
  NOR2_X1 U9937 ( .A1(n8283), .A2(n8247), .ZN(n8274) );
  NAND3_X1 U9938 ( .A1(n8285), .A2(n8248), .A3(n8406), .ZN(n8279) );
  NOR2_X1 U9939 ( .A1(n8279), .A2(n8249), .ZN(n8273) );
  AND2_X1 U9940 ( .A1(n8253), .A2(n8250), .ZN(n8252) );
  OAI21_X1 U9941 ( .B1(n8252), .B2(n8251), .A(n8256), .ZN(n8259) );
  INV_X1 U9942 ( .A(n8253), .ZN(n8255) );
  NAND2_X1 U9943 ( .A1(n8255), .A2(n8254), .ZN(n8257) );
  AND2_X1 U9944 ( .A1(n8257), .A2(n8256), .ZN(n8258) );
  MUX2_X1 U9945 ( .A(n8259), .B(n8258), .S(n8406), .Z(n8269) );
  NAND2_X1 U9946 ( .A1(n8261), .A2(n8260), .ZN(n8265) );
  NAND2_X1 U9947 ( .A1(n8263), .A2(n8262), .ZN(n8264) );
  MUX2_X1 U9948 ( .A(n8265), .B(n8264), .S(n8406), .Z(n8266) );
  INV_X1 U9949 ( .A(n8266), .ZN(n8267) );
  OAI21_X1 U9950 ( .B1(n8269), .B2(n8268), .A(n8267), .ZN(n8271) );
  AND2_X1 U9951 ( .A1(n8271), .A2(n8270), .ZN(n8272) );
  OAI21_X1 U9952 ( .B1(n8274), .B2(n8273), .A(n8272), .ZN(n8296) );
  NAND2_X1 U9953 ( .A1(n8306), .A2(n8303), .ZN(n8301) );
  NAND2_X1 U9954 ( .A1(n8301), .A2(n8402), .ZN(n8276) );
  AND2_X1 U9955 ( .A1(n8299), .A2(n8298), .ZN(n8275) );
  AND2_X1 U9956 ( .A1(n8276), .A2(n8275), .ZN(n8302) );
  AOI21_X1 U9957 ( .B1(n8277), .B2(n8402), .A(n9990), .ZN(n8292) );
  AOI21_X1 U9958 ( .B1(n8590), .B2(n8406), .A(n8278), .ZN(n8291) );
  INV_X1 U9959 ( .A(n8287), .ZN(n8282) );
  AND2_X1 U9960 ( .A1(n8592), .A2(n9978), .ZN(n8281) );
  INV_X1 U9961 ( .A(n8279), .ZN(n8280) );
  OAI21_X1 U9962 ( .B1(n8282), .B2(n8281), .A(n8280), .ZN(n8290) );
  INV_X1 U9963 ( .A(n8283), .ZN(n8288) );
  NAND2_X1 U9964 ( .A1(n8285), .A2(n8284), .ZN(n8286) );
  NAND3_X1 U9965 ( .A1(n8288), .A2(n8287), .A3(n8286), .ZN(n8289) );
  OAI211_X1 U9966 ( .C1(n8292), .C2(n8291), .A(n8290), .B(n8289), .ZN(n8293)
         );
  INV_X1 U9967 ( .A(n8293), .ZN(n8295) );
  NAND4_X1 U9968 ( .A1(n8296), .A2(n8302), .A3(n8295), .A4(n8294), .ZN(n8312)
         );
  AND2_X1 U9969 ( .A1(n8298), .A2(n8297), .ZN(n8300) );
  OAI211_X1 U9970 ( .C1(n8301), .C2(n8300), .A(n8315), .B(n8299), .ZN(n8311)
         );
  INV_X1 U9971 ( .A(n8302), .ZN(n8309) );
  OAI21_X1 U9972 ( .B1(n8304), .B2(n8589), .A(n8303), .ZN(n8305) );
  INV_X1 U9973 ( .A(n8305), .ZN(n8308) );
  OAI211_X1 U9974 ( .C1(n8309), .C2(n8308), .A(n8307), .B(n8306), .ZN(n8310)
         );
  NAND2_X1 U9975 ( .A1(n8316), .A2(n8313), .ZN(n8314) );
  NAND2_X1 U9976 ( .A1(n8314), .A2(n8317), .ZN(n8322) );
  INV_X1 U9977 ( .A(n8317), .ZN(n8318) );
  AOI21_X1 U9978 ( .B1(n8320), .B2(n8319), .A(n8318), .ZN(n8321) );
  MUX2_X1 U9979 ( .A(n8324), .B(n8323), .S(n8406), .Z(n8325) );
  INV_X1 U9980 ( .A(n8328), .ZN(n8329) );
  MUX2_X1 U9981 ( .A(n8330), .B(n8329), .S(n8406), .Z(n8331) );
  NOR2_X1 U9982 ( .A1(n8332), .A2(n8331), .ZN(n8333) );
  MUX2_X1 U9983 ( .A(n8335), .B(n8334), .S(n8406), .Z(n8336) );
  NAND2_X1 U9984 ( .A1(n8337), .A2(n8905), .ZN(n8349) );
  NAND3_X1 U9985 ( .A1(n8349), .A2(n8338), .A3(n8350), .ZN(n8339) );
  NAND2_X1 U9986 ( .A1(n8343), .A2(n8342), .ZN(n8344) );
  NAND2_X1 U9987 ( .A1(n8344), .A2(n8406), .ZN(n8345) );
  NAND3_X1 U9988 ( .A1(n8353), .A2(n8358), .A3(n8354), .ZN(n8346) );
  NAND2_X1 U9989 ( .A1(n8349), .A2(n8348), .ZN(n8351) );
  NAND3_X1 U9990 ( .A1(n8351), .A2(n8402), .A3(n8350), .ZN(n8352) );
  NAND2_X1 U9991 ( .A1(n8353), .A2(n8352), .ZN(n8356) );
  NAND3_X1 U9992 ( .A1(n8356), .A2(n8355), .A3(n8354), .ZN(n8357) );
  NAND2_X1 U9993 ( .A1(n8842), .A2(n8358), .ZN(n8361) );
  NAND2_X1 U9994 ( .A1(n8828), .A2(n8359), .ZN(n8360) );
  MUX2_X1 U9995 ( .A(n8361), .B(n8360), .S(n8406), .Z(n8362) );
  OR2_X1 U9996 ( .A1(n8363), .A2(n8406), .ZN(n8364) );
  AOI21_X1 U9997 ( .B1(n8366), .B2(n8365), .A(n8402), .ZN(n8369) );
  NOR2_X1 U9998 ( .A1(n8367), .A2(n8402), .ZN(n8368) );
  NAND2_X1 U9999 ( .A1(n8371), .A2(n8370), .ZN(n8375) );
  NAND2_X1 U10000 ( .A1(n8375), .A2(n8785), .ZN(n8372) );
  NAND2_X1 U10001 ( .A1(n8372), .A2(n8786), .ZN(n8378) );
  INV_X1 U10002 ( .A(n8784), .ZN(n8373) );
  OAI211_X1 U10003 ( .C1(n8375), .C2(n8374), .A(n8786), .B(n8373), .ZN(n8377)
         );
  MUX2_X1 U10004 ( .A(n8380), .B(n8379), .S(n8406), .Z(n8381) );
  MUX2_X1 U10005 ( .A(n8384), .B(n8383), .S(n8406), .Z(n8385) );
  NOR2_X1 U10006 ( .A1(n8386), .A2(n8385), .ZN(n8387) );
  MUX2_X1 U10007 ( .A(n8389), .B(n8388), .S(n8402), .Z(n8390) );
  INV_X1 U10008 ( .A(n8393), .ZN(n8391) );
  MUX2_X1 U10009 ( .A(n8443), .B(n8401), .S(n8402), .Z(n8392) );
  INV_X1 U10010 ( .A(n8409), .ZN(n8400) );
  INV_X1 U10011 ( .A(n8407), .ZN(n8398) );
  INV_X1 U10012 ( .A(n8395), .ZN(n8396) );
  NAND3_X1 U10013 ( .A1(n8398), .A2(n8397), .A3(n8396), .ZN(n8399) );
  AOI21_X1 U10014 ( .B1(n8401), .B2(n8400), .A(n8399), .ZN(n8414) );
  NOR2_X1 U10015 ( .A1(n8403), .A2(n8402), .ZN(n8404) );
  OAI22_X1 U10016 ( .A1(n8748), .A2(n8404), .B1(n8406), .B2(n8578), .ZN(n8413)
         );
  NOR3_X1 U10017 ( .A1(n8407), .A2(n8406), .A3(n8405), .ZN(n8408) );
  OAI21_X1 U10018 ( .B1(n8580), .B2(n8409), .A(n8408), .ZN(n8412) );
  INV_X1 U10019 ( .A(n8410), .ZN(n8411) );
  OAI211_X1 U10020 ( .C1(n8414), .C2(n8413), .A(n8412), .B(n8411), .ZN(n8416)
         );
  OAI22_X1 U10021 ( .A1(n8419), .A2(n8418), .B1(n4412), .B2(n8417), .ZN(n8421)
         );
  XNOR2_X1 U10022 ( .A(n8421), .B(n8420), .ZN(n8428) );
  NAND3_X1 U10023 ( .A1(n8423), .A2(n8422), .A3(n6107), .ZN(n8424) );
  OAI211_X1 U10024 ( .C1(n8425), .C2(n8427), .A(n8424), .B(P2_B_REG_SCAN_IN), 
        .ZN(n8426) );
  OAI21_X1 U10025 ( .B1(n8428), .B2(n8427), .A(n8426), .ZN(P2_U3296) );
  INV_X1 U10026 ( .A(n8429), .ZN(n8434) );
  OAI222_X1 U10027 ( .A1(n9824), .A2(n10303), .B1(n9822), .B2(n8434), .C1(
        P1_U3086), .C2(n5021), .ZN(P1_U3325) );
  OAI222_X1 U10028 ( .A1(n8435), .A2(n9821), .B1(n8431), .B2(P2_U3151), .C1(
        n8430), .C2(n8437), .ZN(P2_U3266) );
  OAI222_X1 U10029 ( .A1(n8437), .A2(n8436), .B1(n8435), .B2(n8434), .C1(
        P2_U3151), .C2(n8432), .ZN(P2_U3265) );
  AOI21_X1 U10030 ( .B1(n8438), .B2(n8439), .A(n8571), .ZN(n8441) );
  NAND2_X1 U10031 ( .A1(n8441), .A2(n8440), .ZN(n8446) );
  AOI22_X1 U10032 ( .A1(n8775), .A2(n8568), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3151), .ZN(n8442) );
  OAI21_X1 U10033 ( .B1(n8443), .B2(n8566), .A(n8442), .ZN(n8444) );
  AOI21_X1 U10034 ( .B1(n8757), .B2(n8558), .A(n8444), .ZN(n8445) );
  OAI211_X1 U10035 ( .C1(n8759), .C2(n8554), .A(n8446), .B(n8445), .ZN(
        P2_U3154) );
  OAI21_X1 U10036 ( .B1(n8449), .B2(n8448), .A(n8447), .ZN(n8450) );
  NAND2_X1 U10037 ( .A1(n8450), .A2(n8545), .ZN(n8458) );
  INV_X1 U10038 ( .A(n8451), .ZN(n8456) );
  INV_X1 U10039 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n8452) );
  NOR2_X1 U10040 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8452), .ZN(n8655) );
  AOI21_X1 U10041 ( .B1(n8568), .B2(n8584), .A(n8655), .ZN(n8453) );
  OAI21_X1 U10042 ( .B1(n8454), .B2(n8566), .A(n8453), .ZN(n8455) );
  AOI21_X1 U10043 ( .B1(n8456), .B2(n8558), .A(n8455), .ZN(n8457) );
  OAI211_X1 U10044 ( .C1(n8459), .C2(n8554), .A(n8458), .B(n8457), .ZN(
        P2_U3155) );
  XNOR2_X1 U10045 ( .A(n8460), .B(n8819), .ZN(n8465) );
  AOI22_X1 U10046 ( .A1(n8807), .A2(n8568), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3151), .ZN(n8462) );
  NAND2_X1 U10047 ( .A1(n8558), .A2(n8810), .ZN(n8461) );
  OAI211_X1 U10048 ( .C1(n8777), .C2(n8566), .A(n8462), .B(n8461), .ZN(n8463)
         );
  OAI21_X1 U10049 ( .B1(n8465), .B2(n8571), .A(n8464), .ZN(P2_U3156) );
  INV_X1 U10050 ( .A(n8952), .ZN(n8477) );
  INV_X1 U10051 ( .A(n8466), .ZN(n8546) );
  INV_X1 U10052 ( .A(n8467), .ZN(n8469) );
  NOR3_X1 U10053 ( .A1(n8546), .A2(n8469), .A3(n8468), .ZN(n8471) );
  INV_X1 U10054 ( .A(n8470), .ZN(n8525) );
  OAI21_X1 U10055 ( .B1(n8471), .B2(n8525), .A(n8545), .ZN(n8476) );
  NAND2_X1 U10056 ( .A1(n8568), .A2(n8881), .ZN(n8473) );
  OAI211_X1 U10057 ( .C1(n8566), .C2(n8856), .A(n8473), .B(n8472), .ZN(n8474)
         );
  AOI21_X1 U10058 ( .B1(n8861), .B2(n8558), .A(n8474), .ZN(n8475) );
  OAI211_X1 U10059 ( .C1(n8477), .C2(n8554), .A(n8476), .B(n8475), .ZN(
        P2_U3159) );
  INV_X1 U10060 ( .A(n8479), .ZN(n8526) );
  NOR3_X1 U10061 ( .A1(n8526), .A2(n4933), .A3(n8481), .ZN(n8482) );
  OAI21_X1 U10062 ( .B1(n8482), .B2(n4931), .A(n8545), .ZN(n8486) );
  AOI22_X1 U10063 ( .A1(n8568), .A2(n8581), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3151), .ZN(n8483) );
  OAI21_X1 U10064 ( .B1(n8827), .B2(n8566), .A(n8483), .ZN(n8484) );
  AOI21_X1 U10065 ( .B1(n8832), .B2(n8558), .A(n8484), .ZN(n8485) );
  OAI211_X1 U10066 ( .C1(n9009), .C2(n8554), .A(n8486), .B(n8485), .ZN(
        P2_U3163) );
  XOR2_X1 U10067 ( .A(n8488), .B(n8487), .Z(n8493) );
  AOI22_X1 U10068 ( .A1(n8775), .A2(n8548), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3151), .ZN(n8490) );
  NAND2_X1 U10069 ( .A1(n8782), .A2(n8558), .ZN(n8489) );
  OAI211_X1 U10070 ( .C1(n8777), .C2(n8550), .A(n8490), .B(n8489), .ZN(n8491)
         );
  AOI21_X1 U10071 ( .B1(n8985), .B2(n8576), .A(n8491), .ZN(n8492) );
  OAI21_X1 U10072 ( .B1(n8493), .B2(n8571), .A(n8492), .ZN(P2_U3165) );
  INV_X1 U10073 ( .A(n9031), .ZN(n8503) );
  AOI21_X1 U10074 ( .B1(n4965), .B2(n8496), .A(n8495), .ZN(n8497) );
  OAI21_X1 U10075 ( .B1(n8497), .B2(n4495), .A(n8545), .ZN(n8502) );
  INV_X1 U10076 ( .A(n8498), .ZN(n8900) );
  NAND2_X1 U10077 ( .A1(n8568), .A2(n8894), .ZN(n8499) );
  NAND2_X1 U10078 ( .A1(P2_U3151), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8689) );
  OAI211_X1 U10079 ( .C1(n8566), .C2(n8896), .A(n8499), .B(n8689), .ZN(n8500)
         );
  AOI21_X1 U10080 ( .B1(n8900), .B2(n8558), .A(n8500), .ZN(n8501) );
  OAI211_X1 U10081 ( .C1(n8503), .C2(n8554), .A(n8502), .B(n8501), .ZN(
        P2_U3166) );
  INV_X1 U10082 ( .A(n9025), .ZN(n8513) );
  NOR3_X1 U10083 ( .A1(n4495), .A2(n8505), .A3(n8504), .ZN(n8506) );
  OAI21_X1 U10084 ( .B1(n4496), .B2(n8506), .A(n8545), .ZN(n8512) );
  INV_X1 U10085 ( .A(n8507), .ZN(n8884) );
  NAND2_X1 U10086 ( .A1(n8568), .A2(n8910), .ZN(n8508) );
  NAND2_X1 U10087 ( .A1(P2_U3151), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n8710) );
  OAI211_X1 U10088 ( .C1(n8566), .C2(n8509), .A(n8508), .B(n8710), .ZN(n8510)
         );
  AOI21_X1 U10089 ( .B1(n8884), .B2(n8558), .A(n8510), .ZN(n8511) );
  OAI211_X1 U10090 ( .C1(n8513), .C2(n8554), .A(n8512), .B(n8511), .ZN(
        P2_U3168) );
  XOR2_X1 U10091 ( .A(n8515), .B(n8514), .Z(n8520) );
  AOI22_X1 U10092 ( .A1(n8793), .A2(n8548), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3151), .ZN(n8517) );
  NAND2_X1 U10093 ( .A1(n8797), .A2(n8558), .ZN(n8516) );
  OAI211_X1 U10094 ( .C1(n8539), .C2(n8550), .A(n8517), .B(n8516), .ZN(n8518)
         );
  AOI21_X1 U10095 ( .B1(n8991), .B2(n8576), .A(n8518), .ZN(n8519) );
  OAI21_X1 U10096 ( .B1(n8520), .B2(n8571), .A(n8519), .ZN(P2_U3169) );
  INV_X1 U10097 ( .A(n8522), .ZN(n8524) );
  NOR3_X1 U10098 ( .A1(n8525), .A2(n8524), .A3(n8523), .ZN(n8527) );
  OAI21_X1 U10099 ( .B1(n8527), .B2(n8526), .A(n8545), .ZN(n8531) );
  AOI22_X1 U10100 ( .A1(n8548), .A2(n8818), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3151), .ZN(n8528) );
  OAI21_X1 U10101 ( .B1(n8868), .B2(n8550), .A(n8528), .ZN(n8529) );
  AOI21_X1 U10102 ( .B1(n8844), .B2(n8558), .A(n8529), .ZN(n8530) );
  OAI211_X1 U10103 ( .C1(n9014), .C2(n8554), .A(n8531), .B(n8530), .ZN(
        P2_U3173) );
  INV_X1 U10104 ( .A(n8532), .ZN(n8534) );
  NAND2_X1 U10105 ( .A1(n8534), .A2(n8533), .ZN(n8535) );
  XNOR2_X1 U10106 ( .A(n8536), .B(n8535), .ZN(n8542) );
  AOI22_X1 U10107 ( .A1(n8818), .A2(n8568), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3151), .ZN(n8538) );
  NAND2_X1 U10108 ( .A1(n8558), .A2(n8822), .ZN(n8537) );
  OAI211_X1 U10109 ( .C1(n8539), .C2(n8566), .A(n8538), .B(n8537), .ZN(n8540)
         );
  AOI21_X1 U10110 ( .B1(n9002), .B2(n8576), .A(n8540), .ZN(n8541) );
  OAI21_X1 U10111 ( .B1(n8542), .B2(n8571), .A(n8541), .ZN(P2_U3175) );
  INV_X1 U10112 ( .A(n8956), .ZN(n8555) );
  NOR3_X1 U10113 ( .A1(n4496), .A2(n4963), .A3(n8544), .ZN(n8547) );
  OAI21_X1 U10114 ( .B1(n8547), .B2(n8546), .A(n8545), .ZN(n8553) );
  AND2_X1 U10115 ( .A1(P2_U3151), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8728) );
  AOI21_X1 U10116 ( .B1(n8548), .B2(n8582), .A(n8728), .ZN(n8549) );
  OAI21_X1 U10117 ( .B1(n8896), .B2(n8550), .A(n8549), .ZN(n8551) );
  AOI21_X1 U10118 ( .B1(n8873), .B2(n8558), .A(n8551), .ZN(n8552) );
  OAI211_X1 U10119 ( .C1(n8555), .C2(n8554), .A(n8553), .B(n8552), .ZN(
        P2_U3178) );
  XOR2_X1 U10120 ( .A(n8557), .B(n8556), .Z(n8564) );
  AOI22_X1 U10121 ( .A1(n8793), .A2(n8568), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3151), .ZN(n8560) );
  NAND2_X1 U10122 ( .A1(n8771), .A2(n8558), .ZN(n8559) );
  OAI211_X1 U10123 ( .C1(n8561), .C2(n8566), .A(n8560), .B(n8559), .ZN(n8562)
         );
  AOI21_X1 U10124 ( .B1(n8979), .B2(n8576), .A(n8562), .ZN(n8563) );
  OAI21_X1 U10125 ( .B1(n8564), .B2(n8571), .A(n8563), .ZN(P2_U3180) );
  NAND2_X1 U10126 ( .A1(P2_U3151), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8675) );
  OAI21_X1 U10127 ( .B1(n8566), .B2(n8565), .A(n8675), .ZN(n8567) );
  AOI21_X1 U10128 ( .B1(n8568), .B2(n8908), .A(n8567), .ZN(n8569) );
  OAI21_X1 U10129 ( .B1(n8915), .B2(n8570), .A(n8569), .ZN(n8575) );
  AOI211_X1 U10130 ( .C1(n8573), .C2(n8572), .A(n8571), .B(n8494), .ZN(n8574)
         );
  AOI211_X1 U10131 ( .C1(n9037), .C2(n8576), .A(n8575), .B(n8574), .ZN(n8577)
         );
  INV_X1 U10132 ( .A(n8577), .ZN(P2_U3181) );
  MUX2_X1 U10133 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n8742), .S(P2_U3893), .Z(
        P2_U3522) );
  MUX2_X1 U10134 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n8578), .S(P2_U3893), .Z(
        P2_U3521) );
  MUX2_X1 U10135 ( .A(n8579), .B(P2_DATAO_REG_29__SCAN_IN), .S(n8727), .Z(
        P2_U3520) );
  MUX2_X1 U10136 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n8580), .S(P2_U3893), .Z(
        P2_U3519) );
  MUX2_X1 U10137 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8768), .S(P2_U3893), .Z(
        P2_U3518) );
  MUX2_X1 U10138 ( .A(n8775), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8727), .Z(
        P2_U3517) );
  MUX2_X1 U10139 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8793), .S(P2_U3893), .Z(
        P2_U3516) );
  MUX2_X1 U10140 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n8806), .S(P2_U3893), .Z(
        P2_U3515) );
  MUX2_X1 U10141 ( .A(n8819), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8727), .Z(
        P2_U3514) );
  MUX2_X1 U10142 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8807), .S(P2_U3893), .Z(
        P2_U3513) );
  MUX2_X1 U10143 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8818), .S(P2_U3893), .Z(
        P2_U3512) );
  MUX2_X1 U10144 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8581), .S(P2_U3893), .Z(
        P2_U3511) );
  MUX2_X1 U10145 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8582), .S(P2_U3893), .Z(
        P2_U3510) );
  MUX2_X1 U10146 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n8881), .S(P2_U3893), .Z(
        P2_U3509) );
  MUX2_X1 U10147 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8583), .S(P2_U3893), .Z(
        P2_U3508) );
  MUX2_X1 U10148 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8910), .S(P2_U3893), .Z(
        P2_U3507) );
  MUX2_X1 U10149 ( .A(n8894), .B(P2_DATAO_REG_15__SCAN_IN), .S(n8727), .Z(
        P2_U3506) );
  MUX2_X1 U10150 ( .A(n8908), .B(P2_DATAO_REG_14__SCAN_IN), .S(n8727), .Z(
        P2_U3505) );
  MUX2_X1 U10151 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n8584), .S(P2_U3893), .Z(
        P2_U3504) );
  MUX2_X1 U10152 ( .A(n8585), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8727), .Z(
        P2_U3503) );
  MUX2_X1 U10153 ( .A(n8586), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8727), .Z(
        P2_U3501) );
  MUX2_X1 U10154 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n8587), .S(P2_U3893), .Z(
        P2_U3500) );
  MUX2_X1 U10155 ( .A(n8588), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8727), .Z(
        P2_U3499) );
  MUX2_X1 U10156 ( .A(n8589), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8727), .Z(
        P2_U3498) );
  MUX2_X1 U10157 ( .A(n8590), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8727), .Z(
        P2_U3497) );
  MUX2_X1 U10158 ( .A(n8591), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8727), .Z(
        P2_U3496) );
  MUX2_X1 U10159 ( .A(n8592), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8727), .Z(
        P2_U3495) );
  MUX2_X1 U10160 ( .A(n5772), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8727), .Z(
        P2_U3494) );
  MUX2_X1 U10161 ( .A(n5755), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8727), .Z(
        P2_U3493) );
  MUX2_X1 U10162 ( .A(n5739), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8727), .Z(
        P2_U3492) );
  OAI21_X1 U10163 ( .B1(n8595), .B2(n8594), .A(n8593), .ZN(n8596) );
  NAND2_X1 U10164 ( .A1(n8596), .A2(n9918), .ZN(n8614) );
  OAI21_X1 U10165 ( .B1(n9938), .B2(n8598), .A(n8597), .ZN(n8599) );
  AOI21_X1 U10166 ( .B1(n9934), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n8599), .ZN(
        n8613) );
  INV_X1 U10167 ( .A(n8600), .ZN(n8602) );
  NOR3_X1 U10168 ( .A1(n8603), .A2(n8602), .A3(n8601), .ZN(n8605) );
  OAI21_X1 U10169 ( .B1(n8605), .B2(n8604), .A(n8737), .ZN(n8612) );
  AND3_X1 U10170 ( .A1(n7311), .A2(n8607), .A3(n8606), .ZN(n8609) );
  OAI21_X1 U10171 ( .B1(n8610), .B2(n8609), .A(n8608), .ZN(n8611) );
  NAND4_X1 U10172 ( .A1(n8614), .A2(n8613), .A3(n8612), .A4(n8611), .ZN(
        P2_U3190) );
  AOI21_X1 U10173 ( .B1(n8617), .B2(n8616), .A(n8615), .ZN(n8632) );
  OAI21_X1 U10174 ( .B1(n8620), .B2(n8619), .A(n8618), .ZN(n8630) );
  AOI21_X1 U10175 ( .B1(n8623), .B2(n8622), .A(n8621), .ZN(n8624) );
  NOR2_X1 U10176 ( .A1(n9929), .A2(n8624), .ZN(n8625) );
  AOI211_X1 U10177 ( .C1(n8627), .C2(n8709), .A(n8626), .B(n8625), .ZN(n8628)
         );
  OAI21_X1 U10178 ( .B1(n10071), .B2(n8735), .A(n8628), .ZN(n8629) );
  AOI21_X1 U10179 ( .B1(n9918), .B2(n8630), .A(n8629), .ZN(n8631) );
  OAI21_X1 U10180 ( .B1(n8632), .B2(n9930), .A(n8631), .ZN(P2_U3194) );
  AOI21_X1 U10181 ( .B1(n5898), .B2(n8634), .A(n8633), .ZN(n8649) );
  OAI21_X1 U10182 ( .B1(n8637), .B2(n8636), .A(n8635), .ZN(n8647) );
  AOI21_X1 U10183 ( .B1(n8639), .B2(n5903), .A(n8638), .ZN(n8640) );
  NOR2_X1 U10184 ( .A1(n9929), .A2(n8640), .ZN(n8641) );
  AOI211_X1 U10185 ( .C1(n8643), .C2(n8709), .A(n8642), .B(n8641), .ZN(n8644)
         );
  OAI21_X1 U10186 ( .B1(n8645), .B2(n8735), .A(n8644), .ZN(n8646) );
  AOI21_X1 U10187 ( .B1(n9918), .B2(n8647), .A(n8646), .ZN(n8648) );
  OAI21_X1 U10188 ( .B1(n8649), .B2(n9930), .A(n8648), .ZN(P2_U3195) );
  AOI21_X1 U10189 ( .B1(n4506), .B2(n8651), .A(n8650), .ZN(n8665) );
  OAI21_X1 U10190 ( .B1(n8654), .B2(n8653), .A(n8652), .ZN(n8663) );
  AOI21_X1 U10191 ( .B1(n8709), .B2(n8656), .A(n8655), .ZN(n8657) );
  OAI21_X1 U10192 ( .B1(n10342), .B2(n8735), .A(n8657), .ZN(n8662) );
  AOI21_X1 U10193 ( .B1(n4503), .B2(n8659), .A(n8658), .ZN(n8660) );
  NOR2_X1 U10194 ( .A1(n8660), .A2(n9929), .ZN(n8661) );
  AOI211_X1 U10195 ( .C1(n9918), .C2(n8663), .A(n8662), .B(n8661), .ZN(n8664)
         );
  OAI21_X1 U10196 ( .B1(n8665), .B2(n9930), .A(n8664), .ZN(P2_U3196) );
  AOI21_X1 U10197 ( .B1(n8965), .B2(n8667), .A(n8666), .ZN(n8682) );
  OAI21_X1 U10198 ( .B1(n8670), .B2(n8669), .A(n8668), .ZN(n8680) );
  AOI21_X1 U10199 ( .B1(n8672), .B2(n8914), .A(n8671), .ZN(n8673) );
  NOR2_X1 U10200 ( .A1(n9929), .A2(n8673), .ZN(n8679) );
  NAND2_X1 U10201 ( .A1(n8709), .A2(n8674), .ZN(n8676) );
  OAI211_X1 U10202 ( .C1(n8677), .C2(n8735), .A(n8676), .B(n8675), .ZN(n8678)
         );
  AOI211_X1 U10203 ( .C1(n9918), .C2(n8680), .A(n8679), .B(n8678), .ZN(n8681)
         );
  OAI21_X1 U10204 ( .B1(n8682), .B2(n9930), .A(n8681), .ZN(P2_U3197) );
  AOI21_X1 U10205 ( .B1(n4462), .B2(n8684), .A(n8683), .ZN(n8698) );
  OAI21_X1 U10206 ( .B1(n8687), .B2(n8686), .A(n8685), .ZN(n8696) );
  NAND2_X1 U10207 ( .A1(n8709), .A2(n8688), .ZN(n8690) );
  OAI211_X1 U10208 ( .C1(n8691), .C2(n8735), .A(n8690), .B(n8689), .ZN(n8695)
         );
  NOR2_X1 U10209 ( .A1(n8693), .A2(n9930), .ZN(n8694) );
  AOI211_X1 U10210 ( .C1(n9918), .C2(n8696), .A(n8695), .B(n8694), .ZN(n8697)
         );
  OAI21_X1 U10211 ( .B1(n8698), .B2(n9929), .A(n8697), .ZN(P2_U3198) );
  AOI21_X1 U10212 ( .B1(n8959), .B2(n8700), .A(n8699), .ZN(n8718) );
  OAI21_X1 U10213 ( .B1(n8703), .B2(n8702), .A(n8701), .ZN(n8716) );
  NOR2_X1 U10214 ( .A1(n8735), .A2(n8704), .ZN(n8715) );
  NAND2_X1 U10215 ( .A1(n8709), .A2(n8708), .ZN(n8711) );
  OAI21_X1 U10216 ( .B1(n8713), .B2(n9929), .A(n8712), .ZN(n8714) );
  AOI211_X1 U10217 ( .C1(n9918), .C2(n8716), .A(n8715), .B(n8714), .ZN(n8717)
         );
  OAI21_X1 U10218 ( .B1(n8718), .B2(n9930), .A(n8717), .ZN(P2_U3199) );
  AOI21_X1 U10219 ( .B1(n8721), .B2(n8720), .A(n8719), .ZN(n8740) );
  OAI21_X1 U10220 ( .B1(n4464), .B2(n4537), .A(n8724), .ZN(n8738) );
  NAND2_X1 U10221 ( .A1(n8726), .A2(n8725), .ZN(n8732) );
  OAI21_X1 U10222 ( .B1(n8727), .B2(n8732), .A(n9938), .ZN(n8729) );
  AOI21_X1 U10223 ( .B1(n8730), .B2(n8729), .A(n8728), .ZN(n8734) );
  NAND3_X1 U10224 ( .A1(n8732), .A2(n9918), .A3(n8731), .ZN(n8733) );
  OAI211_X1 U10225 ( .C1(n8735), .C2(n10099), .A(n8734), .B(n8733), .ZN(n8736)
         );
  AOI21_X1 U10226 ( .B1(n8738), .B2(n8737), .A(n8736), .ZN(n8739) );
  OAI21_X1 U10227 ( .B1(n8740), .B2(n9929), .A(n8739), .ZN(P2_U3200) );
  NAND2_X1 U10228 ( .A1(n8923), .A2(n8918), .ZN(n8745) );
  NAND2_X1 U10229 ( .A1(n8743), .A2(n8917), .ZN(n8751) );
  INV_X1 U10230 ( .A(n8751), .ZN(n8744) );
  OAI21_X1 U10231 ( .B1(n8970), .B2(n8744), .A(n8913), .ZN(n8746) );
  OAI211_X1 U10232 ( .C1(n8205), .C2(n8913), .A(n8745), .B(n8746), .ZN(
        P2_U3202) );
  NAND2_X1 U10233 ( .A1(n9960), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n8747) );
  OAI211_X1 U10234 ( .C1(n8748), .C2(n8846), .A(n8747), .B(n8746), .ZN(
        P2_U3203) );
  NAND2_X1 U10235 ( .A1(n8749), .A2(n8913), .ZN(n8754) );
  NAND2_X1 U10236 ( .A1(n9960), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n8750) );
  NAND2_X1 U10237 ( .A1(n8751), .A2(n8750), .ZN(n8752) );
  AOI21_X1 U10238 ( .B1(n6395), .B2(n8918), .A(n8752), .ZN(n8753) );
  OAI211_X1 U10239 ( .C1(n8755), .C2(n9956), .A(n8754), .B(n8753), .ZN(
        P2_U3204) );
  INV_X1 U10240 ( .A(n8756), .ZN(n8763) );
  AOI22_X1 U10241 ( .A1(n8757), .A2(n8917), .B1(n9960), .B2(
        P2_REG2_REG_27__SCAN_IN), .ZN(n8758) );
  OAI21_X1 U10242 ( .B1(n8759), .B2(n8846), .A(n8758), .ZN(n8760) );
  AOI21_X1 U10243 ( .B1(n8761), .B2(n8848), .A(n8760), .ZN(n8762) );
  OAI21_X1 U10244 ( .B1(n8763), .B2(n9960), .A(n8762), .ZN(P2_U3206) );
  XNOR2_X1 U10245 ( .A(n8765), .B(n8764), .ZN(n8982) );
  XNOR2_X1 U10246 ( .A(n8767), .B(n8766), .ZN(n8769) );
  AOI222_X1 U10247 ( .A1(n8912), .A2(n8769), .B1(n8768), .B2(n8909), .C1(n8793), .C2(n8907), .ZN(n8977) );
  MUX2_X1 U10248 ( .A(n8770), .B(n8977), .S(n8913), .Z(n8773) );
  AOI22_X1 U10249 ( .A1(n8979), .A2(n8918), .B1(n8917), .B2(n8771), .ZN(n8772)
         );
  OAI211_X1 U10250 ( .C1(n8922), .C2(n8982), .A(n8773), .B(n8772), .ZN(
        P2_U3207) );
  NOR2_X1 U10251 ( .A1(n4671), .A2(n9944), .ZN(n8781) );
  XNOR2_X1 U10252 ( .A(n4488), .B(n8774), .ZN(n8779) );
  NAND2_X1 U10253 ( .A1(n8775), .A2(n8909), .ZN(n8776) );
  OAI21_X1 U10254 ( .B1(n8777), .B2(n9951), .A(n8776), .ZN(n8778) );
  AOI21_X1 U10255 ( .B1(n8779), .B2(n8912), .A(n8778), .ZN(n8983) );
  INV_X1 U10256 ( .A(n8983), .ZN(n8780) );
  AOI211_X1 U10257 ( .C1(n8917), .C2(n8782), .A(n8781), .B(n8780), .ZN(n8791)
         );
  OR2_X1 U10258 ( .A1(n8783), .A2(n8784), .ZN(n8799) );
  NAND2_X1 U10259 ( .A1(n8799), .A2(n8785), .ZN(n8787) );
  NAND2_X1 U10260 ( .A1(n8787), .A2(n8786), .ZN(n8789) );
  XNOR2_X1 U10261 ( .A(n8789), .B(n8788), .ZN(n8986) );
  AOI22_X1 U10262 ( .A1(n8986), .A2(n8848), .B1(P2_REG2_REG_25__SCAN_IN), .B2(
        n9960), .ZN(n8790) );
  OAI21_X1 U10263 ( .B1(n8791), .B2(n9960), .A(n8790), .ZN(P2_U3208) );
  INV_X1 U10264 ( .A(n8991), .ZN(n8792) );
  NOR2_X1 U10265 ( .A1(n8792), .A2(n9944), .ZN(n8796) );
  XNOR2_X1 U10266 ( .A(n4484), .B(n8801), .ZN(n8794) );
  AOI222_X1 U10267 ( .A1(n8912), .A2(n8794), .B1(n8819), .B2(n8907), .C1(n8793), .C2(n8909), .ZN(n8989) );
  INV_X1 U10268 ( .A(n8989), .ZN(n8795) );
  AOI211_X1 U10269 ( .C1(n8917), .C2(n8797), .A(n8796), .B(n8795), .ZN(n8803)
         );
  NAND2_X1 U10270 ( .A1(n8799), .A2(n8798), .ZN(n8800) );
  XOR2_X1 U10271 ( .A(n8801), .B(n8800), .Z(n8992) );
  AOI22_X1 U10272 ( .A1(n8992), .A2(n8848), .B1(P2_REG2_REG_24__SCAN_IN), .B2(
        n9960), .ZN(n8802) );
  OAI21_X1 U10273 ( .B1(n8803), .B2(n9960), .A(n8802), .ZN(P2_U3209) );
  XNOR2_X1 U10274 ( .A(n8783), .B(n8804), .ZN(n8997) );
  INV_X1 U10275 ( .A(n8997), .ZN(n8813) );
  INV_X1 U10276 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n8809) );
  XNOR2_X1 U10277 ( .A(n8805), .B(n8804), .ZN(n8808) );
  AOI222_X1 U10278 ( .A1(n8912), .A2(n8808), .B1(n8807), .B2(n8907), .C1(n8806), .C2(n8909), .ZN(n8995) );
  MUX2_X1 U10279 ( .A(n8809), .B(n8995), .S(n8913), .Z(n8812) );
  OAI211_X1 U10280 ( .C1(n8922), .C2(n8813), .A(n8812), .B(n8811), .ZN(
        P2_U3210) );
  XNOR2_X1 U10281 ( .A(n8815), .B(n8814), .ZN(n9005) );
  INV_X1 U10282 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n8821) );
  XNOR2_X1 U10283 ( .A(n8816), .B(n8817), .ZN(n8820) );
  AOI222_X1 U10284 ( .A1(n8912), .A2(n8820), .B1(n8819), .B2(n8909), .C1(n8818), .C2(n8907), .ZN(n9000) );
  MUX2_X1 U10285 ( .A(n8821), .B(n9000), .S(n8913), .Z(n8824) );
  AOI22_X1 U10286 ( .A1(n9002), .A2(n8918), .B1(n8917), .B2(n8822), .ZN(n8823)
         );
  OAI211_X1 U10287 ( .C1(n8922), .C2(n9005), .A(n8824), .B(n8823), .ZN(
        P2_U3211) );
  XNOR2_X1 U10288 ( .A(n8825), .B(n8830), .ZN(n8826) );
  OAI222_X1 U10289 ( .A1(n9953), .A2(n8827), .B1(n9951), .B2(n8856), .C1(n9949), .C2(n8826), .ZN(n8943) );
  INV_X1 U10290 ( .A(n8943), .ZN(n8836) );
  NAND2_X1 U10291 ( .A1(n8829), .A2(n8828), .ZN(n8831) );
  XNOR2_X1 U10292 ( .A(n8831), .B(n8830), .ZN(n8944) );
  AOI22_X1 U10293 ( .A1(n9960), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n8917), .B2(
        n8832), .ZN(n8833) );
  OAI21_X1 U10294 ( .B1(n9009), .B2(n8846), .A(n8833), .ZN(n8834) );
  AOI21_X1 U10295 ( .B1(n8944), .B2(n8848), .A(n8834), .ZN(n8835) );
  OAI21_X1 U10296 ( .B1(n8836), .B2(n9960), .A(n8835), .ZN(P2_U3212) );
  INV_X1 U10297 ( .A(n8837), .ZN(n8838) );
  AOI21_X1 U10298 ( .B1(n8842), .B2(n8839), .A(n8838), .ZN(n8840) );
  OAI222_X1 U10299 ( .A1(n9951), .A2(n8868), .B1(n9953), .B2(n8841), .C1(n9949), .C2(n8840), .ZN(n8947) );
  INV_X1 U10300 ( .A(n8947), .ZN(n8850) );
  XOR2_X1 U10301 ( .A(n8842), .B(n8843), .Z(n8948) );
  AOI22_X1 U10302 ( .A1(n9960), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n8917), .B2(
        n8844), .ZN(n8845) );
  OAI21_X1 U10303 ( .B1(n9014), .B2(n8846), .A(n8845), .ZN(n8847) );
  AOI21_X1 U10304 ( .B1(n8948), .B2(n8848), .A(n8847), .ZN(n8849) );
  OAI21_X1 U10305 ( .B1(n8850), .B2(n9960), .A(n8849), .ZN(P2_U3213) );
  OAI211_X1 U10306 ( .C1(n4659), .C2(n8853), .A(n8912), .B(n8852), .ZN(n8855)
         );
  NAND2_X1 U10307 ( .A1(n8881), .A2(n8907), .ZN(n8854) );
  OAI211_X1 U10308 ( .C1(n8856), .C2(n9953), .A(n8855), .B(n8854), .ZN(n8951)
         );
  OR2_X1 U10309 ( .A1(n8858), .A2(n8857), .ZN(n8859) );
  NAND2_X1 U10310 ( .A1(n8860), .A2(n8859), .ZN(n9018) );
  AOI22_X1 U10311 ( .A1(n9960), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n8917), .B2(
        n8861), .ZN(n8863) );
  NAND2_X1 U10312 ( .A1(n8952), .A2(n8918), .ZN(n8862) );
  OAI211_X1 U10313 ( .C1(n9018), .C2(n8922), .A(n8863), .B(n8862), .ZN(n8864)
         );
  AOI21_X1 U10314 ( .B1(n8951), .B2(n8913), .A(n8864), .ZN(n8865) );
  INV_X1 U10315 ( .A(n8865), .ZN(P2_U3214) );
  XNOR2_X1 U10316 ( .A(n8866), .B(n8870), .ZN(n8867) );
  OAI222_X1 U10317 ( .A1(n9953), .A2(n8868), .B1(n9951), .B2(n8896), .C1(n8867), .C2(n9949), .ZN(n8955) );
  NAND2_X1 U10318 ( .A1(n8869), .A2(n8870), .ZN(n8871) );
  NAND2_X1 U10319 ( .A1(n8872), .A2(n8871), .ZN(n9023) );
  AOI22_X1 U10320 ( .A1(n9960), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n8917), .B2(
        n8873), .ZN(n8875) );
  NAND2_X1 U10321 ( .A1(n8956), .A2(n8918), .ZN(n8874) );
  OAI211_X1 U10322 ( .C1(n9023), .C2(n8922), .A(n8875), .B(n8874), .ZN(n8876)
         );
  AOI21_X1 U10323 ( .B1(n8955), .B2(n8913), .A(n8876), .ZN(n8877) );
  INV_X1 U10324 ( .A(n8877), .ZN(P2_U3215) );
  XNOR2_X1 U10325 ( .A(n8878), .B(n8880), .ZN(n9026) );
  INV_X1 U10326 ( .A(n9026), .ZN(n8887) );
  XNOR2_X1 U10327 ( .A(n8879), .B(n8880), .ZN(n8882) );
  AOI222_X1 U10328 ( .A1(n8912), .A2(n8882), .B1(n8881), .B2(n8909), .C1(n8910), .C2(n8907), .ZN(n9024) );
  MUX2_X1 U10329 ( .A(n8883), .B(n9024), .S(n8913), .Z(n8886) );
  AOI22_X1 U10330 ( .A1(n9025), .A2(n8918), .B1(n8917), .B2(n8884), .ZN(n8885)
         );
  OAI211_X1 U10331 ( .C1(n8922), .C2(n8887), .A(n8886), .B(n8885), .ZN(
        P2_U3216) );
  XNOR2_X1 U10332 ( .A(n8889), .B(n8888), .ZN(n9032) );
  INV_X1 U10333 ( .A(n9032), .ZN(n8903) );
  NAND2_X1 U10334 ( .A1(n8891), .A2(n8890), .ZN(n8893) );
  XNOR2_X1 U10335 ( .A(n8893), .B(n8892), .ZN(n8898) );
  NAND2_X1 U10336 ( .A1(n8894), .A2(n8907), .ZN(n8895) );
  OAI21_X1 U10337 ( .B1(n8896), .B2(n9953), .A(n8895), .ZN(n8897) );
  AOI21_X1 U10338 ( .B1(n8898), .B2(n8912), .A(n8897), .ZN(n9029) );
  MUX2_X1 U10339 ( .A(n8899), .B(n9029), .S(n8913), .Z(n8902) );
  AOI22_X1 U10340 ( .A1(n9031), .A2(n8918), .B1(n8917), .B2(n8900), .ZN(n8901)
         );
  OAI211_X1 U10341 ( .C1(n8922), .C2(n8903), .A(n8902), .B(n8901), .ZN(
        P2_U3217) );
  XNOR2_X1 U10342 ( .A(n8904), .B(n8905), .ZN(n9039) );
  INV_X1 U10343 ( .A(n9039), .ZN(n8921) );
  XOR2_X1 U10344 ( .A(n8906), .B(n8905), .Z(n8911) );
  AOI222_X1 U10345 ( .A1(n8912), .A2(n8911), .B1(n8910), .B2(n8909), .C1(n8908), .C2(n8907), .ZN(n9035) );
  MUX2_X1 U10346 ( .A(n8914), .B(n9035), .S(n8913), .Z(n8920) );
  INV_X1 U10347 ( .A(n8915), .ZN(n8916) );
  AOI22_X1 U10348 ( .A1(n9037), .A2(n8918), .B1(n8917), .B2(n8916), .ZN(n8919)
         );
  OAI211_X1 U10349 ( .C1(n8922), .C2(n8921), .A(n8920), .B(n8919), .ZN(
        P2_U3218) );
  NAND2_X1 U10350 ( .A1(n8923), .A2(n8966), .ZN(n8924) );
  NAND2_X1 U10351 ( .A1(n8970), .A2(n10029), .ZN(n8925) );
  OAI211_X1 U10352 ( .C1(n10029), .C2(n8209), .A(n8924), .B(n8925), .ZN(
        P2_U3490) );
  NAND2_X1 U10353 ( .A1(n8973), .A2(n8966), .ZN(n8926) );
  OAI211_X1 U10354 ( .C1(n10029), .C2(n8927), .A(n8926), .B(n8925), .ZN(
        P2_U3489) );
  INV_X1 U10355 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n8928) );
  MUX2_X1 U10356 ( .A(n8928), .B(n8977), .S(n10029), .Z(n8930) );
  NAND2_X1 U10357 ( .A1(n8979), .A2(n8966), .ZN(n8929) );
  OAI211_X1 U10358 ( .C1(n8982), .C2(n8958), .A(n8930), .B(n8929), .ZN(
        P2_U3485) );
  MUX2_X1 U10359 ( .A(n8931), .B(n8983), .S(n10029), .Z(n8933) );
  AOI22_X1 U10360 ( .A1(n8986), .A2(n8967), .B1(n8966), .B2(n8985), .ZN(n8932)
         );
  NAND2_X1 U10361 ( .A1(n8933), .A2(n8932), .ZN(P2_U3484) );
  INV_X1 U10362 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n8934) );
  MUX2_X1 U10363 ( .A(n8934), .B(n8989), .S(n10029), .Z(n8936) );
  AOI22_X1 U10364 ( .A1(n8992), .A2(n8967), .B1(n8966), .B2(n8991), .ZN(n8935)
         );
  NAND2_X1 U10365 ( .A1(n8936), .A2(n8935), .ZN(P2_U3483) );
  MUX2_X1 U10366 ( .A(n8937), .B(n8995), .S(n10029), .Z(n8939) );
  NAND2_X1 U10367 ( .A1(n8939), .A2(n8938), .ZN(P2_U3482) );
  INV_X1 U10368 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n8940) );
  MUX2_X1 U10369 ( .A(n8940), .B(n9000), .S(n10029), .Z(n8942) );
  NAND2_X1 U10370 ( .A1(n9002), .A2(n8966), .ZN(n8941) );
  OAI211_X1 U10371 ( .C1(n9005), .C2(n8958), .A(n8942), .B(n8941), .ZN(
        P2_U3481) );
  INV_X1 U10372 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n8945) );
  AOI21_X1 U10373 ( .B1(n8944), .B2(n9970), .A(n8943), .ZN(n9006) );
  MUX2_X1 U10374 ( .A(n8945), .B(n9006), .S(n10029), .Z(n8946) );
  OAI21_X1 U10375 ( .B1(n9009), .B2(n8950), .A(n8946), .ZN(P2_U3480) );
  AOI21_X1 U10376 ( .B1(n9970), .B2(n8948), .A(n8947), .ZN(n9010) );
  MUX2_X1 U10377 ( .A(n10195), .B(n9010), .S(n10029), .Z(n8949) );
  OAI21_X1 U10378 ( .B1(n9014), .B2(n8950), .A(n8949), .ZN(P2_U3479) );
  AOI21_X1 U10379 ( .B1(n10015), .B2(n8952), .A(n8951), .ZN(n9015) );
  MUX2_X1 U10380 ( .A(n8953), .B(n9015), .S(n10029), .Z(n8954) );
  OAI21_X1 U10381 ( .B1(n8958), .B2(n9018), .A(n8954), .ZN(P2_U3478) );
  AOI21_X1 U10382 ( .B1(n10015), .B2(n8956), .A(n8955), .ZN(n9019) );
  MUX2_X1 U10383 ( .A(n10276), .B(n9019), .S(n10029), .Z(n8957) );
  OAI21_X1 U10384 ( .B1(n8958), .B2(n9023), .A(n8957), .ZN(P2_U3477) );
  MUX2_X1 U10385 ( .A(n8959), .B(n9024), .S(n10029), .Z(n8961) );
  AOI22_X1 U10386 ( .A1(n9026), .A2(n8967), .B1(n8966), .B2(n9025), .ZN(n8960)
         );
  NAND2_X1 U10387 ( .A1(n8961), .A2(n8960), .ZN(P2_U3476) );
  MUX2_X1 U10388 ( .A(n8962), .B(n9029), .S(n10029), .Z(n8964) );
  AOI22_X1 U10389 ( .A1(n9032), .A2(n8967), .B1(n8966), .B2(n9031), .ZN(n8963)
         );
  NAND2_X1 U10390 ( .A1(n8964), .A2(n8963), .ZN(P2_U3475) );
  MUX2_X1 U10391 ( .A(n8965), .B(n9035), .S(n10029), .Z(n8969) );
  AOI22_X1 U10392 ( .A1(n9039), .A2(n8967), .B1(n8966), .B2(n9037), .ZN(n8968)
         );
  NAND2_X1 U10393 ( .A1(n8969), .A2(n8968), .ZN(P2_U3474) );
  NAND2_X1 U10394 ( .A1(n8970), .A2(n10016), .ZN(n8974) );
  NAND2_X1 U10395 ( .A1(n10017), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n8971) );
  OAI211_X1 U10396 ( .C1(n8972), .C2(n9013), .A(n8974), .B(n8971), .ZN(
        P2_U3458) );
  INV_X1 U10397 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n8976) );
  NAND2_X1 U10398 ( .A1(n8973), .A2(n6396), .ZN(n8975) );
  OAI211_X1 U10399 ( .C1(n8976), .C2(n10016), .A(n8975), .B(n8974), .ZN(
        P2_U3457) );
  INV_X1 U10400 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n8978) );
  MUX2_X1 U10401 ( .A(n8978), .B(n8977), .S(n10016), .Z(n8981) );
  NAND2_X1 U10402 ( .A1(n8979), .A2(n6396), .ZN(n8980) );
  OAI211_X1 U10403 ( .C1(n8982), .C2(n9022), .A(n8981), .B(n8980), .ZN(
        P2_U3453) );
  INV_X1 U10404 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n8984) );
  MUX2_X1 U10405 ( .A(n8984), .B(n8983), .S(n10016), .Z(n8988) );
  AOI22_X1 U10406 ( .A1(n8986), .A2(n9038), .B1(n6396), .B2(n8985), .ZN(n8987)
         );
  NAND2_X1 U10407 ( .A1(n8988), .A2(n8987), .ZN(P2_U3452) );
  INV_X1 U10408 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n8990) );
  MUX2_X1 U10409 ( .A(n8990), .B(n8989), .S(n10016), .Z(n8994) );
  AOI22_X1 U10410 ( .A1(n8992), .A2(n9038), .B1(n6396), .B2(n8991), .ZN(n8993)
         );
  NAND2_X1 U10411 ( .A1(n8994), .A2(n8993), .ZN(P2_U3451) );
  INV_X1 U10412 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n8996) );
  MUX2_X1 U10413 ( .A(n8996), .B(n8995), .S(n10016), .Z(n8999) );
  NAND2_X1 U10414 ( .A1(n8999), .A2(n8998), .ZN(P2_U3450) );
  INV_X1 U10415 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n9001) );
  MUX2_X1 U10416 ( .A(n9001), .B(n9000), .S(n10016), .Z(n9004) );
  NAND2_X1 U10417 ( .A1(n9002), .A2(n6396), .ZN(n9003) );
  OAI211_X1 U10418 ( .C1(n9005), .C2(n9022), .A(n9004), .B(n9003), .ZN(
        P2_U3449) );
  INV_X1 U10419 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n9007) );
  MUX2_X1 U10420 ( .A(n9007), .B(n9006), .S(n10016), .Z(n9008) );
  OAI21_X1 U10421 ( .B1(n9009), .B2(n9013), .A(n9008), .ZN(P2_U3448) );
  MUX2_X1 U10422 ( .A(n9011), .B(n9010), .S(n10016), .Z(n9012) );
  OAI21_X1 U10423 ( .B1(n9014), .B2(n9013), .A(n9012), .ZN(P2_U3447) );
  MUX2_X1 U10424 ( .A(n9016), .B(n9015), .S(n10016), .Z(n9017) );
  OAI21_X1 U10425 ( .B1(n9018), .B2(n9022), .A(n9017), .ZN(P2_U3446) );
  MUX2_X1 U10426 ( .A(n9020), .B(n9019), .S(n10016), .Z(n9021) );
  OAI21_X1 U10427 ( .B1(n9023), .B2(n9022), .A(n9021), .ZN(P2_U3444) );
  MUX2_X1 U10428 ( .A(n10086), .B(n9024), .S(n10016), .Z(n9028) );
  AOI22_X1 U10429 ( .A1(n9026), .A2(n9038), .B1(n6396), .B2(n9025), .ZN(n9027)
         );
  NAND2_X1 U10430 ( .A1(n9028), .A2(n9027), .ZN(P2_U3441) );
  INV_X1 U10431 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n9030) );
  MUX2_X1 U10432 ( .A(n9030), .B(n9029), .S(n10016), .Z(n9034) );
  AOI22_X1 U10433 ( .A1(n9032), .A2(n9038), .B1(n6396), .B2(n9031), .ZN(n9033)
         );
  NAND2_X1 U10434 ( .A1(n9034), .A2(n9033), .ZN(P2_U3438) );
  INV_X1 U10435 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n9036) );
  MUX2_X1 U10436 ( .A(n9036), .B(n9035), .S(n10016), .Z(n9041) );
  AOI22_X1 U10437 ( .A1(n9039), .A2(n9038), .B1(n6396), .B2(n9037), .ZN(n9040)
         );
  NAND2_X1 U10438 ( .A1(n9041), .A2(n9040), .ZN(P2_U3435) );
  NAND3_X1 U10439 ( .A1(n9042), .A2(P2_STATE_REG_SCAN_IN), .A3(
        P2_IR_REG_31__SCAN_IN), .ZN(n9047) );
  NAND2_X1 U10440 ( .A1(n9812), .A2(n9043), .ZN(n9046) );
  NAND2_X1 U10441 ( .A1(n9044), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n9045) );
  OAI211_X1 U10442 ( .C1(n9048), .C2(n9047), .A(n9046), .B(n9045), .ZN(
        P2_U3264) );
  MUX2_X1 U10443 ( .A(n9049), .B(n9911), .S(P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  INV_X1 U10444 ( .A(n9051), .ZN(n9052) );
  AOI21_X1 U10445 ( .B1(n9053), .B2(n9050), .A(n9052), .ZN(n9061) );
  NOR2_X1 U10446 ( .A1(n9227), .A2(n9134), .ZN(n9054) );
  AOI211_X1 U10447 ( .C1(n9225), .C2(n9253), .A(n9055), .B(n9054), .ZN(n9056)
         );
  OAI21_X1 U10448 ( .B1(n9057), .B2(n9239), .A(n9056), .ZN(n9058) );
  AOI21_X1 U10449 ( .B1(n9059), .B2(n9209), .A(n9058), .ZN(n9060) );
  OAI21_X1 U10450 ( .B1(n9061), .B2(n9205), .A(n9060), .ZN(P1_U3215) );
  NAND2_X1 U10451 ( .A1(n4504), .A2(n9062), .ZN(n9063) );
  XNOR2_X1 U10452 ( .A(n9064), .B(n9063), .ZN(n9069) );
  AOI22_X1 U10453 ( .A1(n9244), .A2(n9469), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        P1_U3086), .ZN(n9066) );
  NAND2_X1 U10454 ( .A1(n9225), .A2(n9532), .ZN(n9065) );
  OAI211_X1 U10455 ( .C1(n9503), .C2(n9239), .A(n9066), .B(n9065), .ZN(n9067)
         );
  AOI21_X1 U10456 ( .B1(n9685), .B2(n9209), .A(n9067), .ZN(n9068) );
  OAI21_X1 U10457 ( .B1(n9069), .B2(n9205), .A(n9068), .ZN(P1_U3216) );
  XNOR2_X1 U10458 ( .A(n9070), .B(n9071), .ZN(n9213) );
  NAND2_X1 U10459 ( .A1(n9213), .A2(n9214), .ZN(n9212) );
  NAND2_X1 U10460 ( .A1(n9070), .A2(n9072), .ZN(n9076) );
  AND2_X1 U10461 ( .A1(n9212), .A2(n9076), .ZN(n9078) );
  INV_X1 U10462 ( .A(n9073), .ZN(n9074) );
  XNOR2_X1 U10463 ( .A(n9075), .B(n9074), .ZN(n9077) );
  NAND3_X1 U10464 ( .A1(n9212), .A2(n9077), .A3(n9076), .ZN(n9176) );
  OAI211_X1 U10465 ( .C1(n9078), .C2(n9077), .A(n9236), .B(n9176), .ZN(n9082)
         );
  NAND2_X1 U10466 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9390) );
  OAI21_X1 U10467 ( .B1(n9227), .B2(n9524), .A(n9390), .ZN(n9080) );
  NOR2_X1 U10468 ( .A1(n9239), .A2(n9568), .ZN(n9079) );
  AOI211_X1 U10469 ( .C1(n9225), .C2(n9610), .A(n9080), .B(n9079), .ZN(n9081)
         );
  OAI211_X1 U10470 ( .C1(n9571), .C2(n9247), .A(n9082), .B(n9081), .ZN(
        P1_U3219) );
  NAND2_X1 U10471 ( .A1(n9649), .A2(n6587), .ZN(n9084) );
  OR2_X1 U10472 ( .A1(n6589), .A2(n9432), .ZN(n9083) );
  NAND2_X1 U10473 ( .A1(n9084), .A2(n9083), .ZN(n9086) );
  XNOR2_X1 U10474 ( .A(n9086), .B(n9085), .ZN(n9090) );
  NAND2_X1 U10475 ( .A1(n9649), .A2(n9087), .ZN(n9088) );
  OAI21_X1 U10476 ( .B1(n9432), .B2(n6418), .A(n9088), .ZN(n9089) );
  XNOR2_X1 U10477 ( .A(n9090), .B(n9089), .ZN(n9097) );
  INV_X1 U10478 ( .A(n9097), .ZN(n9092) );
  INV_X1 U10479 ( .A(n9098), .ZN(n9091) );
  NAND3_X1 U10480 ( .A1(n9093), .A2(n9236), .A3(n9097), .ZN(n9101) );
  AOI22_X1 U10481 ( .A1(n9244), .A2(n9410), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3086), .ZN(n9095) );
  NAND2_X1 U10482 ( .A1(n9225), .A2(n9648), .ZN(n9094) );
  OAI211_X1 U10483 ( .C1(n9239), .C2(n9413), .A(n9095), .B(n9094), .ZN(n9096)
         );
  AOI21_X1 U10484 ( .B1(n9649), .B2(n9209), .A(n9096), .ZN(n9100) );
  NAND3_X1 U10485 ( .A1(n9098), .A2(n9236), .A3(n9097), .ZN(n9099) );
  NAND4_X1 U10486 ( .A1(n9102), .A2(n9101), .A3(n9100), .A4(n9099), .ZN(
        P1_U3220) );
  AOI22_X1 U10487 ( .A1(n4417), .A2(n9209), .B1(n9244), .B2(n9264), .ZN(n9110)
         );
  AOI22_X1 U10488 ( .A1(n9225), .A2(n6414), .B1(n9104), .B2(
        P1_REG3_REG_1__SCAN_IN), .ZN(n9109) );
  OAI21_X1 U10489 ( .B1(n9106), .B2(n4999), .A(n9105), .ZN(n9107) );
  NAND2_X1 U10490 ( .A1(n9107), .A2(n9236), .ZN(n9108) );
  NAND3_X1 U10491 ( .A1(n9110), .A2(n9109), .A3(n9108), .ZN(P1_U3222) );
  OAI21_X1 U10492 ( .B1(n9113), .B2(n9112), .A(n9111), .ZN(n9114) );
  NAND2_X1 U10493 ( .A1(n9114), .A2(n9236), .ZN(n9119) );
  INV_X1 U10494 ( .A(n9537), .ZN(n9117) );
  AOI22_X1 U10495 ( .A1(n9244), .A2(n9532), .B1(P1_REG3_REG_21__SCAN_IN), .B2(
        P1_U3086), .ZN(n9115) );
  OAI21_X1 U10496 ( .B1(n9524), .B2(n9241), .A(n9115), .ZN(n9116) );
  AOI21_X1 U10497 ( .B1(n9117), .B2(n9229), .A(n9116), .ZN(n9118) );
  OAI211_X1 U10498 ( .C1(n9536), .C2(n9247), .A(n9119), .B(n9118), .ZN(
        P1_U3223) );
  OAI21_X1 U10499 ( .B1(n9121), .B2(n9120), .A(n9221), .ZN(n9122) );
  NAND2_X1 U10500 ( .A1(n9122), .A2(n9236), .ZN(n9126) );
  OAI22_X1 U10501 ( .A1(n9227), .A2(n9657), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10058), .ZN(n9124) );
  NOR2_X1 U10502 ( .A1(n9239), .A2(n9466), .ZN(n9123) );
  AOI211_X1 U10503 ( .C1(n9225), .C2(n9469), .A(n9124), .B(n9123), .ZN(n9125)
         );
  OAI211_X1 U10504 ( .C1(n9669), .C2(n9247), .A(n9126), .B(n9125), .ZN(
        P1_U3225) );
  NAND2_X1 U10505 ( .A1(n4734), .A2(n9129), .ZN(n9130) );
  XNOR2_X1 U10506 ( .A(n9127), .B(n9130), .ZN(n9137) );
  NOR2_X1 U10507 ( .A1(n9131), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9351) );
  AOI21_X1 U10508 ( .B1(n9244), .B2(n9625), .A(n9351), .ZN(n9133) );
  NAND2_X1 U10509 ( .A1(n9229), .A2(n9631), .ZN(n9132) );
  OAI211_X1 U10510 ( .C1(n9241), .C2(n9134), .A(n9133), .B(n9132), .ZN(n9135)
         );
  AOI21_X1 U10511 ( .B1(n9801), .B2(n9209), .A(n9135), .ZN(n9136) );
  OAI21_X1 U10512 ( .B1(n9137), .B2(n9205), .A(n9136), .ZN(P1_U3226) );
  XNOR2_X1 U10513 ( .A(n9139), .B(n9138), .ZN(n9140) );
  XNOR2_X1 U10514 ( .A(n4437), .B(n9140), .ZN(n9151) );
  NAND2_X1 U10515 ( .A1(n9229), .A2(n9141), .ZN(n9145) );
  NAND2_X1 U10516 ( .A1(n9142), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9144) );
  MUX2_X1 U10517 ( .A(n9145), .B(n9144), .S(n9143), .Z(n9148) );
  NAND2_X1 U10518 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9873) );
  INV_X1 U10519 ( .A(n9873), .ZN(n9146) );
  AOI21_X1 U10520 ( .B1(n9244), .B2(n9610), .A(n9146), .ZN(n9147) );
  OAI211_X1 U10521 ( .C1(n9607), .C2(n9241), .A(n9148), .B(n9147), .ZN(n9149)
         );
  AOI21_X1 U10522 ( .B1(n9724), .B2(n9209), .A(n9149), .ZN(n9150) );
  OAI21_X1 U10523 ( .B1(n9151), .B2(n9205), .A(n9150), .ZN(P1_U3228) );
  OAI21_X1 U10524 ( .B1(n9154), .B2(n9153), .A(n9152), .ZN(n9155) );
  NAND2_X1 U10525 ( .A1(n9155), .A2(n9236), .ZN(n9159) );
  OAI22_X1 U10526 ( .A1(n9227), .A2(n9478), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10098), .ZN(n9157) );
  NOR2_X1 U10527 ( .A1(n9239), .A2(n9484), .ZN(n9156) );
  AOI211_X1 U10528 ( .C1(n9225), .C2(n9675), .A(n9157), .B(n9156), .ZN(n9158)
         );
  OAI211_X1 U10529 ( .C1(n4683), .C2(n9247), .A(n9159), .B(n9158), .ZN(
        P1_U3229) );
  NAND2_X1 U10530 ( .A1(n9244), .A2(n9256), .ZN(n9163) );
  NAND2_X1 U10531 ( .A1(n9225), .A2(n9258), .ZN(n9162) );
  NAND2_X1 U10532 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_U3086), .ZN(n9836) );
  NAND2_X1 U10533 ( .A1(n9229), .A2(n9160), .ZN(n9161) );
  NAND4_X1 U10534 ( .A1(n9163), .A2(n9162), .A3(n9836), .A4(n9161), .ZN(n9172)
         );
  AOI21_X1 U10535 ( .B1(n9165), .B2(n7836), .A(n9164), .ZN(n9169) );
  XNOR2_X1 U10536 ( .A(n9167), .B(n9166), .ZN(n9168) );
  XNOR2_X1 U10537 ( .A(n9169), .B(n9168), .ZN(n9170) );
  NOR2_X1 U10538 ( .A1(n9170), .A2(n9205), .ZN(n9171) );
  AOI211_X1 U10539 ( .C1(n9173), .C2(n9209), .A(n9172), .B(n9171), .ZN(n9174)
         );
  INV_X1 U10540 ( .A(n9174), .ZN(P1_U3231) );
  NAND2_X1 U10541 ( .A1(n9176), .A2(n9175), .ZN(n9180) );
  NOR2_X1 U10542 ( .A1(n9178), .A2(n9177), .ZN(n9179) );
  XNOR2_X1 U10543 ( .A(n9180), .B(n9179), .ZN(n9185) );
  AOI22_X1 U10544 ( .A1(n9244), .A2(n9545), .B1(P1_REG3_REG_20__SCAN_IN), .B2(
        P1_U3086), .ZN(n9182) );
  NAND2_X1 U10545 ( .A1(n9225), .A2(n9554), .ZN(n9181) );
  OAI211_X1 U10546 ( .C1(n9239), .C2(n9551), .A(n9182), .B(n9181), .ZN(n9183)
         );
  AOI21_X1 U10547 ( .B1(n9703), .B2(n9209), .A(n9183), .ZN(n9184) );
  OAI21_X1 U10548 ( .B1(n9185), .B2(n9205), .A(n9184), .ZN(P1_U3233) );
  NOR2_X1 U10549 ( .A1(n9186), .A2(n4450), .ZN(n9188) );
  XNOR2_X1 U10550 ( .A(n9188), .B(n9187), .ZN(n9193) );
  AOI22_X1 U10551 ( .A1(n9244), .A2(n9675), .B1(P1_REG3_REG_22__SCAN_IN), .B2(
        P1_U3086), .ZN(n9190) );
  NAND2_X1 U10552 ( .A1(n9225), .A2(n9545), .ZN(n9189) );
  OAI211_X1 U10553 ( .C1(n9239), .C2(n9510), .A(n9190), .B(n9189), .ZN(n9191)
         );
  AOI21_X1 U10554 ( .B1(n9509), .B2(n9209), .A(n9191), .ZN(n9192) );
  OAI21_X1 U10555 ( .B1(n9193), .B2(n9205), .A(n9192), .ZN(P1_U3235) );
  NAND2_X1 U10556 ( .A1(n9244), .A2(n9254), .ZN(n9198) );
  NAND2_X1 U10557 ( .A1(n9225), .A2(n9256), .ZN(n9197) );
  NAND2_X1 U10558 ( .A1(n9229), .A2(n9194), .ZN(n9195) );
  NAND4_X1 U10559 ( .A1(n9198), .A2(n9197), .A3(n9196), .A4(n9195), .ZN(n9208)
         );
  OAI21_X1 U10560 ( .B1(n7909), .B2(n9200), .A(n9199), .ZN(n9204) );
  XNOR2_X1 U10561 ( .A(n9202), .B(n9201), .ZN(n9203) );
  XNOR2_X1 U10562 ( .A(n9204), .B(n9203), .ZN(n9206) );
  NOR2_X1 U10563 ( .A1(n9206), .A2(n9205), .ZN(n9207) );
  AOI211_X1 U10564 ( .C1(n9210), .C2(n9209), .A(n9208), .B(n9207), .ZN(n9211)
         );
  INV_X1 U10565 ( .A(n9211), .ZN(P1_U3236) );
  OAI21_X1 U10566 ( .B1(n9214), .B2(n9213), .A(n9212), .ZN(n9215) );
  NAND2_X1 U10567 ( .A1(n9215), .A2(n9236), .ZN(n9219) );
  NAND2_X1 U10568 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9362) );
  OAI21_X1 U10569 ( .B1(n9227), .B2(n9706), .A(n9362), .ZN(n9217) );
  NOR2_X1 U10570 ( .A1(n9239), .A2(n9582), .ZN(n9216) );
  AOI211_X1 U10571 ( .C1(n9225), .C2(n9625), .A(n9217), .B(n9216), .ZN(n9218)
         );
  OAI211_X1 U10572 ( .C1(n9586), .C2(n9247), .A(n9219), .B(n9218), .ZN(
        P1_U3238) );
  AND2_X1 U10573 ( .A1(n9221), .A2(n9220), .ZN(n9224) );
  OAI211_X1 U10574 ( .C1(n9224), .C2(n9223), .A(n9236), .B(n9222), .ZN(n9232)
         );
  INV_X1 U10575 ( .A(n9448), .ZN(n9230) );
  AOI22_X1 U10576 ( .A1(n9225), .A2(n9251), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3086), .ZN(n9226) );
  OAI21_X1 U10577 ( .B1(n9441), .B2(n9227), .A(n9226), .ZN(n9228) );
  AOI21_X1 U10578 ( .B1(n9230), .B2(n9229), .A(n9228), .ZN(n9231) );
  OAI211_X1 U10579 ( .C1(n9452), .C2(n9247), .A(n9232), .B(n9231), .ZN(
        P1_U3240) );
  OAI21_X1 U10580 ( .B1(n9235), .B2(n9234), .A(n9233), .ZN(n9237) );
  NAND2_X1 U10581 ( .A1(n9237), .A2(n9236), .ZN(n9246) );
  NOR2_X1 U10582 ( .A1(n9239), .A2(n9238), .ZN(n9243) );
  NAND2_X1 U10583 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9327) );
  OAI21_X1 U10584 ( .B1(n9241), .B2(n9240), .A(n9327), .ZN(n9242) );
  AOI211_X1 U10585 ( .C1(n9244), .C2(n9722), .A(n9243), .B(n9242), .ZN(n9245)
         );
  OAI211_X1 U10586 ( .C1(n9248), .C2(n9247), .A(n9246), .B(n9245), .ZN(
        P1_U3241) );
  MUX2_X1 U10587 ( .A(n9394), .B(P1_DATAO_REG_31__SCAN_IN), .S(n10054), .Z(
        P1_U3585) );
  MUX2_X1 U10588 ( .A(n9249), .B(P1_DATAO_REG_30__SCAN_IN), .S(n10054), .Z(
        P1_U3584) );
  MUX2_X1 U10589 ( .A(n9410), .B(P1_DATAO_REG_29__SCAN_IN), .S(n10054), .Z(
        P1_U3583) );
  MUX2_X1 U10590 ( .A(n9250), .B(P1_DATAO_REG_28__SCAN_IN), .S(n10054), .Z(
        P1_U3582) );
  MUX2_X1 U10591 ( .A(n9648), .B(P1_DATAO_REG_27__SCAN_IN), .S(n10054), .Z(
        P1_U3581) );
  MUX2_X1 U10592 ( .A(n5524), .B(P1_DATAO_REG_26__SCAN_IN), .S(n10054), .Z(
        P1_U3580) );
  MUX2_X1 U10593 ( .A(n9251), .B(P1_DATAO_REG_25__SCAN_IN), .S(n10054), .Z(
        P1_U3579) );
  MUX2_X1 U10594 ( .A(n9469), .B(P1_DATAO_REG_24__SCAN_IN), .S(n10054), .Z(
        P1_U3578) );
  MUX2_X1 U10595 ( .A(n9675), .B(P1_DATAO_REG_23__SCAN_IN), .S(n10054), .Z(
        P1_U3577) );
  MUX2_X1 U10596 ( .A(n9532), .B(P1_DATAO_REG_22__SCAN_IN), .S(n10054), .Z(
        P1_U3576) );
  MUX2_X1 U10597 ( .A(n9545), .B(P1_DATAO_REG_21__SCAN_IN), .S(n10054), .Z(
        P1_U3575) );
  MUX2_X1 U10598 ( .A(n9695), .B(P1_DATAO_REG_20__SCAN_IN), .S(n10054), .Z(
        P1_U3574) );
  MUX2_X1 U10599 ( .A(n9554), .B(P1_DATAO_REG_19__SCAN_IN), .S(n10054), .Z(
        P1_U3573) );
  MUX2_X1 U10600 ( .A(n9625), .B(P1_DATAO_REG_17__SCAN_IN), .S(n10054), .Z(
        P1_U3571) );
  MUX2_X1 U10601 ( .A(n9722), .B(P1_DATAO_REG_16__SCAN_IN), .S(n10054), .Z(
        P1_U3570) );
  MUX2_X1 U10602 ( .A(n9624), .B(P1_DATAO_REG_15__SCAN_IN), .S(n10054), .Z(
        P1_U3569) );
  MUX2_X1 U10603 ( .A(n9252), .B(P1_DATAO_REG_14__SCAN_IN), .S(n10054), .Z(
        P1_U3568) );
  MUX2_X1 U10604 ( .A(n9253), .B(P1_DATAO_REG_13__SCAN_IN), .S(n10054), .Z(
        P1_U3567) );
  MUX2_X1 U10605 ( .A(n9254), .B(P1_DATAO_REG_12__SCAN_IN), .S(n10054), .Z(
        P1_U3566) );
  MUX2_X1 U10606 ( .A(n9255), .B(P1_DATAO_REG_11__SCAN_IN), .S(n10054), .Z(
        P1_U3565) );
  MUX2_X1 U10607 ( .A(n9256), .B(P1_DATAO_REG_10__SCAN_IN), .S(n10054), .Z(
        P1_U3564) );
  MUX2_X1 U10608 ( .A(n9257), .B(P1_DATAO_REG_9__SCAN_IN), .S(n10054), .Z(
        P1_U3563) );
  MUX2_X1 U10609 ( .A(n9258), .B(P1_DATAO_REG_8__SCAN_IN), .S(n10054), .Z(
        P1_U3562) );
  MUX2_X1 U10610 ( .A(n9259), .B(P1_DATAO_REG_7__SCAN_IN), .S(n10054), .Z(
        P1_U3561) );
  MUX2_X1 U10611 ( .A(n9260), .B(P1_DATAO_REG_6__SCAN_IN), .S(n10054), .Z(
        P1_U3560) );
  MUX2_X1 U10612 ( .A(n9261), .B(P1_DATAO_REG_5__SCAN_IN), .S(n10054), .Z(
        P1_U3559) );
  MUX2_X1 U10613 ( .A(n9262), .B(P1_DATAO_REG_4__SCAN_IN), .S(n10054), .Z(
        P1_U3558) );
  MUX2_X1 U10614 ( .A(n9263), .B(P1_DATAO_REG_3__SCAN_IN), .S(n10054), .Z(
        P1_U3557) );
  MUX2_X1 U10615 ( .A(n9264), .B(P1_DATAO_REG_2__SCAN_IN), .S(n10054), .Z(
        P1_U3556) );
  MUX2_X1 U10616 ( .A(n6427), .B(P1_DATAO_REG_1__SCAN_IN), .S(n10054), .Z(
        P1_U3555) );
  MUX2_X1 U10617 ( .A(n6414), .B(P1_DATAO_REG_0__SCAN_IN), .S(n10054), .Z(
        P1_U3554) );
  INV_X1 U10618 ( .A(n9265), .ZN(n9268) );
  NOR2_X1 U10619 ( .A1(n9866), .A2(n9266), .ZN(n9267) );
  AOI211_X1 U10620 ( .C1(n9352), .C2(P1_ADDR_REG_5__SCAN_IN), .A(n9268), .B(
        n9267), .ZN(n9278) );
  OAI211_X1 U10621 ( .C1(n9271), .C2(n9270), .A(n9872), .B(n9269), .ZN(n9277)
         );
  INV_X1 U10622 ( .A(n9272), .ZN(n9288) );
  NAND3_X1 U10623 ( .A1(n9846), .A2(n9274), .A3(n9273), .ZN(n9275) );
  NAND3_X1 U10624 ( .A1(n9386), .A2(n9288), .A3(n9275), .ZN(n9276) );
  NAND3_X1 U10625 ( .A1(n9278), .A2(n9277), .A3(n9276), .ZN(P1_U3248) );
  NOR2_X1 U10626 ( .A1(n9866), .A2(n9285), .ZN(n9279) );
  AOI211_X1 U10627 ( .C1(n9352), .C2(P1_ADDR_REG_6__SCAN_IN), .A(n9280), .B(
        n9279), .ZN(n9292) );
  OAI211_X1 U10628 ( .C1(n9283), .C2(n9282), .A(n9872), .B(n9281), .ZN(n9291)
         );
  INV_X1 U10629 ( .A(n9284), .ZN(n9287) );
  MUX2_X1 U10630 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n6998), .S(n9285), .Z(n9286)
         );
  NAND3_X1 U10631 ( .A1(n9288), .A2(n9287), .A3(n9286), .ZN(n9289) );
  NAND3_X1 U10632 ( .A1(n9386), .A2(n9302), .A3(n9289), .ZN(n9290) );
  NAND3_X1 U10633 ( .A1(n9292), .A2(n9291), .A3(n9290), .ZN(P1_U3249) );
  INV_X1 U10634 ( .A(n9293), .ZN(n9296) );
  NOR2_X1 U10635 ( .A1(n9866), .A2(n9294), .ZN(n9295) );
  AOI211_X1 U10636 ( .C1(n9352), .C2(P1_ADDR_REG_7__SCAN_IN), .A(n9296), .B(
        n9295), .ZN(n9307) );
  OAI211_X1 U10637 ( .C1(n9299), .C2(n9298), .A(n9297), .B(n9872), .ZN(n9306)
         );
  INV_X1 U10638 ( .A(n9317), .ZN(n9304) );
  NAND3_X1 U10639 ( .A1(n9302), .A2(n9301), .A3(n9300), .ZN(n9303) );
  NAND3_X1 U10640 ( .A1(n9386), .A2(n9304), .A3(n9303), .ZN(n9305) );
  NAND3_X1 U10641 ( .A1(n9307), .A2(n9306), .A3(n9305), .ZN(P1_U3250) );
  INV_X1 U10642 ( .A(n9308), .ZN(n9311) );
  NOR2_X1 U10643 ( .A1(n9866), .A2(n9309), .ZN(n9310) );
  AOI211_X1 U10644 ( .C1(n9352), .C2(P1_ADDR_REG_8__SCAN_IN), .A(n9311), .B(
        n9310), .ZN(n9322) );
  OAI211_X1 U10645 ( .C1(n9314), .C2(n9313), .A(n9312), .B(n9872), .ZN(n9321)
         );
  OR3_X1 U10646 ( .A1(n9317), .A2(n9316), .A3(n9315), .ZN(n9318) );
  NAND3_X1 U10647 ( .A1(n9386), .A2(n9319), .A3(n9318), .ZN(n9320) );
  NAND3_X1 U10648 ( .A1(n9322), .A2(n9321), .A3(n9320), .ZN(P1_U3251) );
  INV_X1 U10649 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n10251) );
  NOR2_X1 U10650 ( .A1(n10251), .A2(n9325), .ZN(n9345) );
  AOI211_X1 U10651 ( .C1(n10251), .C2(n9325), .A(n9345), .B(n9844), .ZN(n9326)
         );
  INV_X1 U10652 ( .A(n9326), .ZN(n9336) );
  INV_X1 U10653 ( .A(n9866), .ZN(n9329) );
  OAI21_X1 U10654 ( .B1(n9875), .B2(n7722), .A(n9327), .ZN(n9328) );
  AOI21_X1 U10655 ( .B1(n9338), .B2(n9329), .A(n9328), .ZN(n9335) );
  OAI21_X1 U10656 ( .B1(n9332), .B2(n9331), .A(n9330), .ZN(n9337) );
  XNOR2_X1 U10657 ( .A(n9343), .B(n9337), .ZN(n9333) );
  NAND2_X1 U10658 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(n9333), .ZN(n9339) );
  OAI211_X1 U10659 ( .C1(P1_REG1_REG_15__SCAN_IN), .C2(n9333), .A(n9386), .B(
        n9339), .ZN(n9334) );
  NAND3_X1 U10660 ( .A1(n9336), .A2(n9335), .A3(n9334), .ZN(P1_U3258) );
  NAND2_X1 U10661 ( .A1(n9338), .A2(n9337), .ZN(n9340) );
  NAND2_X1 U10662 ( .A1(n9340), .A2(n9339), .ZN(n9342) );
  XNOR2_X1 U10663 ( .A(n9365), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n9341) );
  NOR2_X1 U10664 ( .A1(n9341), .A2(n9342), .ZN(n9356) );
  AOI21_X1 U10665 ( .B1(n9342), .B2(n9341), .A(n9356), .ZN(n9355) );
  NOR2_X1 U10666 ( .A1(n9344), .A2(n9343), .ZN(n9346) );
  NOR2_X1 U10667 ( .A1(n9346), .A2(n9345), .ZN(n9348) );
  AOI22_X1 U10668 ( .A1(n9365), .A2(n10147), .B1(P1_REG2_REG_16__SCAN_IN), 
        .B2(n9358), .ZN(n9347) );
  NOR2_X1 U10669 ( .A1(n9348), .A2(n9347), .ZN(n9364) );
  AOI211_X1 U10670 ( .C1(n9348), .C2(n9347), .A(n9364), .B(n9844), .ZN(n9349)
         );
  INV_X1 U10671 ( .A(n9349), .ZN(n9354) );
  NOR2_X1 U10672 ( .A1(n9866), .A2(n9358), .ZN(n9350) );
  AOI211_X1 U10673 ( .C1(n9352), .C2(P1_ADDR_REG_16__SCAN_IN), .A(n9351), .B(
        n9350), .ZN(n9353) );
  OAI211_X1 U10674 ( .C1(n9355), .C2(n9869), .A(n9354), .B(n9353), .ZN(
        P1_U3259) );
  INV_X1 U10675 ( .A(n9381), .ZN(n9376) );
  XNOR2_X1 U10676 ( .A(n9381), .B(P1_REG1_REG_18__SCAN_IN), .ZN(n9361) );
  XNOR2_X1 U10677 ( .A(n9859), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n9864) );
  AOI21_X1 U10678 ( .B1(n9358), .B2(n9357), .A(n9356), .ZN(n9865) );
  NOR2_X1 U10679 ( .A1(n9864), .A2(n9865), .ZN(n9863) );
  NOR2_X1 U10680 ( .A1(n9859), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n9359) );
  OR2_X1 U10681 ( .A1(n9863), .A2(n9359), .ZN(n9360) );
  NOR3_X1 U10682 ( .A1(n9863), .A2(n9361), .A3(n9359), .ZN(n9380) );
  AOI211_X1 U10683 ( .C1(n9361), .C2(n9360), .A(n9380), .B(n9869), .ZN(n9374)
         );
  INV_X1 U10684 ( .A(n9362), .ZN(n9373) );
  INV_X1 U10685 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n9363) );
  NOR2_X1 U10686 ( .A1(n9875), .A2(n9363), .ZN(n9372) );
  NAND2_X1 U10687 ( .A1(n9861), .A2(n4596), .ZN(n9366) );
  NAND2_X1 U10688 ( .A1(n9367), .A2(n9366), .ZN(n9370) );
  NAND2_X1 U10689 ( .A1(n9381), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9377) );
  OR2_X1 U10690 ( .A1(n9381), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9368) );
  NAND2_X1 U10691 ( .A1(n9377), .A2(n9368), .ZN(n9369) );
  AOI211_X1 U10692 ( .C1(n9370), .C2(n9369), .A(n9378), .B(n9844), .ZN(n9371)
         );
  NOR4_X1 U10693 ( .A1(n9374), .A2(n9373), .A3(n9372), .A4(n9371), .ZN(n9375)
         );
  OAI21_X1 U10694 ( .B1(n9376), .B2(n9866), .A(n9375), .ZN(P1_U3261) );
  AOI21_X1 U10695 ( .B1(P1_REG1_REG_18__SCAN_IN), .B2(n9381), .A(n9380), .ZN(
        n9382) );
  XNOR2_X1 U10696 ( .A(n9382), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n9385) );
  OAI21_X1 U10697 ( .B1(n9385), .B2(n9869), .A(n9866), .ZN(n9383) );
  AOI21_X1 U10698 ( .B1(n9384), .B2(n9872), .A(n9383), .ZN(n9389) );
  AOI22_X1 U10699 ( .A1(n9387), .A2(n9872), .B1(n9386), .B2(n9385), .ZN(n9388)
         );
  MUX2_X1 U10700 ( .A(n9389), .B(n9388), .S(n4519), .Z(n9391) );
  OAI211_X1 U10701 ( .C1(n4852), .C2(n9875), .A(n9391), .B(n9390), .ZN(
        P1_U3262) );
  XNOR2_X1 U10702 ( .A(n9399), .B(n9752), .ZN(n9392) );
  NOR2_X1 U10703 ( .A1(n9392), .A2(n9567), .ZN(n9638) );
  NAND2_X1 U10704 ( .A1(n9638), .A2(n9578), .ZN(n9398) );
  AND2_X1 U10705 ( .A1(n9394), .A2(n9393), .ZN(n9395) );
  AND2_X1 U10706 ( .A1(n9881), .A2(n9395), .ZN(n9641) );
  INV_X1 U10707 ( .A(n9641), .ZN(n9396) );
  NOR2_X1 U10708 ( .A1(n9889), .A2(n9396), .ZN(n9402) );
  AOI21_X1 U10709 ( .B1(n9889), .B2(P1_REG2_REG_31__SCAN_IN), .A(n9402), .ZN(
        n9397) );
  OAI211_X1 U10710 ( .C1(n9752), .C2(n9585), .A(n9398), .B(n9397), .ZN(
        P1_U3263) );
  AOI211_X1 U10711 ( .C1(n9401), .C2(n9400), .A(n9567), .B(n9399), .ZN(n9642)
         );
  NAND2_X1 U10712 ( .A1(n9642), .A2(n9578), .ZN(n9404) );
  AOI21_X1 U10713 ( .B1(n9889), .B2(P1_REG2_REG_30__SCAN_IN), .A(n9402), .ZN(
        n9403) );
  OAI211_X1 U10714 ( .C1(n9756), .C2(n9585), .A(n9404), .B(n9403), .ZN(
        P1_U3264) );
  NAND2_X1 U10715 ( .A1(n9429), .A2(n9405), .ZN(n9408) );
  INV_X1 U10716 ( .A(n9406), .ZN(n9407) );
  AOI211_X1 U10717 ( .C1(n9411), .C2(n9408), .A(n9498), .B(n9407), .ZN(n9409)
         );
  AOI21_X1 U10718 ( .B1(n9881), .B2(n9410), .A(n9409), .ZN(n9647) );
  NAND3_X1 U10719 ( .A1(n9646), .A2(n9645), .A3(n9446), .ZN(n9421) );
  INV_X1 U10720 ( .A(n9413), .ZN(n9414) );
  AOI22_X1 U10721 ( .A1(n9889), .A2(P1_REG2_REG_28__SCAN_IN), .B1(n9414), .B2(
        n9632), .ZN(n9415) );
  OAI21_X1 U10722 ( .B1(n9441), .B2(n9606), .A(n9415), .ZN(n9419) );
  INV_X1 U10723 ( .A(n9416), .ZN(n9417) );
  OAI211_X1 U10724 ( .C1(n4679), .C2(n4444), .A(n9417), .B(n9628), .ZN(n9651)
         );
  NOR2_X1 U10725 ( .A1(n9651), .A2(n9489), .ZN(n9418) );
  AOI211_X1 U10726 ( .C1(n9620), .C2(n9649), .A(n9419), .B(n9418), .ZN(n9420)
         );
  OAI211_X1 U10727 ( .C1(n9889), .C2(n9647), .A(n9421), .B(n9420), .ZN(
        P1_U3265) );
  XNOR2_X1 U10728 ( .A(n9422), .B(n4457), .ZN(n9761) );
  INV_X1 U10729 ( .A(n9423), .ZN(n9451) );
  AOI211_X1 U10730 ( .C1(n9424), .C2(n9451), .A(n9567), .B(n4444), .ZN(n9661)
         );
  NAND2_X1 U10731 ( .A1(n9424), .A2(n9620), .ZN(n9427) );
  AOI22_X1 U10732 ( .A1(n9889), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n9425), .B2(
        n9632), .ZN(n9426) );
  OAI211_X1 U10733 ( .C1(n9657), .C2(n9606), .A(n9427), .B(n9426), .ZN(n9428)
         );
  AOI21_X1 U10734 ( .B1(n9661), .B2(n9578), .A(n9428), .ZN(n9436) );
  OAI21_X1 U10735 ( .B1(n4457), .B2(n9430), .A(n9429), .ZN(n9431) );
  NAND2_X1 U10736 ( .A1(n9431), .A2(n9893), .ZN(n9434) );
  OR2_X1 U10737 ( .A1(n9432), .A2(n9591), .ZN(n9433) );
  NAND2_X1 U10738 ( .A1(n9434), .A2(n9433), .ZN(n9660) );
  NAND2_X1 U10739 ( .A1(n9660), .A2(n9560), .ZN(n9435) );
  OAI211_X1 U10740 ( .C1(n9761), .C2(n9637), .A(n9436), .B(n9435), .ZN(
        P1_U3266) );
  NAND2_X1 U10741 ( .A1(n9459), .A2(n9437), .ZN(n9438) );
  NAND2_X1 U10742 ( .A1(n9438), .A2(n9444), .ZN(n9440) );
  NAND2_X1 U10743 ( .A1(n9440), .A2(n9439), .ZN(n9443) );
  OAI22_X1 U10744 ( .A1(n9705), .A2(n9478), .B1(n9441), .B2(n9591), .ZN(n9442)
         );
  AOI21_X1 U10745 ( .B1(n9443), .B2(n9893), .A(n9442), .ZN(n9665) );
  XOR2_X1 U10746 ( .A(n9445), .B(n9444), .Z(n9766) );
  INV_X1 U10747 ( .A(n9766), .ZN(n9447) );
  NAND2_X1 U10748 ( .A1(n9447), .A2(n9446), .ZN(n9456) );
  OAI22_X1 U10749 ( .A1(n9560), .A2(n9449), .B1(n9448), .B2(n9886), .ZN(n9454)
         );
  INV_X1 U10750 ( .A(n9450), .ZN(n9463) );
  OAI211_X1 U10751 ( .C1(n9452), .C2(n9463), .A(n9451), .B(n9628), .ZN(n9664)
         );
  NOR2_X1 U10752 ( .A1(n9664), .A2(n9489), .ZN(n9453) );
  AOI211_X1 U10753 ( .C1(n9620), .C2(n9764), .A(n9454), .B(n9453), .ZN(n9455)
         );
  OAI211_X1 U10754 ( .C1(n9889), .C2(n9665), .A(n9456), .B(n9455), .ZN(
        P1_U3267) );
  XNOR2_X1 U10755 ( .A(n9458), .B(n9457), .ZN(n9770) );
  OAI211_X1 U10756 ( .C1(n9461), .C2(n9460), .A(n9459), .B(n9893), .ZN(n9462)
         );
  OAI21_X1 U10757 ( .B1(n9657), .B2(n9591), .A(n9462), .ZN(n9671) );
  INV_X1 U10758 ( .A(n9483), .ZN(n9464) );
  AOI211_X1 U10759 ( .C1(n9465), .C2(n9464), .A(n9567), .B(n9463), .ZN(n9672)
         );
  NAND2_X1 U10760 ( .A1(n9672), .A2(n9578), .ZN(n9471) );
  OAI22_X1 U10761 ( .A1(n9560), .A2(n9467), .B1(n9466), .B2(n9886), .ZN(n9468)
         );
  AOI21_X1 U10762 ( .B1(n9555), .B2(n9469), .A(n9468), .ZN(n9470) );
  OAI211_X1 U10763 ( .C1(n9669), .C2(n9585), .A(n9471), .B(n9470), .ZN(n9472)
         );
  AOI21_X1 U10764 ( .B1(n9560), .B2(n9671), .A(n9472), .ZN(n9473) );
  OAI21_X1 U10765 ( .B1(n9770), .B2(n9637), .A(n9473), .ZN(P1_U3268) );
  XNOR2_X1 U10766 ( .A(n9474), .B(n9476), .ZN(n9774) );
  OR2_X1 U10767 ( .A1(n9494), .A2(n9475), .ZN(n9477) );
  XNOR2_X1 U10768 ( .A(n9477), .B(n9476), .ZN(n9480) );
  NOR2_X1 U10769 ( .A1(n9478), .A2(n9591), .ZN(n9479) );
  AOI21_X1 U10770 ( .B1(n9480), .B2(n9893), .A(n9479), .ZN(n9680) );
  INV_X1 U10771 ( .A(n9680), .ZN(n9491) );
  NAND2_X1 U10772 ( .A1(n9676), .A2(n9501), .ZN(n9481) );
  NAND2_X1 U10773 ( .A1(n9481), .A2(n9628), .ZN(n9482) );
  OR2_X1 U10774 ( .A1(n9483), .A2(n9482), .ZN(n9678) );
  NOR2_X1 U10775 ( .A1(n9606), .A2(n9519), .ZN(n9487) );
  OAI22_X1 U10776 ( .A1(n9560), .A2(n9485), .B1(n9484), .B2(n9886), .ZN(n9486)
         );
  AOI211_X1 U10777 ( .C1(n9676), .C2(n9620), .A(n9487), .B(n9486), .ZN(n9488)
         );
  OAI21_X1 U10778 ( .B1(n9678), .B2(n9489), .A(n9488), .ZN(n9490) );
  AOI21_X1 U10779 ( .B1(n9491), .B2(n9560), .A(n9490), .ZN(n9492) );
  OAI21_X1 U10780 ( .B1(n9774), .B2(n9637), .A(n9492), .ZN(P1_U3269) );
  XNOR2_X1 U10781 ( .A(n9493), .B(n9496), .ZN(n9687) );
  AOI22_X1 U10782 ( .A1(n9685), .A2(n9620), .B1(n9889), .B2(
        P1_REG2_REG_23__SCAN_IN), .ZN(n9507) );
  AOI21_X1 U10783 ( .B1(n9496), .B2(n9495), .A(n9494), .ZN(n9497) );
  OAI222_X1 U10784 ( .A1(n9591), .A2(n9668), .B1(n9705), .B2(n9499), .C1(n9498), .C2(n9497), .ZN(n9683) );
  INV_X1 U10785 ( .A(n9501), .ZN(n9502) );
  AOI211_X1 U10786 ( .C1(n9685), .C2(n4687), .A(n9567), .B(n9502), .ZN(n9684)
         );
  INV_X1 U10787 ( .A(n9684), .ZN(n9504) );
  OAI22_X1 U10788 ( .A1(n9504), .A2(n5666), .B1(n9503), .B2(n9886), .ZN(n9505)
         );
  OAI21_X1 U10789 ( .B1(n9683), .B2(n9505), .A(n9560), .ZN(n9506) );
  OAI211_X1 U10790 ( .C1(n9687), .C2(n9637), .A(n9507), .B(n9506), .ZN(
        P1_U3270) );
  XNOR2_X1 U10791 ( .A(n9508), .B(n9517), .ZN(n9779) );
  AOI211_X1 U10792 ( .C1(n9509), .C2(n9535), .A(n9567), .B(n9500), .ZN(n9692)
         );
  NAND2_X1 U10793 ( .A1(n9509), .A2(n9620), .ZN(n9513) );
  INV_X1 U10794 ( .A(n9510), .ZN(n9511) );
  AOI22_X1 U10795 ( .A1(n9889), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n9511), .B2(
        n9632), .ZN(n9512) );
  OAI211_X1 U10796 ( .C1(n9688), .C2(n9606), .A(n9513), .B(n9512), .ZN(n9514)
         );
  AOI21_X1 U10797 ( .B1(n9692), .B2(n9615), .A(n9514), .ZN(n9521) );
  OAI211_X1 U10798 ( .C1(n9517), .C2(n9516), .A(n9515), .B(n9893), .ZN(n9518)
         );
  OAI21_X1 U10799 ( .B1(n9519), .B2(n9591), .A(n9518), .ZN(n9691) );
  NAND2_X1 U10800 ( .A1(n9691), .A2(n9560), .ZN(n9520) );
  OAI211_X1 U10801 ( .C1(n9779), .C2(n9637), .A(n9521), .B(n9520), .ZN(
        P1_U3271) );
  XOR2_X1 U10802 ( .A(n9528), .B(n9522), .Z(n9783) );
  OAI22_X1 U10803 ( .A1(n9606), .A2(n9524), .B1(n9523), .B2(n9560), .ZN(n9525)
         );
  AOI21_X1 U10804 ( .B1(n9696), .B2(n9620), .A(n9525), .ZN(n9540) );
  NAND2_X1 U10805 ( .A1(n9544), .A2(n9543), .ZN(n9542) );
  NAND2_X1 U10806 ( .A1(n9542), .A2(n9527), .ZN(n9530) );
  INV_X1 U10807 ( .A(n9528), .ZN(n9529) );
  XNOR2_X1 U10808 ( .A(n9530), .B(n9529), .ZN(n9531) );
  NAND2_X1 U10809 ( .A1(n9531), .A2(n9893), .ZN(n9534) );
  NAND2_X1 U10810 ( .A1(n9881), .A2(n9532), .ZN(n9533) );
  NAND2_X1 U10811 ( .A1(n9534), .A2(n9533), .ZN(n9700) );
  OAI211_X1 U10812 ( .C1(n9536), .C2(n9550), .A(n9628), .B(n9535), .ZN(n9698)
         );
  OAI22_X1 U10813 ( .A1(n9698), .A2(n5666), .B1(n9886), .B2(n9537), .ZN(n9538)
         );
  OAI21_X1 U10814 ( .B1(n9700), .B2(n9538), .A(n9560), .ZN(n9539) );
  OAI211_X1 U10815 ( .C1(n9783), .C2(n9637), .A(n9540), .B(n9539), .ZN(
        P1_U3272) );
  XNOR2_X1 U10816 ( .A(n9541), .B(n9543), .ZN(n9787) );
  INV_X1 U10817 ( .A(n9787), .ZN(n9562) );
  OAI211_X1 U10818 ( .C1(n9544), .C2(n9543), .A(n9542), .B(n9893), .ZN(n9547)
         );
  NAND2_X1 U10819 ( .A1(n9881), .A2(n9545), .ZN(n9546) );
  NAND2_X1 U10820 ( .A1(n9547), .A2(n9546), .ZN(n9709) );
  NAND2_X1 U10821 ( .A1(n9565), .A2(n9703), .ZN(n9548) );
  NAND2_X1 U10822 ( .A1(n9548), .A2(n9628), .ZN(n9549) );
  NOR2_X1 U10823 ( .A1(n9550), .A2(n9549), .ZN(n9708) );
  NAND2_X1 U10824 ( .A1(n9708), .A2(n9578), .ZN(n9557) );
  OAI22_X1 U10825 ( .A1(n9560), .A2(n9552), .B1(n9551), .B2(n9886), .ZN(n9553)
         );
  AOI21_X1 U10826 ( .B1(n9555), .B2(n9554), .A(n9553), .ZN(n9556) );
  OAI211_X1 U10827 ( .C1(n9558), .C2(n9585), .A(n9557), .B(n9556), .ZN(n9559)
         );
  AOI21_X1 U10828 ( .B1(n9709), .B2(n9560), .A(n9559), .ZN(n9561) );
  OAI21_X1 U10829 ( .B1(n9562), .B2(n9637), .A(n9561), .ZN(P1_U3273) );
  XNOR2_X1 U10830 ( .A(n9563), .B(n9564), .ZN(n9717) );
  INV_X1 U10831 ( .A(n9565), .ZN(n9566) );
  AOI211_X1 U10832 ( .C1(n9714), .C2(n9581), .A(n9567), .B(n9566), .ZN(n9713)
         );
  INV_X1 U10833 ( .A(n9568), .ZN(n9569) );
  AOI22_X1 U10834 ( .A1(n9889), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9569), .B2(
        n9632), .ZN(n9570) );
  OAI21_X1 U10835 ( .B1(n9571), .B2(n9585), .A(n9570), .ZN(n9577) );
  OAI21_X1 U10836 ( .B1(n9574), .B2(n9573), .A(n9572), .ZN(n9575) );
  AOI222_X1 U10837 ( .A1(n9893), .A2(n9575), .B1(n9695), .B2(n9881), .C1(n9610), .C2(n9723), .ZN(n9716) );
  NOR2_X1 U10838 ( .A1(n9716), .A2(n9889), .ZN(n9576) );
  AOI211_X1 U10839 ( .C1(n9713), .C2(n9578), .A(n9577), .B(n9576), .ZN(n9579)
         );
  OAI21_X1 U10840 ( .B1(n9717), .B2(n9637), .A(n9579), .ZN(P1_U3274) );
  XNOR2_X1 U10841 ( .A(n9580), .B(n9587), .ZN(n9794) );
  OAI211_X1 U10842 ( .C1(n9586), .C2(n9601), .A(n9581), .B(n9628), .ZN(n9718)
         );
  INV_X1 U10843 ( .A(n9718), .ZN(n9597) );
  INV_X1 U10844 ( .A(n9582), .ZN(n9583) );
  AOI22_X1 U10845 ( .A1(n9889), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9583), .B2(
        n9632), .ZN(n9584) );
  OAI21_X1 U10846 ( .B1(n9586), .B2(n9585), .A(n9584), .ZN(n9596) );
  NAND2_X1 U10847 ( .A1(n9588), .A2(n9587), .ZN(n9589) );
  NAND2_X1 U10848 ( .A1(n9590), .A2(n9589), .ZN(n9594) );
  OAI22_X1 U10849 ( .A1(n9705), .A2(n9592), .B1(n9706), .B2(n9591), .ZN(n9593)
         );
  AOI21_X1 U10850 ( .B1(n9594), .B2(n9893), .A(n9593), .ZN(n9719) );
  NOR2_X1 U10851 ( .A1(n9719), .A2(n9889), .ZN(n9595) );
  AOI211_X1 U10852 ( .C1(n9597), .C2(n9615), .A(n9596), .B(n9595), .ZN(n9598)
         );
  OAI21_X1 U10853 ( .B1(n9794), .B2(n9637), .A(n9598), .ZN(P1_U3275) );
  XNOR2_X1 U10854 ( .A(n9599), .B(n9608), .ZN(n9798) );
  OAI21_X1 U10855 ( .B1(n4497), .B2(n9600), .A(n9628), .ZN(n9602) );
  OR2_X1 U10856 ( .A1(n9602), .A2(n9601), .ZN(n9725) );
  INV_X1 U10857 ( .A(n9725), .ZN(n9616) );
  NAND2_X1 U10858 ( .A1(n9724), .A2(n9620), .ZN(n9605) );
  AOI22_X1 U10859 ( .A1(n9889), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9603), .B2(
        n9632), .ZN(n9604) );
  OAI211_X1 U10860 ( .C1(n9607), .C2(n9606), .A(n9605), .B(n9604), .ZN(n9614)
         );
  XNOR2_X1 U10861 ( .A(n9609), .B(n9608), .ZN(n9612) );
  AND2_X1 U10862 ( .A1(n9610), .A2(n9881), .ZN(n9611) );
  AOI21_X1 U10863 ( .B1(n9612), .B2(n9893), .A(n9611), .ZN(n9727) );
  NOR2_X1 U10864 ( .A1(n9727), .A2(n9889), .ZN(n9613) );
  AOI211_X1 U10865 ( .C1(n9616), .C2(n9615), .A(n9614), .B(n9613), .ZN(n9617)
         );
  OAI21_X1 U10866 ( .B1(n9798), .B2(n9637), .A(n9617), .ZN(P1_U3276) );
  XNOR2_X1 U10867 ( .A(n9619), .B(n9618), .ZN(n9804) );
  AOI22_X1 U10868 ( .A1(n9801), .A2(n9620), .B1(n9889), .B2(
        P1_REG2_REG_16__SCAN_IN), .ZN(n9636) );
  OAI21_X1 U10869 ( .B1(n9623), .B2(n9622), .A(n9621), .ZN(n9626) );
  AOI222_X1 U10870 ( .A1(n9893), .A2(n9626), .B1(n9625), .B2(n9881), .C1(n9624), .C2(n9723), .ZN(n9732) );
  NAND2_X1 U10871 ( .A1(n9627), .A2(n9801), .ZN(n9629) );
  NAND2_X1 U10872 ( .A1(n9629), .A2(n9628), .ZN(n9630) );
  NOR2_X1 U10873 ( .A1(n4497), .A2(n9630), .ZN(n9730) );
  AOI22_X1 U10874 ( .A1(n9730), .A2(n4519), .B1(n9632), .B2(n9631), .ZN(n9633)
         );
  AOI21_X1 U10875 ( .B1(n9732), .B2(n9633), .A(n9889), .ZN(n9634) );
  INV_X1 U10876 ( .A(n9634), .ZN(n9635) );
  OAI211_X1 U10877 ( .C1(n9804), .C2(n9637), .A(n9636), .B(n9635), .ZN(
        P1_U3277) );
  NOR2_X1 U10878 ( .A1(n9638), .A2(n9641), .ZN(n9749) );
  MUX2_X1 U10879 ( .A(n9639), .B(n9749), .S(n9910), .Z(n9640) );
  OAI21_X1 U10880 ( .B1(n9752), .B2(n9644), .A(n9640), .ZN(P1_U3553) );
  NOR2_X1 U10881 ( .A1(n9642), .A2(n9641), .ZN(n9753) );
  MUX2_X1 U10882 ( .A(n5645), .B(n9753), .S(n9910), .Z(n9643) );
  OAI21_X1 U10883 ( .B1(n9756), .B2(n9644), .A(n9643), .ZN(P1_U3552) );
  INV_X1 U10884 ( .A(n9645), .ZN(n9656) );
  AOI22_X1 U10885 ( .A1(n9649), .A2(n9745), .B1(n9723), .B2(n9648), .ZN(n9650)
         );
  OAI21_X1 U10886 ( .B1(n9656), .B2(n9655), .A(n9654), .ZN(n9757) );
  MUX2_X1 U10887 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9757), .S(n9910), .Z(
        P1_U3550) );
  OAI22_X1 U10888 ( .A1(n9658), .A2(n9899), .B1(n9657), .B2(n9705), .ZN(n9659)
         );
  NOR3_X1 U10889 ( .A1(n9661), .A2(n9660), .A3(n9659), .ZN(n9758) );
  MUX2_X1 U10890 ( .A(n9662), .B(n9758), .S(n9910), .Z(n9663) );
  OAI21_X1 U10891 ( .B1(n9761), .B2(n9736), .A(n9663), .ZN(P1_U3549) );
  NAND2_X1 U10892 ( .A1(n9665), .A2(n9664), .ZN(n9762) );
  MUX2_X1 U10893 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9762), .S(n9910), .Z(n9666) );
  AOI21_X1 U10894 ( .B1(n9734), .B2(n9764), .A(n9666), .ZN(n9667) );
  OAI21_X1 U10895 ( .B1(n9766), .B2(n9736), .A(n9667), .ZN(P1_U3548) );
  OAI22_X1 U10896 ( .A1(n9669), .A2(n9899), .B1(n9668), .B2(n9705), .ZN(n9670)
         );
  NOR3_X1 U10897 ( .A1(n9672), .A2(n9671), .A3(n9670), .ZN(n9767) );
  MUX2_X1 U10898 ( .A(n9673), .B(n9767), .S(n9910), .Z(n9674) );
  OAI21_X1 U10899 ( .B1(n9770), .B2(n9736), .A(n9674), .ZN(P1_U3547) );
  AOI22_X1 U10900 ( .A1(n9676), .A2(n9745), .B1(n9723), .B2(n9675), .ZN(n9677)
         );
  AND2_X1 U10901 ( .A1(n9678), .A2(n9677), .ZN(n9679) );
  AND2_X1 U10902 ( .A1(n9680), .A2(n9679), .ZN(n9772) );
  MUX2_X1 U10903 ( .A(n9772), .B(n9681), .S(n9908), .Z(n9682) );
  OAI21_X1 U10904 ( .B1(n9774), .B2(n9736), .A(n9682), .ZN(P1_U3546) );
  INV_X1 U10905 ( .A(n9903), .ZN(n9747) );
  AOI211_X1 U10906 ( .C1(n9745), .C2(n9685), .A(n9684), .B(n9683), .ZN(n9686)
         );
  OAI21_X1 U10907 ( .B1(n9687), .B2(n9747), .A(n9686), .ZN(n9775) );
  MUX2_X1 U10908 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9775), .S(n9910), .Z(
        P1_U3545) );
  INV_X1 U10909 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n9693) );
  OAI22_X1 U10910 ( .A1(n9689), .A2(n9899), .B1(n9688), .B2(n9705), .ZN(n9690)
         );
  NOR3_X1 U10911 ( .A1(n9692), .A2(n9691), .A3(n9690), .ZN(n9776) );
  MUX2_X1 U10912 ( .A(n9693), .B(n9776), .S(n9910), .Z(n9694) );
  OAI21_X1 U10913 ( .B1(n9779), .B2(n9736), .A(n9694), .ZN(P1_U3544) );
  AOI22_X1 U10914 ( .A1(n9696), .A2(n9745), .B1(n9723), .B2(n9695), .ZN(n9697)
         );
  NAND2_X1 U10915 ( .A1(n9698), .A2(n9697), .ZN(n9699) );
  NOR2_X1 U10916 ( .A1(n9700), .A2(n9699), .ZN(n9780) );
  MUX2_X1 U10917 ( .A(n9701), .B(n9780), .S(n9910), .Z(n9702) );
  OAI21_X1 U10918 ( .B1(n9783), .B2(n9736), .A(n9702), .ZN(P1_U3543) );
  NAND2_X1 U10919 ( .A1(n9703), .A2(n9745), .ZN(n9704) );
  OAI21_X1 U10920 ( .B1(n9706), .B2(n9705), .A(n9704), .ZN(n9707) );
  MUX2_X1 U10921 ( .A(n9784), .B(P1_REG1_REG_20__SCAN_IN), .S(n9908), .Z(n9710) );
  AOI21_X1 U10922 ( .B1(n9787), .B2(n9711), .A(n9710), .ZN(n9712) );
  INV_X1 U10923 ( .A(n9712), .ZN(P1_U3542) );
  AOI21_X1 U10924 ( .B1(n9745), .B2(n9714), .A(n9713), .ZN(n9715) );
  OAI211_X1 U10925 ( .C1(n9717), .C2(n9747), .A(n9716), .B(n9715), .ZN(n9789)
         );
  MUX2_X1 U10926 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9789), .S(n9910), .Z(
        P1_U3541) );
  NAND2_X1 U10927 ( .A1(n9719), .A2(n9718), .ZN(n9790) );
  MUX2_X1 U10928 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9790), .S(n9910), .Z(n9720) );
  AOI21_X1 U10929 ( .B1(n9734), .B2(n9792), .A(n9720), .ZN(n9721) );
  OAI21_X1 U10930 ( .B1(n9794), .B2(n9736), .A(n9721), .ZN(P1_U3540) );
  AOI22_X1 U10931 ( .A1(n9724), .A2(n9745), .B1(n9723), .B2(n9722), .ZN(n9726)
         );
  AND3_X1 U10932 ( .A1(n9727), .A2(n9726), .A3(n9725), .ZN(n9795) );
  MUX2_X1 U10933 ( .A(n9728), .B(n9795), .S(n9910), .Z(n9729) );
  OAI21_X1 U10934 ( .B1(n9798), .B2(n9736), .A(n9729), .ZN(P1_U3539) );
  INV_X1 U10935 ( .A(n9730), .ZN(n9731) );
  NAND2_X1 U10936 ( .A1(n9732), .A2(n9731), .ZN(n9799) );
  MUX2_X1 U10937 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9799), .S(n9910), .Z(n9733) );
  AOI21_X1 U10938 ( .B1(n9734), .B2(n9801), .A(n9733), .ZN(n9735) );
  OAI21_X1 U10939 ( .B1(n9804), .B2(n9736), .A(n9735), .ZN(P1_U3538) );
  AOI211_X1 U10940 ( .C1(n9745), .C2(n9739), .A(n9738), .B(n9737), .ZN(n9740)
         );
  OAI21_X1 U10941 ( .B1(n9741), .B2(n9747), .A(n9740), .ZN(n9805) );
  MUX2_X1 U10942 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n9805), .S(n9910), .Z(
        P1_U3537) );
  AOI211_X1 U10943 ( .C1(n9745), .C2(n9744), .A(n9743), .B(n9742), .ZN(n9746)
         );
  OAI21_X1 U10944 ( .B1(n9748), .B2(n9747), .A(n9746), .ZN(n9806) );
  MUX2_X1 U10945 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n9806), .S(n9910), .Z(
        P1_U3535) );
  INV_X1 U10946 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n9750) );
  MUX2_X1 U10947 ( .A(n9750), .B(n9749), .S(n9906), .Z(n9751) );
  OAI21_X1 U10948 ( .B1(n9752), .B2(n9755), .A(n9751), .ZN(P1_U3521) );
  INV_X1 U10949 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n10166) );
  MUX2_X1 U10950 ( .A(n10166), .B(n9753), .S(n9906), .Z(n9754) );
  OAI21_X1 U10951 ( .B1(n9756), .B2(n9755), .A(n9754), .ZN(P1_U3520) );
  MUX2_X1 U10952 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n9757), .S(n9906), .Z(
        P1_U3518) );
  MUX2_X1 U10953 ( .A(n9759), .B(n9758), .S(n9906), .Z(n9760) );
  OAI21_X1 U10954 ( .B1(n9761), .B2(n9803), .A(n9760), .ZN(P1_U3517) );
  MUX2_X1 U10955 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9762), .S(n9906), .Z(n9763) );
  AOI21_X1 U10956 ( .B1(n5657), .B2(n9764), .A(n9763), .ZN(n9765) );
  OAI21_X1 U10957 ( .B1(n9766), .B2(n9803), .A(n9765), .ZN(P1_U3516) );
  INV_X1 U10958 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n9768) );
  MUX2_X1 U10959 ( .A(n9768), .B(n9767), .S(n9906), .Z(n9769) );
  OAI21_X1 U10960 ( .B1(n9770), .B2(n9803), .A(n9769), .ZN(P1_U3515) );
  INV_X1 U10961 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n9771) );
  MUX2_X1 U10962 ( .A(n9772), .B(n9771), .S(n9905), .Z(n9773) );
  OAI21_X1 U10963 ( .B1(n9774), .B2(n9803), .A(n9773), .ZN(P1_U3514) );
  MUX2_X1 U10964 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9775), .S(n9906), .Z(
        P1_U3513) );
  MUX2_X1 U10965 ( .A(n9777), .B(n9776), .S(n9906), .Z(n9778) );
  OAI21_X1 U10966 ( .B1(n9779), .B2(n9803), .A(n9778), .ZN(P1_U3512) );
  INV_X1 U10967 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n9781) );
  MUX2_X1 U10968 ( .A(n9781), .B(n9780), .S(n9906), .Z(n9782) );
  OAI21_X1 U10969 ( .B1(n9783), .B2(n9803), .A(n9782), .ZN(P1_U3511) );
  MUX2_X1 U10970 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9784), .S(n9906), .Z(n9785) );
  AOI21_X1 U10971 ( .B1(n9787), .B2(n9786), .A(n9785), .ZN(n9788) );
  INV_X1 U10972 ( .A(n9788), .ZN(P1_U3510) );
  MUX2_X1 U10973 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9789), .S(n9906), .Z(
        P1_U3509) );
  MUX2_X1 U10974 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9790), .S(n9906), .Z(n9791) );
  AOI21_X1 U10975 ( .B1(n5657), .B2(n9792), .A(n9791), .ZN(n9793) );
  OAI21_X1 U10976 ( .B1(n9794), .B2(n9803), .A(n9793), .ZN(P1_U3507) );
  INV_X1 U10977 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n9796) );
  MUX2_X1 U10978 ( .A(n9796), .B(n9795), .S(n9906), .Z(n9797) );
  OAI21_X1 U10979 ( .B1(n9798), .B2(n9803), .A(n9797), .ZN(P1_U3504) );
  MUX2_X1 U10980 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n9799), .S(n9906), .Z(n9800) );
  AOI21_X1 U10981 ( .B1(n5657), .B2(n9801), .A(n9800), .ZN(n9802) );
  OAI21_X1 U10982 ( .B1(n9804), .B2(n9803), .A(n9802), .ZN(P1_U3501) );
  MUX2_X1 U10983 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n9805), .S(n9906), .Z(
        P1_U3498) );
  MUX2_X1 U10984 ( .A(P1_REG0_REG_13__SCAN_IN), .B(n9806), .S(n9906), .Z(
        P1_U3492) );
  INV_X1 U10985 ( .A(n9807), .ZN(n9808) );
  MUX2_X1 U10986 ( .A(P1_D_REG_1__SCAN_IN), .B(n9810), .S(n9891), .Z(P1_U3440)
         );
  MUX2_X1 U10987 ( .A(P1_D_REG_0__SCAN_IN), .B(n9811), .S(n9891), .Z(P1_U3439)
         );
  INV_X1 U10988 ( .A(n9812), .ZN(n9819) );
  NOR4_X1 U10989 ( .A1(n9813), .A2(P1_IR_REG_30__SCAN_IN), .A3(n9815), .A4(
        P1_U3086), .ZN(n9816) );
  AOI21_X1 U10990 ( .B1(n9817), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9816), .ZN(
        n9818) );
  OAI21_X1 U10991 ( .B1(n9819), .B2(n9822), .A(n9818), .ZN(P1_U3324) );
  OAI222_X1 U10992 ( .A1(n9824), .A2(n9823), .B1(n9822), .B2(n9821), .C1(n9820), .C2(P1_U3086), .ZN(P1_U3326) );
  MUX2_X1 U10993 ( .A(n9825), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  OAI21_X1 U10994 ( .B1(n9828), .B2(n9827), .A(n9826), .ZN(n9835) );
  AOI21_X1 U10995 ( .B1(n9831), .B2(n9830), .A(n9829), .ZN(n9833) );
  OAI22_X1 U10996 ( .A1(n9833), .A2(n9869), .B1(n9832), .B2(n9866), .ZN(n9834)
         );
  AOI21_X1 U10997 ( .B1(n9872), .B2(n9835), .A(n9834), .ZN(n9837) );
  OAI211_X1 U10998 ( .C1(n9875), .C2(n9838), .A(n9837), .B(n9836), .ZN(
        P1_U3252) );
  XNOR2_X1 U10999 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U11000 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  NOR3_X1 U11001 ( .A1(n9841), .A2(n9840), .A3(n4581), .ZN(n9842) );
  NOR3_X1 U11002 ( .A1(n9844), .A2(n9843), .A3(n9842), .ZN(n9854) );
  NOR2_X1 U11003 ( .A1(n9866), .A2(n9845), .ZN(n9853) );
  INV_X1 U11004 ( .A(n9846), .ZN(n9851) );
  NOR3_X1 U11005 ( .A1(n9849), .A2(n9848), .A3(n9847), .ZN(n9850) );
  NOR3_X1 U11006 ( .A1(n9869), .A2(n9851), .A3(n9850), .ZN(n9852) );
  NOR4_X1 U11007 ( .A1(n9855), .A2(n9854), .A3(n9853), .A4(n9852), .ZN(n9857)
         );
  OAI211_X1 U11008 ( .C1(n9858), .C2(n9875), .A(n9857), .B(n9856), .ZN(
        P1_U3247) );
  MUX2_X1 U11009 ( .A(P1_REG2_REG_17__SCAN_IN), .B(n4596), .S(n9859), .Z(n9862) );
  NAND2_X1 U11010 ( .A1(n9861), .A2(n9862), .ZN(n9860) );
  OAI21_X1 U11011 ( .B1(n9862), .B2(n9861), .A(n9860), .ZN(n9871) );
  AOI21_X1 U11012 ( .B1(n9865), .B2(n9864), .A(n9863), .ZN(n9868) );
  OAI22_X1 U11013 ( .A1(n9869), .A2(n9868), .B1(n9867), .B2(n9866), .ZN(n9870)
         );
  AOI21_X1 U11014 ( .B1(n9872), .B2(n9871), .A(n9870), .ZN(n9874) );
  OAI211_X1 U11015 ( .C1(n9875), .C2(n10181), .A(n9874), .B(n9873), .ZN(
        P1_U3260) );
  NAND3_X1 U11016 ( .A1(n9892), .A2(n9877), .A3(n9876), .ZN(n9885) );
  INV_X1 U11017 ( .A(n9877), .ZN(n9878) );
  NAND2_X1 U11018 ( .A1(n9879), .A2(n9878), .ZN(n9895) );
  INV_X1 U11019 ( .A(n9880), .ZN(n9882) );
  NAND2_X1 U11020 ( .A1(n9881), .A2(n6427), .ZN(n9894) );
  OAI21_X1 U11021 ( .B1(n9895), .B2(n9882), .A(n9894), .ZN(n9883) );
  INV_X1 U11022 ( .A(n9883), .ZN(n9884) );
  OAI211_X1 U11023 ( .C1(n7144), .C2(n9886), .A(n9885), .B(n9884), .ZN(n9887)
         );
  INV_X1 U11024 ( .A(n9887), .ZN(n9888) );
  AOI22_X1 U11025 ( .A1(n9889), .A2(n5137), .B1(n9888), .B2(n9560), .ZN(
        P1_U3293) );
  INV_X1 U11026 ( .A(P1_D_REG_31__SCAN_IN), .ZN(n10096) );
  NOR2_X1 U11027 ( .A1(n9891), .A2(n10096), .ZN(P1_U3294) );
  INV_X1 U11028 ( .A(P1_D_REG_30__SCAN_IN), .ZN(n10308) );
  NOR2_X1 U11029 ( .A1(n9891), .A2(n10308), .ZN(P1_U3295) );
  INV_X1 U11030 ( .A(P1_D_REG_29__SCAN_IN), .ZN(n10211) );
  NOR2_X1 U11031 ( .A1(n9891), .A2(n10211), .ZN(P1_U3296) );
  AND2_X1 U11032 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n9890), .ZN(P1_U3297) );
  AND2_X1 U11033 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n9890), .ZN(P1_U3298) );
  NOR2_X1 U11034 ( .A1(n9891), .A2(n10159), .ZN(P1_U3299) );
  AND2_X1 U11035 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n9890), .ZN(P1_U3300) );
  AND2_X1 U11036 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9890), .ZN(P1_U3301) );
  INV_X1 U11037 ( .A(P1_D_REG_23__SCAN_IN), .ZN(n10210) );
  NOR2_X1 U11038 ( .A1(n9891), .A2(n10210), .ZN(P1_U3302) );
  AND2_X1 U11039 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n9890), .ZN(P1_U3303) );
  AND2_X1 U11040 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n9890), .ZN(P1_U3304) );
  INV_X1 U11041 ( .A(P1_D_REG_20__SCAN_IN), .ZN(n10324) );
  NOR2_X1 U11042 ( .A1(n9891), .A2(n10324), .ZN(P1_U3305) );
  AND2_X1 U11043 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n9890), .ZN(P1_U3306) );
  NOR2_X1 U11044 ( .A1(n9891), .A2(n10237), .ZN(P1_U3307) );
  AND2_X1 U11045 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n9890), .ZN(P1_U3308) );
  AND2_X1 U11046 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n9890), .ZN(P1_U3309) );
  AND2_X1 U11047 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n9890), .ZN(P1_U3310) );
  INV_X1 U11048 ( .A(P1_D_REG_14__SCAN_IN), .ZN(n10247) );
  NOR2_X1 U11049 ( .A1(n9891), .A2(n10247), .ZN(P1_U3311) );
  AND2_X1 U11050 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n9890), .ZN(P1_U3312) );
  INV_X1 U11051 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n10184) );
  NOR2_X1 U11052 ( .A1(n9891), .A2(n10184), .ZN(P1_U3313) );
  AND2_X1 U11053 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n9890), .ZN(P1_U3314) );
  AND2_X1 U11054 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n9890), .ZN(P1_U3315) );
  AND2_X1 U11055 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n9890), .ZN(P1_U3316) );
  INV_X1 U11056 ( .A(P1_D_REG_8__SCAN_IN), .ZN(n10223) );
  NOR2_X1 U11057 ( .A1(n9891), .A2(n10223), .ZN(P1_U3317) );
  AND2_X1 U11058 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n9890), .ZN(P1_U3318) );
  AND2_X1 U11059 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n9890), .ZN(P1_U3319) );
  AND2_X1 U11060 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n9890), .ZN(P1_U3320) );
  NOR2_X1 U11061 ( .A1(n9891), .A2(n10238), .ZN(P1_U3321) );
  NOR2_X1 U11062 ( .A1(n9891), .A2(n10064), .ZN(P1_U3322) );
  INV_X1 U11063 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n10325) );
  NOR2_X1 U11064 ( .A1(n9891), .A2(n10325), .ZN(P1_U3323) );
  OAI21_X1 U11065 ( .B1(n9893), .B2(n9903), .A(n9892), .ZN(n9896) );
  AND3_X1 U11066 ( .A1(n9896), .A2(n9895), .A3(n9894), .ZN(n9907) );
  AOI22_X1 U11067 ( .A1(n9906), .A2(n9907), .B1(n5136), .B2(n9905), .ZN(
        P1_U3453) );
  INV_X1 U11068 ( .A(n9897), .ZN(n9898) );
  OAI21_X1 U11069 ( .B1(n9900), .B2(n9899), .A(n9898), .ZN(n9901) );
  AOI211_X1 U11070 ( .C1(n9904), .C2(n9903), .A(n9902), .B(n9901), .ZN(n9909)
         );
  INV_X1 U11071 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n10326) );
  AOI22_X1 U11072 ( .A1(n9906), .A2(n9909), .B1(n10326), .B2(n9905), .ZN(
        P1_U3468) );
  AOI22_X1 U11073 ( .A1(n9910), .A2(n9907), .B1(n6876), .B2(n9908), .ZN(
        P1_U3522) );
  AOI22_X1 U11074 ( .A1(n9910), .A2(n9909), .B1(n5196), .B2(n9908), .ZN(
        P1_U3527) );
  INV_X1 U11075 ( .A(n9911), .ZN(n9917) );
  AOI22_X1 U11076 ( .A1(P2_ADDR_REG_0__SCAN_IN), .A2(n9934), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3151), .ZN(n9916) );
  XNOR2_X1 U11077 ( .A(n9912), .B(n9911), .ZN(n9913) );
  OAI21_X1 U11078 ( .B1(n9914), .B2(n9918), .A(n9913), .ZN(n9915) );
  OAI211_X1 U11079 ( .C1(n9938), .C2(n9917), .A(n9916), .B(n9915), .ZN(
        P2_U3182) );
  OAI211_X1 U11080 ( .C1(n9921), .C2(n9920), .A(n9919), .B(n9918), .ZN(n9922)
         );
  INV_X1 U11081 ( .A(n9922), .ZN(n9933) );
  AOI21_X1 U11082 ( .B1(n9924), .B2(n9923), .A(n4518), .ZN(n9931) );
  AOI21_X1 U11083 ( .B1(n9927), .B2(n9926), .A(n9925), .ZN(n9928) );
  OAI22_X1 U11084 ( .A1(n9931), .A2(n9930), .B1(n9929), .B2(n9928), .ZN(n9932)
         );
  AOI211_X1 U11085 ( .C1(P2_ADDR_REG_4__SCAN_IN), .C2(n9934), .A(n9933), .B(
        n9932), .ZN(n9936) );
  OAI211_X1 U11086 ( .C1(n9938), .C2(n9937), .A(n9936), .B(n9935), .ZN(
        P2_U3186) );
  INV_X1 U11087 ( .A(n9939), .ZN(n9955) );
  OAI21_X1 U11088 ( .B1(n9941), .B2(n9946), .A(n9940), .ZN(n9969) );
  OAI22_X1 U11089 ( .A1(n9966), .A2(n9944), .B1(n9943), .B2(n9942), .ZN(n9954)
         );
  INV_X1 U11090 ( .A(n5739), .ZN(n9950) );
  NAND3_X1 U11091 ( .A1(n7534), .A2(n9946), .A3(n9945), .ZN(n9947) );
  AND2_X1 U11092 ( .A1(n7376), .A2(n9947), .ZN(n9948) );
  OAI222_X1 U11093 ( .A1(n9953), .A2(n9952), .B1(n9951), .B2(n9950), .C1(n9949), .C2(n9948), .ZN(n9967) );
  AOI211_X1 U11094 ( .C1(n9955), .C2(n9969), .A(n9954), .B(n9967), .ZN(n9959)
         );
  INV_X1 U11095 ( .A(n9956), .ZN(n9957) );
  AOI22_X1 U11096 ( .A1(n9969), .A2(n9957), .B1(n9960), .B2(
        P2_REG2_REG_2__SCAN_IN), .ZN(n9958) );
  OAI21_X1 U11097 ( .B1(n9960), .B2(n9959), .A(n9958), .ZN(P2_U3231) );
  INV_X1 U11098 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n9965) );
  NOR2_X1 U11099 ( .A1(n9961), .A2(n10005), .ZN(n9963) );
  AOI211_X1 U11100 ( .C1(n9970), .C2(n9964), .A(n9963), .B(n9962), .ZN(n10018)
         );
  AOI22_X1 U11101 ( .A1(n10017), .A2(n9965), .B1(n10018), .B2(n10016), .ZN(
        P2_U3393) );
  NOR2_X1 U11102 ( .A1(n9966), .A2(n10005), .ZN(n9968) );
  AOI211_X1 U11103 ( .C1(n9970), .C2(n9969), .A(n9968), .B(n9967), .ZN(n10019)
         );
  AOI22_X1 U11104 ( .A1(n10017), .A2(n5741), .B1(n10019), .B2(n10016), .ZN(
        P2_U3396) );
  INV_X1 U11105 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n9976) );
  INV_X1 U11106 ( .A(n9971), .ZN(n9975) );
  OAI22_X1 U11107 ( .A1(n9973), .A2(n10010), .B1(n9972), .B2(n10005), .ZN(
        n9974) );
  NOR2_X1 U11108 ( .A1(n9975), .A2(n9974), .ZN(n10020) );
  AOI22_X1 U11109 ( .A1(n10017), .A2(n9976), .B1(n10020), .B2(n10016), .ZN(
        P2_U3399) );
  INV_X1 U11110 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n9982) );
  INV_X1 U11111 ( .A(n9977), .ZN(n9981) );
  OAI22_X1 U11112 ( .A1(n9979), .A2(n10010), .B1(n9978), .B2(n10005), .ZN(
        n9980) );
  NOR2_X1 U11113 ( .A1(n9981), .A2(n9980), .ZN(n10021) );
  AOI22_X1 U11114 ( .A1(n10017), .A2(n9982), .B1(n10021), .B2(n10016), .ZN(
        P2_U3402) );
  INV_X1 U11115 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n9988) );
  INV_X1 U11116 ( .A(n9983), .ZN(n9987) );
  OAI22_X1 U11117 ( .A1(n9985), .A2(n10010), .B1(n9984), .B2(n10005), .ZN(
        n9986) );
  NOR2_X1 U11118 ( .A1(n9987), .A2(n9986), .ZN(n10022) );
  AOI22_X1 U11119 ( .A1(n10017), .A2(n9988), .B1(n10022), .B2(n10016), .ZN(
        P2_U3405) );
  INV_X1 U11120 ( .A(n9989), .ZN(n9993) );
  OAI22_X1 U11121 ( .A1(n9991), .A2(n10010), .B1(n9990), .B2(n10005), .ZN(
        n9992) );
  NOR2_X1 U11122 ( .A1(n9993), .A2(n9992), .ZN(n10023) );
  AOI22_X1 U11123 ( .A1(n10017), .A2(n5798), .B1(n10023), .B2(n10016), .ZN(
        P2_U3408) );
  OAI22_X1 U11124 ( .A1(n9995), .A2(n10010), .B1(n9994), .B2(n10005), .ZN(
        n9998) );
  INV_X1 U11125 ( .A(n9996), .ZN(n9997) );
  NOR2_X1 U11126 ( .A1(n9998), .A2(n9997), .ZN(n10024) );
  AOI22_X1 U11127 ( .A1(n10017), .A2(n5826), .B1(n10024), .B2(n10016), .ZN(
        P2_U3414) );
  INV_X1 U11128 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n10004) );
  OAI22_X1 U11129 ( .A1(n10001), .A2(n10000), .B1(n9999), .B2(n10005), .ZN(
        n10002) );
  NOR2_X1 U11130 ( .A1(n10003), .A2(n10002), .ZN(n10025) );
  AOI22_X1 U11131 ( .A1(n10017), .A2(n10004), .B1(n10025), .B2(n10016), .ZN(
        P2_U3420) );
  INV_X1 U11132 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n10327) );
  OAI22_X1 U11133 ( .A1(n10007), .A2(n10010), .B1(n10006), .B2(n10005), .ZN(
        n10008) );
  NOR2_X1 U11134 ( .A1(n10009), .A2(n10008), .ZN(n10026) );
  AOI22_X1 U11135 ( .A1(n10017), .A2(n10327), .B1(n10026), .B2(n10016), .ZN(
        P2_U3423) );
  INV_X1 U11136 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n10111) );
  NOR2_X1 U11137 ( .A1(n10011), .A2(n10010), .ZN(n10013) );
  AOI211_X1 U11138 ( .C1(n10015), .C2(n10014), .A(n10013), .B(n10012), .ZN(
        n10028) );
  AOI22_X1 U11139 ( .A1(n10017), .A2(n10111), .B1(n10028), .B2(n10016), .ZN(
        P2_U3426) );
  AOI22_X1 U11140 ( .A1(n10029), .A2(n10018), .B1(n6256), .B2(n10027), .ZN(
        P2_U3460) );
  AOI22_X1 U11141 ( .A1(n10029), .A2(n10019), .B1(n6214), .B2(n10027), .ZN(
        P2_U3461) );
  AOI22_X1 U11142 ( .A1(n10029), .A2(n10020), .B1(n5758), .B2(n10027), .ZN(
        P2_U3462) );
  AOI22_X1 U11143 ( .A1(n10029), .A2(n10021), .B1(n6217), .B2(n10027), .ZN(
        P2_U3463) );
  AOI22_X1 U11144 ( .A1(n10029), .A2(n10022), .B1(n5787), .B2(n10027), .ZN(
        P2_U3464) );
  AOI22_X1 U11145 ( .A1(n10029), .A2(n10023), .B1(n5801), .B2(n10027), .ZN(
        P2_U3465) );
  AOI22_X1 U11146 ( .A1(n10029), .A2(n10024), .B1(n6226), .B2(n10027), .ZN(
        P2_U3467) );
  AOI22_X1 U11147 ( .A1(n10029), .A2(n10025), .B1(n5855), .B2(n10027), .ZN(
        P2_U3469) );
  AOI22_X1 U11148 ( .A1(n10029), .A2(n10026), .B1(n5870), .B2(n10027), .ZN(
        P2_U3470) );
  AOI22_X1 U11149 ( .A1(n10029), .A2(n10028), .B1(n5889), .B2(n10027), .ZN(
        P2_U3471) );
  NOR2_X1 U11150 ( .A1(n10031), .A2(n10030), .ZN(n10032) );
  XOR2_X1 U11151 ( .A(n10032), .B(P2_ADDR_REG_1__SCAN_IN), .Z(ADD_1068_U5) );
  AOI21_X1 U11152 ( .B1(n6968), .B2(n10034), .A(n10033), .ZN(ADD_1068_U46) );
  OAI21_X1 U11153 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n10036), .A(n10035), 
        .ZN(n10037) );
  XOR2_X1 U11154 ( .A(n10037), .B(n10099), .Z(ADD_1068_U55) );
  XNOR2_X1 U11155 ( .A(n10039), .B(n10038), .ZN(ADD_1068_U56) );
  XNOR2_X1 U11156 ( .A(n10041), .B(n10040), .ZN(ADD_1068_U57) );
  XNOR2_X1 U11157 ( .A(n10043), .B(n10042), .ZN(ADD_1068_U58) );
  XNOR2_X1 U11158 ( .A(n10045), .B(n10044), .ZN(ADD_1068_U59) );
  XNOR2_X1 U11159 ( .A(n10047), .B(n10046), .ZN(ADD_1068_U60) );
  XNOR2_X1 U11160 ( .A(n10049), .B(n10048), .ZN(ADD_1068_U61) );
  XNOR2_X1 U11161 ( .A(n10051), .B(n10050), .ZN(ADD_1068_U62) );
  XNOR2_X1 U11162 ( .A(n10053), .B(n10052), .ZN(ADD_1068_U63) );
  MUX2_X1 U11163 ( .A(n10056), .B(n10055), .S(n10054), .Z(n10269) );
  AOI22_X1 U11164 ( .A1(n10339), .A2(keyinput61), .B1(n10058), .B2(keyinput98), 
        .ZN(n10057) );
  OAI221_X1 U11165 ( .B1(n10339), .B2(keyinput61), .C1(n10058), .C2(keyinput98), .A(n10057), .ZN(n10069) );
  AOI22_X1 U11166 ( .A1(n8770), .A2(keyinput119), .B1(n10060), .B2(keyinput85), 
        .ZN(n10059) );
  OAI221_X1 U11167 ( .B1(n8770), .B2(keyinput119), .C1(n10060), .C2(keyinput85), .A(n10059), .ZN(n10068) );
  AOI22_X1 U11168 ( .A1(n10062), .A2(keyinput62), .B1(n10344), .B2(keyinput67), 
        .ZN(n10061) );
  OAI221_X1 U11169 ( .B1(n10062), .B2(keyinput62), .C1(n10344), .C2(keyinput67), .A(n10061), .ZN(n10067) );
  AOI22_X1 U11170 ( .A1(n10065), .A2(keyinput69), .B1(n10064), .B2(keyinput80), 
        .ZN(n10063) );
  OAI221_X1 U11171 ( .B1(n10065), .B2(keyinput69), .C1(n10064), .C2(keyinput80), .A(n10063), .ZN(n10066) );
  NOR4_X1 U11172 ( .A1(n10069), .A2(n10068), .A3(n10067), .A4(n10066), .ZN(
        n10109) );
  AOI22_X1 U11173 ( .A1(n10071), .A2(keyinput72), .B1(n10343), .B2(keyinput127), .ZN(n10070) );
  OAI221_X1 U11174 ( .B1(n10071), .B2(keyinput72), .C1(n10343), .C2(
        keyinput127), .A(n10070), .ZN(n10080) );
  INV_X1 U11175 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n10073) );
  AOI22_X1 U11176 ( .A1(n10073), .A2(keyinput109), .B1(keyinput106), .B2(
        n10342), .ZN(n10072) );
  OAI221_X1 U11177 ( .B1(n10073), .B2(keyinput109), .C1(n10342), .C2(
        keyinput106), .A(n10072), .ZN(n10079) );
  AOI22_X1 U11178 ( .A1(n5826), .A2(keyinput92), .B1(n7905), .B2(keyinput121), 
        .ZN(n10074) );
  OAI221_X1 U11179 ( .B1(n5826), .B2(keyinput92), .C1(n7905), .C2(keyinput121), 
        .A(n10074), .ZN(n10078) );
  AOI22_X1 U11180 ( .A1(n6998), .A2(keyinput91), .B1(n10076), .B2(keyinput15), 
        .ZN(n10075) );
  OAI221_X1 U11181 ( .B1(n6998), .B2(keyinput91), .C1(n10076), .C2(keyinput15), 
        .A(n10075), .ZN(n10077) );
  NOR4_X1 U11182 ( .A1(n10080), .A2(n10079), .A3(n10078), .A4(n10077), .ZN(
        n10108) );
  AOI22_X1 U11183 ( .A1(n8209), .A2(keyinput102), .B1(n10082), .B2(keyinput20), 
        .ZN(n10081) );
  OAI221_X1 U11184 ( .B1(n8209), .B2(keyinput102), .C1(n10082), .C2(keyinput20), .A(n10081), .ZN(n10091) );
  AOI22_X1 U11185 ( .A1(n10333), .A2(keyinput105), .B1(n7567), .B2(keyinput24), 
        .ZN(n10083) );
  OAI221_X1 U11186 ( .B1(n10333), .B2(keyinput105), .C1(n7567), .C2(keyinput24), .A(n10083), .ZN(n10090) );
  INV_X1 U11187 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n10332) );
  AOI22_X1 U11188 ( .A1(n10332), .A2(keyinput5), .B1(n10340), .B2(keyinput82), 
        .ZN(n10084) );
  OAI221_X1 U11189 ( .B1(n10332), .B2(keyinput5), .C1(n10340), .C2(keyinput82), 
        .A(n10084), .ZN(n10089) );
  AOI22_X1 U11190 ( .A1(n10087), .A2(keyinput84), .B1(keyinput46), .B2(n10086), 
        .ZN(n10085) );
  OAI221_X1 U11191 ( .B1(n10087), .B2(keyinput84), .C1(n10086), .C2(keyinput46), .A(n10085), .ZN(n10088) );
  NOR4_X1 U11192 ( .A1(n10091), .A2(n10090), .A3(n10089), .A4(n10088), .ZN(
        n10107) );
  INV_X1 U11193 ( .A(SI_19_), .ZN(n10094) );
  AOI22_X1 U11194 ( .A1(n10094), .A2(keyinput22), .B1(n10093), .B2(keyinput66), 
        .ZN(n10092) );
  OAI221_X1 U11195 ( .B1(n10094), .B2(keyinput22), .C1(n10093), .C2(keyinput66), .A(n10092), .ZN(n10105) );
  AOI22_X1 U11196 ( .A1(n10334), .A2(keyinput90), .B1(n10096), .B2(keyinput71), 
        .ZN(n10095) );
  OAI221_X1 U11197 ( .B1(n10334), .B2(keyinput90), .C1(n10096), .C2(keyinput71), .A(n10095), .ZN(n10104) );
  AOI22_X1 U11198 ( .A1(n10099), .A2(keyinput81), .B1(n10098), .B2(keyinput2), 
        .ZN(n10097) );
  OAI221_X1 U11199 ( .B1(n10099), .B2(keyinput81), .C1(n10098), .C2(keyinput2), 
        .A(n10097), .ZN(n10103) );
  XNOR2_X1 U11200 ( .A(P1_REG3_REG_13__SCAN_IN), .B(keyinput33), .ZN(n10101)
         );
  XNOR2_X1 U11201 ( .A(P1_IR_REG_17__SCAN_IN), .B(keyinput10), .ZN(n10100) );
  NAND2_X1 U11202 ( .A1(n10101), .A2(n10100), .ZN(n10102) );
  NOR4_X1 U11203 ( .A1(n10105), .A2(n10104), .A3(n10103), .A4(n10102), .ZN(
        n10106) );
  NAND4_X1 U11204 ( .A1(n10109), .A2(n10108), .A3(n10107), .A4(n10106), .ZN(
        n10267) );
  AOI22_X1 U11205 ( .A1(n10308), .A2(keyinput3), .B1(keyinput56), .B2(n10312), 
        .ZN(n10110) );
  OAI221_X1 U11206 ( .B1(n10308), .B2(keyinput3), .C1(n10312), .C2(keyinput56), 
        .A(n10110), .ZN(n10119) );
  XOR2_X1 U11207 ( .A(P2_IR_REG_26__SCAN_IN), .B(keyinput19), .Z(n10118) );
  XNOR2_X1 U11208 ( .A(keyinput36), .B(n10111), .ZN(n10117) );
  XNOR2_X1 U11209 ( .A(P1_IR_REG_18__SCAN_IN), .B(keyinput54), .ZN(n10115) );
  XNOR2_X1 U11210 ( .A(SI_12_), .B(keyinput93), .ZN(n10114) );
  XNOR2_X1 U11211 ( .A(P2_IR_REG_11__SCAN_IN), .B(keyinput108), .ZN(n10113) );
  XNOR2_X1 U11212 ( .A(P1_IR_REG_20__SCAN_IN), .B(keyinput116), .ZN(n10112) );
  NAND4_X1 U11213 ( .A1(n10115), .A2(n10114), .A3(n10113), .A4(n10112), .ZN(
        n10116) );
  NOR4_X1 U11214 ( .A1(n10119), .A2(n10118), .A3(n10117), .A4(n10116), .ZN(
        n10157) );
  AOI22_X1 U11215 ( .A1(n10271), .A2(keyinput77), .B1(n10121), .B2(keyinput11), 
        .ZN(n10120) );
  OAI221_X1 U11216 ( .B1(n10271), .B2(keyinput77), .C1(n10121), .C2(keyinput11), .A(n10120), .ZN(n10130) );
  XNOR2_X1 U11217 ( .A(P2_REG1_REG_16__SCAN_IN), .B(keyinput23), .ZN(n10125)
         );
  XNOR2_X1 U11218 ( .A(SI_5_), .B(keyinput94), .ZN(n10124) );
  XNOR2_X1 U11219 ( .A(P1_IR_REG_26__SCAN_IN), .B(keyinput126), .ZN(n10123) );
  XNOR2_X1 U11220 ( .A(P2_IR_REG_19__SCAN_IN), .B(keyinput50), .ZN(n10122) );
  NAND4_X1 U11221 ( .A1(n10125), .A2(n10124), .A3(n10123), .A4(n10122), .ZN(
        n10129) );
  XNOR2_X1 U11222 ( .A(n10314), .B(keyinput124), .ZN(n10128) );
  XNOR2_X1 U11223 ( .A(keyinput6), .B(n10126), .ZN(n10127) );
  NOR4_X1 U11224 ( .A1(n10130), .A2(n10129), .A3(n10128), .A4(n10127), .ZN(
        n10156) );
  AOI22_X1 U11225 ( .A1(n10133), .A2(keyinput73), .B1(n10132), .B2(keyinput26), 
        .ZN(n10131) );
  OAI221_X1 U11226 ( .B1(n10133), .B2(keyinput73), .C1(n10132), .C2(keyinput26), .A(n10131), .ZN(n10141) );
  INV_X1 U11227 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n10282) );
  AOI22_X1 U11228 ( .A1(n10282), .A2(keyinput123), .B1(n10277), .B2(keyinput13), .ZN(n10134) );
  OAI221_X1 U11229 ( .B1(n10282), .B2(keyinput123), .C1(n10277), .C2(
        keyinput13), .A(n10134), .ZN(n10140) );
  AOI22_X1 U11230 ( .A1(n10280), .A2(keyinput53), .B1(n10281), .B2(keyinput97), 
        .ZN(n10135) );
  OAI221_X1 U11231 ( .B1(n10280), .B2(keyinput53), .C1(n10281), .C2(keyinput97), .A(n10135), .ZN(n10139) );
  XNOR2_X1 U11232 ( .A(P2_IR_REG_8__SCAN_IN), .B(keyinput12), .ZN(n10137) );
  XNOR2_X1 U11233 ( .A(P1_REG3_REG_16__SCAN_IN), .B(keyinput115), .ZN(n10136)
         );
  NAND2_X1 U11234 ( .A1(n10137), .A2(n10136), .ZN(n10138) );
  NOR4_X1 U11235 ( .A1(n10141), .A2(n10140), .A3(n10139), .A4(n10138), .ZN(
        n10155) );
  AOI22_X1 U11236 ( .A1(n10143), .A2(keyinput48), .B1(keyinput1), .B2(n10317), 
        .ZN(n10142) );
  OAI221_X1 U11237 ( .B1(n10143), .B2(keyinput48), .C1(n10317), .C2(keyinput1), 
        .A(n10142), .ZN(n10153) );
  AOI22_X1 U11238 ( .A1(n7405), .A2(keyinput63), .B1(n10145), .B2(keyinput42), 
        .ZN(n10144) );
  OAI221_X1 U11239 ( .B1(n7405), .B2(keyinput63), .C1(n10145), .C2(keyinput42), 
        .A(n10144), .ZN(n10152) );
  AOI22_X1 U11240 ( .A1(n6968), .A2(keyinput74), .B1(n10147), .B2(keyinput14), 
        .ZN(n10146) );
  OAI221_X1 U11241 ( .B1(n6968), .B2(keyinput74), .C1(n10147), .C2(keyinput14), 
        .A(n10146), .ZN(n10151) );
  XNOR2_X1 U11242 ( .A(P2_REG1_REG_18__SCAN_IN), .B(keyinput60), .ZN(n10149)
         );
  XNOR2_X1 U11243 ( .A(P2_IR_REG_2__SCAN_IN), .B(keyinput32), .ZN(n10148) );
  NAND2_X1 U11244 ( .A1(n10149), .A2(n10148), .ZN(n10150) );
  NOR4_X1 U11245 ( .A1(n10153), .A2(n10152), .A3(n10151), .A4(n10150), .ZN(
        n10154) );
  NAND4_X1 U11246 ( .A1(n10157), .A2(n10156), .A3(n10155), .A4(n10154), .ZN(
        n10266) );
  AOI22_X1 U11247 ( .A1(n7290), .A2(keyinput0), .B1(n10324), .B2(keyinput107), 
        .ZN(n10158) );
  OAI221_X1 U11248 ( .B1(n7290), .B2(keyinput0), .C1(n10324), .C2(keyinput107), 
        .A(n10158), .ZN(n10162) );
  XNOR2_X1 U11249 ( .A(n4695), .B(keyinput16), .ZN(n10161) );
  XNOR2_X1 U11250 ( .A(n10159), .B(keyinput7), .ZN(n10160) );
  OR3_X1 U11251 ( .A1(n10162), .A2(n10161), .A3(n10160), .ZN(n10169) );
  AOI22_X1 U11252 ( .A1(n10164), .A2(keyinput104), .B1(keyinput110), .B2(
        n10327), .ZN(n10163) );
  OAI221_X1 U11253 ( .B1(n10164), .B2(keyinput104), .C1(n10327), .C2(
        keyinput110), .A(n10163), .ZN(n10168) );
  AOI22_X1 U11254 ( .A1(n10166), .A2(keyinput76), .B1(n6339), .B2(keyinput49), 
        .ZN(n10165) );
  OAI221_X1 U11255 ( .B1(n10166), .B2(keyinput76), .C1(n6339), .C2(keyinput49), 
        .A(n10165), .ZN(n10167) );
  NOR3_X1 U11256 ( .A1(n10169), .A2(n10168), .A3(n10167), .ZN(n10207) );
  AOI22_X1 U11257 ( .A1(n10325), .A2(keyinput118), .B1(keyinput86), .B2(n7004), 
        .ZN(n10170) );
  OAI221_X1 U11258 ( .B1(n10325), .B2(keyinput118), .C1(n7004), .C2(keyinput86), .A(n10170), .ZN(n10179) );
  AOI22_X1 U11259 ( .A1(n5836), .A2(keyinput44), .B1(n5889), .B2(keyinput125), 
        .ZN(n10171) );
  OAI221_X1 U11260 ( .B1(n5836), .B2(keyinput44), .C1(n5889), .C2(keyinput125), 
        .A(n10171), .ZN(n10178) );
  AOI22_X1 U11261 ( .A1(n10173), .A2(keyinput40), .B1(keyinput9), .B2(n9552), 
        .ZN(n10172) );
  OAI221_X1 U11262 ( .B1(n10173), .B2(keyinput40), .C1(n9552), .C2(keyinput9), 
        .A(n10172), .ZN(n10177) );
  XOR2_X1 U11263 ( .A(n10326), .B(keyinput114), .Z(n10175) );
  XNOR2_X1 U11264 ( .A(P1_IR_REG_12__SCAN_IN), .B(keyinput4), .ZN(n10174) );
  NAND2_X1 U11265 ( .A1(n10175), .A2(n10174), .ZN(n10176) );
  NOR4_X1 U11266 ( .A1(n10179), .A2(n10178), .A3(n10177), .A4(n10176), .ZN(
        n10206) );
  AOI22_X1 U11267 ( .A1(n10302), .A2(keyinput88), .B1(keyinput35), .B2(n10181), 
        .ZN(n10180) );
  OAI221_X1 U11268 ( .B1(n10302), .B2(keyinput88), .C1(n10181), .C2(keyinput35), .A(n10180), .ZN(n10190) );
  INV_X1 U11269 ( .A(SI_6_), .ZN(n10299) );
  AOI22_X1 U11270 ( .A1(n7350), .A2(keyinput29), .B1(n10299), .B2(keyinput18), 
        .ZN(n10182) );
  OAI221_X1 U11271 ( .B1(n7350), .B2(keyinput29), .C1(n10299), .C2(keyinput18), 
        .A(n10182), .ZN(n10189) );
  AOI22_X1 U11272 ( .A1(n10184), .A2(keyinput39), .B1(n10301), .B2(keyinput79), 
        .ZN(n10183) );
  OAI221_X1 U11273 ( .B1(n10184), .B2(keyinput39), .C1(n10301), .C2(keyinput79), .A(n10183), .ZN(n10188) );
  XOR2_X1 U11274 ( .A(n6040), .B(keyinput122), .Z(n10186) );
  XNOR2_X1 U11275 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(keyinput78), .ZN(n10185)
         );
  NAND2_X1 U11276 ( .A1(n10186), .A2(n10185), .ZN(n10187) );
  NOR4_X1 U11277 ( .A1(n10190), .A2(n10189), .A3(n10188), .A4(n10187), .ZN(
        n10205) );
  AOI22_X1 U11278 ( .A1(n5461), .A2(keyinput52), .B1(n10192), .B2(keyinput95), 
        .ZN(n10191) );
  OAI221_X1 U11279 ( .B1(n5461), .B2(keyinput52), .C1(n10192), .C2(keyinput95), 
        .A(n10191), .ZN(n10198) );
  INV_X1 U11280 ( .A(SI_30_), .ZN(n10194) );
  AOI22_X1 U11281 ( .A1(n10195), .A2(keyinput89), .B1(keyinput64), .B2(n10194), 
        .ZN(n10193) );
  OAI221_X1 U11282 ( .B1(n10195), .B2(keyinput89), .C1(n10194), .C2(keyinput64), .A(n10193), .ZN(n10197) );
  INV_X1 U11283 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n10311) );
  XNOR2_X1 U11284 ( .A(n10311), .B(keyinput87), .ZN(n10196) );
  OR3_X1 U11285 ( .A1(n10198), .A2(n10197), .A3(n10196), .ZN(n10203) );
  AOI22_X1 U11286 ( .A1(n10300), .A2(keyinput37), .B1(keyinput47), .B2(n7386), 
        .ZN(n10199) );
  OAI221_X1 U11287 ( .B1(n10300), .B2(keyinput37), .C1(n7386), .C2(keyinput47), 
        .A(n10199), .ZN(n10202) );
  XNOR2_X1 U11288 ( .A(n10200), .B(keyinput38), .ZN(n10201) );
  NOR3_X1 U11289 ( .A1(n10203), .A2(n10202), .A3(n10201), .ZN(n10204) );
  NAND4_X1 U11290 ( .A1(n10207), .A2(n10206), .A3(n10205), .A4(n10204), .ZN(
        n10265) );
  AOI22_X1 U11291 ( .A1(n10210), .A2(keyinput27), .B1(keyinput100), .B2(n10209), .ZN(n10208) );
  OAI221_X1 U11292 ( .B1(n10210), .B2(keyinput27), .C1(n10209), .C2(
        keyinput100), .A(n10208), .ZN(n10214) );
  XNOR2_X1 U11293 ( .A(n10211), .B(keyinput65), .ZN(n10213) );
  XOR2_X1 U11294 ( .A(P1_IR_REG_6__SCAN_IN), .B(keyinput117), .Z(n10212) );
  OR3_X1 U11295 ( .A1(n10214), .A2(n10213), .A3(n10212), .ZN(n10220) );
  AOI22_X1 U11296 ( .A1(n9449), .A2(keyinput99), .B1(n5304), .B2(keyinput68), 
        .ZN(n10215) );
  OAI221_X1 U11297 ( .B1(n9449), .B2(keyinput99), .C1(n5304), .C2(keyinput68), 
        .A(n10215), .ZN(n10219) );
  INV_X1 U11298 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n10217) );
  AOI22_X1 U11299 ( .A1(n6226), .A2(keyinput45), .B1(keyinput21), .B2(n10217), 
        .ZN(n10216) );
  OAI221_X1 U11300 ( .B1(n6226), .B2(keyinput45), .C1(n10217), .C2(keyinput21), 
        .A(n10216), .ZN(n10218) );
  NOR3_X1 U11301 ( .A1(n10220), .A2(n10219), .A3(n10218), .ZN(n10263) );
  XOR2_X1 U11302 ( .A(P1_REG1_REG_16__SCAN_IN), .B(keyinput58), .Z(n10227) );
  XNOR2_X1 U11303 ( .A(P1_IR_REG_2__SCAN_IN), .B(keyinput113), .ZN(n10222) );
  XNOR2_X1 U11304 ( .A(P1_IR_REG_28__SCAN_IN), .B(keyinput83), .ZN(n10221) );
  NAND2_X1 U11305 ( .A1(n10222), .A2(n10221), .ZN(n10226) );
  XNOR2_X1 U11306 ( .A(n10272), .B(keyinput103), .ZN(n10225) );
  XNOR2_X1 U11307 ( .A(keyinput111), .B(n10223), .ZN(n10224) );
  OR4_X1 U11308 ( .A1(n10227), .A2(n10226), .A3(n10225), .A4(n10224), .ZN(
        n10233) );
  AOI22_X1 U11309 ( .A1(n5985), .A2(keyinput8), .B1(n10229), .B2(keyinput41), 
        .ZN(n10228) );
  OAI221_X1 U11310 ( .B1(n5985), .B2(keyinput8), .C1(n10229), .C2(keyinput41), 
        .A(n10228), .ZN(n10232) );
  INV_X1 U11311 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n10230) );
  XNOR2_X1 U11312 ( .A(n10230), .B(keyinput34), .ZN(n10231) );
  NOR3_X1 U11313 ( .A1(n10233), .A2(n10232), .A3(n10231), .ZN(n10262) );
  AOI22_X1 U11314 ( .A1(n10297), .A2(keyinput70), .B1(n10235), .B2(keyinput112), .ZN(n10234) );
  OAI221_X1 U11315 ( .B1(n10297), .B2(keyinput70), .C1(n10235), .C2(
        keyinput112), .A(n10234), .ZN(n10245) );
  AOI22_X1 U11316 ( .A1(n10238), .A2(keyinput120), .B1(keyinput17), .B2(n10237), .ZN(n10236) );
  OAI221_X1 U11317 ( .B1(n10238), .B2(keyinput120), .C1(n10237), .C2(
        keyinput17), .A(n10236), .ZN(n10244) );
  AOI22_X1 U11318 ( .A1(n6345), .A2(keyinput96), .B1(n10298), .B2(keyinput57), 
        .ZN(n10239) );
  OAI221_X1 U11319 ( .B1(n6345), .B2(keyinput96), .C1(n10298), .C2(keyinput57), 
        .A(n10239), .ZN(n10243) );
  INV_X1 U11320 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n10241) );
  AOI22_X1 U11321 ( .A1(n10241), .A2(keyinput28), .B1(keyinput43), .B2(n10285), 
        .ZN(n10240) );
  OAI221_X1 U11322 ( .B1(n10241), .B2(keyinput28), .C1(n10285), .C2(keyinput43), .A(n10240), .ZN(n10242) );
  NOR4_X1 U11323 ( .A1(n10245), .A2(n10244), .A3(n10243), .A4(n10242), .ZN(
        n10261) );
  AOI22_X1 U11324 ( .A1(n10248), .A2(keyinput75), .B1(keyinput31), .B2(n10247), 
        .ZN(n10246) );
  OAI221_X1 U11325 ( .B1(n10248), .B2(keyinput75), .C1(n10247), .C2(keyinput31), .A(n10246), .ZN(n10259) );
  INV_X1 U11326 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n10250) );
  AOI22_X1 U11327 ( .A1(n10251), .A2(keyinput59), .B1(keyinput51), .B2(n10250), 
        .ZN(n10249) );
  OAI221_X1 U11328 ( .B1(n10251), .B2(keyinput59), .C1(n10250), .C2(keyinput51), .A(n10249), .ZN(n10258) );
  AOI22_X1 U11329 ( .A1(n10253), .A2(keyinput30), .B1(keyinput55), .B2(n10284), 
        .ZN(n10252) );
  OAI221_X1 U11330 ( .B1(n10253), .B2(keyinput30), .C1(n10284), .C2(keyinput55), .A(n10252), .ZN(n10257) );
  XNOR2_X1 U11331 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(keyinput25), .ZN(n10255)
         );
  XNOR2_X1 U11332 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(keyinput101), .ZN(n10254)
         );
  NAND2_X1 U11333 ( .A1(n10255), .A2(n10254), .ZN(n10256) );
  NOR4_X1 U11334 ( .A1(n10259), .A2(n10258), .A3(n10257), .A4(n10256), .ZN(
        n10260) );
  NAND4_X1 U11335 ( .A1(n10263), .A2(n10262), .A3(n10261), .A4(n10260), .ZN(
        n10264) );
  NOR4_X1 U11336 ( .A1(n10267), .A2(n10266), .A3(n10265), .A4(n10264), .ZN(
        n10268) );
  XNOR2_X1 U11337 ( .A(n10269), .B(n10268), .ZN(n10356) );
  AND4_X1 U11338 ( .A1(n10271), .A2(n10270), .A3(P1_IR_REG_17__SCAN_IN), .A4(
        P1_IR_REG_20__SCAN_IN), .ZN(n10274) );
  NOR2_X1 U11339 ( .A1(P1_REG0_REG_18__SCAN_IN), .A2(P1_REG1_REG_16__SCAN_IN), 
        .ZN(n10273) );
  NAND4_X1 U11340 ( .A1(n10274), .A2(SI_5_), .A3(n10273), .A4(n10272), .ZN(
        n10295) );
  NAND4_X1 U11341 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_1__SCAN_IN), .A3(
        n6226), .A4(n9449), .ZN(n10294) );
  NOR4_X1 U11342 ( .A1(n10275), .A2(n5015), .A3(P1_IR_REG_6__SCAN_IN), .A4(
        P1_IR_REG_18__SCAN_IN), .ZN(n10292) );
  NOR4_X1 U11343 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .A3(
        n10277), .A4(n10276), .ZN(n10279) );
  NAND3_X1 U11344 ( .A1(n5985), .A2(n10279), .A3(n10278), .ZN(n10289) );
  NOR4_X1 U11345 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(n10282), .A3(n10281), .A4(
        n10280), .ZN(n10283) );
  NAND2_X1 U11346 ( .A1(n7386), .A2(n10283), .ZN(n10288) );
  NAND4_X1 U11347 ( .A1(P2_REG3_REG_26__SCAN_IN), .A2(P2_IR_REG_23__SCAN_IN), 
        .A3(n10285), .A4(n10284), .ZN(n10286) );
  NOR4_X1 U11348 ( .A1(n10289), .A2(n10288), .A3(n10287), .A4(n10286), .ZN(
        n10291) );
  NAND4_X1 U11349 ( .A1(n10292), .A2(SI_30_), .A3(n10291), .A4(n10290), .ZN(
        n10293) );
  OR4_X1 U11350 ( .A1(n10296), .A2(n10295), .A3(n10294), .A4(n10293), .ZN(
        n10310) );
  NAND4_X1 U11351 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n6345), .A3(n10298), 
        .A4(n10297), .ZN(n10309) );
  NAND4_X1 U11352 ( .A1(n10301), .A2(n10300), .A3(n10299), .A4(n5461), .ZN(
        n10306) );
  NAND4_X1 U11353 ( .A1(P2_DATAO_REG_2__SCAN_IN), .A2(P2_REG2_REG_24__SCAN_IN), 
        .A3(P1_ADDR_REG_17__SCAN_IN), .A4(n10302), .ZN(n10305) );
  NAND4_X1 U11354 ( .A1(n10303), .A2(P2_REG1_REG_16__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P2_D_REG_15__SCAN_IN), .ZN(n10304) );
  OR3_X1 U11355 ( .A1(n10306), .A2(n10305), .A3(n10304), .ZN(n10307) );
  NOR4_X1 U11356 ( .A1(n10310), .A2(n10309), .A3(n10308), .A4(n10307), .ZN(
        n10323) );
  NAND4_X1 U11357 ( .A1(n10312), .A2(n10311), .A3(P1_IR_REG_12__SCAN_IN), .A4(
        P1_REG2_REG_15__SCAN_IN), .ZN(n10316) );
  INV_X1 U11358 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n10313) );
  NAND4_X1 U11359 ( .A1(n10314), .A2(n10313), .A3(P2_IR_REG_19__SCAN_IN), .A4(
        P2_REG1_REG_20__SCAN_IN), .ZN(n10315) );
  NOR3_X1 U11360 ( .A1(n10317), .A2(n10316), .A3(n10315), .ZN(n10321) );
  AND4_X1 U11361 ( .A1(n10319), .A2(P2_ADDR_REG_6__SCAN_IN), .A3(n10318), .A4(
        P1_ADDR_REG_0__SCAN_IN), .ZN(n10320) );
  NAND4_X1 U11362 ( .A1(n10323), .A2(n10322), .A3(n10321), .A4(n10320), .ZN(
        n10352) );
  NOR4_X1 U11363 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(P1_REG0_REG_30__SCAN_IN), 
        .A3(n6339), .A4(n10324), .ZN(n10331) );
  NOR4_X1 U11364 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(P1_REG2_REG_16__SCAN_IN), 
        .A3(P1_REG2_REG_12__SCAN_IN), .A4(P1_REG2_REG_3__SCAN_IN), .ZN(n10330)
         );
  NOR4_X1 U11365 ( .A1(P2_REG1_REG_12__SCAN_IN), .A2(P1_REG2_REG_20__SCAN_IN), 
        .A3(P1_REG1_REG_9__SCAN_IN), .A4(n10325), .ZN(n10329) );
  NOR4_X1 U11366 ( .A1(P1_DATAO_REG_1__SCAN_IN), .A2(P2_REG2_REG_9__SCAN_IN), 
        .A3(n10327), .A4(n10326), .ZN(n10328) );
  NAND4_X1 U11367 ( .A1(n10331), .A2(n10330), .A3(n10329), .A4(n10328), .ZN(
        n10351) );
  NOR4_X1 U11368 ( .A1(P2_REG3_REG_21__SCAN_IN), .A2(n7567), .A3(n10333), .A4(
        n10332), .ZN(n10338) );
  NOR4_X1 U11369 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P1_REG0_REG_15__SCAN_IN), 
        .A3(P1_REG1_REG_6__SCAN_IN), .A4(P2_REG1_REG_31__SCAN_IN), .ZN(n10337)
         );
  NOR4_X1 U11370 ( .A1(P2_IR_REG_26__SCAN_IN), .A2(SI_19_), .A3(SI_12_), .A4(
        P2_REG0_REG_12__SCAN_IN), .ZN(n10336) );
  NOR4_X1 U11371 ( .A1(P2_REG0_REG_17__SCAN_IN), .A2(P1_REG3_REG_24__SCAN_IN), 
        .A3(P2_ADDR_REG_18__SCAN_IN), .A4(n10334), .ZN(n10335) );
  NAND4_X1 U11372 ( .A1(n10338), .A2(n10337), .A3(n10336), .A4(n10335), .ZN(
        n10350) );
  NOR4_X1 U11373 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(P1_REG3_REG_16__SCAN_IN), 
        .A3(n10340), .A4(n10339), .ZN(n10348) );
  NOR4_X1 U11374 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_REG3_REG_10__SCAN_IN), 
        .A3(n5304), .A4(n10341), .ZN(n10347) );
  NOR4_X1 U11375 ( .A1(P2_REG0_REG_8__SCAN_IN), .A2(n7905), .A3(n10343), .A4(
        n10342), .ZN(n10346) );
  NOR4_X1 U11376 ( .A1(P2_REG2_REG_26__SCAN_IN), .A2(SI_8_), .A3(
        P1_REG3_REG_25__SCAN_IN), .A4(n10344), .ZN(n10345) );
  NAND4_X1 U11377 ( .A1(n10348), .A2(n10347), .A3(n10346), .A4(n10345), .ZN(
        n10349) );
  NOR4_X1 U11378 ( .A1(n10352), .A2(n10351), .A3(n10350), .A4(n10349), .ZN(
        n10354) );
  NAND2_X1 U11379 ( .A1(n10354), .A2(n10353), .ZN(n10355) );
  XNOR2_X1 U11380 ( .A(n10356), .B(n10355), .ZN(P1_U3572) );
  XNOR2_X1 U11381 ( .A(n10358), .B(n10357), .ZN(ADD_1068_U50) );
  XNOR2_X1 U11382 ( .A(n10360), .B(n10359), .ZN(ADD_1068_U51) );
  XNOR2_X1 U11383 ( .A(n10362), .B(n10361), .ZN(ADD_1068_U47) );
  XNOR2_X1 U11384 ( .A(n10364), .B(n10363), .ZN(ADD_1068_U49) );
  XNOR2_X1 U11385 ( .A(n10366), .B(n10365), .ZN(ADD_1068_U48) );
  XOR2_X1 U11386 ( .A(n10368), .B(n10367), .Z(ADD_1068_U54) );
  XOR2_X1 U11387 ( .A(n10370), .B(n10369), .Z(ADD_1068_U53) );
  XNOR2_X1 U11388 ( .A(n10372), .B(n10371), .ZN(ADD_1068_U52) );
  CLKBUF_X1 U4928 ( .A(n7196), .Z(n8250) );
  CLKBUF_X1 U4951 ( .A(n6418), .Z(n6590) );
  CLKBUF_X1 U5143 ( .A(n5446), .Z(n5572) );
  CLKBUF_X1 U6776 ( .A(n5369), .Z(n5649) );
endmodule

