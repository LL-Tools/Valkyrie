

module b20_C_AntiSAT_k_128_9 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, 
        ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58, 
        ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63, 
        ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51, 
        ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46, 
        U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, 
        P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, 
        P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, 
        P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, 
        P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439, P1_U3440, 
        P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, 
        P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, 
        P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, 
        P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, 
        P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462, P1_U3465, 
        P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, 
        P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, 
        P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, 
        P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, 
        P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, 
        P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, 
        P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, 
        P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, 
        P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291, P1_U3290, 
        P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, 
        P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, 
        P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, 
        P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, 
        P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, 
        P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, 
        P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3554, 
        P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, 
        P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, 
        P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, 
        P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, 
        P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240, P1_U3239, 
        P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, 
        P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, 
        P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, 
        P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, 
        P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, 
        P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, 
        P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, 
        P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, 
        P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376, P2_U3377, 
        P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, 
        P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, 
        P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, 
        P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, 
        P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399, P2_U3402, 
        P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420, P2_U3423, 
        P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441, P2_U3444, 
        P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451, P2_U3452, 
        P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458, P2_U3459, 
        P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465, P2_U3466, 
        P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472, P2_U3473, 
        P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479, P2_U3480, 
        P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486, P2_U3487, 
        P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, 
        P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, 
        P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, 
        P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, 
        P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3491, 
        P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, 
        P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, 
        P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, 
        P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, 
        P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180, P2_U3179, 
        P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, 
        P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, 
        P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, 
        P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151, P2_U3150, 
        P2_U3893 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324,
         n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334,
         n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344,
         n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354,
         n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364,
         n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374,
         n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384,
         n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394,
         n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404,
         n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414,
         n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424,
         n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434,
         n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444,
         n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454,
         n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464,
         n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474,
         n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484,
         n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494,
         n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504,
         n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514,
         n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524,
         n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534,
         n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544,
         n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554,
         n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564,
         n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574,
         n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584,
         n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594,
         n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604,
         n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614,
         n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624,
         n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634,
         n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644,
         n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654,
         n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664,
         n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674,
         n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684,
         n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694,
         n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704,
         n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714,
         n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724,
         n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734,
         n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744,
         n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754,
         n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764,
         n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774,
         n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784,
         n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794,
         n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804,
         n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814,
         n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824,
         n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834,
         n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844,
         n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854,
         n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864,
         n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874,
         n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884,
         n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894,
         n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904,
         n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914,
         n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924,
         n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934,
         n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944,
         n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954,
         n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964,
         n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974,
         n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984,
         n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994,
         n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004,
         n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014,
         n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024,
         n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034,
         n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044,
         n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054,
         n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064,
         n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074,
         n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084,
         n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094,
         n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104,
         n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114,
         n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124,
         n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134,
         n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144,
         n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154,
         n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164,
         n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174,
         n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184,
         n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194,
         n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204,
         n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214,
         n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224,
         n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234,
         n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244,
         n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254,
         n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264,
         n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274,
         n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284,
         n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294,
         n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304,
         n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314,
         n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324,
         n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334,
         n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344,
         n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354,
         n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364,
         n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374,
         n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384,
         n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394,
         n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404,
         n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414,
         n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424,
         n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434,
         n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444,
         n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454,
         n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464,
         n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474,
         n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484,
         n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494,
         n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504,
         n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514,
         n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524,
         n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534,
         n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544,
         n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554,
         n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564,
         n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574,
         n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584,
         n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594,
         n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604,
         n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614,
         n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624,
         n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634,
         n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644,
         n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654,
         n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664,
         n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674,
         n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684,
         n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694,
         n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704,
         n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714,
         n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724,
         n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734,
         n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744,
         n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754,
         n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764,
         n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774,
         n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784,
         n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794,
         n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804,
         n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814,
         n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824,
         n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834,
         n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844,
         n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854,
         n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864,
         n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874,
         n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884,
         n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894,
         n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904,
         n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914,
         n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924,
         n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934,
         n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944,
         n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954,
         n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964,
         n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974,
         n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984,
         n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994,
         n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004,
         n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014,
         n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024,
         n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034,
         n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044,
         n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054,
         n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064,
         n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074,
         n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084,
         n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094,
         n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104,
         n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114,
         n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124,
         n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134,
         n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144,
         n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154,
         n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164,
         n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174,
         n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184,
         n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194,
         n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204,
         n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214,
         n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224,
         n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234,
         n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244,
         n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254,
         n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264,
         n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274,
         n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284,
         n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294,
         n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304,
         n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314,
         n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324,
         n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334,
         n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344,
         n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354,
         n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364,
         n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374,
         n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384,
         n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394,
         n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404,
         n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414,
         n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424,
         n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434,
         n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444,
         n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454,
         n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464,
         n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474,
         n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484,
         n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494,
         n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504,
         n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514,
         n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524,
         n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534,
         n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544,
         n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554,
         n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564,
         n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574,
         n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584,
         n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594,
         n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604,
         n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614,
         n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624,
         n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634,
         n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644,
         n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654,
         n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664,
         n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674,
         n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684,
         n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694,
         n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704,
         n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714,
         n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724,
         n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734,
         n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744,
         n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754,
         n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764,
         n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774,
         n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784,
         n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794,
         n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804,
         n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814,
         n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824,
         n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834,
         n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844,
         n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854,
         n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864,
         n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874,
         n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884,
         n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894,
         n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904,
         n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914,
         n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924,
         n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934,
         n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944,
         n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954,
         n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964,
         n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974,
         n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984,
         n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994,
         n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004,
         n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014,
         n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024,
         n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034,
         n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044,
         n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054,
         n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064,
         n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074,
         n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084,
         n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094,
         n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104,
         n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114,
         n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124,
         n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134,
         n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144,
         n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154,
         n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164,
         n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174,
         n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184,
         n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194,
         n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204,
         n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214,
         n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224,
         n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234,
         n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244,
         n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254,
         n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264,
         n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274,
         n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284,
         n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294,
         n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304,
         n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314,
         n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324,
         n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334,
         n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344,
         n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354,
         n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364,
         n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374,
         n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384,
         n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394,
         n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404,
         n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414,
         n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424,
         n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434,
         n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444,
         n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454,
         n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464,
         n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474,
         n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484,
         n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494,
         n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504,
         n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514,
         n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524,
         n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534,
         n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544,
         n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554,
         n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564,
         n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574,
         n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584,
         n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594,
         n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604,
         n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614,
         n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624,
         n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634,
         n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644,
         n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654,
         n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664,
         n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674,
         n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684,
         n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694,
         n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704,
         n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714,
         n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724,
         n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734,
         n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744,
         n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754,
         n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764,
         n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774,
         n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784,
         n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794,
         n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804,
         n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814,
         n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824,
         n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834,
         n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844,
         n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854,
         n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864,
         n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874,
         n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884,
         n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894,
         n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904,
         n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914,
         n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924,
         n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934,
         n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944,
         n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954,
         n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964,
         n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974,
         n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984,
         n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994,
         n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004,
         n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014,
         n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024,
         n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034,
         n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044,
         n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054,
         n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064,
         n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074,
         n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084,
         n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094,
         n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104,
         n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114,
         n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124,
         n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134,
         n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144,
         n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154,
         n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164,
         n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174,
         n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184,
         n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194,
         n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204,
         n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214,
         n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224,
         n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234,
         n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244,
         n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254,
         n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264,
         n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274,
         n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284,
         n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294,
         n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304,
         n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314,
         n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324,
         n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334,
         n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344,
         n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354,
         n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364,
         n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374,
         n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384,
         n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394,
         n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404,
         n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414,
         n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424,
         n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434,
         n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444,
         n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454,
         n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464,
         n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474,
         n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484,
         n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494,
         n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504,
         n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514,
         n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524,
         n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534,
         n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544,
         n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554,
         n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564,
         n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574,
         n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584,
         n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594,
         n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604,
         n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614,
         n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624,
         n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634,
         n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644,
         n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654,
         n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664,
         n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674,
         n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684,
         n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694,
         n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704,
         n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714,
         n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724,
         n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734,
         n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744,
         n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754,
         n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764,
         n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774,
         n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784,
         n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794,
         n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804,
         n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814,
         n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824,
         n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834,
         n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844,
         n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854,
         n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864,
         n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874,
         n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884,
         n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894,
         n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904,
         n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914,
         n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924,
         n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934,
         n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944,
         n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954,
         n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964,
         n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974,
         n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984,
         n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994,
         n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004,
         n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014,
         n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024,
         n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034,
         n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044,
         n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054,
         n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064,
         n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074,
         n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084,
         n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094,
         n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104,
         n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114,
         n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124,
         n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134,
         n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144,
         n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154,
         n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164,
         n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174,
         n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184,
         n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194,
         n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204,
         n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214,
         n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224,
         n9225, n9226, n9227, n9228, n9230, n9231, n9232, n9233, n9234, n9235,
         n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245,
         n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255,
         n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265,
         n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275,
         n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285,
         n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295,
         n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305,
         n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315,
         n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325,
         n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335,
         n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345,
         n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355,
         n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365,
         n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375,
         n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385,
         n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395,
         n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405,
         n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415,
         n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425,
         n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435,
         n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445,
         n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455,
         n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465,
         n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475,
         n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485,
         n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495,
         n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505,
         n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515,
         n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525,
         n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535,
         n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545,
         n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555,
         n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565,
         n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575,
         n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585,
         n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595,
         n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605,
         n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615,
         n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625,
         n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635,
         n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645,
         n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655,
         n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665,
         n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675,
         n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685,
         n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695,
         n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705,
         n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715,
         n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725,
         n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735,
         n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745,
         n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755,
         n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765,
         n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775,
         n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785,
         n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795,
         n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805,
         n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815,
         n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825,
         n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835,
         n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845,
         n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855,
         n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865,
         n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875,
         n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885,
         n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895,
         n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905,
         n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915,
         n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925,
         n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935,
         n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945,
         n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955,
         n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965,
         n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975,
         n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985,
         n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995,
         n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004,
         n10005, n10006, n10007, n10008, n10009, n10010, n10011, n10012,
         n10013, n10014, n10015, n10016, n10017, n10018, n10019, n10020,
         n10021, n10022, n10023, n10024, n10025, n10026, n10027, n10028,
         n10029, n10030, n10031, n10032, n10033, n10034, n10035, n10036,
         n10037, n10038, n10039, n10040, n10042, n10043, n10044, n10045,
         n10046, n10047, n10048, n10049, n10050, n10051, n10052, n10053,
         n10054, n10055, n10056, n10057, n10058, n10059, n10060, n10061,
         n10062, n10063, n10064, n10065, n10066, n10067, n10068, n10069,
         n10070, n10071, n10072, n10073, n10074, n10075, n10076, n10077,
         n10078, n10079, n10080, n10081, n10082, n10083, n10084, n10085,
         n10086, n10087, n10088, n10089, n10090, n10091, n10092, n10093,
         n10094, n10095, n10096, n10097, n10098, n10099, n10100, n10101,
         n10102, n10103, n10104, n10105, n10106, n10107, n10108, n10109,
         n10110, n10111, n10112, n10113, n10114, n10115, n10116, n10117,
         n10118, n10119, n10120, n10121, n10122, n10123, n10124, n10125,
         n10126, n10127, n10128, n10129, n10130, n10131, n10132, n10133,
         n10134, n10135, n10136, n10137, n10138, n10139, n10140, n10141,
         n10142, n10143, n10144, n10145, n10146, n10147, n10148, n10149,
         n10150, n10151, n10152, n10153, n10154, n10155, n10156, n10157,
         n10158, n10159, n10160, n10161, n10162, n10163, n10164, n10165,
         n10166, n10167, n10168, n10169, n10170, n10171, n10172, n10173,
         n10174, n10175, n10176, n10177, n10178, n10179, n10180, n10181,
         n10182, n10183, n10184, n10185, n10186, n10187, n10188, n10189,
         n10190, n10191, n10192, n10193, n10194, n10195, n10196;

  OAI21_X1 U4821 ( .B1(n9027), .B2(n4855), .A(n4852), .ZN(n9236) );
  AOI21_X1 U4822 ( .B1(n8476), .B2(n8843), .A(n8475), .ZN(n8883) );
  NAND2_X1 U4823 ( .A1(n8752), .A2(n8751), .ZN(n8750) );
  OAI21_X1 U4824 ( .B1(n9069), .B2(n9067), .A(n9066), .ZN(n8126) );
  OR2_X1 U4825 ( .A1(n7733), .A2(n9221), .ZN(n9891) );
  OR2_X1 U4826 ( .A1(n9005), .A2(n8853), .ZN(n8330) );
  INV_X1 U4827 ( .A(n9113), .ZN(n9033) );
  NAND2_X1 U4828 ( .A1(n7654), .A2(n8290), .ZN(n10078) );
  XNOR2_X1 U4829 ( .A(n5804), .B(n5805), .ZN(n6350) );
  INV_X1 U4830 ( .A(n7366), .ZN(n10112) );
  NAND2_X1 U4831 ( .A1(n5799), .A2(n5801), .ZN(n5803) );
  NAND2_X1 U4832 ( .A1(n5983), .A2(n4405), .ZN(n7366) );
  INV_X1 U4833 ( .A(n6013), .ZN(n8409) );
  CLKBUF_X2 U4834 ( .A(n5986), .Z(n6111) );
  INV_X1 U4835 ( .A(n5948), .ZN(n6128) );
  AND3_X1 U4836 ( .A1(n5941), .A2(n5940), .A3(n5939), .ZN(n10097) );
  NAND2_X2 U4837 ( .A1(n8457), .A2(n6272), .ZN(n8226) );
  AND3_X1 U4838 ( .A1(n4815), .A2(n4814), .A3(n4435), .ZN(n4434) );
  INV_X4 U4839 ( .A(n9611), .ZN(n4315) );
  AOI21_X1 U4840 ( .B1(n6783), .B2(n6781), .A(n6782), .ZN(n6899) );
  INV_X1 U4841 ( .A(n5951), .ZN(n6297) );
  INV_X1 U4842 ( .A(n6193), .ZN(n6013) );
  INV_X1 U4843 ( .A(n8226), .ZN(n6127) );
  AOI21_X1 U4844 ( .B1(n9076), .B2(n9201), .A(n4806), .ZN(n4805) );
  OR2_X1 U4845 ( .A1(n7020), .A2(n4947), .ZN(n4810) );
  INV_X1 U4846 ( .A(n5648), .ZN(n5616) );
  NOR2_X1 U4847 ( .A1(n5137), .A2(n4437), .ZN(n5104) );
  NAND2_X1 U4848 ( .A1(n5260), .A2(n6552), .ZN(n5295) );
  XNOR2_X1 U4849 ( .A(n8642), .B(n10017), .ZN(n10024) );
  INV_X1 U4850 ( .A(n8374), .ZN(n8388) );
  NAND2_X1 U4851 ( .A1(n8226), .A2(n6364), .ZN(n5964) );
  OR2_X1 U4852 ( .A1(n9027), .A2(n4851), .ZN(n4425) );
  INV_X1 U4853 ( .A(n5259), .ZN(n5308) );
  CLKBUF_X2 U4854 ( .A(n5283), .Z(n5648) );
  NAND2_X1 U4855 ( .A1(n9430), .A2(n9651), .ZN(n9417) );
  INV_X1 U4856 ( .A(n7600), .ZN(n9927) );
  XNOR2_X1 U4857 ( .A(n5083), .B(n5084), .ZN(n5149) );
  AND4_X1 U4858 ( .A1(n5972), .A2(n5971), .A3(n5970), .A4(n5969), .ZN(n7319)
         );
  AND2_X1 U4859 ( .A1(n7016), .A2(n7015), .ZN(n7021) );
  AND4_X1 U4860 ( .A1(n5323), .A2(n5322), .A3(n5321), .A4(n5320), .ZN(n7597)
         );
  OAI21_X1 U4861 ( .B1(n9453), .B2(n9398), .A(n4944), .ZN(n9439) );
  OR2_X1 U4862 ( .A1(n5799), .A2(n5801), .ZN(n5802) );
  CLKBUF_X3 U4863 ( .A(n8077), .Z(n4316) );
  AND2_X1 U4864 ( .A1(n5570), .A2(n5569), .ZN(n9473) );
  OAI211_X2 U4865 ( .C1(n4862), .C2(n5656), .A(n4858), .B(n4367), .ZN(n4861)
         );
  AOI21_X2 U4866 ( .B1(P2_REG2_REG_12__SCAN_IN), .B2(n8637), .A(n8636), .ZN(
        n8638) );
  AOI21_X2 U4867 ( .B1(n10071), .B2(n8295), .A(n8287), .ZN(n7656) );
  NAND2_X2 U4868 ( .A1(n7391), .A2(n10070), .ZN(n10071) );
  OAI21_X2 U4869 ( .B1(n9086), .B2(n8007), .A(n8006), .ZN(n8117) );
  NAND2_X2 U4870 ( .A1(n4831), .A2(n4830), .ZN(n9086) );
  NAND3_X4 U4871 ( .A1(n6821), .A2(n6820), .A3(n6819), .ZN(n9030) );
  OAI21_X2 U4872 ( .B1(n8765), .B2(n8955), .A(n8750), .ZN(n8739) );
  AOI21_X2 U4873 ( .B1(n8784), .B2(n8244), .A(n8218), .ZN(n8776) );
  NAND2_X2 U4874 ( .A1(n8217), .A2(n8343), .ZN(n8784) );
  XNOR2_X2 U4875 ( .A(n8399), .B(n8451), .ZN(n8727) );
  AOI21_X2 U4876 ( .B1(P2_REG2_REG_14__SCAN_IN), .B2(n8641), .A(n10010), .ZN(
        n8642) );
  OR2_X1 U4877 ( .A1(n8027), .A2(n4658), .ZN(n4654) );
  NAND2_X1 U4878 ( .A1(n5901), .A2(n5900), .ZN(n7822) );
  NAND2_X1 U4879 ( .A1(n7746), .A2(n7600), .ZN(n7504) );
  NAND2_X2 U4880 ( .A1(n7444), .A2(n9270), .ZN(n5768) );
  INV_X2 U4881 ( .A(n6889), .ZN(n5582) );
  INV_X1 U4882 ( .A(n7247), .ZN(n7072) );
  INV_X1 U4883 ( .A(n7228), .ZN(n7467) );
  INV_X1 U4884 ( .A(n8619), .ZN(n7359) );
  INV_X1 U4885 ( .A(n7242), .ZN(n8622) );
  AND4_X1 U4886 ( .A1(n6021), .A2(n6020), .A3(n6019), .A4(n6018), .ZN(n7396)
         );
  NOR2_X1 U4887 ( .A1(n7063), .A2(n7048), .ZN(n8252) );
  AND2_X1 U4888 ( .A1(n5129), .A2(n5166), .ZN(n5375) );
  INV_X4 U4889 ( .A(n6864), .ZN(n9049) );
  NAND2_X1 U4891 ( .A1(n5808), .A2(n5807), .ZN(n6820) );
  XNOR2_X1 U4892 ( .A(n5144), .B(P1_IR_REG_21__SCAN_IN), .ZN(n6814) );
  NAND2_X1 U4893 ( .A1(n5827), .A2(n4353), .ZN(n5867) );
  AND2_X1 U4894 ( .A1(n4460), .A2(n4456), .ZN(n5814) );
  NAND2_X1 U4895 ( .A1(n4425), .A2(n4849), .ZN(n9116) );
  OAI21_X1 U4896 ( .B1(n9439), .B2(n4692), .A(n4690), .ZN(n4685) );
  AND2_X1 U4897 ( .A1(n9638), .A2(n9637), .ZN(n9753) );
  NAND2_X1 U4898 ( .A1(n5646), .A2(n5645), .ZN(n9381) );
  NAND2_X1 U4899 ( .A1(n8209), .A2(n8208), .ZN(n8879) );
  INV_X1 U4900 ( .A(n9077), .ZN(n4806) );
  NAND2_X1 U4901 ( .A1(n5082), .A2(n5081), .ZN(n5083) );
  AND2_X1 U4902 ( .A1(n4654), .A2(n4652), .ZN(n8088) );
  AOI21_X1 U4903 ( .B1(P2_REG2_REG_16__SCAN_IN), .B2(n8646), .A(n10042), .ZN(
        n8647) );
  AND2_X1 U4904 ( .A1(n9886), .A2(n9885), .ZN(n9888) );
  NAND2_X1 U4905 ( .A1(n6143), .A2(n6142), .ZN(n8979) );
  NAND2_X1 U4906 ( .A1(n6130), .A2(n6129), .ZN(n8986) );
  AND2_X1 U4907 ( .A1(n5523), .A2(n5522), .ZN(n9770) );
  NAND2_X1 U4908 ( .A1(n5191), .A2(n5190), .ZN(n9541) );
  OAI211_X1 U4909 ( .C1(n4377), .C2(n5434), .A(n4473), .B(n4471), .ZN(n5481)
         );
  NOR2_X1 U4910 ( .A1(n4653), .A2(n4661), .ZN(n4652) );
  NAND2_X1 U4911 ( .A1(n5508), .A2(n5507), .ZN(n9560) );
  NAND2_X1 U4912 ( .A1(n6140), .A2(n6139), .ZN(n8913) );
  NAND2_X1 U4913 ( .A1(n6120), .A2(n6119), .ZN(n8992) );
  NAND2_X1 U4914 ( .A1(n6098), .A2(n6097), .ZN(n8998) );
  CLKBUF_X1 U4915 ( .A(n9005), .Z(n4431) );
  AND2_X1 U4916 ( .A1(n9606), .A2(n9263), .ZN(n4661) );
  NAND2_X1 U4917 ( .A1(n7486), .A2(n7487), .ZN(n8626) );
  NAND2_X2 U4918 ( .A1(n5898), .A2(n5897), .ZN(n8588) );
  NAND2_X1 U4919 ( .A1(n5467), .A2(n5466), .ZN(n9749) );
  NAND2_X1 U4920 ( .A1(n7276), .A2(n7275), .ZN(n7490) );
  NAND2_X1 U4921 ( .A1(n5451), .A2(n5450), .ZN(n9958) );
  OR2_X1 U4922 ( .A1(n7182), .A2(n7181), .ZN(n7276) );
  NAND2_X1 U4923 ( .A1(n7387), .A2(n7388), .ZN(n10070) );
  NAND2_X1 U4924 ( .A1(n5422), .A2(n5421), .ZN(n9221) );
  NOR2_X1 U4925 ( .A1(n7128), .A2(n7127), .ZN(n7134) );
  OR2_X1 U4926 ( .A1(n5402), .A2(n5401), .ZN(n5403) );
  NAND2_X1 U4927 ( .A1(n5374), .A2(n5373), .ZN(n7984) );
  NAND2_X1 U4928 ( .A1(n7119), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n7185) );
  NAND2_X1 U4929 ( .A1(n4535), .A2(n6027), .ZN(n10134) );
  NAND2_X1 U4930 ( .A1(n6012), .A2(n6011), .ZN(n10125) );
  XNOR2_X1 U4931 ( .A(n4802), .B(n5352), .ZN(n6399) );
  NAND2_X1 U4932 ( .A1(n5001), .A2(n5000), .ZN(n5370) );
  OR2_X1 U4933 ( .A1(n6372), .A2(n5964), .ZN(n5997) );
  NAND2_X1 U4934 ( .A1(n5242), .A2(n5243), .ZN(n6372) );
  NAND2_X1 U4935 ( .A1(n5346), .A2(n5345), .ZN(n6375) );
  CLKBUF_X1 U4936 ( .A(n7129), .Z(n4406) );
  AND2_X1 U4937 ( .A1(n5965), .A2(n4929), .ZN(n6853) );
  NAND2_X1 U4938 ( .A1(n5344), .A2(n5343), .ZN(n5346) );
  AND4_X1 U4939 ( .A1(n5288), .A2(n5287), .A3(n5286), .A4(n5285), .ZN(n7330)
         );
  OAI211_X1 U4940 ( .C1(n5308), .C2(n6365), .A(n5299), .B(n5298), .ZN(n7228)
         );
  NAND2_X1 U4941 ( .A1(n5303), .A2(n4980), .ZN(n5325) );
  NAND4_X2 U4942 ( .A1(n5990), .A2(n5989), .A3(n5988), .A4(n5987), .ZN(n8619)
         );
  INV_X1 U4943 ( .A(n6330), .ZN(n8082) );
  AND2_X1 U4944 ( .A1(n8076), .A2(n5129), .ZN(n5284) );
  NAND4_X1 U4945 ( .A1(n5931), .A2(n5930), .A3(n5929), .A4(n5928), .ZN(n7063)
         );
  OR2_X1 U4946 ( .A1(n8402), .A2(n4428), .ZN(n5982) );
  NAND2_X1 U4947 ( .A1(n5506), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5142) );
  INV_X2 U4948 ( .A(n8412), .ZN(n6264) );
  CLKBUF_X1 U4949 ( .A(n5810), .Z(n8467) );
  NAND2_X2 U4950 ( .A1(n8468), .A2(n9018), .ZN(n8412) );
  NAND2_X1 U4951 ( .A1(n5873), .A2(n9018), .ZN(n6017) );
  INV_X2 U4952 ( .A(n6590), .ZN(n8697) );
  AND2_X1 U4953 ( .A1(n4974), .A2(n4975), .ZN(n5289) );
  NAND2_X1 U4954 ( .A1(n5825), .A2(n5867), .ZN(n8457) );
  NAND2_X1 U4955 ( .A1(n5870), .A2(n5869), .ZN(n9018) );
  NAND2_X1 U4956 ( .A1(n5803), .A2(n5802), .ZN(n7902) );
  NAND2_X1 U4957 ( .A1(n5803), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4808) );
  MUX2_X1 U4958 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5823), .S(
        P2_IR_REG_28__SCAN_IN), .Z(n5825) );
  NAND2_X1 U4959 ( .A1(n4937), .A2(n4935), .ZN(n5850) );
  OR2_X1 U4960 ( .A1(n6243), .A2(n5826), .ZN(n4937) );
  NAND2_X1 U4961 ( .A1(n6243), .A2(n5820), .ZN(n6240) );
  INV_X1 U4962 ( .A(n4826), .ZN(n4825) );
  AND3_X1 U4963 ( .A1(n4436), .A2(n4814), .A3(n5097), .ZN(n5133) );
  NOR2_X1 U4964 ( .A1(n4703), .A2(n4702), .ZN(n4701) );
  INV_X1 U4965 ( .A(n5295), .ZN(n4815) );
  NAND2_X1 U4966 ( .A1(n5105), .A2(n5146), .ZN(n4829) );
  AND2_X1 U4967 ( .A1(n4712), .A2(n4711), .ZN(n5937) );
  INV_X1 U4968 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n4707) );
  NOR2_X1 U4969 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n4704) );
  INV_X1 U4970 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5993) );
  INV_X4 U4971 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  INV_X1 U4972 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n5961) );
  INV_X1 U4973 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n4709) );
  NOR2_X1 U4974 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), .ZN(
        n4435) );
  INV_X1 U4975 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n4711) );
  INV_X1 U4976 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5141) );
  INV_X1 U4977 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n6552) );
  INV_X1 U4978 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n5096) );
  INV_X1 U4979 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5134) );
  NOR2_X2 U4980 ( .A1(n6976), .A2(n6975), .ZN(n6874) );
  INV_X2 U4981 ( .A(n5282), .ZN(n7219) );
  XNOR2_X1 U4982 ( .A(n4754), .B(P2_IR_REG_2__SCAN_IN), .ZN(n8077) );
  NOR2_X2 U4983 ( .A1(n7591), .A2(n7590), .ZN(n7742) );
  NOR2_X2 U4984 ( .A1(n7416), .A2(n7417), .ZN(n7591) );
  OAI22_X2 U4985 ( .A1(n9193), .A2(n9192), .B1(n8123), .B2(n8122), .ZN(n9069)
         );
  AOI21_X2 U4986 ( .B1(n8117), .B2(n8116), .A(n4940), .ZN(n9193) );
  AOI21_X1 U4987 ( .B1(n4670), .B2(n4668), .A(n4369), .ZN(n4667) );
  INV_X1 U4988 ( .A(n4671), .ZN(n4668) );
  AOI21_X1 U4989 ( .B1(n4821), .B2(n4822), .A(n4359), .ZN(n4819) );
  INV_X1 U4990 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n4954) );
  BUF_X1 U4991 ( .A(n5871), .Z(n5873) );
  INV_X1 U4992 ( .A(n9018), .ZN(n5872) );
  NOR2_X1 U4993 ( .A1(n4318), .A2(n4349), .ZN(n4738) );
  NOR2_X1 U4994 ( .A1(n8618), .A2(n7393), .ZN(n4726) );
  NAND2_X1 U4995 ( .A1(n4701), .A2(n5819), .ZN(n4619) );
  AND2_X1 U4996 ( .A1(n5267), .A2(n6363), .ZN(n5259) );
  NAND2_X1 U4997 ( .A1(n8459), .A2(n8453), .ZN(n8374) );
  AND2_X1 U4998 ( .A1(n6820), .A2(n7303), .ZN(n6816) );
  AOI21_X1 U4999 ( .B1(n4667), .B2(n4669), .A(n4358), .ZN(n4664) );
  OAI21_X1 U5000 ( .B1(n5519), .B2(n4887), .A(n4884), .ZN(n5554) );
  INV_X1 U5001 ( .A(n4888), .ZN(n4887) );
  AOI21_X1 U5002 ( .B1(n4888), .B2(n4886), .A(n4885), .ZN(n4884) );
  INV_X1 U5003 ( .A(n5551), .ZN(n4885) );
  OAI21_X1 U5004 ( .B1(n5335), .B2(n4441), .A(n5334), .ZN(n4440) );
  NAND2_X1 U5005 ( .A1(n5737), .A2(n4445), .ZN(n4441) );
  INV_X1 U5006 ( .A(n5736), .ZN(n4445) );
  NAND2_X1 U5007 ( .A1(n5432), .A2(n5431), .ZN(n4472) );
  NAND2_X1 U5008 ( .A1(n4735), .A2(n4737), .ZN(n4732) );
  NOR2_X1 U5009 ( .A1(n4734), .A2(n8206), .ZN(n4733) );
  INV_X1 U5010 ( .A(n4735), .ZN(n4734) );
  INV_X1 U5011 ( .A(n8358), .ZN(n8419) );
  NOR2_X1 U5012 ( .A1(n8624), .A2(n7055), .ZN(n8253) );
  OR2_X1 U5013 ( .A1(n8944), .A2(n8583), .ZN(n8370) );
  OR2_X1 U5014 ( .A1(n8962), .A2(n8774), .ZN(n8360) );
  INV_X1 U5015 ( .A(n4720), .ZN(n4718) );
  NOR2_X1 U5016 ( .A1(n4745), .A2(n8862), .ZN(n4744) );
  NOR2_X1 U5017 ( .A1(n7955), .A2(n4748), .ZN(n4745) );
  OR2_X1 U5018 ( .A1(n8047), .A2(n8596), .ZN(n8324) );
  OR2_X1 U5019 ( .A1(n10134), .A2(n7675), .ZN(n8294) );
  AND2_X1 U5020 ( .A1(n8177), .A2(n8176), .ZN(n8179) );
  NAND2_X1 U5021 ( .A1(n4379), .A2(n4839), .ZN(n4836) );
  NAND2_X1 U5022 ( .A1(n7741), .A2(n7740), .ZN(n4838) );
  OAI21_X1 U5023 ( .B1(n4898), .B2(n5787), .A(n4897), .ZN(n4896) );
  NAND2_X1 U5024 ( .A1(n4859), .A2(n5789), .ZN(n4897) );
  AND2_X1 U5025 ( .A1(n5788), .A2(n9528), .ZN(n4898) );
  OR2_X1 U5026 ( .A1(n9661), .A2(n9242), .ZN(n5723) );
  OR2_X1 U5027 ( .A1(n8096), .A2(n9681), .ZN(n9385) );
  OR2_X1 U5028 ( .A1(n9583), .A2(n9571), .ZN(n5731) );
  NAND2_X1 U5029 ( .A1(n9090), .A2(n4589), .ZN(n7733) );
  NAND2_X1 U5030 ( .A1(n5078), .A2(n5077), .ZN(n5623) );
  AND2_X1 U5031 ( .A1(n5072), .A2(n5071), .ZN(n5597) );
  AND2_X1 U5032 ( .A1(n5067), .A2(n5066), .ZN(n5584) );
  AND2_X1 U5033 ( .A1(n4901), .A2(n4899), .ZN(n5224) );
  INV_X1 U5034 ( .A(n4902), .ZN(n4899) );
  OAI211_X1 U5035 ( .C1(n4958), .C2(n4959), .A(n4905), .B(n4904), .ZN(n4962)
         );
  AND2_X1 U5036 ( .A1(n6050), .A2(n6024), .ZN(n4490) );
  OR2_X1 U5037 ( .A1(n6257), .A2(n8453), .ZN(n4502) );
  AND2_X1 U5038 ( .A1(n6223), .A2(n4500), .ZN(n4499) );
  NAND2_X1 U5039 ( .A1(n6131), .A2(n8570), .ZN(n4927) );
  OR2_X1 U5040 ( .A1(n6131), .A2(n8570), .ZN(n4928) );
  NOR2_X1 U5041 ( .A1(n4621), .A2(n4623), .ZN(n4620) );
  INV_X1 U5042 ( .A(n4938), .ZN(n4623) );
  INV_X1 U5043 ( .A(n4621), .ZN(n4618) );
  AND2_X1 U5044 ( .A1(n6209), .A2(n6208), .ZN(n8576) );
  NAND3_X1 U5045 ( .A1(n6239), .A2(n6238), .A3(n6237), .ZN(n6580) );
  INV_X1 U5046 ( .A(n8039), .ZN(n6237) );
  NAND2_X1 U5047 ( .A1(n8651), .A2(n8652), .ZN(n8708) );
  OR2_X1 U5048 ( .A1(n8986), .A2(n8570), .ZN(n8348) );
  NAND2_X1 U5049 ( .A1(n7660), .A2(n7659), .ZN(n7674) );
  NAND2_X1 U5050 ( .A1(n4723), .A2(n4346), .ZN(n7660) );
  OR2_X1 U5051 ( .A1(n7395), .A2(n4727), .ZN(n4723) );
  NAND2_X1 U5052 ( .A1(n4728), .A2(n10078), .ZN(n4727) );
  INV_X1 U5053 ( .A(n7394), .ZN(n4728) );
  AND2_X1 U5054 ( .A1(n8588), .A2(n8609), .ZN(n4748) );
  OR2_X1 U5055 ( .A1(n8459), .A2(n8453), .ZN(n10118) );
  AND2_X1 U5056 ( .A1(n8076), .A2(n5167), .ZN(n5283) );
  OR2_X1 U5057 ( .A1(n7021), .A2(n7020), .ZN(n4812) );
  AND2_X1 U5058 ( .A1(n8148), .A2(n8151), .ZN(n4432) );
  OR2_X1 U5059 ( .A1(n5600), .A2(n9240), .ZN(n5626) );
  OAI22_X1 U5060 ( .A1(n5721), .A2(n6891), .B1(n6814), .B2(n9373), .ZN(n4459)
         );
  AND2_X1 U5061 ( .A1(n9755), .A2(n6388), .ZN(n5790) );
  AOI21_X1 U5062 ( .B1(n4582), .B2(n4588), .A(n4581), .ZN(n4580) );
  INV_X1 U5063 ( .A(n9391), .ZN(n4581) );
  NOR2_X1 U5064 ( .A1(n8093), .A2(n4672), .ZN(n4671) );
  INV_X1 U5065 ( .A(n4948), .ZN(n4672) );
  AOI21_X1 U5066 ( .B1(n4645), .B2(n4647), .A(n4360), .ZN(n4643) );
  NAND2_X1 U5067 ( .A1(n4660), .A2(n4659), .ZN(n4658) );
  INV_X1 U5068 ( .A(n8087), .ZN(n4659) );
  INV_X1 U5069 ( .A(n8026), .ZN(n4660) );
  NAND2_X1 U5070 ( .A1(n9958), .A2(n9881), .ZN(n4662) );
  BUF_X1 U5071 ( .A(n5310), .Z(n5613) );
  AND2_X1 U5072 ( .A1(n5167), .A2(n5166), .ZN(n5310) );
  AND2_X1 U5073 ( .A1(n5543), .A2(n5542), .ZN(n9693) );
  CLKBUF_X2 U5074 ( .A(n5259), .Z(n5353) );
  NAND2_X1 U5075 ( .A1(n5042), .A2(n5041), .ZN(n5519) );
  NAND2_X1 U5076 ( .A1(n5133), .A2(n5104), .ZN(n5145) );
  NAND2_X1 U5077 ( .A1(n5445), .A2(n5444), .ZN(n5447) );
  NAND3_X1 U5078 ( .A1(n4519), .A2(n4963), .A3(n4517), .ZN(n5258) );
  INV_X1 U5079 ( .A(n4966), .ZN(n4517) );
  AND2_X1 U5080 ( .A1(n4967), .A2(SI_0_), .ZN(n4519) );
  INV_X1 U5081 ( .A(n8941), .ZN(n8887) );
  AND2_X1 U5082 ( .A1(n5806), .A2(n6350), .ZN(n5807) );
  AND2_X1 U5083 ( .A1(n6808), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6316) );
  INV_X1 U5084 ( .A(n4440), .ZN(n4439) );
  AOI21_X1 U5085 ( .B1(n8441), .B2(n8388), .A(n4534), .ZN(n4533) );
  NOR2_X1 U5086 ( .A1(n8330), .A2(n8374), .ZN(n4534) );
  NAND2_X1 U5087 ( .A1(n4472), .A2(n4338), .ZN(n4471) );
  OAI21_X1 U5088 ( .B1(n4531), .B2(n4530), .A(n4529), .ZN(n4528) );
  INV_X1 U5089 ( .A(n8366), .ZN(n4529) );
  NOR2_X1 U5090 ( .A1(n8362), .A2(n8374), .ZN(n4531) );
  OAI21_X1 U5091 ( .B1(n8363), .B2(n8388), .A(n8748), .ZN(n4530) );
  NAND2_X1 U5092 ( .A1(n8369), .A2(n8728), .ZN(n4526) );
  INV_X1 U5093 ( .A(n8740), .ZN(n4527) );
  NAND2_X1 U5094 ( .A1(n8243), .A2(n8242), .ZN(n8376) );
  NAND2_X1 U5095 ( .A1(n5539), .A2(n5582), .ZN(n4479) );
  INV_X1 U5096 ( .A(n5581), .ZN(n4476) );
  AND2_X1 U5097 ( .A1(n5020), .A2(n5027), .ZN(n4865) );
  AND2_X1 U5098 ( .A1(n4453), .A2(n4384), .ZN(n4450) );
  NAND2_X1 U5099 ( .A1(n4452), .A2(n5582), .ZN(n4451) );
  NAND2_X1 U5100 ( .A1(n4955), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n4956) );
  INV_X1 U5101 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4955) );
  NOR2_X1 U5102 ( .A1(n4918), .A2(n4510), .ZN(n4509) );
  INV_X1 U5103 ( .A(n4513), .ZN(n4510) );
  INV_X1 U5104 ( .A(n4919), .ZN(n4918) );
  NOR2_X1 U5105 ( .A1(n4920), .A2(n8502), .ZN(n4919) );
  INV_X1 U5106 ( .A(n4923), .ZN(n4920) );
  OR2_X1 U5107 ( .A1(n6164), .A2(n8607), .ZN(n6165) );
  INV_X1 U5108 ( .A(n7840), .ZN(n4913) );
  AND2_X1 U5109 ( .A1(n6241), .A2(n5820), .ZN(n4938) );
  NOR2_X1 U5110 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), .ZN(
        n5828) );
  OAI21_X1 U5111 ( .B1(n7280), .B2(n7193), .A(n7279), .ZN(n7482) );
  AND2_X1 U5112 ( .A1(n8342), .A2(n8794), .ZN(n8443) );
  AND2_X1 U5113 ( .A1(n8618), .A2(n10119), .ZN(n8281) );
  OR2_X1 U5114 ( .A1(n8973), .A2(n8801), .ZN(n8246) );
  OR2_X1 U5115 ( .A1(n8992), .A2(n8852), .ZN(n8338) );
  NAND2_X1 U5116 ( .A1(n4431), .A2(n8608), .ZN(n4746) );
  AND2_X1 U5117 ( .A1(n7865), .A2(n7864), .ZN(n7866) );
  INV_X1 U5118 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n6241) );
  INV_X1 U5119 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5820) );
  INV_X1 U5120 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n5857) );
  AOI21_X1 U5121 ( .B1(n4836), .B2(n4834), .A(n4372), .ZN(n4833) );
  INV_X1 U5122 ( .A(n4837), .ZN(n4834) );
  INV_X1 U5123 ( .A(n4836), .ZN(n4835) );
  INV_X1 U5124 ( .A(n8148), .ZN(n4845) );
  NOR2_X1 U5125 ( .A1(n4845), .A2(n4842), .ZN(n4841) );
  INV_X1 U5126 ( .A(n8143), .ZN(n4842) );
  OAI21_X1 U5127 ( .B1(n5657), .B2(n9381), .A(n4860), .ZN(n4862) );
  NAND2_X1 U5128 ( .A1(n9381), .A2(n6889), .ZN(n4860) );
  OR2_X1 U5129 ( .A1(n9401), .A2(n9658), .ZN(n5722) );
  INV_X1 U5130 ( .A(n9669), .ZN(n6331) );
  AND2_X1 U5131 ( .A1(n9458), .A2(n9665), .ZN(n9388) );
  OR2_X1 U5132 ( .A1(n9499), .A2(n9680), .ZN(n8100) );
  OR2_X1 U5133 ( .A1(n9514), .A2(n9531), .ZN(n5728) );
  INV_X1 U5134 ( .A(n8098), .ZN(n4566) );
  NAND2_X1 U5135 ( .A1(n9552), .A2(n4418), .ZN(n4417) );
  INV_X1 U5136 ( .A(n5782), .ZN(n4418) );
  OR2_X1 U5137 ( .A1(n4795), .A2(n5750), .ZN(n5771) );
  AND2_X1 U5138 ( .A1(n5747), .A2(n4380), .ZN(n4795) );
  INV_X1 U5139 ( .A(n8076), .ZN(n5166) );
  INV_X1 U5140 ( .A(n9473), .ZN(n8096) );
  NAND2_X1 U5141 ( .A1(n7455), .A2(n7270), .ZN(n7146) );
  NAND2_X1 U5142 ( .A1(n4868), .A2(n4866), .ZN(n5609) );
  AOI21_X1 U5143 ( .B1(n4870), .B2(n4872), .A(n4867), .ZN(n4866) );
  NAND2_X1 U5144 ( .A1(n5585), .A2(n4870), .ZN(n4868) );
  INV_X1 U5145 ( .A(n5072), .ZN(n4867) );
  AND2_X1 U5146 ( .A1(n5061), .A2(n5060), .ZN(n5567) );
  NAND2_X1 U5147 ( .A1(n4828), .A2(n4827), .ZN(n4826) );
  INV_X1 U5148 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n4827) );
  INV_X1 U5149 ( .A(n4829), .ZN(n4828) );
  NAND2_X1 U5150 ( .A1(n5212), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5491) );
  INV_X1 U5151 ( .A(n5418), .ZN(n4875) );
  AOI21_X1 U5152 ( .B1(n4880), .B2(n4878), .A(n4877), .ZN(n4876) );
  INV_X1 U5153 ( .A(n5009), .ZN(n4877) );
  INV_X1 U5154 ( .A(n5369), .ZN(n4878) );
  NAND2_X1 U5155 ( .A1(n5346), .A2(n4352), .ZN(n5001) );
  INV_X1 U5156 ( .A(n4816), .ZN(n4814) );
  OR2_X1 U5157 ( .A1(n6121), .A2(n8825), .ZN(n4513) );
  INV_X1 U5158 ( .A(n8528), .ZN(n4512) );
  AND2_X1 U5159 ( .A1(n7840), .A2(n8613), .ZN(n4915) );
  NAND2_X1 U5160 ( .A1(n6093), .A2(n8853), .ZN(n4931) );
  NOR2_X1 U5161 ( .A1(n8521), .A2(n4934), .ZN(n4930) );
  XNOR2_X1 U5162 ( .A(n6853), .B(n5951), .ZN(n5977) );
  NAND2_X1 U5163 ( .A1(n8547), .A2(n4924), .ZN(n4923) );
  INV_X1 U5164 ( .A(n4927), .ZN(n4924) );
  NAND2_X1 U5165 ( .A1(n7964), .A2(n7965), .ZN(n7963) );
  NAND2_X1 U5166 ( .A1(n4483), .A2(n4488), .ZN(n7605) );
  NAND2_X1 U5167 ( .A1(n6049), .A2(n8614), .ZN(n4488) );
  NAND2_X1 U5168 ( .A1(n7208), .A2(n4325), .ZN(n4483) );
  NAND2_X1 U5169 ( .A1(n4914), .A2(n4913), .ZN(n4910) );
  AND3_X1 U5170 ( .A1(n8407), .A2(n8876), .A3(n8406), .ZN(n4410) );
  AND2_X1 U5171 ( .A1(n6270), .A2(n6269), .ZN(n8382) );
  AND4_X1 U5172 ( .A1(n6087), .A2(n6086), .A3(n6085), .A4(n6084), .ZN(n8596)
         );
  AND4_X1 U5173 ( .A1(n5956), .A2(n5955), .A3(n5954), .A4(n5953), .ZN(n7315)
         );
  NAND2_X1 U5174 ( .A1(n6713), .A2(n6712), .ZN(n6711) );
  NAND2_X1 U5175 ( .A1(n6711), .A2(n4751), .ZN(n4750) );
  NOR2_X1 U5176 ( .A1(n4752), .A2(n6626), .ZN(n4751) );
  INV_X1 U5177 ( .A(n6625), .ZN(n4752) );
  NAND2_X1 U5178 ( .A1(n4753), .A2(n6626), .ZN(n6725) );
  NAND2_X1 U5179 ( .A1(n6711), .A2(n6625), .ZN(n4753) );
  NAND2_X1 U5180 ( .A1(n6725), .A2(n4749), .ZN(n6730) );
  AND2_X1 U5181 ( .A1(n4750), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n4749) );
  NAND2_X1 U5182 ( .A1(n10035), .A2(n10036), .ZN(n10034) );
  CLKBUF_X1 U5183 ( .A(n6272), .Z(n6590) );
  AOI21_X1 U5184 ( .B1(n4612), .B2(n4614), .A(n4609), .ZN(n4608) );
  INV_X1 U5185 ( .A(n8370), .ZN(n4609) );
  AOI21_X1 U5186 ( .B1(n4738), .B2(n4736), .A(n4363), .ZN(n4735) );
  INV_X1 U5187 ( .A(n8204), .ZN(n4736) );
  AOI21_X1 U5188 ( .B1(n4717), .B2(n4718), .A(n4362), .ZN(n4714) );
  INV_X1 U5189 ( .A(n8443), .ZN(n8817) );
  NOR2_X1 U5190 ( .A1(n4626), .A2(n4625), .ZN(n4624) );
  INV_X1 U5191 ( .A(n8307), .ZN(n4625) );
  AND4_X1 U5192 ( .A1(n6033), .A2(n6032), .A3(n6031), .A4(n6030), .ZN(n7675)
         );
  AOI21_X1 U5193 ( .B1(n10078), .B2(n4726), .A(n4365), .ZN(n4725) );
  AND2_X1 U5194 ( .A1(n7655), .A2(n8291), .ZN(n8429) );
  NAND2_X1 U5195 ( .A1(n4697), .A2(n4694), .ZN(n7368) );
  NAND2_X1 U5196 ( .A1(n4698), .A2(n4695), .ZN(n4694) );
  AND2_X1 U5197 ( .A1(n8277), .A2(n8270), .ZN(n7311) );
  NAND2_X1 U5198 ( .A1(n8455), .A2(n8452), .ZN(n6257) );
  NAND2_X1 U5199 ( .A1(n8256), .A2(n8252), .ZN(n4635) );
  NAND2_X1 U5200 ( .A1(n8265), .A2(n8256), .ZN(n7056) );
  NAND2_X1 U5201 ( .A1(n7044), .A2(n7407), .ZN(n7045) );
  AND2_X1 U5202 ( .A1(n8809), .A2(n8817), .ZN(n8807) );
  AND2_X1 U5203 ( .A1(n8370), .A2(n8371), .ZN(n8728) );
  NOR2_X1 U5204 ( .A1(n8222), .A2(n8365), .ZN(n4615) );
  OR2_X1 U5205 ( .A1(n8950), .A2(n8576), .ZN(n8367) );
  NAND2_X1 U5206 ( .A1(n6190), .A2(n6189), .ZN(n8201) );
  OR2_X1 U5207 ( .A1(n8898), .A2(n8774), .ZN(n4943) );
  INV_X1 U5208 ( .A(n8748), .ZN(n8751) );
  NOR2_X1 U5209 ( .A1(n4630), .A2(n4629), .ZN(n4628) );
  INV_X1 U5210 ( .A(n8357), .ZN(n4629) );
  AOI21_X1 U5211 ( .B1(n8797), .B2(n8798), .A(n4364), .ZN(n4720) );
  NAND2_X1 U5212 ( .A1(n8807), .A2(n8797), .ZN(n4716) );
  AOI21_X1 U5213 ( .B1(n4720), .B2(n8444), .A(n8783), .ZN(n4717) );
  OR2_X1 U5214 ( .A1(n8807), .A2(n4718), .ZN(n4713) );
  AND2_X1 U5215 ( .A1(n8348), .A2(n8342), .ZN(n4632) );
  AND2_X1 U5216 ( .A1(n8348), .A2(n8347), .ZN(n8823) );
  NAND2_X1 U5217 ( .A1(n5840), .A2(n5839), .ZN(n9005) );
  AND4_X1 U5218 ( .A1(n6105), .A2(n6104), .A3(n6103), .A4(n6102), .ZN(n8864)
         );
  AND2_X1 U5219 ( .A1(n7956), .A2(n7955), .ZN(n8195) );
  OAI21_X1 U5220 ( .B1(n7956), .B2(n4748), .A(n4744), .ZN(n4747) );
  AND2_X1 U5221 ( .A1(n7062), .A2(n8388), .ZN(n8838) );
  AND2_X1 U5222 ( .A1(n7823), .A2(n4345), .ZN(n7850) );
  INV_X1 U5223 ( .A(n10074), .ZN(n8840) );
  AND2_X1 U5224 ( .A1(n7710), .A2(n7711), .ZN(n8433) );
  OR2_X1 U5225 ( .A1(n7062), .A2(n8374), .ZN(n10074) );
  INV_X1 U5226 ( .A(n8843), .ZN(n10080) );
  INV_X1 U5227 ( .A(n7393), .ZN(n10119) );
  OR2_X1 U5228 ( .A1(n6257), .A2(n8459), .ZN(n10136) );
  AND2_X1 U5229 ( .A1(n6276), .A2(n7039), .ZN(n6752) );
  NOR2_X1 U5230 ( .A1(n6284), .A2(n8458), .ZN(n6754) );
  NAND2_X1 U5231 ( .A1(n4500), .A2(n6757), .ZN(n8843) );
  AND2_X1 U5232 ( .A1(n5852), .A2(n5851), .ZN(n6239) );
  AND2_X1 U5233 ( .A1(n5843), .A2(n5845), .ZN(n6238) );
  XNOR2_X1 U5234 ( .A(n5863), .B(P2_IR_REG_21__SCAN_IN), .ZN(n8453) );
  NOR2_X1 U5235 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n5815) );
  NOR2_X1 U5236 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .ZN(
        n4706) );
  NOR2_X1 U5237 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n4705) );
  NAND2_X1 U5238 ( .A1(n5858), .A2(n5857), .ZN(n4514) );
  AND2_X1 U5239 ( .A1(n5915), .A2(n6065), .ZN(n7492) );
  INV_X1 U5240 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5962) );
  NAND2_X1 U5241 ( .A1(n9058), .A2(n9140), .ZN(n4851) );
  NAND2_X1 U5242 ( .A1(n4322), .A2(n4823), .ZN(n4822) );
  INV_X1 U5243 ( .A(n8155), .ZN(n4823) );
  NAND2_X1 U5244 ( .A1(n4378), .A2(n4322), .ZN(n4821) );
  INV_X1 U5245 ( .A(n9271), .ZN(n7418) );
  AND2_X1 U5246 ( .A1(n9026), .A2(n8182), .ZN(n8186) );
  OR2_X1 U5247 ( .A1(n5524), .A2(n9133), .ZN(n5544) );
  AND2_X1 U5248 ( .A1(n9040), .A2(n4853), .ZN(n4852) );
  AND2_X1 U5249 ( .A1(n9238), .A2(n9235), .ZN(n9040) );
  NAND2_X1 U5250 ( .A1(n9140), .A2(n4854), .ZN(n4853) );
  INV_X1 U5251 ( .A(n9026), .ZN(n4854) );
  AND2_X1 U5252 ( .A1(n6803), .A2(n6802), .ZN(n6828) );
  NAND2_X1 U5253 ( .A1(n4892), .A2(n5791), .ZN(n5792) );
  NAND2_X1 U5254 ( .A1(n4371), .A2(n4893), .ZN(n4892) );
  NAND2_X1 U5255 ( .A1(n4896), .A2(n4894), .ZN(n4893) );
  XNOR2_X1 U5256 ( .A(n6641), .B(n6635), .ZN(n9276) );
  NOR2_X1 U5257 ( .A1(n6926), .A2(n4335), .ZN(n9290) );
  OR2_X1 U5258 ( .A1(n9290), .A2(n9289), .ZN(n4545) );
  OR2_X1 U5259 ( .A1(n9304), .A2(n9303), .ZN(n4541) );
  AND2_X1 U5260 ( .A1(n4541), .A2(n4540), .ZN(n9318) );
  NAND2_X1 U5261 ( .A1(n9309), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n4540) );
  OR2_X1 U5262 ( .A1(n9318), .A2(n9317), .ZN(n4539) );
  NOR2_X1 U5263 ( .A1(n9330), .A2(n4546), .ZN(n6637) );
  NOR2_X1 U5264 ( .A1(n4548), .A2(n4547), .ZN(n4546) );
  INV_X1 U5265 ( .A(n9336), .ZN(n4548) );
  NOR2_X1 U5266 ( .A1(n6637), .A2(n6636), .ZN(n6695) );
  NOR2_X1 U5267 ( .A1(n9804), .A2(n4398), .ZN(n9818) );
  NOR2_X1 U5268 ( .A1(n9843), .A2(n4554), .ZN(n7905) );
  AND2_X1 U5269 ( .A1(n9837), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n4554) );
  NAND2_X1 U5270 ( .A1(n9428), .A2(n4693), .ZN(n4692) );
  INV_X1 U5271 ( .A(n9400), .ZN(n4693) );
  AOI21_X1 U5272 ( .B1(n9428), .B2(n4691), .A(n4370), .ZN(n4690) );
  INV_X1 U5273 ( .A(n9399), .ZN(n4691) );
  NOR2_X1 U5274 ( .A1(n9400), .A2(n4684), .ZN(n4683) );
  OAI21_X1 U5275 ( .B1(n9400), .B2(n4681), .A(n9399), .ZN(n4680) );
  NAND2_X1 U5276 ( .A1(n4944), .A2(n9398), .ZN(n4681) );
  OAI21_X1 U5277 ( .B1(n9461), .B2(n9388), .A(n9387), .ZN(n9442) );
  AND2_X1 U5278 ( .A1(n5724), .A2(n9389), .ZN(n9441) );
  AOI21_X1 U5279 ( .B1(n4671), .B2(n4673), .A(n4356), .ZN(n4670) );
  INV_X1 U5280 ( .A(n9527), .ZN(n4673) );
  AND2_X1 U5281 ( .A1(n5728), .A2(n5727), .ZN(n9508) );
  INV_X1 U5282 ( .A(n9552), .ZN(n4784) );
  AND2_X1 U5283 ( .A1(n4323), .A2(n8090), .ZN(n4649) );
  NAND2_X1 U5284 ( .A1(n4323), .A2(n4361), .ZN(n4648) );
  AND2_X1 U5285 ( .A1(n5729), .A2(n5785), .ZN(n9539) );
  NAND2_X1 U5286 ( .A1(n9563), .A2(n5781), .ZN(n5783) );
  AND2_X1 U5287 ( .A1(n5730), .A2(n5784), .ZN(n9552) );
  AND2_X1 U5288 ( .A1(n4605), .A2(n9719), .ZN(n8089) );
  NAND2_X1 U5289 ( .A1(n4569), .A2(n4568), .ZN(n9563) );
  AOI21_X1 U5290 ( .B1(n4317), .B2(n4571), .A(n5485), .ZN(n4568) );
  NAND2_X1 U5291 ( .A1(n4317), .A2(n4792), .ZN(n4569) );
  INV_X1 U5292 ( .A(n9597), .ZN(n4792) );
  NAND2_X1 U5293 ( .A1(n5215), .A2(n5214), .ZN(n9583) );
  NOR2_X1 U5294 ( .A1(n4657), .A2(n4656), .ZN(n4655) );
  NOR2_X1 U5295 ( .A1(n8087), .A2(n4662), .ZN(n4657) );
  NOR2_X1 U5296 ( .A1(n9631), .A2(n9955), .ZN(n4656) );
  NAND2_X1 U5297 ( .A1(n4792), .A2(n4791), .ZN(n9599) );
  INV_X1 U5298 ( .A(n9596), .ZN(n4791) );
  NOR2_X1 U5299 ( .A1(n9888), .A2(n8025), .ZN(n8027) );
  OR2_X1 U5300 ( .A1(n8027), .A2(n8026), .ZN(n4663) );
  AND2_X1 U5301 ( .A1(n5733), .A2(n9614), .ZN(n8026) );
  NAND2_X1 U5302 ( .A1(n7689), .A2(n7688), .ZN(n7691) );
  AOI21_X1 U5303 ( .B1(n9913), .B2(n6349), .A(n6806), .ZN(n7259) );
  AND2_X1 U5304 ( .A1(n4639), .A2(n7626), .ZN(n4638) );
  NAND3_X1 U5305 ( .A1(n7511), .A2(n7353), .A3(n7352), .ZN(n4640) );
  NAND2_X1 U5306 ( .A1(n6399), .A2(n5353), .ZN(n4801) );
  AND4_X1 U5307 ( .A1(n5252), .A2(n5251), .A3(n5250), .A4(n5249), .ZN(n7746)
         );
  OAI211_X1 U5308 ( .C1(n4463), .C2(n4468), .A(n5739), .B(n4462), .ZN(n7328)
         );
  NAND3_X1 U5309 ( .A1(n4461), .A2(n5670), .A3(n5738), .ZN(n4462) );
  NAND2_X1 U5310 ( .A1(n5738), .A2(n5670), .ZN(n4463) );
  INV_X1 U5311 ( .A(n4466), .ZN(n4461) );
  NAND2_X1 U5312 ( .A1(n4464), .A2(n5670), .ZN(n7224) );
  NAND2_X1 U5313 ( .A1(n4468), .A2(n4466), .ZN(n4464) );
  INV_X1 U5314 ( .A(n9645), .ZN(n4798) );
  INV_X1 U5315 ( .A(n9643), .ZN(n4797) );
  AND2_X1 U5316 ( .A1(n5607), .A2(n5606), .ZN(n9657) );
  AND2_X1 U5317 ( .A1(n5579), .A2(n5578), .ZN(n9681) );
  NAND2_X1 U5318 ( .A1(n5556), .A2(n5555), .ZN(n9684) );
  INV_X1 U5319 ( .A(n9954), .ZN(n9880) );
  INV_X1 U5320 ( .A(n7339), .ZN(n9921) );
  INV_X1 U5321 ( .A(n6802), .ZN(n7260) );
  OAI21_X1 U5322 ( .B1(n5267), .B2(n6641), .A(n4433), .ZN(n6330) );
  NAND2_X1 U5323 ( .A1(n5267), .A2(n4599), .ZN(n4433) );
  OAI22_X1 U5324 ( .A1(n4602), .A2(n6364), .B1(n4600), .B2(n6363), .ZN(n4599)
         );
  NAND2_X1 U5325 ( .A1(n7148), .A2(n7147), .ZN(n9952) );
  NAND2_X1 U5326 ( .A1(n8467), .A2(n7147), .ZN(n9954) );
  NAND2_X1 U5327 ( .A1(n9620), .A2(n9914), .ZN(n9964) );
  INV_X1 U5328 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5119) );
  XNOR2_X1 U5329 ( .A(n5643), .B(n5642), .ZN(n8464) );
  XNOR2_X1 U5330 ( .A(n5609), .B(n5610), .ZN(n8072) );
  XNOR2_X1 U5331 ( .A(n5596), .B(n5597), .ZN(n8065) );
  NAND2_X1 U5332 ( .A1(n4869), .A2(n5067), .ZN(n5596) );
  AOI21_X1 U5333 ( .B1(n4890), .B2(n5045), .A(n4889), .ZN(n4888) );
  INV_X1 U5334 ( .A(n5050), .ZN(n4889) );
  NOR2_X1 U5335 ( .A1(n5541), .A2(n4891), .ZN(n4890) );
  INV_X1 U5336 ( .A(n5044), .ZN(n4891) );
  OAI21_X1 U5337 ( .B1(n5519), .B2(n5045), .A(n5044), .ZN(n5540) );
  OR2_X1 U5338 ( .A1(n5448), .A2(P1_IR_REG_13__SCAN_IN), .ZN(n5225) );
  NAND2_X1 U5339 ( .A1(n5403), .A2(n5012), .ZN(n5445) );
  AND2_X1 U5340 ( .A1(n5017), .A2(n5016), .ZN(n5444) );
  AND2_X1 U5341 ( .A1(n5408), .A2(n5448), .ZN(n7910) );
  NOR2_X1 U5342 ( .A1(n5383), .A2(n5004), .ZN(n4880) );
  XNOR2_X1 U5343 ( .A(n5370), .B(n5369), .ZN(n6600) );
  INV_X1 U5344 ( .A(n4990), .ZN(n4786) );
  NAND2_X1 U5345 ( .A1(n5325), .A2(n5324), .ZN(n5327) );
  NAND2_X1 U5346 ( .A1(n5096), .A2(n4817), .ZN(n4816) );
  INV_X1 U5347 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n4817) );
  NAND2_X1 U5348 ( .A1(n4970), .A2(n4777), .ZN(n5275) );
  NAND2_X1 U5349 ( .A1(n4779), .A2(n4778), .ZN(n4777) );
  INV_X1 U5350 ( .A(SI_2_), .ZN(n4778) );
  INV_X1 U5351 ( .A(n4968), .ZN(n4779) );
  NAND2_X1 U5352 ( .A1(n5258), .A2(n4967), .ZN(n5274) );
  NAND2_X1 U5353 ( .A1(n4961), .A2(n4960), .ZN(n4963) );
  INV_X1 U5354 ( .A(n4962), .ZN(n4961) );
  NAND2_X1 U5355 ( .A1(n4520), .A2(n4515), .ZN(n4966) );
  NAND2_X1 U5356 ( .A1(n4518), .A2(n4516), .ZN(n4515) );
  OR2_X1 U5357 ( .A1(n4518), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n4520) );
  NAND2_X1 U5358 ( .A1(n7963), .A2(n4492), .ZN(n8040) );
  NAND2_X1 U5359 ( .A1(n4493), .A2(n8045), .ZN(n4492) );
  INV_X1 U5360 ( .A(n6077), .ZN(n4493) );
  NAND2_X1 U5361 ( .A1(n6167), .A2(n6166), .ZN(n8489) );
  NAND2_X1 U5362 ( .A1(n4511), .A2(n4513), .ZN(n8493) );
  AND4_X1 U5363 ( .A1(n5888), .A2(n5887), .A3(n5886), .A4(n5885), .ZN(n8863)
         );
  AND3_X1 U5364 ( .A1(n6126), .A2(n6125), .A3(n6124), .ZN(n8570) );
  INV_X1 U5365 ( .A(n7675), .ZN(n8615) );
  NAND2_X1 U5366 ( .A1(n8708), .A2(n8707), .ZN(n4773) );
  AOI21_X1 U5367 ( .B1(n4326), .B2(n10057), .A(n4769), .ZN(n4413) );
  NAND2_X1 U5368 ( .A1(n6064), .A2(n6063), .ZN(n10140) );
  INV_X1 U5369 ( .A(n8819), .ZN(n8872) );
  OR2_X1 U5370 ( .A1(n5964), .A2(n6362), .ZN(n5922) );
  NAND2_X1 U5371 ( .A1(n4337), .A2(n10104), .ZN(n8882) );
  AND2_X1 U5372 ( .A1(n6296), .A2(n6295), .ZN(n8941) );
  INV_X1 U5373 ( .A(n7127), .ZN(n4416) );
  NAND2_X1 U5374 ( .A1(n8152), .A2(n9225), .ZN(n9104) );
  AND3_X1 U5375 ( .A1(n5184), .A2(n5183), .A3(n5182), .ZN(n9709) );
  INV_X1 U5376 ( .A(n9762), .ZN(n9458) );
  OR2_X1 U5377 ( .A1(n6846), .A2(n5308), .ZN(n5451) );
  NAND2_X1 U5378 ( .A1(n4407), .A2(n9076), .ZN(n9200) );
  NAND2_X1 U5379 ( .A1(n4420), .A2(n4419), .ZN(n4407) );
  INV_X1 U5380 ( .A(n8164), .ZN(n4419) );
  NAND2_X1 U5381 ( .A1(n5231), .A2(n5230), .ZN(n9606) );
  XNOR2_X1 U5382 ( .A(n5143), .B(P1_IR_REG_22__SCAN_IN), .ZN(n6884) );
  INV_X1 U5383 ( .A(n9556), .ZN(n9719) );
  INV_X1 U5384 ( .A(n9092), .ZN(n9266) );
  AND2_X1 U5385 ( .A1(n4543), .A2(n4542), .ZN(n6944) );
  INV_X1 U5386 ( .A(n6945), .ZN(n4542) );
  OR2_X1 U5387 ( .A1(n6658), .A2(n6920), .ZN(n9857) );
  INV_X1 U5388 ( .A(n9861), .ZN(n9842) );
  INV_X1 U5389 ( .A(n4676), .ZN(n4675) );
  OAI21_X1 U5390 ( .B1(n4799), .B2(n9962), .A(n4403), .ZN(n9644) );
  OAI21_X1 U5391 ( .B1(n4580), .B2(n9403), .A(n4573), .ZN(n4572) );
  NAND2_X1 U5392 ( .A1(n6831), .A2(n6830), .ZN(n9532) );
  AND2_X1 U5393 ( .A1(n5117), .A2(n5116), .ZN(n9755) );
  NAND2_X1 U5394 ( .A1(n4595), .A2(n9573), .ZN(n9638) );
  XNOR2_X1 U5395 ( .A(n9376), .B(n9755), .ZN(n4595) );
  NOR2_X1 U5396 ( .A1(n9966), .A2(n4598), .ZN(n4597) );
  INV_X1 U5397 ( .A(n9637), .ZN(n4598) );
  NAND2_X1 U5398 ( .A1(n5392), .A2(n5391), .ZN(n8000) );
  NAND2_X1 U5399 ( .A1(n9968), .A2(n9959), .ZN(n9788) );
  NAND2_X1 U5400 ( .A1(n5333), .A2(n4447), .ZN(n4446) );
  NOR2_X1 U5401 ( .A1(n5677), .A2(n4392), .ZN(n4447) );
  OR3_X1 U5402 ( .A1(n5735), .A2(n9264), .A3(n6889), .ZN(n5437) );
  NAND2_X1 U5403 ( .A1(n8335), .A2(n4340), .ZN(n8350) );
  NAND2_X1 U5404 ( .A1(n4470), .A2(n4469), .ZN(n5477) );
  AND2_X1 U5405 ( .A1(n5777), .A2(n6889), .ZN(n4469) );
  OAI21_X1 U5406 ( .B1(n5481), .B2(n5476), .A(n5776), .ZN(n4470) );
  OAI21_X1 U5407 ( .B1(n4537), .B2(n4536), .A(n8355), .ZN(n8359) );
  OAI21_X1 U5408 ( .B1(n8354), .B2(n8388), .A(n8783), .ZN(n4536) );
  AOI21_X1 U5409 ( .B1(n8345), .B2(n8344), .A(n8374), .ZN(n4537) );
  NOR2_X1 U5410 ( .A1(n4525), .A2(n4524), .ZN(n8373) );
  INV_X1 U5411 ( .A(n8372), .ZN(n4524) );
  AOI21_X1 U5412 ( .B1(n4528), .B2(n4527), .A(n4526), .ZN(n4525) );
  INV_X1 U5413 ( .A(n5583), .ZN(n4474) );
  INV_X1 U5414 ( .A(n5722), .ZN(n4452) );
  AND2_X1 U5415 ( .A1(n5723), .A2(n6889), .ZN(n4454) );
  NOR2_X1 U5416 ( .A1(n8384), .A2(n8383), .ZN(n8389) );
  NOR2_X1 U5417 ( .A1(n8979), .A2(n8560), .ZN(n8351) );
  NAND2_X1 U5418 ( .A1(n7926), .A2(n7925), .ZN(n4839) );
  INV_X1 U5419 ( .A(n5067), .ZN(n4872) );
  INV_X1 U5420 ( .A(n4871), .ZN(n4870) );
  OAI21_X1 U5421 ( .B1(n5584), .B2(n4872), .A(n5597), .ZN(n4871) );
  INV_X1 U5422 ( .A(n5520), .ZN(n5043) );
  INV_X1 U5423 ( .A(SI_19_), .ZN(n5028) );
  NAND2_X1 U5424 ( .A1(n4393), .A2(n5027), .ZN(n4864) );
  INV_X1 U5425 ( .A(SI_15_), .ZN(n4900) );
  NOR2_X1 U5426 ( .A1(n5459), .A2(SI_14_), .ZN(n4902) );
  NAND2_X1 U5427 ( .A1(n5447), .A2(n4391), .ZN(n4901) );
  NAND2_X1 U5428 ( .A1(n5459), .A2(SI_14_), .ZN(n4903) );
  OR2_X1 U5429 ( .A1(n6199), .A2(n8741), .ZN(n6200) );
  NAND2_X1 U5430 ( .A1(n4710), .A2(n4622), .ZN(n4621) );
  INV_X1 U5431 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n4622) );
  AND2_X1 U5432 ( .A1(n7002), .A2(n7001), .ZN(n7003) );
  INV_X1 U5433 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n6320) );
  INV_X1 U5434 ( .A(n7003), .ZN(n4761) );
  INV_X1 U5435 ( .A(n7496), .ZN(n4758) );
  NAND2_X1 U5436 ( .A1(n8626), .A2(n8627), .ZN(n8628) );
  INV_X1 U5437 ( .A(n4613), .ZN(n4612) );
  OAI21_X1 U5438 ( .B1(n4615), .B2(n4614), .A(n8371), .ZN(n4613) );
  INV_X1 U5439 ( .A(n8367), .ZN(n4614) );
  NOR2_X1 U5440 ( .A1(n6216), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n6260) );
  NOR2_X1 U5441 ( .A1(n6170), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6179) );
  NOR2_X1 U5442 ( .A1(n6122), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n6133) );
  AND2_X1 U5443 ( .A1(n5877), .A2(n5876), .ZN(n6099) );
  NOR2_X1 U5444 ( .A1(n6083), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5877) );
  NOR2_X1 U5445 ( .A1(n6069), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5902) );
  INV_X1 U5446 ( .A(n8302), .ZN(n4626) );
  OR2_X1 U5447 ( .A1(n6051), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n6053) );
  AND2_X1 U5448 ( .A1(n6014), .A2(n6320), .ZN(n6028) );
  NAND2_X1 U5449 ( .A1(n4700), .A2(n4699), .ZN(n4698) );
  INV_X1 U5450 ( .A(n7362), .ZN(n4699) );
  INV_X1 U5451 ( .A(n7364), .ZN(n4700) );
  OR2_X1 U5452 ( .A1(n7364), .A2(n4696), .ZN(n4695) );
  INV_X1 U5453 ( .A(n7365), .ZN(n4696) );
  AND2_X1 U5454 ( .A1(n6225), .A2(n6376), .ZN(n7037) );
  INV_X1 U5455 ( .A(n8418), .ZN(n4630) );
  INV_X1 U5456 ( .A(n8351), .ZN(n8343) );
  OR2_X1 U5457 ( .A1(n8998), .A2(n8864), .ZN(n8333) );
  OR2_X1 U5458 ( .A1(n8588), .A2(n8863), .ZN(n8331) );
  NAND2_X1 U5459 ( .A1(n4953), .A2(n7710), .ZN(n7823) );
  INV_X1 U5460 ( .A(n4936), .ZN(n4935) );
  OAI21_X1 U5461 ( .B1(n4938), .B2(n5826), .A(n5830), .ZN(n4936) );
  OR2_X1 U5462 ( .A1(n5827), .A2(n5826), .ZN(n5842) );
  AND2_X1 U5463 ( .A1(n4839), .A2(n7740), .ZN(n4837) );
  INV_X2 U5464 ( .A(n7129), .ZN(n9044) );
  NOR2_X1 U5465 ( .A1(n5790), .A2(n4895), .ZN(n4894) );
  AND2_X1 U5466 ( .A1(n9381), .A2(n5654), .ZN(n4895) );
  NAND2_X1 U5467 ( .A1(n5658), .A2(n4857), .ZN(n4856) );
  NOR2_X1 U5468 ( .A1(n9381), .A2(n5582), .ZN(n4857) );
  NAND2_X1 U5469 ( .A1(n4689), .A2(n4333), .ZN(n4688) );
  INV_X1 U5470 ( .A(n4692), .ZN(n4689) );
  INV_X1 U5471 ( .A(n9415), .ZN(n4584) );
  OR2_X1 U5472 ( .A1(n6331), .A2(n9657), .ZN(n5724) );
  INV_X1 U5473 ( .A(n4670), .ZN(n4669) );
  OR2_X1 U5474 ( .A1(n9705), .A2(n9709), .ZN(n8098) );
  INV_X1 U5475 ( .A(n4648), .ZN(n4647) );
  INV_X1 U5476 ( .A(n4646), .ZN(n4645) );
  OAI21_X1 U5477 ( .B1(n4649), .B2(n4647), .A(n8091), .ZN(n4646) );
  OR2_X1 U5478 ( .A1(n9541), .A2(n9718), .ZN(n8091) );
  NOR2_X1 U5479 ( .A1(n9606), .A2(n9749), .ZN(n4604) );
  INV_X1 U5480 ( .A(n4655), .ZN(n4653) );
  INV_X1 U5481 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n5452) );
  OR2_X1 U5482 ( .A1(n5453), .A2(n5452), .ZN(n5469) );
  AND2_X1 U5483 ( .A1(n6815), .A2(n7147), .ZN(n6806) );
  INV_X1 U5484 ( .A(n7509), .ZN(n4641) );
  INV_X1 U5485 ( .A(n7328), .ZN(n4563) );
  NOR2_X1 U5486 ( .A1(n5268), .A2(n4467), .ZN(n4466) );
  OR2_X1 U5487 ( .A1(n9684), .A2(n9494), .ZN(n9481) );
  INV_X1 U5488 ( .A(n9770), .ZN(n9514) );
  NOR2_X1 U5489 ( .A1(n4592), .A2(n4594), .ZN(n7646) );
  AND2_X1 U5490 ( .A1(n6884), .A2(n6814), .ZN(n7147) );
  AND2_X1 U5491 ( .A1(n5077), .A2(n5076), .ZN(n5610) );
  INV_X1 U5492 ( .A(n4890), .ZN(n4886) );
  INV_X1 U5493 ( .A(SI_20_), .ZN(n5173) );
  INV_X1 U5494 ( .A(n5039), .ZN(n5503) );
  INV_X1 U5495 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n6529) );
  OAI21_X1 U5496 ( .B1(n6363), .B2(n4412), .A(n4411), .ZN(n4986) );
  NAND2_X1 U5497 ( .A1(n6363), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n4411) );
  OAI21_X1 U5498 ( .B1(n6363), .B2(n4428), .A(n4427), .ZN(n4981) );
  NAND2_X1 U5499 ( .A1(n6363), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n4427) );
  OAI211_X1 U5500 ( .C1(n4958), .C2(n4776), .A(n4775), .B(n4774), .ZN(n4968)
         );
  NAND2_X1 U5501 ( .A1(n4906), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n4775) );
  AOI21_X1 U5502 ( .B1(n4926), .B2(n4919), .A(n4917), .ZN(n4916) );
  INV_X1 U5503 ( .A(n8501), .ZN(n4917) );
  AOI21_X1 U5504 ( .B1(n8536), .B2(n8788), .A(n4507), .ZN(n4504) );
  INV_X1 U5505 ( .A(n8537), .ZN(n4507) );
  OAI21_X1 U5506 ( .B1(n4914), .B2(n4912), .A(n4911), .ZN(n7964) );
  AOI21_X1 U5507 ( .B1(n4908), .B2(n7883), .A(n4334), .ZN(n4911) );
  NAND2_X1 U5508 ( .A1(n8499), .A2(n6154), .ZN(n8556) );
  INV_X1 U5509 ( .A(n4490), .ZN(n4487) );
  INV_X1 U5510 ( .A(n7606), .ZN(n4486) );
  XNOR2_X1 U5511 ( .A(n7241), .B(n5951), .ZN(n5957) );
  NAND2_X1 U5512 ( .A1(n4932), .A2(n4351), .ZN(n6108) );
  NAND2_X1 U5513 ( .A1(n8408), .A2(n8932), .ZN(n4409) );
  XNOR2_X1 U5514 ( .A(n4316), .B(n7174), .ZN(n6713) );
  OAI21_X1 U5515 ( .B1(n4316), .B2(n6619), .A(n4421), .ZN(n6709) );
  NAND2_X1 U5516 ( .A1(n4316), .A2(n6619), .ZN(n4421) );
  NAND2_X1 U5517 ( .A1(n6678), .A2(n6789), .ZN(n6781) );
  OR2_X1 U5518 ( .A1(n6680), .A2(n6679), .ZN(n6783) );
  NOR2_X1 U5519 ( .A1(n6901), .A2(n10090), .ZN(n7004) );
  NOR2_X1 U5520 ( .A1(n7004), .A2(n7003), .ZN(n7006) );
  XNOR2_X1 U5521 ( .A(n7183), .B(n7177), .ZN(n7119) );
  OAI21_X1 U5522 ( .B1(n7004), .B2(n4760), .A(n4759), .ZN(n7176) );
  NAND2_X1 U5523 ( .A1(n7005), .A2(n4762), .ZN(n4759) );
  NAND2_X1 U5524 ( .A1(n4761), .A2(n4762), .ZN(n4760) );
  NAND2_X1 U5525 ( .A1(n7104), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n4762) );
  INV_X1 U5526 ( .A(n7490), .ZN(n7491) );
  NAND2_X1 U5527 ( .A1(n4755), .A2(n4757), .ZN(n8636) );
  NAND2_X1 U5528 ( .A1(n7494), .A2(n4758), .ZN(n4757) );
  OR2_X1 U5529 ( .A1(n7277), .A2(n4756), .ZN(n4755) );
  NAND2_X1 U5530 ( .A1(n4758), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n4756) );
  XNOR2_X1 U5531 ( .A(n8638), .B(n9984), .ZN(n9996) );
  OR2_X1 U5532 ( .A1(n6065), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n5891) );
  OAI21_X1 U5533 ( .B1(n9996), .B2(n4764), .A(n4763), .ZN(n10010) );
  NAND2_X1 U5534 ( .A1(n4765), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n4764) );
  NAND2_X1 U5535 ( .A1(n8639), .A2(n4765), .ZN(n4763) );
  INV_X1 U5536 ( .A(n10011), .ZN(n4765) );
  NOR2_X1 U5537 ( .A1(n9996), .A2(n9995), .ZN(n9994) );
  NAND2_X1 U5538 ( .A1(n4768), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n4767) );
  NAND2_X1 U5539 ( .A1(n8644), .A2(n4768), .ZN(n4766) );
  INV_X1 U5540 ( .A(n10043), .ZN(n4768) );
  NAND2_X1 U5541 ( .A1(n4415), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n8650) );
  NAND2_X1 U5542 ( .A1(n8650), .A2(n8649), .ZN(n8651) );
  NAND2_X1 U5543 ( .A1(n10034), .A2(n4402), .ZN(n8634) );
  NAND2_X1 U5544 ( .A1(n10049), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n4770) );
  INV_X1 U5545 ( .A(n4731), .ZN(n4730) );
  OAI22_X1 U5546 ( .A1(n4732), .A2(n8206), .B1(n8941), .B2(n8382), .ZN(n4731)
         );
  AND2_X1 U5547 ( .A1(n8416), .A2(n6305), .ZN(n8474) );
  INV_X1 U5548 ( .A(n4738), .ZN(n4737) );
  OR2_X1 U5549 ( .A1(n6157), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6170) );
  NAND2_X1 U5550 ( .A1(n6099), .A2(n6529), .ZN(n6109) );
  OAI21_X1 U5551 ( .B1(n7395), .B2(n7394), .A(n4724), .ZN(n10079) );
  INV_X1 U5552 ( .A(n4726), .ZN(n4724) );
  AND4_X1 U5553 ( .A1(n6040), .A2(n6039), .A3(n6038), .A4(n6037), .ZN(n10075)
         );
  NAND2_X1 U5554 ( .A1(n4637), .A2(n4636), .ZN(n7388) );
  AND2_X1 U5555 ( .A1(n8271), .A2(n8277), .ZN(n4636) );
  NAND2_X1 U5556 ( .A1(n7164), .A2(n7163), .ZN(n7251) );
  OR2_X1 U5557 ( .A1(n8807), .A2(n8798), .ZN(n4719) );
  AND2_X1 U5558 ( .A1(n7043), .A2(n7042), .ZN(n7407) );
  AND2_X1 U5559 ( .A1(n8202), .A2(n8220), .ZN(n8748) );
  AOI22_X1 U5560 ( .A1(n8772), .A2(n8200), .B1(n8561), .B2(n8970), .ZN(n8762)
         );
  NAND2_X1 U5561 ( .A1(n4746), .A2(n4743), .ZN(n4742) );
  INV_X1 U5562 ( .A(n4748), .ZN(n4743) );
  NOR2_X1 U5563 ( .A1(n8850), .A2(n8851), .ZN(n8849) );
  AND4_X1 U5564 ( .A1(n6115), .A2(n6114), .A3(n6113), .A4(n6112), .ZN(n8852)
         );
  INV_X1 U5565 ( .A(n8441), .ZN(n8851) );
  NAND2_X1 U5566 ( .A1(n7859), .A2(n4722), .ZN(n7867) );
  AND2_X1 U5567 ( .A1(n7860), .A2(n7866), .ZN(n4722) );
  NAND2_X1 U5568 ( .A1(n7853), .A2(n7852), .ZN(n7860) );
  NAND2_X1 U5569 ( .A1(n4721), .A2(n8321), .ZN(n7954) );
  INV_X1 U5570 ( .A(n7867), .ZN(n4721) );
  NAND2_X1 U5571 ( .A1(n6240), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6242) );
  INV_X1 U5572 ( .A(n8458), .ZN(n7039) );
  XNOR2_X1 U5573 ( .A(n5866), .B(P2_IR_REG_30__SCAN_IN), .ZN(n5871) );
  NAND2_X1 U5574 ( .A1(n5869), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5866) );
  INV_X1 U5575 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n4739) );
  NAND2_X1 U5576 ( .A1(n5817), .A2(n4710), .ZN(n4617) );
  XNOR2_X1 U5577 ( .A(n5859), .B(P2_IR_REG_19__SCAN_IN), .ZN(n8455) );
  NAND2_X1 U5578 ( .A1(n6117), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5859) );
  OR2_X1 U5579 ( .A1(n5856), .A2(P2_IR_REG_16__SCAN_IN), .ZN(n6094) );
  AND2_X1 U5580 ( .A1(n6062), .A2(n6061), .ZN(n7280) );
  AND2_X1 U5581 ( .A1(n6010), .A2(n6009), .ZN(n6995) );
  OR2_X1 U5582 ( .A1(n5979), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n5992) );
  AND2_X1 U5583 ( .A1(n5937), .A2(n5938), .ZN(n5946) );
  AND2_X1 U5584 ( .A1(n8184), .A2(n8174), .ZN(n9077) );
  OR2_X1 U5585 ( .A1(n5396), .A2(n9919), .ZN(n5273) );
  NAND2_X1 U5586 ( .A1(n9027), .A2(n9026), .ZN(n9139) );
  OR2_X1 U5587 ( .A1(n5471), .A2(n5232), .ZN(n5234) );
  INV_X1 U5588 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n8059) );
  NAND2_X1 U5589 ( .A1(n4832), .A2(n4836), .ZN(n9169) );
  NAND2_X1 U5590 ( .A1(n7742), .A2(n4837), .ZN(n4832) );
  INV_X1 U5591 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n5376) );
  OR2_X1 U5592 ( .A1(n5194), .A2(n9186), .ZN(n5524) );
  AOI21_X1 U5593 ( .B1(n4833), .B2(n4835), .A(n4373), .ZN(n4830) );
  NAND2_X1 U5594 ( .A1(n4840), .A2(n4843), .ZN(n9224) );
  INV_X1 U5595 ( .A(n4844), .ZN(n4843) );
  OAI21_X1 U5596 ( .B1(n4336), .B2(n4845), .A(n8150), .ZN(n4844) );
  OR2_X1 U5597 ( .A1(n5494), .A2(n8059), .ZN(n5510) );
  NAND2_X1 U5598 ( .A1(n4545), .A2(n4544), .ZN(n4543) );
  NAND2_X1 U5599 ( .A1(n9295), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n4544) );
  NAND2_X1 U5600 ( .A1(n9323), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n4538) );
  NOR2_X1 U5601 ( .A1(n6695), .A2(n4388), .ZN(n6698) );
  NAND2_X1 U5602 ( .A1(n6698), .A2(n6697), .ZN(n7084) );
  NOR2_X1 U5603 ( .A1(n9818), .A2(n9817), .ZN(n9816) );
  NOR2_X1 U5604 ( .A1(n9816), .A2(n4549), .ZN(n7088) );
  NOR2_X1 U5605 ( .A1(n4551), .A2(n4550), .ZN(n4549) );
  INV_X1 U5606 ( .A(n9821), .ZN(n4551) );
  NAND2_X1 U5607 ( .A1(n7088), .A2(n7087), .ZN(n7904) );
  NOR2_X1 U5608 ( .A1(n9825), .A2(n4555), .ZN(n9844) );
  AND2_X1 U5609 ( .A1(n9833), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n4555) );
  NOR2_X1 U5610 ( .A1(n9844), .A2(n9845), .ZN(n9843) );
  XNOR2_X1 U5611 ( .A(n7905), .B(n9856), .ZN(n9860) );
  NAND2_X1 U5612 ( .A1(n5140), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5504) );
  INV_X1 U5613 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5139) );
  NOR2_X1 U5614 ( .A1(n4688), .A2(n4684), .ZN(n4678) );
  OAI21_X1 U5615 ( .B1(n4688), .B2(n4677), .A(n4686), .ZN(n4676) );
  NAND2_X1 U5616 ( .A1(n4944), .A2(n9398), .ZN(n4677) );
  NAND2_X1 U5617 ( .A1(n4687), .A2(n4333), .ZN(n4686) );
  NAND2_X1 U5618 ( .A1(n4690), .A2(n9402), .ZN(n4687) );
  NAND2_X1 U5619 ( .A1(n4580), .A2(n4574), .ZN(n4573) );
  NAND2_X1 U5620 ( .A1(n4583), .A2(n4577), .ZN(n4574) );
  OR2_X1 U5621 ( .A1(n9440), .A2(n4579), .ZN(n4578) );
  NAND2_X1 U5622 ( .A1(n4582), .A2(n9403), .ZN(n4579) );
  AND2_X1 U5623 ( .A1(n4580), .A2(n4577), .ZN(n4576) );
  NAND2_X1 U5624 ( .A1(n9428), .A2(n9390), .ZN(n4586) );
  AND2_X1 U5625 ( .A1(n5620), .A2(n5619), .ZN(n9242) );
  INV_X1 U5626 ( .A(n6332), .ZN(n9443) );
  AND2_X1 U5627 ( .A1(n9385), .A2(n5660), .ZN(n8105) );
  AOI21_X1 U5628 ( .B1(n9480), .B2(n9479), .A(n4800), .ZN(n8104) );
  INV_X1 U5629 ( .A(n8103), .ZN(n4800) );
  AND2_X1 U5630 ( .A1(n5726), .A2(n8103), .ZN(n9479) );
  NOR2_X1 U5631 ( .A1(n9522), .A2(n9514), .ZN(n9513) );
  NAND2_X1 U5632 ( .A1(n9513), .A2(n9693), .ZN(n9494) );
  NAND2_X1 U5633 ( .A1(n9506), .A2(n8099), .ZN(n9493) );
  AND3_X1 U5634 ( .A1(n5528), .A2(n5527), .A3(n5526), .ZN(n9531) );
  OAI211_X1 U5635 ( .C1(n4783), .C2(n4780), .A(n9539), .B(n4781), .ZN(n5786)
         );
  NAND2_X1 U5636 ( .A1(n4782), .A2(n4784), .ZN(n4781) );
  NAND2_X1 U5637 ( .A1(n4607), .A2(n9525), .ZN(n9522) );
  AND2_X1 U5638 ( .A1(n5781), .A2(n5782), .ZN(n9565) );
  NAND2_X1 U5639 ( .A1(n9624), .A2(n4604), .ZN(n9604) );
  NAND2_X1 U5640 ( .A1(n9624), .A2(n9631), .ZN(n9625) );
  AOI21_X1 U5641 ( .B1(n8024), .B2(n8023), .A(n8022), .ZN(n9886) );
  NAND2_X1 U5642 ( .A1(n5772), .A2(n5771), .ZN(n7687) );
  NAND2_X1 U5643 ( .A1(n4794), .A2(n4793), .ZN(n7724) );
  INV_X1 U5644 ( .A(n7690), .ZN(n4793) );
  INV_X1 U5645 ( .A(n7687), .ZN(n4794) );
  NAND2_X1 U5646 ( .A1(n7691), .A2(n7690), .ZN(n7722) );
  NAND2_X1 U5647 ( .A1(n7632), .A2(n7631), .ZN(n7689) );
  NAND2_X1 U5648 ( .A1(n4590), .A2(n7437), .ZN(n7645) );
  AND4_X1 U5649 ( .A1(n5363), .A2(n5362), .A3(n5361), .A4(n5360), .ZN(n9174)
         );
  NAND2_X1 U5650 ( .A1(n7437), .A2(n9927), .ZN(n7517) );
  AND4_X1 U5651 ( .A1(n5342), .A2(n5341), .A3(n5340), .A4(n5339), .ZN(n7940)
         );
  NAND2_X1 U5652 ( .A1(n7433), .A2(n7435), .ZN(n7432) );
  NAND2_X1 U5653 ( .A1(n4449), .A2(n5737), .ZN(n7434) );
  NAND2_X1 U5654 ( .A1(n4563), .A2(n5736), .ZN(n4449) );
  NAND2_X1 U5655 ( .A1(n5737), .A2(n5736), .ZN(n7333) );
  NAND2_X1 U5656 ( .A1(n6887), .A2(n6886), .ZN(n9620) );
  NOR2_X1 U5657 ( .A1(n6330), .A2(n7270), .ZN(n7305) );
  NAND2_X1 U5658 ( .A1(n5269), .A2(n7153), .ZN(n4468) );
  INV_X1 U5659 ( .A(n5268), .ZN(n4465) );
  AND2_X1 U5660 ( .A1(n5634), .A2(n5633), .ZN(n9658) );
  OR2_X1 U5661 ( .A1(n9419), .A2(n5628), .ZN(n5634) );
  AND2_X1 U5662 ( .A1(n6891), .A2(n6890), .ZN(n9962) );
  OR2_X1 U5663 ( .A1(n6889), .A2(n6888), .ZN(n9914) );
  AND2_X1 U5664 ( .A1(n7259), .A2(n6352), .ZN(n6356) );
  NAND2_X1 U5665 ( .A1(n6815), .A2(n7262), .ZN(n9947) );
  INV_X1 U5666 ( .A(n9947), .ZN(n9959) );
  MUX2_X1 U5667 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5114), .S(
        P1_IR_REG_28__SCAN_IN), .Z(n5115) );
  INV_X1 U5668 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5107) );
  INV_X1 U5669 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5800) );
  INV_X1 U5670 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5801) );
  XNOR2_X1 U5671 ( .A(n5798), .B(n5797), .ZN(n6808) );
  NAND2_X1 U5672 ( .A1(n4396), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5798) );
  XNOR2_X1 U5673 ( .A(n5206), .B(n5205), .ZN(n7236) );
  AOI21_X1 U5674 ( .B1(n4319), .B2(n4879), .A(n4376), .ZN(n4874) );
  INV_X1 U5675 ( .A(n4985), .ZN(n4790) );
  INV_X1 U5676 ( .A(n5295), .ZN(n4436) );
  INV_X1 U5677 ( .A(n5275), .ZN(n4969) );
  NAND2_X1 U5678 ( .A1(n7027), .A2(n6006), .ZN(n7209) );
  AOI21_X1 U5679 ( .B1(n8767), .B2(n6111), .A(n6184), .ZN(n8774) );
  INV_X1 U5680 ( .A(n8485), .ZN(n4506) );
  NAND2_X1 U5681 ( .A1(n4950), .A2(n8536), .ZN(n8485) );
  NAND2_X1 U5682 ( .A1(n7208), .A2(n4490), .ZN(n4484) );
  AND3_X1 U5683 ( .A1(n6138), .A2(n6137), .A3(n6136), .ZN(n8802) );
  AND4_X1 U5684 ( .A1(n5912), .A2(n5911), .A3(n5910), .A4(n5909), .ZN(n7887)
         );
  NAND2_X1 U5685 ( .A1(n4910), .A2(n4909), .ZN(n7881) );
  INV_X1 U5686 ( .A(n4912), .ZN(n4909) );
  NAND2_X1 U5687 ( .A1(n8590), .A2(n4933), .ZN(n8520) );
  NAND2_X1 U5688 ( .A1(n6849), .A2(n5978), .ZN(n6953) );
  AND2_X1 U5689 ( .A1(n4932), .A2(n4931), .ZN(n8529) );
  AND2_X1 U5690 ( .A1(n5966), .A2(n4339), .ZN(n4929) );
  NAND2_X1 U5691 ( .A1(n4921), .A2(n4923), .ZN(n8500) );
  NAND2_X1 U5692 ( .A1(n8493), .A2(n4925), .ZN(n4921) );
  NAND2_X1 U5693 ( .A1(n4922), .A2(n4927), .ZN(n8548) );
  NAND2_X1 U5694 ( .A1(n8493), .A2(n4928), .ZN(n4922) );
  NOR2_X1 U5695 ( .A1(n4482), .A2(n7605), .ZN(n7841) );
  AOI21_X1 U5696 ( .B1(n4481), .B2(n4489), .A(n4480), .ZN(n4482) );
  INV_X1 U5697 ( .A(n4485), .ZN(n4480) );
  AOI21_X1 U5698 ( .B1(n4489), .B2(n4487), .A(n4486), .ZN(n4485) );
  INV_X1 U5699 ( .A(n4910), .ZN(n7839) );
  NAND2_X1 U5700 ( .A1(n6275), .A2(n7062), .ZN(n8595) );
  NAND2_X1 U5701 ( .A1(n6108), .A2(n8528), .ZN(n8566) );
  NAND2_X1 U5702 ( .A1(n4496), .A2(n4494), .ZN(n7027) );
  AND3_X1 U5703 ( .A1(n4495), .A2(n4375), .A3(n7028), .ZN(n4494) );
  AND2_X1 U5704 ( .A1(n4496), .A2(n4497), .ZN(n7029) );
  AND2_X1 U5705 ( .A1(n6222), .A2(n6221), .ZN(n8583) );
  INV_X1 U5706 ( .A(n8602), .ZN(n8585) );
  AOI22_X1 U5707 ( .A1(n8040), .A2(n8041), .B1(n6089), .B2(n8596), .ZN(n8592)
         );
  NAND2_X1 U5708 ( .A1(n8592), .A2(n8591), .ZN(n8590) );
  NAND2_X1 U5709 ( .A1(n6250), .A2(n6249), .ZN(n8589) );
  NAND2_X1 U5710 ( .A1(n6580), .A2(n6379), .ZN(n8458) );
  XNOR2_X1 U5711 ( .A(n6245), .B(P2_IR_REG_22__SCAN_IN), .ZN(n8459) );
  INV_X1 U5712 ( .A(n6243), .ZN(n6244) );
  INV_X1 U5713 ( .A(n8583), .ZN(n8742) );
  INV_X1 U5714 ( .A(n8576), .ZN(n8753) );
  INV_X1 U5715 ( .A(n8765), .ZN(n8741) );
  INV_X1 U5716 ( .A(n8802), .ZN(n8826) );
  INV_X1 U5717 ( .A(n8852), .ZN(n8825) );
  INV_X1 U5718 ( .A(n8864), .ZN(n8839) );
  INV_X1 U5719 ( .A(n7887), .ZN(n8613) );
  INV_X1 U5720 ( .A(n7315), .ZN(n8621) );
  NAND2_X1 U5721 ( .A1(n6264), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n5925) );
  OR2_X1 U5722 ( .A1(n6580), .A2(n6329), .ZN(n8623) );
  OR2_X1 U5723 ( .A1(n8412), .A2(n5927), .ZN(n5931) );
  NAND2_X1 U5724 ( .A1(n6725), .A2(n4750), .ZN(n6628) );
  XNOR2_X1 U5725 ( .A(n7176), .B(n7177), .ZN(n7105) );
  NOR2_X1 U5726 ( .A1(n7667), .A2(n7105), .ZN(n7178) );
  XNOR2_X1 U5727 ( .A(n7490), .B(n7483), .ZN(n7277) );
  NOR2_X1 U5728 ( .A1(n7277), .A2(n7278), .ZN(n7493) );
  NOR2_X1 U5729 ( .A1(n10024), .A2(n8643), .ZN(n10028) );
  AND2_X1 U5730 ( .A1(n6747), .A2(n6590), .ZN(n10058) );
  AND2_X1 U5731 ( .A1(n6118), .A2(n6117), .ZN(n8688) );
  INV_X1 U5732 ( .A(n8709), .ZN(n4772) );
  NAND2_X1 U5733 ( .A1(n4631), .A2(n8418), .ZN(n8768) );
  NAND2_X1 U5734 ( .A1(n4633), .A2(n8348), .ZN(n8818) );
  NAND2_X1 U5735 ( .A1(n6068), .A2(n6067), .ZN(n8312) );
  NAND2_X1 U5736 ( .A1(n6600), .A2(n8404), .ZN(n4535) );
  NAND2_X1 U5737 ( .A1(n4723), .A2(n4725), .ZN(n7657) );
  INV_X1 U5738 ( .A(n6853), .ZN(n7382) );
  NAND2_X1 U5739 ( .A1(n4637), .A2(n8277), .ZN(n7376) );
  AND2_X1 U5740 ( .A1(n10091), .A2(n7246), .ZN(n8819) );
  NAND2_X1 U5741 ( .A1(n4634), .A2(n8265), .ZN(n7160) );
  INV_X1 U5742 ( .A(n4635), .ZN(n4634) );
  INV_X1 U5743 ( .A(n8779), .ZN(n10085) );
  INV_X1 U5744 ( .A(n8813), .ZN(n10087) );
  AND2_X1 U5745 ( .A1(n8379), .A2(n8378), .ZN(n8876) );
  INV_X1 U5746 ( .A(n8979), .ZN(n8910) );
  NAND2_X1 U5747 ( .A1(n6215), .A2(n6214), .ZN(n8944) );
  NAND2_X1 U5748 ( .A1(n4611), .A2(n8367), .ZN(n8729) );
  NAND2_X1 U5749 ( .A1(n8221), .A2(n4615), .ZN(n4611) );
  NAND2_X1 U5750 ( .A1(n6202), .A2(n6201), .ZN(n8950) );
  NAND2_X1 U5751 ( .A1(n8221), .A2(n8220), .ZN(n8738) );
  INV_X1 U5752 ( .A(n8201), .ZN(n8955) );
  NAND2_X1 U5753 ( .A1(n6178), .A2(n6177), .ZN(n8962) );
  INV_X1 U5754 ( .A(n8489), .ZN(n8970) );
  NAND2_X1 U5755 ( .A1(n6156), .A2(n6155), .ZN(n8973) );
  NAND2_X1 U5756 ( .A1(n4713), .A2(n4717), .ZN(n8785) );
  NAND2_X1 U5757 ( .A1(n4716), .A2(n4720), .ZN(n8787) );
  NOR2_X1 U5758 ( .A1(n8195), .A2(n4748), .ZN(n8861) );
  NAND2_X1 U5759 ( .A1(n6080), .A2(n6079), .ZN(n8047) );
  NAND2_X1 U5760 ( .A1(n4627), .A2(n8302), .ZN(n7759) );
  NAND2_X1 U5761 ( .A1(n5917), .A2(n5916), .ZN(n7844) );
  INV_X2 U5762 ( .A(n10144), .ZN(n10142) );
  AND2_X1 U5763 ( .A1(n6579), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6379) );
  INV_X1 U5764 ( .A(n6239), .ZN(n8067) );
  XNOR2_X1 U5765 ( .A(n5847), .B(n5846), .ZN(n8039) );
  INV_X1 U5766 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n5846) );
  NAND2_X1 U5767 ( .A1(n5845), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5847) );
  INV_X1 U5768 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7801) );
  INV_X1 U5769 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7703) );
  INV_X1 U5770 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7473) );
  INV_X1 U5771 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n7386) );
  INV_X1 U5772 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n7295) );
  INV_X1 U5773 ( .A(n10002), .ZN(n8641) );
  INV_X1 U5774 ( .A(n7488), .ZN(n8637) );
  INV_X1 U5775 ( .A(n7492), .ZN(n7483) );
  INV_X1 U5776 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6605) );
  NAND2_X1 U5777 ( .A1(n4850), .A2(n9058), .ZN(n4849) );
  INV_X1 U5778 ( .A(n4852), .ZN(n4850) );
  AND2_X1 U5779 ( .A1(n9051), .A2(n9050), .ZN(n9121) );
  NAND2_X1 U5780 ( .A1(n5625), .A2(n5624), .ZN(n9401) );
  NAND2_X1 U5781 ( .A1(n4424), .A2(n4422), .ZN(n9126) );
  NOR2_X1 U5782 ( .A1(n9122), .A2(n4423), .ZN(n4422) );
  INV_X1 U5783 ( .A(n9116), .ZN(n4424) );
  OR2_X1 U5784 ( .A1(n9121), .A2(n9259), .ZN(n4423) );
  NAND2_X1 U5785 ( .A1(n4818), .A2(n4821), .ZN(n9129) );
  OR2_X1 U5786 ( .A1(n9104), .A2(n4822), .ZN(n4818) );
  OAI211_X1 U5787 ( .C1(n5308), .C2(n6370), .A(n5332), .B(n5331), .ZN(n9900)
         );
  NOR2_X1 U5788 ( .A1(n4846), .A2(n8142), .ZN(n9161) );
  INV_X1 U5789 ( .A(n4848), .ZN(n4846) );
  INV_X1 U5790 ( .A(n7131), .ZN(n4811) );
  OAI211_X1 U5791 ( .C1(n5308), .C2(n6367), .A(n5307), .B(n5306), .ZN(n7339)
         );
  INV_X1 U5792 ( .A(n7270), .ZN(n7150) );
  NAND2_X1 U5793 ( .A1(n4824), .A2(n8154), .ZN(n9127) );
  OR2_X1 U5794 ( .A1(n9104), .A2(n8155), .ZN(n4824) );
  AND4_X1 U5795 ( .A1(n5416), .A2(n5415), .A3(n5414), .A4(n5413), .ZN(n9953)
         );
  INV_X1 U5796 ( .A(n9201), .ZN(n4803) );
  INV_X1 U5797 ( .A(n9200), .ZN(n4804) );
  INV_X1 U5798 ( .A(n9693), .ZN(n9499) );
  AND4_X1 U5799 ( .A1(n5400), .A2(n5399), .A3(n5398), .A4(n5397), .ZN(n9219)
         );
  OAI211_X1 U5800 ( .C1(n5308), .C2(n6372), .A(n5246), .B(n5245), .ZN(n7600)
         );
  AND2_X1 U5801 ( .A1(n5626), .A2(n5601), .ZN(n9445) );
  NAND2_X1 U5802 ( .A1(n6813), .A2(n6812), .ZN(n9252) );
  INV_X1 U5803 ( .A(n9237), .ZN(n9259) );
  INV_X1 U5804 ( .A(n9601), .ZN(n9955) );
  NAND2_X1 U5805 ( .A1(n6832), .A2(n9532), .ZN(n9257) );
  NAND2_X1 U5806 ( .A1(n4458), .A2(n5793), .ZN(n4457) );
  AOI21_X1 U5807 ( .B1(n5795), .B2(n5796), .A(n5794), .ZN(n4460) );
  INV_X1 U5808 ( .A(n9658), .ZN(n9434) );
  NAND2_X1 U5809 ( .A1(n5595), .A2(n5594), .ZN(n9665) );
  OR2_X1 U5810 ( .A1(n9455), .A2(n5628), .ZN(n5595) );
  AND2_X1 U5811 ( .A1(n5550), .A2(n5549), .ZN(n9680) );
  INV_X1 U5812 ( .A(n9953), .ZN(n9264) );
  NAND2_X1 U5813 ( .A1(n5314), .A2(n4949), .ZN(n9271) );
  CLKBUF_X1 U5814 ( .A(n6835), .Z(n9274) );
  INV_X1 U5815 ( .A(n4545), .ZN(n9288) );
  INV_X1 U5816 ( .A(n4543), .ZN(n6946) );
  INV_X1 U5817 ( .A(n4541), .ZN(n9302) );
  INV_X1 U5818 ( .A(n4539), .ZN(n9316) );
  NAND2_X1 U5819 ( .A1(n9375), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n4559) );
  INV_X1 U5820 ( .A(n9374), .ZN(n4558) );
  OAI21_X1 U5821 ( .B1(n9370), .B2(n9857), .A(n4355), .ZN(n4562) );
  OAI22_X1 U5822 ( .A1(n9372), .A2(n9857), .B1(n9371), .B2(n9861), .ZN(n4560)
         );
  INV_X1 U5823 ( .A(n9401), .ZN(n9651) );
  INV_X1 U5824 ( .A(n4685), .ZN(n9414) );
  NAND2_X1 U5825 ( .A1(n4682), .A2(n4679), .ZN(n9429) );
  INV_X1 U5826 ( .A(n4680), .ZN(n4679) );
  NAND2_X1 U5827 ( .A1(n9440), .A2(n9389), .ZN(n9427) );
  INV_X1 U5828 ( .A(n9242), .ZN(n9666) );
  AOI21_X1 U5829 ( .B1(n9465), .B2(n9876), .A(n9464), .ZN(n9675) );
  INV_X1 U5830 ( .A(n9681), .ZN(n9486) );
  NAND2_X1 U5831 ( .A1(n5565), .A2(n5564), .ZN(n9690) );
  NAND2_X1 U5832 ( .A1(n4666), .A2(n4670), .ZN(n9492) );
  NAND2_X1 U5833 ( .A1(n8092), .A2(n4671), .ZN(n4666) );
  OAI21_X1 U5834 ( .B1(n8092), .B2(n4673), .A(n4948), .ZN(n9504) );
  OAI21_X1 U5835 ( .B1(n5783), .B2(n4784), .A(n4782), .ZN(n9538) );
  NAND2_X1 U5836 ( .A1(n4644), .A2(n4648), .ZN(n9537) );
  NAND2_X1 U5837 ( .A1(n9566), .A2(n4649), .ZN(n4644) );
  NOR2_X1 U5838 ( .A1(n4315), .A2(n9962), .ZN(n9549) );
  NAND2_X1 U5839 ( .A1(n5783), .A2(n5782), .ZN(n9551) );
  INV_X1 U5840 ( .A(n8089), .ZN(n4650) );
  NAND2_X1 U5841 ( .A1(n9566), .A2(n8090), .ZN(n4651) );
  AND4_X1 U5842 ( .A1(n5221), .A2(n5220), .A3(n5219), .A4(n5218), .ZN(n9571)
         );
  NAND2_X1 U5843 ( .A1(n9599), .A2(n5779), .ZN(n9589) );
  OAI21_X1 U5844 ( .B1(n4792), .B2(n4571), .A(n4317), .ZN(n9588) );
  NAND2_X1 U5845 ( .A1(n4654), .A2(n4655), .ZN(n9595) );
  AND2_X1 U5846 ( .A1(n4663), .A2(n4662), .ZN(n9619) );
  NAND2_X1 U5847 ( .A1(n5410), .A2(n5409), .ZN(n9890) );
  AND4_X1 U5848 ( .A1(n5382), .A2(n5381), .A3(n5380), .A4(n5379), .ZN(n9092)
         );
  NAND2_X1 U5849 ( .A1(n7261), .A2(n9532), .ZN(n9611) );
  NAND2_X1 U5850 ( .A1(n7512), .A2(n7511), .ZN(n7627) );
  NAND2_X1 U5851 ( .A1(n7510), .A2(n7509), .ZN(n7512) );
  INV_X1 U5852 ( .A(n9907), .ZN(n9894) );
  OR2_X1 U5853 ( .A1(n4315), .A2(n7269), .ZN(n9630) );
  NAND4_X1 U5854 ( .A1(n5265), .A2(n5264), .A3(n5263), .A4(n5262), .ZN(n7455)
         );
  INV_X1 U5855 ( .A(n9630), .ZN(n9901) );
  NAND2_X1 U5856 ( .A1(n9983), .A2(n9959), .ZN(n9747) );
  INV_X2 U5857 ( .A(n9981), .ZN(n9983) );
  NOR2_X1 U5858 ( .A1(n9644), .A2(n4796), .ZN(n9646) );
  NAND2_X1 U5859 ( .A1(n4798), .A2(n4797), .ZN(n4796) );
  NAND2_X1 U5860 ( .A1(n5587), .A2(n5586), .ZN(n9762) );
  INV_X1 U5861 ( .A(n9541), .ZN(n9775) );
  INV_X1 U5862 ( .A(n9606), .ZN(n9789) );
  INV_X1 U5863 ( .A(n9900), .ZN(n7444) );
  XNOR2_X1 U5864 ( .A(n5122), .B(n5121), .ZN(n5129) );
  NAND2_X1 U5865 ( .A1(n5127), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5122) );
  NAND2_X1 U5866 ( .A1(n5128), .A2(n5127), .ZN(n8076) );
  NAND2_X1 U5867 ( .A1(n5126), .A2(n5125), .ZN(n5128) );
  NAND2_X1 U5868 ( .A1(n4883), .A2(n4888), .ZN(n5552) );
  INV_X1 U5869 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7804) );
  INV_X1 U5870 ( .A(n6884), .ZN(n7802) );
  INV_X1 U5871 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7701) );
  INV_X1 U5872 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n8472) );
  INV_X1 U5873 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n7425) );
  INV_X1 U5874 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n7294) );
  AND2_X1 U5875 ( .A1(n5465), .A2(n5464), .ZN(n9837) );
  OR2_X1 U5876 ( .A1(n5445), .A2(n5444), .ZN(n5446) );
  NAND2_X1 U5877 ( .A1(n4881), .A2(n4880), .ZN(n5385) );
  AND2_X1 U5878 ( .A1(n5390), .A2(n5419), .ZN(n9809) );
  NAND2_X1 U5879 ( .A1(n5346), .A2(n4995), .ZN(n4802) );
  AOI22_X1 U5880 ( .A1(n4374), .A2(n9799), .B1(n4553), .B2(n9793), .ZN(n4552)
         );
  INV_X1 U5881 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n4553) );
  OR2_X1 U5882 ( .A1(n4966), .A2(n4965), .ZN(n4564) );
  NAND2_X1 U5883 ( .A1(n4967), .A2(n4963), .ZN(n5257) );
  CLKBUF_X1 U5884 ( .A(P1_IR_REG_0__SCAN_IN), .Z(n9799) );
  NAND2_X1 U5885 ( .A1(n4414), .A2(n4354), .ZN(P2_U3201) );
  NAND2_X1 U5886 ( .A1(n4771), .A2(n10026), .ZN(n4414) );
  XNOR2_X1 U5887 ( .A(n4773), .B(n4772), .ZN(n4771) );
  NAND2_X1 U5888 ( .A1(n10156), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n8884) );
  MUX2_X1 U5889 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n8938), .S(n10142), .Z(n8939) );
  INV_X1 U5890 ( .A(n6316), .ZN(n6317) );
  NAND2_X1 U5891 ( .A1(n4561), .A2(n4556), .ZN(P1_U3262) );
  AOI21_X1 U5892 ( .B1(n4560), .B2(n9373), .A(n4557), .ZN(n4556) );
  NAND2_X1 U5893 ( .A1(n4562), .A2(n7268), .ZN(n4561) );
  NAND2_X1 U5894 ( .A1(n4559), .A2(n4558), .ZN(n4557) );
  NAND2_X1 U5895 ( .A1(n4596), .A2(n4330), .ZN(n9754) );
  NAND2_X1 U5896 ( .A1(n9638), .A2(n4597), .ZN(n4596) );
  AND2_X1 U5897 ( .A1(n9590), .A2(n4570), .ZN(n4317) );
  INV_X1 U5898 ( .A(n5284), .ZN(n5396) );
  NOR2_X1 U5899 ( .A1(n8203), .A2(n8576), .ZN(n4318) );
  AND2_X1 U5900 ( .A1(n4876), .A2(n4875), .ZN(n4319) );
  NAND2_X1 U5901 ( .A1(n5148), .A2(n5653), .ZN(n4320) );
  INV_X2 U5902 ( .A(n4601), .ZN(n5644) );
  INV_X2 U5903 ( .A(n4601), .ZN(n5293) );
  AND2_X1 U5904 ( .A1(n4506), .A2(n8561), .ZN(n4321) );
  OR2_X1 U5905 ( .A1(n8160), .A2(n9128), .ZN(n4322) );
  AOI21_X1 U5906 ( .B1(n8401), .B2(n8404), .A(n8403), .ZN(n8932) );
  INV_X1 U5907 ( .A(n8932), .ZN(n4523) );
  NAND2_X1 U5908 ( .A1(n4586), .A2(n4584), .ZN(n4583) );
  INV_X1 U5909 ( .A(n5779), .ZN(n4571) );
  OR2_X1 U5910 ( .A1(n9560), .A2(n9727), .ZN(n4323) );
  NAND4_X1 U5911 ( .A1(n5819), .A2(n5946), .A3(n5817), .A4(n4366), .ZN(n4324)
         );
  AND2_X1 U5912 ( .A1(n4490), .A2(n8614), .ZN(n4325) );
  AND2_X1 U5913 ( .A1(n4491), .A2(n7838), .ZN(n4489) );
  XOR2_X1 U5914 ( .A(n8699), .B(n8698), .Z(n4326) );
  INV_X1 U5915 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n9793) );
  NAND2_X1 U5916 ( .A1(n4881), .A2(n4882), .ZN(n4327) );
  AND2_X1 U5917 ( .A1(n4604), .A2(n4603), .ZN(n4328) );
  NAND2_X2 U5918 ( .A1(n4956), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n4957) );
  NAND2_X1 U5919 ( .A1(n8343), .A2(n8344), .ZN(n8797) );
  INV_X1 U5920 ( .A(n8797), .ZN(n8444) );
  AND2_X1 U5921 ( .A1(n6022), .A2(n6006), .ZN(n4329) );
  NAND2_X1 U5922 ( .A1(n5860), .A2(n5862), .ZN(n8452) );
  INV_X1 U5923 ( .A(n8452), .ZN(n4501) );
  OR2_X1 U5924 ( .A1(n9968), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n4330) );
  OR2_X1 U5925 ( .A1(n6815), .A2(n6884), .ZN(n4331) );
  AND2_X1 U5926 ( .A1(n5946), .A2(n5817), .ZN(n5889) );
  OR2_X1 U5927 ( .A1(n4619), .A2(n4617), .ZN(n5860) );
  NAND2_X1 U5928 ( .A1(n5267), .A2(n6364), .ZN(n4601) );
  AND2_X1 U5929 ( .A1(n4804), .A2(n4803), .ZN(n4332) );
  NAND2_X1 U5930 ( .A1(n9401), .A2(n9434), .ZN(n4333) );
  INV_X1 U5931 ( .A(n9560), .ZN(n9779) );
  NAND2_X1 U5932 ( .A1(n4815), .A2(n5096), .ZN(n5294) );
  NOR2_X1 U5933 ( .A1(n6076), .A2(n8612), .ZN(n4334) );
  NAND2_X1 U5934 ( .A1(n5659), .A2(n5711), .ZN(n9403) );
  INV_X1 U5935 ( .A(n9403), .ZN(n4577) );
  AND2_X1 U5936 ( .A1(n6644), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n4335) );
  INV_X1 U5937 ( .A(n4944), .ZN(n4684) );
  NAND2_X1 U5938 ( .A1(n4665), .A2(n4664), .ZN(n9478) );
  AND2_X1 U5939 ( .A1(n4847), .A2(n9160), .ZN(n4336) );
  NAND2_X1 U5940 ( .A1(n8480), .A2(n8479), .ZN(n4337) );
  INV_X1 U5941 ( .A(n8560), .ZN(n8810) );
  INV_X1 U5942 ( .A(n9140), .ZN(n4855) );
  AND4_X1 U5943 ( .A1(n5734), .A2(n5582), .A3(n5749), .A4(n9873), .ZN(n4338)
         );
  INV_X1 U5944 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n5938) );
  INV_X1 U5945 ( .A(n9583), .ZN(n4603) );
  OR2_X1 U5946 ( .A1(n8226), .A2(n6676), .ZN(n4339) );
  NOR2_X1 U5947 ( .A1(n5295), .A2(n4816), .ZN(n5328) );
  NAND2_X1 U5948 ( .A1(n5178), .A2(n5177), .ZN(n9705) );
  AND3_X1 U5949 ( .A1(n8336), .A2(n4533), .A3(n4532), .ZN(n4340) );
  AND2_X1 U5950 ( .A1(n9560), .A2(n9727), .ZN(n4341) );
  AND2_X1 U5951 ( .A1(n4539), .A2(n4538), .ZN(n4342) );
  OR2_X1 U5952 ( .A1(n7658), .A2(n8616), .ZN(n4343) );
  AND2_X1 U5953 ( .A1(n4719), .A2(n8797), .ZN(n4344) );
  NAND2_X1 U5954 ( .A1(n8312), .A2(n8612), .ZN(n4345) );
  AND2_X1 U5955 ( .A1(n4725), .A2(n4343), .ZN(n4346) );
  OR2_X1 U5956 ( .A1(n5145), .A2(n4829), .ZN(n4347) );
  INV_X1 U5957 ( .A(n4861), .ZN(n5721) );
  NOR2_X1 U5958 ( .A1(n10028), .A2(n8644), .ZN(n4348) );
  AND2_X1 U5959 ( .A1(n8944), .A2(n8742), .ZN(n4349) );
  AND2_X1 U5960 ( .A1(n5580), .A2(n8105), .ZN(n4350) );
  AND2_X1 U5961 ( .A1(n8527), .A2(n4931), .ZN(n4351) );
  INV_X1 U5962 ( .A(n8321), .ZN(n8437) );
  AND2_X1 U5963 ( .A1(n4996), .A2(n4995), .ZN(n4352) );
  AND2_X1 U5964 ( .A1(n5822), .A2(n4739), .ZN(n4353) );
  AND2_X1 U5965 ( .A1(n8713), .A2(n4413), .ZN(n4354) );
  INV_X1 U5966 ( .A(n4588), .ZN(n4587) );
  NAND2_X1 U5967 ( .A1(n9390), .A2(n9389), .ZN(n4588) );
  INV_X1 U5968 ( .A(n4934), .ZN(n4933) );
  AND2_X1 U5969 ( .A1(n9369), .A2(n9851), .ZN(n4355) );
  AND2_X1 U5970 ( .A1(n9770), .A2(n9531), .ZN(n4356) );
  OR2_X1 U5971 ( .A1(n7503), .A2(n6889), .ZN(n4357) );
  AND2_X1 U5972 ( .A1(n9693), .A2(n9680), .ZN(n4358) );
  INV_X1 U5973 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5146) );
  NAND2_X1 U5974 ( .A1(n5261), .A2(n4552), .ZN(n6641) );
  NOR2_X1 U5975 ( .A1(n8162), .A2(n8161), .ZN(n4359) );
  NOR2_X1 U5976 ( .A1(n9775), .A2(n9530), .ZN(n4360) );
  OR2_X1 U5977 ( .A1(n8089), .A2(n4341), .ZN(n4361) );
  AND2_X1 U5978 ( .A1(n8199), .A2(n8801), .ZN(n4362) );
  INV_X1 U5979 ( .A(n5737), .ZN(n4448) );
  INV_X1 U5980 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n6553) );
  AND2_X1 U5981 ( .A1(n8205), .A2(n8583), .ZN(n4363) );
  NOR2_X1 U5982 ( .A1(n8979), .A2(n8810), .ZN(n4364) );
  AND2_X1 U5983 ( .A1(n7397), .A2(n7396), .ZN(n4365) );
  INV_X1 U5984 ( .A(n8365), .ZN(n8220) );
  AND2_X1 U5985 ( .A1(n8201), .A2(n8765), .ZN(n8365) );
  INV_X1 U5986 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n5797) );
  AND4_X1 U5987 ( .A1(n4708), .A2(n4709), .A3(n4707), .A4(n5857), .ZN(n4366)
         );
  AND2_X1 U5988 ( .A1(n4856), .A2(n4320), .ZN(n4367) );
  OR2_X1 U5989 ( .A1(n7991), .A2(n9170), .ZN(n4368) );
  NOR2_X1 U5990 ( .A1(n9693), .A2(n9680), .ZN(n4369) );
  NOR2_X1 U5991 ( .A1(n9661), .A2(n9666), .ZN(n4370) );
  AND2_X1 U5992 ( .A1(n4320), .A2(n7147), .ZN(n4371) );
  NAND2_X1 U5993 ( .A1(n7986), .A2(n7985), .ZN(n4372) );
  NAND2_X1 U5994 ( .A1(n7992), .A2(n4368), .ZN(n4373) );
  AND2_X1 U5995 ( .A1(n8246), .A2(n8244), .ZN(n8783) );
  AND2_X2 U5996 ( .A1(n9113), .A2(n9030), .ZN(n7129) );
  NAND2_X1 U5997 ( .A1(n5723), .A2(n9390), .ZN(n9428) );
  AND2_X1 U5998 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n4374) );
  INV_X1 U5999 ( .A(n4926), .ZN(n4925) );
  NAND2_X1 U6000 ( .A1(n8547), .A2(n4928), .ZN(n4926) );
  NAND2_X1 U6001 ( .A1(n5991), .A2(n7359), .ZN(n4375) );
  NOR2_X1 U6002 ( .A1(n5010), .A2(SI_11_), .ZN(n4376) );
  AND2_X1 U6003 ( .A1(n5436), .A2(n5435), .ZN(n4377) );
  NAND2_X1 U6004 ( .A1(n4942), .A2(n8154), .ZN(n4378) );
  NAND2_X1 U6005 ( .A1(n7927), .A2(n4838), .ZN(n4379) );
  INV_X1 U6006 ( .A(n4783), .ZN(n4782) );
  NAND2_X1 U6007 ( .A1(n4417), .A2(n5784), .ZN(n4783) );
  INV_X1 U6008 ( .A(n4583), .ZN(n4582) );
  AND2_X1 U6009 ( .A1(n7616), .A2(n7503), .ZN(n4380) );
  AND2_X1 U6010 ( .A1(n4651), .A2(n4650), .ZN(n4381) );
  AND2_X1 U6011 ( .A1(n8100), .A2(n8101), .ZN(n4382) );
  INV_X1 U6012 ( .A(n9381), .ZN(n4859) );
  NOR2_X1 U6013 ( .A1(n8567), .A2(n4512), .ZN(n4383) );
  AND2_X1 U6014 ( .A1(n5493), .A2(n5492), .ZN(n9783) );
  INV_X1 U6015 ( .A(n9783), .ZN(n4605) );
  AND2_X1 U6016 ( .A1(n4577), .A2(n4451), .ZN(n4384) );
  OR2_X1 U6017 ( .A1(n5145), .A2(P1_IR_REG_20__SCAN_IN), .ZN(n4385) );
  OR2_X1 U6018 ( .A1(n8913), .A2(n8802), .ZN(n8342) );
  INV_X1 U6019 ( .A(n4947), .ZN(n4813) );
  OR2_X1 U6020 ( .A1(n5335), .A2(n4448), .ZN(n4386) );
  INV_X1 U6021 ( .A(n5004), .ZN(n4882) );
  INV_X1 U6022 ( .A(n4880), .ZN(n4879) );
  INV_X1 U6023 ( .A(n5375), .ZN(n5631) );
  INV_X1 U6024 ( .A(n7838), .ZN(n8614) );
  INV_X1 U6025 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n4516) );
  NAND2_X1 U6026 ( .A1(n8590), .A2(n4930), .ZN(n4932) );
  INV_X1 U6027 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n4428) );
  AND2_X1 U6028 ( .A1(n9624), .A2(n4328), .ZN(n4387) );
  INV_X1 U6029 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n4430) );
  INV_X1 U6030 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n4776) );
  AND2_X1 U6031 ( .A1(n6696), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n4388) );
  NAND2_X1 U6032 ( .A1(n5612), .A2(n5611), .ZN(n9661) );
  INV_X1 U6033 ( .A(n9661), .ZN(n4606) );
  NAND2_X1 U6034 ( .A1(n5889), .A2(n5819), .ZN(n5856) );
  NOR2_X1 U6035 ( .A1(n7494), .A2(n7493), .ZN(n4389) );
  NOR2_X1 U6036 ( .A1(n9994), .A2(n8639), .ZN(n4390) );
  INV_X1 U6037 ( .A(n8142), .ZN(n4847) );
  AND2_X1 U6038 ( .A1(n5017), .A2(n4903), .ZN(n4391) );
  INV_X1 U6039 ( .A(n4607), .ZN(n9540) );
  INV_X1 U6040 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n5832) );
  NAND2_X1 U6041 ( .A1(n5736), .A2(n5767), .ZN(n4392) );
  INV_X1 U6042 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n4708) );
  NAND2_X1 U6043 ( .A1(n5026), .A2(n5487), .ZN(n4393) );
  AND4_X1 U6044 ( .A1(n6057), .A2(n6056), .A3(n6055), .A4(n6054), .ZN(n7838)
         );
  NOR2_X1 U6045 ( .A1(n4902), .A2(n4900), .ZN(n4394) );
  AND2_X1 U6046 ( .A1(n5857), .A2(n4708), .ZN(n4395) );
  NAND2_X1 U6047 ( .A1(n7268), .A2(n7802), .ZN(n6889) );
  AND2_X1 U6048 ( .A1(n7208), .A2(n6024), .ZN(n6318) );
  INV_X1 U6049 ( .A(n4812), .ZN(n7132) );
  AND2_X1 U6050 ( .A1(n8468), .A2(n5872), .ZN(n6193) );
  INV_X2 U6051 ( .A(n9966), .ZN(n9968) );
  NAND2_X1 U6052 ( .A1(n6818), .A2(n7526), .ZN(n6815) );
  AND2_X1 U6053 ( .A1(n6176), .A2(n6175), .ZN(n8561) );
  AOI21_X1 U6054 ( .B1(n5855), .B2(n5854), .A(n6378), .ZN(n6223) );
  XNOR2_X1 U6055 ( .A(n4808), .B(n5800), .ZN(n6336) );
  OR2_X1 U6056 ( .A1(n5145), .A2(n4826), .ZN(n4396) );
  NAND2_X1 U6057 ( .A1(n4907), .A2(n7883), .ZN(n4912) );
  NOR2_X1 U6058 ( .A1(n7006), .A2(n7005), .ZN(n4397) );
  AND2_X1 U6059 ( .A1(n9809), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n4398) );
  NAND2_X1 U6060 ( .A1(n9927), .A2(n7743), .ZN(n4594) );
  INV_X1 U6061 ( .A(n4594), .ZN(n4590) );
  AND2_X1 U6062 ( .A1(n4484), .A2(n4489), .ZN(n4399) );
  NAND2_X1 U6063 ( .A1(n4812), .A2(n4811), .ZN(n4400) );
  AND2_X1 U6064 ( .A1(n4468), .A2(n4465), .ZN(n4401) );
  NAND2_X1 U6065 ( .A1(n4801), .A2(n5356), .ZN(n7938) );
  INV_X1 U6066 ( .A(n7938), .ZN(n4593) );
  NAND2_X1 U6067 ( .A1(n4501), .A2(n8453), .ZN(n4500) );
  OR2_X1 U6068 ( .A1(n10033), .A2(n8926), .ZN(n4402) );
  NAND2_X1 U6069 ( .A1(n4635), .A2(n8265), .ZN(n7240) );
  INV_X1 U6070 ( .A(n7220), .ZN(n7225) );
  OR2_X1 U6071 ( .A1(n9393), .A2(n9392), .ZN(n4403) );
  OR2_X1 U6072 ( .A1(n8712), .A2(n8711), .ZN(n4404) );
  INV_X1 U6073 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n4550) );
  INV_X1 U6074 ( .A(n7526), .ZN(n6888) );
  INV_X1 U6075 ( .A(n4602), .ZN(n6362) );
  NAND2_X1 U6076 ( .A1(n5258), .A2(n4565), .ZN(n4602) );
  INV_X1 U6077 ( .A(n6818), .ZN(n7268) );
  INV_X1 U6078 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n4412) );
  INV_X1 U6079 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n4600) );
  INV_X1 U6080 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n4547) );
  NAND2_X2 U6081 ( .A1(n6363), .A2(P2_U3151), .ZN(n9015) );
  OAI21_X2 U6082 ( .B1(n8848), .B2(n8216), .A(n8337), .ZN(n8832) );
  NAND2_X1 U6083 ( .A1(n5301), .A2(n5300), .ZN(n5303) );
  NAND2_X1 U6084 ( .A1(n7707), .A2(n7706), .ZN(n4627) );
  NAND2_X1 U6085 ( .A1(n7821), .A2(n8314), .ZN(n7847) );
  NAND2_X1 U6086 ( .A1(n4633), .A2(n4632), .ZN(n8795) );
  NAND2_X1 U6087 ( .A1(n8219), .A2(n8360), .ZN(n8749) );
  NAND2_X1 U6088 ( .A1(n8224), .A2(n8223), .ZN(n8480) );
  NAND2_X1 U6089 ( .A1(n8776), .A2(n8419), .ZN(n4631) );
  AND2_X1 U6090 ( .A1(n5982), .A2(n5981), .ZN(n4405) );
  NAND2_X1 U6091 ( .A1(n8822), .A2(n8823), .ZN(n4633) );
  NAND2_X1 U6092 ( .A1(n7656), .A2(n8430), .ZN(n7707) );
  INV_X1 U6093 ( .A(n8281), .ZN(n8273) );
  NAND2_X2 U6094 ( .A1(n5997), .A2(n5996), .ZN(n7393) );
  NAND2_X1 U6095 ( .A1(n9147), .A2(n8143), .ZN(n4848) );
  OAI21_X1 U6096 ( .B1(n7415), .B2(n7414), .A(n7589), .ZN(n7416) );
  OAI21_X2 U6097 ( .B1(n7021), .B2(n4810), .A(n4809), .ZN(n7414) );
  NAND2_X1 U6098 ( .A1(n7312), .A2(n7311), .ZN(n4637) );
  NAND2_X1 U6099 ( .A1(n4408), .A2(n4523), .ZN(n4522) );
  NAND2_X1 U6100 ( .A1(n8405), .A2(n8408), .ZN(n4408) );
  AOI21_X1 U6101 ( .B1(n8399), .B2(n8398), .A(n8397), .ZN(n8407) );
  OAI211_X1 U6102 ( .C1(n5850), .C2(n5836), .A(n5835), .B(n5834), .ZN(n5837)
         );
  INV_X1 U6103 ( .A(n4789), .ZN(n4788) );
  OAI21_X1 U6104 ( .B1(n4410), .B2(n4409), .A(n8417), .ZN(n4521) );
  NAND2_X1 U6105 ( .A1(n5289), .A2(n5290), .ZN(n5292) );
  NAND2_X1 U6106 ( .A1(n8102), .A2(n8101), .ZN(n9480) );
  NAND2_X1 U6107 ( .A1(n8104), .A2(n8105), .ZN(n9386) );
  NAND2_X1 U6108 ( .A1(n6363), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n4429) );
  OAI21_X1 U6109 ( .B1(n6363), .B2(n4430), .A(n4429), .ZN(n4971) );
  AOI21_X1 U6110 ( .B1(n4567), .B2(n8097), .A(n4566), .ZN(n9507) );
  INV_X1 U6111 ( .A(n8650), .ZN(n10060) );
  INV_X1 U6112 ( .A(n10062), .ZN(n4415) );
  NOR2_X1 U6113 ( .A1(n5937), .A2(n5826), .ZN(n4754) );
  OR2_X1 U6114 ( .A1(n6872), .A2(n6871), .ZN(n7015) );
  NAND2_X1 U6115 ( .A1(n4820), .A2(n4819), .ZN(n8165) );
  NAND2_X1 U6116 ( .A1(n4863), .A2(n4864), .ZN(n5039) );
  NAND2_X1 U6117 ( .A1(n4715), .A2(n4714), .ZN(n8772) );
  NAND2_X1 U6118 ( .A1(n4906), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n4905) );
  OAI211_X2 U6119 ( .C1(n8727), .C2(n8236), .A(n8235), .B(n8237), .ZN(n8720)
         );
  XNOR2_X1 U6120 ( .A(n7126), .B(n4416), .ZN(n7020) );
  XNOR2_X1 U6121 ( .A(n7019), .B(n9030), .ZN(n7126) );
  INV_X1 U6122 ( .A(n8165), .ZN(n4420) );
  NAND2_X1 U6123 ( .A1(n9507), .A2(n9508), .ZN(n9506) );
  NAND2_X1 U6124 ( .A1(n9139), .A2(n9140), .ZN(n9138) );
  INV_X1 U6125 ( .A(n9528), .ZN(n4567) );
  NAND2_X1 U6126 ( .A1(n9159), .A2(n4432), .ZN(n9225) );
  NAND2_X1 U6127 ( .A1(n4585), .A2(n4586), .ZN(n9416) );
  NAND2_X1 U6128 ( .A1(n8215), .A2(n8330), .ZN(n8848) );
  XNOR2_X1 U6129 ( .A(n4426), .B(n8711), .ZN(n8463) );
  NAND3_X1 U6130 ( .A1(n4521), .A2(n4522), .A3(n4952), .ZN(n4426) );
  NAND2_X1 U6131 ( .A1(n4610), .A2(n4608), .ZN(n8477) );
  NAND2_X1 U6132 ( .A1(n4457), .A2(n6888), .ZN(n4456) );
  INV_X1 U6133 ( .A(n5443), .ZN(n4473) );
  NAND2_X1 U6134 ( .A1(n5538), .A2(n6889), .ZN(n4478) );
  NAND2_X1 U6135 ( .A1(n4459), .A2(n5791), .ZN(n4458) );
  NAND2_X1 U6136 ( .A1(n4477), .A2(n4476), .ZN(n4475) );
  NAND2_X1 U6137 ( .A1(n5639), .A2(n4450), .ZN(n5641) );
  OAI21_X1 U6138 ( .B1(n5324), .B2(n4790), .A(n5240), .ZN(n4789) );
  AOI21_X1 U6139 ( .B1(n4788), .B2(n4790), .A(n4786), .ZN(n4785) );
  INV_X1 U6140 ( .A(n4744), .ZN(n4741) );
  NAND2_X1 U6141 ( .A1(n4741), .A2(n4746), .ZN(n4740) );
  NAND2_X1 U6142 ( .A1(n4807), .A2(n4805), .ZN(n8185) );
  INV_X2 U6143 ( .A(n5267), .ZN(n5305) );
  NAND3_X1 U6144 ( .A1(n5104), .A2(n4825), .A3(n4434), .ZN(n5109) );
  NAND4_X1 U6146 ( .A1(n5103), .A2(n5102), .A3(n5134), .A4(n6523), .ZN(n4437)
         );
  NAND4_X1 U6147 ( .A1(n5099), .A2(n5098), .A3(n5101), .A4(n5100), .ZN(n5137)
         );
  NAND2_X1 U6148 ( .A1(n7503), .A2(n5768), .ZN(n4438) );
  NAND2_X1 U6149 ( .A1(n7504), .A2(n4438), .ZN(n4444) );
  OAI21_X1 U6150 ( .B1(n4563), .B2(n4386), .A(n4439), .ZN(n4442) );
  NAND3_X1 U6151 ( .A1(n4443), .A2(n4442), .A3(n4357), .ZN(n5351) );
  NAND3_X1 U6152 ( .A1(n4446), .A2(n6889), .A3(n4444), .ZN(n4443) );
  NAND3_X1 U6153 ( .A1(n4455), .A2(n5722), .A3(n4454), .ZN(n4453) );
  NAND3_X1 U6154 ( .A1(n5621), .A2(n9390), .A3(n9389), .ZN(n4455) );
  INV_X1 U6155 ( .A(n5740), .ZN(n4467) );
  AOI21_X2 U6156 ( .B1(n4475), .B2(n4350), .A(n4474), .ZN(n5636) );
  NAND3_X1 U6157 ( .A1(n4479), .A2(n4478), .A3(n4382), .ZN(n4477) );
  INV_X1 U6158 ( .A(n7208), .ZN(n4481) );
  INV_X1 U6159 ( .A(n6049), .ZN(n4491) );
  AND2_X1 U6160 ( .A1(n4495), .A2(n4375), .ZN(n4497) );
  NAND2_X1 U6161 ( .A1(n4498), .A2(n6954), .ZN(n4495) );
  NAND3_X1 U6162 ( .A1(n6847), .A2(n5976), .A3(n6954), .ZN(n4496) );
  INV_X1 U6163 ( .A(n5978), .ZN(n4498) );
  NAND2_X1 U6164 ( .A1(n5976), .A2(n6847), .ZN(n6849) );
  NAND2_X2 U6165 ( .A1(n4502), .A2(n4499), .ZN(n5951) );
  INV_X1 U6166 ( .A(n4950), .ZN(n4503) );
  NAND2_X1 U6167 ( .A1(n4503), .A2(n8536), .ZN(n4505) );
  NAND2_X1 U6168 ( .A1(n4505), .A2(n4504), .ZN(n8539) );
  NAND2_X1 U6169 ( .A1(n6108), .A2(n4383), .ZN(n4511) );
  NAND2_X1 U6170 ( .A1(n4511), .A2(n4509), .ZN(n4508) );
  NAND2_X1 U6171 ( .A1(n4508), .A2(n4916), .ZN(n8499) );
  NAND2_X1 U6172 ( .A1(n5858), .A2(n4395), .ZN(n6117) );
  NAND2_X1 U6173 ( .A1(n4514), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6116) );
  NAND2_X1 U6174 ( .A1(n6096), .A2(n4514), .ZN(n8678) );
  INV_X8 U6175 ( .A(n4518), .ZN(n6363) );
  NAND2_X2 U6176 ( .A1(n4958), .A2(n4957), .ZN(n4518) );
  NAND2_X1 U6177 ( .A1(n4962), .A2(SI_1_), .ZN(n4967) );
  NAND4_X1 U6178 ( .A1(n8327), .A2(n8325), .A3(n8388), .A4(n8326), .ZN(n4532)
         );
  OAI21_X4 U6179 ( .B1(P1_ADDR_REG_19__SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(
        n4954), .ZN(n4958) );
  NAND2_X1 U6180 ( .A1(n4564), .A2(n5257), .ZN(n4565) );
  NAND2_X1 U6181 ( .A1(n9596), .A2(n5779), .ZN(n4570) );
  NAND2_X1 U6182 ( .A1(n9440), .A2(n4576), .ZN(n4575) );
  NAND2_X1 U6183 ( .A1(n9440), .A2(n4587), .ZN(n4585) );
  NAND3_X1 U6184 ( .A1(n4578), .A2(n4575), .A3(n4572), .ZN(n4799) );
  NAND2_X1 U6185 ( .A1(n7437), .A2(n4593), .ZN(n4592) );
  INV_X1 U6186 ( .A(n4592), .ZN(n4591) );
  AND3_X1 U6187 ( .A1(n4591), .A2(n9940), .A3(n4590), .ZN(n4589) );
  AND3_X2 U6188 ( .A1(n9783), .A2(n4328), .A3(n9624), .ZN(n9572) );
  NOR2_X2 U6189 ( .A1(n9417), .A2(n6333), .ZN(n9405) );
  AND2_X2 U6190 ( .A1(n6332), .A2(n4606), .ZN(n9430) );
  NOR2_X2 U6191 ( .A1(n9557), .A2(n9541), .ZN(n4607) );
  NAND2_X1 U6192 ( .A1(n8221), .A2(n4612), .ZN(n4610) );
  NAND2_X1 U6193 ( .A1(n4618), .A2(n5817), .ZN(n4616) );
  NOR2_X2 U6194 ( .A1(n4616), .A2(n4619), .ZN(n6243) );
  AND4_X2 U6195 ( .A1(n4701), .A2(n4620), .A3(n5819), .A4(n5817), .ZN(n5827)
         );
  NAND2_X1 U6196 ( .A1(n4627), .A2(n4624), .ZN(n7708) );
  NAND2_X1 U6197 ( .A1(n4631), .A2(n4628), .ZN(n8219) );
  OR2_X2 U6198 ( .A1(n8832), .A2(n8836), .ZN(n8833) );
  NAND2_X1 U6199 ( .A1(n7511), .A2(n4641), .ZN(n4639) );
  NAND2_X1 U6200 ( .A1(n7353), .A2(n7352), .ZN(n7510) );
  NAND2_X1 U6201 ( .A1(n4640), .A2(n4638), .ZN(n7640) );
  INV_X1 U6202 ( .A(n5109), .ZN(n5113) );
  NAND2_X1 U6203 ( .A1(n9566), .A2(n4645), .ZN(n4642) );
  NAND2_X1 U6204 ( .A1(n4642), .A2(n4643), .ZN(n9521) );
  INV_X1 U6205 ( .A(n4663), .ZN(n8086) );
  NAND2_X1 U6206 ( .A1(n8092), .A2(n4667), .ZN(n4665) );
  NAND2_X1 U6207 ( .A1(n4674), .A2(n4675), .ZN(n9404) );
  NAND2_X1 U6208 ( .A1(n9453), .A2(n4678), .ZN(n4674) );
  NAND2_X1 U6209 ( .A1(n9453), .A2(n4683), .ZN(n4682) );
  OR2_X1 U6210 ( .A1(n6375), .A2(n5964), .ZN(n6012) );
  OAI211_X2 U6211 ( .C1(n6597), .C2(n8226), .A(n5922), .B(n5921), .ZN(n7055)
         );
  NAND2_X1 U6212 ( .A1(n8480), .A2(n8225), .ZN(n8399) );
  AOI21_X1 U6213 ( .B1(n9789), .B2(n9736), .A(n8088), .ZN(n9582) );
  OAI21_X2 U6214 ( .B1(n9478), .B2(n8095), .A(n8094), .ZN(n9395) );
  NAND2_X1 U6215 ( .A1(n7640), .A2(n7639), .ZN(n7638) );
  NAND2_X1 U6216 ( .A1(n5113), .A2(n4939), .ZN(n5118) );
  NAND2_X1 U6217 ( .A1(n7222), .A2(n7223), .ZN(n7332) );
  OR2_X1 U6218 ( .A1(n9395), .A2(n9394), .ZN(n9397) );
  NAND2_X1 U6219 ( .A1(n7350), .A2(n7349), .ZN(n7433) );
  INV_X1 U6220 ( .A(n9521), .ZN(n8092) );
  XNOR2_X1 U6221 ( .A(n6835), .B(n8082), .ZN(n7145) );
  NAND2_X1 U6222 ( .A1(n7722), .A2(n7721), .ZN(n8024) );
  NAND2_X1 U6223 ( .A1(n7432), .A2(n7351), .ZN(n7353) );
  XNOR2_X1 U6224 ( .A(n5108), .B(n5107), .ZN(n5809) );
  NAND2_X1 U6225 ( .A1(n9580), .A2(n4941), .ZN(n9566) );
  NAND2_X1 U6226 ( .A1(n7334), .A2(n7333), .ZN(n7350) );
  NAND2_X1 U6227 ( .A1(n5327), .A2(n4985), .ZN(n5241) );
  NAND3_X1 U6228 ( .A1(n7363), .A2(n8420), .A3(n4698), .ZN(n4697) );
  NAND3_X1 U6229 ( .A1(n4708), .A2(n5857), .A3(n5938), .ZN(n4702) );
  NAND4_X1 U6230 ( .A1(n4707), .A2(n4709), .A3(n4712), .A4(n4711), .ZN(n4703)
         );
  AND4_X2 U6231 ( .A1(n5818), .A2(n4706), .A3(n4705), .A4(n4704), .ZN(n5819)
         );
  INV_X2 U6232 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n4712) );
  INV_X1 U6233 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n4710) );
  NAND2_X1 U6234 ( .A1(n8807), .A2(n4717), .ZN(n4715) );
  NAND2_X1 U6235 ( .A1(n8739), .A2(n4733), .ZN(n4729) );
  OAI21_X1 U6236 ( .B1(n8739), .B2(n4737), .A(n4735), .ZN(n8473) );
  NAND2_X1 U6237 ( .A1(n4729), .A2(n4730), .ZN(n8211) );
  AOI21_X1 U6238 ( .B1(n8739), .B2(n8204), .A(n4318), .ZN(n8731) );
  NAND2_X1 U6239 ( .A1(n5827), .A2(n5822), .ZN(n5824) );
  INV_X1 U6240 ( .A(n5867), .ZN(n5865) );
  NAND2_X1 U6241 ( .A1(n5867), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5868) );
  OAI21_X1 U6242 ( .B1(n7956), .B2(n4742), .A(n4740), .ZN(n8850) );
  INV_X1 U6243 ( .A(n4747), .ZN(n8860) );
  OAI21_X1 U6244 ( .B1(n10024), .B2(n4767), .A(n4766), .ZN(n10042) );
  NAND3_X1 U6245 ( .A1(n4404), .A2(n8710), .A3(n4770), .ZN(n4769) );
  NAND3_X1 U6246 ( .A1(n4958), .A2(n4957), .A3(P2_DATAO_REG_2__SCAN_IN), .ZN(
        n4774) );
  INV_X1 U6247 ( .A(n5783), .ZN(n4780) );
  OAI21_X1 U6248 ( .B1(n5325), .B2(n4790), .A(n4788), .ZN(n5243) );
  NAND2_X1 U6249 ( .A1(n4787), .A2(n4785), .ZN(n5344) );
  NAND2_X1 U6250 ( .A1(n5325), .A2(n4788), .ZN(n4787) );
  NAND2_X1 U6251 ( .A1(n9200), .A2(n9076), .ZN(n4807) );
  NAND2_X1 U6252 ( .A1(n8185), .A2(n8184), .ZN(n8187) );
  NAND2_X1 U6253 ( .A1(n7131), .A2(n4813), .ZN(n4809) );
  NAND2_X1 U6254 ( .A1(n9104), .A2(n4821), .ZN(n4820) );
  NAND2_X1 U6255 ( .A1(n7742), .A2(n4833), .ZN(n4831) );
  OAI21_X1 U6256 ( .B1(n7742), .B2(n7741), .A(n7740), .ZN(n7928) );
  NAND2_X1 U6257 ( .A1(n9147), .A2(n4841), .ZN(n4840) );
  NAND2_X1 U6258 ( .A1(n4848), .A2(n4336), .ZN(n9159) );
  NAND3_X1 U6259 ( .A1(n5658), .A2(n5657), .A3(n9381), .ZN(n4858) );
  NAND3_X1 U6260 ( .A1(n5203), .A2(n4865), .A3(n5202), .ZN(n4863) );
  NAND3_X1 U6261 ( .A1(n5203), .A2(n5202), .A3(n5020), .ZN(n5488) );
  NAND2_X1 U6262 ( .A1(n5585), .A2(n5584), .ZN(n4869) );
  NAND2_X1 U6263 ( .A1(n5370), .A2(n4319), .ZN(n4873) );
  NAND2_X1 U6264 ( .A1(n4873), .A2(n4874), .ZN(n5402) );
  OAI21_X1 U6265 ( .B1(n5370), .B2(n4879), .A(n4876), .ZN(n5417) );
  NAND2_X1 U6266 ( .A1(n5370), .A2(n5369), .ZN(n4881) );
  NAND2_X1 U6267 ( .A1(n5519), .A2(n4890), .ZN(n4883) );
  NAND2_X1 U6268 ( .A1(n4901), .A2(n4394), .ZN(n5019) );
  NAND2_X1 U6269 ( .A1(n5447), .A2(n5017), .ZN(n5461) );
  NAND3_X1 U6270 ( .A1(n4958), .A2(n4957), .A3(P2_DATAO_REG_1__SCAN_IN), .ZN(
        n4904) );
  INV_X1 U6271 ( .A(n4957), .ZN(n4906) );
  INV_X1 U6272 ( .A(n4915), .ZN(n4907) );
  NOR2_X1 U6273 ( .A1(n4915), .A2(n4913), .ZN(n4908) );
  NOR2_X1 U6274 ( .A1(n7839), .A2(n4915), .ZN(n7882) );
  INV_X1 U6275 ( .A(n7841), .ZN(n4914) );
  NAND2_X1 U6276 ( .A1(n7027), .A2(n4329), .ZN(n7208) );
  XNOR2_X1 U6277 ( .A(n7319), .B(n5977), .ZN(n6852) );
  INV_X1 U6278 ( .A(n4932), .ZN(n8519) );
  NOR2_X1 U6279 ( .A1(n6091), .A2(n8863), .ZN(n4934) );
  NAND2_X1 U6280 ( .A1(n5136), .A2(n5135), .ZN(n5354) );
  INV_X1 U6281 ( .A(n5347), .ZN(n5136) );
  NAND2_X1 U6282 ( .A1(n8477), .A2(n8478), .ZN(n8479) );
  AND2_X2 U6283 ( .A1(n7439), .A2(n7444), .ZN(n7437) );
  NAND2_X1 U6284 ( .A1(n6338), .A2(n6350), .ZN(n6800) );
  INV_X1 U6285 ( .A(n5207), .ZN(n5371) );
  INV_X1 U6286 ( .A(n5871), .ZN(n8468) );
  OR2_X1 U6287 ( .A1(n7304), .A2(n7228), .ZN(n7227) );
  NAND2_X1 U6288 ( .A1(n8885), .A2(n8884), .ZN(n8886) );
  NAND2_X1 U6289 ( .A1(n8938), .A2(n10158), .ZN(n8885) );
  NAND2_X1 U6290 ( .A1(n5123), .A2(n5115), .ZN(n5810) );
  OAI21_X1 U6291 ( .B1(n7129), .B2(n8082), .A(n6862), .ZN(n6863) );
  OR2_X1 U6292 ( .A1(n8402), .A2(n6213), .ZN(n6214) );
  INV_X1 U6293 ( .A(n9504), .ZN(n9505) );
  XNOR2_X1 U6294 ( .A(n6863), .B(n9111), .ZN(n6868) );
  NAND2_X1 U6295 ( .A1(n7850), .A2(n7861), .ZN(n7855) );
  OR2_X1 U6296 ( .A1(n6846), .A2(n5964), .ZN(n5901) );
  CLKBUF_X1 U6297 ( .A(n5809), .Z(n8084) );
  NAND2_X1 U6298 ( .A1(n5792), .A2(n9373), .ZN(n5793) );
  NAND2_X1 U6299 ( .A1(n5842), .A2(n5841), .ZN(n5845) );
  OR2_X1 U6300 ( .A1(n5842), .A2(n5841), .ZN(n5843) );
  NAND4_X2 U6301 ( .A1(n5926), .A2(n5925), .A3(n5924), .A4(n5923), .ZN(n8624)
         );
  INV_X2 U6302 ( .A(n5396), .ZN(n5649) );
  NAND3_X1 U6303 ( .A1(n6255), .A2(n6254), .A3(n6253), .ZN(n6315) );
  XNOR2_X1 U6304 ( .A(n7055), .B(n5951), .ZN(n5934) );
  NAND2_X1 U6305 ( .A1(n8575), .A2(n8576), .ZN(n6255) );
  XNOR2_X1 U6306 ( .A(n6212), .B(n6210), .ZN(n8575) );
  OR2_X1 U6307 ( .A1(n5948), .A2(n6366), .ZN(n5965) );
  NAND2_X1 U6308 ( .A1(n6169), .A2(n6168), .ZN(n8536) );
  AND2_X1 U6309 ( .A1(n6273), .A2(n8226), .ZN(n7062) );
  AOI21_X1 U6310 ( .B1(n6822), .B2(P1_REG1_REG_0__SCAN_IN), .A(n6859), .ZN(
        n6861) );
  AND2_X1 U6311 ( .A1(n6363), .A2(P1_U3086), .ZN(n6398) );
  INV_X1 U6312 ( .A(n6363), .ZN(n6364) );
  INV_X1 U6313 ( .A(n8801), .ZN(n8607) );
  AND2_X1 U6314 ( .A1(n6163), .A2(n6162), .ZN(n8801) );
  AND2_X1 U6315 ( .A1(n5112), .A2(n5111), .ZN(n4939) );
  INV_X1 U6316 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n4959) );
  AND2_X1 U6317 ( .A1(n8115), .A2(n8114), .ZN(n4940) );
  OR2_X1 U6318 ( .A1(n4603), .A2(n9571), .ZN(n4941) );
  NOR2_X1 U6319 ( .A1(n9185), .A2(n8160), .ZN(n4942) );
  OR2_X1 U6320 ( .A1(n9458), .A2(n9447), .ZN(n4944) );
  NOR2_X1 U6321 ( .A1(n5185), .A2(n5037), .ZN(n4945) );
  AND2_X1 U6322 ( .A1(n5119), .A2(n6553), .ZN(n4946) );
  AND2_X1 U6323 ( .A1(n7412), .A2(n7411), .ZN(n4947) );
  OR2_X1 U6324 ( .A1(n9525), .A2(n9709), .ZN(n4948) );
  INV_X1 U6325 ( .A(n9727), .ZN(n9708) );
  AND3_X1 U6326 ( .A1(n5313), .A2(n5312), .A3(n5311), .ZN(n4949) );
  INV_X1 U6327 ( .A(n9015), .ZN(n9020) );
  INV_X1 U6328 ( .A(n8973), .ZN(n8199) );
  OR2_X1 U6329 ( .A1(n6169), .A2(n6168), .ZN(n4950) );
  INV_X1 U6330 ( .A(n10158), .ZN(n10156) );
  AND2_X1 U6331 ( .A1(n8236), .A2(n10136), .ZN(n10120) );
  AND3_X1 U6332 ( .A1(n6301), .A2(n8589), .A3(n6309), .ZN(n4951) );
  NAND2_X1 U6333 ( .A1(n7045), .A2(n8813), .ZN(n8867) );
  AOI222_X1 U6334 ( .A1(n7455), .A2(n9033), .B1(n7270), .B2(n9049), .C1(n6822), 
        .C2(n9799), .ZN(n6860) );
  OR3_X1 U6335 ( .A1(n8454), .A2(n8453), .A3(n8452), .ZN(n4952) );
  NAND2_X1 U6336 ( .A1(n7755), .A2(n7711), .ZN(n4953) );
  INV_X1 U6337 ( .A(n8455), .ZN(n8711) );
  AND2_X1 U6338 ( .A1(n9391), .A2(n9390), .ZN(n5706) );
  INV_X1 U6339 ( .A(n7855), .ZN(n7853) );
  INV_X1 U6340 ( .A(n5789), .ZN(n5654) );
  INV_X1 U6341 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5105) );
  INV_X1 U6342 ( .A(n7210), .ZN(n6022) );
  NAND2_X1 U6343 ( .A1(n5655), .A2(n5654), .ZN(n5656) );
  AND2_X1 U6344 ( .A1(n5959), .A2(n7076), .ZN(n5960) );
  NAND2_X1 U6345 ( .A1(n5850), .A2(n5831), .ZN(n5835) );
  OR2_X1 U6346 ( .A1(n6224), .A2(P2_D_REG_1__SCAN_IN), .ZN(n6225) );
  INV_X1 U6347 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n5826) );
  INV_X1 U6348 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n5232) );
  OR2_X1 U6349 ( .A1(n6800), .A2(P1_D_REG_1__SCAN_IN), .ZN(n6351) );
  INV_X1 U6350 ( .A(SI_27_), .ZN(n5073) );
  INV_X1 U6351 ( .A(SI_26_), .ZN(n5068) );
  INV_X1 U6352 ( .A(SI_23_), .ZN(n5052) );
  AND2_X1 U6353 ( .A1(n5035), .A2(n5186), .ZN(n5036) );
  INV_X1 U6354 ( .A(SI_17_), .ZN(n5021) );
  INV_X1 U6355 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n5135) );
  INV_X1 U6356 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n5097) );
  OR2_X1 U6357 ( .A1(n6053), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6069) );
  INV_X1 U6358 ( .A(n8478), .ZN(n8223) );
  OR2_X1 U6359 ( .A1(n6191), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n6203) );
  AND2_X1 U6360 ( .A1(n6133), .A2(n6132), .ZN(n6145) );
  NOR2_X1 U6361 ( .A1(n6224), .A2(n6236), .ZN(n7041) );
  AOI21_X1 U6362 ( .B1(n8839), .B2(n8998), .A(n8849), .ZN(n8837) );
  OR2_X1 U6363 ( .A1(n8195), .A2(n7957), .ZN(n7959) );
  INV_X1 U6364 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5864) );
  INV_X1 U6365 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5841) );
  INV_X1 U6366 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n6059) );
  OR2_X1 U6367 ( .A1(n5393), .A2(n9093), .ZN(n5424) );
  OR2_X1 U6368 ( .A1(n7134), .A2(n7133), .ZN(n7131) );
  INV_X1 U6369 ( .A(n9241), .ZN(n9251) );
  INV_X1 U6370 ( .A(n9030), .ZN(n9111) );
  CLKBUF_X1 U6371 ( .A(n5741), .Z(n5670) );
  AND2_X1 U6372 ( .A1(n9890), .A2(n9264), .ZN(n8025) );
  NAND2_X1 U6373 ( .A1(n6351), .A2(n9791), .ZN(n7257) );
  AND2_X1 U6374 ( .A1(n5056), .A2(n5055), .ZN(n5551) );
  NOR2_X1 U6375 ( .A1(n5037), .A2(n5036), .ZN(n5038) );
  AND2_X1 U6376 ( .A1(n5386), .A2(n5208), .ZN(n5405) );
  INV_X1 U6377 ( .A(n8608), .ZN(n8853) );
  INV_X1 U6378 ( .A(n8593), .ZN(n8582) );
  OR2_X1 U6379 ( .A1(n9988), .A2(n9987), .ZN(n9991) );
  AND2_X1 U6380 ( .A1(n6260), .A2(n6259), .ZN(n8716) );
  OR2_X1 U6381 ( .A1(n6203), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n6216) );
  NAND2_X1 U6382 ( .A1(n6145), .A2(n6144), .ZN(n6157) );
  OR2_X1 U6383 ( .A1(n6109), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n6122) );
  OR2_X1 U6384 ( .A1(n6081), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n6083) );
  OR2_X1 U6385 ( .A1(n5999), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n6015) );
  INV_X1 U6386 ( .A(n8456), .ZN(n7049) );
  NAND2_X1 U6387 ( .A1(n8883), .A2(n8882), .ZN(n8938) );
  INV_X1 U6388 ( .A(n8838), .ZN(n10076) );
  NAND2_X1 U6389 ( .A1(n5849), .A2(n5832), .ZN(n5852) );
  OR2_X1 U6390 ( .A1(n6061), .A2(P2_IR_REG_11__SCAN_IN), .ZN(n6065) );
  INV_X1 U6391 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n9093) );
  OR2_X1 U6392 ( .A1(n5572), .A2(n5571), .ZN(n5589) );
  OR2_X1 U6393 ( .A1(n5377), .A2(n5376), .ZN(n5393) );
  INV_X1 U6394 ( .A(n9665), .ZN(n9447) );
  NAND2_X1 U6395 ( .A1(n6879), .A2(n7148), .ZN(n9255) );
  INV_X1 U6396 ( .A(n5613), .ZN(n5628) );
  INV_X1 U6397 ( .A(n8467), .ZN(n7148) );
  AND2_X1 U6398 ( .A1(n7802), .A2(n7702), .ZN(n7262) );
  NOR2_X1 U6399 ( .A1(n9770), .A2(n9531), .ZN(n8093) );
  INV_X1 U6400 ( .A(n9718), .ZN(n9530) );
  OR2_X1 U6401 ( .A1(n4315), .A2(n7303), .ZN(n9632) );
  OR2_X1 U6402 ( .A1(n6800), .A2(P1_D_REG_0__SCAN_IN), .ZN(n6353) );
  INV_X1 U6403 ( .A(n5755), .ZN(n9618) );
  INV_X1 U6404 ( .A(n9573), .ZN(n9889) );
  AND2_X1 U6405 ( .A1(n7627), .A2(n7513), .ZN(n7771) );
  NAND2_X1 U6406 ( .A1(n6553), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5125) );
  INV_X1 U6407 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n5805) );
  NAND2_X1 U6408 ( .A1(n5504), .A2(n6523), .ZN(n5506) );
  OAI21_X1 U6409 ( .B1(n8205), .B2(n8602), .A(n6289), .ZN(n6290) );
  OR2_X1 U6410 ( .A1(n8252), .A2(n5933), .ZN(n6961) );
  AND2_X1 U6411 ( .A1(n6275), .A2(n6274), .ZN(n8593) );
  NAND2_X1 U6412 ( .A1(n7039), .A2(n7401), .ZN(n8813) );
  AND2_X1 U6413 ( .A1(n6198), .A2(n6197), .ZN(n8765) );
  INV_X1 U6414 ( .A(n9989), .ZN(n10057) );
  INV_X1 U6415 ( .A(n8654), .ZN(n10049) );
  INV_X1 U6416 ( .A(n8760), .ZN(n7046) );
  INV_X1 U6417 ( .A(n8289), .ZN(n8430) );
  INV_X1 U6418 ( .A(n5964), .ZN(n8404) );
  AND2_X1 U6419 ( .A1(n10158), .A2(n10141), .ZN(n8927) );
  AND2_X1 U6420 ( .A1(n8715), .A2(n8714), .ZN(n8933) );
  INV_X1 U6421 ( .A(n8440), .ZN(n8862) );
  INV_X1 U6422 ( .A(n8969), .ZN(n9004) );
  INV_X1 U6423 ( .A(n10118), .ZN(n10141) );
  INV_X1 U6424 ( .A(n10120), .ZN(n10104) );
  XNOR2_X1 U6425 ( .A(n6242), .B(n6241), .ZN(n6579) );
  XNOR2_X1 U6426 ( .A(n5896), .B(P2_IR_REG_15__SCAN_IN), .ZN(n10017) );
  INV_X1 U6427 ( .A(n9255), .ZN(n9228) );
  AND2_X1 U6428 ( .A1(n6828), .A2(n6825), .ZN(n9237) );
  AND2_X1 U6429 ( .A1(n5172), .A2(n5171), .ZN(n9261) );
  AND4_X1 U6430 ( .A1(n5499), .A2(n5498), .A3(n5497), .A4(n5496), .ZN(n9556)
         );
  AND4_X1 U6431 ( .A1(n5458), .A2(n5457), .A3(n5456), .A4(n5455), .ZN(n9617)
         );
  OR2_X1 U6432 ( .A1(n6658), .A2(n7148), .ZN(n9851) );
  INV_X1 U6433 ( .A(n6652), .ZN(n9309) );
  INV_X1 U6434 ( .A(n7915), .ZN(n8054) );
  AND2_X1 U6435 ( .A1(n7262), .A2(n7526), .ZN(n9573) );
  INV_X1 U6436 ( .A(n9532), .ZN(n9898) );
  NAND2_X1 U6437 ( .A1(n9632), .A2(n7335), .ZN(n9907) );
  INV_X1 U6438 ( .A(n9962), .ZN(n9876) );
  AND2_X1 U6439 ( .A1(n6353), .A2(n9792), .ZN(n6802) );
  INV_X1 U6440 ( .A(n9964), .ZN(n9741) );
  AND2_X1 U6441 ( .A1(n6820), .A2(n6316), .ZN(n6831) );
  INV_X1 U6442 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n7538) );
  INV_X1 U6443 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n7547) );
  INV_X1 U6444 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n7554) );
  INV_X1 U6445 ( .A(n6290), .ZN(n6291) );
  NAND2_X1 U6446 ( .A1(n6315), .A2(n4951), .ZN(n6313) );
  INV_X1 U6447 ( .A(n8962), .ZN(n8898) );
  INV_X1 U6448 ( .A(n8589), .ZN(n8573) );
  AND2_X1 U6449 ( .A1(n6258), .A2(n8813), .ZN(n8602) );
  INV_X1 U6450 ( .A(n8382), .ZN(n8732) );
  INV_X1 U6451 ( .A(n8561), .ZN(n8788) );
  INV_X1 U6452 ( .A(n8596), .ZN(n8610) );
  INV_X1 U6453 ( .A(n10075), .ZN(n8616) );
  OR2_X1 U6454 ( .A1(n6583), .A2(n6590), .ZN(n10064) );
  NAND2_X1 U6455 ( .A1(n7047), .A2(n7046), .ZN(n8779) );
  INV_X1 U6456 ( .A(n8867), .ZN(n10092) );
  INV_X1 U6457 ( .A(n10092), .ZN(n10091) );
  INV_X1 U6458 ( .A(n8927), .ZN(n8909) );
  NAND2_X1 U6459 ( .A1(n10158), .A2(n10104), .ZN(n8930) );
  AND2_X2 U6460 ( .A1(n7408), .A2(n7407), .ZN(n10158) );
  OR2_X1 U6461 ( .A1(n10144), .A2(n10118), .ZN(n8969) );
  OR2_X1 U6462 ( .A1(n10144), .A2(n10120), .ZN(n9008) );
  AND2_X1 U6463 ( .A1(n6756), .A2(n6755), .ZN(n10144) );
  AND2_X1 U6464 ( .A1(n8067), .A2(n7950), .ZN(n6378) );
  NAND2_X1 U6465 ( .A1(n7039), .A2(n6224), .ZN(n6380) );
  INV_X1 U6466 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n7820) );
  INV_X1 U6467 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n7237) );
  INV_X1 U6468 ( .A(n7118), .ZN(n7104) );
  INV_X1 U6469 ( .A(n9257), .ZN(n9247) );
  AND3_X1 U6470 ( .A1(n5652), .A2(n5651), .A3(n5650), .ZN(n9393) );
  INV_X1 U6471 ( .A(n9617), .ZN(n9881) );
  OR2_X1 U6472 ( .A1(n6658), .A2(n6919), .ZN(n9861) );
  INV_X1 U6473 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n9855) );
  INV_X1 U6474 ( .A(n9635), .ZN(n9904) );
  AND2_X1 U6475 ( .A1(n9883), .A2(n9882), .ZN(n9946) );
  NAND2_X1 U6476 ( .A1(n6356), .A2(n6802), .ZN(n9981) );
  NAND2_X1 U6477 ( .A1(n6356), .A2(n7260), .ZN(n9966) );
  NAND2_X2 U6478 ( .A1(n6800), .A2(n6831), .ZN(n9913) );
  INV_X1 U6479 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n8070) );
  XNOR2_X1 U6480 ( .A(n5147), .B(n5146), .ZN(n7526) );
  INV_X1 U6481 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n7239) );
  INV_X1 U6482 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n6601) );
  INV_X2 U6483 ( .A(n6398), .ZN(n9797) );
  INV_X2 U6484 ( .A(n8623), .ZN(P2_U3893) );
  NOR2_X2 U6485 ( .A1(n6820), .A2(n6317), .ZN(P1_U3973) );
  INV_X1 U6486 ( .A(SI_1_), .ZN(n4960) );
  INV_X1 U6487 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n4964) );
  INV_X1 U6488 ( .A(SI_0_), .ZN(n4965) );
  NAND2_X1 U6489 ( .A1(n4968), .A2(SI_2_), .ZN(n4970) );
  NAND2_X1 U6490 ( .A1(n5274), .A2(n4969), .ZN(n5277) );
  NAND2_X1 U6491 ( .A1(n5277), .A2(n4970), .ZN(n5290) );
  NAND2_X1 U6492 ( .A1(n4971), .A2(SI_3_), .ZN(n4975) );
  INV_X1 U6493 ( .A(n4971), .ZN(n4973) );
  INV_X1 U6494 ( .A(SI_3_), .ZN(n4972) );
  NAND2_X1 U6495 ( .A1(n4973), .A2(n4972), .ZN(n4974) );
  NAND2_X1 U6496 ( .A1(n5292), .A2(n4975), .ZN(n5301) );
  MUX2_X1 U6497 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .S(n6363), .Z(n4976) );
  NAND2_X1 U6498 ( .A1(n4976), .A2(SI_4_), .ZN(n4980) );
  INV_X1 U6499 ( .A(n4976), .ZN(n4978) );
  INV_X1 U6500 ( .A(SI_4_), .ZN(n4977) );
  NAND2_X1 U6501 ( .A1(n4978), .A2(n4977), .ZN(n4979) );
  AND2_X1 U6502 ( .A1(n4980), .A2(n4979), .ZN(n5300) );
  NAND2_X1 U6503 ( .A1(n4981), .A2(SI_5_), .ZN(n4985) );
  INV_X1 U6504 ( .A(n4981), .ZN(n4983) );
  INV_X1 U6505 ( .A(SI_5_), .ZN(n4982) );
  NAND2_X1 U6506 ( .A1(n4983), .A2(n4982), .ZN(n4984) );
  AND2_X1 U6507 ( .A1(n4985), .A2(n4984), .ZN(n5324) );
  NAND2_X1 U6508 ( .A1(n4986), .A2(SI_6_), .ZN(n4990) );
  INV_X1 U6509 ( .A(n4986), .ZN(n4988) );
  INV_X1 U6510 ( .A(SI_6_), .ZN(n4987) );
  NAND2_X1 U6511 ( .A1(n4988), .A2(n4987), .ZN(n4989) );
  AND2_X1 U6512 ( .A1(n4989), .A2(n4990), .ZN(n5240) );
  MUX2_X1 U6513 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n6363), .Z(n4991) );
  NAND2_X1 U6514 ( .A1(n4991), .A2(SI_7_), .ZN(n4995) );
  INV_X1 U6515 ( .A(n4991), .ZN(n4993) );
  INV_X1 U6516 ( .A(SI_7_), .ZN(n4992) );
  NAND2_X1 U6517 ( .A1(n4993), .A2(n4992), .ZN(n4994) );
  AND2_X1 U6518 ( .A1(n4995), .A2(n4994), .ZN(n5343) );
  MUX2_X1 U6519 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .S(n6363), .Z(n4997) );
  XNOR2_X1 U6520 ( .A(n4997), .B(SI_8_), .ZN(n5352) );
  INV_X1 U6521 ( .A(n5352), .ZN(n4996) );
  INV_X1 U6522 ( .A(n4997), .ZN(n4999) );
  INV_X1 U6523 ( .A(SI_8_), .ZN(n4998) );
  NAND2_X1 U6524 ( .A1(n4999), .A2(n4998), .ZN(n5000) );
  MUX2_X1 U6525 ( .A(n6605), .B(n6601), .S(n6363), .Z(n5002) );
  XNOR2_X1 U6526 ( .A(n5002), .B(SI_9_), .ZN(n5369) );
  INV_X1 U6527 ( .A(n5002), .ZN(n5003) );
  NOR2_X1 U6528 ( .A1(n5003), .A2(SI_9_), .ZN(n5004) );
  MUX2_X1 U6529 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .S(n6363), .Z(n5005) );
  NAND2_X1 U6530 ( .A1(n5005), .A2(SI_10_), .ZN(n5009) );
  INV_X1 U6531 ( .A(n5005), .ZN(n5007) );
  INV_X1 U6532 ( .A(SI_10_), .ZN(n5006) );
  NAND2_X1 U6533 ( .A1(n5007), .A2(n5006), .ZN(n5008) );
  NAND2_X1 U6534 ( .A1(n5009), .A2(n5008), .ZN(n5383) );
  MUX2_X1 U6535 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .S(n6363), .Z(n5010) );
  XNOR2_X1 U6536 ( .A(n5010), .B(SI_11_), .ZN(n5418) );
  MUX2_X1 U6537 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .S(n6363), .Z(n5011) );
  NAND2_X1 U6538 ( .A1(n5011), .A2(SI_12_), .ZN(n5012) );
  OAI21_X1 U6539 ( .B1(n5011), .B2(SI_12_), .A(n5012), .ZN(n5401) );
  MUX2_X1 U6540 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n6363), .Z(n5013) );
  NAND2_X1 U6541 ( .A1(n5013), .A2(SI_13_), .ZN(n5017) );
  INV_X1 U6542 ( .A(n5013), .ZN(n5015) );
  INV_X1 U6543 ( .A(SI_13_), .ZN(n5014) );
  NAND2_X1 U6544 ( .A1(n5015), .A2(n5014), .ZN(n5016) );
  MUX2_X1 U6545 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n6363), .Z(n5459) );
  OR2_X2 U6546 ( .A1(n5224), .A2(SI_15_), .ZN(n5203) );
  MUX2_X1 U6547 ( .A(n7237), .B(n7239), .S(n6363), .Z(n5204) );
  INV_X1 U6548 ( .A(n5204), .ZN(n5025) );
  OR2_X1 U6549 ( .A1(n5025), .A2(SI_16_), .ZN(n5020) );
  MUX2_X1 U6550 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .S(n6363), .Z(n5222) );
  INV_X1 U6551 ( .A(n5222), .ZN(n5018) );
  NAND2_X1 U6552 ( .A1(n5019), .A2(n5018), .ZN(n5202) );
  MUX2_X1 U6553 ( .A(n7295), .B(n7294), .S(n6363), .Z(n5022) );
  NAND2_X1 U6554 ( .A1(n5022), .A2(n5021), .ZN(n5027) );
  INV_X1 U6555 ( .A(n5022), .ZN(n5023) );
  NAND2_X1 U6556 ( .A1(n5023), .A2(SI_17_), .ZN(n5024) );
  NAND2_X1 U6557 ( .A1(n5027), .A2(n5024), .ZN(n5489) );
  INV_X1 U6558 ( .A(n5489), .ZN(n5026) );
  NAND2_X1 U6559 ( .A1(n5025), .A2(SI_16_), .ZN(n5487) );
  MUX2_X1 U6560 ( .A(n7386), .B(n7425), .S(n6363), .Z(n5033) );
  XNOR2_X1 U6561 ( .A(n5033), .B(SI_18_), .ZN(n5502) );
  INV_X1 U6562 ( .A(n5502), .ZN(n5185) );
  MUX2_X1 U6563 ( .A(n7473), .B(n8472), .S(n6363), .Z(n5029) );
  NAND2_X1 U6564 ( .A1(n5029), .A2(n5028), .ZN(n5032) );
  INV_X1 U6565 ( .A(n5032), .ZN(n5037) );
  INV_X1 U6566 ( .A(n5029), .ZN(n5030) );
  NAND2_X1 U6567 ( .A1(n5030), .A2(SI_19_), .ZN(n5031) );
  NAND2_X1 U6568 ( .A1(n5032), .A2(n5031), .ZN(n5188) );
  INV_X1 U6569 ( .A(n5188), .ZN(n5035) );
  INV_X1 U6570 ( .A(n5033), .ZN(n5034) );
  NAND2_X1 U6571 ( .A1(n5034), .A2(SI_18_), .ZN(n5186) );
  AOI21_X2 U6572 ( .B1(n5039), .B2(n4945), .A(n5038), .ZN(n5176) );
  MUX2_X1 U6573 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(P2_DATAO_REG_20__SCAN_IN), 
        .S(n6363), .Z(n5174) );
  INV_X1 U6574 ( .A(n5174), .ZN(n5040) );
  OAI21_X1 U6575 ( .B1(n5176), .B2(n5173), .A(n5040), .ZN(n5042) );
  NAND2_X1 U6576 ( .A1(n5176), .A2(n5173), .ZN(n5041) );
  MUX2_X1 U6577 ( .A(n7703), .B(n7701), .S(n6363), .Z(n5520) );
  NOR2_X1 U6578 ( .A1(n5043), .A2(SI_21_), .ZN(n5045) );
  NAND2_X1 U6579 ( .A1(n5043), .A2(SI_21_), .ZN(n5044) );
  MUX2_X1 U6580 ( .A(n7801), .B(n7804), .S(n6363), .Z(n5047) );
  INV_X1 U6581 ( .A(SI_22_), .ZN(n5046) );
  NAND2_X1 U6582 ( .A1(n5047), .A2(n5046), .ZN(n5050) );
  INV_X1 U6583 ( .A(n5047), .ZN(n5048) );
  NAND2_X1 U6584 ( .A1(n5048), .A2(SI_22_), .ZN(n5049) );
  NAND2_X1 U6585 ( .A1(n5050), .A2(n5049), .ZN(n5541) );
  INV_X1 U6586 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n5051) );
  MUX2_X1 U6587 ( .A(n7820), .B(n5051), .S(n6363), .Z(n5053) );
  NAND2_X1 U6588 ( .A1(n5053), .A2(n5052), .ZN(n5056) );
  INV_X1 U6589 ( .A(n5053), .ZN(n5054) );
  NAND2_X1 U6590 ( .A1(n5054), .A2(SI_23_), .ZN(n5055) );
  NAND2_X1 U6591 ( .A1(n5554), .A2(n5056), .ZN(n5568) );
  INV_X1 U6592 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7948) );
  INV_X1 U6593 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7901) );
  MUX2_X1 U6594 ( .A(n7948), .B(n7901), .S(n6363), .Z(n5058) );
  INV_X1 U6595 ( .A(SI_24_), .ZN(n5057) );
  NAND2_X1 U6596 ( .A1(n5058), .A2(n5057), .ZN(n5061) );
  INV_X1 U6597 ( .A(n5058), .ZN(n5059) );
  NAND2_X1 U6598 ( .A1(n5059), .A2(SI_24_), .ZN(n5060) );
  NAND2_X1 U6599 ( .A1(n5568), .A2(n5567), .ZN(n5062) );
  NAND2_X1 U6600 ( .A1(n5062), .A2(n5061), .ZN(n5585) );
  INV_X1 U6601 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n8037) );
  INV_X1 U6602 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n8036) );
  MUX2_X1 U6603 ( .A(n8037), .B(n8036), .S(n6363), .Z(n5064) );
  INV_X1 U6604 ( .A(SI_25_), .ZN(n5063) );
  NAND2_X1 U6605 ( .A1(n5064), .A2(n5063), .ZN(n5067) );
  INV_X1 U6606 ( .A(n5064), .ZN(n5065) );
  NAND2_X1 U6607 ( .A1(n5065), .A2(SI_25_), .ZN(n5066) );
  INV_X1 U6608 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n8066) );
  MUX2_X1 U6609 ( .A(n8066), .B(n8070), .S(n6363), .Z(n5069) );
  NAND2_X1 U6610 ( .A1(n5069), .A2(n5068), .ZN(n5072) );
  INV_X1 U6611 ( .A(n5069), .ZN(n5070) );
  NAND2_X1 U6612 ( .A1(n5070), .A2(SI_26_), .ZN(n5071) );
  INV_X1 U6613 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n6213) );
  INV_X1 U6614 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n8083) );
  MUX2_X1 U6615 ( .A(n6213), .B(n8083), .S(n6363), .Z(n5074) );
  NAND2_X1 U6616 ( .A1(n5074), .A2(n5073), .ZN(n5077) );
  INV_X1 U6617 ( .A(n5074), .ZN(n5075) );
  NAND2_X1 U6618 ( .A1(n5075), .A2(SI_27_), .ZN(n5076) );
  NAND2_X1 U6619 ( .A1(n5609), .A2(n5610), .ZN(n5078) );
  INV_X1 U6620 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n6294) );
  INV_X1 U6621 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n8466) );
  MUX2_X1 U6622 ( .A(n6294), .B(n8466), .S(n6363), .Z(n5080) );
  XNOR2_X1 U6623 ( .A(n5080), .B(SI_28_), .ZN(n5622) );
  NAND2_X1 U6624 ( .A1(n5623), .A2(n5622), .ZN(n5082) );
  INV_X1 U6625 ( .A(SI_28_), .ZN(n5079) );
  NAND2_X1 U6626 ( .A1(n5080), .A2(n5079), .ZN(n5081) );
  INV_X1 U6627 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n9016) );
  INV_X1 U6628 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n8075) );
  MUX2_X1 U6629 ( .A(n9016), .B(n8075), .S(n6363), .Z(n5084) );
  INV_X1 U6630 ( .A(SI_29_), .ZN(n5086) );
  OR2_X1 U6631 ( .A1(n5084), .A2(n5083), .ZN(n5085) );
  OAI21_X1 U6632 ( .B1(n5149), .B2(n5086), .A(n5085), .ZN(n5643) );
  INV_X1 U6633 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n8465) );
  INV_X1 U6634 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n8470) );
  MUX2_X1 U6635 ( .A(n8465), .B(n8470), .S(n6364), .Z(n5088) );
  INV_X1 U6636 ( .A(SI_30_), .ZN(n5087) );
  NAND2_X1 U6637 ( .A1(n5088), .A2(n5087), .ZN(n5091) );
  INV_X1 U6638 ( .A(n5088), .ZN(n5089) );
  NAND2_X1 U6639 ( .A1(n5089), .A2(SI_30_), .ZN(n5090) );
  NAND2_X1 U6640 ( .A1(n5091), .A2(n5090), .ZN(n5642) );
  OAI21_X1 U6641 ( .B1(n5643), .B2(n5642), .A(n5091), .ZN(n5095) );
  INV_X1 U6642 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n5092) );
  INV_X1 U6643 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n9011) );
  MUX2_X1 U6644 ( .A(n5092), .B(n9011), .S(n6364), .Z(n5093) );
  XNOR2_X1 U6645 ( .A(n5093), .B(SI_31_), .ZN(n5094) );
  XNOR2_X1 U6646 ( .A(n5095), .B(n5094), .ZN(n8401) );
  NOR2_X4 U6647 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5260) );
  NOR2_X1 U6648 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n5101) );
  NOR2_X1 U6649 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n5100) );
  NOR2_X1 U6650 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n5099) );
  NOR2_X1 U6651 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n5098) );
  NOR2_X1 U6652 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n5103) );
  NOR2_X1 U6653 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n5102) );
  INV_X2 U6654 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n6523) );
  NAND2_X1 U6655 ( .A1(n5801), .A2(n5800), .ZN(n5110) );
  NAND2_X1 U6656 ( .A1(n5110), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5106) );
  NAND2_X1 U6657 ( .A1(n5799), .A2(n5106), .ZN(n5804) );
  OAI21_X2 U6658 ( .B1(n5804), .B2(P1_IR_REG_26__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5108) );
  INV_X1 U6659 ( .A(n5110), .ZN(n5112) );
  NOR2_X1 U6660 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), .ZN(
        n5111) );
  NAND2_X1 U6661 ( .A1(n5120), .A2(n5119), .ZN(n5123) );
  NAND2_X1 U6662 ( .A1(n5118), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5114) );
  NAND2_X2 U6663 ( .A1(n5809), .A2(n5810), .ZN(n5267) );
  NAND2_X1 U6664 ( .A1(n8401), .A2(n5353), .ZN(n5117) );
  NAND2_X1 U6665 ( .A1(n5293), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n5116) );
  INV_X1 U6666 ( .A(n5118), .ZN(n5120) );
  NAND2_X1 U6667 ( .A1(n5120), .A2(n4946), .ZN(n5127) );
  INV_X1 U6668 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n5121) );
  NAND2_X1 U6669 ( .A1(n5123), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5124) );
  NAND2_X1 U6670 ( .A1(n5124), .A2(P1_IR_REG_29__SCAN_IN), .ZN(n5126) );
  NAND2_X1 U6671 ( .A1(n5647), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n5132) );
  INV_X1 U6672 ( .A(n5129), .ZN(n5167) );
  NAND2_X1 U6673 ( .A1(n5648), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n5131) );
  NAND2_X1 U6674 ( .A1(n5649), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n5130) );
  NAND3_X1 U6675 ( .A1(n5132), .A2(n5131), .A3(n5130), .ZN(n6388) );
  NAND2_X1 U6676 ( .A1(n5133), .A2(n5134), .ZN(n5347) );
  NOR2_X2 U6677 ( .A1(n5354), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n5207) );
  INV_X1 U6678 ( .A(n5137), .ZN(n5138) );
  NAND2_X1 U6679 ( .A1(n5207), .A2(n5138), .ZN(n5212) );
  NAND2_X1 U6680 ( .A1(n5491), .A2(n5139), .ZN(n5140) );
  XNOR2_X2 U6681 ( .A(n5142), .B(n5141), .ZN(n6818) );
  NAND2_X1 U6682 ( .A1(n4347), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5143) );
  NAND2_X1 U6683 ( .A1(n4385), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5144) );
  NAND2_X1 U6684 ( .A1(n5145), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5147) );
  NAND2_X1 U6685 ( .A1(n6814), .A2(n6888), .ZN(n6890) );
  AOI211_X1 U6686 ( .C1(n5790), .C2(n7268), .A(n6884), .B(n6890), .ZN(n5796)
         );
  INV_X1 U6687 ( .A(n9755), .ZN(n5148) );
  INV_X1 U6688 ( .A(n6388), .ZN(n5653) );
  INV_X1 U6689 ( .A(n7268), .ZN(n9373) );
  XNOR2_X2 U6690 ( .A(n5149), .B(SI_29_), .ZN(n8207) );
  NAND2_X1 U6691 ( .A1(n8207), .A2(n5353), .ZN(n5151) );
  NAND2_X1 U6692 ( .A1(n5644), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n5150) );
  NAND2_X2 U6693 ( .A1(n5151), .A2(n5150), .ZN(n6333) );
  NAND3_X1 U6694 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n5318) );
  INV_X1 U6695 ( .A(n5318), .ZN(n5152) );
  NAND2_X1 U6696 ( .A1(n5152), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5337) );
  INV_X1 U6697 ( .A(n5337), .ZN(n5153) );
  NAND2_X1 U6698 ( .A1(n5153), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5358) );
  INV_X1 U6699 ( .A(n5358), .ZN(n5154) );
  NAND2_X1 U6700 ( .A1(n5154), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5377) );
  INV_X1 U6701 ( .A(n5424), .ZN(n5155) );
  NAND2_X1 U6702 ( .A1(n5155), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5426) );
  INV_X1 U6703 ( .A(n5426), .ZN(n5156) );
  NAND2_X1 U6704 ( .A1(n5156), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n5453) );
  INV_X1 U6705 ( .A(n5469), .ZN(n5157) );
  NAND2_X1 U6706 ( .A1(n5157), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n5471) );
  INV_X1 U6707 ( .A(n5234), .ZN(n5158) );
  NAND2_X1 U6708 ( .A1(n5158), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n5494) );
  INV_X1 U6709 ( .A(n5510), .ZN(n5159) );
  NAND2_X1 U6710 ( .A1(n5159), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n5512) );
  INV_X1 U6711 ( .A(n5512), .ZN(n5160) );
  NAND2_X1 U6712 ( .A1(n5160), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n5194) );
  INV_X1 U6713 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n9186) );
  INV_X1 U6714 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n9133) );
  INV_X1 U6715 ( .A(n5544), .ZN(n5161) );
  NAND2_X1 U6716 ( .A1(n5161), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n5558) );
  INV_X1 U6717 ( .A(n5558), .ZN(n5162) );
  NAND2_X1 U6718 ( .A1(n5162), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n5572) );
  INV_X1 U6719 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n5571) );
  INV_X1 U6720 ( .A(n5589), .ZN(n5163) );
  NAND2_X1 U6721 ( .A1(n5163), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n5600) );
  INV_X1 U6722 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n9240) );
  INV_X1 U6723 ( .A(n5626), .ZN(n5165) );
  AND2_X1 U6724 ( .A1(P1_REG3_REG_28__SCAN_IN), .A2(P1_REG3_REG_27__SCAN_IN), 
        .ZN(n5164) );
  NAND2_X1 U6725 ( .A1(n5165), .A2(n5164), .ZN(n9407) );
  OR2_X1 U6726 ( .A1(n9407), .A2(n5628), .ZN(n5172) );
  INV_X1 U6727 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n9406) );
  NAND2_X1 U6728 ( .A1(n5649), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n5169) );
  NAND2_X1 U6729 ( .A1(n5647), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n5168) );
  OAI211_X1 U6730 ( .C1(n9406), .C2(n5616), .A(n5169), .B(n5168), .ZN(n5170)
         );
  INV_X1 U6731 ( .A(n5170), .ZN(n5171) );
  OR2_X2 U6732 ( .A1(n6333), .A2(n9261), .ZN(n5659) );
  NAND2_X1 U6733 ( .A1(n6333), .A2(n9261), .ZN(n5711) );
  XNOR2_X1 U6734 ( .A(n5174), .B(n5173), .ZN(n5175) );
  XNOR2_X1 U6735 ( .A(n5176), .B(n5175), .ZN(n7524) );
  NAND2_X1 U6736 ( .A1(n7524), .A2(n5353), .ZN(n5178) );
  NAND2_X1 U6737 ( .A1(n5293), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n5177) );
  NAND2_X1 U6738 ( .A1(n5647), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n5180) );
  NAND2_X1 U6739 ( .A1(n5648), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n5179) );
  AND2_X1 U6740 ( .A1(n5180), .A2(n5179), .ZN(n5184) );
  NAND2_X1 U6741 ( .A1(n5194), .A2(n9186), .ZN(n5181) );
  NAND2_X1 U6742 ( .A1(n5524), .A2(n5181), .ZN(n9533) );
  OR2_X1 U6743 ( .A1(n9533), .A2(n5628), .ZN(n5183) );
  NAND2_X1 U6744 ( .A1(n5649), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n5182) );
  NAND2_X1 U6745 ( .A1(n9705), .A2(n9709), .ZN(n8097) );
  NAND2_X1 U6746 ( .A1(n8098), .A2(n8097), .ZN(n9527) );
  OR2_X1 U6747 ( .A1(n5503), .A2(n5185), .ZN(n5187) );
  NAND2_X1 U6748 ( .A1(n5187), .A2(n5186), .ZN(n5189) );
  XNOR2_X1 U6749 ( .A(n5189), .B(n5188), .ZN(n7472) );
  NAND2_X1 U6750 ( .A1(n7472), .A2(n5353), .ZN(n5191) );
  AOI22_X1 U6751 ( .A1(n5644), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n7268), .B2(
        n5305), .ZN(n5190) );
  NAND2_X1 U6752 ( .A1(n8098), .A2(n5582), .ZN(n5192) );
  OAI21_X1 U6753 ( .B1(n9527), .B2(n9541), .A(n5192), .ZN(n5199) );
  INV_X1 U6754 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n9105) );
  NAND2_X1 U6755 ( .A1(n5512), .A2(n9105), .ZN(n5193) );
  AND2_X1 U6756 ( .A1(n5194), .A2(n5193), .ZN(n9542) );
  NAND2_X1 U6757 ( .A1(n9542), .A2(n5613), .ZN(n5198) );
  NAND2_X1 U6758 ( .A1(n5647), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n5197) );
  NAND2_X1 U6759 ( .A1(n5649), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n5196) );
  NAND2_X1 U6760 ( .A1(n5648), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n5195) );
  NAND4_X1 U6761 ( .A1(n5198), .A2(n5197), .A3(n5196), .A4(n5195), .ZN(n9718)
         );
  OR2_X1 U6762 ( .A1(n9541), .A2(n9530), .ZN(n5729) );
  NAND2_X1 U6763 ( .A1(n5199), .A2(n5729), .ZN(n5201) );
  NAND3_X1 U6764 ( .A1(n8097), .A2(n9718), .A3(n6889), .ZN(n5200) );
  NAND2_X1 U6765 ( .A1(n5201), .A2(n5200), .ZN(n5535) );
  NAND2_X1 U6766 ( .A1(n5203), .A2(n5202), .ZN(n5206) );
  XNOR2_X1 U6767 ( .A(n5204), .B(SI_16_), .ZN(n5205) );
  NAND2_X1 U6768 ( .A1(n7236), .A2(n5353), .ZN(n5215) );
  NOR2_X1 U6769 ( .A1(n5371), .A2(P1_IR_REG_9__SCAN_IN), .ZN(n5386) );
  NOR2_X1 U6770 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n5208) );
  INV_X1 U6771 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n5209) );
  NAND2_X1 U6772 ( .A1(n5405), .A2(n5209), .ZN(n5448) );
  INV_X1 U6773 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5226) );
  INV_X1 U6774 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n5227) );
  NAND2_X1 U6775 ( .A1(n5226), .A2(n5227), .ZN(n5210) );
  OAI21_X1 U6776 ( .B1(n5225), .B2(n5210), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n5211) );
  MUX2_X1 U6777 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5211), .S(
        P1_IR_REG_16__SCAN_IN), .Z(n5213) );
  NAND2_X1 U6778 ( .A1(n5213), .A2(n5212), .ZN(n7915) );
  AOI22_X1 U6779 ( .A1(n5644), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n5305), .B2(
        n8054), .ZN(n5214) );
  INV_X2 U6780 ( .A(n5631), .ZN(n5647) );
  NAND2_X1 U6781 ( .A1(n5647), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n5221) );
  NAND2_X1 U6782 ( .A1(n5648), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n5220) );
  INV_X1 U6783 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n5216) );
  NAND2_X1 U6784 ( .A1(n5234), .A2(n5216), .ZN(n5217) );
  AND2_X1 U6785 ( .A1(n5494), .A2(n5217), .ZN(n9584) );
  NAND2_X1 U6786 ( .A1(n5613), .A2(n9584), .ZN(n5219) );
  NAND2_X1 U6787 ( .A1(n5649), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n5218) );
  XNOR2_X1 U6788 ( .A(n5222), .B(SI_15_), .ZN(n5223) );
  XNOR2_X1 U6789 ( .A(n5224), .B(n5223), .ZN(n7141) );
  NAND2_X1 U6790 ( .A1(n7141), .A2(n5353), .ZN(n5231) );
  INV_X1 U6791 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n7144) );
  NAND2_X1 U6792 ( .A1(n5225), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5462) );
  NAND2_X1 U6793 ( .A1(n5462), .A2(n5226), .ZN(n5464) );
  NAND2_X1 U6794 ( .A1(n5464), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5228) );
  XNOR2_X1 U6795 ( .A(n5228), .B(n5227), .ZN(n9856) );
  OAI22_X1 U6796 ( .A1(n4601), .A2(n7144), .B1(n9856), .B2(n5267), .ZN(n5229)
         );
  INV_X1 U6797 ( .A(n5229), .ZN(n5230) );
  NAND2_X1 U6798 ( .A1(n5647), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n5238) );
  NAND2_X1 U6799 ( .A1(n5649), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n5237) );
  NAND2_X1 U6800 ( .A1(n5471), .A2(n5232), .ZN(n5233) );
  AND2_X1 U6801 ( .A1(n5234), .A2(n5233), .ZN(n9607) );
  NAND2_X1 U6802 ( .A1(n5613), .A2(n9607), .ZN(n5236) );
  NAND2_X1 U6803 ( .A1(n5648), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n5235) );
  NAND4_X1 U6804 ( .A1(n5238), .A2(n5237), .A3(n5236), .A4(n5235), .ZN(n9263)
         );
  INV_X1 U6805 ( .A(n9263), .ZN(n9736) );
  NAND2_X1 U6806 ( .A1(n9606), .A2(n9736), .ZN(n5779) );
  NOR2_X1 U6807 ( .A1(n9606), .A2(n6889), .ZN(n5239) );
  AOI21_X1 U6808 ( .B1(n5731), .B2(n4571), .A(n5239), .ZN(n5479) );
  NAND2_X1 U6809 ( .A1(n9583), .A2(n9571), .ZN(n5780) );
  AOI21_X1 U6810 ( .B1(n5780), .B2(n9263), .A(n6889), .ZN(n5478) );
  OR2_X1 U6811 ( .A1(n9606), .A2(n9736), .ZN(n5732) );
  NAND2_X1 U6812 ( .A1(n5731), .A2(n5732), .ZN(n5688) );
  OR2_X1 U6813 ( .A1(n5241), .A2(n5240), .ZN(n5242) );
  NAND2_X1 U6814 ( .A1(n5644), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n5246) );
  OR2_X1 U6815 ( .A1(n5133), .A2(n9793), .ZN(n5244) );
  XNOR2_X1 U6816 ( .A(n5244), .B(P1_IR_REG_6__SCAN_IN), .ZN(n9323) );
  NAND2_X1 U6817 ( .A1(n5305), .A2(n9323), .ZN(n5245) );
  NAND2_X1 U6818 ( .A1(n5647), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n5252) );
  NAND2_X1 U6819 ( .A1(n5649), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5251) );
  INV_X1 U6820 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n5247) );
  NAND2_X1 U6821 ( .A1(n5318), .A2(n5247), .ZN(n5248) );
  AND2_X1 U6822 ( .A1(n5337), .A2(n5248), .ZN(n7601) );
  NAND2_X1 U6823 ( .A1(n5613), .A2(n7601), .ZN(n5250) );
  NAND2_X1 U6824 ( .A1(n5648), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n5249) );
  INV_X1 U6825 ( .A(n7746), .ZN(n9269) );
  NAND2_X1 U6826 ( .A1(n9927), .A2(n9269), .ZN(n7503) );
  NAND2_X1 U6827 ( .A1(n5375), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5256) );
  NAND2_X1 U6828 ( .A1(n5310), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n5255) );
  NAND2_X1 U6829 ( .A1(n5284), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n5254) );
  NAND2_X1 U6830 ( .A1(n5283), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5253) );
  NAND4_X1 U6831 ( .A1(n5256), .A2(n5255), .A3(n5254), .A4(n5253), .ZN(n6835)
         );
  INV_X1 U6832 ( .A(n5260), .ZN(n5261) );
  INV_X1 U6833 ( .A(n6641), .ZN(n9281) );
  INV_X1 U6834 ( .A(n7145), .ZN(n5269) );
  NAND2_X1 U6835 ( .A1(n5375), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5265) );
  NAND2_X1 U6836 ( .A1(n5284), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5264) );
  NAND2_X1 U6837 ( .A1(n5310), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n5263) );
  NAND2_X1 U6838 ( .A1(n5283), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n5262) );
  NAND2_X1 U6839 ( .A1(n6363), .A2(SI_0_), .ZN(n5266) );
  XNOR2_X1 U6840 ( .A(n5266), .B(P2_DATAO_REG_0__SCAN_IN), .ZN(n9800) );
  MUX2_X1 U6841 ( .A(n9799), .B(n9800), .S(n5267), .Z(n7270) );
  NOR2_X1 U6842 ( .A1(n7455), .A2(n7150), .ZN(n7153) );
  NOR2_X1 U6843 ( .A1(n8082), .A2(n9274), .ZN(n5268) );
  INV_X1 U6844 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n9919) );
  NAND2_X1 U6845 ( .A1(n5283), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5272) );
  NAND2_X1 U6846 ( .A1(n5375), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5271) );
  NAND2_X1 U6847 ( .A1(n5310), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n5270) );
  INV_X1 U6849 ( .A(n5274), .ZN(n5276) );
  NAND2_X1 U6850 ( .A1(n5276), .A2(n5275), .ZN(n5278) );
  NAND2_X1 U6851 ( .A1(n5278), .A2(n5277), .ZN(n8078) );
  NAND2_X1 U6852 ( .A1(n5293), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n5281) );
  OR2_X1 U6853 ( .A1(n5260), .A2(n9793), .ZN(n5279) );
  XNOR2_X1 U6854 ( .A(n5279), .B(P1_IR_REG_2__SCAN_IN), .ZN(n6644) );
  NAND2_X1 U6855 ( .A1(n5305), .A2(n6644), .ZN(n5280) );
  OAI211_X1 U6856 ( .C1(n5308), .C2(n8078), .A(n5281), .B(n5280), .ZN(n5282)
         );
  NAND2_X1 U6857 ( .A1(n7220), .A2(n5282), .ZN(n5740) );
  NAND2_X1 U6858 ( .A1(n7225), .A2(n7219), .ZN(n5741) );
  INV_X1 U6859 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n7464) );
  NAND2_X1 U6860 ( .A1(n5310), .A2(n7464), .ZN(n5288) );
  NAND2_X1 U6861 ( .A1(n5375), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n5287) );
  NAND2_X1 U6862 ( .A1(n5283), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5286) );
  NAND2_X1 U6863 ( .A1(n5284), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5285) );
  OR2_X1 U6864 ( .A1(n5290), .A2(n5289), .ZN(n5291) );
  NAND2_X1 U6865 ( .A1(n5292), .A2(n5291), .ZN(n6365) );
  NAND2_X1 U6866 ( .A1(n5293), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n5299) );
  NAND2_X1 U6867 ( .A1(n5295), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5296) );
  MUX2_X1 U6868 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5296), .S(
        P1_IR_REG_3__SCAN_IN), .Z(n5297) );
  AND2_X1 U6869 ( .A1(n5294), .A2(n5297), .ZN(n9295) );
  NAND2_X1 U6870 ( .A1(n5305), .A2(n9295), .ZN(n5298) );
  NAND2_X1 U6871 ( .A1(n7330), .A2(n7228), .ZN(n5739) );
  NAND2_X1 U6872 ( .A1(n7224), .A2(n5739), .ZN(n5667) );
  INV_X1 U6873 ( .A(n7330), .ZN(n9272) );
  NAND2_X1 U6874 ( .A1(n7467), .A2(n9272), .ZN(n5738) );
  OR2_X1 U6875 ( .A1(n5301), .A2(n5300), .ZN(n5302) );
  NAND2_X1 U6876 ( .A1(n5303), .A2(n5302), .ZN(n6367) );
  NAND2_X1 U6877 ( .A1(n5644), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n5307) );
  NAND2_X1 U6878 ( .A1(n5294), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5304) );
  XNOR2_X1 U6879 ( .A(n5304), .B(P1_IR_REG_4__SCAN_IN), .ZN(n6650) );
  NAND2_X1 U6880 ( .A1(n5305), .A2(n6650), .ZN(n5306) );
  NAND2_X1 U6881 ( .A1(n5648), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n5314) );
  NAND2_X1 U6882 ( .A1(n5284), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5313) );
  INV_X1 U6883 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n5309) );
  XNOR2_X1 U6884 ( .A(n5309), .B(P1_REG3_REG_3__SCAN_IN), .ZN(n7338) );
  NAND2_X1 U6885 ( .A1(n5310), .A2(n7338), .ZN(n5312) );
  NAND2_X1 U6886 ( .A1(n5375), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5311) );
  NAND2_X1 U6887 ( .A1(n9921), .A2(n9271), .ZN(n5737) );
  NAND3_X1 U6888 ( .A1(n5667), .A2(n5738), .A3(n5737), .ZN(n5333) );
  NAND2_X1 U6889 ( .A1(n7418), .A2(n7339), .ZN(n5736) );
  NAND2_X1 U6890 ( .A1(n5375), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5323) );
  INV_X1 U6891 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n5316) );
  NAND2_X1 U6892 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n5315) );
  NAND2_X1 U6893 ( .A1(n5316), .A2(n5315), .ZN(n5317) );
  AND2_X1 U6894 ( .A1(n5318), .A2(n5317), .ZN(n9899) );
  NAND2_X1 U6895 ( .A1(n5613), .A2(n9899), .ZN(n5322) );
  NAND2_X1 U6896 ( .A1(n5648), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n5321) );
  INV_X1 U6897 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n5319) );
  OR2_X1 U6898 ( .A1(n5396), .A2(n5319), .ZN(n5320) );
  OR2_X1 U6899 ( .A1(n5325), .A2(n5324), .ZN(n5326) );
  NAND2_X1 U6900 ( .A1(n5327), .A2(n5326), .ZN(n6370) );
  NAND2_X1 U6901 ( .A1(n5644), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n5332) );
  NOR2_X1 U6902 ( .A1(n5328), .A2(n9793), .ZN(n5329) );
  MUX2_X1 U6903 ( .A(n9793), .B(n5329), .S(P1_IR_REG_5__SCAN_IN), .Z(n5330) );
  OR2_X1 U6904 ( .A1(n5330), .A2(n5133), .ZN(n6652) );
  NAND2_X1 U6905 ( .A1(n5305), .A2(n9309), .ZN(n5331) );
  NAND2_X1 U6906 ( .A1(n7597), .A2(n9900), .ZN(n5767) );
  INV_X1 U6907 ( .A(n7597), .ZN(n9270) );
  INV_X1 U6908 ( .A(n7504), .ZN(n5677) );
  INV_X1 U6909 ( .A(n5768), .ZN(n5335) );
  AND3_X1 U6910 ( .A1(n7504), .A2(n5767), .A3(n5582), .ZN(n5334) );
  NAND2_X1 U6911 ( .A1(n5649), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5342) );
  NAND2_X1 U6912 ( .A1(n5647), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5341) );
  INV_X1 U6913 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n5336) );
  NAND2_X1 U6914 ( .A1(n5337), .A2(n5336), .ZN(n5338) );
  AND2_X1 U6915 ( .A1(n5358), .A2(n5338), .ZN(n7749) );
  NAND2_X1 U6916 ( .A1(n5613), .A2(n7749), .ZN(n5340) );
  NAND2_X1 U6917 ( .A1(n5648), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n5339) );
  OR2_X1 U6918 ( .A1(n5344), .A2(n5343), .ZN(n5345) );
  OR2_X1 U6919 ( .A1(n6375), .A2(n5308), .ZN(n5350) );
  NAND2_X1 U6920 ( .A1(n5347), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5348) );
  XNOR2_X1 U6921 ( .A(n5348), .B(P1_IR_REG_7__SCAN_IN), .ZN(n9336) );
  AOI22_X1 U6922 ( .A1(n5644), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n5305), .B2(
        n9336), .ZN(n5349) );
  NAND2_X1 U6923 ( .A1(n5350), .A2(n5349), .ZN(n7767) );
  NAND2_X1 U6924 ( .A1(n7940), .A2(n7767), .ZN(n7635) );
  INV_X1 U6925 ( .A(n7767), .ZN(n7743) );
  INV_X1 U6926 ( .A(n7940), .ZN(n9268) );
  NAND2_X1 U6927 ( .A1(n7743), .A2(n9268), .ZN(n5364) );
  NAND2_X1 U6928 ( .A1(n7635), .A2(n5364), .ZN(n7511) );
  INV_X1 U6929 ( .A(n7511), .ZN(n7508) );
  NAND2_X1 U6930 ( .A1(n5351), .A2(n7508), .ZN(n5366) );
  NAND2_X1 U6931 ( .A1(n5354), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5355) );
  XNOR2_X1 U6932 ( .A(n5355), .B(P1_IR_REG_8__SCAN_IN), .ZN(n6696) );
  AOI22_X1 U6933 ( .A1(n5293), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n5305), .B2(
        n6696), .ZN(n5356) );
  NAND2_X1 U6934 ( .A1(n5647), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5363) );
  NAND2_X1 U6935 ( .A1(n5648), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n5362) );
  INV_X1 U6936 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n5357) );
  NAND2_X1 U6937 ( .A1(n5358), .A2(n5357), .ZN(n5359) );
  AND2_X1 U6938 ( .A1(n5377), .A2(n5359), .ZN(n7939) );
  NAND2_X1 U6939 ( .A1(n5613), .A2(n7939), .ZN(n5361) );
  NAND2_X1 U6940 ( .A1(n5649), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n5360) );
  OR2_X1 U6941 ( .A1(n7938), .A2(n9174), .ZN(n7629) );
  AND2_X1 U6942 ( .A1(n7629), .A2(n5364), .ZN(n5747) );
  NAND2_X1 U6943 ( .A1(n7938), .A2(n9174), .ZN(n7628) );
  NAND2_X1 U6944 ( .A1(n7628), .A2(n7635), .ZN(n5675) );
  INV_X1 U6945 ( .A(n5675), .ZN(n7618) );
  MUX2_X1 U6946 ( .A(n5747), .B(n7618), .S(n6889), .Z(n5365) );
  NAND2_X1 U6947 ( .A1(n5366), .A2(n5365), .ZN(n5368) );
  MUX2_X1 U6948 ( .A(n7628), .B(n7629), .S(n6889), .Z(n5367) );
  NAND2_X1 U6949 ( .A1(n5368), .A2(n5367), .ZN(n5433) );
  NAND2_X1 U6950 ( .A1(n6600), .A2(n5353), .ZN(n5374) );
  NAND2_X1 U6951 ( .A1(n5371), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5372) );
  XNOR2_X1 U6952 ( .A(n5372), .B(P1_IR_REG_9__SCAN_IN), .ZN(n7085) );
  AOI22_X1 U6953 ( .A1(n5644), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n5305), .B2(
        n7085), .ZN(n5373) );
  NAND2_X1 U6954 ( .A1(n5375), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n5382) );
  NAND2_X1 U6955 ( .A1(n5649), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5381) );
  NAND2_X1 U6956 ( .A1(n5377), .A2(n5376), .ZN(n5378) );
  AND2_X1 U6957 ( .A1(n5393), .A2(n5378), .ZN(n9180) );
  NAND2_X1 U6958 ( .A1(n5613), .A2(n9180), .ZN(n5380) );
  INV_X1 U6959 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n7622) );
  OR2_X1 U6960 ( .A1(n5616), .A2(n7622), .ZN(n5379) );
  OR2_X1 U6961 ( .A1(n7984), .A2(n9092), .ZN(n7616) );
  NAND2_X1 U6962 ( .A1(n5433), .A2(n7616), .ZN(n5432) );
  NAND2_X1 U6963 ( .A1(n4327), .A2(n5383), .ZN(n5384) );
  NAND2_X1 U6964 ( .A1(n5385), .A2(n5384), .ZN(n6603) );
  OR2_X1 U6965 ( .A1(n6603), .A2(n5308), .ZN(n5392) );
  NOR2_X1 U6966 ( .A1(n5386), .A2(n9793), .ZN(n5387) );
  NAND2_X1 U6967 ( .A1(n5387), .A2(P1_IR_REG_10__SCAN_IN), .ZN(n5390) );
  INV_X1 U6968 ( .A(n5387), .ZN(n5389) );
  INV_X1 U6969 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5388) );
  NAND2_X1 U6970 ( .A1(n5389), .A2(n5388), .ZN(n5419) );
  AOI22_X1 U6971 ( .A1(n5293), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n5305), .B2(
        n9809), .ZN(n5391) );
  NAND2_X1 U6972 ( .A1(n5647), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n5400) );
  NAND2_X1 U6973 ( .A1(n5393), .A2(n9093), .ZN(n5394) );
  AND2_X1 U6974 ( .A1(n5424), .A2(n5394), .ZN(n9091) );
  NAND2_X1 U6975 ( .A1(n5613), .A2(n9091), .ZN(n5399) );
  NAND2_X1 U6976 ( .A1(n5648), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n5398) );
  INV_X1 U6977 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n5395) );
  OR2_X1 U6978 ( .A1(n5396), .A2(n5395), .ZN(n5397) );
  NAND2_X1 U6979 ( .A1(n8000), .A2(n9219), .ZN(n7723) );
  NAND2_X1 U6980 ( .A1(n7984), .A2(n9092), .ZN(n7615) );
  AND2_X1 U6981 ( .A1(n7723), .A2(n7615), .ZN(n5431) );
  NAND2_X1 U6982 ( .A1(n5402), .A2(n5401), .ZN(n5404) );
  NAND2_X1 U6983 ( .A1(n5404), .A2(n5403), .ZN(n6768) );
  OR2_X1 U6984 ( .A1(n6768), .A2(n5308), .ZN(n5410) );
  NOR2_X1 U6985 ( .A1(n5405), .A2(n9793), .ZN(n5406) );
  MUX2_X1 U6986 ( .A(n9793), .B(n5406), .S(P1_IR_REG_12__SCAN_IN), .Z(n5407)
         );
  INV_X1 U6987 ( .A(n5407), .ZN(n5408) );
  AOI22_X1 U6988 ( .A1(n5293), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n5305), .B2(
        n7910), .ZN(n5409) );
  INV_X1 U6989 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n5411) );
  NAND2_X1 U6990 ( .A1(n5426), .A2(n5411), .ZN(n5412) );
  AND2_X1 U6991 ( .A1(n5453), .A2(n5412), .ZN(n9884) );
  NAND2_X1 U6992 ( .A1(n5613), .A2(n9884), .ZN(n5416) );
  NAND2_X1 U6993 ( .A1(n5647), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n5415) );
  NAND2_X1 U6994 ( .A1(n5648), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n5414) );
  NAND2_X1 U6995 ( .A1(n5649), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5413) );
  OR2_X1 U6996 ( .A1(n9890), .A2(n9953), .ZN(n5734) );
  OR2_X1 U6997 ( .A1(n8000), .A2(n9219), .ZN(n5749) );
  XNOR2_X1 U6998 ( .A(n5417), .B(n5418), .ZN(n5913) );
  NAND2_X1 U6999 ( .A1(n5913), .A2(n5353), .ZN(n5422) );
  NAND2_X1 U7000 ( .A1(n5419), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5420) );
  XNOR2_X1 U7001 ( .A(n5420), .B(P1_IR_REG_11__SCAN_IN), .ZN(n9821) );
  AOI22_X1 U7002 ( .A1(n5644), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n5305), .B2(
        n9821), .ZN(n5421) );
  NAND2_X1 U7003 ( .A1(n5647), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n5430) );
  NAND2_X1 U7004 ( .A1(n5648), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n5429) );
  INV_X1 U7005 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n5423) );
  NAND2_X1 U7006 ( .A1(n5424), .A2(n5423), .ZN(n5425) );
  AND2_X1 U7007 ( .A1(n5426), .A2(n5425), .ZN(n9216) );
  NAND2_X1 U7008 ( .A1(n5613), .A2(n9216), .ZN(n5428) );
  NAND2_X1 U7009 ( .A1(n5649), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5427) );
  NAND4_X1 U7010 ( .A1(n5430), .A2(n5429), .A3(n5428), .A4(n5427), .ZN(n9878)
         );
  INV_X1 U7011 ( .A(n9878), .ZN(n9094) );
  OR2_X1 U7012 ( .A1(n9221), .A2(n9094), .ZN(n9873) );
  NAND2_X1 U7013 ( .A1(n5433), .A2(n7615), .ZN(n5436) );
  AND2_X1 U7014 ( .A1(n5749), .A2(n7616), .ZN(n5435) );
  NAND2_X1 U7015 ( .A1(n9890), .A2(n9953), .ZN(n8017) );
  NAND2_X1 U7016 ( .A1(n8017), .A2(n6889), .ZN(n5442) );
  NAND2_X1 U7017 ( .A1(n9221), .A2(n9094), .ZN(n5735) );
  AND2_X1 U7018 ( .A1(n5735), .A2(n7723), .ZN(n5773) );
  INV_X1 U7019 ( .A(n5773), .ZN(n5680) );
  OR2_X1 U7020 ( .A1(n5442), .A2(n5680), .ZN(n5434) );
  OR3_X1 U7021 ( .A1(n9890), .A2(n9953), .A3(n5582), .ZN(n5438) );
  AND2_X1 U7022 ( .A1(n5438), .A2(n5437), .ZN(n5441) );
  NAND2_X1 U7023 ( .A1(n5735), .A2(n9264), .ZN(n5439) );
  NAND3_X1 U7024 ( .A1(n9890), .A2(n5439), .A3(n5582), .ZN(n5440) );
  OAI211_X1 U7025 ( .C1(n5442), .C2(n9873), .A(n5441), .B(n5440), .ZN(n5443)
         );
  NAND2_X1 U7026 ( .A1(n5447), .A2(n5446), .ZN(n6846) );
  NAND2_X1 U7027 ( .A1(n5448), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5449) );
  XNOR2_X1 U7028 ( .A(n5449), .B(P1_IR_REG_13__SCAN_IN), .ZN(n9833) );
  AOI22_X1 U7029 ( .A1(n5644), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n5305), .B2(
        n9833), .ZN(n5450) );
  NAND2_X1 U7030 ( .A1(n5647), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n5458) );
  NAND2_X1 U7031 ( .A1(n5648), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n5457) );
  NAND2_X1 U7032 ( .A1(n5453), .A2(n5452), .ZN(n5454) );
  AND2_X1 U7033 ( .A1(n5469), .A2(n5454), .ZN(n9194) );
  NAND2_X1 U7034 ( .A1(n5613), .A2(n9194), .ZN(n5456) );
  NAND2_X1 U7035 ( .A1(n5649), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n5455) );
  OR2_X1 U7036 ( .A1(n9958), .A2(n9617), .ZN(n5733) );
  INV_X1 U7037 ( .A(n5733), .ZN(n5476) );
  XNOR2_X1 U7038 ( .A(n5459), .B(SI_14_), .ZN(n5460) );
  XNOR2_X1 U7039 ( .A(n5461), .B(n5460), .ZN(n6896) );
  NAND2_X1 U7040 ( .A1(n6896), .A2(n5353), .ZN(n5467) );
  INV_X1 U7041 ( .A(n5462), .ZN(n5463) );
  NAND2_X1 U7042 ( .A1(n5463), .A2(P1_IR_REG_14__SCAN_IN), .ZN(n5465) );
  AOI22_X1 U7043 ( .A1(n5293), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n5305), .B2(
        n9837), .ZN(n5466) );
  NAND2_X1 U7044 ( .A1(n5649), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5475) );
  NAND2_X1 U7045 ( .A1(n5647), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n5474) );
  INV_X1 U7046 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n5468) );
  NAND2_X1 U7047 ( .A1(n5469), .A2(n5468), .ZN(n5470) );
  AND2_X1 U7048 ( .A1(n5471), .A2(n5470), .ZN(n9628) );
  NAND2_X1 U7049 ( .A1(n5613), .A2(n9628), .ZN(n5473) );
  NAND2_X1 U7050 ( .A1(n5648), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n5472) );
  NAND4_X1 U7051 ( .A1(n5475), .A2(n5474), .A3(n5473), .A4(n5472), .ZN(n9601)
         );
  OR2_X1 U7052 ( .A1(n9749), .A2(n9955), .ZN(n5777) );
  NAND2_X1 U7053 ( .A1(n9749), .A2(n9955), .ZN(n5482) );
  NAND2_X1 U7054 ( .A1(n5777), .A2(n5482), .ZN(n5755) );
  NAND2_X1 U7055 ( .A1(n9958), .A2(n9617), .ZN(n9614) );
  INV_X1 U7056 ( .A(n9614), .ZN(n5480) );
  NOR2_X1 U7057 ( .A1(n5755), .A2(n5480), .ZN(n5776) );
  OAI22_X1 U7058 ( .A1(n5479), .A2(n5478), .B1(n5688), .B2(n5477), .ZN(n5501)
         );
  OAI211_X1 U7059 ( .C1(n5481), .C2(n5480), .A(n9618), .B(n5733), .ZN(n5483)
         );
  AND2_X1 U7060 ( .A1(n5779), .A2(n5482), .ZN(n5684) );
  NAND3_X1 U7061 ( .A1(n5780), .A2(n5483), .A3(n5684), .ZN(n5484) );
  NAND2_X1 U7062 ( .A1(n5484), .A2(n5731), .ZN(n5486) );
  INV_X1 U7063 ( .A(n5780), .ZN(n5485) );
  MUX2_X1 U7064 ( .A(n5486), .B(n5485), .S(n6889), .Z(n5500) );
  NAND2_X1 U7065 ( .A1(n5488), .A2(n5487), .ZN(n5490) );
  XNOR2_X1 U7066 ( .A(n5490), .B(n5489), .ZN(n7293) );
  NAND2_X1 U7067 ( .A1(n7293), .A2(n5353), .ZN(n5493) );
  XNOR2_X1 U7068 ( .A(n5491), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9349) );
  AOI22_X1 U7069 ( .A1(n5293), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n5305), .B2(
        n9349), .ZN(n5492) );
  NAND2_X1 U7070 ( .A1(n5649), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n5499) );
  NAND2_X1 U7071 ( .A1(n5647), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n5498) );
  NAND2_X1 U7072 ( .A1(n5494), .A2(n8059), .ZN(n5495) );
  AND2_X1 U7073 ( .A1(n5510), .A2(n5495), .ZN(n9567) );
  NAND2_X1 U7074 ( .A1(n5613), .A2(n9567), .ZN(n5497) );
  NAND2_X1 U7075 ( .A1(n5648), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n5496) );
  OR2_X1 U7076 ( .A1(n4605), .A2(n9556), .ZN(n5781) );
  NAND2_X1 U7077 ( .A1(n4605), .A2(n9556), .ZN(n5782) );
  OAI21_X1 U7078 ( .B1(n5501), .B2(n5500), .A(n9565), .ZN(n5532) );
  XNOR2_X1 U7079 ( .A(n5503), .B(n5502), .ZN(n7385) );
  NAND2_X1 U7080 ( .A1(n7385), .A2(n5353), .ZN(n5508) );
  OR2_X1 U7081 ( .A1(n5504), .A2(n6523), .ZN(n5505) );
  AND2_X1 U7082 ( .A1(n5506), .A2(n5505), .ZN(n9358) );
  AOI22_X1 U7083 ( .A1(n5644), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n5305), .B2(
        n9358), .ZN(n5507) );
  NAND2_X1 U7084 ( .A1(n5647), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n5516) );
  NAND2_X1 U7085 ( .A1(n5648), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n5515) );
  INV_X1 U7086 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n5509) );
  NAND2_X1 U7087 ( .A1(n5510), .A2(n5509), .ZN(n5511) );
  AND2_X1 U7088 ( .A1(n5512), .A2(n5511), .ZN(n9553) );
  NAND2_X1 U7089 ( .A1(n5613), .A2(n9553), .ZN(n5514) );
  NAND2_X1 U7090 ( .A1(n5649), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n5513) );
  NAND4_X1 U7091 ( .A1(n5516), .A2(n5515), .A3(n5514), .A4(n5513), .ZN(n9727)
         );
  OR2_X1 U7092 ( .A1(n9560), .A2(n9708), .ZN(n5730) );
  AND2_X1 U7093 ( .A1(n5781), .A2(n5730), .ZN(n5692) );
  NAND2_X1 U7094 ( .A1(n5532), .A2(n5692), .ZN(n5517) );
  NAND2_X1 U7095 ( .A1(n9541), .A2(n9530), .ZN(n5785) );
  NAND2_X1 U7096 ( .A1(n9560), .A2(n9708), .ZN(n5784) );
  NAND3_X1 U7097 ( .A1(n5517), .A2(n5785), .A3(n5784), .ZN(n5518) );
  NAND2_X1 U7098 ( .A1(n5535), .A2(n5518), .ZN(n5531) );
  XNOR2_X1 U7099 ( .A(n5520), .B(SI_21_), .ZN(n5521) );
  XNOR2_X1 U7100 ( .A(n5519), .B(n5521), .ZN(n7700) );
  NAND2_X1 U7101 ( .A1(n7700), .A2(n5353), .ZN(n5523) );
  NAND2_X1 U7102 ( .A1(n5293), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n5522) );
  NAND2_X1 U7103 ( .A1(n5524), .A2(n9133), .ZN(n5525) );
  AND2_X1 U7104 ( .A1(n5544), .A2(n5525), .ZN(n9515) );
  NAND2_X1 U7105 ( .A1(n9515), .A2(n5613), .ZN(n5528) );
  AOI22_X1 U7106 ( .A1(n5649), .A2(P1_REG0_REG_21__SCAN_IN), .B1(n5647), .B2(
        P1_REG1_REG_21__SCAN_IN), .ZN(n5527) );
  NAND2_X1 U7107 ( .A1(n5648), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n5526) );
  NAND2_X1 U7108 ( .A1(n9514), .A2(n9531), .ZN(n5727) );
  NAND2_X1 U7109 ( .A1(n5727), .A2(n8097), .ZN(n5697) );
  INV_X1 U7110 ( .A(n5697), .ZN(n5530) );
  INV_X1 U7111 ( .A(n5728), .ZN(n5529) );
  AOI21_X1 U7112 ( .B1(n5531), .B2(n5530), .A(n5529), .ZN(n5539) );
  AND2_X1 U7113 ( .A1(n5729), .A2(n5730), .ZN(n5693) );
  AND2_X1 U7114 ( .A1(n5784), .A2(n5782), .ZN(n5689) );
  NAND2_X1 U7115 ( .A1(n5532), .A2(n5689), .ZN(n5533) );
  NAND2_X1 U7116 ( .A1(n5693), .A2(n5533), .ZN(n5534) );
  NAND2_X1 U7117 ( .A1(n5535), .A2(n5534), .ZN(n5537) );
  AND2_X1 U7118 ( .A1(n5728), .A2(n8098), .ZN(n5665) );
  INV_X1 U7119 ( .A(n5727), .ZN(n5536) );
  AOI21_X1 U7120 ( .B1(n5537), .B2(n5665), .A(n5536), .ZN(n5538) );
  XNOR2_X1 U7121 ( .A(n5540), .B(n5541), .ZN(n7800) );
  NAND2_X1 U7122 ( .A1(n7800), .A2(n5353), .ZN(n5543) );
  NAND2_X1 U7123 ( .A1(n5293), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n5542) );
  INV_X1 U7124 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n9202) );
  NAND2_X1 U7125 ( .A1(n5544), .A2(n9202), .ZN(n5545) );
  NAND2_X1 U7126 ( .A1(n5558), .A2(n5545), .ZN(n9495) );
  OR2_X1 U7127 ( .A1(n9495), .A2(n5628), .ZN(n5550) );
  INV_X1 U7128 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n9496) );
  NAND2_X1 U7129 ( .A1(n5647), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n5547) );
  NAND2_X1 U7130 ( .A1(n5649), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n5546) );
  OAI211_X1 U7131 ( .C1(n9496), .C2(n5616), .A(n5547), .B(n5546), .ZN(n5548)
         );
  INV_X1 U7132 ( .A(n5548), .ZN(n5549) );
  NAND2_X1 U7133 ( .A1(n9499), .A2(n9680), .ZN(n8101) );
  OR2_X1 U7134 ( .A1(n5552), .A2(n5551), .ZN(n5553) );
  NAND2_X1 U7135 ( .A1(n5554), .A2(n5553), .ZN(n7817) );
  NAND2_X1 U7136 ( .A1(n7817), .A2(n5353), .ZN(n5556) );
  NAND2_X1 U7137 ( .A1(n5644), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n5555) );
  INV_X1 U7138 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n5557) );
  NAND2_X1 U7139 ( .A1(n5558), .A2(n5557), .ZN(n5559) );
  NAND2_X1 U7140 ( .A1(n5572), .A2(n5559), .ZN(n9081) );
  OR2_X1 U7141 ( .A1(n9081), .A2(n5628), .ZN(n5565) );
  INV_X1 U7142 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n5562) );
  NAND2_X1 U7143 ( .A1(n5647), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n5561) );
  NAND2_X1 U7144 ( .A1(n5649), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n5560) );
  OAI211_X1 U7145 ( .C1(n5616), .C2(n5562), .A(n5561), .B(n5560), .ZN(n5563)
         );
  INV_X1 U7146 ( .A(n5563), .ZN(n5564) );
  INV_X1 U7147 ( .A(n9690), .ZN(n8191) );
  OR2_X1 U7148 ( .A1(n9684), .A2(n8191), .ZN(n5726) );
  NAND2_X1 U7149 ( .A1(n5726), .A2(n8100), .ZN(n5661) );
  NAND2_X1 U7150 ( .A1(n9684), .A2(n8191), .ZN(n8103) );
  NAND2_X1 U7151 ( .A1(n8103), .A2(n8101), .ZN(n5566) );
  MUX2_X1 U7152 ( .A(n5661), .B(n5566), .S(n6889), .Z(n5581) );
  XNOR2_X1 U7153 ( .A(n5568), .B(n5567), .ZN(n7900) );
  NAND2_X1 U7154 ( .A1(n7900), .A2(n5353), .ZN(n5570) );
  NAND2_X1 U7155 ( .A1(n5644), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n5569) );
  NAND2_X1 U7156 ( .A1(n5572), .A2(n5571), .ZN(n5573) );
  AND2_X1 U7157 ( .A1(n5589), .A2(n5573), .ZN(n9470) );
  NAND2_X1 U7158 ( .A1(n9470), .A2(n5613), .ZN(n5579) );
  INV_X1 U7159 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n5576) );
  NAND2_X1 U7160 ( .A1(n5649), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n5575) );
  NAND2_X1 U7161 ( .A1(n5647), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n5574) );
  OAI211_X1 U7162 ( .C1(n5576), .C2(n5616), .A(n5575), .B(n5574), .ZN(n5577)
         );
  INV_X1 U7163 ( .A(n5577), .ZN(n5578) );
  NAND2_X1 U7164 ( .A1(n8096), .A2(n9681), .ZN(n5660) );
  MUX2_X1 U7165 ( .A(n8103), .B(n5726), .S(n6889), .Z(n5580) );
  MUX2_X1 U7166 ( .A(n5660), .B(n9385), .S(n5582), .Z(n5583) );
  INV_X1 U7167 ( .A(n5636), .ZN(n5608) );
  XNOR2_X1 U7168 ( .A(n5585), .B(n5584), .ZN(n8035) );
  NAND2_X1 U7169 ( .A1(n8035), .A2(n5353), .ZN(n5587) );
  NAND2_X1 U7170 ( .A1(n5293), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n5586) );
  INV_X1 U7171 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n5588) );
  NAND2_X1 U7172 ( .A1(n5589), .A2(n5588), .ZN(n5590) );
  NAND2_X1 U7173 ( .A1(n5600), .A2(n5590), .ZN(n9455) );
  INV_X1 U7174 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n9454) );
  NAND2_X1 U7175 ( .A1(n5649), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n5592) );
  NAND2_X1 U7176 ( .A1(n5647), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n5591) );
  OAI211_X1 U7177 ( .C1(n9454), .C2(n5616), .A(n5592), .B(n5591), .ZN(n5593)
         );
  INV_X1 U7178 ( .A(n5593), .ZN(n5594) );
  NAND2_X1 U7179 ( .A1(n9762), .A2(n9447), .ZN(n9387) );
  INV_X1 U7180 ( .A(n9387), .ZN(n5725) );
  NAND2_X1 U7181 ( .A1(n8065), .A2(n5353), .ZN(n5599) );
  NAND2_X1 U7182 ( .A1(n5644), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n5598) );
  AND2_X2 U7183 ( .A1(n5599), .A2(n5598), .ZN(n9669) );
  NAND2_X1 U7184 ( .A1(n5600), .A2(n9240), .ZN(n5601) );
  NAND2_X1 U7185 ( .A1(n9445), .A2(n5613), .ZN(n5607) );
  INV_X1 U7186 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n5604) );
  NAND2_X1 U7187 ( .A1(n5647), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n5603) );
  NAND2_X1 U7188 ( .A1(n5649), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n5602) );
  OAI211_X1 U7189 ( .C1(n5616), .C2(n5604), .A(n5603), .B(n5602), .ZN(n5605)
         );
  INV_X1 U7190 ( .A(n5605), .ZN(n5606) );
  INV_X1 U7191 ( .A(n9388), .ZN(n5635) );
  OAI211_X1 U7192 ( .C1(n5608), .C2(n5725), .A(n5724), .B(n5635), .ZN(n5621)
         );
  NAND2_X1 U7193 ( .A1(n6331), .A2(n9657), .ZN(n9389) );
  NAND2_X1 U7194 ( .A1(n8072), .A2(n5353), .ZN(n5612) );
  NAND2_X1 U7195 ( .A1(n5293), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n5611) );
  XNOR2_X1 U7196 ( .A(n5626), .B(P1_REG3_REG_27__SCAN_IN), .ZN(n9431) );
  NAND2_X1 U7197 ( .A1(n9431), .A2(n5613), .ZN(n5620) );
  INV_X1 U7198 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n5617) );
  NAND2_X1 U7199 ( .A1(n5649), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n5615) );
  NAND2_X1 U7200 ( .A1(n5647), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n5614) );
  OAI211_X1 U7201 ( .C1(n5617), .C2(n5616), .A(n5615), .B(n5614), .ZN(n5618)
         );
  INV_X1 U7202 ( .A(n5618), .ZN(n5619) );
  NAND2_X1 U7203 ( .A1(n9661), .A2(n9242), .ZN(n9390) );
  XNOR2_X1 U7204 ( .A(n5623), .B(n5622), .ZN(n6293) );
  NAND2_X1 U7205 ( .A1(n6293), .A2(n5353), .ZN(n5625) );
  NAND2_X1 U7206 ( .A1(n5644), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n5624) );
  INV_X1 U7207 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n9060) );
  INV_X1 U7208 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n9117) );
  OAI21_X1 U7209 ( .B1(n5626), .B2(n9060), .A(n9117), .ZN(n5627) );
  NAND2_X1 U7210 ( .A1(n5627), .A2(n9407), .ZN(n9419) );
  INV_X1 U7211 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n6405) );
  NAND2_X1 U7212 ( .A1(n5648), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n5630) );
  NAND2_X1 U7213 ( .A1(n5649), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n5629) );
  OAI211_X1 U7214 ( .C1(n5631), .C2(n6405), .A(n5630), .B(n5629), .ZN(n5632)
         );
  INV_X1 U7215 ( .A(n5632), .ZN(n5633) );
  NAND2_X1 U7216 ( .A1(n9389), .A2(n9387), .ZN(n5701) );
  AOI21_X1 U7217 ( .B1(n5636), .B2(n5635), .A(n5701), .ZN(n5637) );
  NAND2_X1 U7218 ( .A1(n5723), .A2(n5724), .ZN(n5704) );
  NAND2_X1 U7219 ( .A1(n9401), .A2(n9658), .ZN(n9391) );
  OAI21_X1 U7220 ( .B1(n5637), .B2(n5704), .A(n5706), .ZN(n5638) );
  MUX2_X1 U7221 ( .A(n5638), .B(n9391), .S(n6889), .Z(n5639) );
  MUX2_X1 U7222 ( .A(n5711), .B(n5659), .S(n6889), .Z(n5640) );
  NAND2_X1 U7223 ( .A1(n5641), .A2(n5640), .ZN(n5657) );
  NAND2_X1 U7224 ( .A1(n8464), .A2(n5353), .ZN(n5646) );
  NAND2_X1 U7225 ( .A1(n5644), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n5645) );
  INV_X1 U7226 ( .A(n5790), .ZN(n5655) );
  NAND2_X1 U7227 ( .A1(n5647), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n5652) );
  NAND2_X1 U7228 ( .A1(n5648), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n5651) );
  NAND2_X1 U7229 ( .A1(n5649), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n5650) );
  NOR2_X1 U7230 ( .A1(n9393), .A2(n5653), .ZN(n5789) );
  NOR2_X1 U7231 ( .A1(n9755), .A2(n9393), .ZN(n5658) );
  OAI21_X1 U7232 ( .B1(n4320), .B2(n9373), .A(n4861), .ZN(n5795) );
  INV_X1 U7233 ( .A(n6815), .ZN(n5720) );
  NOR2_X1 U7234 ( .A1(n9373), .A2(n6888), .ZN(n5719) );
  NAND2_X1 U7235 ( .A1(n5659), .A2(n5722), .ZN(n5710) );
  NAND2_X1 U7236 ( .A1(n5660), .A2(n8103), .ZN(n5700) );
  INV_X1 U7237 ( .A(n5661), .ZN(n5662) );
  NOR2_X1 U7238 ( .A1(n5700), .A2(n5662), .ZN(n5664) );
  INV_X1 U7239 ( .A(n9385), .ZN(n5663) );
  OR3_X1 U7240 ( .A1(n5664), .A2(n9388), .A3(n5663), .ZN(n5696) );
  INV_X1 U7241 ( .A(n5665), .ZN(n5666) );
  NOR4_X1 U7242 ( .A1(n5710), .A2(n5704), .A3(n5696), .A4(n5666), .ZN(n5788)
         );
  INV_X1 U7243 ( .A(n5667), .ZN(n5672) );
  AND2_X1 U7244 ( .A1(n7150), .A2(n7455), .ZN(n5742) );
  INV_X1 U7245 ( .A(n5742), .ZN(n5669) );
  NAND2_X1 U7246 ( .A1(n8082), .A2(n9274), .ZN(n5668) );
  NAND4_X1 U7247 ( .A1(n5670), .A2(n5669), .A3(n6814), .A4(n5668), .ZN(n5671)
         );
  NAND2_X1 U7248 ( .A1(n5672), .A2(n5671), .ZN(n5674) );
  AND3_X1 U7249 ( .A1(n5737), .A2(n5738), .A3(n5768), .ZN(n5673) );
  AOI22_X1 U7250 ( .A1(n5674), .A2(n5673), .B1(n5768), .B2(n4392), .ZN(n5679)
         );
  NAND3_X1 U7251 ( .A1(n7616), .A2(n5675), .A3(n7629), .ZN(n5676) );
  NAND2_X1 U7252 ( .A1(n5676), .A2(n7615), .ZN(n5750) );
  NOR2_X1 U7253 ( .A1(n5750), .A2(n5677), .ZN(n5770) );
  NAND2_X1 U7254 ( .A1(n5771), .A2(n5749), .ZN(n5678) );
  AOI21_X1 U7255 ( .B1(n5679), .B2(n5770), .A(n5678), .ZN(n5681) );
  AND2_X1 U7256 ( .A1(n5734), .A2(n9873), .ZN(n5774) );
  OAI21_X1 U7257 ( .B1(n5681), .B2(n5680), .A(n5774), .ZN(n5682) );
  NAND3_X1 U7258 ( .A1(n5682), .A2(n8017), .A3(n9614), .ZN(n5683) );
  AND2_X1 U7259 ( .A1(n5683), .A2(n5733), .ZN(n5686) );
  INV_X1 U7260 ( .A(n5684), .ZN(n5685) );
  AOI21_X1 U7261 ( .B1(n5686), .B2(n5777), .A(n5685), .ZN(n5687) );
  OAI21_X1 U7262 ( .B1(n5688), .B2(n5687), .A(n5780), .ZN(n5691) );
  INV_X1 U7263 ( .A(n5689), .ZN(n5690) );
  AOI21_X1 U7264 ( .B1(n5692), .B2(n5691), .A(n5690), .ZN(n5695) );
  INV_X1 U7265 ( .A(n5693), .ZN(n5694) );
  OAI21_X1 U7266 ( .B1(n5695), .B2(n5694), .A(n5785), .ZN(n5714) );
  NAND2_X1 U7267 ( .A1(n9381), .A2(n9393), .ZN(n5763) );
  INV_X1 U7268 ( .A(n5763), .ZN(n5713) );
  INV_X1 U7269 ( .A(n5696), .ZN(n5703) );
  INV_X1 U7270 ( .A(n8101), .ZN(n5699) );
  NAND2_X1 U7271 ( .A1(n5697), .A2(n5728), .ZN(n8099) );
  INV_X1 U7272 ( .A(n8099), .ZN(n5698) );
  OR3_X1 U7273 ( .A1(n5700), .A2(n5699), .A3(n5698), .ZN(n5702) );
  AOI21_X1 U7274 ( .B1(n5703), .B2(n5702), .A(n5701), .ZN(n5705) );
  NOR2_X1 U7275 ( .A1(n5705), .A2(n5704), .ZN(n5708) );
  INV_X1 U7276 ( .A(n5706), .ZN(n5707) );
  NOR2_X1 U7277 ( .A1(n5708), .A2(n5707), .ZN(n5709) );
  OR2_X1 U7278 ( .A1(n5710), .A2(n5709), .ZN(n5712) );
  NAND2_X1 U7279 ( .A1(n5712), .A2(n5711), .ZN(n5787) );
  AOI211_X1 U7280 ( .C1(n5788), .C2(n5714), .A(n5713), .B(n5787), .ZN(n5716)
         );
  OR2_X1 U7281 ( .A1(n9381), .A2(n9393), .ZN(n5764) );
  INV_X1 U7282 ( .A(n5764), .ZN(n5715) );
  NOR2_X1 U7283 ( .A1(n5716), .A2(n5715), .ZN(n5717) );
  OAI21_X1 U7284 ( .B1(n5717), .B2(n5790), .A(n4320), .ZN(n5718) );
  MUX2_X1 U7285 ( .A(n5720), .B(n5719), .S(n5718), .Z(n5794) );
  NAND2_X1 U7286 ( .A1(n7268), .A2(n6884), .ZN(n6891) );
  NAND2_X1 U7287 ( .A1(n5722), .A2(n9391), .ZN(n9415) );
  NOR2_X1 U7288 ( .A1(n9388), .A2(n5725), .ZN(n9463) );
  INV_X1 U7289 ( .A(n9565), .ZN(n9564) );
  NAND2_X1 U7290 ( .A1(n5731), .A2(n5780), .ZN(n9581) );
  NAND2_X1 U7291 ( .A1(n5732), .A2(n5779), .ZN(n9596) );
  NAND2_X1 U7292 ( .A1(n5734), .A2(n8017), .ZN(n9885) );
  NAND2_X1 U7293 ( .A1(n9873), .A2(n5735), .ZN(n7725) );
  NAND2_X1 U7294 ( .A1(n5767), .A2(n5768), .ZN(n7435) );
  NOR2_X1 U7295 ( .A1(n7435), .A2(n7333), .ZN(n5745) );
  NAND2_X1 U7296 ( .A1(n5739), .A2(n5738), .ZN(n7223) );
  INV_X1 U7297 ( .A(n7223), .ZN(n5744) );
  NAND2_X1 U7298 ( .A1(n5741), .A2(n5740), .ZN(n7218) );
  NOR2_X1 U7299 ( .A1(n7218), .A2(n6814), .ZN(n5743) );
  NOR2_X1 U7300 ( .A1(n7153), .A2(n5742), .ZN(n7264) );
  AND4_X1 U7301 ( .A1(n5745), .A2(n5744), .A3(n5743), .A4(n7264), .ZN(n5748)
         );
  NAND2_X1 U7302 ( .A1(n7504), .A2(n7503), .ZN(n7352) );
  NOR2_X1 U7303 ( .A1(n7145), .A2(n7352), .ZN(n5746) );
  NAND4_X1 U7304 ( .A1(n5748), .A2(n5747), .A3(n5746), .A4(n7616), .ZN(n5751)
         );
  NAND2_X1 U7305 ( .A1(n5749), .A2(n7723), .ZN(n7690) );
  OR3_X1 U7306 ( .A1(n5751), .A2(n7690), .A3(n5750), .ZN(n5752) );
  NOR3_X1 U7307 ( .A1(n9885), .A2(n7725), .A3(n5752), .ZN(n5753) );
  NAND2_X1 U7308 ( .A1(n8026), .A2(n5753), .ZN(n5754) );
  OR4_X1 U7309 ( .A1(n9581), .A2(n5755), .A3(n9596), .A4(n5754), .ZN(n5756) );
  NOR2_X1 U7310 ( .A1(n9564), .A2(n5756), .ZN(n5757) );
  NAND3_X1 U7311 ( .A1(n9539), .A2(n9552), .A3(n5757), .ZN(n5758) );
  NOR2_X1 U7312 ( .A1(n9527), .A2(n5758), .ZN(n5759) );
  AND4_X1 U7313 ( .A1(n9479), .A2(n4382), .A3(n9508), .A4(n5759), .ZN(n5760)
         );
  NAND4_X1 U7314 ( .A1(n9441), .A2(n9463), .A3(n8105), .A4(n5760), .ZN(n5761)
         );
  OR3_X1 U7315 ( .A1(n9415), .A2(n9428), .A3(n5761), .ZN(n5762) );
  NOR2_X1 U7316 ( .A1(n9403), .A2(n5762), .ZN(n5766) );
  AND2_X1 U7317 ( .A1(n5764), .A2(n5763), .ZN(n5765) );
  NAND4_X1 U7318 ( .A1(n5655), .A2(n4320), .A3(n5766), .A4(n5765), .ZN(n5791)
         );
  NAND2_X1 U7319 ( .A1(n7434), .A2(n5767), .ZN(n5769) );
  NAND2_X1 U7320 ( .A1(n5769), .A2(n5768), .ZN(n7506) );
  NAND2_X1 U7321 ( .A1(n7506), .A2(n5770), .ZN(n5772) );
  NAND2_X1 U7322 ( .A1(n7724), .A2(n5773), .ZN(n9874) );
  NAND2_X1 U7323 ( .A1(n9874), .A2(n5774), .ZN(n8020) );
  NAND2_X1 U7324 ( .A1(n8020), .A2(n8017), .ZN(n5775) );
  NAND2_X1 U7325 ( .A1(n5775), .A2(n8026), .ZN(n9615) );
  NAND2_X1 U7326 ( .A1(n5776), .A2(n9615), .ZN(n5778) );
  NAND2_X1 U7327 ( .A1(n5778), .A2(n5777), .ZN(n9597) );
  INV_X1 U7328 ( .A(n9581), .ZN(n9590) );
  NAND2_X1 U7329 ( .A1(n5786), .A2(n5785), .ZN(n9528) );
  INV_X4 U7330 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  OR2_X1 U7331 ( .A1(n6808), .A2(P1_U3086), .ZN(n7814) );
  INV_X1 U7332 ( .A(n6336), .ZN(n5808) );
  INV_X1 U7333 ( .A(n7902), .ZN(n5806) );
  INV_X1 U7334 ( .A(n6831), .ZN(n6824) );
  INV_X1 U7335 ( .A(n8084), .ZN(n6920) );
  NAND2_X1 U7336 ( .A1(n6920), .A2(n7148), .ZN(n6919) );
  INV_X1 U7337 ( .A(n7147), .ZN(n6804) );
  OR2_X1 U7338 ( .A1(n6815), .A2(n6804), .ZN(n6887) );
  NOR3_X1 U7339 ( .A1(n6824), .A2(n6919), .A3(n6887), .ZN(n5812) );
  OAI21_X1 U7340 ( .B1(n7814), .B2(n6884), .A(P1_B_REG_SCAN_IN), .ZN(n5811) );
  OR2_X1 U7341 ( .A1(n5812), .A2(n5811), .ZN(n5813) );
  OAI21_X1 U7342 ( .B1(n5814), .B2(n7814), .A(n5813), .ZN(P1_U3242) );
  NAND4_X1 U7343 ( .A1(n5815), .A2(n5962), .A3(n5961), .A4(n5993), .ZN(n5816)
         );
  INV_X1 U7344 ( .A(n5816), .ZN(n5817) );
  NOR2_X1 U7345 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(P2_IR_REG_13__SCAN_IN), .ZN(
        n5818) );
  NOR2_X1 U7346 ( .A1(P2_IR_REG_26__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), .ZN(
        n5821) );
  AND2_X1 U7347 ( .A1(n5828), .A2(n5821), .ZN(n5822) );
  NAND2_X1 U7348 ( .A1(n5824), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5823) );
  INV_X1 U7349 ( .A(n5828), .ZN(n5829) );
  NAND2_X1 U7350 ( .A1(n5829), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5830) );
  NAND2_X1 U7351 ( .A1(n5832), .A2(P2_IR_REG_27__SCAN_IN), .ZN(n5836) );
  INV_X1 U7352 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5831) );
  OAI21_X1 U7353 ( .B1(n5832), .B2(P2_IR_REG_27__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5833) );
  OAI21_X1 U7354 ( .B1(P2_IR_REG_31__SCAN_IN), .B2(P2_IR_REG_27__SCAN_IN), .A(
        n5833), .ZN(n5834) );
  INV_X1 U7355 ( .A(n5837), .ZN(n6272) );
  NAND2_X1 U7356 ( .A1(n7236), .A2(n8404), .ZN(n5840) );
  NAND2_X1 U7357 ( .A1(n8226), .A2(n6363), .ZN(n5948) );
  NAND2_X1 U7358 ( .A1(n5856), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5838) );
  XNOR2_X1 U7359 ( .A(n5838), .B(P2_IR_REG_16__SCAN_IN), .ZN(n10033) );
  AOI22_X1 U7360 ( .A1(n6128), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n6127), .B2(
        n10033), .ZN(n5839) );
  INV_X1 U7361 ( .A(P2_B_REG_SCAN_IN), .ZN(n5844) );
  XNOR2_X1 U7362 ( .A(n6238), .B(n5844), .ZN(n5848) );
  NAND2_X1 U7363 ( .A1(n5848), .A2(n8039), .ZN(n5853) );
  INV_X1 U7364 ( .A(n5850), .ZN(n5849) );
  NAND2_X1 U7365 ( .A1(n5850), .A2(P2_IR_REG_26__SCAN_IN), .ZN(n5851) );
  NAND2_X1 U7366 ( .A1(n5853), .A2(n6239), .ZN(n6224) );
  INV_X1 U7367 ( .A(n6224), .ZN(n5855) );
  INV_X1 U7368 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n5854) );
  INV_X1 U7369 ( .A(n6238), .ZN(n7950) );
  INV_X1 U7370 ( .A(n6094), .ZN(n5858) );
  NAND2_X1 U7371 ( .A1(n4324), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5861) );
  MUX2_X1 U7372 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5861), .S(
        P2_IR_REG_20__SCAN_IN), .Z(n5862) );
  NAND2_X1 U7373 ( .A1(n5860), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5863) );
  XNOR2_X1 U7374 ( .A(n4431), .B(n5951), .ZN(n6092) );
  INV_X1 U7375 ( .A(n6092), .ZN(n6093) );
  NAND2_X1 U7376 ( .A1(n5865), .A2(n5864), .ZN(n5869) );
  MUX2_X1 U7377 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5868), .S(
        P2_IR_REG_29__SCAN_IN), .Z(n5870) );
  INV_X2 U7378 ( .A(n6013), .ZN(n8229) );
  NAND2_X1 U7379 ( .A1(n8229), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n5882) );
  INV_X2 U7380 ( .A(n6017), .ZN(n8228) );
  NAND2_X1 U7381 ( .A1(n8228), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n5881) );
  AND2_X2 U7382 ( .A1(n5873), .A2(n5872), .ZN(n5986) );
  NOR2_X1 U7383 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n5967) );
  INV_X1 U7384 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n6682) );
  NAND2_X1 U7385 ( .A1(n5967), .A2(n6682), .ZN(n5999) );
  NOR2_X1 U7386 ( .A1(n6015), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n6014) );
  INV_X1 U7387 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5874) );
  NAND2_X1 U7388 ( .A1(n6028), .A2(n5874), .ZN(n6051) );
  INV_X1 U7389 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n5875) );
  NAND2_X1 U7390 ( .A1(n5902), .A2(n5875), .ZN(n6081) );
  INV_X1 U7391 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n5876) );
  INV_X1 U7392 ( .A(n6099), .ZN(n6100) );
  INV_X1 U7393 ( .A(n5877), .ZN(n5884) );
  NAND2_X1 U7394 ( .A1(n5884), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5878) );
  NAND2_X1 U7395 ( .A1(n6100), .A2(n5878), .ZN(n8869) );
  NAND2_X1 U7396 ( .A1(n6111), .A2(n8869), .ZN(n5880) );
  NAND2_X1 U7397 ( .A1(n6264), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n5879) );
  NAND4_X1 U7398 ( .A1(n5882), .A2(n5881), .A3(n5880), .A4(n5879), .ZN(n8608)
         );
  NAND2_X1 U7399 ( .A1(n8229), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n5888) );
  NAND2_X1 U7400 ( .A1(n6083), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5883) );
  NAND2_X1 U7401 ( .A1(n5884), .A2(n5883), .ZN(n8599) );
  NAND2_X1 U7402 ( .A1(n6111), .A2(n8599), .ZN(n5887) );
  NAND2_X1 U7403 ( .A1(n6264), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n5886) );
  INV_X1 U7404 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n8643) );
  OR2_X1 U7405 ( .A1(n6017), .A2(n8643), .ZN(n5885) );
  NAND2_X1 U7406 ( .A1(n7141), .A2(n8404), .ZN(n5898) );
  INV_X1 U7407 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n5890) );
  NAND2_X1 U7408 ( .A1(n5889), .A2(n5890), .ZN(n6025) );
  NOR2_X1 U7409 ( .A1(n6025), .A2(P2_IR_REG_9__SCAN_IN), .ZN(n6058) );
  NAND2_X1 U7410 ( .A1(n6058), .A2(n6059), .ZN(n6061) );
  NAND2_X1 U7411 ( .A1(n5891), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5899) );
  INV_X1 U7412 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5892) );
  NAND2_X1 U7413 ( .A1(n5899), .A2(n5892), .ZN(n5893) );
  NAND2_X1 U7414 ( .A1(n5893), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6078) );
  INV_X1 U7415 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5894) );
  NAND2_X1 U7416 ( .A1(n6078), .A2(n5894), .ZN(n5895) );
  NAND2_X1 U7417 ( .A1(n5895), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5896) );
  AOI22_X1 U7418 ( .A1(n6128), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n6127), .B2(
        n10017), .ZN(n5897) );
  XNOR2_X1 U7419 ( .A(n8588), .B(n5951), .ZN(n6090) );
  INV_X1 U7420 ( .A(n6090), .ZN(n6091) );
  XNOR2_X1 U7421 ( .A(n5899), .B(P2_IR_REG_13__SCAN_IN), .ZN(n9984) );
  AOI22_X1 U7422 ( .A1(n6128), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6127), .B2(
        n9984), .ZN(n5900) );
  XNOR2_X1 U7423 ( .A(n7822), .B(n5951), .ZN(n6077) );
  NAND2_X1 U7424 ( .A1(n8228), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n5907) );
  NAND2_X1 U7425 ( .A1(n8229), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n5906) );
  INV_X1 U7426 ( .A(n5902), .ZN(n6071) );
  NAND2_X1 U7427 ( .A1(n6071), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n5903) );
  NAND2_X1 U7428 ( .A1(n6081), .A2(n5903), .ZN(n7969) );
  NAND2_X1 U7429 ( .A1(n6111), .A2(n7969), .ZN(n5905) );
  NAND2_X1 U7430 ( .A1(n6264), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5904) );
  NAND4_X1 U7431 ( .A1(n5907), .A2(n5906), .A3(n5905), .A4(n5904), .ZN(n8611)
         );
  NAND2_X1 U7432 ( .A1(n8228), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n5912) );
  NAND2_X1 U7433 ( .A1(n8229), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n5911) );
  NAND2_X1 U7434 ( .A1(n6053), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5908) );
  NAND2_X1 U7435 ( .A1(n6069), .A2(n5908), .ZN(n7835) );
  NAND2_X1 U7436 ( .A1(n6111), .A2(n7835), .ZN(n5910) );
  NAND2_X1 U7437 ( .A1(n6264), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5909) );
  NAND2_X1 U7438 ( .A1(n5913), .A2(n8404), .ZN(n5917) );
  NAND2_X1 U7439 ( .A1(n6061), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5914) );
  MUX2_X1 U7440 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5914), .S(
        P2_IR_REG_11__SCAN_IN), .Z(n5915) );
  AOI22_X1 U7441 ( .A1(n6128), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n6127), .B2(
        n7492), .ZN(n5916) );
  OR2_X1 U7442 ( .A1(n7844), .A2(n8613), .ZN(n7710) );
  NAND2_X1 U7443 ( .A1(n7844), .A2(n8613), .ZN(n7711) );
  XNOR2_X1 U7444 ( .A(n8433), .B(n6297), .ZN(n7840) );
  NAND2_X1 U7445 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5918) );
  MUX2_X1 U7446 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5918), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n5920) );
  INV_X1 U7447 ( .A(n5937), .ZN(n5919) );
  NAND2_X1 U7448 ( .A1(n5920), .A2(n5919), .ZN(n6608) );
  INV_X1 U7449 ( .A(n6608), .ZN(n6597) );
  OR2_X1 U7450 ( .A1(n5948), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n5921) );
  INV_X2 U7451 ( .A(n6017), .ZN(n5998) );
  NAND2_X1 U7452 ( .A1(n5998), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n5926) );
  NAND2_X1 U7453 ( .A1(n5986), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n5924) );
  NAND2_X1 U7454 ( .A1(n6193), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5923) );
  XNOR2_X1 U7455 ( .A(n5934), .B(n8624), .ZN(n6960) );
  INV_X1 U7456 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n5927) );
  NAND2_X1 U7457 ( .A1(n5986), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n5930) );
  NAND2_X1 U7458 ( .A1(n6193), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5929) );
  NAND2_X1 U7459 ( .A1(n5998), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5928) );
  NAND2_X1 U7460 ( .A1(n6364), .A2(SI_0_), .ZN(n5932) );
  XNOR2_X1 U7461 ( .A(n5932), .B(n4516), .ZN(n9024) );
  MUX2_X1 U7462 ( .A(n4712), .B(n9024), .S(n8226), .Z(n7048) );
  AND2_X1 U7463 ( .A1(n5951), .A2(n7048), .ZN(n5933) );
  NAND2_X1 U7464 ( .A1(n6960), .A2(n6961), .ZN(n5936) );
  INV_X1 U7465 ( .A(n8624), .ZN(n7162) );
  NAND2_X1 U7466 ( .A1(n5934), .A2(n7162), .ZN(n5935) );
  NAND2_X1 U7467 ( .A1(n5936), .A2(n5935), .ZN(n6967) );
  OR2_X1 U7468 ( .A1(n5948), .A2(n4776), .ZN(n5941) );
  OR2_X1 U7469 ( .A1(n5964), .A2(n8078), .ZN(n5940) );
  OR2_X1 U7470 ( .A1(n8226), .A2(n4316), .ZN(n5939) );
  INV_X1 U7471 ( .A(n10097), .ZN(n7241) );
  NAND2_X1 U7472 ( .A1(n5986), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n5945) );
  NAND2_X1 U7473 ( .A1(n6264), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5944) );
  NAND2_X1 U7474 ( .A1(n8228), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n5943) );
  NAND2_X1 U7475 ( .A1(n6193), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5942) );
  AND4_X2 U7476 ( .A1(n5945), .A2(n5944), .A3(n5943), .A4(n5942), .ZN(n7242)
         );
  XNOR2_X1 U7477 ( .A(n5957), .B(n7242), .ZN(n6966) );
  NAND2_X1 U7478 ( .A1(n6967), .A2(n6966), .ZN(n7077) );
  OR2_X1 U7479 ( .A1(n5946), .A2(n5826), .ZN(n5947) );
  XNOR2_X1 U7480 ( .A(n5947), .B(n5961), .ZN(n6626) );
  OR2_X1 U7481 ( .A1(n5948), .A2(n4430), .ZN(n5950) );
  OR2_X1 U7482 ( .A1(n5964), .A2(n6365), .ZN(n5949) );
  OAI211_X1 U7483 ( .C1(n8226), .C2(n6626), .A(n5950), .B(n5949), .ZN(n7247)
         );
  XNOR2_X1 U7484 ( .A(n5951), .B(n7072), .ZN(n5973) );
  INV_X1 U7485 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n5952) );
  NAND2_X1 U7486 ( .A1(n5986), .A2(n5952), .ZN(n5956) );
  NAND2_X1 U7487 ( .A1(n5998), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n5955) );
  NAND2_X1 U7488 ( .A1(n6264), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5954) );
  NAND2_X1 U7489 ( .A1(n6193), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5953) );
  XNOR2_X1 U7490 ( .A(n5973), .B(n7315), .ZN(n7080) );
  INV_X1 U7491 ( .A(n7080), .ZN(n5959) );
  INV_X1 U7492 ( .A(n5957), .ZN(n5958) );
  NAND2_X1 U7493 ( .A1(n5958), .A2(n7242), .ZN(n7076) );
  NAND2_X1 U7494 ( .A1(n7077), .A2(n5960), .ZN(n6847) );
  NAND2_X1 U7495 ( .A1(n5946), .A2(n5961), .ZN(n5979) );
  NAND2_X1 U7496 ( .A1(n5979), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5963) );
  XNOR2_X1 U7497 ( .A(n5963), .B(n5962), .ZN(n6676) );
  OR2_X1 U7498 ( .A1(n5964), .A2(n6367), .ZN(n5966) );
  INV_X1 U7499 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6366) );
  NAND2_X1 U7500 ( .A1(n5998), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5972) );
  NAND2_X1 U7501 ( .A1(n8229), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5971) );
  INV_X1 U7502 ( .A(n5967), .ZN(n5984) );
  NAND2_X1 U7503 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n5968) );
  NAND2_X1 U7504 ( .A1(n5984), .A2(n5968), .ZN(n7381) );
  NAND2_X1 U7505 ( .A1(n5986), .A2(n7381), .ZN(n5970) );
  NAND2_X1 U7506 ( .A1(n6264), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n5969) );
  INV_X1 U7507 ( .A(n5973), .ZN(n5974) );
  NAND2_X1 U7508 ( .A1(n5974), .A2(n8621), .ZN(n6848) );
  INV_X1 U7509 ( .A(n6848), .ZN(n5975) );
  NOR2_X1 U7510 ( .A1(n6852), .A2(n5975), .ZN(n5976) );
  NAND2_X1 U7511 ( .A1(n5977), .A2(n7319), .ZN(n5978) );
  OR2_X1 U7512 ( .A1(n6370), .A2(n5964), .ZN(n5983) );
  NAND2_X1 U7513 ( .A1(n5992), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5980) );
  XNOR2_X1 U7514 ( .A(n5980), .B(n5993), .ZN(n6789) );
  OR2_X1 U7515 ( .A1(n8226), .A2(n6789), .ZN(n5981) );
  XNOR2_X1 U7516 ( .A(n5951), .B(n10112), .ZN(n5991) );
  NAND2_X1 U7517 ( .A1(n5998), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n5990) );
  NAND2_X1 U7518 ( .A1(n8229), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n5989) );
  NAND2_X1 U7519 ( .A1(n5984), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5985) );
  NAND2_X1 U7520 ( .A1(n5999), .A2(n5985), .ZN(n7325) );
  NAND2_X1 U7521 ( .A1(n5986), .A2(n7325), .ZN(n5988) );
  NAND2_X1 U7522 ( .A1(n6264), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5987) );
  XNOR2_X1 U7523 ( .A(n5991), .B(n8619), .ZN(n6954) );
  INV_X1 U7524 ( .A(n5992), .ZN(n5994) );
  NAND2_X1 U7525 ( .A1(n5994), .A2(n5993), .ZN(n6007) );
  NAND2_X1 U7526 ( .A1(n6007), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5995) );
  XNOR2_X1 U7527 ( .A(n5995), .B(P2_IR_REG_6__SCAN_IN), .ZN(n6796) );
  AOI22_X1 U7528 ( .A1(n6128), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n6127), .B2(
        n6796), .ZN(n5996) );
  XNOR2_X1 U7529 ( .A(n5951), .B(n7393), .ZN(n6005) );
  NAND2_X1 U7530 ( .A1(n5998), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n6004) );
  NAND2_X1 U7531 ( .A1(n8229), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6003) );
  NAND2_X1 U7532 ( .A1(n5999), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n6000) );
  NAND2_X1 U7533 ( .A1(n6015), .A2(n6000), .ZN(n7372) );
  NAND2_X1 U7534 ( .A1(n6111), .A2(n7372), .ZN(n6002) );
  NAND2_X1 U7535 ( .A1(n6264), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n6001) );
  AND4_X2 U7536 ( .A1(n6004), .A2(n6003), .A3(n6002), .A4(n6001), .ZN(n10077)
         );
  XNOR2_X1 U7537 ( .A(n6005), .B(n10077), .ZN(n7028) );
  INV_X1 U7538 ( .A(n10077), .ZN(n8618) );
  NAND2_X1 U7539 ( .A1(n6005), .A2(n8618), .ZN(n6006) );
  OAI21_X1 U7540 ( .B1(n6007), .B2(P2_IR_REG_6__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n6008) );
  MUX2_X1 U7541 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6008), .S(
        P2_IR_REG_7__SCAN_IN), .Z(n6010) );
  INV_X1 U7542 ( .A(n5889), .ZN(n6009) );
  AOI22_X1 U7543 ( .A1(n6128), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n6127), .B2(
        n6995), .ZN(n6011) );
  XNOR2_X1 U7544 ( .A(n10125), .B(n6297), .ZN(n6023) );
  NAND2_X1 U7545 ( .A1(n8409), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6021) );
  INV_X1 U7546 ( .A(n6014), .ZN(n6034) );
  NAND2_X1 U7547 ( .A1(n6015), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n6016) );
  NAND2_X1 U7548 ( .A1(n6034), .A2(n6016), .ZN(n10088) );
  NAND2_X1 U7549 ( .A1(n6111), .A2(n10088), .ZN(n6020) );
  NAND2_X1 U7550 ( .A1(n6264), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n6019) );
  NAND2_X1 U7551 ( .A1(n5998), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n6018) );
  XNOR2_X1 U7552 ( .A(n6023), .B(n7396), .ZN(n7210) );
  NAND2_X1 U7553 ( .A1(n6023), .A2(n7396), .ZN(n6024) );
  NAND2_X1 U7554 ( .A1(n6025), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6026) );
  XNOR2_X1 U7555 ( .A(n6026), .B(P2_IR_REG_9__SCAN_IN), .ZN(n7177) );
  AOI22_X1 U7556 ( .A1(n6128), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6127), .B2(
        n7177), .ZN(n6027) );
  XNOR2_X1 U7557 ( .A(n10134), .B(n6297), .ZN(n7577) );
  NAND2_X1 U7558 ( .A1(n8229), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n6033) );
  NAND2_X1 U7559 ( .A1(n6264), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n6032) );
  INV_X1 U7560 ( .A(n6028), .ZN(n6036) );
  NAND2_X1 U7561 ( .A1(n6036), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n6029) );
  NAND2_X1 U7562 ( .A1(n6051), .A2(n6029), .ZN(n7665) );
  NAND2_X1 U7563 ( .A1(n6111), .A2(n7665), .ZN(n6031) );
  NAND2_X1 U7564 ( .A1(n8228), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n6030) );
  NAND2_X1 U7565 ( .A1(n8228), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n6040) );
  NAND2_X1 U7566 ( .A1(n8229), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n6039) );
  NAND2_X1 U7567 ( .A1(n6034), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n6035) );
  NAND2_X1 U7568 ( .A1(n6036), .A2(n6035), .ZN(n7428) );
  NAND2_X1 U7569 ( .A1(n6111), .A2(n7428), .ZN(n6038) );
  NAND2_X1 U7570 ( .A1(n6264), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n6037) );
  NAND2_X1 U7571 ( .A1(n6399), .A2(n8404), .ZN(n6043) );
  OR2_X1 U7572 ( .A1(n5889), .A2(n5826), .ZN(n6041) );
  XNOR2_X1 U7573 ( .A(n6041), .B(P2_IR_REG_8__SCAN_IN), .ZN(n7118) );
  AOI22_X1 U7574 ( .A1(n6128), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n6127), .B2(
        n7118), .ZN(n6042) );
  NAND2_X1 U7575 ( .A1(n6043), .A2(n6042), .ZN(n7658) );
  XNOR2_X1 U7576 ( .A(n7658), .B(n6297), .ZN(n6046) );
  AOI22_X1 U7577 ( .A1(n7577), .A2(n7675), .B1(n10075), .B2(n6046), .ZN(n6050)
         );
  INV_X1 U7578 ( .A(n7577), .ZN(n6045) );
  OAI21_X1 U7579 ( .B1(n6046), .B2(n10075), .A(n7675), .ZN(n6044) );
  NAND2_X1 U7580 ( .A1(n6045), .A2(n6044), .ZN(n6048) );
  INV_X1 U7581 ( .A(n6046), .ZN(n7575) );
  NAND3_X1 U7582 ( .A1(n7575), .A2(n8616), .A3(n8615), .ZN(n6047) );
  NAND2_X1 U7583 ( .A1(n6048), .A2(n6047), .ZN(n6049) );
  NAND2_X1 U7584 ( .A1(n8228), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n6057) );
  NAND2_X1 U7585 ( .A1(n8229), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n6056) );
  NAND2_X1 U7586 ( .A1(n6051), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n6052) );
  NAND2_X1 U7587 ( .A1(n6053), .A2(n6052), .ZN(n7680) );
  NAND2_X1 U7588 ( .A1(n6111), .A2(n7680), .ZN(n6055) );
  NAND2_X1 U7589 ( .A1(n6264), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n6054) );
  OR2_X1 U7590 ( .A1(n6603), .A2(n5964), .ZN(n6064) );
  OR2_X1 U7591 ( .A1(n6058), .A2(n5826), .ZN(n6060) );
  MUX2_X1 U7592 ( .A(n6060), .B(P2_IR_REG_31__SCAN_IN), .S(n6059), .Z(n6062)
         );
  AOI22_X1 U7593 ( .A1(n6128), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6127), .B2(
        n7280), .ZN(n6063) );
  XNOR2_X1 U7594 ( .A(n10140), .B(n5951), .ZN(n7606) );
  OR2_X1 U7595 ( .A1(n6768), .A2(n5964), .ZN(n6068) );
  NAND2_X1 U7596 ( .A1(n6065), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6066) );
  XNOR2_X1 U7597 ( .A(n6066), .B(P2_IR_REG_12__SCAN_IN), .ZN(n7488) );
  AOI22_X1 U7598 ( .A1(n6128), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6127), .B2(
        n7488), .ZN(n6067) );
  XNOR2_X1 U7599 ( .A(n8312), .B(n5951), .ZN(n6076) );
  NAND2_X1 U7600 ( .A1(n8409), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n6075) );
  NAND2_X1 U7601 ( .A1(n8228), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n6074) );
  NAND2_X1 U7602 ( .A1(n6069), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n6070) );
  NAND2_X1 U7603 ( .A1(n6071), .A2(n6070), .ZN(n7889) );
  NAND2_X1 U7604 ( .A1(n6111), .A2(n7889), .ZN(n6073) );
  NAND2_X1 U7605 ( .A1(n6264), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n6072) );
  NAND4_X1 U7606 ( .A1(n6075), .A2(n6074), .A3(n6073), .A4(n6072), .ZN(n8612)
         );
  INV_X1 U7607 ( .A(n8612), .ZN(n8311) );
  XNOR2_X1 U7608 ( .A(n6076), .B(n8311), .ZN(n7883) );
  INV_X1 U7609 ( .A(n8611), .ZN(n8045) );
  XNOR2_X1 U7610 ( .A(n6077), .B(n8045), .ZN(n7965) );
  NAND2_X1 U7611 ( .A1(n6896), .A2(n8404), .ZN(n6080) );
  XNOR2_X1 U7612 ( .A(n6078), .B(P2_IR_REG_14__SCAN_IN), .ZN(n10002) );
  AOI22_X1 U7613 ( .A1(n6128), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n6127), .B2(
        n10002), .ZN(n6079) );
  XNOR2_X1 U7614 ( .A(n8047), .B(n5951), .ZN(n6088) );
  NAND2_X1 U7615 ( .A1(n8228), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n6087) );
  NAND2_X1 U7616 ( .A1(n8409), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n6086) );
  NAND2_X1 U7617 ( .A1(n6081), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n6082) );
  NAND2_X1 U7618 ( .A1(n6083), .A2(n6082), .ZN(n8042) );
  NAND2_X1 U7619 ( .A1(n6111), .A2(n8042), .ZN(n6085) );
  NAND2_X1 U7620 ( .A1(n6264), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n6084) );
  XNOR2_X1 U7621 ( .A(n6088), .B(n8596), .ZN(n8041) );
  INV_X1 U7622 ( .A(n6088), .ZN(n6089) );
  XNOR2_X1 U7623 ( .A(n6090), .B(n8863), .ZN(n8591) );
  XNOR2_X1 U7624 ( .A(n6092), .B(n8608), .ZN(n8521) );
  NAND2_X1 U7625 ( .A1(n7293), .A2(n8404), .ZN(n6098) );
  NAND2_X1 U7626 ( .A1(n6094), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6095) );
  MUX2_X1 U7627 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6095), .S(
        P2_IR_REG_17__SCAN_IN), .Z(n6096) );
  INV_X1 U7628 ( .A(n8678), .ZN(n10050) );
  AOI22_X1 U7629 ( .A1(n6128), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n6127), .B2(
        n10050), .ZN(n6097) );
  XNOR2_X1 U7630 ( .A(n8998), .B(n6297), .ZN(n6106) );
  NAND2_X1 U7631 ( .A1(n8228), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n6105) );
  NAND2_X1 U7632 ( .A1(n8409), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n6104) );
  NAND2_X1 U7633 ( .A1(n6100), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n6101) );
  NAND2_X1 U7634 ( .A1(n6109), .A2(n6101), .ZN(n8856) );
  NAND2_X1 U7635 ( .A1(n6111), .A2(n8856), .ZN(n6103) );
  NAND2_X1 U7636 ( .A1(n6264), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n6102) );
  NAND2_X1 U7637 ( .A1(n6106), .A2(n8864), .ZN(n8527) );
  INV_X1 U7638 ( .A(n6106), .ZN(n6107) );
  NAND2_X1 U7639 ( .A1(n6107), .A2(n8839), .ZN(n8528) );
  NAND2_X1 U7640 ( .A1(n5998), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n6115) );
  NAND2_X1 U7641 ( .A1(n6109), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n6110) );
  NAND2_X1 U7642 ( .A1(n6122), .A2(n6110), .ZN(n8845) );
  NAND2_X1 U7643 ( .A1(n8845), .A2(n6111), .ZN(n6114) );
  NAND2_X1 U7644 ( .A1(n8409), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n6113) );
  NAND2_X1 U7645 ( .A1(n6264), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n6112) );
  NAND2_X1 U7646 ( .A1(n7385), .A2(n8404), .ZN(n6120) );
  MUX2_X1 U7647 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6116), .S(
        P2_IR_REG_18__SCAN_IN), .Z(n6118) );
  AOI22_X1 U7648 ( .A1(n6128), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6127), .B2(
        n8688), .ZN(n6119) );
  XNOR2_X1 U7649 ( .A(n8992), .B(n5951), .ZN(n6121) );
  XOR2_X1 U7650 ( .A(n8852), .B(n6121), .Z(n8567) );
  INV_X1 U7651 ( .A(n6133), .ZN(n6134) );
  NAND2_X1 U7652 ( .A1(n6122), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n6123) );
  NAND2_X1 U7653 ( .A1(n6134), .A2(n6123), .ZN(n8829) );
  NAND2_X1 U7654 ( .A1(n8829), .A2(n6111), .ZN(n6126) );
  AOI22_X1 U7655 ( .A1(n5998), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n6193), .B2(
        P2_REG1_REG_19__SCAN_IN), .ZN(n6125) );
  NAND2_X1 U7656 ( .A1(n6264), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n6124) );
  NAND2_X1 U7657 ( .A1(n7472), .A2(n8404), .ZN(n6130) );
  AOI22_X1 U7658 ( .A1(n6128), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n8455), .B2(
        n6127), .ZN(n6129) );
  XOR2_X1 U7659 ( .A(n5951), .B(n8986), .Z(n6131) );
  INV_X1 U7660 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n6132) );
  INV_X1 U7661 ( .A(n6145), .ZN(n6146) );
  NAND2_X1 U7662 ( .A1(n6134), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n6135) );
  NAND2_X1 U7663 ( .A1(n6146), .A2(n6135), .ZN(n8812) );
  NAND2_X1 U7664 ( .A1(n8812), .A2(n6111), .ZN(n6138) );
  AOI22_X1 U7665 ( .A1(n6264), .A2(P2_REG0_REG_20__SCAN_IN), .B1(n6193), .B2(
        P2_REG1_REG_20__SCAN_IN), .ZN(n6137) );
  NAND2_X1 U7666 ( .A1(n5998), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n6136) );
  NAND2_X1 U7667 ( .A1(n7524), .A2(n8404), .ZN(n6140) );
  INV_X1 U7668 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7587) );
  OR2_X1 U7669 ( .A1(n5948), .A2(n7587), .ZN(n6139) );
  XNOR2_X1 U7670 ( .A(n8913), .B(n5951), .ZN(n6141) );
  NOR2_X1 U7671 ( .A1(n6141), .A2(n8826), .ZN(n8502) );
  AOI21_X1 U7672 ( .B1(n8826), .B2(n6141), .A(n8502), .ZN(n8547) );
  NAND2_X1 U7673 ( .A1(n7700), .A2(n8404), .ZN(n6143) );
  OR2_X1 U7674 ( .A1(n8402), .A2(n7703), .ZN(n6142) );
  XNOR2_X1 U7675 ( .A(n8979), .B(n6297), .ZN(n6151) );
  INV_X1 U7676 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n6144) );
  NAND2_X1 U7677 ( .A1(n6146), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n6147) );
  NAND2_X1 U7678 ( .A1(n6157), .A2(n6147), .ZN(n8804) );
  INV_X1 U7679 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n8978) );
  NAND2_X1 U7680 ( .A1(n8409), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n6149) );
  NAND2_X1 U7681 ( .A1(n5998), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n6148) );
  OAI211_X1 U7682 ( .C1(n8978), .C2(n8412), .A(n6149), .B(n6148), .ZN(n6150)
         );
  AOI21_X1 U7683 ( .B1(n8804), .B2(n6111), .A(n6150), .ZN(n8560) );
  NAND2_X1 U7684 ( .A1(n6151), .A2(n8560), .ZN(n6154) );
  INV_X1 U7685 ( .A(n6151), .ZN(n6152) );
  NAND2_X1 U7686 ( .A1(n6152), .A2(n8810), .ZN(n6153) );
  AND2_X1 U7687 ( .A1(n6154), .A2(n6153), .ZN(n8501) );
  NAND2_X1 U7688 ( .A1(n7800), .A2(n8404), .ZN(n6156) );
  OR2_X1 U7689 ( .A1(n5948), .A2(n7801), .ZN(n6155) );
  XNOR2_X1 U7690 ( .A(n8973), .B(n5951), .ZN(n6164) );
  NAND2_X1 U7691 ( .A1(n6157), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6158) );
  NAND2_X1 U7692 ( .A1(n6170), .A2(n6158), .ZN(n8791) );
  NAND2_X1 U7693 ( .A1(n8791), .A2(n6111), .ZN(n6163) );
  INV_X1 U7694 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n8972) );
  NAND2_X1 U7695 ( .A1(n8229), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n6160) );
  NAND2_X1 U7696 ( .A1(n8228), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n6159) );
  OAI211_X1 U7697 ( .C1(n8972), .C2(n8412), .A(n6160), .B(n6159), .ZN(n6161)
         );
  INV_X1 U7698 ( .A(n6161), .ZN(n6162) );
  XNOR2_X1 U7699 ( .A(n6164), .B(n8801), .ZN(n8557) );
  NAND2_X1 U7700 ( .A1(n8556), .A2(n8557), .ZN(n8555) );
  NAND2_X1 U7701 ( .A1(n8555), .A2(n6165), .ZN(n6169) );
  NAND2_X1 U7702 ( .A1(n7817), .A2(n8404), .ZN(n6167) );
  OR2_X1 U7703 ( .A1(n8402), .A2(n7820), .ZN(n6166) );
  XNOR2_X1 U7704 ( .A(n8970), .B(n5951), .ZN(n6168) );
  INV_X1 U7705 ( .A(n6179), .ZN(n6180) );
  NAND2_X1 U7706 ( .A1(n6170), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6171) );
  NAND2_X1 U7707 ( .A1(n6180), .A2(n6171), .ZN(n8777) );
  NAND2_X1 U7708 ( .A1(n8777), .A2(n5986), .ZN(n6176) );
  INV_X1 U7709 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n8967) );
  NAND2_X1 U7710 ( .A1(n8228), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n6173) );
  NAND2_X1 U7711 ( .A1(n8409), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n6172) );
  OAI211_X1 U7712 ( .C1(n8967), .C2(n8412), .A(n6173), .B(n6172), .ZN(n6174)
         );
  INV_X1 U7713 ( .A(n6174), .ZN(n6175) );
  NAND2_X1 U7714 ( .A1(n7900), .A2(n8404), .ZN(n6178) );
  OR2_X1 U7715 ( .A1(n5948), .A2(n7948), .ZN(n6177) );
  XNOR2_X1 U7716 ( .A(n8962), .B(n6297), .ZN(n6185) );
  INV_X1 U7717 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n8542) );
  NAND2_X1 U7718 ( .A1(n6179), .A2(n8542), .ZN(n6191) );
  NAND2_X1 U7719 ( .A1(n6180), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n6181) );
  NAND2_X1 U7720 ( .A1(n6191), .A2(n6181), .ZN(n8767) );
  INV_X1 U7721 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n8961) );
  NAND2_X1 U7722 ( .A1(n5998), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n6183) );
  NAND2_X1 U7723 ( .A1(n8409), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n6182) );
  OAI211_X1 U7724 ( .C1(n8961), .C2(n8412), .A(n6183), .B(n6182), .ZN(n6184)
         );
  NAND2_X1 U7725 ( .A1(n6185), .A2(n8774), .ZN(n6188) );
  INV_X1 U7726 ( .A(n6185), .ZN(n6186) );
  INV_X1 U7727 ( .A(n8774), .ZN(n8606) );
  NAND2_X1 U7728 ( .A1(n6186), .A2(n8606), .ZN(n6187) );
  AND2_X1 U7729 ( .A1(n6188), .A2(n6187), .ZN(n8537) );
  NAND2_X1 U7730 ( .A1(n8539), .A2(n6188), .ZN(n8510) );
  NAND2_X1 U7731 ( .A1(n8035), .A2(n8404), .ZN(n6190) );
  OR2_X1 U7732 ( .A1(n8402), .A2(n8037), .ZN(n6189) );
  XNOR2_X1 U7733 ( .A(n8201), .B(n5951), .ZN(n6199) );
  NAND2_X1 U7734 ( .A1(n6191), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n6192) );
  NAND2_X1 U7735 ( .A1(n6203), .A2(n6192), .ZN(n8513) );
  NAND2_X1 U7736 ( .A1(n8513), .A2(n6111), .ZN(n6198) );
  INV_X1 U7737 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n6561) );
  NAND2_X1 U7738 ( .A1(n8228), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n6195) );
  NAND2_X1 U7739 ( .A1(n6264), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n6194) );
  OAI211_X1 U7740 ( .C1(n6013), .C2(n6561), .A(n6195), .B(n6194), .ZN(n6196)
         );
  INV_X1 U7741 ( .A(n6196), .ZN(n6197) );
  XNOR2_X1 U7742 ( .A(n6199), .B(n8765), .ZN(n8511) );
  NAND2_X1 U7743 ( .A1(n8510), .A2(n8511), .ZN(n8509) );
  NAND2_X1 U7744 ( .A1(n8509), .A2(n6200), .ZN(n6212) );
  NAND2_X1 U7745 ( .A1(n8065), .A2(n8404), .ZN(n6202) );
  OR2_X1 U7746 ( .A1(n5948), .A2(n8066), .ZN(n6201) );
  XNOR2_X1 U7747 ( .A(n8950), .B(n5951), .ZN(n6210) );
  NAND2_X1 U7748 ( .A1(n6203), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n6204) );
  NAND2_X1 U7749 ( .A1(n6216), .A2(n6204), .ZN(n8745) );
  NAND2_X1 U7750 ( .A1(n8745), .A2(n5986), .ZN(n6209) );
  INV_X1 U7751 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n8949) );
  NAND2_X1 U7752 ( .A1(n8228), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n6206) );
  NAND2_X1 U7753 ( .A1(n8409), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n6205) );
  OAI211_X1 U7754 ( .C1(n8949), .C2(n8412), .A(n6206), .B(n6205), .ZN(n6207)
         );
  INV_X1 U7755 ( .A(n6207), .ZN(n6208) );
  INV_X1 U7756 ( .A(n6255), .ZN(n8577) );
  INV_X1 U7757 ( .A(n6210), .ZN(n6211) );
  AND2_X1 U7758 ( .A1(n6212), .A2(n6211), .ZN(n6251) );
  NAND2_X1 U7759 ( .A1(n8072), .A2(n8404), .ZN(n6215) );
  XNOR2_X1 U7760 ( .A(n8944), .B(n6297), .ZN(n6308) );
  INV_X1 U7761 ( .A(n6260), .ZN(n6261) );
  NAND2_X1 U7762 ( .A1(n6216), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n6217) );
  NAND2_X1 U7763 ( .A1(n6261), .A2(n6217), .ZN(n8735) );
  NAND2_X1 U7764 ( .A1(n8735), .A2(n6111), .ZN(n6222) );
  INV_X1 U7765 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n8943) );
  NAND2_X1 U7766 ( .A1(n5998), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n6219) );
  NAND2_X1 U7767 ( .A1(n8409), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n6218) );
  OAI211_X1 U7768 ( .C1(n8943), .C2(n8412), .A(n6219), .B(n6218), .ZN(n6220)
         );
  INV_X1 U7769 ( .A(n6220), .ZN(n6221) );
  XNOR2_X1 U7770 ( .A(n6308), .B(n8583), .ZN(n6252) );
  OAI21_X1 U7771 ( .B1(n8577), .B2(n6251), .A(n6252), .ZN(n6256) );
  NAND2_X1 U7772 ( .A1(n8039), .A2(n8067), .ZN(n6376) );
  NAND2_X1 U7773 ( .A1(n6223), .A2(n7037), .ZN(n7043) );
  NOR2_X1 U7774 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .ZN(
        n6229) );
  NOR4_X1 U7775 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_18__SCAN_IN), .ZN(n6228) );
  NOR4_X1 U7776 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_26__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n6227) );
  NOR4_X1 U7777 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_22__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n6226) );
  NAND4_X1 U7778 ( .A1(n6229), .A2(n6228), .A3(n6227), .A4(n6226), .ZN(n6235)
         );
  NOR4_X1 U7779 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_21__SCAN_IN), .ZN(n6233) );
  NOR4_X1 U7780 ( .A1(P2_D_REG_25__SCAN_IN), .A2(P2_D_REG_24__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_17__SCAN_IN), .ZN(n6232) );
  NOR4_X1 U7781 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n6231) );
  NOR4_X1 U7782 ( .A1(P2_D_REG_8__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_19__SCAN_IN), .ZN(n6230) );
  NAND4_X1 U7783 ( .A1(n6233), .A2(n6232), .A3(n6231), .A4(n6230), .ZN(n6234)
         );
  NOR2_X1 U7784 ( .A1(n6235), .A2(n6234), .ZN(n6236) );
  NOR2_X1 U7785 ( .A1(n7043), .A2(n7041), .ZN(n6276) );
  NAND2_X1 U7786 ( .A1(n6244), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6245) );
  NAND2_X1 U7787 ( .A1(n8459), .A2(n8455), .ZN(n6757) );
  OR2_X1 U7788 ( .A1(n6757), .A2(n8452), .ZN(n6248) );
  AND3_X1 U7789 ( .A1(n6248), .A2(n8374), .A3(n10118), .ZN(n6277) );
  NAND2_X1 U7790 ( .A1(n6752), .A2(n6277), .ZN(n6250) );
  INV_X1 U7791 ( .A(n6223), .ZN(n6247) );
  INV_X1 U7792 ( .A(n7037), .ZN(n7400) );
  INV_X1 U7793 ( .A(n7041), .ZN(n6246) );
  NAND3_X1 U7794 ( .A1(n6247), .A2(n7400), .A3(n6246), .ZN(n6284) );
  NOR2_X1 U7795 ( .A1(n6248), .A2(n8453), .ZN(n6750) );
  NAND2_X1 U7796 ( .A1(n6754), .A2(n6750), .ZN(n6249) );
  INV_X1 U7797 ( .A(n6251), .ZN(n6254) );
  INV_X1 U7798 ( .A(n6252), .ZN(n6253) );
  NAND3_X1 U7799 ( .A1(n6256), .A2(n8589), .A3(n6315), .ZN(n6292) );
  INV_X1 U7800 ( .A(n8944), .ZN(n8205) );
  NAND2_X1 U7801 ( .A1(n10141), .A2(n6257), .ZN(n8760) );
  NAND2_X1 U7802 ( .A1(n6752), .A2(n7046), .ZN(n6258) );
  NOR2_X1 U7803 ( .A1(n10118), .A2(n6257), .ZN(n7401) );
  INV_X1 U7804 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n6259) );
  INV_X1 U7805 ( .A(n8716), .ZN(n6263) );
  NAND2_X1 U7806 ( .A1(n6261), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n6262) );
  NAND2_X1 U7807 ( .A1(n6263), .A2(n6262), .ZN(n8481) );
  NAND2_X1 U7808 ( .A1(n8481), .A2(n5986), .ZN(n6270) );
  INV_X1 U7809 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n6267) );
  NAND2_X1 U7810 ( .A1(n5998), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n6266) );
  NAND2_X1 U7811 ( .A1(n6264), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n6265) );
  OAI211_X1 U7812 ( .C1(n6013), .C2(n6267), .A(n6266), .B(n6265), .ZN(n6268)
         );
  INV_X1 U7813 ( .A(n6268), .ZN(n6269) );
  INV_X1 U7814 ( .A(n6754), .ZN(n6271) );
  NAND2_X1 U7815 ( .A1(n8711), .A2(n8452), .ZN(n6758) );
  OR2_X1 U7816 ( .A1(n8374), .A2(n6758), .ZN(n8456) );
  NOR2_X1 U7817 ( .A1(n6271), .A2(n8456), .ZN(n6275) );
  INV_X1 U7818 ( .A(n8457), .ZN(n6577) );
  NAND2_X1 U7819 ( .A1(n8697), .A2(n6577), .ZN(n6273) );
  INV_X1 U7820 ( .A(n7062), .ZN(n6274) );
  INV_X1 U7821 ( .A(n6276), .ZN(n6279) );
  INV_X1 U7822 ( .A(n6277), .ZN(n6278) );
  NAND2_X1 U7823 ( .A1(n6278), .A2(n8760), .ZN(n6753) );
  NAND2_X1 U7824 ( .A1(n6279), .A2(n6753), .ZN(n6282) );
  NAND2_X1 U7825 ( .A1(n8388), .A2(n6758), .ZN(n7038) );
  NAND3_X1 U7826 ( .A1(n6580), .A2(n6579), .A3(n7038), .ZN(n6280) );
  AOI21_X1 U7827 ( .B1(n6284), .B2(n6750), .A(n6280), .ZN(n6281) );
  NAND2_X1 U7828 ( .A1(n6282), .A2(n6281), .ZN(n6283) );
  NAND2_X1 U7829 ( .A1(n6283), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6286) );
  NAND3_X1 U7830 ( .A1(n6284), .A2(n7049), .A3(n7039), .ZN(n6285) );
  NAND2_X2 U7831 ( .A1(n6286), .A2(n6285), .ZN(n8598) );
  AOI22_X1 U7832 ( .A1(n8735), .A2(n8598), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3151), .ZN(n6287) );
  OAI21_X1 U7833 ( .B1(n8576), .B2(n8595), .A(n6287), .ZN(n6288) );
  AOI21_X1 U7834 ( .B1(n8732), .B2(n8593), .A(n6288), .ZN(n6289) );
  NAND2_X1 U7835 ( .A1(n6292), .A2(n6291), .ZN(P2_U3154) );
  NAND2_X1 U7836 ( .A1(n6293), .A2(n8404), .ZN(n6296) );
  OR2_X1 U7837 ( .A1(n8402), .A2(n6294), .ZN(n6295) );
  XNOR2_X1 U7838 ( .A(n8382), .B(n6297), .ZN(n6298) );
  XNOR2_X1 U7839 ( .A(n8941), .B(n6298), .ZN(n6309) );
  INV_X1 U7840 ( .A(n6309), .ZN(n6299) );
  NAND2_X1 U7841 ( .A1(n6299), .A2(n8589), .ZN(n6314) );
  INV_X1 U7842 ( .A(n6308), .ZN(n6300) );
  NAND2_X1 U7843 ( .A1(n6300), .A2(n8742), .ZN(n6301) );
  NAND2_X1 U7844 ( .A1(n8716), .A2(n5986), .ZN(n8416) );
  INV_X1 U7845 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n8239) );
  NAND2_X1 U7846 ( .A1(n8409), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n6303) );
  NAND2_X1 U7847 ( .A1(n8228), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n6302) );
  OAI211_X1 U7848 ( .C1(n8412), .C2(n8239), .A(n6303), .B(n6302), .ZN(n6304)
         );
  INV_X1 U7849 ( .A(n6304), .ZN(n6305) );
  INV_X1 U7850 ( .A(n8474), .ZN(n8605) );
  NAND2_X1 U7851 ( .A1(n8605), .A2(n8593), .ZN(n6307) );
  AOI22_X1 U7852 ( .A1(n8481), .A2(n8598), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3151), .ZN(n6306) );
  OAI211_X1 U7853 ( .C1(n8583), .C2(n8595), .A(n6307), .B(n6306), .ZN(n6311)
         );
  NOR4_X1 U7854 ( .A1(n6309), .A2(n8583), .A3(n6308), .A4(n8573), .ZN(n6310)
         );
  AOI211_X1 U7855 ( .C1(n8887), .C2(n8585), .A(n6311), .B(n6310), .ZN(n6312)
         );
  OAI211_X1 U7856 ( .C1(n6315), .C2(n6314), .A(n6313), .B(n6312), .ZN(P2_U3160) );
  XNOR2_X1 U7857 ( .A(n6318), .B(n7575), .ZN(n7576) );
  XNOR2_X1 U7858 ( .A(n7576), .B(n10075), .ZN(n6319) );
  NOR2_X1 U7859 ( .A1(n6319), .A2(n8573), .ZN(n6326) );
  INV_X1 U7860 ( .A(n7658), .ZN(n7459) );
  NOR2_X1 U7861 ( .A1(n8602), .A2(n7459), .ZN(n6325) );
  AND2_X1 U7862 ( .A1(n8598), .A2(n7428), .ZN(n6324) );
  NAND2_X1 U7863 ( .A1(n8593), .A2(n8615), .ZN(n6322) );
  NOR2_X1 U7864 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6320), .ZN(n7008) );
  INV_X1 U7865 ( .A(n7008), .ZN(n6321) );
  OAI211_X1 U7866 ( .C1(n7396), .C2(n8595), .A(n6322), .B(n6321), .ZN(n6323)
         );
  OR4_X1 U7867 ( .A1(n6326), .A2(n6325), .A3(n6324), .A4(n6323), .ZN(P2_U3161)
         );
  NAND2_X1 U7868 ( .A1(n6580), .A2(n8374), .ZN(n6327) );
  NAND2_X1 U7869 ( .A1(n6327), .A2(n6579), .ZN(n6582) );
  NAND2_X1 U7870 ( .A1(n6582), .A2(n8226), .ZN(n6328) );
  NAND2_X1 U7871 ( .A1(n6328), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3150) );
  INV_X1 U7872 ( .A(n6379), .ZN(n6329) );
  NAND2_X1 U7873 ( .A1(n7305), .A2(n7219), .ZN(n7304) );
  NOR2_X2 U7874 ( .A1(n7227), .A2(n7339), .ZN(n7439) );
  INV_X1 U7875 ( .A(n8000), .ZN(n9090) );
  INV_X1 U7876 ( .A(n7984), .ZN(n9940) );
  OR2_X2 U7877 ( .A1(n9891), .A2(n9890), .ZN(n9892) );
  NOR2_X4 U7878 ( .A1(n9892), .A2(n9958), .ZN(n9624) );
  INV_X1 U7879 ( .A(n9749), .ZN(n9631) );
  NAND2_X1 U7880 ( .A1(n9779), .A2(n9572), .ZN(n9557) );
  NOR2_X2 U7881 ( .A1(n8096), .A2(n9481), .ZN(n9457) );
  NAND2_X1 U7882 ( .A1(n9458), .A2(n9457), .ZN(n9456) );
  NOR2_X2 U7883 ( .A1(n9456), .A2(n6331), .ZN(n6332) );
  INV_X1 U7884 ( .A(n6814), .ZN(n7702) );
  NAND2_X1 U7885 ( .A1(n4859), .A2(n9405), .ZN(n9376) );
  OAI211_X1 U7886 ( .C1(n4859), .C2(n9405), .A(n9573), .B(n9376), .ZN(n9384)
         );
  NAND2_X1 U7887 ( .A1(n6920), .A2(P1_B_REG_SCAN_IN), .ZN(n6334) );
  NAND2_X1 U7888 ( .A1(n6334), .A2(n9880), .ZN(n9392) );
  INV_X1 U7889 ( .A(n9392), .ZN(n6335) );
  NAND2_X1 U7890 ( .A1(n6388), .A2(n6335), .ZN(n9637) );
  NAND2_X1 U7891 ( .A1(n9384), .A2(n9637), .ZN(n6357) );
  NAND2_X1 U7892 ( .A1(n6336), .A2(P1_B_REG_SCAN_IN), .ZN(n6337) );
  MUX2_X1 U7893 ( .A(P1_B_REG_SCAN_IN), .B(n6337), .S(n7902), .Z(n6338) );
  NOR2_X1 U7894 ( .A1(P1_D_REG_19__SCAN_IN), .A2(P1_D_REG_2__SCAN_IN), .ZN(
        n6342) );
  NOR4_X1 U7895 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_3__SCAN_IN), .A4(P1_D_REG_4__SCAN_IN), .ZN(n6341) );
  NOR4_X1 U7896 ( .A1(P1_D_REG_9__SCAN_IN), .A2(P1_D_REG_10__SCAN_IN), .A3(
        P1_D_REG_11__SCAN_IN), .A4(P1_D_REG_12__SCAN_IN), .ZN(n6340) );
  NOR4_X1 U7897 ( .A1(P1_D_REG_5__SCAN_IN), .A2(P1_D_REG_6__SCAN_IN), .A3(
        P1_D_REG_7__SCAN_IN), .A4(P1_D_REG_8__SCAN_IN), .ZN(n6339) );
  NAND4_X1 U7898 ( .A1(n6342), .A2(n6341), .A3(n6340), .A4(n6339), .ZN(n6348)
         );
  NOR4_X1 U7899 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_18__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n6346) );
  NOR4_X1 U7900 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_13__SCAN_IN), .A3(
        P1_D_REG_14__SCAN_IN), .A4(P1_D_REG_16__SCAN_IN), .ZN(n6345) );
  NOR4_X1 U7901 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n6344) );
  NOR4_X1 U7902 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n6343) );
  NAND4_X1 U7903 ( .A1(n6346), .A2(n6345), .A3(n6344), .A4(n6343), .ZN(n6347)
         );
  NOR2_X1 U7904 ( .A1(n6348), .A2(n6347), .ZN(n6799) );
  NAND2_X1 U7905 ( .A1(n6831), .A2(n6799), .ZN(n6349) );
  INV_X1 U7906 ( .A(n6350), .ZN(n8069) );
  NAND2_X1 U7907 ( .A1(n8069), .A2(n6336), .ZN(n9791) );
  NAND2_X1 U7908 ( .A1(n7268), .A2(n9573), .ZN(n6829) );
  AND2_X1 U7909 ( .A1(n7257), .A2(n6829), .ZN(n6352) );
  NAND2_X1 U7910 ( .A1(n8069), .A2(n7902), .ZN(n9792) );
  MUX2_X1 U7911 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n6357), .S(n9968), .Z(n6355)
         );
  INV_X1 U7912 ( .A(n9788), .ZN(n9763) );
  AND2_X1 U7913 ( .A1(n9381), .A2(n9763), .ZN(n6354) );
  OR2_X1 U7914 ( .A1(n6355), .A2(n6354), .ZN(P1_U3520) );
  MUX2_X1 U7915 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n6357), .S(n9983), .Z(n6359)
         );
  INV_X1 U7916 ( .A(n9747), .ZN(n9678) );
  AND2_X1 U7917 ( .A1(n9381), .A2(n9678), .ZN(n6358) );
  OR2_X1 U7918 ( .A1(n6359), .A2(n6358), .ZN(P1_U3552) );
  NAND2_X1 U7919 ( .A1(n6364), .A2(P1_U3086), .ZN(n8071) );
  INV_X1 U7920 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6360) );
  INV_X1 U7921 ( .A(n6644), .ZN(n6935) );
  OAI222_X1 U7922 ( .A1(n8071), .A2(n6360), .B1(n6935), .B2(P1_U3086), .C1(
        n9797), .C2(n8078), .ZN(P1_U3353) );
  INV_X1 U7923 ( .A(n8071), .ZN(n9795) );
  AOI22_X1 U7924 ( .A1(n9295), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_3__SCAN_IN), .B2(n9795), .ZN(n6361) );
  OAI21_X1 U7925 ( .B1(n6365), .B2(n9797), .A(n6361), .ZN(P1_U3352) );
  OAI222_X1 U7926 ( .A1(n8071), .A2(n4600), .B1(n6641), .B2(P1_U3086), .C1(
        n9797), .C2(n4602), .ZN(P1_U3354) );
  AND2_X1 U7927 ( .A1(n6364), .A2(P2_U3151), .ZN(n7816) );
  INV_X2 U7928 ( .A(n7816), .ZN(n9022) );
  OAI222_X1 U7929 ( .A1(n9015), .A2(n4430), .B1(n9022), .B2(n6365), .C1(
        P2_U3151), .C2(n6626), .ZN(P2_U3292) );
  OAI222_X1 U7930 ( .A1(P2_U3151), .A2(n6676), .B1(n9022), .B2(n6367), .C1(
        n6366), .C2(n9015), .ZN(P2_U3291) );
  INV_X1 U7931 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6368) );
  INV_X1 U7932 ( .A(n6650), .ZN(n6948) );
  OAI222_X1 U7933 ( .A1(n8071), .A2(n6368), .B1(n6948), .B2(P1_U3086), .C1(
        n9797), .C2(n6367), .ZN(P1_U3351) );
  OAI222_X1 U7934 ( .A1(n6608), .A2(P2_U3151), .B1(n9015), .B2(n4959), .C1(
        n9022), .C2(n4602), .ZN(P2_U3294) );
  INV_X1 U7935 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6369) );
  OAI222_X1 U7936 ( .A1(n9797), .A2(n6370), .B1(n6652), .B2(P1_U3086), .C1(
        n6369), .C2(n8071), .ZN(P1_U3350) );
  OAI222_X1 U7937 ( .A1(P2_U3151), .A2(n6789), .B1(n9022), .B2(n6370), .C1(
        n4428), .C2(n9015), .ZN(P2_U3290) );
  AOI22_X1 U7938 ( .A1(n9323), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n9795), .ZN(n6371) );
  OAI21_X1 U7939 ( .B1(n6372), .B2(n9797), .A(n6371), .ZN(P1_U3349) );
  INV_X1 U7940 ( .A(n6796), .ZN(n6900) );
  OAI222_X1 U7941 ( .A1(P2_U3151), .A2(n6900), .B1(n9022), .B2(n6372), .C1(
        n4412), .C2(n9015), .ZN(P2_U3289) );
  AOI22_X1 U7942 ( .A1(n9336), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n9795), .ZN(n6373) );
  OAI21_X1 U7943 ( .B1(n6375), .B2(n9797), .A(n6373), .ZN(P1_U3348) );
  INV_X1 U7944 ( .A(n6995), .ZN(n7001) );
  INV_X1 U7945 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6374) );
  OAI222_X1 U7946 ( .A1(P2_U3151), .A2(n7001), .B1(n9022), .B2(n6375), .C1(
        n6374), .C2(n9015), .ZN(P2_U3288) );
  INV_X1 U7947 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n6428) );
  INV_X1 U7948 ( .A(n6376), .ZN(n6377) );
  AOI22_X1 U7949 ( .A1(n6380), .A2(n6428), .B1(n6379), .B2(n6377), .ZN(
        P2_U3377) );
  AOI22_X1 U7950 ( .A1(n6380), .A2(n5854), .B1(n6379), .B2(n6378), .ZN(
        P2_U3376) );
  AND2_X1 U7951 ( .A1(n6380), .A2(P2_D_REG_30__SCAN_IN), .ZN(P2_U3235) );
  AND2_X1 U7952 ( .A1(n6380), .A2(P2_D_REG_29__SCAN_IN), .ZN(P2_U3236) );
  AND2_X1 U7953 ( .A1(n6380), .A2(P2_D_REG_15__SCAN_IN), .ZN(P2_U3250) );
  AND2_X1 U7954 ( .A1(n6380), .A2(P2_D_REG_17__SCAN_IN), .ZN(P2_U3248) );
  AND2_X1 U7955 ( .A1(n6380), .A2(P2_D_REG_16__SCAN_IN), .ZN(P2_U3249) );
  AND2_X1 U7956 ( .A1(n6380), .A2(P2_D_REG_9__SCAN_IN), .ZN(P2_U3256) );
  AND2_X1 U7957 ( .A1(n6380), .A2(P2_D_REG_8__SCAN_IN), .ZN(P2_U3257) );
  AND2_X1 U7958 ( .A1(n6380), .A2(P2_D_REG_7__SCAN_IN), .ZN(P2_U3258) );
  AND2_X1 U7959 ( .A1(n6380), .A2(P2_D_REG_6__SCAN_IN), .ZN(P2_U3259) );
  AND2_X1 U7960 ( .A1(n6380), .A2(P2_D_REG_5__SCAN_IN), .ZN(P2_U3260) );
  AND2_X1 U7961 ( .A1(n6380), .A2(P2_D_REG_4__SCAN_IN), .ZN(P2_U3261) );
  AND2_X1 U7962 ( .A1(n6380), .A2(P2_D_REG_3__SCAN_IN), .ZN(P2_U3262) );
  AND2_X1 U7963 ( .A1(n6380), .A2(P2_D_REG_2__SCAN_IN), .ZN(P2_U3263) );
  AND2_X1 U7964 ( .A1(n6380), .A2(P2_D_REG_14__SCAN_IN), .ZN(P2_U3251) );
  AND2_X1 U7965 ( .A1(n6380), .A2(P2_D_REG_13__SCAN_IN), .ZN(P2_U3252) );
  AND2_X1 U7966 ( .A1(n6380), .A2(P2_D_REG_12__SCAN_IN), .ZN(P2_U3253) );
  AND2_X1 U7967 ( .A1(n6380), .A2(P2_D_REG_10__SCAN_IN), .ZN(P2_U3255) );
  AND2_X1 U7968 ( .A1(n6380), .A2(P2_D_REG_27__SCAN_IN), .ZN(P2_U3238) );
  AND2_X1 U7969 ( .A1(n6380), .A2(P2_D_REG_26__SCAN_IN), .ZN(P2_U3239) );
  AND2_X1 U7970 ( .A1(n6380), .A2(P2_D_REG_25__SCAN_IN), .ZN(P2_U3240) );
  AND2_X1 U7971 ( .A1(n6380), .A2(P2_D_REG_24__SCAN_IN), .ZN(P2_U3241) );
  AND2_X1 U7972 ( .A1(n6380), .A2(P2_D_REG_22__SCAN_IN), .ZN(P2_U3243) );
  AND2_X1 U7973 ( .A1(n6380), .A2(P2_D_REG_21__SCAN_IN), .ZN(P2_U3244) );
  AND2_X1 U7974 ( .A1(n6380), .A2(P2_D_REG_20__SCAN_IN), .ZN(P2_U3245) );
  AND2_X1 U7975 ( .A1(n6380), .A2(P2_D_REG_19__SCAN_IN), .ZN(P2_U3246) );
  AND2_X1 U7976 ( .A1(n6380), .A2(P2_D_REG_31__SCAN_IN), .ZN(P2_U3234) );
  INV_X1 U7977 ( .A(n6380), .ZN(n6382) );
  INV_X1 U7978 ( .A(P2_D_REG_23__SCAN_IN), .ZN(n6381) );
  NOR2_X1 U7979 ( .A1(n6382), .A2(n6381), .ZN(P2_U3242) );
  INV_X1 U7980 ( .A(P2_D_REG_28__SCAN_IN), .ZN(n6421) );
  NOR2_X1 U7981 ( .A1(n6382), .A2(n6421), .ZN(P2_U3237) );
  INV_X1 U7982 ( .A(P2_D_REG_18__SCAN_IN), .ZN(n6544) );
  NOR2_X1 U7983 ( .A1(n6382), .A2(n6544), .ZN(P2_U3247) );
  INV_X1 U7984 ( .A(P2_D_REG_11__SCAN_IN), .ZN(n6435) );
  NOR2_X1 U7985 ( .A1(n6382), .A2(n6435), .ZN(P2_U3254) );
  NAND2_X1 U7986 ( .A1(n6824), .A2(n7814), .ZN(n6392) );
  NAND2_X1 U7987 ( .A1(n6808), .A2(n7147), .ZN(n6383) );
  NAND2_X1 U7988 ( .A1(n5267), .A2(n6383), .ZN(n6390) );
  NAND2_X1 U7989 ( .A1(n6392), .A2(n6390), .ZN(n9872) );
  INV_X1 U7990 ( .A(n9872), .ZN(n9375) );
  NOR2_X1 U7991 ( .A1(n9375), .A2(P1_U3973), .ZN(P1_U3085) );
  INV_X1 U7992 ( .A(n6399), .ZN(n6384) );
  INV_X1 U7993 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6429) );
  OAI222_X1 U7994 ( .A1(n7104), .A2(P2_U3151), .B1(n9022), .B2(n6384), .C1(
        n6429), .C2(n9015), .ZN(P2_U3287) );
  NAND2_X1 U7995 ( .A1(n7063), .A2(P2_U3893), .ZN(n6385) );
  OAI21_X1 U7996 ( .B1(P2_U3893), .B2(n4964), .A(n6385), .ZN(P2_U3491) );
  NAND2_X1 U7997 ( .A1(n7455), .A2(P1_U3973), .ZN(n6386) );
  OAI21_X1 U7998 ( .B1(P1_U3973), .B2(n4516), .A(n6386), .ZN(P1_U3554) );
  INV_X2 U7999 ( .A(P1_U3973), .ZN(n9273) );
  NAND2_X1 U8000 ( .A1(n9273), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n6387) );
  OAI21_X1 U8001 ( .B1(n9393), .B2(n9273), .A(n6387), .ZN(P1_U3584) );
  NAND2_X1 U8002 ( .A1(n6388), .A2(P1_U3973), .ZN(n6389) );
  OAI21_X1 U8003 ( .B1(P1_U3973), .B2(n9011), .A(n6389), .ZN(P1_U3585) );
  INV_X1 U8004 ( .A(n6390), .ZN(n6391) );
  NAND2_X1 U8005 ( .A1(n6392), .A2(n6391), .ZN(n6658) );
  INV_X1 U8006 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n6394) );
  OR2_X1 U8007 ( .A1(n8084), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n6393) );
  NAND2_X1 U8008 ( .A1(n6393), .A2(n7148), .ZN(n6924) );
  AOI21_X1 U8009 ( .B1(n8084), .B2(n6394), .A(n6924), .ZN(n6395) );
  XNOR2_X1 U8010 ( .A(n6395), .B(n9799), .ZN(n6397) );
  AOI22_X1 U8011 ( .A1(n9375), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n6396) );
  OAI21_X1 U8012 ( .B1(n6658), .B2(n6397), .A(n6396), .ZN(P1_U3243) );
  AOI222_X1 U8013 ( .A1(n6399), .A2(n6398), .B1(P2_DATAO_REG_8__SCAN_IN), .B2(
        n9795), .C1(P1_STATE_REG_SCAN_IN), .C2(n6696), .ZN(n6574) );
  INV_X1 U8014 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6767) );
  INV_X1 U8015 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6974) );
  AOI22_X1 U8016 ( .A1(n6767), .A2(keyinput74), .B1(n6974), .B2(keyinput70), 
        .ZN(n6400) );
  OAI221_X1 U8017 ( .B1(n6767), .B2(keyinput74), .C1(n6974), .C2(keyinput70), 
        .A(n6400), .ZN(n6409) );
  XNOR2_X1 U8018 ( .A(P2_REG3_REG_17__SCAN_IN), .B(keyinput72), .ZN(n6404) );
  XNOR2_X1 U8019 ( .A(SI_3_), .B(keyinput117), .ZN(n6403) );
  XNOR2_X1 U8020 ( .A(P1_IR_REG_29__SCAN_IN), .B(keyinput104), .ZN(n6402) );
  XNOR2_X1 U8021 ( .A(P1_REG3_REG_2__SCAN_IN), .B(keyinput95), .ZN(n6401) );
  NAND4_X1 U8022 ( .A1(n6404), .A2(n6403), .A3(n6402), .A4(n6401), .ZN(n6408)
         );
  XNOR2_X1 U8023 ( .A(n6405), .B(keyinput98), .ZN(n6407) );
  INV_X1 U8024 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n7249) );
  XNOR2_X1 U8025 ( .A(keyinput64), .B(n7249), .ZN(n6406) );
  NOR4_X1 U8026 ( .A1(n6409), .A2(n6408), .A3(n6407), .A4(n6406), .ZN(n6449)
         );
  XOR2_X1 U8027 ( .A(P1_IR_REG_9__SCAN_IN), .B(keyinput73), .Z(n6415) );
  XOR2_X1 U8028 ( .A(P2_REG3_REG_1__SCAN_IN), .B(keyinput110), .Z(n6414) );
  INV_X1 U8029 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n7054) );
  XNOR2_X1 U8030 ( .A(keyinput82), .B(n7054), .ZN(n6413) );
  XNOR2_X1 U8031 ( .A(P2_REG1_REG_25__SCAN_IN), .B(keyinput125), .ZN(n6411) );
  XNOR2_X1 U8032 ( .A(P2_IR_REG_1__SCAN_IN), .B(keyinput96), .ZN(n6410) );
  NAND2_X1 U8033 ( .A1(n6411), .A2(n6410), .ZN(n6412) );
  OR4_X1 U8034 ( .A1(n6415), .A2(n6414), .A3(n6413), .A4(n6412), .ZN(n6419) );
  AOI22_X1 U8035 ( .A1(n5562), .A2(keyinput100), .B1(n8070), .B2(keyinput75), 
        .ZN(n6416) );
  OAI221_X1 U8036 ( .B1(n5562), .B2(keyinput100), .C1(n8070), .C2(keyinput75), 
        .A(n6416), .ZN(n6418) );
  XNOR2_X1 U8037 ( .A(n7554), .B(keyinput118), .ZN(n6417) );
  NOR3_X1 U8038 ( .A1(n6419), .A2(n6418), .A3(n6417), .ZN(n6448) );
  INV_X1 U8039 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n9973) );
  AOI22_X1 U8040 ( .A1(n9105), .A2(keyinput87), .B1(keyinput123), .B2(n9973), 
        .ZN(n6420) );
  OAI221_X1 U8041 ( .B1(n9105), .B2(keyinput87), .C1(n9973), .C2(keyinput123), 
        .A(n6420), .ZN(n6423) );
  XNOR2_X1 U8042 ( .A(n6421), .B(keyinput107), .ZN(n6422) );
  NOR2_X1 U8043 ( .A1(n6423), .A2(n6422), .ZN(n6434) );
  INV_X1 U8044 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n10111) );
  INV_X1 U8045 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n6425) );
  AOI22_X1 U8046 ( .A1(n10111), .A2(keyinput114), .B1(n6425), .B2(keyinput68), 
        .ZN(n6424) );
  OAI221_X1 U8047 ( .B1(n10111), .B2(keyinput114), .C1(n6425), .C2(keyinput68), 
        .A(n6424), .ZN(n6426) );
  INV_X1 U8048 ( .A(n6426), .ZN(n6433) );
  AOI22_X1 U8049 ( .A1(n6429), .A2(keyinput78), .B1(keyinput84), .B2(n6428), 
        .ZN(n6427) );
  OAI221_X1 U8050 ( .B1(n6429), .B2(keyinput78), .C1(n6428), .C2(keyinput84), 
        .A(n6427), .ZN(n6430) );
  INV_X1 U8051 ( .A(n6430), .ZN(n6432) );
  XNOR2_X1 U8052 ( .A(P2_REG2_REG_2__SCAN_IN), .B(keyinput76), .ZN(n6431) );
  AND4_X1 U8053 ( .A1(n6434), .A2(n6433), .A3(n6432), .A4(n6431), .ZN(n6447)
         );
  XOR2_X1 U8054 ( .A(keyinput66), .B(n6435), .Z(n6439) );
  XNOR2_X1 U8055 ( .A(P1_IR_REG_2__SCAN_IN), .B(keyinput79), .ZN(n6438) );
  XNOR2_X1 U8056 ( .A(P2_IR_REG_30__SCAN_IN), .B(keyinput94), .ZN(n6437) );
  XNOR2_X1 U8057 ( .A(P1_REG2_REG_0__SCAN_IN), .B(keyinput89), .ZN(n6436) );
  NAND4_X1 U8058 ( .A1(n6439), .A2(n6438), .A3(n6437), .A4(n6436), .ZN(n6445)
         );
  INV_X1 U8059 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n6843) );
  AOI22_X1 U8060 ( .A1(n5395), .A2(keyinput109), .B1(n6843), .B2(keyinput122), 
        .ZN(n6440) );
  OAI221_X1 U8061 ( .B1(n5395), .B2(keyinput109), .C1(n6843), .C2(keyinput122), 
        .A(n6440), .ZN(n6444) );
  INV_X1 U8062 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n6442) );
  INV_X1 U8063 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n8985) );
  AOI22_X1 U8064 ( .A1(n6442), .A2(keyinput80), .B1(keyinput71), .B2(n8985), 
        .ZN(n6441) );
  OAI221_X1 U8065 ( .B1(n6442), .B2(keyinput80), .C1(n8985), .C2(keyinput71), 
        .A(n6441), .ZN(n6443) );
  NOR3_X1 U8066 ( .A1(n6445), .A2(n6444), .A3(n6443), .ZN(n6446) );
  AND4_X1 U8067 ( .A1(n6449), .A2(n6448), .A3(n6447), .A4(n6446), .ZN(n6572)
         );
  OAI22_X1 U8068 ( .A1(P2_REG1_REG_28__SCAN_IN), .A2(keyinput86), .B1(
        P2_ADDR_REG_3__SCAN_IN), .B2(keyinput90), .ZN(n6450) );
  AOI221_X1 U8069 ( .B1(P2_REG1_REG_28__SCAN_IN), .B2(keyinput86), .C1(
        keyinput90), .C2(P2_ADDR_REG_3__SCAN_IN), .A(n6450), .ZN(n6457) );
  OAI22_X1 U8070 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(keyinput65), .B1(
        P2_IR_REG_10__SCAN_IN), .B2(keyinput101), .ZN(n6451) );
  AOI221_X1 U8071 ( .B1(P1_DATAO_REG_17__SCAN_IN), .B2(keyinput65), .C1(
        keyinput101), .C2(P2_IR_REG_10__SCAN_IN), .A(n6451), .ZN(n6456) );
  OAI22_X1 U8072 ( .A1(P1_D_REG_19__SCAN_IN), .A2(keyinput99), .B1(
        P1_REG2_REG_29__SCAN_IN), .B2(keyinput124), .ZN(n6452) );
  AOI221_X1 U8073 ( .B1(P1_D_REG_19__SCAN_IN), .B2(keyinput99), .C1(
        keyinput124), .C2(P1_REG2_REG_29__SCAN_IN), .A(n6452), .ZN(n6455) );
  OAI22_X1 U8074 ( .A1(P2_DATAO_REG_9__SCAN_IN), .A2(keyinput88), .B1(
        keyinput112), .B2(P1_REG1_REG_1__SCAN_IN), .ZN(n6453) );
  AOI221_X1 U8075 ( .B1(P2_DATAO_REG_9__SCAN_IN), .B2(keyinput88), .C1(
        P1_REG1_REG_1__SCAN_IN), .C2(keyinput112), .A(n6453), .ZN(n6454) );
  NAND4_X1 U8076 ( .A1(n6457), .A2(n6456), .A3(n6455), .A4(n6454), .ZN(n6485)
         );
  OAI22_X1 U8077 ( .A1(P1_D_REG_1__SCAN_IN), .A2(keyinput106), .B1(
        P1_REG0_REG_5__SCAN_IN), .B2(keyinput111), .ZN(n6458) );
  AOI221_X1 U8078 ( .B1(P1_D_REG_1__SCAN_IN), .B2(keyinput106), .C1(
        keyinput111), .C2(P1_REG0_REG_5__SCAN_IN), .A(n6458), .ZN(n6465) );
  OAI22_X1 U8079 ( .A1(P2_DATAO_REG_23__SCAN_IN), .A2(keyinput126), .B1(
        keyinput91), .B2(P2_REG0_REG_23__SCAN_IN), .ZN(n6459) );
  AOI221_X1 U8080 ( .B1(P2_DATAO_REG_23__SCAN_IN), .B2(keyinput126), .C1(
        P2_REG0_REG_23__SCAN_IN), .C2(keyinput91), .A(n6459), .ZN(n6464) );
  OAI22_X1 U8081 ( .A1(P2_D_REG_18__SCAN_IN), .A2(keyinput108), .B1(
        P2_REG3_REG_24__SCAN_IN), .B2(keyinput67), .ZN(n6460) );
  AOI221_X1 U8082 ( .B1(P2_D_REG_18__SCAN_IN), .B2(keyinput108), .C1(
        keyinput67), .C2(P2_REG3_REG_24__SCAN_IN), .A(n6460), .ZN(n6463) );
  OAI22_X1 U8083 ( .A1(P2_D_REG_23__SCAN_IN), .A2(keyinput92), .B1(
        P1_REG1_REG_30__SCAN_IN), .B2(keyinput120), .ZN(n6461) );
  AOI221_X1 U8084 ( .B1(P2_D_REG_23__SCAN_IN), .B2(keyinput92), .C1(
        keyinput120), .C2(P1_REG1_REG_30__SCAN_IN), .A(n6461), .ZN(n6462) );
  NAND4_X1 U8085 ( .A1(n6465), .A2(n6464), .A3(n6463), .A4(n6462), .ZN(n6484)
         );
  OAI22_X1 U8086 ( .A1(P1_REG3_REG_16__SCAN_IN), .A2(keyinput69), .B1(
        keyinput115), .B2(P1_REG3_REG_12__SCAN_IN), .ZN(n6466) );
  AOI221_X1 U8087 ( .B1(P1_REG3_REG_16__SCAN_IN), .B2(keyinput69), .C1(
        P1_REG3_REG_12__SCAN_IN), .C2(keyinput115), .A(n6466), .ZN(n6473) );
  OAI22_X1 U8088 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(keyinput102), .B1(
        P1_REG3_REG_5__SCAN_IN), .B2(keyinput81), .ZN(n6467) );
  AOI221_X1 U8089 ( .B1(P1_REG3_REG_6__SCAN_IN), .B2(keyinput102), .C1(
        keyinput81), .C2(P1_REG3_REG_5__SCAN_IN), .A(n6467), .ZN(n6472) );
  OAI22_X1 U8090 ( .A1(n6523), .A2(keyinput105), .B1(keyinput85), .B2(
        P2_DATAO_REG_3__SCAN_IN), .ZN(n6468) );
  AOI221_X1 U8091 ( .B1(n6523), .B2(keyinput105), .C1(P2_DATAO_REG_3__SCAN_IN), 
        .C2(keyinput85), .A(n6468), .ZN(n6471) );
  OAI22_X1 U8092 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(keyinput77), .B1(
        P1_ADDR_REG_10__SCAN_IN), .B2(keyinput93), .ZN(n6469) );
  AOI221_X1 U8093 ( .B1(P1_IR_REG_12__SCAN_IN), .B2(keyinput77), .C1(
        keyinput93), .C2(P1_ADDR_REG_10__SCAN_IN), .A(n6469), .ZN(n6470) );
  NAND4_X1 U8094 ( .A1(n6473), .A2(n6472), .A3(n6471), .A4(n6470), .ZN(n6483)
         );
  OAI22_X1 U8095 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(keyinput113), .B1(
        keyinput97), .B2(P2_REG0_REG_15__SCAN_IN), .ZN(n6474) );
  AOI221_X1 U8096 ( .B1(P1_DATAO_REG_21__SCAN_IN), .B2(keyinput113), .C1(
        P2_REG0_REG_15__SCAN_IN), .C2(keyinput97), .A(n6474), .ZN(n6481) );
  OAI22_X1 U8097 ( .A1(P1_REG2_REG_7__SCAN_IN), .A2(keyinput83), .B1(
        P1_ADDR_REG_9__SCAN_IN), .B2(keyinput121), .ZN(n6475) );
  AOI221_X1 U8098 ( .B1(P1_REG2_REG_7__SCAN_IN), .B2(keyinput83), .C1(
        keyinput121), .C2(P1_ADDR_REG_9__SCAN_IN), .A(n6475), .ZN(n6480) );
  OAI22_X1 U8099 ( .A1(P2_DATAO_REG_2__SCAN_IN), .A2(keyinput127), .B1(
        P1_ADDR_REG_11__SCAN_IN), .B2(keyinput103), .ZN(n6476) );
  AOI221_X1 U8100 ( .B1(P2_DATAO_REG_2__SCAN_IN), .B2(keyinput127), .C1(
        keyinput103), .C2(P1_ADDR_REG_11__SCAN_IN), .A(n6476), .ZN(n6479) );
  OAI22_X1 U8101 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(keyinput116), .B1(
        keyinput119), .B2(P2_ADDR_REG_5__SCAN_IN), .ZN(n6477) );
  AOI221_X1 U8102 ( .B1(P2_IR_REG_18__SCAN_IN), .B2(keyinput116), .C1(
        P2_ADDR_REG_5__SCAN_IN), .C2(keyinput119), .A(n6477), .ZN(n6478) );
  NAND4_X1 U8103 ( .A1(n6481), .A2(n6480), .A3(n6479), .A4(n6478), .ZN(n6482)
         );
  NOR4_X1 U8104 ( .A1(n6485), .A2(n6484), .A3(n6483), .A4(n6482), .ZN(n6571)
         );
  AOI22_X1 U8105 ( .A1(P1_REG3_REG_16__SCAN_IN), .A2(keyinput5), .B1(
        P1_IR_REG_9__SCAN_IN), .B2(keyinput9), .ZN(n6486) );
  OAI221_X1 U8106 ( .B1(P1_REG3_REG_16__SCAN_IN), .B2(keyinput5), .C1(
        P1_IR_REG_9__SCAN_IN), .C2(keyinput9), .A(n6486), .ZN(n6493) );
  AOI22_X1 U8107 ( .A1(P2_REG3_REG_24__SCAN_IN), .A2(keyinput3), .B1(
        P1_REG3_REG_12__SCAN_IN), .B2(keyinput51), .ZN(n6487) );
  OAI221_X1 U8108 ( .B1(P2_REG3_REG_24__SCAN_IN), .B2(keyinput3), .C1(
        P1_REG3_REG_12__SCAN_IN), .C2(keyinput51), .A(n6487), .ZN(n6492) );
  AOI22_X1 U8109 ( .A1(P1_REG1_REG_30__SCAN_IN), .A2(keyinput56), .B1(
        P1_REG1_REG_28__SCAN_IN), .B2(keyinput34), .ZN(n6488) );
  OAI221_X1 U8110 ( .B1(P1_REG1_REG_30__SCAN_IN), .B2(keyinput56), .C1(
        P1_REG1_REG_28__SCAN_IN), .C2(keyinput34), .A(n6488), .ZN(n6491) );
  AOI22_X1 U8111 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(keyinput16), .B1(
        P2_D_REG_11__SCAN_IN), .B2(keyinput2), .ZN(n6489) );
  OAI221_X1 U8112 ( .B1(P2_REG3_REG_14__SCAN_IN), .B2(keyinput16), .C1(
        P2_D_REG_11__SCAN_IN), .C2(keyinput2), .A(n6489), .ZN(n6490) );
  NOR4_X1 U8113 ( .A1(n6493), .A2(n6492), .A3(n6491), .A4(n6490), .ZN(n6521)
         );
  AOI22_X1 U8114 ( .A1(P2_REG2_REG_0__SCAN_IN), .A2(keyinput18), .B1(SI_3_), 
        .B2(keyinput53), .ZN(n6494) );
  OAI221_X1 U8115 ( .B1(P2_REG2_REG_0__SCAN_IN), .B2(keyinput18), .C1(SI_3_), 
        .C2(keyinput53), .A(n6494), .ZN(n6501) );
  AOI22_X1 U8116 ( .A1(P2_REG2_REG_3__SCAN_IN), .A2(keyinput0), .B1(
        P2_IR_REG_18__SCAN_IN), .B2(keyinput52), .ZN(n6495) );
  OAI221_X1 U8117 ( .B1(P2_REG2_REG_3__SCAN_IN), .B2(keyinput0), .C1(
        P2_IR_REG_18__SCAN_IN), .C2(keyinput52), .A(n6495), .ZN(n6500) );
  AOI22_X1 U8118 ( .A1(P1_DATAO_REG_14__SCAN_IN), .A2(keyinput6), .B1(
        P2_DATAO_REG_23__SCAN_IN), .B2(keyinput62), .ZN(n6496) );
  OAI221_X1 U8119 ( .B1(P1_DATAO_REG_14__SCAN_IN), .B2(keyinput6), .C1(
        P2_DATAO_REG_23__SCAN_IN), .C2(keyinput62), .A(n6496), .ZN(n6499) );
  AOI22_X1 U8120 ( .A1(P2_D_REG_23__SCAN_IN), .A2(keyinput28), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(keyinput31), .ZN(n6497) );
  OAI221_X1 U8121 ( .B1(P2_D_REG_23__SCAN_IN), .B2(keyinput28), .C1(
        P1_REG3_REG_2__SCAN_IN), .C2(keyinput31), .A(n6497), .ZN(n6498) );
  NOR4_X1 U8122 ( .A1(n6501), .A2(n6500), .A3(n6499), .A4(n6498), .ZN(n6520)
         );
  AOI22_X1 U8123 ( .A1(P1_REG2_REG_0__SCAN_IN), .A2(keyinput25), .B1(
        P1_REG3_REG_6__SCAN_IN), .B2(keyinput38), .ZN(n6502) );
  OAI221_X1 U8124 ( .B1(P1_REG2_REG_0__SCAN_IN), .B2(keyinput25), .C1(
        P1_REG3_REG_6__SCAN_IN), .C2(keyinput38), .A(n6502), .ZN(n6509) );
  AOI22_X1 U8125 ( .A1(P2_REG1_REG_28__SCAN_IN), .A2(keyinput22), .B1(
        P2_IR_REG_30__SCAN_IN), .B2(keyinput30), .ZN(n6503) );
  OAI221_X1 U8126 ( .B1(P2_REG1_REG_28__SCAN_IN), .B2(keyinput22), .C1(
        P2_IR_REG_30__SCAN_IN), .C2(keyinput30), .A(n6503), .ZN(n6508) );
  AOI22_X1 U8127 ( .A1(P2_REG2_REG_25__SCAN_IN), .A2(keyinput4), .B1(
        P1_IR_REG_12__SCAN_IN), .B2(keyinput13), .ZN(n6504) );
  OAI221_X1 U8128 ( .B1(P2_REG2_REG_25__SCAN_IN), .B2(keyinput4), .C1(
        P1_IR_REG_12__SCAN_IN), .C2(keyinput13), .A(n6504), .ZN(n6507) );
  AOI22_X1 U8129 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(keyinput54), .B1(
        P2_D_REG_1__SCAN_IN), .B2(keyinput20), .ZN(n6505) );
  OAI221_X1 U8130 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(keyinput54), .C1(
        P2_D_REG_1__SCAN_IN), .C2(keyinput20), .A(n6505), .ZN(n6506) );
  NOR4_X1 U8131 ( .A1(n6509), .A2(n6508), .A3(n6507), .A4(n6506), .ZN(n6519)
         );
  AOI22_X1 U8132 ( .A1(P2_REG2_REG_2__SCAN_IN), .A2(keyinput12), .B1(
        P1_D_REG_1__SCAN_IN), .B2(keyinput42), .ZN(n6510) );
  OAI221_X1 U8133 ( .B1(P2_REG2_REG_2__SCAN_IN), .B2(keyinput12), .C1(
        P1_D_REG_1__SCAN_IN), .C2(keyinput42), .A(n6510), .ZN(n6517) );
  AOI22_X1 U8134 ( .A1(P2_REG0_REG_23__SCAN_IN), .A2(keyinput27), .B1(
        P1_REG2_REG_7__SCAN_IN), .B2(keyinput19), .ZN(n6511) );
  OAI221_X1 U8135 ( .B1(P2_REG0_REG_23__SCAN_IN), .B2(keyinput27), .C1(
        P1_REG2_REG_7__SCAN_IN), .C2(keyinput19), .A(n6511), .ZN(n6516) );
  AOI22_X1 U8136 ( .A1(P2_REG3_REG_1__SCAN_IN), .A2(keyinput46), .B1(
        P1_REG0_REG_10__SCAN_IN), .B2(keyinput45), .ZN(n6512) );
  OAI221_X1 U8137 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(keyinput46), .C1(
        P1_REG0_REG_10__SCAN_IN), .C2(keyinput45), .A(n6512), .ZN(n6515) );
  AOI22_X1 U8138 ( .A1(P2_REG0_REG_4__SCAN_IN), .A2(keyinput50), .B1(
        P1_DATAO_REG_8__SCAN_IN), .B2(keyinput14), .ZN(n6513) );
  OAI221_X1 U8139 ( .B1(P2_REG0_REG_4__SCAN_IN), .B2(keyinput50), .C1(
        P1_DATAO_REG_8__SCAN_IN), .C2(keyinput14), .A(n6513), .ZN(n6514) );
  NOR4_X1 U8140 ( .A1(n6517), .A2(n6516), .A3(n6515), .A4(n6514), .ZN(n6518)
         );
  NAND4_X1 U8141 ( .A1(n6521), .A2(n6520), .A3(n6519), .A4(n6518), .ZN(n6570)
         );
  AOI22_X1 U8142 ( .A1(n6523), .A2(keyinput41), .B1(keyinput24), .B2(n6601), 
        .ZN(n6522) );
  OAI221_X1 U8143 ( .B1(n6523), .B2(keyinput41), .C1(n6601), .C2(keyinput24), 
        .A(n6522), .ZN(n6526) );
  INV_X1 U8144 ( .A(P1_D_REG_19__SCAN_IN), .ZN(n9911) );
  XNOR2_X1 U8145 ( .A(n9911), .B(keyinput35), .ZN(n6525) );
  XOR2_X1 U8146 ( .A(P2_IR_REG_1__SCAN_IN), .B(keyinput32), .Z(n6524) );
  OR3_X1 U8147 ( .A1(n6526), .A2(n6525), .A3(n6524), .ZN(n6532) );
  INV_X1 U8148 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n9812) );
  AOI22_X1 U8149 ( .A1(n9812), .A2(keyinput29), .B1(n9406), .B2(keyinput60), 
        .ZN(n6527) );
  OAI221_X1 U8150 ( .B1(n9812), .B2(keyinput29), .C1(n9406), .C2(keyinput60), 
        .A(n6527), .ZN(n6531) );
  AOI22_X1 U8151 ( .A1(n6529), .A2(keyinput8), .B1(n5316), .B2(keyinput17), 
        .ZN(n6528) );
  OAI221_X1 U8152 ( .B1(n6529), .B2(keyinput8), .C1(n5316), .C2(keyinput17), 
        .A(n6528), .ZN(n6530) );
  NOR3_X1 U8153 ( .A1(n6532), .A2(n6531), .A3(n6530), .ZN(n6568) );
  AOI22_X1 U8154 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(keyinput1), .B1(n5319), 
        .B2(keyinput47), .ZN(n6533) );
  OAI221_X1 U8155 ( .B1(P1_DATAO_REG_17__SCAN_IN), .B2(keyinput1), .C1(n5319), 
        .C2(keyinput47), .A(n6533), .ZN(n6541) );
  AOI22_X1 U8156 ( .A1(n7703), .A2(keyinput49), .B1(keyinput23), .B2(n9105), 
        .ZN(n6534) );
  OAI221_X1 U8157 ( .B1(n7703), .B2(keyinput49), .C1(n9105), .C2(keyinput23), 
        .A(n6534), .ZN(n6540) );
  AOI22_X1 U8158 ( .A1(P2_REG0_REG_19__SCAN_IN), .A2(keyinput7), .B1(
        P2_D_REG_28__SCAN_IN), .B2(keyinput43), .ZN(n6535) );
  OAI221_X1 U8159 ( .B1(P2_REG0_REG_19__SCAN_IN), .B2(keyinput7), .C1(
        P2_D_REG_28__SCAN_IN), .C2(keyinput43), .A(n6535), .ZN(n6539) );
  XNOR2_X1 U8160 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(keyinput63), .ZN(n6537) );
  XNOR2_X1 U8161 ( .A(P1_REG1_REG_1__SCAN_IN), .B(keyinput48), .ZN(n6536) );
  NAND2_X1 U8162 ( .A1(n6537), .A2(n6536), .ZN(n6538) );
  NOR4_X1 U8163 ( .A1(n6541), .A2(n6540), .A3(n6539), .A4(n6538), .ZN(n6567)
         );
  AOI22_X1 U8164 ( .A1(n5562), .A2(keyinput36), .B1(keyinput55), .B2(n7538), 
        .ZN(n6542) );
  OAI221_X1 U8165 ( .B1(n5562), .B2(keyinput36), .C1(n7538), .C2(keyinput55), 
        .A(n6542), .ZN(n6551) );
  INV_X1 U8166 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n9824) );
  AOI22_X1 U8167 ( .A1(n6544), .A2(keyinput44), .B1(keyinput39), .B2(n9824), 
        .ZN(n6543) );
  OAI221_X1 U8168 ( .B1(n6544), .B2(keyinput44), .C1(n9824), .C2(keyinput39), 
        .A(n6543), .ZN(n6550) );
  INV_X1 U8169 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n7551) );
  AOI22_X1 U8170 ( .A1(n7551), .A2(keyinput57), .B1(n8070), .B2(keyinput11), 
        .ZN(n6545) );
  OAI221_X1 U8171 ( .B1(n7551), .B2(keyinput57), .C1(n8070), .C2(keyinput11), 
        .A(n6545), .ZN(n6549) );
  XNOR2_X1 U8172 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(keyinput21), .ZN(n6547) );
  XNOR2_X1 U8173 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(keyinput58), .ZN(n6546) );
  NAND2_X1 U8174 ( .A1(n6547), .A2(n6546), .ZN(n6548) );
  NOR4_X1 U8175 ( .A1(n6551), .A2(n6550), .A3(n6549), .A4(n6548), .ZN(n6566)
         );
  XOR2_X1 U8176 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(keyinput10), .Z(n6556) );
  XNOR2_X1 U8177 ( .A(n6552), .B(keyinput15), .ZN(n6555) );
  XNOR2_X1 U8178 ( .A(n6553), .B(keyinput40), .ZN(n6554) );
  NOR3_X1 U8179 ( .A1(n6556), .A2(n6555), .A3(n6554), .ZN(n6559) );
  XNOR2_X1 U8180 ( .A(P2_REG0_REG_15__SCAN_IN), .B(keyinput33), .ZN(n6558) );
  XNOR2_X1 U8181 ( .A(P2_IR_REG_10__SCAN_IN), .B(keyinput37), .ZN(n6557) );
  NAND3_X1 U8182 ( .A1(n6559), .A2(n6558), .A3(n6557), .ZN(n6564) );
  AOI22_X1 U8183 ( .A1(n6561), .A2(keyinput61), .B1(n9973), .B2(keyinput59), 
        .ZN(n6560) );
  OAI221_X1 U8184 ( .B1(n6561), .B2(keyinput61), .C1(n9973), .C2(keyinput59), 
        .A(n6560), .ZN(n6563) );
  INV_X1 U8185 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n7527) );
  XNOR2_X1 U8186 ( .A(n7527), .B(keyinput26), .ZN(n6562) );
  NOR3_X1 U8187 ( .A1(n6564), .A2(n6563), .A3(n6562), .ZN(n6565) );
  NAND4_X1 U8188 ( .A1(n6568), .A2(n6567), .A3(n6566), .A4(n6565), .ZN(n6569)
         );
  AOI211_X1 U8189 ( .C1(n6572), .C2(n6571), .A(n6570), .B(n6569), .ZN(n6573)
         );
  XNOR2_X1 U8190 ( .A(n6574), .B(n6573), .ZN(P1_U3347) );
  AOI22_X1 U8191 ( .A1(n9809), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n9795), .ZN(n6575) );
  OAI21_X1 U8192 ( .B1(n6603), .B2(n9797), .A(n6575), .ZN(P1_U3345) );
  NAND2_X1 U8193 ( .A1(P2_U3893), .A2(n8457), .ZN(n9989) );
  MUX2_X1 U8194 ( .A(P2_REG1_REG_1__SCAN_IN), .B(P2_REG2_REG_1__SCAN_IN), .S(
        n8697), .Z(n6609) );
  XNOR2_X1 U8195 ( .A(n6609), .B(n6597), .ZN(n6607) );
  INV_X1 U8196 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n6576) );
  MUX2_X1 U8197 ( .A(n6576), .B(n7054), .S(n8697), .Z(n6745) );
  NAND2_X1 U8198 ( .A1(n6745), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n6744) );
  XNOR2_X1 U8199 ( .A(n6607), .B(n6744), .ZN(n6599) );
  AND2_X1 U8200 ( .A1(n8697), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8073) );
  NAND2_X1 U8201 ( .A1(n6582), .A2(n8073), .ZN(n6578) );
  MUX2_X1 U8202 ( .A(n6578), .B(n8623), .S(n6577), .Z(n8712) );
  INV_X1 U8203 ( .A(n8712), .ZN(n10051) );
  INV_X1 U8204 ( .A(n6579), .ZN(n7818) );
  NOR2_X1 U8205 ( .A1(n6580), .A2(n7818), .ZN(n6581) );
  OR2_X1 U8206 ( .A1(P2_U3150), .A2(n6581), .ZN(n8654) );
  INV_X1 U8207 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n6589) );
  NOR2_X1 U8208 ( .A1(n8457), .A2(P2_U3151), .ZN(n9019) );
  AND2_X1 U8209 ( .A1(n6582), .A2(n9019), .ZN(n6747) );
  INV_X1 U8210 ( .A(n6747), .ZN(n6583) );
  INV_X1 U8211 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n6587) );
  AND2_X1 U8212 ( .A1(n4712), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6584) );
  NAND2_X1 U8213 ( .A1(n5937), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6623) );
  OAI21_X1 U8214 ( .B1(n6608), .B2(n6584), .A(n6623), .ZN(n6586) );
  OR2_X1 U8215 ( .A1(n6586), .A2(n6587), .ZN(n6624) );
  INV_X1 U8216 ( .A(n6624), .ZN(n6585) );
  AOI21_X1 U8217 ( .B1(n6587), .B2(n6586), .A(n6585), .ZN(n6588) );
  OAI22_X1 U8218 ( .A1(n8654), .A2(n6589), .B1(n10064), .B2(n6588), .ZN(n6596)
         );
  INV_X1 U8219 ( .A(n10058), .ZN(n8693) );
  NAND2_X1 U8220 ( .A1(n5937), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6621) );
  NAND2_X1 U8221 ( .A1(n6608), .A2(n6621), .ZN(n6593) );
  NAND2_X1 U8222 ( .A1(n4712), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6591) );
  OR2_X1 U8223 ( .A1(n6591), .A2(n5937), .ZN(n6592) );
  NAND2_X1 U8224 ( .A1(n6593), .A2(n6592), .ZN(n6620) );
  XOR2_X1 U8225 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n6620), .Z(n6594) );
  INV_X1 U8226 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n7059) );
  OAI22_X1 U8227 ( .A1(n8693), .A2(n6594), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7059), .ZN(n6595) );
  AOI211_X1 U8228 ( .C1(n6597), .C2(n10051), .A(n6596), .B(n6595), .ZN(n6598)
         );
  OAI21_X1 U8229 ( .B1(n9989), .B2(n6599), .A(n6598), .ZN(P2_U3183) );
  INV_X1 U8230 ( .A(n6600), .ZN(n6606) );
  INV_X1 U8231 ( .A(n7085), .ZN(n7094) );
  OAI222_X1 U8232 ( .A1(n9797), .A2(n6606), .B1(n7094), .B2(P1_U3086), .C1(
        n6601), .C2(n8071), .ZN(P1_U3346) );
  INV_X1 U8233 ( .A(n7280), .ZN(n7274) );
  INV_X1 U8234 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6602) );
  OAI222_X1 U8235 ( .A1(P2_U3151), .A2(n7274), .B1(n9022), .B2(n6603), .C1(
        n6602), .C2(n9015), .ZN(P2_U3285) );
  NAND2_X1 U8236 ( .A1(n9273), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n6604) );
  OAI21_X1 U8237 ( .B1(n9680), .B2(n9273), .A(n6604), .ZN(P1_U3576) );
  INV_X1 U8238 ( .A(n7177), .ZN(n7184) );
  OAI222_X1 U8239 ( .A1(P2_U3151), .A2(n7184), .B1(n9022), .B2(n6606), .C1(
        n6605), .C2(n9015), .ZN(P2_U3286) );
  MUX2_X1 U8240 ( .A(P2_REG1_REG_3__SCAN_IN), .B(P2_REG2_REG_3__SCAN_IN), .S(
        n8697), .Z(n6664) );
  XNOR2_X1 U8241 ( .A(n6664), .B(n6626), .ZN(n6618) );
  NAND2_X1 U8242 ( .A1(n6607), .A2(n6744), .ZN(n6611) );
  NAND2_X1 U8243 ( .A1(n6609), .A2(n6608), .ZN(n6610) );
  NAND2_X1 U8244 ( .A1(n6611), .A2(n6610), .ZN(n6704) );
  MUX2_X1 U8245 ( .A(P2_REG1_REG_2__SCAN_IN), .B(P2_REG2_REG_2__SCAN_IN), .S(
        n8697), .Z(n6613) );
  INV_X1 U8246 ( .A(n4316), .ZN(n6612) );
  XNOR2_X1 U8247 ( .A(n6613), .B(n6612), .ZN(n6705) );
  NAND2_X1 U8248 ( .A1(n6704), .A2(n6705), .ZN(n6615) );
  NAND2_X1 U8249 ( .A1(n6613), .A2(n4316), .ZN(n6614) );
  NAND2_X1 U8250 ( .A1(n6615), .A2(n6614), .ZN(n6617) );
  OR2_X1 U8251 ( .A1(n6617), .A2(n6618), .ZN(n6724) );
  INV_X1 U8252 ( .A(n6724), .ZN(n6616) );
  AOI21_X1 U8253 ( .B1(n6618), .B2(n6617), .A(n6616), .ZN(n6634) );
  INV_X1 U8254 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n6619) );
  NAND2_X1 U8255 ( .A1(n6620), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n6622) );
  NAND2_X1 U8256 ( .A1(n6622), .A2(n6621), .ZN(n6708) );
  AND2_X1 U8257 ( .A1(n6709), .A2(n6708), .ZN(n6706) );
  AOI21_X1 U8258 ( .B1(P2_REG1_REG_2__SCAN_IN), .B2(n4316), .A(n6706), .ZN(
        n6669) );
  INV_X1 U8259 ( .A(n6626), .ZN(n6670) );
  XNOR2_X1 U8260 ( .A(n6669), .B(n6670), .ZN(n6672) );
  XOR2_X1 U8261 ( .A(n6672), .B(P2_REG1_REG_3__SCAN_IN), .Z(n6631) );
  NOR2_X1 U8262 ( .A1(n5952), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7073) );
  NAND2_X1 U8263 ( .A1(n6624), .A2(n6623), .ZN(n6712) );
  INV_X1 U8264 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n7174) );
  NAND2_X1 U8265 ( .A1(n4316), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6625) );
  INV_X1 U8266 ( .A(n6730), .ZN(n6627) );
  AOI21_X1 U8267 ( .B1(n7249), .B2(n6628), .A(n6627), .ZN(n6629) );
  OAI22_X1 U8268 ( .A1(n8654), .A2(n7527), .B1(n10064), .B2(n6629), .ZN(n6630)
         );
  AOI211_X1 U8269 ( .C1(n10058), .C2(n6631), .A(n7073), .B(n6630), .ZN(n6633)
         );
  NAND2_X1 U8270 ( .A1(n10051), .A2(n6670), .ZN(n6632) );
  OAI211_X1 U8271 ( .C1(n6634), .C2(n9989), .A(n6633), .B(n6632), .ZN(P2_U3185) );
  INV_X1 U8272 ( .A(n9851), .ZN(n9868) );
  NAND2_X1 U8273 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n7936) );
  OAI21_X1 U8274 ( .B1(n9872), .B2(n7547), .A(n7936), .ZN(n6639) );
  INV_X1 U8275 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n6635) );
  INV_X1 U8276 ( .A(n9799), .ZN(n6925) );
  NOR3_X1 U8277 ( .A1(n9276), .A2(n6394), .A3(n6925), .ZN(n9275) );
  AOI21_X1 U8278 ( .B1(n9281), .B2(P1_REG1_REG_1__SCAN_IN), .A(n9275), .ZN(
        n6928) );
  XNOR2_X1 U8279 ( .A(n6644), .B(P1_REG1_REG_2__SCAN_IN), .ZN(n6927) );
  NOR2_X1 U8280 ( .A1(n6928), .A2(n6927), .ZN(n6926) );
  XNOR2_X1 U8281 ( .A(n9295), .B(P1_REG1_REG_3__SCAN_IN), .ZN(n9289) );
  XNOR2_X1 U8282 ( .A(n6650), .B(P1_REG1_REG_4__SCAN_IN), .ZN(n6945) );
  AOI21_X1 U8283 ( .B1(P1_REG1_REG_4__SCAN_IN), .B2(n6650), .A(n6944), .ZN(
        n9304) );
  XNOR2_X1 U8284 ( .A(n9309), .B(P1_REG1_REG_5__SCAN_IN), .ZN(n9303) );
  XNOR2_X1 U8285 ( .A(n9323), .B(P1_REG1_REG_6__SCAN_IN), .ZN(n9317) );
  XNOR2_X1 U8286 ( .A(n9336), .B(P1_REG1_REG_7__SCAN_IN), .ZN(n9331) );
  NOR2_X1 U8287 ( .A1(n4342), .A2(n9331), .ZN(n9330) );
  XNOR2_X1 U8288 ( .A(n6696), .B(P1_REG1_REG_8__SCAN_IN), .ZN(n6636) );
  AOI211_X1 U8289 ( .C1(n6637), .C2(n6636), .A(n9857), .B(n6695), .ZN(n6638)
         );
  AOI211_X1 U8290 ( .C1(n9868), .C2(n6696), .A(n6639), .B(n6638), .ZN(n6662)
         );
  INV_X1 U8291 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n6640) );
  XNOR2_X1 U8292 ( .A(n6696), .B(n6640), .ZN(n6660) );
  XNOR2_X1 U8293 ( .A(n6641), .B(P1_REG2_REG_1__SCAN_IN), .ZN(n9283) );
  NAND2_X1 U8294 ( .A1(n9799), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n6918) );
  INV_X1 U8295 ( .A(n6918), .ZN(n9284) );
  NAND2_X1 U8296 ( .A1(n9283), .A2(n9284), .ZN(n9282) );
  NAND2_X1 U8297 ( .A1(n9281), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6642) );
  NAND2_X1 U8298 ( .A1(n9282), .A2(n6642), .ZN(n6929) );
  INV_X1 U8299 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n6643) );
  XNOR2_X1 U8300 ( .A(n6644), .B(n6643), .ZN(n6930) );
  AND2_X1 U8301 ( .A1(n6929), .A2(n6930), .ZN(n6931) );
  INV_X1 U8302 ( .A(n6931), .ZN(n6646) );
  NAND2_X1 U8303 ( .A1(n6644), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6645) );
  NAND2_X1 U8304 ( .A1(n6646), .A2(n6645), .ZN(n9297) );
  INV_X1 U8305 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n6647) );
  XNOR2_X1 U8306 ( .A(n9295), .B(n6647), .ZN(n9298) );
  NAND2_X1 U8307 ( .A1(n9297), .A2(n9298), .ZN(n9296) );
  NAND2_X1 U8308 ( .A1(n9295), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6648) );
  NAND2_X1 U8309 ( .A1(n9296), .A2(n6648), .ZN(n6939) );
  INV_X1 U8310 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6649) );
  XNOR2_X1 U8311 ( .A(n6650), .B(n6649), .ZN(n6940) );
  AND2_X1 U8312 ( .A1(n6939), .A2(n6940), .ZN(n6941) );
  AND2_X1 U8313 ( .A1(n6650), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n6651) );
  OR2_X1 U8314 ( .A1(n6941), .A2(n6651), .ZN(n9311) );
  XNOR2_X1 U8315 ( .A(n6652), .B(P1_REG2_REG_5__SCAN_IN), .ZN(n9312) );
  NAND2_X1 U8316 ( .A1(n9311), .A2(n9312), .ZN(n9310) );
  NAND2_X1 U8317 ( .A1(n9309), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n6653) );
  NAND2_X1 U8318 ( .A1(n9310), .A2(n6653), .ZN(n9325) );
  INV_X1 U8319 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n6654) );
  XNOR2_X1 U8320 ( .A(n9323), .B(n6654), .ZN(n9326) );
  NAND2_X1 U8321 ( .A1(n9325), .A2(n9326), .ZN(n9324) );
  NAND2_X1 U8322 ( .A1(n9323), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6655) );
  NAND2_X1 U8323 ( .A1(n9324), .A2(n6655), .ZN(n9338) );
  INV_X1 U8324 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n6656) );
  XNOR2_X1 U8325 ( .A(n9336), .B(n6656), .ZN(n9339) );
  NAND2_X1 U8326 ( .A1(n9338), .A2(n9339), .ZN(n9337) );
  NAND2_X1 U8327 ( .A1(n9336), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n6657) );
  NAND2_X1 U8328 ( .A1(n9337), .A2(n6657), .ZN(n6659) );
  NAND2_X1 U8329 ( .A1(n6659), .A2(n6660), .ZN(n6691) );
  OAI211_X1 U8330 ( .C1(n6660), .C2(n6659), .A(n9842), .B(n6691), .ZN(n6661)
         );
  NAND2_X1 U8331 ( .A1(n6662), .A2(n6661), .ZN(P1_U3251) );
  INV_X1 U8332 ( .A(n5913), .ZN(n6765) );
  AOI22_X1 U8333 ( .A1(n9821), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n9795), .ZN(n6663) );
  OAI21_X1 U8334 ( .B1(n6765), .B2(n9797), .A(n6663), .ZN(P1_U3344) );
  MUX2_X1 U8335 ( .A(P2_REG1_REG_4__SCAN_IN), .B(P2_REG2_REG_4__SCAN_IN), .S(
        n8697), .Z(n6667) );
  INV_X1 U8336 ( .A(n6676), .ZN(n6740) );
  XNOR2_X1 U8337 ( .A(n6667), .B(n6740), .ZN(n6722) );
  INV_X1 U8338 ( .A(n6664), .ZN(n6665) );
  NAND2_X1 U8339 ( .A1(n6665), .A2(n6670), .ZN(n6723) );
  AND2_X1 U8340 ( .A1(n6722), .A2(n6723), .ZN(n6666) );
  NAND2_X1 U8341 ( .A1(n6724), .A2(n6666), .ZN(n6721) );
  NAND2_X1 U8342 ( .A1(n6667), .A2(n6676), .ZN(n6668) );
  NAND2_X1 U8343 ( .A1(n6721), .A2(n6668), .ZN(n6770) );
  MUX2_X1 U8344 ( .A(P2_REG1_REG_5__SCAN_IN), .B(P2_REG2_REG_5__SCAN_IN), .S(
        n8697), .Z(n6771) );
  INV_X1 U8345 ( .A(n6789), .ZN(n6673) );
  XNOR2_X1 U8346 ( .A(n6771), .B(n6673), .ZN(n6769) );
  XNOR2_X1 U8347 ( .A(n6770), .B(n6769), .ZN(n6689) );
  INV_X1 U8348 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n10149) );
  INV_X1 U8349 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n6671) );
  OAI22_X1 U8350 ( .A1(n6672), .A2(n6671), .B1(n6670), .B2(n6669), .ZN(n6733)
         );
  MUX2_X1 U8351 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n10149), .S(n6676), .Z(n6734)
         );
  NAND2_X1 U8352 ( .A1(n6733), .A2(n6734), .ZN(n6732) );
  OAI21_X1 U8353 ( .B1(n6740), .B2(n10149), .A(n6732), .ZN(n6788) );
  XNOR2_X1 U8354 ( .A(n6788), .B(n6673), .ZN(n6790) );
  XNOR2_X1 U8355 ( .A(n6790), .B(P2_REG1_REG_5__SCAN_IN), .ZN(n6687) );
  INV_X1 U8356 ( .A(n10064), .ZN(n10026) );
  NAND2_X1 U8357 ( .A1(n6730), .A2(n6725), .ZN(n6675) );
  INV_X1 U8358 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n6674) );
  MUX2_X1 U8359 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n6674), .S(n6676), .Z(n6726)
         );
  NAND2_X1 U8360 ( .A1(n6675), .A2(n6726), .ZN(n6728) );
  NAND2_X1 U8361 ( .A1(n6676), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n6677) );
  NAND2_X1 U8362 ( .A1(n6728), .A2(n6677), .ZN(n6678) );
  OAI21_X1 U8363 ( .B1(n6678), .B2(n6789), .A(n6781), .ZN(n6680) );
  INV_X1 U8364 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n6679) );
  NAND2_X1 U8365 ( .A1(n6680), .A2(n6679), .ZN(n6681) );
  NAND2_X1 U8366 ( .A1(n6783), .A2(n6681), .ZN(n6683) );
  NOR2_X1 U8367 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6682), .ZN(n6956) );
  AOI21_X1 U8368 ( .B1(n10026), .B2(n6683), .A(n6956), .ZN(n6685) );
  NAND2_X1 U8369 ( .A1(n10049), .A2(P2_ADDR_REG_5__SCAN_IN), .ZN(n6684) );
  OAI211_X1 U8370 ( .C1(n8712), .C2(n6789), .A(n6685), .B(n6684), .ZN(n6686)
         );
  AOI21_X1 U8371 ( .B1(n10058), .B2(n6687), .A(n6686), .ZN(n6688) );
  OAI21_X1 U8372 ( .B1(n6689), .B2(n9989), .A(n6688), .ZN(P2_U3187) );
  XNOR2_X1 U8373 ( .A(n7085), .B(P1_REG2_REG_9__SCAN_IN), .ZN(n6694) );
  NAND2_X1 U8374 ( .A1(n6696), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6690) );
  NAND2_X1 U8375 ( .A1(n6691), .A2(n6690), .ZN(n6693) );
  OR2_X1 U8376 ( .A1(n6693), .A2(n6694), .ZN(n7096) );
  INV_X1 U8377 ( .A(n7096), .ZN(n6692) );
  AOI21_X1 U8378 ( .B1(n6694), .B2(n6693), .A(n6692), .ZN(n6703) );
  MUX2_X1 U8379 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n9977), .S(n7085), .Z(n6697)
         );
  OAI21_X1 U8380 ( .B1(n6698), .B2(n6697), .A(n7084), .ZN(n6701) );
  INV_X1 U8381 ( .A(n9857), .ZN(n9847) );
  AND2_X1 U8382 ( .A1(P1_U3086), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n9175) );
  AOI21_X1 U8383 ( .B1(n9375), .B2(P1_ADDR_REG_9__SCAN_IN), .A(n9175), .ZN(
        n6699) );
  OAI21_X1 U8384 ( .B1(n7094), .B2(n9851), .A(n6699), .ZN(n6700) );
  AOI21_X1 U8385 ( .B1(n6701), .B2(n9847), .A(n6700), .ZN(n6702) );
  OAI21_X1 U8386 ( .B1(n6703), .B2(n9861), .A(n6702), .ZN(P1_U3252) );
  XOR2_X1 U8387 ( .A(n6705), .B(n6704), .Z(n6719) );
  INV_X1 U8388 ( .A(n6706), .ZN(n6707) );
  OAI21_X1 U8389 ( .B1(n6709), .B2(n6708), .A(n6707), .ZN(n6710) );
  AOI22_X1 U8390 ( .A1(n10049), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(n10058), .B2(
        n6710), .ZN(n6717) );
  OAI21_X1 U8391 ( .B1(n6713), .B2(n6712), .A(n6711), .ZN(n6715) );
  INV_X1 U8392 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n7171) );
  NOR2_X1 U8393 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7171), .ZN(n6714) );
  AOI21_X1 U8394 ( .B1(n10026), .B2(n6715), .A(n6714), .ZN(n6716) );
  OAI211_X1 U8395 ( .C1(n4316), .C2(n8712), .A(n6717), .B(n6716), .ZN(n6718)
         );
  AOI21_X1 U8396 ( .B1(n6719), .B2(n10057), .A(n6718), .ZN(n6720) );
  INV_X1 U8397 ( .A(n6720), .ZN(P2_U3184) );
  NAND2_X1 U8398 ( .A1(n6721), .A2(n10057), .ZN(n6743) );
  AOI21_X1 U8399 ( .B1(n6724), .B2(n6723), .A(n6722), .ZN(n6742) );
  INV_X1 U8400 ( .A(n6725), .ZN(n6727) );
  NOR2_X1 U8401 ( .A1(n6727), .A2(n6726), .ZN(n6731) );
  INV_X1 U8402 ( .A(n6728), .ZN(n6729) );
  AOI21_X1 U8403 ( .B1(n6731), .B2(n6730), .A(n6729), .ZN(n6738) );
  OAI21_X1 U8404 ( .B1(n6734), .B2(n6733), .A(n6732), .ZN(n6735) );
  AOI22_X1 U8405 ( .A1(n10049), .A2(P2_ADDR_REG_4__SCAN_IN), .B1(n10058), .B2(
        n6735), .ZN(n6737) );
  NAND2_X1 U8406 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3151), .ZN(n6736) );
  OAI211_X1 U8407 ( .C1(n6738), .C2(n10064), .A(n6737), .B(n6736), .ZN(n6739)
         );
  AOI21_X1 U8408 ( .B1(n6740), .B2(n10051), .A(n6739), .ZN(n6741) );
  OAI21_X1 U8409 ( .B1(n6743), .B2(n6742), .A(n6741), .ZN(P2_U3186) );
  AOI22_X1 U8410 ( .A1(n10049), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3151), .ZN(n6749) );
  OAI21_X1 U8411 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(n6745), .A(n6744), .ZN(n6746) );
  OAI21_X1 U8412 ( .B1(n10057), .B2(n6747), .A(n6746), .ZN(n6748) );
  OAI211_X1 U8413 ( .C1(n8712), .C2(n4712), .A(n6749), .B(n6748), .ZN(P2_U3182) );
  OR2_X1 U8414 ( .A1(n7049), .A2(n6750), .ZN(n6751) );
  NAND2_X1 U8415 ( .A1(n6752), .A2(n6751), .ZN(n6756) );
  NAND2_X1 U8416 ( .A1(n6754), .A2(n6753), .ZN(n6755) );
  NOR2_X1 U8417 ( .A1(n7162), .A2(n10074), .ZN(n7050) );
  INV_X1 U8418 ( .A(n7050), .ZN(n6762) );
  AND2_X1 U8419 ( .A1(n4501), .A2(n8453), .ZN(n8406) );
  NAND2_X1 U8420 ( .A1(n8711), .A2(n8459), .ZN(n6759) );
  NAND2_X1 U8421 ( .A1(n6759), .A2(n6758), .ZN(n6760) );
  NAND3_X1 U8422 ( .A1(n6760), .A2(n8456), .A3(n10118), .ZN(n8236) );
  INV_X1 U8423 ( .A(n8252), .ZN(n7057) );
  NAND2_X1 U8424 ( .A1(n7063), .A2(n7048), .ZN(n8255) );
  NAND2_X1 U8425 ( .A1(n7057), .A2(n8255), .ZN(n6839) );
  OAI21_X1 U8426 ( .B1(n8843), .B2(n10104), .A(n6839), .ZN(n6761) );
  OAI211_X1 U8427 ( .C1(n10118), .C2(n7048), .A(n6762), .B(n6761), .ZN(n8931)
         );
  NAND2_X1 U8428 ( .A1(n10142), .A2(n8931), .ZN(n6763) );
  OAI21_X1 U8429 ( .B1(n10142), .B2(n5927), .A(n6763), .ZN(P2_U3390) );
  INV_X1 U8430 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6764) );
  OAI222_X1 U8431 ( .A1(n7483), .A2(P2_U3151), .B1(n9022), .B2(n6765), .C1(
        n6764), .C2(n9015), .ZN(P2_U3284) );
  INV_X1 U8432 ( .A(n7910), .ZN(n7090) );
  INV_X1 U8433 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n6766) );
  OAI222_X1 U8434 ( .A1(n9797), .A2(n6768), .B1(n7090), .B2(P1_U3086), .C1(
        n6766), .C2(n8071), .ZN(P1_U3343) );
  OAI222_X1 U8435 ( .A1(P2_U3151), .A2(n8637), .B1(n9022), .B2(n6768), .C1(
        n6767), .C2(n9015), .ZN(P2_U3283) );
  NAND2_X1 U8436 ( .A1(n6770), .A2(n6769), .ZN(n6773) );
  NAND2_X1 U8437 ( .A1(n6771), .A2(n6789), .ZN(n6772) );
  NAND2_X1 U8438 ( .A1(n6773), .A2(n6772), .ZN(n6780) );
  INV_X1 U8439 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n6774) );
  INV_X1 U8440 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n7371) );
  MUX2_X1 U8441 ( .A(n6774), .B(n7371), .S(n8697), .Z(n6775) );
  NAND2_X1 U8442 ( .A1(n6775), .A2(n6796), .ZN(n6911) );
  INV_X1 U8443 ( .A(n6775), .ZN(n6776) );
  NAND2_X1 U8444 ( .A1(n6776), .A2(n6900), .ZN(n6777) );
  NAND2_X1 U8445 ( .A1(n6911), .A2(n6777), .ZN(n6779) );
  OR2_X1 U8446 ( .A1(n6780), .A2(n6779), .ZN(n6912) );
  INV_X1 U8447 ( .A(n6912), .ZN(n6778) );
  AOI21_X1 U8448 ( .B1(n6780), .B2(n6779), .A(n6778), .ZN(n6798) );
  INV_X1 U8449 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n7541) );
  XNOR2_X1 U8450 ( .A(n6796), .B(n7371), .ZN(n6782) );
  INV_X1 U8451 ( .A(n6899), .ZN(n6785) );
  NAND3_X1 U8452 ( .A1(n6783), .A2(n6782), .A3(n6781), .ZN(n6784) );
  NAND2_X1 U8453 ( .A1(n6785), .A2(n6784), .ZN(n6786) );
  NAND2_X1 U8454 ( .A1(n10026), .A2(n6786), .ZN(n6787) );
  NAND2_X1 U8455 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3151), .ZN(n7030) );
  OAI211_X1 U8456 ( .C1(n8654), .C2(n7541), .A(n6787), .B(n7030), .ZN(n6795)
         );
  MUX2_X1 U8457 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n6774), .S(n6796), .Z(n6792)
         );
  AOI22_X1 U8458 ( .A1(n6790), .A2(P2_REG1_REG_5__SCAN_IN), .B1(n6789), .B2(
        n6788), .ZN(n6791) );
  NOR2_X1 U8459 ( .A1(n6791), .A2(n6792), .ZN(n6898) );
  AOI21_X1 U8460 ( .B1(n6792), .B2(n6791), .A(n6898), .ZN(n6793) );
  NOR2_X1 U8461 ( .A1(n6793), .A2(n8693), .ZN(n6794) );
  AOI211_X1 U8462 ( .C1(n10051), .C2(n6796), .A(n6795), .B(n6794), .ZN(n6797)
         );
  OAI21_X1 U8463 ( .B1(n6798), .B2(n9989), .A(n6797), .ZN(P2_U3188) );
  NOR2_X1 U8464 ( .A1(n6800), .A2(n6799), .ZN(n6801) );
  NOR2_X1 U8465 ( .A1(n7257), .A2(n6801), .ZN(n6803) );
  INV_X1 U8466 ( .A(n6828), .ZN(n6834) );
  NAND2_X1 U8467 ( .A1(n9947), .A2(n6804), .ZN(n6823) );
  INV_X1 U8468 ( .A(n6823), .ZN(n6805) );
  NAND2_X1 U8469 ( .A1(n6834), .A2(n6805), .ZN(n6809) );
  INV_X1 U8470 ( .A(n6806), .ZN(n6807) );
  NAND4_X1 U8471 ( .A1(n6809), .A2(n6820), .A3(n6808), .A4(n6807), .ZN(n6810)
         );
  NAND2_X1 U8472 ( .A1(n6810), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6813) );
  NAND2_X1 U8473 ( .A1(n7262), .A2(n6888), .ZN(n7269) );
  INV_X1 U8474 ( .A(n6887), .ZN(n7263) );
  NAND2_X1 U8475 ( .A1(n7263), .A2(n6831), .ZN(n6833) );
  OAI21_X1 U8476 ( .B1(n7269), .B2(P1_U3086), .A(n6833), .ZN(n6811) );
  NAND2_X1 U8477 ( .A1(n6834), .A2(n6811), .ZN(n6812) );
  NOR2_X1 U8478 ( .A1(n9252), .A2(P1_U3086), .ZN(n6977) );
  INV_X1 U8479 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n6838) );
  NAND2_X1 U8480 ( .A1(n6814), .A2(n7526), .ZN(n6819) );
  OR2_X1 U8481 ( .A1(n6818), .A2(n6819), .ZN(n7303) );
  NAND2_X4 U8482 ( .A1(n6816), .A2(n4331), .ZN(n9113) );
  INV_X1 U8483 ( .A(n6819), .ZN(n6817) );
  NAND2_X2 U8484 ( .A1(n6820), .A2(n6817), .ZN(n6864) );
  INV_X1 U8485 ( .A(n6820), .ZN(n6822) );
  INV_X1 U8486 ( .A(n7455), .ZN(n7149) );
  NAND2_X1 U8487 ( .A1(n6818), .A2(n6884), .ZN(n6821) );
  OAI22_X1 U8488 ( .A1(n7149), .A2(n6864), .B1(n7129), .B2(n7150), .ZN(n6859)
         );
  XOR2_X1 U8489 ( .A(n6860), .B(n6861), .Z(n6921) );
  NOR2_X1 U8490 ( .A1(n6824), .A2(n6823), .ZN(n6825) );
  INV_X1 U8491 ( .A(n7269), .ZN(n6826) );
  AND2_X1 U8492 ( .A1(n6831), .A2(n6826), .ZN(n6827) );
  NAND2_X1 U8493 ( .A1(n6828), .A2(n6827), .ZN(n6832) );
  INV_X1 U8494 ( .A(n6829), .ZN(n6830) );
  NOR2_X1 U8495 ( .A1(n6834), .A2(n6833), .ZN(n6879) );
  NAND2_X1 U8496 ( .A1(n6879), .A2(n8467), .ZN(n9241) );
  INV_X1 U8497 ( .A(n6835), .ZN(n7299) );
  OAI22_X1 U8498 ( .A1(n9247), .A2(n7150), .B1(n9241), .B2(n7299), .ZN(n6836)
         );
  AOI21_X1 U8499 ( .B1(n6921), .B2(n9237), .A(n6836), .ZN(n6837) );
  OAI21_X1 U8500 ( .B1(n6977), .B2(n6838), .A(n6837), .ZN(P1_U3232) );
  NOR2_X1 U8501 ( .A1(n8598), .A2(P2_U3151), .ZN(n6968) );
  INV_X1 U8502 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n6842) );
  INV_X1 U8503 ( .A(n6839), .ZN(n8422) );
  OAI22_X1 U8504 ( .A1(n8573), .A2(n8422), .B1(n8602), .B2(n7048), .ZN(n6840)
         );
  AOI21_X1 U8505 ( .B1(n8593), .B2(n8624), .A(n6840), .ZN(n6841) );
  OAI21_X1 U8506 ( .B1(n6968), .B2(n6842), .A(n6841), .ZN(P2_U3172) );
  INV_X1 U8507 ( .A(n9833), .ZN(n6844) );
  OAI222_X1 U8508 ( .A1(n9797), .A2(n6846), .B1(n6844), .B2(P1_U3086), .C1(
        n6843), .C2(n8071), .ZN(P1_U3342) );
  INV_X1 U8509 ( .A(n9984), .ZN(n8662) );
  INV_X1 U8510 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6845) );
  OAI222_X1 U8511 ( .A1(P2_U3151), .A2(n8662), .B1(n9022), .B2(n6846), .C1(
        n6845), .C2(n9015), .ZN(P2_U3282) );
  NAND2_X1 U8512 ( .A1(n6847), .A2(n6848), .ZN(n6851) );
  INV_X1 U8513 ( .A(n6849), .ZN(n6850) );
  AOI21_X1 U8514 ( .B1(n6852), .B2(n6851), .A(n6850), .ZN(n6858) );
  OAI22_X1 U8515 ( .A1(n8582), .A2(n7359), .B1(n7315), .B2(n8595), .ZN(n6856)
         );
  INV_X1 U8516 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n6854) );
  OAI22_X1 U8517 ( .A1(n8602), .A2(n6853), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6854), .ZN(n6855) );
  AOI211_X1 U8518 ( .C1(n7381), .C2(n8598), .A(n6856), .B(n6855), .ZN(n6857)
         );
  OAI21_X1 U8519 ( .B1(n6858), .B2(n8573), .A(n6857), .ZN(P2_U3170) );
  INV_X1 U8520 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n6883) );
  OAI22_X1 U8521 ( .A1(n6861), .A2(n6860), .B1(n9030), .B2(n6859), .ZN(n6976)
         );
  NAND2_X1 U8522 ( .A1(n9274), .A2(n9049), .ZN(n6862) );
  OR2_X1 U8523 ( .A1(n8082), .A2(n6864), .ZN(n6866) );
  NAND2_X1 U8524 ( .A1(n9274), .A2(n9033), .ZN(n6865) );
  AND2_X1 U8525 ( .A1(n6866), .A2(n6865), .ZN(n6867) );
  NAND2_X1 U8526 ( .A1(n6868), .A2(n6867), .ZN(n6869) );
  OAI21_X1 U8527 ( .B1(n6868), .B2(n6867), .A(n6869), .ZN(n6975) );
  INV_X1 U8528 ( .A(n6869), .ZN(n6876) );
  OAI22_X1 U8529 ( .A1(n7129), .A2(n7219), .B1(n7220), .B2(n6864), .ZN(n6870)
         );
  XNOR2_X1 U8530 ( .A(n6870), .B(n9030), .ZN(n6872) );
  OAI22_X1 U8531 ( .A1(n7220), .A2(n9113), .B1(n7219), .B2(n6864), .ZN(n6871)
         );
  NAND2_X1 U8532 ( .A1(n6872), .A2(n6871), .ZN(n6873) );
  AND2_X1 U8533 ( .A1(n7015), .A2(n6873), .ZN(n6875) );
  OAI21_X1 U8534 ( .B1(n6874), .B2(n6876), .A(n6875), .ZN(n7016) );
  INV_X1 U8535 ( .A(n7016), .ZN(n6878) );
  NOR3_X1 U8536 ( .A1(n6874), .A2(n6876), .A3(n6875), .ZN(n6877) );
  OAI21_X1 U8537 ( .B1(n6878), .B2(n6877), .A(n9237), .ZN(n6882) );
  OAI22_X1 U8538 ( .A1(n7219), .A2(n9247), .B1(n9241), .B2(n7330), .ZN(n6880)
         );
  AOI21_X1 U8539 ( .B1(n9228), .B2(n9274), .A(n6880), .ZN(n6881) );
  OAI211_X1 U8540 ( .C1(n6977), .C2(n6883), .A(n6882), .B(n6881), .ZN(P1_U3237) );
  INV_X1 U8541 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n6895) );
  INV_X1 U8542 ( .A(n7262), .ZN(n6893) );
  OAI21_X1 U8543 ( .B1(n6884), .B2(n7526), .A(n6893), .ZN(n6885) );
  NOR2_X1 U8544 ( .A1(n7268), .A2(n6885), .ZN(n6886) );
  NOR2_X1 U8545 ( .A1(n9964), .A2(n9876), .ZN(n6892) );
  OAI222_X1 U8546 ( .A1(n7150), .A2(n6893), .B1(n7264), .B2(n6892), .C1(n9954), 
        .C2(n7299), .ZN(n6982) );
  NAND2_X1 U8547 ( .A1(n6982), .A2(n9968), .ZN(n6894) );
  OAI21_X1 U8548 ( .B1(n9968), .B2(n6895), .A(n6894), .ZN(P1_U3453) );
  INV_X1 U8549 ( .A(n6896), .ZN(n6973) );
  AOI22_X1 U8550 ( .A1(n9837), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n9795), .ZN(n6897) );
  OAI21_X1 U8551 ( .B1(n6973), .B2(n9797), .A(n6897), .ZN(P1_U3341) );
  AOI21_X1 U8552 ( .B1(P2_REG1_REG_6__SCAN_IN), .B2(n6900), .A(n6898), .ZN(
        n6994) );
  XNOR2_X1 U8553 ( .A(n6994), .B(n6995), .ZN(n6997) );
  INV_X1 U8554 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n6996) );
  XNOR2_X1 U8555 ( .A(n6997), .B(n6996), .ZN(n6916) );
  INV_X1 U8556 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n10090) );
  AOI21_X1 U8557 ( .B1(P2_REG2_REG_6__SCAN_IN), .B2(n6900), .A(n6899), .ZN(
        n7000) );
  XNOR2_X1 U8558 ( .A(n7000), .B(n6995), .ZN(n6901) );
  AOI21_X1 U8559 ( .B1(n10090), .B2(n6901), .A(n7004), .ZN(n6904) );
  AND2_X1 U8560 ( .A1(P2_U3151), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n7212) );
  INV_X1 U8561 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n7544) );
  NOR2_X1 U8562 ( .A1(n8654), .A2(n7544), .ZN(n6902) );
  AOI211_X1 U8563 ( .C1(n10051), .C2(n6995), .A(n7212), .B(n6902), .ZN(n6903)
         );
  OAI21_X1 U8564 ( .B1(n6904), .B2(n10064), .A(n6903), .ZN(n6915) );
  NAND2_X1 U8565 ( .A1(n6912), .A2(n6911), .ZN(n6908) );
  MUX2_X1 U8566 ( .A(n6996), .B(n10090), .S(n8697), .Z(n6905) );
  NAND2_X1 U8567 ( .A1(n6905), .A2(n6995), .ZN(n6989) );
  INV_X1 U8568 ( .A(n6905), .ZN(n6906) );
  NAND2_X1 U8569 ( .A1(n6906), .A2(n7001), .ZN(n6907) );
  AND2_X1 U8570 ( .A1(n6989), .A2(n6907), .ZN(n6909) );
  NAND2_X1 U8571 ( .A1(n6908), .A2(n6909), .ZN(n6992) );
  INV_X1 U8572 ( .A(n6909), .ZN(n6910) );
  NAND3_X1 U8573 ( .A1(n6912), .A2(n6911), .A3(n6910), .ZN(n6913) );
  AOI21_X1 U8574 ( .B1(n6992), .B2(n6913), .A(n9989), .ZN(n6914) );
  AOI211_X1 U8575 ( .C1(n10058), .C2(n6916), .A(n6915), .B(n6914), .ZN(n6917)
         );
  INV_X1 U8576 ( .A(n6917), .ZN(P2_U3189) );
  OAI21_X1 U8577 ( .B1(n6919), .B2(n6918), .A(P1_U3973), .ZN(n6923) );
  NOR3_X1 U8578 ( .A1(n6921), .A2(n6920), .A3(n8467), .ZN(n6922) );
  AOI211_X1 U8579 ( .C1(n6925), .C2(n6924), .A(n6923), .B(n6922), .ZN(n6952)
         );
  AOI211_X1 U8580 ( .C1(n6928), .C2(n6927), .A(n6926), .B(n9857), .ZN(n6938)
         );
  INV_X1 U8581 ( .A(n6929), .ZN(n6933) );
  INV_X1 U8582 ( .A(n6930), .ZN(n6932) );
  AOI211_X1 U8583 ( .C1(n6933), .C2(n6932), .A(n6931), .B(n9861), .ZN(n6937)
         );
  AOI22_X1 U8584 ( .A1(n9375), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n6934) );
  OAI21_X1 U8585 ( .B1(n6935), .B2(n9851), .A(n6934), .ZN(n6936) );
  OR4_X1 U8586 ( .A1(n6952), .A2(n6938), .A3(n6937), .A4(n6936), .ZN(P1_U3245)
         );
  INV_X1 U8587 ( .A(n6939), .ZN(n6943) );
  INV_X1 U8588 ( .A(n6940), .ZN(n6942) );
  AOI211_X1 U8589 ( .C1(n6943), .C2(n6942), .A(n6941), .B(n9861), .ZN(n6951)
         );
  AOI211_X1 U8590 ( .C1(n6946), .C2(n6945), .A(n6944), .B(n9857), .ZN(n6950)
         );
  AND2_X1 U8591 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n7137) );
  AOI21_X1 U8592 ( .B1(n9375), .B2(P1_ADDR_REG_4__SCAN_IN), .A(n7137), .ZN(
        n6947) );
  OAI21_X1 U8593 ( .B1(n6948), .B2(n9851), .A(n6947), .ZN(n6949) );
  OR4_X1 U8594 ( .A1(n6952), .A2(n6951), .A3(n6950), .A4(n6949), .ZN(P1_U3247)
         );
  XOR2_X1 U8595 ( .A(n6954), .B(n6953), .Z(n6959) );
  OAI22_X1 U8596 ( .A1(n8582), .A2(n10077), .B1(n7319), .B2(n8595), .ZN(n6955)
         );
  AOI211_X1 U8597 ( .C1(n7366), .C2(n8585), .A(n6956), .B(n6955), .ZN(n6958)
         );
  NAND2_X1 U8598 ( .A1(n8598), .A2(n7325), .ZN(n6957) );
  OAI211_X1 U8599 ( .C1(n6959), .C2(n8573), .A(n6958), .B(n6957), .ZN(P2_U3167) );
  XOR2_X1 U8600 ( .A(n6960), .B(n6961), .Z(n6965) );
  INV_X1 U8601 ( .A(n8595), .ZN(n8579) );
  OAI22_X1 U8602 ( .A1(n8602), .A2(n7055), .B1(n8582), .B2(n7242), .ZN(n6963)
         );
  NOR2_X1 U8603 ( .A1(n6968), .A2(n7059), .ZN(n6962) );
  AOI211_X1 U8604 ( .C1(n8579), .C2(n7063), .A(n6963), .B(n6962), .ZN(n6964)
         );
  OAI21_X1 U8605 ( .B1(n8573), .B2(n6965), .A(n6964), .ZN(P2_U3162) );
  XOR2_X1 U8606 ( .A(n6967), .B(n6966), .Z(n6972) );
  OAI22_X1 U8607 ( .A1(n10097), .A2(n8602), .B1(n8582), .B2(n7315), .ZN(n6970)
         );
  NOR2_X1 U8608 ( .A1(n6968), .A2(n7171), .ZN(n6969) );
  AOI211_X1 U8609 ( .C1(n8579), .C2(n8624), .A(n6970), .B(n6969), .ZN(n6971)
         );
  OAI21_X1 U8610 ( .B1(n8573), .B2(n6972), .A(n6971), .ZN(P2_U3177) );
  OAI222_X1 U8611 ( .A1(n9015), .A2(n6974), .B1(n9022), .B2(n6973), .C1(n8641), 
        .C2(P2_U3151), .ZN(P2_U3281) );
  AOI21_X1 U8612 ( .B1(n6976), .B2(n6975), .A(n6874), .ZN(n6981) );
  OAI22_X1 U8613 ( .A1(n8082), .A2(n9247), .B1(n9241), .B2(n7220), .ZN(n6979)
         );
  INV_X1 U8614 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n9279) );
  NOR2_X1 U8615 ( .A1(n6977), .A2(n9279), .ZN(n6978) );
  AOI211_X1 U8616 ( .C1(n9228), .C2(n7455), .A(n6979), .B(n6978), .ZN(n6980)
         );
  OAI21_X1 U8617 ( .B1(n6981), .B2(n9259), .A(n6980), .ZN(P1_U3222) );
  NAND2_X1 U8618 ( .A1(n6982), .A2(n9983), .ZN(n6983) );
  OAI21_X1 U8619 ( .B1(n9983), .B2(n6394), .A(n6983), .ZN(P1_U3522) );
  INV_X1 U8620 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n6984) );
  INV_X1 U8621 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7427) );
  MUX2_X1 U8622 ( .A(n6984), .B(n7427), .S(n8697), .Z(n6985) );
  NAND2_X1 U8623 ( .A1(n6985), .A2(n7118), .ZN(n7112) );
  INV_X1 U8624 ( .A(n6985), .ZN(n6986) );
  NAND2_X1 U8625 ( .A1(n6986), .A2(n7104), .ZN(n6987) );
  AND2_X1 U8626 ( .A1(n7112), .A2(n6987), .ZN(n6990) );
  INV_X1 U8627 ( .A(n6989), .ZN(n6988) );
  NOR2_X1 U8628 ( .A1(n6990), .A2(n6988), .ZN(n6993) );
  NAND2_X1 U8629 ( .A1(n6992), .A2(n6989), .ZN(n6991) );
  NAND2_X1 U8630 ( .A1(n6991), .A2(n6990), .ZN(n7113) );
  INV_X1 U8631 ( .A(n7113), .ZN(n7111) );
  AOI21_X1 U8632 ( .B1(n6993), .B2(n6992), .A(n7111), .ZN(n7014) );
  OAI22_X1 U8633 ( .A1(n6997), .A2(n6996), .B1(n6995), .B2(n6994), .ZN(n6999)
         );
  AOI22_X1 U8634 ( .A1(n7118), .A2(n6984), .B1(P2_REG1_REG_8__SCAN_IN), .B2(
        n7104), .ZN(n6998) );
  NAND2_X1 U8635 ( .A1(n6998), .A2(n6999), .ZN(n7117) );
  OAI21_X1 U8636 ( .B1(n6999), .B2(n6998), .A(n7117), .ZN(n7012) );
  INV_X1 U8637 ( .A(n7000), .ZN(n7002) );
  AOI22_X1 U8638 ( .A1(n7118), .A2(P2_REG2_REG_8__SCAN_IN), .B1(n7427), .B2(
        n7104), .ZN(n7005) );
  AOI21_X1 U8639 ( .B1(n7006), .B2(n7005), .A(n4397), .ZN(n7010) );
  NOR2_X1 U8640 ( .A1(n8712), .A2(n7104), .ZN(n7007) );
  AOI211_X1 U8641 ( .C1(n10049), .C2(P2_ADDR_REG_8__SCAN_IN), .A(n7008), .B(
        n7007), .ZN(n7009) );
  OAI21_X1 U8642 ( .B1(n7010), .B2(n10064), .A(n7009), .ZN(n7011) );
  AOI21_X1 U8643 ( .B1(n7012), .B2(n10058), .A(n7011), .ZN(n7013) );
  OAI21_X1 U8644 ( .B1(n7014), .B2(n9989), .A(n7013), .ZN(P2_U3190) );
  OR2_X1 U8645 ( .A1(n7330), .A2(n9113), .ZN(n7018) );
  NAND2_X1 U8646 ( .A1(n7228), .A2(n9049), .ZN(n7017) );
  NAND2_X1 U8647 ( .A1(n7018), .A2(n7017), .ZN(n7127) );
  AOI22_X1 U8648 ( .A1(n9272), .A2(n9049), .B1(n7228), .B2(n9044), .ZN(n7019)
         );
  AOI21_X1 U8649 ( .B1(n7021), .B2(n7020), .A(n7132), .ZN(n7026) );
  NAND2_X1 U8650 ( .A1(P1_U3086), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n9292) );
  INV_X1 U8651 ( .A(n9292), .ZN(n7023) );
  OAI22_X1 U8652 ( .A1(n7220), .A2(n9255), .B1(n9241), .B2(n7418), .ZN(n7022)
         );
  AOI211_X1 U8653 ( .C1(n7228), .C2(n9257), .A(n7023), .B(n7022), .ZN(n7025)
         );
  NAND2_X1 U8654 ( .A1(n9252), .A2(n7464), .ZN(n7024) );
  OAI211_X1 U8655 ( .C1(n7026), .C2(n9259), .A(n7025), .B(n7024), .ZN(P1_U3218) );
  INV_X1 U8656 ( .A(n7372), .ZN(n7035) );
  INV_X1 U8657 ( .A(n8598), .ZN(n8515) );
  OAI211_X1 U8658 ( .C1(n7029), .C2(n7028), .A(n7027), .B(n8589), .ZN(n7034)
         );
  INV_X1 U8659 ( .A(n7030), .ZN(n7032) );
  OAI22_X1 U8660 ( .A1(n8582), .A2(n7396), .B1(n7359), .B2(n8595), .ZN(n7031)
         );
  AOI211_X1 U8661 ( .C1(n7393), .C2(n8585), .A(n7032), .B(n7031), .ZN(n7033)
         );
  OAI211_X1 U8662 ( .C1(n7035), .C2(n8515), .A(n7034), .B(n7033), .ZN(P2_U3179) );
  NAND3_X1 U8663 ( .A1(n8711), .A2(n8459), .A3(n4501), .ZN(n7036) );
  NAND2_X1 U8664 ( .A1(n7036), .A2(n8374), .ZN(n7399) );
  INV_X1 U8665 ( .A(n7399), .ZN(n7403) );
  MUX2_X1 U8666 ( .A(n6223), .B(n7037), .S(n7403), .Z(n7044) );
  NAND2_X1 U8667 ( .A1(n7039), .A2(n7038), .ZN(n7040) );
  NOR2_X1 U8668 ( .A1(n7041), .A2(n7040), .ZN(n7042) );
  INV_X1 U8669 ( .A(n7045), .ZN(n7047) );
  INV_X1 U8670 ( .A(n7048), .ZN(n7060) );
  AOI22_X1 U8671 ( .A1(n10085), .A2(n7060), .B1(P2_REG3_REG_0__SCAN_IN), .B2(
        n10087), .ZN(n7053) );
  NOR3_X1 U8672 ( .A1(n8422), .A2(n7049), .A3(n10141), .ZN(n7051) );
  OAI21_X1 U8673 ( .B1(n7051), .B2(n7050), .A(n8867), .ZN(n7052) );
  OAI211_X1 U8674 ( .C1(n7054), .C2(n10091), .A(n7053), .B(n7052), .ZN(
        P2_U3233) );
  INV_X1 U8675 ( .A(n8453), .ZN(n7705) );
  NOR2_X1 U8676 ( .A1(n6257), .A2(n7705), .ZN(n7244) );
  NAND2_X1 U8677 ( .A1(n8867), .A2(n7244), .ZN(n8726) );
  INV_X1 U8678 ( .A(n8726), .ZN(n10086) );
  INV_X1 U8679 ( .A(n8253), .ZN(n8265) );
  NAND2_X1 U8680 ( .A1(n8624), .A2(n7055), .ZN(n8256) );
  NAND2_X1 U8681 ( .A1(n7057), .A2(n7056), .ZN(n7058) );
  NAND2_X1 U8682 ( .A1(n7160), .A2(n7058), .ZN(n10095) );
  OAI22_X1 U8683 ( .A1(n8779), .A2(n7055), .B1(n7059), .B2(n8813), .ZN(n7070)
         );
  INV_X1 U8684 ( .A(n8236), .ZN(n10084) );
  NAND2_X1 U8685 ( .A1(n10095), .A2(n10084), .ZN(n7068) );
  NAND2_X1 U8686 ( .A1(n7063), .A2(n7060), .ZN(n7061) );
  NAND2_X1 U8687 ( .A1(n7056), .A2(n7061), .ZN(n7166) );
  OAI21_X1 U8688 ( .B1(n7061), .B2(n7056), .A(n7166), .ZN(n7066) );
  NAND2_X1 U8689 ( .A1(n7063), .A2(n8838), .ZN(n7064) );
  OAI21_X1 U8690 ( .B1(n7242), .B2(n10074), .A(n7064), .ZN(n7065) );
  AOI21_X1 U8691 ( .B1(n7066), .B2(n8843), .A(n7065), .ZN(n7067) );
  NAND2_X1 U8692 ( .A1(n7068), .A2(n7067), .ZN(n10093) );
  MUX2_X1 U8693 ( .A(n10093), .B(P2_REG2_REG_1__SCAN_IN), .S(n10092), .Z(n7069) );
  AOI211_X1 U8694 ( .C1(n10086), .C2(n10095), .A(n7070), .B(n7069), .ZN(n7071)
         );
  INV_X1 U8695 ( .A(n7071), .ZN(P2_U3232) );
  INV_X1 U8696 ( .A(n7319), .ZN(n8620) );
  AOI22_X1 U8697 ( .A1(n8579), .A2(n8622), .B1(n8593), .B2(n8620), .ZN(n7075)
         );
  INV_X1 U8698 ( .A(n7073), .ZN(n7074) );
  OAI211_X1 U8699 ( .C1(n7072), .C2(n8602), .A(n7075), .B(n7074), .ZN(n7082)
         );
  NAND2_X1 U8700 ( .A1(n7077), .A2(n7076), .ZN(n7079) );
  INV_X1 U8701 ( .A(n6847), .ZN(n7078) );
  AOI211_X1 U8702 ( .C1(n7080), .C2(n7079), .A(n8573), .B(n7078), .ZN(n7081)
         );
  AOI211_X1 U8703 ( .C1(n5952), .C2(n8598), .A(n7082), .B(n7081), .ZN(n7083)
         );
  INV_X1 U8704 ( .A(n7083), .ZN(P2_U3158) );
  OAI21_X1 U8705 ( .B1(n7085), .B2(P1_REG1_REG_9__SCAN_IN), .A(n7084), .ZN(
        n9805) );
  INV_X1 U8706 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n7086) );
  MUX2_X1 U8707 ( .A(n7086), .B(P1_REG1_REG_10__SCAN_IN), .S(n9809), .Z(n9806)
         );
  NOR2_X1 U8708 ( .A1(n9805), .A2(n9806), .ZN(n9804) );
  MUX2_X1 U8709 ( .A(n4550), .B(P1_REG1_REG_11__SCAN_IN), .S(n9821), .Z(n9817)
         );
  INV_X1 U8710 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n9979) );
  AOI22_X1 U8711 ( .A1(P1_REG1_REG_12__SCAN_IN), .A2(n7910), .B1(n7090), .B2(
        n9979), .ZN(n7087) );
  OAI21_X1 U8712 ( .B1(n7088), .B2(n7087), .A(n7904), .ZN(n7092) );
  NAND2_X1 U8713 ( .A1(n9375), .A2(P1_ADDR_REG_12__SCAN_IN), .ZN(n7089) );
  NAND2_X1 U8714 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n8011) );
  OAI211_X1 U8715 ( .C1(n9851), .C2(n7090), .A(n7089), .B(n8011), .ZN(n7091)
         );
  AOI21_X1 U8716 ( .B1(n7092), .B2(n9847), .A(n7091), .ZN(n7103) );
  NOR2_X1 U8717 ( .A1(P1_REG2_REG_12__SCAN_IN), .A2(n7910), .ZN(n7093) );
  AOI21_X1 U8718 ( .B1(n7910), .B2(P1_REG2_REG_12__SCAN_IN), .A(n7093), .ZN(
        n7100) );
  NAND2_X1 U8719 ( .A1(n7094), .A2(n7622), .ZN(n7095) );
  NAND2_X1 U8720 ( .A1(n7096), .A2(n7095), .ZN(n9803) );
  NAND2_X1 U8721 ( .A1(n9809), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n7097) );
  OAI21_X1 U8722 ( .B1(n9809), .B2(P1_REG2_REG_10__SCAN_IN), .A(n7097), .ZN(
        n9802) );
  NOR2_X1 U8723 ( .A1(n9803), .A2(n9802), .ZN(n9801) );
  AOI21_X1 U8724 ( .B1(P1_REG2_REG_10__SCAN_IN), .B2(n9809), .A(n9801), .ZN(
        n9815) );
  NAND2_X1 U8725 ( .A1(n9821), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n7098) );
  OAI21_X1 U8726 ( .B1(n9821), .B2(P1_REG2_REG_11__SCAN_IN), .A(n7098), .ZN(
        n9814) );
  NOR2_X1 U8727 ( .A1(n9815), .A2(n9814), .ZN(n9813) );
  AOI21_X1 U8728 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n9821), .A(n9813), .ZN(
        n7099) );
  NAND2_X1 U8729 ( .A1(n7100), .A2(n7099), .ZN(n7909) );
  OAI21_X1 U8730 ( .B1(n7100), .B2(n7099), .A(n7909), .ZN(n7101) );
  NAND2_X1 U8731 ( .A1(n7101), .A2(n9842), .ZN(n7102) );
  NAND2_X1 U8732 ( .A1(n7103), .A2(n7102), .ZN(P1_U3255) );
  INV_X1 U8733 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7667) );
  AOI21_X1 U8734 ( .B1(n7667), .B2(n7105), .A(n7178), .ZN(n7125) );
  INV_X1 U8735 ( .A(n7112), .ZN(n7110) );
  INV_X1 U8736 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n7106) );
  MUX2_X1 U8737 ( .A(n7106), .B(n7667), .S(n8697), .Z(n7107) );
  NAND2_X1 U8738 ( .A1(n7107), .A2(n7177), .ZN(n7199) );
  INV_X1 U8739 ( .A(n7107), .ZN(n7108) );
  NAND2_X1 U8740 ( .A1(n7108), .A2(n7184), .ZN(n7109) );
  AND2_X1 U8741 ( .A1(n7199), .A2(n7109), .ZN(n7114) );
  NOR3_X1 U8742 ( .A1(n7111), .A2(n7110), .A3(n7114), .ZN(n7116) );
  NAND2_X1 U8743 ( .A1(n7113), .A2(n7112), .ZN(n7115) );
  NAND2_X1 U8744 ( .A1(n7115), .A2(n7114), .ZN(n7200) );
  INV_X1 U8745 ( .A(n7200), .ZN(n7198) );
  OAI21_X1 U8746 ( .B1(n7116), .B2(n7198), .A(n10057), .ZN(n7124) );
  OAI21_X1 U8747 ( .B1(n7118), .B2(n6984), .A(n7117), .ZN(n7183) );
  OAI21_X1 U8748 ( .B1(P2_REG1_REG_9__SCAN_IN), .B2(n7119), .A(n7185), .ZN(
        n7122) );
  INV_X1 U8749 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n7552) );
  NAND2_X1 U8750 ( .A1(n10051), .A2(n7177), .ZN(n7120) );
  NAND2_X1 U8751 ( .A1(P2_U3151), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n7580) );
  OAI211_X1 U8752 ( .C1(n7552), .C2(n8654), .A(n7120), .B(n7580), .ZN(n7121)
         );
  AOI21_X1 U8753 ( .B1(n7122), .B2(n10058), .A(n7121), .ZN(n7123) );
  OAI211_X1 U8754 ( .C1(n7125), .C2(n10064), .A(n7124), .B(n7123), .ZN(
        P2_U3191) );
  INV_X1 U8755 ( .A(n9252), .ZN(n9205) );
  INV_X1 U8756 ( .A(n7338), .ZN(n7140) );
  INV_X1 U8757 ( .A(n7126), .ZN(n7128) );
  OAI22_X1 U8758 ( .A1(n7418), .A2(n6864), .B1(n9921), .B2(n7129), .ZN(n7130)
         );
  XNOR2_X1 U8759 ( .A(n7130), .B(n9030), .ZN(n7412) );
  OAI22_X1 U8760 ( .A1(n7418), .A2(n9113), .B1(n9921), .B2(n6864), .ZN(n7411)
         );
  XNOR2_X1 U8761 ( .A(n7412), .B(n7411), .ZN(n7133) );
  OAI21_X1 U8762 ( .B1(n7132), .B2(n7134), .A(n7133), .ZN(n7135) );
  NAND3_X1 U8763 ( .A1(n4400), .A2(n9237), .A3(n7135), .ZN(n7139) );
  OAI22_X1 U8764 ( .A1(n7330), .A2(n9255), .B1(n9241), .B2(n7597), .ZN(n7136)
         );
  AOI211_X1 U8765 ( .C1(n7339), .C2(n9257), .A(n7137), .B(n7136), .ZN(n7138)
         );
  OAI211_X1 U8766 ( .C1(n9205), .C2(n7140), .A(n7139), .B(n7138), .ZN(P1_U3230) );
  INV_X1 U8767 ( .A(n10017), .ZN(n8631) );
  INV_X1 U8768 ( .A(n7141), .ZN(n7143) );
  INV_X1 U8769 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n7142) );
  OAI222_X1 U8770 ( .A1(n8631), .A2(P2_U3151), .B1(n9022), .B2(n7143), .C1(
        n7142), .C2(n9015), .ZN(P2_U3280) );
  OAI222_X1 U8771 ( .A1(n8071), .A2(n7144), .B1(n9797), .B2(n7143), .C1(
        P1_U3086), .C2(n9856), .ZN(P1_U3340) );
  NAND2_X1 U8772 ( .A1(n7145), .A2(n7146), .ZN(n7217) );
  OAI21_X1 U8773 ( .B1(n7145), .B2(n7146), .A(n7217), .ZN(n7449) );
  OAI22_X1 U8774 ( .A1(n7149), .A2(n9952), .B1(n7220), .B2(n9954), .ZN(n7152)
         );
  OAI21_X1 U8775 ( .B1(n8082), .B2(n7150), .A(n9573), .ZN(n7151) );
  NOR2_X1 U8776 ( .A1(n7151), .A2(n7305), .ZN(n7450) );
  AOI211_X1 U8777 ( .C1(n7449), .C2(n9964), .A(n7152), .B(n7450), .ZN(n7156)
         );
  INV_X1 U8778 ( .A(n7153), .ZN(n7154) );
  XNOR2_X1 U8779 ( .A(n7145), .B(n7154), .ZN(n7155) );
  NAND2_X1 U8780 ( .A1(n7155), .A2(n9876), .ZN(n7457) );
  NAND2_X1 U8781 ( .A1(n7156), .A2(n7457), .ZN(n8079) );
  INV_X1 U8782 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n7157) );
  OAI22_X1 U8783 ( .A1(n9788), .A2(n8082), .B1(n9968), .B2(n7157), .ZN(n7158)
         );
  AOI21_X1 U8784 ( .B1(n8079), .B2(n9968), .A(n7158), .ZN(n7159) );
  INV_X1 U8785 ( .A(n7159), .ZN(P1_U3456) );
  NAND2_X1 U8786 ( .A1(n7242), .A2(n10097), .ZN(n7250) );
  NAND2_X1 U8787 ( .A1(n8622), .A2(n7241), .ZN(n7161) );
  NAND2_X1 U8788 ( .A1(n7250), .A2(n7161), .ZN(n8421) );
  INV_X1 U8789 ( .A(n8421), .ZN(n7164) );
  XNOR2_X1 U8790 ( .A(n7240), .B(n7164), .ZN(n10098) );
  AOI22_X1 U8791 ( .A1(n8621), .A2(n8840), .B1(n8838), .B2(n8624), .ZN(n7170)
         );
  NAND2_X1 U8792 ( .A1(n7162), .A2(n7055), .ZN(n7165) );
  NAND2_X1 U8793 ( .A1(n7166), .A2(n7165), .ZN(n7163) );
  INV_X1 U8794 ( .A(n7251), .ZN(n7168) );
  AND3_X1 U8795 ( .A1(n7166), .A2(n8421), .A3(n7165), .ZN(n7167) );
  OAI21_X1 U8796 ( .B1(n7168), .B2(n7167), .A(n8843), .ZN(n7169) );
  OAI211_X1 U8797 ( .C1(n10098), .C2(n8236), .A(n7170), .B(n7169), .ZN(n10100)
         );
  OAI22_X1 U8798 ( .A1(n10097), .A2(n8760), .B1(n8813), .B2(n7171), .ZN(n7172)
         );
  NOR2_X1 U8799 ( .A1(n10100), .A2(n7172), .ZN(n7173) );
  MUX2_X1 U8800 ( .A(n7174), .B(n7173), .S(n10091), .Z(n7175) );
  OAI21_X1 U8801 ( .B1(n10098), .B2(n8726), .A(n7175), .ZN(P2_U3231) );
  NOR2_X1 U8802 ( .A1(n7177), .A2(n7176), .ZN(n7179) );
  NOR2_X1 U8803 ( .A1(n7179), .A2(n7178), .ZN(n7182) );
  INV_X1 U8804 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7682) );
  MUX2_X1 U8805 ( .A(P2_REG2_REG_10__SCAN_IN), .B(n7682), .S(n7280), .Z(n7181)
         );
  INV_X1 U8806 ( .A(n7276), .ZN(n7180) );
  AOI21_X1 U8807 ( .B1(n7182), .B2(n7181), .A(n7180), .ZN(n7207) );
  NAND2_X1 U8808 ( .A1(n7184), .A2(n7183), .ZN(n7186) );
  NAND2_X1 U8809 ( .A1(n7186), .A2(n7185), .ZN(n7188) );
  INV_X1 U8810 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n7193) );
  MUX2_X1 U8811 ( .A(n7193), .B(P2_REG1_REG_10__SCAN_IN), .S(n7280), .Z(n7187)
         );
  NAND2_X1 U8812 ( .A1(n7188), .A2(n7187), .ZN(n7279) );
  OAI21_X1 U8813 ( .B1(n7188), .B2(n7187), .A(n7279), .ZN(n7192) );
  NAND2_X1 U8814 ( .A1(n10051), .A2(n7280), .ZN(n7190) );
  INV_X1 U8815 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n7189) );
  OR2_X1 U8816 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7189), .ZN(n7608) );
  OAI211_X1 U8817 ( .C1(n7554), .C2(n8654), .A(n7190), .B(n7608), .ZN(n7191)
         );
  AOI21_X1 U8818 ( .B1(n7192), .B2(n10058), .A(n7191), .ZN(n7206) );
  INV_X1 U8819 ( .A(n7199), .ZN(n7197) );
  MUX2_X1 U8820 ( .A(n7193), .B(n7682), .S(n8697), .Z(n7194) );
  NAND2_X1 U8821 ( .A1(n7194), .A2(n7280), .ZN(n7285) );
  INV_X1 U8822 ( .A(n7194), .ZN(n7195) );
  NAND2_X1 U8823 ( .A1(n7195), .A2(n7274), .ZN(n7196) );
  AND2_X1 U8824 ( .A1(n7285), .A2(n7196), .ZN(n7201) );
  NOR3_X1 U8825 ( .A1(n7198), .A2(n7197), .A3(n7201), .ZN(n7204) );
  NAND2_X1 U8826 ( .A1(n7200), .A2(n7199), .ZN(n7202) );
  NAND2_X1 U8827 ( .A1(n7202), .A2(n7201), .ZN(n7286) );
  INV_X1 U8828 ( .A(n7286), .ZN(n7203) );
  OAI21_X1 U8829 ( .B1(n7204), .B2(n7203), .A(n10057), .ZN(n7205) );
  OAI211_X1 U8830 ( .C1(n7207), .C2(n10064), .A(n7206), .B(n7205), .ZN(
        P2_U3192) );
  AOI21_X1 U8831 ( .B1(n7210), .B2(n7209), .A(n4481), .ZN(n7215) );
  NOR2_X1 U8832 ( .A1(n8595), .A2(n10077), .ZN(n7211) );
  AOI211_X1 U8833 ( .C1(n8593), .C2(n8616), .A(n7212), .B(n7211), .ZN(n7214)
         );
  AOI22_X1 U8834 ( .A1(n8585), .A2(n10125), .B1(n10088), .B2(n8598), .ZN(n7213) );
  OAI211_X1 U8835 ( .C1(n7215), .C2(n8573), .A(n7214), .B(n7213), .ZN(P2_U3153) );
  INV_X1 U8836 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n7232) );
  NAND2_X1 U8837 ( .A1(n7299), .A2(n8082), .ZN(n7216) );
  NAND2_X1 U8838 ( .A1(n7217), .A2(n7216), .ZN(n7297) );
  NAND2_X1 U8839 ( .A1(n7297), .A2(n7218), .ZN(n7298) );
  NAND2_X1 U8840 ( .A1(n7220), .A2(n7219), .ZN(n7221) );
  NAND2_X1 U8841 ( .A1(n7298), .A2(n7221), .ZN(n7222) );
  OAI21_X1 U8842 ( .B1(n7222), .B2(n7223), .A(n7332), .ZN(n7469) );
  INV_X1 U8843 ( .A(n7469), .ZN(n7230) );
  XNOR2_X1 U8844 ( .A(n7224), .B(n7223), .ZN(n7226) );
  INV_X1 U8845 ( .A(n9952), .ZN(n9879) );
  AOI222_X1 U8846 ( .A1(n9876), .A2(n7226), .B1(n9271), .B2(n9880), .C1(n7225), 
        .C2(n9879), .ZN(n7471) );
  INV_X1 U8847 ( .A(n7227), .ZN(n7337) );
  AOI21_X1 U8848 ( .B1(n7228), .B2(n7304), .A(n7337), .ZN(n7463) );
  AOI22_X1 U8849 ( .A1(n7463), .A2(n9573), .B1(n9959), .B2(n7228), .ZN(n7229)
         );
  OAI211_X1 U8850 ( .C1(n9741), .C2(n7230), .A(n7471), .B(n7229), .ZN(n7233)
         );
  NAND2_X1 U8851 ( .A1(n7233), .A2(n9968), .ZN(n7231) );
  OAI21_X1 U8852 ( .B1(n9968), .B2(n7232), .A(n7231), .ZN(P1_U3462) );
  INV_X1 U8853 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n7235) );
  NAND2_X1 U8854 ( .A1(n7233), .A2(n9983), .ZN(n7234) );
  OAI21_X1 U8855 ( .B1(n9983), .B2(n7235), .A(n7234), .ZN(P1_U3525) );
  INV_X1 U8856 ( .A(n7236), .ZN(n7238) );
  INV_X1 U8857 ( .A(n10033), .ZN(n8646) );
  OAI222_X1 U8858 ( .A1(n9015), .A2(n7237), .B1(n9022), .B2(n7238), .C1(
        P2_U3151), .C2(n8646), .ZN(P2_U3279) );
  OAI222_X1 U8859 ( .A1(n8071), .A2(n7239), .B1(n7915), .B2(P1_U3086), .C1(
        n9797), .C2(n7238), .ZN(P1_U3339) );
  NAND2_X1 U8860 ( .A1(n7240), .A2(n8421), .ZN(n7243) );
  NAND2_X1 U8861 ( .A1(n7242), .A2(n7241), .ZN(n8260) );
  NAND2_X1 U8862 ( .A1(n7243), .A2(n8260), .ZN(n7312) );
  NAND2_X1 U8863 ( .A1(n7315), .A2(n7247), .ZN(n8277) );
  NAND2_X1 U8864 ( .A1(n8621), .A2(n7072), .ZN(n8270) );
  XNOR2_X1 U8865 ( .A(n7312), .B(n7311), .ZN(n10105) );
  INV_X1 U8866 ( .A(n7244), .ZN(n7245) );
  NAND2_X1 U8867 ( .A1(n8236), .A2(n7245), .ZN(n7246) );
  AOI22_X1 U8868 ( .A1(n10085), .A2(n7247), .B1(n5952), .B2(n10087), .ZN(n7248) );
  OAI21_X1 U8869 ( .B1(n7249), .B2(n10091), .A(n7248), .ZN(n7255) );
  NAND2_X1 U8870 ( .A1(n7251), .A2(n7250), .ZN(n7363) );
  INV_X1 U8871 ( .A(n7311), .ZN(n8420) );
  NAND2_X1 U8872 ( .A1(n7363), .A2(n8420), .ZN(n7378) );
  NAND3_X1 U8873 ( .A1(n7251), .A2(n7311), .A3(n7250), .ZN(n7252) );
  NAND2_X1 U8874 ( .A1(n7378), .A2(n7252), .ZN(n7253) );
  AOI222_X1 U8875 ( .A1(n8843), .A2(n7253), .B1(n8622), .B2(n8838), .C1(n8620), 
        .C2(n8840), .ZN(n10102) );
  NOR2_X1 U8876 ( .A1(n10102), .A2(n10092), .ZN(n7254) );
  AOI211_X1 U8877 ( .C1(n10105), .C2(n8819), .A(n7255), .B(n7254), .ZN(n7256)
         );
  INV_X1 U8878 ( .A(n7256), .ZN(P2_U3230) );
  INV_X1 U8879 ( .A(n7257), .ZN(n7258) );
  NAND3_X1 U8880 ( .A1(n7260), .A2(n7259), .A3(n7258), .ZN(n7261) );
  NOR2_X1 U8881 ( .A1(n4315), .A2(n9954), .ZN(n9568) );
  INV_X1 U8882 ( .A(n9568), .ZN(n7273) );
  NOR3_X1 U8883 ( .A1(n7264), .A2(n7263), .A3(n7262), .ZN(n7265) );
  AOI21_X1 U8884 ( .B1(n9898), .B2(P1_REG3_REG_0__SCAN_IN), .A(n7265), .ZN(
        n7266) );
  NOR2_X1 U8885 ( .A1(n7266), .A2(n4315), .ZN(n7267) );
  AOI21_X1 U8886 ( .B1(n4315), .B2(P1_REG2_REG_0__SCAN_IN), .A(n7267), .ZN(
        n7272) );
  NOR2_X2 U8887 ( .A1(n4315), .A2(n7268), .ZN(n9635) );
  NOR2_X1 U8888 ( .A1(n9904), .A2(n9889), .ZN(n7522) );
  OAI21_X1 U8889 ( .B1(n7522), .B2(n9901), .A(n7270), .ZN(n7271) );
  OAI211_X1 U8890 ( .C1(n7299), .C2(n7273), .A(n7272), .B(n7271), .ZN(P1_U3293) );
  INV_X1 U8891 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n7278) );
  NAND2_X1 U8892 ( .A1(n7274), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n7275) );
  AOI21_X1 U8893 ( .B1(n7278), .B2(n7277), .A(n7493), .ZN(n7292) );
  XNOR2_X1 U8894 ( .A(n7492), .B(n7482), .ZN(n7281) );
  NAND2_X1 U8895 ( .A1(P2_REG1_REG_11__SCAN_IN), .A2(n7281), .ZN(n7484) );
  OAI21_X1 U8896 ( .B1(P2_REG1_REG_11__SCAN_IN), .B2(n7281), .A(n7484), .ZN(
        n7284) );
  AND2_X1 U8897 ( .A1(P2_U3151), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n7834) );
  AOI21_X1 U8898 ( .B1(n10049), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n7834), .ZN(
        n7282) );
  OAI21_X1 U8899 ( .B1(n7483), .B2(n8712), .A(n7282), .ZN(n7283) );
  AOI21_X1 U8900 ( .B1(n7284), .B2(n10058), .A(n7283), .ZN(n7291) );
  NAND2_X1 U8901 ( .A1(n7286), .A2(n7285), .ZN(n7288) );
  MUX2_X1 U8902 ( .A(P2_REG1_REG_11__SCAN_IN), .B(P2_REG2_REG_11__SCAN_IN), 
        .S(n8697), .Z(n7474) );
  XNOR2_X1 U8903 ( .A(n7474), .B(n7492), .ZN(n7287) );
  NAND2_X1 U8904 ( .A1(n7288), .A2(n7287), .ZN(n7477) );
  OAI21_X1 U8905 ( .B1(n7288), .B2(n7287), .A(n7477), .ZN(n7289) );
  NAND2_X1 U8906 ( .A1(n7289), .A2(n10057), .ZN(n7290) );
  OAI211_X1 U8907 ( .C1(n7292), .C2(n10064), .A(n7291), .B(n7290), .ZN(
        P2_U3193) );
  INV_X1 U8908 ( .A(n7293), .ZN(n7296) );
  INV_X1 U8909 ( .A(n9349), .ZN(n9343) );
  OAI222_X1 U8910 ( .A1(n8071), .A2(n7294), .B1(n9797), .B2(n7296), .C1(
        P1_U3086), .C2(n9343), .ZN(P1_U3338) );
  OAI222_X1 U8911 ( .A1(n8678), .A2(P2_U3151), .B1(n9022), .B2(n7296), .C1(
        n7295), .C2(n9015), .ZN(P2_U3278) );
  XOR2_X1 U8912 ( .A(n7218), .B(n4401), .Z(n7302) );
  OAI21_X1 U8913 ( .B1(n7297), .B2(n7218), .A(n7298), .ZN(n9918) );
  INV_X1 U8914 ( .A(n9620), .ZN(n7641) );
  OAI22_X1 U8915 ( .A1(n7299), .A2(n9952), .B1(n7330), .B2(n9954), .ZN(n7300)
         );
  AOI21_X1 U8916 ( .B1(n9918), .B2(n7641), .A(n7300), .ZN(n7301) );
  OAI21_X1 U8917 ( .B1(n7302), .B2(n9962), .A(n7301), .ZN(n9916) );
  INV_X1 U8918 ( .A(n9916), .ZN(n7310) );
  INV_X1 U8919 ( .A(n9632), .ZN(n7651) );
  OAI211_X1 U8920 ( .C1(n7305), .C2(n7219), .A(n7304), .B(n9573), .ZN(n9915)
         );
  AOI22_X1 U8921 ( .A1(n4315), .A2(P1_REG2_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(n9898), .ZN(n7307) );
  NAND2_X1 U8922 ( .A1(n9901), .A2(n5282), .ZN(n7306) );
  OAI211_X1 U8923 ( .C1(n9904), .C2(n9915), .A(n7307), .B(n7306), .ZN(n7308)
         );
  AOI21_X1 U8924 ( .B1(n7651), .B2(n9918), .A(n7308), .ZN(n7309) );
  OAI21_X1 U8925 ( .B1(n7310), .B2(n4315), .A(n7309), .ZN(P1_U3291) );
  NAND2_X1 U8926 ( .A1(n7319), .A2(n7382), .ZN(n8271) );
  NAND2_X1 U8927 ( .A1(n8620), .A2(n6853), .ZN(n7375) );
  NAND2_X1 U8928 ( .A1(n7388), .A2(n7375), .ZN(n7313) );
  XNOR2_X1 U8929 ( .A(n8619), .B(n10112), .ZN(n8426) );
  XNOR2_X1 U8930 ( .A(n7313), .B(n8426), .ZN(n7314) );
  INV_X1 U8931 ( .A(n7314), .ZN(n10113) );
  NAND2_X1 U8932 ( .A1(n7314), .A2(n10084), .ZN(n7323) );
  NAND2_X1 U8933 ( .A1(n7315), .A2(n7072), .ZN(n7377) );
  NAND2_X1 U8934 ( .A1(n7319), .A2(n6853), .ZN(n7316) );
  AND2_X1 U8935 ( .A1(n7377), .A2(n7316), .ZN(n7365) );
  NAND2_X1 U8936 ( .A1(n7378), .A2(n7365), .ZN(n7317) );
  OR2_X1 U8937 ( .A1(n7319), .A2(n6853), .ZN(n7362) );
  AND2_X1 U8938 ( .A1(n7317), .A2(n7362), .ZN(n7318) );
  XNOR2_X1 U8939 ( .A(n7318), .B(n8426), .ZN(n7321) );
  OAI22_X1 U8940 ( .A1(n10077), .A2(n10074), .B1(n7319), .B2(n10076), .ZN(
        n7320) );
  AOI21_X1 U8941 ( .B1(n7321), .B2(n8843), .A(n7320), .ZN(n7322) );
  NAND2_X1 U8942 ( .A1(n7323), .A2(n7322), .ZN(n10114) );
  MUX2_X1 U8943 ( .A(n10114), .B(P2_REG2_REG_5__SCAN_IN), .S(n10092), .Z(n7324) );
  INV_X1 U8944 ( .A(n7324), .ZN(n7327) );
  AOI22_X1 U8945 ( .A1(n10085), .A2(n7366), .B1(n10087), .B2(n7325), .ZN(n7326) );
  OAI211_X1 U8946 ( .C1(n10113), .C2(n8726), .A(n7327), .B(n7326), .ZN(
        P2_U3228) );
  XNOR2_X1 U8947 ( .A(n7333), .B(n7328), .ZN(n7329) );
  OAI222_X1 U8948 ( .A1(n9954), .A2(n7597), .B1(n9952), .B2(n7330), .C1(n7329), 
        .C2(n9962), .ZN(n9922) );
  INV_X1 U8949 ( .A(n9922), .ZN(n7344) );
  NAND2_X1 U8950 ( .A1(n7330), .A2(n7467), .ZN(n7331) );
  NAND2_X1 U8951 ( .A1(n7332), .A2(n7331), .ZN(n7334) );
  OAI21_X1 U8952 ( .B1(n7334), .B2(n7333), .A(n7350), .ZN(n9924) );
  OR2_X1 U8953 ( .A1(n4315), .A2(n9620), .ZN(n7335) );
  INV_X1 U8954 ( .A(n7439), .ZN(n7336) );
  OAI211_X1 U8955 ( .C1(n9921), .C2(n7337), .A(n7336), .B(n9573), .ZN(n9920)
         );
  AOI22_X1 U8956 ( .A1(n4315), .A2(P1_REG2_REG_4__SCAN_IN), .B1(n7338), .B2(
        n9898), .ZN(n7341) );
  NAND2_X1 U8957 ( .A1(n9901), .A2(n7339), .ZN(n7340) );
  OAI211_X1 U8958 ( .C1(n9920), .C2(n9904), .A(n7341), .B(n7340), .ZN(n7342)
         );
  AOI21_X1 U8959 ( .B1(n9924), .B2(n9907), .A(n7342), .ZN(n7343) );
  OAI21_X1 U8960 ( .B1(n7344), .B2(n4315), .A(n7343), .ZN(P1_U3289) );
  XNOR2_X1 U8961 ( .A(n7506), .B(n7352), .ZN(n7345) );
  NAND2_X1 U8962 ( .A1(n7345), .A2(n9876), .ZN(n7348) );
  OAI22_X1 U8963 ( .A1(n7940), .A2(n9954), .B1(n7597), .B2(n9952), .ZN(n7346)
         );
  INV_X1 U8964 ( .A(n7346), .ZN(n7347) );
  NAND2_X1 U8965 ( .A1(n7348), .A2(n7347), .ZN(n9928) );
  INV_X1 U8966 ( .A(n9928), .ZN(n7358) );
  NAND2_X1 U8967 ( .A1(n7418), .A2(n9921), .ZN(n7349) );
  NAND2_X1 U8968 ( .A1(n7597), .A2(n7444), .ZN(n7351) );
  OAI21_X1 U8969 ( .B1(n7353), .B2(n7352), .A(n7510), .ZN(n9930) );
  OAI211_X1 U8970 ( .C1(n7437), .C2(n9927), .A(n9573), .B(n7517), .ZN(n9926)
         );
  AOI22_X1 U8971 ( .A1(n4315), .A2(P1_REG2_REG_6__SCAN_IN), .B1(n7601), .B2(
        n9898), .ZN(n7355) );
  NAND2_X1 U8972 ( .A1(n9901), .A2(n7600), .ZN(n7354) );
  OAI211_X1 U8973 ( .C1(n9926), .C2(n9904), .A(n7355), .B(n7354), .ZN(n7356)
         );
  AOI21_X1 U8974 ( .B1(n9930), .B2(n9907), .A(n7356), .ZN(n7357) );
  OAI21_X1 U8975 ( .B1(n7358), .B2(n4315), .A(n7357), .ZN(P1_U3287) );
  NAND2_X1 U8976 ( .A1(n8619), .A2(n10112), .ZN(n8275) );
  AND2_X1 U8977 ( .A1(n7375), .A2(n8275), .ZN(n8278) );
  NAND2_X1 U8978 ( .A1(n7388), .A2(n8278), .ZN(n7360) );
  NAND2_X1 U8979 ( .A1(n7359), .A2(n7366), .ZN(n7389) );
  NAND2_X1 U8980 ( .A1(n7360), .A2(n7389), .ZN(n7361) );
  NAND2_X1 U8981 ( .A1(n10077), .A2(n7393), .ZN(n8249) );
  AND2_X1 U8982 ( .A1(n8249), .A2(n8273), .ZN(n7369) );
  INV_X1 U8983 ( .A(n7369), .ZN(n8425) );
  XNOR2_X1 U8984 ( .A(n7361), .B(n8425), .ZN(n10121) );
  NOR2_X1 U8985 ( .A1(n8619), .A2(n7366), .ZN(n7364) );
  NAND2_X1 U8986 ( .A1(n8619), .A2(n7366), .ZN(n7367) );
  NAND2_X1 U8987 ( .A1(n7368), .A2(n7367), .ZN(n7395) );
  XNOR2_X1 U8988 ( .A(n7395), .B(n7369), .ZN(n7370) );
  INV_X1 U8989 ( .A(n7396), .ZN(n8617) );
  AOI222_X1 U8990 ( .A1(n8843), .A2(n7370), .B1(n8617), .B2(n8840), .C1(n8619), 
        .C2(n8838), .ZN(n10117) );
  MUX2_X1 U8991 ( .A(n7371), .B(n10117), .S(n8867), .Z(n7374) );
  AOI22_X1 U8992 ( .A1(n10085), .A2(n7393), .B1(n10087), .B2(n7372), .ZN(n7373) );
  OAI211_X1 U8993 ( .C1(n8872), .C2(n10121), .A(n7374), .B(n7373), .ZN(
        P2_U3227) );
  AND2_X1 U8994 ( .A1(n8271), .A2(n7375), .ZN(n8423) );
  XOR2_X1 U8995 ( .A(n7376), .B(n8423), .Z(n10108) );
  NAND2_X1 U8996 ( .A1(n7378), .A2(n7377), .ZN(n7379) );
  XOR2_X1 U8997 ( .A(n8423), .B(n7379), .Z(n7380) );
  AOI222_X1 U8998 ( .A1(n8843), .A2(n7380), .B1(n8621), .B2(n8838), .C1(n8619), 
        .C2(n8840), .ZN(n10107) );
  MUX2_X1 U8999 ( .A(n6674), .B(n10107), .S(n10091), .Z(n7384) );
  AOI22_X1 U9000 ( .A1(n10085), .A2(n7382), .B1(n10087), .B2(n7381), .ZN(n7383) );
  OAI211_X1 U9001 ( .C1(n8872), .C2(n10108), .A(n7384), .B(n7383), .ZN(
        P2_U3229) );
  INV_X1 U9002 ( .A(n7385), .ZN(n7424) );
  INV_X1 U9003 ( .A(n8688), .ZN(n8700) );
  OAI222_X1 U9004 ( .A1(n9015), .A2(n7386), .B1(n9022), .B2(n7424), .C1(
        P2_U3151), .C2(n8700), .ZN(P2_U3277) );
  AND2_X1 U9005 ( .A1(n8278), .A2(n8273), .ZN(n7387) );
  OR2_X1 U9006 ( .A1(n10125), .A2(n7396), .ZN(n7654) );
  NAND2_X1 U9007 ( .A1(n10125), .A2(n7396), .ZN(n8290) );
  INV_X1 U9008 ( .A(n10078), .ZN(n7390) );
  AND2_X1 U9009 ( .A1(n7389), .A2(n8249), .ZN(n8282) );
  OR2_X1 U9010 ( .A1(n8281), .A2(n8282), .ZN(n10069) );
  AND2_X1 U9011 ( .A1(n10069), .A2(n7390), .ZN(n7391) );
  NAND2_X1 U9012 ( .A1(n10071), .A2(n7654), .ZN(n7392) );
  NOR2_X1 U9013 ( .A1(n7658), .A2(n10075), .ZN(n8286) );
  INV_X1 U9014 ( .A(n8286), .ZN(n7655) );
  AND2_X1 U9015 ( .A1(n7658), .A2(n10075), .ZN(n8287) );
  INV_X1 U9016 ( .A(n8287), .ZN(n8291) );
  XNOR2_X1 U9017 ( .A(n7392), .B(n8429), .ZN(n7431) );
  NOR2_X1 U9018 ( .A1(n10077), .A2(n10119), .ZN(n7394) );
  INV_X1 U9019 ( .A(n10125), .ZN(n7397) );
  XOR2_X1 U9020 ( .A(n8429), .B(n7657), .Z(n7398) );
  AOI222_X1 U9021 ( .A1(n8843), .A2(n7398), .B1(n8617), .B2(n8838), .C1(n8615), 
        .C2(n8840), .ZN(n7426) );
  OAI21_X1 U9022 ( .B1(n10120), .B2(n7431), .A(n7426), .ZN(n7461) );
  INV_X1 U9023 ( .A(n7461), .ZN(n7410) );
  NAND2_X1 U9024 ( .A1(n7400), .A2(n7399), .ZN(n7406) );
  INV_X1 U9025 ( .A(n7401), .ZN(n7402) );
  NAND2_X1 U9026 ( .A1(n6223), .A2(n7402), .ZN(n7404) );
  NAND2_X1 U9027 ( .A1(n7404), .A2(n7403), .ZN(n7405) );
  AND2_X1 U9028 ( .A1(n7406), .A2(n7405), .ZN(n7408) );
  AOI22_X1 U9029 ( .A1(n8927), .A2(n7658), .B1(n10156), .B2(
        P2_REG1_REG_8__SCAN_IN), .ZN(n7409) );
  OAI21_X1 U9030 ( .B1(n7410), .B2(n10156), .A(n7409), .ZN(P2_U3467) );
  OAI22_X1 U9031 ( .A1(n7597), .A2(n9113), .B1(n7444), .B2(n6864), .ZN(n7417)
         );
  AOI22_X1 U9032 ( .A1(n9270), .A2(n9049), .B1(n9900), .B2(n9044), .ZN(n7413)
         );
  XNOR2_X1 U9033 ( .A(n7413), .B(n9030), .ZN(n7415) );
  NAND2_X1 U9034 ( .A1(n7414), .A2(n7415), .ZN(n7589) );
  AOI21_X1 U9035 ( .B1(n7417), .B2(n7416), .A(n7591), .ZN(n7423) );
  NAND2_X1 U9036 ( .A1(P1_U3086), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n9306) );
  INV_X1 U9037 ( .A(n9306), .ZN(n7420) );
  OAI22_X1 U9038 ( .A1(n7746), .A2(n9241), .B1(n9255), .B2(n7418), .ZN(n7419)
         );
  AOI211_X1 U9039 ( .C1(n9900), .C2(n9257), .A(n7420), .B(n7419), .ZN(n7422)
         );
  NAND2_X1 U9040 ( .A1(n9252), .A2(n9899), .ZN(n7421) );
  OAI211_X1 U9041 ( .C1(n7423), .C2(n9259), .A(n7422), .B(n7421), .ZN(P1_U3227) );
  INV_X1 U9042 ( .A(n9358), .ZN(n9346) );
  OAI222_X1 U9043 ( .A1(n8071), .A2(n7425), .B1(n9346), .B2(P1_U3086), .C1(
        n9797), .C2(n7424), .ZN(P1_U3337) );
  MUX2_X1 U9044 ( .A(n7427), .B(n7426), .S(n10091), .Z(n7430) );
  AOI22_X1 U9045 ( .A1(n10085), .A2(n7658), .B1(n10087), .B2(n7428), .ZN(n7429) );
  OAI211_X1 U9046 ( .C1(n7431), .C2(n8872), .A(n7430), .B(n7429), .ZN(P2_U3225) );
  OAI21_X1 U9047 ( .B1(n7433), .B2(n7435), .A(n7432), .ZN(n9908) );
  INV_X1 U9048 ( .A(n9908), .ZN(n7440) );
  XNOR2_X1 U9049 ( .A(n7435), .B(n7434), .ZN(n7436) );
  AOI222_X1 U9050 ( .A1(n9876), .A2(n7436), .B1(n9271), .B2(n9879), .C1(n9269), 
        .C2(n9880), .ZN(n9910) );
  INV_X1 U9051 ( .A(n7437), .ZN(n7438) );
  OAI211_X1 U9052 ( .C1(n7444), .C2(n7439), .A(n7438), .B(n9573), .ZN(n9905)
         );
  OAI211_X1 U9053 ( .C1(n9741), .C2(n7440), .A(n9910), .B(n9905), .ZN(n7446)
         );
  OAI22_X1 U9054 ( .A1(n9788), .A2(n7444), .B1(n9968), .B2(n5319), .ZN(n7441)
         );
  AOI21_X1 U9055 ( .B1(n7446), .B2(n9968), .A(n7441), .ZN(n7442) );
  INV_X1 U9056 ( .A(n7442), .ZN(P1_U3468) );
  INV_X1 U9057 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n7443) );
  OAI22_X1 U9058 ( .A1(n9747), .A2(n7444), .B1(n9983), .B2(n7443), .ZN(n7445)
         );
  AOI21_X1 U9059 ( .B1(n7446), .B2(n9983), .A(n7445), .ZN(n7447) );
  INV_X1 U9060 ( .A(n7447), .ZN(P1_U3527) );
  NOR2_X1 U9061 ( .A1(n4315), .A2(n9952), .ZN(n9421) );
  AOI22_X1 U9062 ( .A1(n4315), .A2(P1_REG2_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(n9898), .ZN(n7448) );
  OAI21_X1 U9063 ( .B1(n9630), .B2(n8082), .A(n7448), .ZN(n7454) );
  INV_X1 U9064 ( .A(n7449), .ZN(n7452) );
  AOI22_X1 U9065 ( .A1(n7450), .A2(n9635), .B1(n9568), .B2(n7225), .ZN(n7451)
         );
  OAI21_X1 U9066 ( .B1(n9894), .B2(n7452), .A(n7451), .ZN(n7453) );
  AOI211_X1 U9067 ( .C1(n9421), .C2(n7455), .A(n7454), .B(n7453), .ZN(n7456)
         );
  OAI21_X1 U9068 ( .B1(n4315), .B2(n7457), .A(n7456), .ZN(P1_U3292) );
  INV_X1 U9069 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n7458) );
  OAI22_X1 U9070 ( .A1(n7459), .A2(n8969), .B1(n10142), .B2(n7458), .ZN(n7460)
         );
  AOI21_X1 U9071 ( .B1(n7461), .B2(n10142), .A(n7460), .ZN(n7462) );
  INV_X1 U9072 ( .A(n7462), .ZN(P2_U3414) );
  NAND2_X1 U9073 ( .A1(n7522), .A2(n7463), .ZN(n7466) );
  AOI22_X1 U9074 ( .A1(n4315), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n9898), .B2(
        n7464), .ZN(n7465) );
  OAI211_X1 U9075 ( .C1(n7467), .C2(n9630), .A(n7466), .B(n7465), .ZN(n7468)
         );
  AOI21_X1 U9076 ( .B1(n9907), .B2(n7469), .A(n7468), .ZN(n7470) );
  OAI21_X1 U9077 ( .B1(n7471), .B2(n4315), .A(n7470), .ZN(P1_U3290) );
  INV_X1 U9078 ( .A(n7472), .ZN(n8471) );
  OAI222_X1 U9079 ( .A1(n8711), .A2(P2_U3151), .B1(n9022), .B2(n8471), .C1(
        n7473), .C2(n9015), .ZN(P2_U3276) );
  INV_X1 U9080 ( .A(n7474), .ZN(n7475) );
  NAND2_X1 U9081 ( .A1(n7475), .A2(n7492), .ZN(n7476) );
  NAND2_X1 U9082 ( .A1(n7477), .A2(n7476), .ZN(n8659) );
  INV_X1 U9083 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n7811) );
  INV_X1 U9084 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n7717) );
  MUX2_X1 U9085 ( .A(n7811), .B(n7717), .S(n8697), .Z(n7478) );
  AND2_X1 U9086 ( .A1(n7478), .A2(n7488), .ZN(n8658) );
  INV_X1 U9087 ( .A(n8658), .ZN(n7480) );
  INV_X1 U9088 ( .A(n7478), .ZN(n7479) );
  NAND2_X1 U9089 ( .A1(n7479), .A2(n8637), .ZN(n8660) );
  NAND2_X1 U9090 ( .A1(n7480), .A2(n8660), .ZN(n7481) );
  XNOR2_X1 U9091 ( .A(n8659), .B(n7481), .ZN(n7502) );
  AOI22_X1 U9092 ( .A1(P2_REG1_REG_12__SCAN_IN), .A2(n8637), .B1(n7488), .B2(
        n7811), .ZN(n7487) );
  NAND2_X1 U9093 ( .A1(n7483), .A2(n7482), .ZN(n7485) );
  NAND2_X1 U9094 ( .A1(n7485), .A2(n7484), .ZN(n7486) );
  OAI21_X1 U9095 ( .B1(n7487), .B2(n7486), .A(n8626), .ZN(n7500) );
  INV_X1 U9096 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n7557) );
  NAND2_X1 U9097 ( .A1(n10051), .A2(n7488), .ZN(n7489) );
  NAND2_X1 U9098 ( .A1(P2_U3151), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n7885) );
  OAI211_X1 U9099 ( .C1(n7557), .C2(n8654), .A(n7489), .B(n7885), .ZN(n7499)
         );
  NOR2_X1 U9100 ( .A1(n7492), .A2(n7491), .ZN(n7494) );
  NAND2_X1 U9101 ( .A1(P2_REG2_REG_12__SCAN_IN), .A2(n8637), .ZN(n7495) );
  OAI21_X1 U9102 ( .B1(P2_REG2_REG_12__SCAN_IN), .B2(n8637), .A(n7495), .ZN(
        n7496) );
  AOI21_X1 U9103 ( .B1(n4389), .B2(n7496), .A(n8636), .ZN(n7497) );
  NOR2_X1 U9104 ( .A1(n7497), .A2(n10064), .ZN(n7498) );
  AOI211_X1 U9105 ( .C1(n10058), .C2(n7500), .A(n7499), .B(n7498), .ZN(n7501)
         );
  OAI21_X1 U9106 ( .B1(n9989), .B2(n7502), .A(n7501), .ZN(P2_U3194) );
  INV_X1 U9107 ( .A(n7503), .ZN(n7505) );
  OAI21_X1 U9108 ( .B1(n7506), .B2(n7505), .A(n7504), .ZN(n7507) );
  NAND2_X1 U9109 ( .A1(n7507), .A2(n7508), .ZN(n7636) );
  OAI21_X1 U9110 ( .B1(n7508), .B2(n7507), .A(n7636), .ZN(n7516) );
  OAI22_X1 U9111 ( .A1(n9174), .A2(n9954), .B1(n7746), .B2(n9952), .ZN(n7515)
         );
  NAND2_X1 U9112 ( .A1(n7746), .A2(n9927), .ZN(n7509) );
  OR2_X1 U9113 ( .A1(n7512), .A2(n7511), .ZN(n7513) );
  NOR2_X1 U9114 ( .A1(n7771), .A2(n9620), .ZN(n7514) );
  AOI211_X1 U9115 ( .C1(n9876), .C2(n7516), .A(n7515), .B(n7514), .ZN(n7770)
         );
  NAND2_X1 U9116 ( .A1(n7517), .A2(n7767), .ZN(n7518) );
  AND2_X1 U9117 ( .A1(n7645), .A2(n7518), .ZN(n7768) );
  AOI22_X1 U9118 ( .A1(n4315), .A2(P1_REG2_REG_7__SCAN_IN), .B1(n7749), .B2(
        n9898), .ZN(n7519) );
  OAI21_X1 U9119 ( .B1(n9630), .B2(n7743), .A(n7519), .ZN(n7521) );
  NOR2_X1 U9120 ( .A1(n7771), .A2(n9632), .ZN(n7520) );
  AOI211_X1 U9121 ( .C1(n7768), .C2(n7522), .A(n7521), .B(n7520), .ZN(n7523)
         );
  OAI21_X1 U9122 ( .B1(n7770), .B2(n4315), .A(n7523), .ZN(P1_U3286) );
  INV_X1 U9123 ( .A(n7524), .ZN(n7588) );
  INV_X1 U9124 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7525) );
  OAI222_X1 U9125 ( .A1(n9797), .A2(n7588), .B1(P1_U3086), .B2(n7526), .C1(
        n7525), .C2(n8071), .ZN(P1_U3335) );
  NOR2_X1 U9126 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n7570) );
  NOR2_X1 U9127 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n7568) );
  NOR2_X1 U9128 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n7566) );
  NOR2_X1 U9129 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n7564) );
  NOR2_X1 U9130 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n7562) );
  NOR2_X1 U9131 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n7560) );
  INV_X1 U9132 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n7556) );
  NOR2_X1 U9133 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n7549) );
  NOR2_X1 U9134 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n7546) );
  NOR2_X1 U9135 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n7543) );
  NOR2_X1 U9136 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n7540) );
  NOR2_X1 U9137 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n7537) );
  NAND2_X1 U9138 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n7535) );
  XNOR2_X1 U9139 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(n7527), .ZN(n10194) );
  NAND2_X1 U9140 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n7533) );
  AOI21_X1 U9141 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(P2_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10159) );
  INV_X1 U9142 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n7529) );
  NAND2_X1 U9143 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .ZN(n7528) );
  NOR2_X1 U9144 ( .A1(n7529), .A2(n7528), .ZN(n10160) );
  NOR2_X1 U9145 ( .A1(P2_ADDR_REG_1__SCAN_IN), .A2(n10160), .ZN(n7530) );
  NOR2_X1 U9146 ( .A1(n10159), .A2(n7530), .ZN(n10192) );
  INV_X1 U9147 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n7531) );
  XNOR2_X1 U9148 ( .A(n7531), .B(P1_ADDR_REG_2__SCAN_IN), .ZN(n10191) );
  NAND2_X1 U9149 ( .A1(n10192), .A2(n10191), .ZN(n7532) );
  NAND2_X1 U9150 ( .A1(n7533), .A2(n7532), .ZN(n10193) );
  NAND2_X1 U9151 ( .A1(n10194), .A2(n10193), .ZN(n7534) );
  NAND2_X1 U9152 ( .A1(n7535), .A2(n7534), .ZN(n10196) );
  XNOR2_X1 U9153 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10195) );
  NOR2_X1 U9154 ( .A1(n10196), .A2(n10195), .ZN(n7536) );
  NOR2_X1 U9155 ( .A1(n7537), .A2(n7536), .ZN(n10184) );
  XOR2_X1 U9156 ( .A(n7538), .B(P1_ADDR_REG_5__SCAN_IN), .Z(n10183) );
  NOR2_X1 U9157 ( .A1(n10184), .A2(n10183), .ZN(n7539) );
  NOR2_X1 U9158 ( .A1(n7540), .A2(n7539), .ZN(n10182) );
  INV_X1 U9159 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n9321) );
  AOI22_X1 U9160 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(n9321), .B1(
        P1_ADDR_REG_6__SCAN_IN), .B2(n7541), .ZN(n10181) );
  NOR2_X1 U9161 ( .A1(n10182), .A2(n10181), .ZN(n7542) );
  NOR2_X1 U9162 ( .A1(n7543), .A2(n7542), .ZN(n10188) );
  INV_X1 U9163 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n9334) );
  AOI22_X1 U9164 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n9334), .B1(
        P1_ADDR_REG_7__SCAN_IN), .B2(n7544), .ZN(n10187) );
  NOR2_X1 U9165 ( .A1(n10188), .A2(n10187), .ZN(n7545) );
  NOR2_X1 U9166 ( .A1(n7546), .A2(n7545), .ZN(n10190) );
  XOR2_X1 U9167 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(n7547), .Z(n10189) );
  NOR2_X1 U9168 ( .A1(n10190), .A2(n10189), .ZN(n7548) );
  NOR2_X1 U9169 ( .A1(n7549), .A2(n7548), .ZN(n10186) );
  AOI22_X1 U9170 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n7551), .B1(
        P1_ADDR_REG_9__SCAN_IN), .B2(n7552), .ZN(n10185) );
  NOR2_X1 U9171 ( .A1(n10186), .A2(n10185), .ZN(n7550) );
  AOI21_X1 U9172 ( .B1(n7552), .B2(n7551), .A(n7550), .ZN(n10180) );
  AOI22_X1 U9173 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(n9812), .B1(
        P1_ADDR_REG_10__SCAN_IN), .B2(n7554), .ZN(n10179) );
  NOR2_X1 U9174 ( .A1(n10180), .A2(n10179), .ZN(n7553) );
  AOI21_X1 U9175 ( .B1(n7554), .B2(n9812), .A(n7553), .ZN(n10178) );
  AOI22_X1 U9176 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(n9824), .B1(
        P1_ADDR_REG_11__SCAN_IN), .B2(n7556), .ZN(n10177) );
  NOR2_X1 U9177 ( .A1(n10178), .A2(n10177), .ZN(n7555) );
  AOI21_X1 U9178 ( .B1(n7556), .B2(n9824), .A(n7555), .ZN(n10176) );
  INV_X1 U9179 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n7558) );
  AOI22_X1 U9180 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(n7558), .B1(
        P1_ADDR_REG_12__SCAN_IN), .B2(n7557), .ZN(n10175) );
  NOR2_X1 U9181 ( .A1(n10176), .A2(n10175), .ZN(n7559) );
  NOR2_X1 U9182 ( .A1(n7560), .A2(n7559), .ZN(n10174) );
  INV_X1 U9183 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n9836) );
  XOR2_X1 U9184 ( .A(P2_ADDR_REG_13__SCAN_IN), .B(n9836), .Z(n10173) );
  NOR2_X1 U9185 ( .A1(n10174), .A2(n10173), .ZN(n7561) );
  NOR2_X1 U9186 ( .A1(n7562), .A2(n7561), .ZN(n10172) );
  XOR2_X1 U9187 ( .A(P2_ADDR_REG_14__SCAN_IN), .B(n9855), .Z(n10171) );
  NOR2_X1 U9188 ( .A1(n10172), .A2(n10171), .ZN(n7563) );
  NOR2_X1 U9189 ( .A1(n7564), .A2(n7563), .ZN(n10170) );
  INV_X1 U9190 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n9871) );
  XOR2_X1 U9191 ( .A(P2_ADDR_REG_15__SCAN_IN), .B(n9871), .Z(n10169) );
  NOR2_X1 U9192 ( .A1(n10170), .A2(n10169), .ZN(n7565) );
  NOR2_X1 U9193 ( .A1(n7566), .A2(n7565), .ZN(n10168) );
  XNOR2_X1 U9194 ( .A(P2_ADDR_REG_16__SCAN_IN), .B(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n10167) );
  NOR2_X1 U9195 ( .A1(n10168), .A2(n10167), .ZN(n7567) );
  NOR2_X1 U9196 ( .A1(n7568), .A2(n7567), .ZN(n10166) );
  XNOR2_X1 U9197 ( .A(P2_ADDR_REG_17__SCAN_IN), .B(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n10165) );
  NOR2_X1 U9198 ( .A1(n10166), .A2(n10165), .ZN(n7569) );
  NOR2_X1 U9199 ( .A1(n7570), .A2(n7569), .ZN(n7571) );
  AND2_X1 U9200 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n7571), .ZN(n10162) );
  NOR2_X1 U9201 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(n10162), .ZN(n7572) );
  NOR2_X1 U9202 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n7571), .ZN(n10163) );
  NOR2_X1 U9203 ( .A1(n7572), .A2(n10163), .ZN(n7574) );
  XNOR2_X1 U9204 ( .A(P1_ADDR_REG_19__SCAN_IN), .B(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n7573) );
  XNOR2_X1 U9205 ( .A(n7574), .B(n7573), .ZN(ADD_1068_U4) );
  OAI22_X1 U9206 ( .A1(n7576), .A2(n8616), .B1(n6318), .B2(n7575), .ZN(n7579)
         );
  XNOR2_X1 U9207 ( .A(n7577), .B(n7675), .ZN(n7578) );
  XNOR2_X1 U9208 ( .A(n7579), .B(n7578), .ZN(n7586) );
  NAND2_X1 U9209 ( .A1(n8598), .A2(n7665), .ZN(n7583) );
  OR2_X1 U9210 ( .A1(n8595), .A2(n10075), .ZN(n7582) );
  NAND2_X1 U9211 ( .A1(n8593), .A2(n8614), .ZN(n7581) );
  NAND4_X1 U9212 ( .A1(n7583), .A2(n7582), .A3(n7581), .A4(n7580), .ZN(n7584)
         );
  AOI21_X1 U9213 ( .B1(n10134), .B2(n8585), .A(n7584), .ZN(n7585) );
  OAI21_X1 U9214 ( .B1(n7586), .B2(n8573), .A(n7585), .ZN(P2_U3171) );
  OAI222_X1 U9215 ( .A1(P2_U3151), .A2(n8452), .B1(n9022), .B2(n7588), .C1(
        n7587), .C2(n9015), .ZN(P2_U3275) );
  INV_X1 U9216 ( .A(n7589), .ZN(n7590) );
  OAI22_X1 U9217 ( .A1(n7746), .A2(n6864), .B1(n9927), .B2(n4406), .ZN(n7592)
         );
  XNOR2_X1 U9218 ( .A(n7592), .B(n9030), .ZN(n7594) );
  OAI22_X1 U9219 ( .A1(n7746), .A2(n9113), .B1(n9927), .B2(n6864), .ZN(n7593)
         );
  OR2_X1 U9220 ( .A1(n7594), .A2(n7593), .ZN(n7740) );
  INV_X1 U9221 ( .A(n7740), .ZN(n7595) );
  AND2_X1 U9222 ( .A1(n7594), .A2(n7593), .ZN(n7741) );
  NOR2_X1 U9223 ( .A1(n7595), .A2(n7741), .ZN(n7596) );
  XNOR2_X1 U9224 ( .A(n7742), .B(n7596), .ZN(n7604) );
  NAND2_X1 U9225 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n9320) );
  INV_X1 U9226 ( .A(n9320), .ZN(n7599) );
  OAI22_X1 U9227 ( .A1(n7940), .A2(n9241), .B1(n9255), .B2(n7597), .ZN(n7598)
         );
  AOI211_X1 U9228 ( .C1(n7600), .C2(n9257), .A(n7599), .B(n7598), .ZN(n7603)
         );
  NAND2_X1 U9229 ( .A1(n9252), .A2(n7601), .ZN(n7602) );
  OAI211_X1 U9230 ( .C1(n7604), .C2(n9259), .A(n7603), .B(n7602), .ZN(P1_U3239) );
  NOR2_X1 U9231 ( .A1(n7605), .A2(n4399), .ZN(n7607) );
  XNOR2_X1 U9232 ( .A(n7607), .B(n7606), .ZN(n7614) );
  NAND2_X1 U9233 ( .A1(n8598), .A2(n7680), .ZN(n7611) );
  OR2_X1 U9234 ( .A1(n8595), .A2(n7675), .ZN(n7610) );
  NAND2_X1 U9235 ( .A1(n8593), .A2(n8613), .ZN(n7609) );
  NAND4_X1 U9236 ( .A1(n7611), .A2(n7610), .A3(n7609), .A4(n7608), .ZN(n7612)
         );
  AOI21_X1 U9237 ( .B1(n10140), .B2(n8585), .A(n7612), .ZN(n7613) );
  OAI21_X1 U9238 ( .B1(n7614), .B2(n8573), .A(n7613), .ZN(P2_U3157) );
  NAND2_X1 U9239 ( .A1(n7616), .A2(n7615), .ZN(n7631) );
  INV_X1 U9240 ( .A(n7629), .ZN(n7617) );
  AOI21_X1 U9241 ( .B1(n7636), .B2(n7618), .A(n7617), .ZN(n7619) );
  XOR2_X1 U9242 ( .A(n7631), .B(n7619), .Z(n7620) );
  INV_X1 U9243 ( .A(n9174), .ZN(n9267) );
  AOI22_X1 U9244 ( .A1(n7620), .A2(n9876), .B1(n9879), .B2(n9267), .ZN(n9939)
         );
  INV_X1 U9245 ( .A(n9180), .ZN(n7621) );
  OAI22_X1 U9246 ( .A1(n9611), .A2(n7622), .B1(n7621), .B2(n9532), .ZN(n7625)
         );
  XNOR2_X1 U9247 ( .A(n7646), .B(n7984), .ZN(n7623) );
  INV_X1 U9248 ( .A(n9219), .ZN(n9265) );
  AOI22_X1 U9249 ( .A1(n7623), .A2(n9573), .B1(n9880), .B2(n9265), .ZN(n9938)
         );
  NOR2_X1 U9250 ( .A1(n9938), .A2(n9904), .ZN(n7624) );
  AOI211_X1 U9251 ( .C1(n9901), .C2(n7984), .A(n7625), .B(n7624), .ZN(n7634)
         );
  NAND2_X1 U9252 ( .A1(n7940), .A2(n7743), .ZN(n7626) );
  NAND2_X1 U9253 ( .A1(n7629), .A2(n7628), .ZN(n7639) );
  OR2_X1 U9254 ( .A1(n7938), .A2(n9267), .ZN(n7630) );
  NAND2_X1 U9255 ( .A1(n7638), .A2(n7630), .ZN(n7632) );
  OAI21_X1 U9256 ( .B1(n7632), .B2(n7631), .A(n7689), .ZN(n9942) );
  NAND2_X1 U9257 ( .A1(n9942), .A2(n9907), .ZN(n7633) );
  OAI211_X1 U9258 ( .C1(n9939), .C2(n4315), .A(n7634), .B(n7633), .ZN(P1_U3284) );
  NAND2_X1 U9259 ( .A1(n7636), .A2(n7635), .ZN(n7637) );
  XNOR2_X1 U9260 ( .A(n7637), .B(n7639), .ZN(n7644) );
  OAI21_X1 U9261 ( .B1(n7640), .B2(n7639), .A(n7638), .ZN(n9935) );
  NAND2_X1 U9262 ( .A1(n9935), .A2(n7641), .ZN(n7643) );
  AOI22_X1 U9263 ( .A1(n9879), .A2(n9268), .B1(n9266), .B2(n9880), .ZN(n7642)
         );
  OAI211_X1 U9264 ( .C1(n9962), .C2(n7644), .A(n7643), .B(n7642), .ZN(n9933)
         );
  INV_X1 U9265 ( .A(n9933), .ZN(n7653) );
  INV_X1 U9266 ( .A(n7645), .ZN(n7647) );
  INV_X1 U9267 ( .A(n7646), .ZN(n7694) );
  OAI211_X1 U9268 ( .C1(n4593), .C2(n7647), .A(n7694), .B(n9573), .ZN(n9932)
         );
  AOI22_X1 U9269 ( .A1(n4315), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n7939), .B2(
        n9898), .ZN(n7649) );
  NAND2_X1 U9270 ( .A1(n9901), .A2(n7938), .ZN(n7648) );
  OAI211_X1 U9271 ( .C1(n9932), .C2(n9904), .A(n7649), .B(n7648), .ZN(n7650)
         );
  AOI21_X1 U9272 ( .B1(n9935), .B2(n7651), .A(n7650), .ZN(n7652) );
  OAI21_X1 U9273 ( .B1(n7653), .B2(n4315), .A(n7652), .ZN(P1_U3285) );
  AND2_X1 U9274 ( .A1(n7655), .A2(n7654), .ZN(n8295) );
  NAND2_X1 U9275 ( .A1(n10134), .A2(n7675), .ZN(n8292) );
  NAND2_X1 U9276 ( .A1(n8294), .A2(n8292), .ZN(n8289) );
  OAI21_X1 U9277 ( .B1(n7656), .B2(n8430), .A(n7707), .ZN(n10131) );
  NAND2_X1 U9278 ( .A1(n7658), .A2(n8616), .ZN(n7659) );
  XNOR2_X1 U9279 ( .A(n7674), .B(n8289), .ZN(n7664) );
  INV_X1 U9280 ( .A(n10131), .ZN(n7662) );
  OAI22_X1 U9281 ( .A1(n10075), .A2(n10076), .B1(n7838), .B2(n10074), .ZN(
        n7661) );
  AOI21_X1 U9282 ( .B1(n7662), .B2(n10084), .A(n7661), .ZN(n7663) );
  OAI21_X1 U9283 ( .B1(n10080), .B2(n7664), .A(n7663), .ZN(n10132) );
  NAND2_X1 U9284 ( .A1(n10132), .A2(n8867), .ZN(n7670) );
  INV_X1 U9285 ( .A(n7665), .ZN(n7666) );
  OAI22_X1 U9286 ( .A1(n8867), .A2(n7667), .B1(n7666), .B2(n8813), .ZN(n7668)
         );
  AOI21_X1 U9287 ( .B1(n10085), .B2(n10134), .A(n7668), .ZN(n7669) );
  OAI211_X1 U9288 ( .C1(n10131), .C2(n8726), .A(n7670), .B(n7669), .ZN(
        P2_U3224) );
  NAND2_X1 U9289 ( .A1(n7707), .A2(n8294), .ZN(n7672) );
  XNOR2_X1 U9290 ( .A(n10140), .B(n8614), .ZN(n8431) );
  INV_X1 U9291 ( .A(n8431), .ZN(n7671) );
  XNOR2_X1 U9292 ( .A(n7672), .B(n7671), .ZN(n7677) );
  INV_X1 U9293 ( .A(n7677), .ZN(n10137) );
  OR2_X1 U9294 ( .A1(n10134), .A2(n8615), .ZN(n7673) );
  NAND2_X1 U9295 ( .A1(n7674), .A2(n7673), .ZN(n7858) );
  NAND2_X1 U9296 ( .A1(n10134), .A2(n8615), .ZN(n7854) );
  NAND2_X1 U9297 ( .A1(n7858), .A2(n7854), .ZN(n7754) );
  XOR2_X1 U9298 ( .A(n8431), .B(n7754), .Z(n7679) );
  OAI22_X1 U9299 ( .A1(n7675), .A2(n10076), .B1(n7887), .B2(n10074), .ZN(n7676) );
  AOI21_X1 U9300 ( .B1(n7677), .B2(n10084), .A(n7676), .ZN(n7678) );
  OAI21_X1 U9301 ( .B1(n7679), .B2(n10080), .A(n7678), .ZN(n10138) );
  NAND2_X1 U9302 ( .A1(n10138), .A2(n8867), .ZN(n7685) );
  INV_X1 U9303 ( .A(n7680), .ZN(n7681) );
  OAI22_X1 U9304 ( .A1(n8867), .A2(n7682), .B1(n7681), .B2(n8813), .ZN(n7683)
         );
  AOI21_X1 U9305 ( .B1(n10140), .B2(n10085), .A(n7683), .ZN(n7684) );
  OAI211_X1 U9306 ( .C1(n10137), .C2(n8726), .A(n7685), .B(n7684), .ZN(
        P2_U3223) );
  INV_X1 U9307 ( .A(n7724), .ZN(n7686) );
  AOI21_X1 U9308 ( .B1(n7690), .B2(n7687), .A(n7686), .ZN(n7778) );
  INV_X1 U9309 ( .A(n9549), .ZN(n9579) );
  OR2_X1 U9310 ( .A1(n7984), .A2(n9266), .ZN(n7688) );
  OAI21_X1 U9311 ( .B1(n7691), .B2(n7690), .A(n7722), .ZN(n7780) );
  NAND2_X1 U9312 ( .A1(n7780), .A2(n9907), .ZN(n7699) );
  INV_X1 U9313 ( .A(n9421), .ZN(n9587) );
  AOI22_X1 U9314 ( .A1(n4315), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n9091), .B2(
        n9898), .ZN(n7693) );
  NAND2_X1 U9315 ( .A1(n9568), .A2(n9878), .ZN(n7692) );
  OAI211_X1 U9316 ( .C1(n9587), .C2(n9092), .A(n7693), .B(n7692), .ZN(n7697)
         );
  OAI21_X1 U9317 ( .B1(n7694), .B2(n7984), .A(n8000), .ZN(n7695) );
  NAND3_X1 U9318 ( .A1(n7695), .A2(n9573), .A3(n7733), .ZN(n7776) );
  NOR2_X1 U9319 ( .A1(n7776), .A2(n9904), .ZN(n7696) );
  AOI211_X1 U9320 ( .C1(n9901), .C2(n8000), .A(n7697), .B(n7696), .ZN(n7698)
         );
  OAI211_X1 U9321 ( .C1(n7778), .C2(n9579), .A(n7699), .B(n7698), .ZN(P1_U3283) );
  INV_X1 U9322 ( .A(n7700), .ZN(n7704) );
  OAI222_X1 U9323 ( .A1(n9797), .A2(n7704), .B1(P1_U3086), .B2(n7702), .C1(
        n7701), .C2(n8071), .ZN(P1_U3334) );
  OAI222_X1 U9324 ( .A1(P2_U3151), .A2(n7705), .B1(n9022), .B2(n7704), .C1(
        n7703), .C2(n9015), .ZN(P2_U3274) );
  OR2_X1 U9325 ( .A1(n10140), .A2(n7838), .ZN(n8303) );
  AND2_X1 U9326 ( .A1(n8294), .A2(n8303), .ZN(n7706) );
  NAND2_X1 U9327 ( .A1(n10140), .A2(n7838), .ZN(n8302) );
  NAND2_X1 U9328 ( .A1(n7844), .A2(n7887), .ZN(n8307) );
  OR2_X1 U9329 ( .A1(n7844), .A2(n7887), .ZN(n8306) );
  NAND2_X1 U9330 ( .A1(n7708), .A2(n8306), .ZN(n7709) );
  XNOR2_X1 U9331 ( .A(n8312), .B(n8612), .ZN(n8435) );
  NAND2_X1 U9332 ( .A1(n7709), .A2(n8435), .ZN(n7821) );
  OAI21_X1 U9333 ( .B1(n7709), .B2(n8435), .A(n7821), .ZN(n7805) );
  OR2_X1 U9334 ( .A1(n10140), .A2(n8614), .ZN(n7753) );
  AND2_X1 U9335 ( .A1(n7753), .A2(n7710), .ZN(n7851) );
  NAND2_X1 U9336 ( .A1(n7754), .A2(n7851), .ZN(n7824) );
  NAND2_X1 U9337 ( .A1(n10140), .A2(n8614), .ZN(n7755) );
  NAND2_X1 U9338 ( .A1(n7824), .A2(n7823), .ZN(n7712) );
  XNOR2_X1 U9339 ( .A(n7712), .B(n8435), .ZN(n7713) );
  NAND2_X1 U9340 ( .A1(n7713), .A2(n8843), .ZN(n7715) );
  AOI22_X1 U9341 ( .A1(n8613), .A2(n8838), .B1(n8840), .B2(n8611), .ZN(n7714)
         );
  NAND2_X1 U9342 ( .A1(n7715), .A2(n7714), .ZN(n7806) );
  NAND2_X1 U9343 ( .A1(n7806), .A2(n8867), .ZN(n7720) );
  INV_X1 U9344 ( .A(n7889), .ZN(n7716) );
  OAI22_X1 U9345 ( .A1(n8867), .A2(n7717), .B1(n7716), .B2(n8813), .ZN(n7718)
         );
  AOI21_X1 U9346 ( .B1(n8312), .B2(n10085), .A(n7718), .ZN(n7719) );
  OAI211_X1 U9347 ( .C1(n7805), .C2(n8872), .A(n7720), .B(n7719), .ZN(P2_U3221) );
  OR2_X1 U9348 ( .A1(n8000), .A2(n9265), .ZN(n7721) );
  XNOR2_X1 U9349 ( .A(n8024), .B(n7725), .ZN(n7794) );
  INV_X1 U9350 ( .A(n7794), .ZN(n7739) );
  NAND2_X1 U9351 ( .A1(n7724), .A2(n7723), .ZN(n7727) );
  INV_X1 U9352 ( .A(n7725), .ZN(n7726) );
  XNOR2_X1 U9353 ( .A(n7727), .B(n7726), .ZN(n7728) );
  NAND2_X1 U9354 ( .A1(n7728), .A2(n9876), .ZN(n7731) );
  OAI22_X1 U9355 ( .A1(n9953), .A2(n9954), .B1(n9219), .B2(n9952), .ZN(n7729)
         );
  INV_X1 U9356 ( .A(n7729), .ZN(n7730) );
  NAND2_X1 U9357 ( .A1(n7731), .A2(n7730), .ZN(n7792) );
  INV_X1 U9358 ( .A(n9221), .ZN(n7736) );
  INV_X1 U9359 ( .A(n9891), .ZN(n7732) );
  AOI211_X1 U9360 ( .C1(n9221), .C2(n7733), .A(n9889), .B(n7732), .ZN(n7793)
         );
  NAND2_X1 U9361 ( .A1(n7793), .A2(n9635), .ZN(n7735) );
  AOI22_X1 U9362 ( .A1(n4315), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n9216), .B2(
        n9898), .ZN(n7734) );
  OAI211_X1 U9363 ( .C1(n7736), .C2(n9630), .A(n7735), .B(n7734), .ZN(n7737)
         );
  AOI21_X1 U9364 ( .B1(n9611), .B2(n7792), .A(n7737), .ZN(n7738) );
  OAI21_X1 U9365 ( .B1(n7739), .B2(n9894), .A(n7738), .ZN(P1_U3282) );
  OAI22_X1 U9366 ( .A1(n7743), .A2(n6864), .B1(n7940), .B2(n9113), .ZN(n7924)
         );
  NAND2_X1 U9367 ( .A1(n7767), .A2(n9044), .ZN(n7744) );
  OAI21_X1 U9368 ( .B1(n7940), .B2(n6864), .A(n7744), .ZN(n7745) );
  XNOR2_X1 U9369 ( .A(n7745), .B(n9030), .ZN(n7923) );
  XOR2_X1 U9370 ( .A(n7924), .B(n7923), .Z(n7927) );
  XOR2_X1 U9371 ( .A(n7928), .B(n7927), .Z(n7752) );
  NAND2_X1 U9372 ( .A1(P1_U3086), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n9333) );
  INV_X1 U9373 ( .A(n9333), .ZN(n7748) );
  OAI22_X1 U9374 ( .A1(n9174), .A2(n9241), .B1(n9255), .B2(n7746), .ZN(n7747)
         );
  AOI211_X1 U9375 ( .C1(n7767), .C2(n9257), .A(n7748), .B(n7747), .ZN(n7751)
         );
  NAND2_X1 U9376 ( .A1(n9252), .A2(n7749), .ZN(n7750) );
  OAI211_X1 U9377 ( .C1(n7752), .C2(n9259), .A(n7751), .B(n7750), .ZN(P1_U3213) );
  NAND2_X1 U9378 ( .A1(n7754), .A2(n7753), .ZN(n7756) );
  NAND2_X1 U9379 ( .A1(n7756), .A2(n7755), .ZN(n7757) );
  XNOR2_X1 U9380 ( .A(n7757), .B(n8433), .ZN(n7758) );
  OAI222_X1 U9381 ( .A1(n10076), .A2(n7838), .B1(n10074), .B2(n8311), .C1(
        n10080), .C2(n7758), .ZN(n7786) );
  INV_X1 U9382 ( .A(n7786), .ZN(n7766) );
  XNOR2_X1 U9383 ( .A(n7759), .B(n8433), .ZN(n7791) );
  INV_X1 U9384 ( .A(n7791), .ZN(n7764) );
  INV_X1 U9385 ( .A(n8930), .ZN(n7763) );
  INV_X1 U9386 ( .A(n7844), .ZN(n7761) );
  INV_X1 U9387 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n7760) );
  OAI22_X1 U9388 ( .A1(n7761), .A2(n8909), .B1(n10158), .B2(n7760), .ZN(n7762)
         );
  AOI21_X1 U9389 ( .B1(n7764), .B2(n7763), .A(n7762), .ZN(n7765) );
  OAI21_X1 U9390 ( .B1(n7766), .B2(n10156), .A(n7765), .ZN(P2_U3470) );
  INV_X1 U9391 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n7773) );
  AOI22_X1 U9392 ( .A1(n7768), .A2(n9573), .B1(n9959), .B2(n7767), .ZN(n7769)
         );
  OAI211_X1 U9393 ( .C1(n7771), .C2(n9914), .A(n7770), .B(n7769), .ZN(n7774)
         );
  NAND2_X1 U9394 ( .A1(n7774), .A2(n9968), .ZN(n7772) );
  OAI21_X1 U9395 ( .B1(n9968), .B2(n7773), .A(n7772), .ZN(P1_U3474) );
  NAND2_X1 U9396 ( .A1(n7774), .A2(n9983), .ZN(n7775) );
  OAI21_X1 U9397 ( .B1(n9983), .B2(n4547), .A(n7775), .ZN(P1_U3529) );
  AOI22_X1 U9398 ( .A1(n9266), .A2(n9879), .B1(n9880), .B2(n9878), .ZN(n7777)
         );
  OAI211_X1 U9399 ( .C1(n7778), .C2(n9962), .A(n7777), .B(n7776), .ZN(n7779)
         );
  AOI21_X1 U9400 ( .B1(n7780), .B2(n9964), .A(n7779), .ZN(n7783) );
  AOI22_X1 U9401 ( .A1(n8000), .A2(n9678), .B1(n9981), .B2(
        P1_REG1_REG_10__SCAN_IN), .ZN(n7781) );
  OAI21_X1 U9402 ( .B1(n7783), .B2(n9981), .A(n7781), .ZN(P1_U3532) );
  AOI22_X1 U9403 ( .A1(n8000), .A2(n9763), .B1(n9966), .B2(
        P1_REG0_REG_10__SCAN_IN), .ZN(n7782) );
  OAI21_X1 U9404 ( .B1(n7783), .B2(n9966), .A(n7782), .ZN(P1_U3483) );
  NAND2_X1 U9405 ( .A1(n7786), .A2(n10142), .ZN(n7785) );
  AOI22_X1 U9406 ( .A1(n7844), .A2(n9004), .B1(P2_REG0_REG_11__SCAN_IN), .B2(
        n10144), .ZN(n7784) );
  OAI211_X1 U9407 ( .C1(n7791), .C2(n9008), .A(n7785), .B(n7784), .ZN(P2_U3423) );
  NAND2_X1 U9408 ( .A1(n7786), .A2(n8867), .ZN(n7790) );
  INV_X1 U9409 ( .A(n7835), .ZN(n7787) );
  OAI22_X1 U9410 ( .A1(n8867), .A2(n7278), .B1(n7787), .B2(n8813), .ZN(n7788)
         );
  AOI21_X1 U9411 ( .B1(n7844), .B2(n10085), .A(n7788), .ZN(n7789) );
  OAI211_X1 U9412 ( .C1(n7791), .C2(n8872), .A(n7790), .B(n7789), .ZN(P2_U3222) );
  AOI211_X1 U9413 ( .C1(n7794), .C2(n9964), .A(n7793), .B(n7792), .ZN(n7799)
         );
  AOI22_X1 U9414 ( .A1(n9221), .A2(n9678), .B1(n9981), .B2(
        P1_REG1_REG_11__SCAN_IN), .ZN(n7795) );
  OAI21_X1 U9415 ( .B1(n7799), .B2(n9981), .A(n7795), .ZN(P1_U3533) );
  INV_X1 U9416 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n7796) );
  NOR2_X1 U9417 ( .A1(n9968), .A2(n7796), .ZN(n7797) );
  AOI21_X1 U9418 ( .B1(n9221), .B2(n9763), .A(n7797), .ZN(n7798) );
  OAI21_X1 U9419 ( .B1(n7799), .B2(n9966), .A(n7798), .ZN(P1_U3486) );
  INV_X1 U9420 ( .A(n8459), .ZN(n8250) );
  INV_X1 U9421 ( .A(n7800), .ZN(n7803) );
  OAI222_X1 U9422 ( .A1(n8250), .A2(P2_U3151), .B1(n9022), .B2(n7803), .C1(
        n7801), .C2(n9015), .ZN(P2_U3273) );
  OAI222_X1 U9423 ( .A1(n8071), .A2(n7804), .B1(n9797), .B2(n7803), .C1(n7802), 
        .C2(P1_U3086), .ZN(P1_U3333) );
  INV_X1 U9424 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n7808) );
  INV_X1 U9425 ( .A(n8312), .ZN(n7892) );
  OAI22_X1 U9426 ( .A1(n7805), .A2(n10120), .B1(n7892), .B2(n10118), .ZN(n7807) );
  NOR2_X1 U9427 ( .A1(n7807), .A2(n7806), .ZN(n7810) );
  MUX2_X1 U9428 ( .A(n7808), .B(n7810), .S(n10142), .Z(n7809) );
  INV_X1 U9429 ( .A(n7809), .ZN(P2_U3426) );
  MUX2_X1 U9430 ( .A(n7811), .B(n7810), .S(n10158), .Z(n7812) );
  INV_X1 U9431 ( .A(n7812), .ZN(P2_U3471) );
  INV_X1 U9432 ( .A(n7817), .ZN(n7815) );
  NAND2_X1 U9433 ( .A1(n9795), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n7813) );
  OAI211_X1 U9434 ( .C1(n7815), .C2(n9797), .A(n7814), .B(n7813), .ZN(P1_U3332) );
  NAND2_X1 U9435 ( .A1(n7817), .A2(n7816), .ZN(n7819) );
  NAND2_X1 U9436 ( .A1(n7818), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8462) );
  OAI211_X1 U9437 ( .C1(n7820), .C2(n9015), .A(n7819), .B(n8462), .ZN(P2_U3272) );
  OR2_X1 U9438 ( .A1(n8312), .A2(n8311), .ZN(n8314) );
  OR2_X1 U9439 ( .A1(n7822), .A2(n8611), .ZN(n7864) );
  NAND2_X1 U9440 ( .A1(n7822), .A2(n8611), .ZN(n7861) );
  NAND2_X1 U9441 ( .A1(n7864), .A2(n7861), .ZN(n8315) );
  XNOR2_X1 U9442 ( .A(n7847), .B(n8315), .ZN(n7896) );
  INV_X1 U9443 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n7828) );
  NAND2_X1 U9444 ( .A1(n7824), .A2(n7850), .ZN(n7825) );
  OR2_X1 U9445 ( .A1(n8312), .A2(n8612), .ZN(n7862) );
  NAND2_X1 U9446 ( .A1(n7825), .A2(n7862), .ZN(n7826) );
  INV_X1 U9447 ( .A(n8315), .ZN(n8434) );
  XNOR2_X1 U9448 ( .A(n7826), .B(n8434), .ZN(n7827) );
  AOI222_X1 U9449 ( .A1(n8843), .A2(n7827), .B1(n8612), .B2(n8838), .C1(n8610), 
        .C2(n8840), .ZN(n7893) );
  MUX2_X1 U9450 ( .A(n7828), .B(n7893), .S(n10142), .Z(n7830) );
  NAND2_X1 U9451 ( .A1(n7822), .A2(n9004), .ZN(n7829) );
  OAI211_X1 U9452 ( .C1(n7896), .C2(n9008), .A(n7830), .B(n7829), .ZN(P2_U3429) );
  INV_X1 U9453 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n7831) );
  MUX2_X1 U9454 ( .A(n7831), .B(n7893), .S(n10158), .Z(n7833) );
  NAND2_X1 U9455 ( .A1(n7822), .A2(n8927), .ZN(n7832) );
  OAI211_X1 U9456 ( .C1(n8930), .C2(n7896), .A(n7833), .B(n7832), .ZN(P2_U3472) );
  AOI21_X1 U9457 ( .B1(n8593), .B2(n8612), .A(n7834), .ZN(n7837) );
  NAND2_X1 U9458 ( .A1(n8598), .A2(n7835), .ZN(n7836) );
  OAI211_X1 U9459 ( .C1(n7838), .C2(n8595), .A(n7837), .B(n7836), .ZN(n7843)
         );
  AOI211_X1 U9460 ( .C1(n7841), .C2(n7840), .A(n8573), .B(n7839), .ZN(n7842)
         );
  AOI211_X1 U9461 ( .C1(n7844), .C2(n8585), .A(n7843), .B(n7842), .ZN(n7845)
         );
  INV_X1 U9462 ( .A(n7845), .ZN(P2_U3176) );
  AND2_X1 U9463 ( .A1(n7822), .A2(n8045), .ZN(n8319) );
  INV_X1 U9464 ( .A(n8319), .ZN(n7846) );
  NAND2_X1 U9465 ( .A1(n7847), .A2(n7846), .ZN(n7849) );
  NOR2_X1 U9466 ( .A1(n7822), .A2(n8045), .ZN(n8318) );
  INV_X1 U9467 ( .A(n8318), .ZN(n7848) );
  NAND2_X1 U9468 ( .A1(n7849), .A2(n7848), .ZN(n7951) );
  NAND2_X1 U9469 ( .A1(n8047), .A2(n8596), .ZN(n8328) );
  NAND2_X1 U9470 ( .A1(n8324), .A2(n8328), .ZN(n8321) );
  XNOR2_X1 U9471 ( .A(n7951), .B(n8437), .ZN(n7880) );
  INV_X1 U9472 ( .A(n8047), .ZN(n7870) );
  INV_X1 U9473 ( .A(n7851), .ZN(n7852) );
  INV_X1 U9474 ( .A(n7854), .ZN(n7856) );
  NOR2_X1 U9475 ( .A1(n7856), .A2(n7855), .ZN(n7857) );
  NAND2_X1 U9476 ( .A1(n7858), .A2(n7857), .ZN(n7859) );
  INV_X1 U9477 ( .A(n7861), .ZN(n7863) );
  OR2_X1 U9478 ( .A1(n7863), .A2(n7862), .ZN(n7865) );
  AOI21_X1 U9479 ( .B1(n7867), .B2(n8437), .A(n10080), .ZN(n7869) );
  OAI22_X1 U9480 ( .A1(n8045), .A2(n10076), .B1(n8863), .B2(n10074), .ZN(n7868) );
  AOI21_X1 U9481 ( .B1(n7869), .B2(n7954), .A(n7868), .ZN(n7876) );
  OAI21_X1 U9482 ( .B1(n7870), .B2(n8760), .A(n7876), .ZN(n7871) );
  NAND2_X1 U9483 ( .A1(n7871), .A2(n8867), .ZN(n7873) );
  AOI22_X1 U9484 ( .A1(n10092), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n10087), 
        .B2(n8042), .ZN(n7872) );
  OAI211_X1 U9485 ( .C1(n7880), .C2(n8872), .A(n7873), .B(n7872), .ZN(P2_U3219) );
  INV_X1 U9486 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n8625) );
  MUX2_X1 U9487 ( .A(n8625), .B(n7876), .S(n10158), .Z(n7875) );
  NAND2_X1 U9488 ( .A1(n8047), .A2(n8927), .ZN(n7874) );
  OAI211_X1 U9489 ( .C1(n7880), .C2(n8930), .A(n7875), .B(n7874), .ZN(P2_U3473) );
  INV_X1 U9490 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n7877) );
  MUX2_X1 U9491 ( .A(n7877), .B(n7876), .S(n10142), .Z(n7879) );
  NAND2_X1 U9492 ( .A1(n8047), .A2(n9004), .ZN(n7878) );
  OAI211_X1 U9493 ( .C1(n7880), .C2(n9008), .A(n7879), .B(n7878), .ZN(P2_U3432) );
  OAI21_X1 U9494 ( .B1(n7883), .B2(n7882), .A(n7881), .ZN(n7884) );
  NAND2_X1 U9495 ( .A1(n7884), .A2(n8589), .ZN(n7891) );
  NAND2_X1 U9496 ( .A1(n8593), .A2(n8611), .ZN(n7886) );
  OAI211_X1 U9497 ( .C1(n7887), .C2(n8595), .A(n7886), .B(n7885), .ZN(n7888)
         );
  AOI21_X1 U9498 ( .B1(n7889), .B2(n8598), .A(n7888), .ZN(n7890) );
  OAI211_X1 U9499 ( .C1(n7892), .C2(n8602), .A(n7891), .B(n7890), .ZN(P2_U3164) );
  INV_X1 U9500 ( .A(n7822), .ZN(n7972) );
  NOR2_X1 U9501 ( .A1(n7972), .A2(n8760), .ZN(n7895) );
  INV_X1 U9502 ( .A(n7893), .ZN(n7894) );
  AOI211_X1 U9503 ( .C1(n10087), .C2(n7969), .A(n7895), .B(n7894), .ZN(n7899)
         );
  INV_X1 U9504 ( .A(n7896), .ZN(n7897) );
  AOI22_X1 U9505 ( .A1(n7897), .A2(n8819), .B1(P2_REG2_REG_13__SCAN_IN), .B2(
        n10092), .ZN(n7898) );
  OAI21_X1 U9506 ( .B1(n7899), .B2(n10092), .A(n7898), .ZN(P2_U3220) );
  INV_X1 U9507 ( .A(n7900), .ZN(n7949) );
  OAI222_X1 U9508 ( .A1(n9797), .A2(n7949), .B1(P1_U3086), .B2(n7902), .C1(
        n7901), .C2(n8071), .ZN(P1_U3331) );
  INV_X1 U9509 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n7903) );
  MUX2_X1 U9510 ( .A(n7903), .B(P1_REG1_REG_13__SCAN_IN), .S(n9833), .Z(n9826)
         );
  OAI21_X1 U9511 ( .B1(P1_REG1_REG_12__SCAN_IN), .B2(n7910), .A(n7904), .ZN(
        n9827) );
  NOR2_X1 U9512 ( .A1(n9826), .A2(n9827), .ZN(n9825) );
  XNOR2_X1 U9513 ( .A(n9837), .B(P1_REG1_REG_14__SCAN_IN), .ZN(n9845) );
  NOR2_X1 U9514 ( .A1(n7905), .A2(n9856), .ZN(n7906) );
  INV_X1 U9515 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n9859) );
  NOR2_X1 U9516 ( .A1(n9859), .A2(n9860), .ZN(n9858) );
  NOR2_X1 U9517 ( .A1(n7906), .A2(n9858), .ZN(n8050) );
  XNOR2_X1 U9518 ( .A(n8054), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n8051) );
  XNOR2_X1 U9519 ( .A(n8050), .B(n8051), .ZN(n7922) );
  INV_X1 U9520 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n7907) );
  NAND2_X1 U9521 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9153) );
  OAI21_X1 U9522 ( .B1(n9872), .B2(n7907), .A(n9153), .ZN(n7920) );
  NAND2_X1 U9523 ( .A1(P1_REG2_REG_13__SCAN_IN), .A2(n9833), .ZN(n7908) );
  OAI21_X1 U9524 ( .B1(P1_REG2_REG_13__SCAN_IN), .B2(n9833), .A(n7908), .ZN(
        n9829) );
  OAI21_X1 U9525 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(n7910), .A(n7909), .ZN(
        n9830) );
  NOR2_X1 U9526 ( .A1(n9829), .A2(n9830), .ZN(n9828) );
  AOI21_X1 U9527 ( .B1(n9833), .B2(P1_REG2_REG_13__SCAN_IN), .A(n9828), .ZN(
        n9839) );
  NAND2_X1 U9528 ( .A1(P1_REG2_REG_14__SCAN_IN), .A2(n9837), .ZN(n7911) );
  OAI21_X1 U9529 ( .B1(P1_REG2_REG_14__SCAN_IN), .B2(n9837), .A(n7911), .ZN(
        n9840) );
  NOR2_X1 U9530 ( .A1(n9839), .A2(n9840), .ZN(n9838) );
  AOI21_X1 U9531 ( .B1(n9837), .B2(P1_REG2_REG_14__SCAN_IN), .A(n9838), .ZN(
        n7912) );
  NOR2_X1 U9532 ( .A1(n7912), .A2(n9856), .ZN(n7913) );
  INV_X1 U9533 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n9863) );
  XNOR2_X1 U9534 ( .A(n9856), .B(n7912), .ZN(n9864) );
  NOR2_X1 U9535 ( .A1(n9863), .A2(n9864), .ZN(n9862) );
  NOR2_X1 U9536 ( .A1(n7913), .A2(n9862), .ZN(n7918) );
  INV_X1 U9537 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n7914) );
  XNOR2_X1 U9538 ( .A(n7915), .B(n7914), .ZN(n7917) );
  OR2_X1 U9539 ( .A1(n7918), .A2(n7917), .ZN(n8056) );
  INV_X1 U9540 ( .A(n8056), .ZN(n7916) );
  AOI211_X1 U9541 ( .C1(n7918), .C2(n7917), .A(n9861), .B(n7916), .ZN(n7919)
         );
  AOI211_X1 U9542 ( .C1(n9868), .C2(n8054), .A(n7920), .B(n7919), .ZN(n7921)
         );
  OAI21_X1 U9543 ( .B1(n7922), .B2(n9857), .A(n7921), .ZN(P1_U3259) );
  INV_X1 U9544 ( .A(n7923), .ZN(n7926) );
  INV_X1 U9545 ( .A(n7924), .ZN(n7925) );
  NAND2_X1 U9546 ( .A1(n7938), .A2(n9044), .ZN(n7930) );
  OR2_X1 U9547 ( .A1(n9174), .A2(n6864), .ZN(n7929) );
  NAND2_X1 U9548 ( .A1(n7930), .A2(n7929), .ZN(n7931) );
  XNOR2_X1 U9549 ( .A(n7931), .B(n9030), .ZN(n9168) );
  XOR2_X1 U9550 ( .A(n9169), .B(n9168), .Z(n7935) );
  NAND2_X1 U9551 ( .A1(n7938), .A2(n9049), .ZN(n7933) );
  OR2_X1 U9552 ( .A1(n9174), .A2(n9113), .ZN(n7932) );
  NAND2_X1 U9553 ( .A1(n7933), .A2(n7932), .ZN(n7987) );
  INV_X1 U9554 ( .A(n7987), .ZN(n7934) );
  NAND2_X1 U9555 ( .A1(n7935), .A2(n7934), .ZN(n9167) );
  OAI21_X1 U9556 ( .B1(n7935), .B2(n7934), .A(n9167), .ZN(n7946) );
  INV_X1 U9557 ( .A(n7936), .ZN(n7937) );
  AOI21_X1 U9558 ( .B1(n9251), .B2(n9266), .A(n7937), .ZN(n7944) );
  NAND2_X1 U9559 ( .A1(n9257), .A2(n7938), .ZN(n7943) );
  NAND2_X1 U9560 ( .A1(n9252), .A2(n7939), .ZN(n7942) );
  OR2_X1 U9561 ( .A1(n9255), .A2(n7940), .ZN(n7941) );
  NAND4_X1 U9562 ( .A1(n7944), .A2(n7943), .A3(n7942), .A4(n7941), .ZN(n7945)
         );
  AOI21_X1 U9563 ( .B1(n7946), .B2(n9237), .A(n7945), .ZN(n7947) );
  INV_X1 U9564 ( .A(n7947), .ZN(P1_U3221) );
  OAI222_X1 U9565 ( .A1(n7950), .A2(P2_U3151), .B1(n9022), .B2(n7949), .C1(
        n7948), .C2(n9015), .ZN(P2_U3271) );
  NAND2_X1 U9566 ( .A1(n7951), .A2(n8328), .ZN(n7952) );
  NAND2_X1 U9567 ( .A1(n7952), .A2(n8324), .ZN(n8213) );
  NAND2_X1 U9568 ( .A1(n8588), .A2(n8863), .ZN(n8326) );
  AND2_X2 U9569 ( .A1(n8331), .A2(n8326), .ZN(n8436) );
  XNOR2_X1 U9570 ( .A(n8213), .B(n8436), .ZN(n7981) );
  NAND2_X1 U9571 ( .A1(n8047), .A2(n8610), .ZN(n7953) );
  NAND2_X1 U9572 ( .A1(n7954), .A2(n7953), .ZN(n7956) );
  INV_X1 U9573 ( .A(n8436), .ZN(n7955) );
  OAI21_X1 U9574 ( .B1(n7956), .B2(n7955), .A(n8843), .ZN(n7957) );
  AOI22_X1 U9575 ( .A1(n8610), .A2(n8838), .B1(n8840), .B2(n8608), .ZN(n7958)
         );
  NAND2_X1 U9576 ( .A1(n7959), .A2(n7958), .ZN(n7973) );
  MUX2_X1 U9577 ( .A(n7973), .B(P2_REG2_REG_15__SCAN_IN), .S(n10092), .Z(n7960) );
  INV_X1 U9578 ( .A(n7960), .ZN(n7962) );
  AOI22_X1 U9579 ( .A1(n8588), .A2(n10085), .B1(n10087), .B2(n8599), .ZN(n7961) );
  OAI211_X1 U9580 ( .C1(n7981), .C2(n8872), .A(n7962), .B(n7961), .ZN(P2_U3218) );
  OAI21_X1 U9581 ( .B1(n7965), .B2(n7964), .A(n7963), .ZN(n7966) );
  NAND2_X1 U9582 ( .A1(n7966), .A2(n8589), .ZN(n7971) );
  AOI22_X1 U9583 ( .A1(n8593), .A2(n8610), .B1(P2_REG3_REG_13__SCAN_IN), .B2(
        P2_U3151), .ZN(n7967) );
  OAI21_X1 U9584 ( .B1(n8311), .B2(n8595), .A(n7967), .ZN(n7968) );
  AOI21_X1 U9585 ( .B1(n7969), .B2(n8598), .A(n7968), .ZN(n7970) );
  OAI211_X1 U9586 ( .C1(n7972), .C2(n8602), .A(n7971), .B(n7970), .ZN(P2_U3174) );
  INV_X1 U9587 ( .A(n7973), .ZN(n7978) );
  INV_X1 U9588 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n7974) );
  MUX2_X1 U9589 ( .A(n7978), .B(n7974), .S(n10156), .Z(n7976) );
  NAND2_X1 U9590 ( .A1(n8588), .A2(n8927), .ZN(n7975) );
  OAI211_X1 U9591 ( .C1(n7981), .C2(n8930), .A(n7976), .B(n7975), .ZN(P2_U3474) );
  INV_X1 U9592 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n7977) );
  MUX2_X1 U9593 ( .A(n7978), .B(n7977), .S(n10144), .Z(n7980) );
  NAND2_X1 U9594 ( .A1(n8588), .A2(n9004), .ZN(n7979) );
  OAI211_X1 U9595 ( .C1(n7981), .C2(n9008), .A(n7980), .B(n7979), .ZN(P2_U3435) );
  AOI22_X1 U9596 ( .A1(n7984), .A2(n9044), .B1(n9049), .B2(n9266), .ZN(n7982)
         );
  XNOR2_X1 U9597 ( .A(n7982), .B(n9030), .ZN(n9171) );
  NOR2_X1 U9598 ( .A1(n9092), .A2(n9113), .ZN(n7983) );
  AOI21_X1 U9599 ( .B1(n7984), .B2(n9049), .A(n7983), .ZN(n9170) );
  NAND2_X1 U9600 ( .A1(n9171), .A2(n9170), .ZN(n7986) );
  OR2_X1 U9601 ( .A1(n9168), .A2(n7987), .ZN(n7985) );
  AND2_X1 U9602 ( .A1(n9168), .A2(n7987), .ZN(n7990) );
  INV_X1 U9603 ( .A(n9170), .ZN(n7989) );
  INV_X1 U9604 ( .A(n9171), .ZN(n7988) );
  OAI21_X1 U9605 ( .B1(n7990), .B2(n7989), .A(n7988), .ZN(n7992) );
  INV_X1 U9606 ( .A(n7990), .ZN(n7991) );
  AOI22_X1 U9607 ( .A1(n9221), .A2(n9044), .B1(n9049), .B2(n9878), .ZN(n7993)
         );
  XOR2_X1 U9608 ( .A(n9030), .B(n7993), .Z(n9213) );
  INV_X1 U9609 ( .A(n9213), .ZN(n8001) );
  NAND2_X1 U9610 ( .A1(n9221), .A2(n9049), .ZN(n7995) );
  NAND2_X1 U9611 ( .A1(n9878), .A2(n9033), .ZN(n7994) );
  NAND2_X1 U9612 ( .A1(n7995), .A2(n7994), .ZN(n9212) );
  INV_X1 U9613 ( .A(n9212), .ZN(n8004) );
  NAND2_X1 U9614 ( .A1(n8000), .A2(n9044), .ZN(n7997) );
  NAND2_X1 U9615 ( .A1(n9265), .A2(n9049), .ZN(n7996) );
  NAND2_X1 U9616 ( .A1(n7997), .A2(n7996), .ZN(n7998) );
  XNOR2_X1 U9617 ( .A(n7998), .B(n9111), .ZN(n9209) );
  NOR2_X1 U9618 ( .A1(n9219), .A2(n9113), .ZN(n7999) );
  AOI21_X1 U9619 ( .B1(n8000), .B2(n9049), .A(n7999), .ZN(n9088) );
  OAI22_X1 U9620 ( .A1(n8001), .A2(n8004), .B1(n9209), .B2(n9088), .ZN(n8007)
         );
  NAND2_X1 U9621 ( .A1(n9209), .A2(n9088), .ZN(n8002) );
  INV_X1 U9622 ( .A(n8002), .ZN(n8005) );
  AOI21_X1 U9623 ( .B1(n9212), .B2(n8002), .A(n9213), .ZN(n8003) );
  AOI21_X1 U9624 ( .B1(n8005), .B2(n8004), .A(n8003), .ZN(n8006) );
  NAND2_X1 U9625 ( .A1(n9890), .A2(n9044), .ZN(n8009) );
  OR2_X1 U9626 ( .A1(n9953), .A2(n6864), .ZN(n8008) );
  NAND2_X1 U9627 ( .A1(n8009), .A2(n8008), .ZN(n8010) );
  XNOR2_X1 U9628 ( .A(n8010), .B(n9030), .ZN(n8113) );
  AOI22_X1 U9629 ( .A1(n9890), .A2(n9049), .B1(n9033), .B2(n9264), .ZN(n8114)
         );
  XNOR2_X1 U9630 ( .A(n8113), .B(n8114), .ZN(n8116) );
  XOR2_X1 U9631 ( .A(n8117), .B(n8116), .Z(n8016) );
  NAND2_X1 U9632 ( .A1(n9251), .A2(n9881), .ZN(n8012) );
  OAI211_X1 U9633 ( .C1(n9094), .C2(n9255), .A(n8012), .B(n8011), .ZN(n8014)
         );
  INV_X1 U9634 ( .A(n9890), .ZN(n9948) );
  NOR2_X1 U9635 ( .A1(n9948), .A2(n9247), .ZN(n8013) );
  AOI211_X1 U9636 ( .C1(n9884), .C2(n9252), .A(n8014), .B(n8013), .ZN(n8015)
         );
  OAI21_X1 U9637 ( .B1(n8016), .B2(n9259), .A(n8015), .ZN(P1_U3224) );
  INV_X1 U9638 ( .A(n8017), .ZN(n8018) );
  NOR2_X1 U9639 ( .A1(n8026), .A2(n8018), .ZN(n8021) );
  INV_X1 U9640 ( .A(n9615), .ZN(n8019) );
  AOI21_X1 U9641 ( .B1(n8021), .B2(n8020), .A(n8019), .ZN(n9961) );
  NAND2_X1 U9642 ( .A1(n9221), .A2(n9878), .ZN(n8023) );
  NOR2_X1 U9643 ( .A1(n9221), .A2(n9878), .ZN(n8022) );
  AOI21_X1 U9644 ( .B1(n8027), .B2(n8026), .A(n8086), .ZN(n9965) );
  NAND2_X1 U9645 ( .A1(n9965), .A2(n9907), .ZN(n8034) );
  AOI211_X1 U9646 ( .C1(n9958), .C2(n9892), .A(n9889), .B(n9624), .ZN(n9956)
         );
  INV_X1 U9647 ( .A(n9958), .ZN(n8031) );
  AOI22_X1 U9648 ( .A1(n4315), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n9194), .B2(
        n9898), .ZN(n8028) );
  OAI21_X1 U9649 ( .B1(n9587), .B2(n9953), .A(n8028), .ZN(n8029) );
  AOI21_X1 U9650 ( .B1(n9568), .B2(n9601), .A(n8029), .ZN(n8030) );
  OAI21_X1 U9651 ( .B1(n8031), .B2(n9630), .A(n8030), .ZN(n8032) );
  AOI21_X1 U9652 ( .B1(n9956), .B2(n9635), .A(n8032), .ZN(n8033) );
  OAI211_X1 U9653 ( .C1(n9961), .C2(n9579), .A(n8034), .B(n8033), .ZN(P1_U3280) );
  INV_X1 U9654 ( .A(n8035), .ZN(n8038) );
  OAI222_X1 U9655 ( .A1(n9797), .A2(n8038), .B1(P1_U3086), .B2(n6336), .C1(
        n8036), .C2(n8071), .ZN(P1_U3330) );
  OAI222_X1 U9656 ( .A1(n8039), .A2(P2_U3151), .B1(n9022), .B2(n8038), .C1(
        n8037), .C2(n9015), .ZN(P2_U3270) );
  XOR2_X1 U9657 ( .A(n8041), .B(n8040), .Z(n8049) );
  INV_X1 U9658 ( .A(n8863), .ZN(n8609) );
  AOI22_X1 U9659 ( .A1(n8593), .A2(n8609), .B1(P2_REG3_REG_14__SCAN_IN), .B2(
        P2_U3151), .ZN(n8044) );
  NAND2_X1 U9660 ( .A1(n8598), .A2(n8042), .ZN(n8043) );
  OAI211_X1 U9661 ( .C1(n8045), .C2(n8595), .A(n8044), .B(n8043), .ZN(n8046)
         );
  AOI21_X1 U9662 ( .B1(n8047), .B2(n8585), .A(n8046), .ZN(n8048) );
  OAI21_X1 U9663 ( .B1(n8049), .B2(n8573), .A(n8048), .ZN(P2_U3155) );
  INV_X1 U9664 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9734) );
  XNOR2_X1 U9665 ( .A(n9349), .B(n9734), .ZN(n9344) );
  INV_X1 U9666 ( .A(n8050), .ZN(n8052) );
  OAI22_X1 U9667 ( .A1(n8052), .A2(n8051), .B1(n8054), .B2(
        P1_REG1_REG_16__SCAN_IN), .ZN(n9345) );
  XOR2_X1 U9668 ( .A(n9344), .B(n9345), .Z(n8064) );
  INV_X1 U9669 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n8053) );
  XNOR2_X1 U9670 ( .A(n9349), .B(n8053), .ZN(n8058) );
  NAND2_X1 U9671 ( .A1(n8054), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n8055) );
  AND2_X1 U9672 ( .A1(n8056), .A2(n8055), .ZN(n8057) );
  NAND2_X1 U9673 ( .A1(n8057), .A2(n8058), .ZN(n9351) );
  OAI21_X1 U9674 ( .B1(n8058), .B2(n8057), .A(n9351), .ZN(n8062) );
  NOR2_X1 U9675 ( .A1(n8059), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9162) );
  AOI21_X1 U9676 ( .B1(n9375), .B2(P1_ADDR_REG_17__SCAN_IN), .A(n9162), .ZN(
        n8060) );
  OAI21_X1 U9677 ( .B1(n9343), .B2(n9851), .A(n8060), .ZN(n8061) );
  AOI21_X1 U9678 ( .B1(n8062), .B2(n9842), .A(n8061), .ZN(n8063) );
  OAI21_X1 U9679 ( .B1(n8064), .B2(n9857), .A(n8063), .ZN(P1_U3260) );
  INV_X1 U9680 ( .A(n8065), .ZN(n8068) );
  OAI222_X1 U9681 ( .A1(n8067), .A2(P2_U3151), .B1(n9022), .B2(n8068), .C1(
        n8066), .C2(n9015), .ZN(P2_U3269) );
  OAI222_X1 U9682 ( .A1(n8071), .A2(n8070), .B1(P1_U3086), .B2(n8069), .C1(
        n9797), .C2(n8068), .ZN(P1_U3329) );
  INV_X1 U9683 ( .A(n8072), .ZN(n8085) );
  AOI21_X1 U9684 ( .B1(n9020), .B2(P1_DATAO_REG_27__SCAN_IN), .A(n8073), .ZN(
        n8074) );
  OAI21_X1 U9685 ( .B1(n8085), .B2(n9022), .A(n8074), .ZN(P2_U3268) );
  INV_X1 U9686 ( .A(n8207), .ZN(n9017) );
  OAI222_X1 U9687 ( .A1(n9797), .A2(n9017), .B1(n8076), .B2(P1_U3086), .C1(
        n8075), .C2(n8071), .ZN(P1_U3326) );
  OAI222_X1 U9688 ( .A1(n9015), .A2(n4776), .B1(n9022), .B2(n8078), .C1(
        P2_U3151), .C2(n4316), .ZN(P2_U3293) );
  NAND2_X1 U9689 ( .A1(n8079), .A2(n9983), .ZN(n8081) );
  NAND2_X1 U9690 ( .A1(n9981), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n8080) );
  OAI211_X1 U9691 ( .C1(n8082), .C2(n9747), .A(n8081), .B(n8080), .ZN(P1_U3523) );
  OAI222_X1 U9692 ( .A1(n9797), .A2(n8085), .B1(n8084), .B2(P1_U3086), .C1(
        n8083), .C2(n8071), .ZN(P1_U3328) );
  INV_X1 U9693 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n8108) );
  NOR2_X1 U9694 ( .A1(n9749), .A2(n9601), .ZN(n8087) );
  NAND2_X1 U9695 ( .A1(n9582), .A2(n9581), .ZN(n9580) );
  NAND2_X1 U9696 ( .A1(n9783), .A2(n9556), .ZN(n8090) );
  INV_X1 U9697 ( .A(n9705), .ZN(n9525) );
  NOR2_X1 U9698 ( .A1(n9684), .A2(n9690), .ZN(n8095) );
  NAND2_X1 U9699 ( .A1(n9684), .A2(n9690), .ZN(n8094) );
  XNOR2_X1 U9700 ( .A(n9395), .B(n8105), .ZN(n9468) );
  AOI211_X1 U9701 ( .C1(n8096), .C2(n9481), .A(n9889), .B(n9457), .ZN(n9469)
         );
  NAND2_X1 U9702 ( .A1(n9493), .A2(n8100), .ZN(n8102) );
  OAI211_X1 U9703 ( .C1(n8105), .C2(n8104), .A(n9386), .B(n9876), .ZN(n8107)
         );
  AOI22_X1 U9704 ( .A1(n9665), .A2(n9880), .B1(n9879), .B2(n9690), .ZN(n8106)
         );
  NAND2_X1 U9705 ( .A1(n8107), .A2(n8106), .ZN(n9475) );
  AOI211_X1 U9706 ( .C1(n9468), .C2(n9964), .A(n9469), .B(n9475), .ZN(n8110)
         );
  MUX2_X1 U9707 ( .A(n8108), .B(n8110), .S(n9968), .Z(n8109) );
  OAI21_X1 U9708 ( .B1(n9473), .B2(n9788), .A(n8109), .ZN(P1_U3514) );
  INV_X1 U9709 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n8111) );
  MUX2_X1 U9710 ( .A(n8111), .B(n8110), .S(n9983), .Z(n8112) );
  OAI21_X1 U9711 ( .B1(n9473), .B2(n9747), .A(n8112), .ZN(P1_U3546) );
  INV_X1 U9712 ( .A(n8113), .ZN(n8115) );
  AOI22_X1 U9713 ( .A1(n9958), .A2(n9049), .B1(n9033), .B2(n9881), .ZN(n8121)
         );
  NAND2_X1 U9714 ( .A1(n9958), .A2(n9044), .ZN(n8119) );
  OR2_X1 U9715 ( .A1(n9617), .A2(n6864), .ZN(n8118) );
  NAND2_X1 U9716 ( .A1(n8119), .A2(n8118), .ZN(n8120) );
  XNOR2_X1 U9717 ( .A(n8120), .B(n9030), .ZN(n8123) );
  XOR2_X1 U9718 ( .A(n8121), .B(n8123), .Z(n9192) );
  INV_X1 U9719 ( .A(n8121), .ZN(n8122) );
  AOI22_X1 U9720 ( .A1(n9749), .A2(n9044), .B1(n9049), .B2(n9601), .ZN(n8124)
         );
  XNOR2_X1 U9721 ( .A(n8124), .B(n9030), .ZN(n9067) );
  AOI22_X1 U9722 ( .A1(n9749), .A2(n9049), .B1(n9033), .B2(n9601), .ZN(n9066)
         );
  NAND2_X1 U9723 ( .A1(n9069), .A2(n9067), .ZN(n8125) );
  NAND2_X1 U9724 ( .A1(n8126), .A2(n8125), .ZN(n9147) );
  NAND2_X1 U9725 ( .A1(n9583), .A2(n9044), .ZN(n8128) );
  OR2_X1 U9726 ( .A1(n9571), .A2(n6864), .ZN(n8127) );
  NAND2_X1 U9727 ( .A1(n8128), .A2(n8127), .ZN(n8129) );
  XNOR2_X1 U9728 ( .A(n8129), .B(n9030), .ZN(n9150) );
  NOR2_X1 U9729 ( .A1(n9571), .A2(n9113), .ZN(n8130) );
  AOI21_X1 U9730 ( .B1(n9583), .B2(n9049), .A(n8130), .ZN(n9149) );
  INV_X1 U9731 ( .A(n9149), .ZN(n8140) );
  NAND2_X1 U9732 ( .A1(n9606), .A2(n9049), .ZN(n8132) );
  NAND2_X1 U9733 ( .A1(n9263), .A2(n9033), .ZN(n8131) );
  AND2_X1 U9734 ( .A1(n8132), .A2(n8131), .ZN(n8137) );
  INV_X1 U9735 ( .A(n8137), .ZN(n9249) );
  NAND2_X1 U9736 ( .A1(n9606), .A2(n9044), .ZN(n8134) );
  NAND2_X1 U9737 ( .A1(n9263), .A2(n9049), .ZN(n8133) );
  NAND2_X1 U9738 ( .A1(n8134), .A2(n8133), .ZN(n8135) );
  XNOR2_X1 U9739 ( .A(n8135), .B(n9111), .ZN(n9148) );
  INV_X1 U9740 ( .A(n9148), .ZN(n8136) );
  AOI22_X1 U9741 ( .A1(n9150), .A2(n8140), .B1(n9249), .B2(n8136), .ZN(n8143)
         );
  AND2_X1 U9742 ( .A1(n9148), .A2(n8137), .ZN(n8138) );
  NOR2_X1 U9743 ( .A1(n8138), .A2(n9149), .ZN(n8141) );
  INV_X1 U9744 ( .A(n8138), .ZN(n8139) );
  OAI22_X1 U9745 ( .A1(n8141), .A2(n9150), .B1(n8140), .B2(n8139), .ZN(n8142)
         );
  AOI22_X1 U9746 ( .A1(n4605), .A2(n9044), .B1(n9049), .B2(n9719), .ZN(n8144)
         );
  XNOR2_X1 U9747 ( .A(n8144), .B(n9030), .ZN(n8145) );
  OAI22_X1 U9748 ( .A1(n9783), .A2(n6864), .B1(n9556), .B2(n9113), .ZN(n8146)
         );
  XNOR2_X1 U9749 ( .A(n8145), .B(n8146), .ZN(n9160) );
  INV_X1 U9750 ( .A(n8145), .ZN(n8147) );
  NAND2_X1 U9751 ( .A1(n8147), .A2(n8146), .ZN(n8148) );
  AOI22_X1 U9752 ( .A1(n9560), .A2(n9044), .B1(n9049), .B2(n9727), .ZN(n8149)
         );
  XOR2_X1 U9753 ( .A(n9030), .B(n8149), .Z(n8150) );
  AOI22_X1 U9754 ( .A1(n9560), .A2(n9049), .B1(n9033), .B2(n9727), .ZN(n9226)
         );
  NAND2_X1 U9755 ( .A1(n9224), .A2(n9226), .ZN(n8152) );
  INV_X1 U9756 ( .A(n8150), .ZN(n8151) );
  AOI22_X1 U9757 ( .A1(n9541), .A2(n9044), .B1(n9049), .B2(n9718), .ZN(n8153)
         );
  XOR2_X1 U9758 ( .A(n9030), .B(n8153), .Z(n9102) );
  OAI22_X1 U9759 ( .A1(n9775), .A2(n6864), .B1(n9530), .B2(n9113), .ZN(n9101)
         );
  NOR2_X1 U9760 ( .A1(n9102), .A2(n9101), .ZN(n8155) );
  NAND2_X1 U9761 ( .A1(n9102), .A2(n9101), .ZN(n8154) );
  OAI22_X1 U9762 ( .A1(n9525), .A2(n4406), .B1(n9709), .B2(n6864), .ZN(n8156)
         );
  XOR2_X1 U9763 ( .A(n9030), .B(n8156), .Z(n8158) );
  INV_X1 U9764 ( .A(n9709), .ZN(n9545) );
  AOI22_X1 U9765 ( .A1(n9705), .A2(n9049), .B1(n9033), .B2(n9545), .ZN(n8157)
         );
  NAND2_X1 U9766 ( .A1(n8158), .A2(n8157), .ZN(n9128) );
  OAI21_X1 U9767 ( .B1(n8158), .B2(n8157), .A(n9128), .ZN(n9185) );
  OAI22_X1 U9768 ( .A1(n9770), .A2(n6864), .B1(n9531), .B2(n9113), .ZN(n8161)
         );
  OAI22_X1 U9769 ( .A1(n9770), .A2(n4406), .B1(n9531), .B2(n6864), .ZN(n8159)
         );
  XNOR2_X1 U9770 ( .A(n8159), .B(n9030), .ZN(n8162) );
  XOR2_X1 U9771 ( .A(n8161), .B(n8162), .Z(n9131) );
  INV_X1 U9772 ( .A(n9131), .ZN(n8160) );
  OAI22_X1 U9773 ( .A1(n9693), .A2(n4406), .B1(n9680), .B2(n6864), .ZN(n8163)
         );
  XOR2_X1 U9774 ( .A(n9030), .B(n8163), .Z(n8164) );
  NAND2_X2 U9775 ( .A1(n8165), .A2(n8164), .ZN(n9076) );
  OAI22_X1 U9776 ( .A1(n9693), .A2(n6864), .B1(n9680), .B2(n9113), .ZN(n9201)
         );
  NAND2_X1 U9777 ( .A1(n9684), .A2(n9044), .ZN(n8167) );
  NAND2_X1 U9778 ( .A1(n9690), .A2(n9049), .ZN(n8166) );
  NAND2_X1 U9779 ( .A1(n8167), .A2(n8166), .ZN(n8168) );
  XNOR2_X1 U9780 ( .A(n8168), .B(n9111), .ZN(n8170) );
  AND2_X1 U9781 ( .A1(n9690), .A2(n9033), .ZN(n8169) );
  AOI21_X1 U9782 ( .B1(n9684), .B2(n9049), .A(n8169), .ZN(n8171) );
  NAND2_X1 U9783 ( .A1(n8170), .A2(n8171), .ZN(n8184) );
  INV_X1 U9784 ( .A(n8170), .ZN(n8173) );
  INV_X1 U9785 ( .A(n8171), .ZN(n8172) );
  NAND2_X1 U9786 ( .A1(n8173), .A2(n8172), .ZN(n8174) );
  INV_X1 U9787 ( .A(n8185), .ZN(n9079) );
  INV_X1 U9788 ( .A(n8184), .ZN(n8183) );
  OAI22_X1 U9789 ( .A1(n9473), .A2(n4406), .B1(n9681), .B2(n6864), .ZN(n8175)
         );
  XNOR2_X1 U9790 ( .A(n8175), .B(n9111), .ZN(n8178) );
  OR2_X1 U9791 ( .A1(n9473), .A2(n6864), .ZN(n8177) );
  NAND2_X1 U9792 ( .A1(n9486), .A2(n9033), .ZN(n8176) );
  NAND2_X1 U9793 ( .A1(n8178), .A2(n8179), .ZN(n9026) );
  INV_X1 U9794 ( .A(n8178), .ZN(n8181) );
  INV_X1 U9795 ( .A(n8179), .ZN(n8180) );
  NAND2_X1 U9796 ( .A1(n8181), .A2(n8180), .ZN(n8182) );
  NOR3_X1 U9797 ( .A1(n9079), .A2(n8183), .A3(n8186), .ZN(n8189) );
  INV_X1 U9799 ( .A(n9027), .ZN(n8188) );
  OAI21_X1 U9800 ( .B1(n8189), .B2(n8188), .A(n9237), .ZN(n8194) );
  AOI22_X1 U9801 ( .A1(n9665), .A2(n9251), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3086), .ZN(n8190) );
  OAI21_X1 U9802 ( .B1(n8191), .B2(n9255), .A(n8190), .ZN(n8192) );
  AOI21_X1 U9803 ( .B1(n9470), .B2(n9252), .A(n8192), .ZN(n8193) );
  OAI211_X1 U9804 ( .C1(n9473), .C2(n9247), .A(n8194), .B(n8193), .ZN(P1_U3229) );
  NAND2_X1 U9805 ( .A1(n9005), .A2(n8853), .ZN(n8325) );
  NAND2_X1 U9806 ( .A1(n8330), .A2(n8325), .ZN(n8440) );
  NAND2_X1 U9807 ( .A1(n8998), .A2(n8864), .ZN(n8337) );
  NAND2_X1 U9808 ( .A1(n8333), .A2(n8337), .ZN(n8441) );
  NOR2_X1 U9809 ( .A1(n8992), .A2(n8825), .ZN(n8197) );
  INV_X1 U9810 ( .A(n8992), .ZN(n8196) );
  OAI22_X1 U9811 ( .A1(n8837), .A2(n8197), .B1(n8852), .B2(n8196), .ZN(n8824)
         );
  NAND2_X1 U9812 ( .A1(n8986), .A2(n8570), .ZN(n8347) );
  INV_X1 U9813 ( .A(n8823), .ZN(n8198) );
  INV_X1 U9814 ( .A(n8570), .ZN(n8841) );
  AOI22_X1 U9815 ( .A1(n8824), .A2(n8198), .B1(n8986), .B2(n8841), .ZN(n8809)
         );
  NAND2_X1 U9816 ( .A1(n8913), .A2(n8802), .ZN(n8794) );
  NOR2_X1 U9817 ( .A1(n8913), .A2(n8826), .ZN(n8798) );
  NAND2_X1 U9818 ( .A1(n8979), .A2(n8560), .ZN(n8344) );
  NAND2_X1 U9819 ( .A1(n8973), .A2(n8801), .ZN(n8244) );
  INV_X1 U9820 ( .A(n8783), .ZN(n8786) );
  NAND2_X1 U9821 ( .A1(n8489), .A2(n8788), .ZN(n8200) );
  NAND2_X1 U9822 ( .A1(n8962), .A2(n8774), .ZN(n8357) );
  NAND2_X1 U9823 ( .A1(n8360), .A2(n8357), .ZN(n8769) );
  NAND2_X1 U9824 ( .A1(n8762), .A2(n8769), .ZN(n8761) );
  NAND2_X1 U9825 ( .A1(n8761), .A2(n4943), .ZN(n8752) );
  NOR2_X1 U9826 ( .A1(n8201), .A2(n8765), .ZN(n8364) );
  INV_X1 U9827 ( .A(n8364), .ZN(n8202) );
  INV_X1 U9828 ( .A(n8950), .ZN(n8203) );
  NAND2_X1 U9829 ( .A1(n8203), .A2(n8576), .ZN(n8204) );
  NOR2_X1 U9830 ( .A1(n8887), .A2(n8732), .ZN(n8206) );
  NAND2_X1 U9831 ( .A1(n8207), .A2(n8404), .ZN(n8209) );
  OR2_X1 U9832 ( .A1(n8402), .A2(n9016), .ZN(n8208) );
  XNOR2_X1 U9833 ( .A(n8879), .B(n8474), .ZN(n8451) );
  INV_X1 U9834 ( .A(n8451), .ZN(n8210) );
  XNOR2_X1 U9835 ( .A(n8211), .B(n8210), .ZN(n8212) );
  NAND2_X1 U9836 ( .A1(n8212), .A2(n8843), .ZN(n8237) );
  NAND2_X1 U9837 ( .A1(n8213), .A2(n8326), .ZN(n8214) );
  NAND2_X1 U9838 ( .A1(n8214), .A2(n8331), .ZN(n8859) );
  NAND2_X1 U9839 ( .A1(n8859), .A2(n8325), .ZN(n8215) );
  INV_X1 U9840 ( .A(n8333), .ZN(n8216) );
  NAND2_X1 U9841 ( .A1(n8992), .A2(n8852), .ZN(n8346) );
  NAND2_X1 U9842 ( .A1(n8338), .A2(n8346), .ZN(n8836) );
  NAND2_X1 U9843 ( .A1(n8833), .A2(n8338), .ZN(n8822) );
  AND2_X1 U9844 ( .A1(n8344), .A2(n8794), .ZN(n8353) );
  NAND2_X1 U9845 ( .A1(n8795), .A2(n8353), .ZN(n8217) );
  INV_X1 U9846 ( .A(n8246), .ZN(n8218) );
  AND2_X1 U9847 ( .A1(n8970), .A2(n8788), .ZN(n8358) );
  NAND2_X1 U9848 ( .A1(n8489), .A2(n8561), .ZN(n8418) );
  OR2_X2 U9849 ( .A1(n8749), .A2(n8364), .ZN(n8221) );
  NAND2_X1 U9850 ( .A1(n8950), .A2(n8576), .ZN(n8368) );
  INV_X1 U9851 ( .A(n8368), .ZN(n8222) );
  NAND2_X1 U9852 ( .A1(n8944), .A2(n8583), .ZN(n8371) );
  INV_X1 U9853 ( .A(n8477), .ZN(n8224) );
  XNOR2_X1 U9854 ( .A(n8887), .B(n8382), .ZN(n8478) );
  NAND2_X1 U9855 ( .A1(n8887), .A2(n8382), .ZN(n8225) );
  AND2_X1 U9856 ( .A1(n8226), .A2(P2_B_REG_SCAN_IN), .ZN(n8227) );
  NOR2_X1 U9857 ( .A1(n10074), .A2(n8227), .ZN(n8714) );
  INV_X1 U9858 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n8232) );
  NAND2_X1 U9859 ( .A1(n8228), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n8231) );
  NAND2_X1 U9860 ( .A1(n8229), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n8230) );
  OAI211_X1 U9861 ( .C1(n8232), .C2(n8412), .A(n8231), .B(n8230), .ZN(n8233)
         );
  INV_X1 U9862 ( .A(n8233), .ZN(n8234) );
  NAND2_X1 U9863 ( .A1(n8416), .A2(n8234), .ZN(n8604) );
  AOI22_X1 U9864 ( .A1(n8732), .A2(n8838), .B1(n8714), .B2(n8604), .ZN(n8235)
         );
  NOR2_X1 U9865 ( .A1(n8727), .A2(n10136), .ZN(n8238) );
  NOR2_X1 U9866 ( .A1(n8720), .A2(n8238), .ZN(n8877) );
  MUX2_X1 U9867 ( .A(n8239), .B(n8877), .S(n10142), .Z(n8241) );
  NAND2_X1 U9868 ( .A1(n8879), .A2(n9004), .ZN(n8240) );
  NAND2_X1 U9869 ( .A1(n8241), .A2(n8240), .ZN(P2_U3456) );
  MUX2_X1 U9870 ( .A(n8374), .B(n8474), .S(n8879), .Z(n8243) );
  OR2_X1 U9871 ( .A1(n8605), .A2(n8388), .ZN(n8242) );
  AND2_X1 U9872 ( .A1(n8418), .A2(n8244), .ZN(n8245) );
  MUX2_X1 U9873 ( .A(n8246), .B(n8245), .S(n8374), .Z(n8355) );
  NOR2_X1 U9874 ( .A1(n8608), .A2(n8388), .ZN(n8247) );
  AND2_X1 U9875 ( .A1(n4431), .A2(n8247), .ZN(n8248) );
  OAI211_X1 U9876 ( .C1(n8441), .C2(n8248), .A(n8338), .B(n8333), .ZN(n8336)
         );
  INV_X1 U9877 ( .A(n8249), .ZN(n8276) );
  AND2_X1 U9878 ( .A1(n8255), .A2(n8250), .ZN(n8251) );
  MUX2_X1 U9879 ( .A(n8252), .B(n8251), .S(n8453), .Z(n8254) );
  OAI21_X1 U9880 ( .B1(n8254), .B2(n8253), .A(n8256), .ZN(n8259) );
  NAND2_X1 U9881 ( .A1(n8256), .A2(n8255), .ZN(n8257) );
  NAND2_X1 U9882 ( .A1(n8257), .A2(n8388), .ZN(n8258) );
  NAND2_X1 U9883 ( .A1(n8259), .A2(n8258), .ZN(n8266) );
  NAND2_X1 U9884 ( .A1(n8277), .A2(n8260), .ZN(n8261) );
  AOI21_X1 U9885 ( .B1(n8266), .B2(n8421), .A(n8261), .ZN(n8264) );
  NAND2_X1 U9886 ( .A1(n8622), .A2(n10097), .ZN(n8262) );
  AND2_X1 U9887 ( .A1(n8270), .A2(n8262), .ZN(n8263) );
  MUX2_X1 U9888 ( .A(n8264), .B(n8263), .S(n8388), .Z(n8268) );
  NAND3_X1 U9889 ( .A1(n8266), .A2(n8421), .A3(n8265), .ZN(n8267) );
  NAND2_X1 U9890 ( .A1(n8268), .A2(n8267), .ZN(n8269) );
  NAND2_X1 U9891 ( .A1(n8269), .A2(n8423), .ZN(n8280) );
  INV_X1 U9892 ( .A(n8270), .ZN(n8272) );
  OAI211_X1 U9893 ( .C1(n8280), .C2(n8272), .A(n8282), .B(n8271), .ZN(n8274)
         );
  OAI211_X1 U9894 ( .C1(n8276), .C2(n8275), .A(n8274), .B(n8273), .ZN(n8285)
         );
  INV_X1 U9895 ( .A(n8277), .ZN(n8279) );
  OAI21_X1 U9896 ( .B1(n8280), .B2(n8279), .A(n8278), .ZN(n8283) );
  AOI21_X1 U9897 ( .B1(n8283), .B2(n8282), .A(n8281), .ZN(n8284) );
  MUX2_X1 U9898 ( .A(n8285), .B(n8284), .S(n8388), .Z(n8301) );
  MUX2_X1 U9899 ( .A(n8287), .B(n8286), .S(n8388), .Z(n8288) );
  OR2_X1 U9900 ( .A1(n8289), .A2(n8288), .ZN(n8296) );
  NOR2_X1 U9901 ( .A1(n8296), .A2(n10078), .ZN(n8300) );
  AND2_X1 U9902 ( .A1(n8291), .A2(n8290), .ZN(n8293) );
  OAI211_X1 U9903 ( .C1(n8296), .C2(n8293), .A(n8302), .B(n8292), .ZN(n8298)
         );
  OAI211_X1 U9904 ( .C1(n8296), .C2(n8295), .A(n8303), .B(n8294), .ZN(n8297)
         );
  MUX2_X1 U9905 ( .A(n8298), .B(n8297), .S(n8374), .Z(n8299) );
  AOI21_X1 U9906 ( .B1(n8301), .B2(n8300), .A(n8299), .ZN(n8310) );
  NAND2_X1 U9907 ( .A1(n8307), .A2(n8302), .ZN(n8305) );
  NAND2_X1 U9908 ( .A1(n8306), .A2(n8303), .ZN(n8304) );
  MUX2_X1 U9909 ( .A(n8305), .B(n8304), .S(n8388), .Z(n8309) );
  MUX2_X1 U9910 ( .A(n8307), .B(n8306), .S(n8374), .Z(n8308) );
  OAI211_X1 U9911 ( .C1(n8310), .C2(n8309), .A(n8308), .B(n8435), .ZN(n8317)
         );
  NAND2_X1 U9912 ( .A1(n8312), .A2(n8311), .ZN(n8313) );
  MUX2_X1 U9913 ( .A(n8314), .B(n8313), .S(n8374), .Z(n8316) );
  NAND3_X1 U9914 ( .A1(n8317), .A2(n8316), .A3(n8315), .ZN(n8323) );
  MUX2_X1 U9915 ( .A(n8319), .B(n8318), .S(n8374), .Z(n8320) );
  NOR2_X1 U9916 ( .A1(n8321), .A2(n8320), .ZN(n8322) );
  NAND2_X1 U9917 ( .A1(n8323), .A2(n8322), .ZN(n8329) );
  NAND3_X1 U9918 ( .A1(n8329), .A2(n8436), .A3(n8324), .ZN(n8327) );
  NAND3_X1 U9919 ( .A1(n8329), .A2(n8436), .A3(n8328), .ZN(n8332) );
  AND4_X1 U9920 ( .A1(n8332), .A2(n8374), .A3(n8331), .A4(n8330), .ZN(n8334)
         );
  NAND3_X1 U9921 ( .A1(n8338), .A2(n8334), .A3(n8333), .ZN(n8335) );
  NAND3_X1 U9922 ( .A1(n8350), .A2(n8337), .A3(n8346), .ZN(n8339) );
  NAND3_X1 U9923 ( .A1(n8339), .A2(n8348), .A3(n8338), .ZN(n8340) );
  NAND3_X1 U9924 ( .A1(n8340), .A2(n8794), .A3(n8347), .ZN(n8341) );
  NAND3_X1 U9925 ( .A1(n8343), .A2(n8342), .A3(n8341), .ZN(n8345) );
  NAND2_X1 U9926 ( .A1(n8347), .A2(n8346), .ZN(n8349) );
  OAI211_X1 U9927 ( .C1(n8350), .C2(n8349), .A(n8443), .B(n8348), .ZN(n8352)
         );
  AOI21_X1 U9928 ( .B1(n8353), .B2(n8352), .A(n8351), .ZN(n8354) );
  NAND3_X1 U9929 ( .A1(n8359), .A2(n8360), .A3(n8419), .ZN(n8356) );
  NAND2_X1 U9930 ( .A1(n8356), .A2(n8357), .ZN(n8363) );
  OAI211_X1 U9931 ( .C1(n8359), .C2(n8358), .A(n8357), .B(n8418), .ZN(n8361)
         );
  NAND2_X1 U9932 ( .A1(n8361), .A2(n8360), .ZN(n8362) );
  MUX2_X1 U9933 ( .A(n8365), .B(n8364), .S(n8388), .Z(n8366) );
  NAND2_X1 U9934 ( .A1(n8367), .A2(n8368), .ZN(n8740) );
  MUX2_X1 U9935 ( .A(n8368), .B(n8367), .S(n8388), .Z(n8369) );
  MUX2_X1 U9936 ( .A(n8371), .B(n8370), .S(n8374), .Z(n8372) );
  NAND2_X1 U9937 ( .A1(n8376), .A2(n8373), .ZN(n8384) );
  MUX2_X1 U9938 ( .A(n8382), .B(n8941), .S(n8374), .Z(n8383) );
  INV_X1 U9939 ( .A(n8383), .ZN(n8375) );
  NAND2_X1 U9940 ( .A1(n8376), .A2(n8375), .ZN(n8377) );
  NAND2_X1 U9941 ( .A1(n8384), .A2(n8377), .ZN(n8387) );
  NAND2_X1 U9942 ( .A1(n8464), .A2(n8404), .ZN(n8379) );
  OR2_X1 U9943 ( .A1(n8402), .A2(n8470), .ZN(n8378) );
  INV_X1 U9944 ( .A(n8876), .ZN(n8935) );
  INV_X1 U9945 ( .A(n8604), .ZN(n8380) );
  AND2_X1 U9946 ( .A1(n8935), .A2(n8380), .ZN(n8385) );
  INV_X1 U9947 ( .A(n8385), .ZN(n8447) );
  NAND2_X1 U9948 ( .A1(n8879), .A2(n8474), .ZN(n8381) );
  NAND2_X1 U9949 ( .A1(n8447), .A2(n8381), .ZN(n8397) );
  AOI21_X1 U9950 ( .B1(n8387), .B2(n8382), .A(n8397), .ZN(n8396) );
  AND2_X1 U9951 ( .A1(n8876), .A2(n8604), .ZN(n8400) );
  NOR2_X1 U9952 ( .A1(n8400), .A2(n8388), .ZN(n8386) );
  INV_X1 U9953 ( .A(n8386), .ZN(n8395) );
  AOI211_X1 U9954 ( .C1(n8389), .C2(n8386), .A(n4501), .B(n8385), .ZN(n8394)
         );
  NAND2_X1 U9955 ( .A1(n8387), .A2(n8941), .ZN(n8392) );
  OR2_X1 U9956 ( .A1(n8879), .A2(n8474), .ZN(n8398) );
  AND2_X1 U9957 ( .A1(n8398), .A2(n8388), .ZN(n8391) );
  INV_X1 U9958 ( .A(n8400), .ZN(n8449) );
  INV_X1 U9959 ( .A(n8389), .ZN(n8390) );
  NAND4_X1 U9960 ( .A1(n8392), .A2(n8391), .A3(n8449), .A4(n8390), .ZN(n8393)
         );
  OAI211_X1 U9961 ( .C1(n8396), .C2(n8395), .A(n8394), .B(n8393), .ZN(n8408)
         );
  OAI21_X1 U9962 ( .B1(n8407), .B2(n8400), .A(n8406), .ZN(n8405) );
  NOR2_X1 U9963 ( .A1(n8402), .A2(n9011), .ZN(n8403) );
  INV_X1 U9964 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n8413) );
  NAND2_X1 U9965 ( .A1(n8228), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n8411) );
  NAND2_X1 U9966 ( .A1(n8409), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n8410) );
  OAI211_X1 U9967 ( .C1(n8413), .C2(n8412), .A(n8411), .B(n8410), .ZN(n8414)
         );
  INV_X1 U9968 ( .A(n8414), .ZN(n8415) );
  NAND2_X1 U9969 ( .A1(n8416), .A2(n8415), .ZN(n8715) );
  INV_X1 U9970 ( .A(n8715), .ZN(n8417) );
  INV_X1 U9971 ( .A(n8728), .ZN(n8730) );
  NAND2_X1 U9972 ( .A1(n8419), .A2(n8418), .ZN(n8775) );
  NOR2_X1 U9973 ( .A1(n8420), .A2(n7056), .ZN(n8424) );
  NAND4_X1 U9974 ( .A1(n8424), .A2(n8423), .A3(n8422), .A4(n8421), .ZN(n8427)
         );
  NOR4_X1 U9975 ( .A1(n8427), .A2(n10078), .A3(n8426), .A4(n8425), .ZN(n8428)
         );
  NAND4_X1 U9976 ( .A1(n8431), .A2(n8430), .A3(n8429), .A4(n8428), .ZN(n8432)
         );
  NOR3_X1 U9977 ( .A1(n8434), .A2(n8433), .A3(n8432), .ZN(n8438) );
  NAND4_X1 U9978 ( .A1(n8438), .A2(n8437), .A3(n8436), .A4(n8435), .ZN(n8439)
         );
  NOR4_X1 U9979 ( .A1(n8836), .A2(n8441), .A3(n8440), .A4(n8439), .ZN(n8442)
         );
  NAND4_X1 U9980 ( .A1(n8444), .A2(n8443), .A3(n8823), .A4(n8442), .ZN(n8445)
         );
  OR4_X1 U9981 ( .A1(n8769), .A2(n8775), .A3(n8786), .A4(n8445), .ZN(n8446) );
  NOR4_X1 U9982 ( .A1(n8730), .A2(n8751), .A3(n8740), .A4(n8446), .ZN(n8448)
         );
  NAND4_X1 U9983 ( .A1(n8449), .A2(n8448), .A3(n8447), .A4(n8223), .ZN(n8450)
         );
  AOI211_X1 U9984 ( .C1(n8932), .C2(n8715), .A(n8451), .B(n8450), .ZN(n8454)
         );
  NOR4_X1 U9985 ( .A1(n8458), .A2(n8697), .A3(n8457), .A4(n8456), .ZN(n8461)
         );
  OAI21_X1 U9986 ( .B1(n8462), .B2(n8459), .A(P2_B_REG_SCAN_IN), .ZN(n8460) );
  OAI22_X1 U9987 ( .A1(n8463), .A2(n8462), .B1(n8461), .B2(n8460), .ZN(
        P2_U3296) );
  INV_X1 U9988 ( .A(n8464), .ZN(n8469) );
  OAI222_X1 U9989 ( .A1(n8071), .A2(n8465), .B1(n9797), .B2(n8469), .C1(
        P1_U3086), .C2(n5129), .ZN(P1_U3325) );
  INV_X1 U9990 ( .A(n6293), .ZN(n9023) );
  OAI222_X1 U9991 ( .A1(n9797), .A2(n9023), .B1(n8467), .B2(P1_U3086), .C1(
        n8466), .C2(n8071), .ZN(P1_U3327) );
  OAI222_X1 U9992 ( .A1(n9015), .A2(n8470), .B1(n9022), .B2(n8469), .C1(n8468), 
        .C2(P2_U3151), .ZN(P2_U3265) );
  OAI222_X1 U9993 ( .A1(n8071), .A2(n8472), .B1(n9797), .B2(n8471), .C1(n9373), 
        .C2(P1_U3086), .ZN(P1_U3336) );
  XNOR2_X1 U9994 ( .A(n8473), .B(n8478), .ZN(n8476) );
  OAI22_X1 U9995 ( .A1(n8474), .A2(n10074), .B1(n8583), .B2(n10076), .ZN(n8475) );
  AOI22_X1 U9996 ( .A1(n8481), .A2(n10087), .B1(n10092), .B2(
        P2_REG2_REG_28__SCAN_IN), .ZN(n8482) );
  OAI21_X1 U9997 ( .B1(n8941), .B2(n8779), .A(n8482), .ZN(n8483) );
  AOI21_X1 U9998 ( .B1(n4337), .B2(n8819), .A(n8483), .ZN(n8484) );
  OAI21_X1 U9999 ( .B1(n8883), .B2(n10092), .A(n8484), .ZN(P2_U3205) );
  AOI21_X1 U10000 ( .B1(n8788), .B2(n8485), .A(n4321), .ZN(n8491) );
  AOI22_X1 U10001 ( .A1(n8607), .A2(n8579), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3151), .ZN(n8487) );
  NAND2_X1 U10002 ( .A1(n8777), .A2(n8598), .ZN(n8486) );
  OAI211_X1 U10003 ( .C1(n8774), .C2(n8582), .A(n8487), .B(n8486), .ZN(n8488)
         );
  AOI21_X1 U10004 ( .B1(n8489), .B2(n8585), .A(n8488), .ZN(n8490) );
  OAI21_X1 U10005 ( .B1(n8491), .B2(n8573), .A(n8490), .ZN(P2_U3156) );
  XNOR2_X1 U10006 ( .A(n8823), .B(n5951), .ZN(n8492) );
  XNOR2_X1 U10007 ( .A(n8493), .B(n8492), .ZN(n8498) );
  NAND2_X1 U10008 ( .A1(n8593), .A2(n8826), .ZN(n8494) );
  NAND2_X1 U10009 ( .A1(P2_U3151), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8710) );
  OAI211_X1 U10010 ( .C1(n8852), .C2(n8595), .A(n8494), .B(n8710), .ZN(n8495)
         );
  AOI21_X1 U10011 ( .B1(n8829), .B2(n8598), .A(n8495), .ZN(n8497) );
  NAND2_X1 U10012 ( .A1(n8986), .A2(n8585), .ZN(n8496) );
  OAI211_X1 U10013 ( .C1(n8498), .C2(n8573), .A(n8497), .B(n8496), .ZN(
        P2_U3159) );
  INV_X1 U10014 ( .A(n8499), .ZN(n8504) );
  NOR3_X1 U10015 ( .A1(n8500), .A2(n8502), .A3(n8501), .ZN(n8503) );
  OAI21_X1 U10016 ( .B1(n8504), .B2(n8503), .A(n8589), .ZN(n8508) );
  AOI22_X1 U10017 ( .A1(n8607), .A2(n8593), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3151), .ZN(n8505) );
  OAI21_X1 U10018 ( .B1(n8802), .B2(n8595), .A(n8505), .ZN(n8506) );
  AOI21_X1 U10019 ( .B1(n8804), .B2(n8598), .A(n8506), .ZN(n8507) );
  OAI211_X1 U10020 ( .C1(n8910), .C2(n8602), .A(n8508), .B(n8507), .ZN(
        P2_U3163) );
  OAI21_X1 U10021 ( .B1(n8511), .B2(n8510), .A(n8509), .ZN(n8512) );
  NAND2_X1 U10022 ( .A1(n8512), .A2(n8589), .ZN(n8518) );
  INV_X1 U10023 ( .A(n8513), .ZN(n8756) );
  AOI22_X1 U10024 ( .A1(n8606), .A2(n8579), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3151), .ZN(n8514) );
  OAI21_X1 U10025 ( .B1(n8756), .B2(n8515), .A(n8514), .ZN(n8516) );
  AOI21_X1 U10026 ( .B1(n8593), .B2(n8753), .A(n8516), .ZN(n8517) );
  OAI211_X1 U10027 ( .C1(n8955), .C2(n8602), .A(n8518), .B(n8517), .ZN(
        P2_U3165) );
  AOI21_X1 U10028 ( .B1(n8521), .B2(n8520), .A(n8519), .ZN(n8526) );
  AOI22_X1 U10029 ( .A1(n8593), .A2(n8839), .B1(P2_REG3_REG_16__SCAN_IN), .B2(
        P2_U3151), .ZN(n8523) );
  NAND2_X1 U10030 ( .A1(n8598), .A2(n8869), .ZN(n8522) );
  OAI211_X1 U10031 ( .C1(n8863), .C2(n8595), .A(n8523), .B(n8522), .ZN(n8524)
         );
  AOI21_X1 U10032 ( .B1(n4431), .B2(n8585), .A(n8524), .ZN(n8525) );
  OAI21_X1 U10033 ( .B1(n8526), .B2(n8573), .A(n8525), .ZN(P2_U3166) );
  NAND2_X1 U10034 ( .A1(n8528), .A2(n8527), .ZN(n8530) );
  XOR2_X1 U10035 ( .A(n8530), .B(n8529), .Z(n8535) );
  NAND2_X1 U10036 ( .A1(n8593), .A2(n8825), .ZN(n8531) );
  NAND2_X1 U10037 ( .A1(P2_U3151), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n10066)
         );
  OAI211_X1 U10038 ( .C1(n8853), .C2(n8595), .A(n8531), .B(n10066), .ZN(n8532)
         );
  AOI21_X1 U10039 ( .B1(n8856), .B2(n8598), .A(n8532), .ZN(n8534) );
  NAND2_X1 U10040 ( .A1(n8998), .A2(n8585), .ZN(n8533) );
  OAI211_X1 U10041 ( .C1(n8535), .C2(n8573), .A(n8534), .B(n8533), .ZN(
        P2_U3168) );
  INV_X1 U10042 ( .A(n8536), .ZN(n8538) );
  NOR3_X1 U10043 ( .A1(n4321), .A2(n8538), .A3(n8537), .ZN(n8541) );
  INV_X1 U10044 ( .A(n8539), .ZN(n8540) );
  OAI21_X1 U10045 ( .B1(n8541), .B2(n8540), .A(n8589), .ZN(n8546) );
  OAI22_X1 U10046 ( .A1(n8561), .A2(n8595), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8542), .ZN(n8544) );
  NOR2_X1 U10047 ( .A1(n8765), .A2(n8582), .ZN(n8543) );
  AOI211_X1 U10048 ( .C1(n8767), .C2(n8598), .A(n8544), .B(n8543), .ZN(n8545)
         );
  OAI211_X1 U10049 ( .C1(n8898), .C2(n8602), .A(n8546), .B(n8545), .ZN(
        P2_U3169) );
  INV_X1 U10050 ( .A(n8913), .ZN(n8554) );
  NOR2_X1 U10051 ( .A1(n8548), .A2(n8547), .ZN(n8549) );
  OAI21_X1 U10052 ( .B1(n8549), .B2(n8500), .A(n8589), .ZN(n8553) );
  AOI22_X1 U10053 ( .A1(n8810), .A2(n8593), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3151), .ZN(n8550) );
  OAI21_X1 U10054 ( .B1(n8570), .B2(n8595), .A(n8550), .ZN(n8551) );
  AOI21_X1 U10055 ( .B1(n8812), .B2(n8598), .A(n8551), .ZN(n8552) );
  OAI211_X1 U10056 ( .C1(n8554), .C2(n8602), .A(n8553), .B(n8552), .ZN(
        P2_U3173) );
  OAI21_X1 U10057 ( .B1(n8557), .B2(n8556), .A(n8555), .ZN(n8558) );
  NAND2_X1 U10058 ( .A1(n8558), .A2(n8589), .ZN(n8565) );
  INV_X1 U10059 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n8559) );
  OAI22_X1 U10060 ( .A1(n8560), .A2(n8595), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8559), .ZN(n8563) );
  NOR2_X1 U10061 ( .A1(n8561), .A2(n8582), .ZN(n8562) );
  AOI211_X1 U10062 ( .C1(n8791), .C2(n8598), .A(n8563), .B(n8562), .ZN(n8564)
         );
  OAI211_X1 U10063 ( .C1(n8199), .C2(n8602), .A(n8565), .B(n8564), .ZN(
        P2_U3175) );
  XOR2_X1 U10064 ( .A(n8567), .B(n8566), .Z(n8574) );
  AND2_X1 U10065 ( .A1(P2_U3151), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8656) );
  AOI21_X1 U10066 ( .B1(n8579), .B2(n8839), .A(n8656), .ZN(n8569) );
  NAND2_X1 U10067 ( .A1(n8598), .A2(n8845), .ZN(n8568) );
  OAI211_X1 U10068 ( .C1(n8570), .C2(n8582), .A(n8569), .B(n8568), .ZN(n8571)
         );
  AOI21_X1 U10069 ( .B1(n8992), .B2(n8585), .A(n8571), .ZN(n8572) );
  OAI21_X1 U10070 ( .B1(n8574), .B2(n8573), .A(n8572), .ZN(P2_U3178) );
  NOR2_X1 U10071 ( .A1(n8575), .A2(n8576), .ZN(n8578) );
  OAI21_X1 U10072 ( .B1(n8578), .B2(n8577), .A(n8589), .ZN(n8587) );
  AOI22_X1 U10073 ( .A1(n8741), .A2(n8579), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3151), .ZN(n8581) );
  NAND2_X1 U10074 ( .A1(n8745), .A2(n8598), .ZN(n8580) );
  OAI211_X1 U10075 ( .C1(n8583), .C2(n8582), .A(n8581), .B(n8580), .ZN(n8584)
         );
  AOI21_X1 U10076 ( .B1(n8950), .B2(n8585), .A(n8584), .ZN(n8586) );
  NAND2_X1 U10077 ( .A1(n8587), .A2(n8586), .ZN(P2_U3180) );
  INV_X1 U10078 ( .A(n8588), .ZN(n8603) );
  OAI211_X1 U10079 ( .C1(n8592), .C2(n8591), .A(n8590), .B(n8589), .ZN(n8601)
         );
  NAND2_X1 U10080 ( .A1(n8593), .A2(n8608), .ZN(n8594) );
  NAND2_X1 U10081 ( .A1(P2_U3151), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n10030)
         );
  OAI211_X1 U10082 ( .C1(n8596), .C2(n8595), .A(n8594), .B(n10030), .ZN(n8597)
         );
  AOI21_X1 U10083 ( .B1(n8599), .B2(n8598), .A(n8597), .ZN(n8600) );
  OAI211_X1 U10084 ( .C1(n8603), .C2(n8602), .A(n8601), .B(n8600), .ZN(
        P2_U3181) );
  MUX2_X1 U10085 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n8715), .S(P2_U3893), .Z(
        P2_U3522) );
  MUX2_X1 U10086 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n8604), .S(P2_U3893), .Z(
        P2_U3521) );
  MUX2_X1 U10087 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n8605), .S(P2_U3893), .Z(
        P2_U3520) );
  MUX2_X1 U10088 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n8732), .S(P2_U3893), .Z(
        P2_U3519) );
  MUX2_X1 U10089 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8742), .S(P2_U3893), .Z(
        P2_U3518) );
  MUX2_X1 U10090 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n8753), .S(P2_U3893), .Z(
        P2_U3517) );
  MUX2_X1 U10091 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8741), .S(P2_U3893), .Z(
        P2_U3516) );
  MUX2_X1 U10092 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n8606), .S(P2_U3893), .Z(
        P2_U3515) );
  MUX2_X1 U10093 ( .A(n8788), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8623), .Z(
        P2_U3514) );
  MUX2_X1 U10094 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8607), .S(P2_U3893), .Z(
        P2_U3513) );
  MUX2_X1 U10095 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8810), .S(P2_U3893), .Z(
        P2_U3512) );
  MUX2_X1 U10096 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8826), .S(P2_U3893), .Z(
        P2_U3511) );
  MUX2_X1 U10097 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8841), .S(P2_U3893), .Z(
        P2_U3510) );
  MUX2_X1 U10098 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n8825), .S(P2_U3893), .Z(
        P2_U3509) );
  MUX2_X1 U10099 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8839), .S(P2_U3893), .Z(
        P2_U3508) );
  MUX2_X1 U10100 ( .A(n8608), .B(P2_DATAO_REG_16__SCAN_IN), .S(n8623), .Z(
        P2_U3507) );
  MUX2_X1 U10101 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n8609), .S(P2_U3893), .Z(
        P2_U3506) );
  MUX2_X1 U10102 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n8610), .S(P2_U3893), .Z(
        P2_U3505) );
  MUX2_X1 U10103 ( .A(n8611), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8623), .Z(
        P2_U3504) );
  MUX2_X1 U10104 ( .A(n8612), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8623), .Z(
        P2_U3503) );
  MUX2_X1 U10105 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n8613), .S(P2_U3893), .Z(
        P2_U3502) );
  MUX2_X1 U10106 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n8614), .S(P2_U3893), .Z(
        P2_U3501) );
  MUX2_X1 U10107 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n8615), .S(P2_U3893), .Z(
        P2_U3500) );
  MUX2_X1 U10108 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n8616), .S(P2_U3893), .Z(
        P2_U3499) );
  MUX2_X1 U10109 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n8617), .S(P2_U3893), .Z(
        P2_U3498) );
  MUX2_X1 U10110 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n8618), .S(P2_U3893), .Z(
        P2_U3497) );
  MUX2_X1 U10111 ( .A(n8619), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8623), .Z(
        P2_U3496) );
  MUX2_X1 U10112 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n8620), .S(P2_U3893), .Z(
        P2_U3495) );
  MUX2_X1 U10113 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(n8621), .S(P2_U3893), .Z(
        P2_U3494) );
  MUX2_X1 U10114 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(n8622), .S(P2_U3893), .Z(
        P2_U3493) );
  MUX2_X1 U10115 ( .A(n8624), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8623), .Z(
        P2_U3492) );
  XNOR2_X1 U10116 ( .A(n8688), .B(P2_REG1_REG_18__SCAN_IN), .ZN(n8701) );
  INV_X1 U10117 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8926) );
  AOI22_X1 U10118 ( .A1(P2_REG1_REG_16__SCAN_IN), .A2(n8646), .B1(n10033), 
        .B2(n8926), .ZN(n10036) );
  NAND2_X1 U10119 ( .A1(P2_REG1_REG_14__SCAN_IN), .A2(n8641), .ZN(n8630) );
  AOI22_X1 U10120 ( .A1(P2_REG1_REG_14__SCAN_IN), .A2(n8641), .B1(n10002), 
        .B2(n8625), .ZN(n10005) );
  NAND2_X1 U10121 ( .A1(P2_REG1_REG_12__SCAN_IN), .A2(n8637), .ZN(n8627) );
  NAND2_X1 U10122 ( .A1(n8662), .A2(n8628), .ZN(n8629) );
  XNOR2_X1 U10123 ( .A(n9984), .B(n8628), .ZN(n9986) );
  NAND2_X1 U10124 ( .A1(P2_REG1_REG_13__SCAN_IN), .A2(n9986), .ZN(n9985) );
  NAND2_X1 U10125 ( .A1(n8629), .A2(n9985), .ZN(n10004) );
  NAND2_X1 U10126 ( .A1(n10005), .A2(n10004), .ZN(n10003) );
  NAND2_X1 U10127 ( .A1(n8630), .A2(n10003), .ZN(n8632) );
  NAND2_X1 U10128 ( .A1(n8631), .A2(n8632), .ZN(n8633) );
  XNOR2_X1 U10129 ( .A(n10017), .B(n8632), .ZN(n10019) );
  NAND2_X1 U10130 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n10019), .ZN(n10018) );
  NAND2_X1 U10131 ( .A1(n8633), .A2(n10018), .ZN(n10035) );
  NAND2_X1 U10132 ( .A1(n8678), .A2(n8634), .ZN(n8635) );
  XNOR2_X1 U10133 ( .A(n10050), .B(n8634), .ZN(n10053) );
  NAND2_X1 U10134 ( .A1(P2_REG1_REG_17__SCAN_IN), .A2(n10053), .ZN(n10052) );
  NAND2_X1 U10135 ( .A1(n8635), .A2(n10052), .ZN(n8702) );
  XOR2_X1 U10136 ( .A(n8701), .B(n8702), .Z(n8694) );
  INV_X1 U10137 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8844) );
  NOR2_X1 U10138 ( .A1(n8688), .A2(n8844), .ZN(n8706) );
  AOI21_X1 U10139 ( .B1(n8688), .B2(n8844), .A(n8706), .ZN(n8652) );
  NOR2_X1 U10140 ( .A1(n9984), .A2(n8638), .ZN(n8639) );
  INV_X1 U10141 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n9995) );
  NAND2_X1 U10142 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n8641), .ZN(n8640) );
  OAI21_X1 U10143 ( .B1(n8641), .B2(P2_REG2_REG_14__SCAN_IN), .A(n8640), .ZN(
        n10011) );
  NOR2_X1 U10144 ( .A1(n10017), .A2(n8642), .ZN(n8644) );
  NAND2_X1 U10145 ( .A1(P2_REG2_REG_16__SCAN_IN), .A2(n8646), .ZN(n8645) );
  OAI21_X1 U10146 ( .B1(n8646), .B2(P2_REG2_REG_16__SCAN_IN), .A(n8645), .ZN(
        n10043) );
  INV_X1 U10147 ( .A(n8647), .ZN(n8648) );
  NAND2_X1 U10148 ( .A1(n8678), .A2(n8648), .ZN(n8649) );
  OAI21_X1 U10149 ( .B1(n8678), .B2(n8648), .A(n8649), .ZN(n10062) );
  INV_X1 U10150 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n10061) );
  OAI21_X1 U10151 ( .B1(n8652), .B2(n8651), .A(n8708), .ZN(n8657) );
  INV_X1 U10152 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n8653) );
  NOR2_X1 U10153 ( .A1(n8654), .A2(n8653), .ZN(n8655) );
  AOI211_X1 U10154 ( .C1(n10026), .C2(n8657), .A(n8656), .B(n8655), .ZN(n8692)
         );
  OR2_X1 U10155 ( .A1(n8659), .A2(n8658), .ZN(n8661) );
  NAND2_X1 U10156 ( .A1(n8661), .A2(n8660), .ZN(n9988) );
  MUX2_X1 U10157 ( .A(P2_REG1_REG_13__SCAN_IN), .B(P2_REG2_REG_13__SCAN_IN), 
        .S(n8697), .Z(n8663) );
  XNOR2_X1 U10158 ( .A(n8663), .B(n8662), .ZN(n9987) );
  INV_X1 U10159 ( .A(n8663), .ZN(n8664) );
  NAND2_X1 U10160 ( .A1(n8664), .A2(n9984), .ZN(n8665) );
  NAND2_X1 U10161 ( .A1(n9991), .A2(n8665), .ZN(n10007) );
  MUX2_X1 U10162 ( .A(P2_REG1_REG_14__SCAN_IN), .B(P2_REG2_REG_14__SCAN_IN), 
        .S(n8697), .Z(n8666) );
  XNOR2_X1 U10163 ( .A(n8666), .B(n10002), .ZN(n10006) );
  NAND2_X1 U10164 ( .A1(n10007), .A2(n10006), .ZN(n8669) );
  INV_X1 U10165 ( .A(n8666), .ZN(n8667) );
  NAND2_X1 U10166 ( .A1(n8667), .A2(n10002), .ZN(n8668) );
  NAND2_X1 U10167 ( .A1(n8669), .A2(n8668), .ZN(n10021) );
  MUX2_X1 U10168 ( .A(P2_REG1_REG_15__SCAN_IN), .B(P2_REG2_REG_15__SCAN_IN), 
        .S(n8697), .Z(n8670) );
  XNOR2_X1 U10169 ( .A(n8670), .B(n10017), .ZN(n10020) );
  NAND2_X1 U10170 ( .A1(n10021), .A2(n10020), .ZN(n8673) );
  INV_X1 U10171 ( .A(n8670), .ZN(n8671) );
  NAND2_X1 U10172 ( .A1(n8671), .A2(n10017), .ZN(n8672) );
  NAND2_X1 U10173 ( .A1(n8673), .A2(n8672), .ZN(n10038) );
  MUX2_X1 U10174 ( .A(P2_REG1_REG_16__SCAN_IN), .B(P2_REG2_REG_16__SCAN_IN), 
        .S(n8697), .Z(n8674) );
  XNOR2_X1 U10175 ( .A(n8674), .B(n10033), .ZN(n10037) );
  NAND2_X1 U10176 ( .A1(n10038), .A2(n10037), .ZN(n8677) );
  INV_X1 U10177 ( .A(n8674), .ZN(n8675) );
  NAND2_X1 U10178 ( .A1(n8675), .A2(n10033), .ZN(n8676) );
  NAND2_X1 U10179 ( .A1(n8677), .A2(n8676), .ZN(n10055) );
  MUX2_X1 U10180 ( .A(P2_REG1_REG_17__SCAN_IN), .B(P2_REG2_REG_17__SCAN_IN), 
        .S(n8697), .Z(n8679) );
  XNOR2_X1 U10181 ( .A(n8679), .B(n10050), .ZN(n10054) );
  NOR2_X1 U10182 ( .A1(n8679), .A2(n8678), .ZN(n8680) );
  AOI21_X1 U10183 ( .B1(n10055), .B2(n10054), .A(n8680), .ZN(n8681) );
  MUX2_X1 U10184 ( .A(P2_REG1_REG_18__SCAN_IN), .B(P2_REG2_REG_18__SCAN_IN), 
        .S(n8697), .Z(n8682) );
  AND2_X1 U10185 ( .A1(n8681), .A2(n8682), .ZN(n8696) );
  INV_X1 U10186 ( .A(n8681), .ZN(n8684) );
  INV_X1 U10187 ( .A(n8682), .ZN(n8683) );
  NAND2_X1 U10188 ( .A1(n8684), .A2(n8683), .ZN(n8695) );
  INV_X1 U10189 ( .A(n8695), .ZN(n8685) );
  OR2_X1 U10190 ( .A1(n8696), .A2(n8685), .ZN(n8686) );
  NAND2_X1 U10191 ( .A1(n8686), .A2(n10057), .ZN(n8690) );
  INV_X1 U10192 ( .A(n8686), .ZN(n8687) );
  AOI21_X1 U10193 ( .B1(n8687), .B2(P2_U3893), .A(n10051), .ZN(n8689) );
  MUX2_X1 U10194 ( .A(n8690), .B(n8689), .S(n8688), .Z(n8691) );
  OAI211_X1 U10195 ( .C1(n8694), .C2(n8693), .A(n8692), .B(n8691), .ZN(
        P2_U3200) );
  OAI21_X1 U10196 ( .B1(n8696), .B2(n8700), .A(n8695), .ZN(n8699) );
  XNOR2_X1 U10197 ( .A(n8711), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n8703) );
  XNOR2_X1 U10198 ( .A(n8711), .B(P2_REG2_REG_19__SCAN_IN), .ZN(n8709) );
  MUX2_X1 U10199 ( .A(n8703), .B(n8709), .S(n8697), .Z(n8698) );
  AOI22_X1 U10200 ( .A1(n8702), .A2(n8701), .B1(P2_REG1_REG_18__SCAN_IN), .B2(
        n8700), .ZN(n8704) );
  XNOR2_X1 U10201 ( .A(n8704), .B(n8703), .ZN(n8705) );
  NAND2_X1 U10202 ( .A1(n8705), .A2(n10058), .ZN(n8713) );
  INV_X1 U10203 ( .A(n8706), .ZN(n8707) );
  AND2_X1 U10204 ( .A1(n8716), .A2(n10087), .ZN(n8723) );
  AOI21_X1 U10205 ( .B1(n8933), .B2(n8867), .A(n8723), .ZN(n8719) );
  NAND2_X1 U10206 ( .A1(n10092), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n8717) );
  OAI211_X1 U10207 ( .C1(n8932), .C2(n8779), .A(n8719), .B(n8717), .ZN(
        P2_U3202) );
  NAND2_X1 U10208 ( .A1(n10092), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n8718) );
  OAI211_X1 U10209 ( .C1(n8876), .C2(n8779), .A(n8719), .B(n8718), .ZN(
        P2_U3203) );
  NAND2_X1 U10210 ( .A1(n8720), .A2(n8867), .ZN(n8725) );
  INV_X1 U10211 ( .A(n8879), .ZN(n8721) );
  NOR2_X1 U10212 ( .A1(n8721), .A2(n8779), .ZN(n8722) );
  AOI211_X1 U10213 ( .C1(n10092), .C2(P2_REG2_REG_29__SCAN_IN), .A(n8723), .B(
        n8722), .ZN(n8724) );
  OAI211_X1 U10214 ( .C1(n8727), .C2(n8726), .A(n8725), .B(n8724), .ZN(
        P2_U3204) );
  XNOR2_X1 U10215 ( .A(n8729), .B(n8728), .ZN(n8947) );
  INV_X1 U10216 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n8734) );
  XNOR2_X1 U10217 ( .A(n8731), .B(n8730), .ZN(n8733) );
  AOI222_X1 U10218 ( .A1(n8843), .A2(n8733), .B1(n8732), .B2(n8840), .C1(n8753), .C2(n8838), .ZN(n8942) );
  MUX2_X1 U10219 ( .A(n8734), .B(n8942), .S(n10091), .Z(n8737) );
  AOI22_X1 U10220 ( .A1(n8944), .A2(n10085), .B1(n10087), .B2(n8735), .ZN(
        n8736) );
  OAI211_X1 U10221 ( .C1(n8947), .C2(n8872), .A(n8737), .B(n8736), .ZN(
        P2_U3206) );
  XNOR2_X1 U10222 ( .A(n8738), .B(n8740), .ZN(n8953) );
  INV_X1 U10223 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n8744) );
  XOR2_X1 U10224 ( .A(n8740), .B(n8739), .Z(n8743) );
  AOI222_X1 U10225 ( .A1(n8843), .A2(n8743), .B1(n8742), .B2(n8840), .C1(n8741), .C2(n8838), .ZN(n8948) );
  MUX2_X1 U10226 ( .A(n8744), .B(n8948), .S(n10091), .Z(n8747) );
  AOI22_X1 U10227 ( .A1(n8950), .A2(n10085), .B1(n10087), .B2(n8745), .ZN(
        n8746) );
  OAI211_X1 U10228 ( .C1(n8953), .C2(n8872), .A(n8747), .B(n8746), .ZN(
        P2_U3207) );
  XNOR2_X1 U10229 ( .A(n8749), .B(n8748), .ZN(n8956) );
  OAI211_X1 U10230 ( .C1(n8752), .C2(n8751), .A(n8750), .B(n8843), .ZN(n8755)
         );
  NAND2_X1 U10231 ( .A1(n8753), .A2(n8840), .ZN(n8754) );
  OAI211_X1 U10232 ( .C1(n8774), .C2(n10076), .A(n8755), .B(n8754), .ZN(n8954)
         );
  OAI22_X1 U10233 ( .A1(n8955), .A2(n8760), .B1(n8756), .B2(n8813), .ZN(n8757)
         );
  OAI21_X1 U10234 ( .B1(n8954), .B2(n8757), .A(n8867), .ZN(n8759) );
  NAND2_X1 U10235 ( .A1(n10092), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n8758) );
  OAI211_X1 U10236 ( .C1(n8956), .C2(n8872), .A(n8759), .B(n8758), .ZN(
        P2_U3208) );
  NOR2_X1 U10237 ( .A1(n8898), .A2(n8760), .ZN(n8766) );
  OAI211_X1 U10238 ( .C1(n8762), .C2(n8769), .A(n8761), .B(n8843), .ZN(n8764)
         );
  NAND2_X1 U10239 ( .A1(n8788), .A2(n8838), .ZN(n8763) );
  OAI211_X1 U10240 ( .C1(n8765), .C2(n10074), .A(n8764), .B(n8763), .ZN(n8959)
         );
  AOI211_X1 U10241 ( .C1(n10087), .C2(n8767), .A(n8766), .B(n8959), .ZN(n8771)
         );
  XOR2_X1 U10242 ( .A(n8769), .B(n8768), .Z(n8897) );
  AOI22_X1 U10243 ( .A1(n8897), .A2(n8819), .B1(P2_REG2_REG_24__SCAN_IN), .B2(
        n10092), .ZN(n8770) );
  OAI21_X1 U10244 ( .B1(n8771), .B2(n10092), .A(n8770), .ZN(P2_U3209) );
  XOR2_X1 U10245 ( .A(n8775), .B(n8772), .Z(n8773) );
  OAI222_X1 U10246 ( .A1(n10074), .A2(n8774), .B1(n10076), .B2(n8801), .C1(
        n10080), .C2(n8773), .ZN(n8901) );
  INV_X1 U10247 ( .A(n8901), .ZN(n8782) );
  XOR2_X1 U10248 ( .A(n8776), .B(n8775), .Z(n8902) );
  AOI22_X1 U10249 ( .A1(n10092), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n8777), 
        .B2(n10087), .ZN(n8778) );
  OAI21_X1 U10250 ( .B1(n8970), .B2(n8779), .A(n8778), .ZN(n8780) );
  AOI21_X1 U10251 ( .B1(n8902), .B2(n8819), .A(n8780), .ZN(n8781) );
  OAI21_X1 U10252 ( .B1(n8782), .B2(n10092), .A(n8781), .ZN(P2_U3210) );
  XNOR2_X1 U10253 ( .A(n8784), .B(n8783), .ZN(n8976) );
  INV_X1 U10254 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n8790) );
  OAI21_X1 U10255 ( .B1(n8787), .B2(n8786), .A(n8785), .ZN(n8789) );
  AOI222_X1 U10256 ( .A1(n8843), .A2(n8789), .B1(n8810), .B2(n8838), .C1(n8788), .C2(n8840), .ZN(n8971) );
  MUX2_X1 U10257 ( .A(n8790), .B(n8971), .S(n10091), .Z(n8793) );
  AOI22_X1 U10258 ( .A1(n8973), .A2(n10085), .B1(n10087), .B2(n8791), .ZN(
        n8792) );
  OAI211_X1 U10259 ( .C1(n8976), .C2(n8872), .A(n8793), .B(n8792), .ZN(
        P2_U3211) );
  NAND2_X1 U10260 ( .A1(n8795), .A2(n8794), .ZN(n8796) );
  XNOR2_X1 U10261 ( .A(n8796), .B(n8797), .ZN(n8982) );
  INV_X1 U10262 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n8803) );
  NOR3_X1 U10263 ( .A1(n8807), .A2(n8798), .A3(n8797), .ZN(n8799) );
  NOR2_X1 U10264 ( .A1(n4344), .A2(n8799), .ZN(n8800) );
  OAI222_X1 U10265 ( .A1(n10076), .A2(n8802), .B1(n10074), .B2(n8801), .C1(
        n10080), .C2(n8800), .ZN(n8908) );
  INV_X1 U10266 ( .A(n8908), .ZN(n8977) );
  MUX2_X1 U10267 ( .A(n8803), .B(n8977), .S(n10091), .Z(n8806) );
  AOI22_X1 U10268 ( .A1(n8979), .A2(n10085), .B1(n10087), .B2(n8804), .ZN(
        n8805) );
  OAI211_X1 U10269 ( .C1(n8982), .C2(n8872), .A(n8806), .B(n8805), .ZN(
        P2_U3212) );
  INV_X1 U10270 ( .A(n8807), .ZN(n8808) );
  OAI21_X1 U10271 ( .B1(n8809), .B2(n8817), .A(n8808), .ZN(n8811) );
  AOI222_X1 U10272 ( .A1(n8843), .A2(n8811), .B1(n8810), .B2(n8840), .C1(n8841), .C2(n8838), .ZN(n8916) );
  INV_X1 U10273 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n8815) );
  INV_X1 U10274 ( .A(n8812), .ZN(n8814) );
  OAI22_X1 U10275 ( .A1(n8867), .A2(n8815), .B1(n8814), .B2(n8813), .ZN(n8816)
         );
  AOI21_X1 U10276 ( .B1(n8913), .B2(n10085), .A(n8816), .ZN(n8821) );
  XNOR2_X1 U10277 ( .A(n8818), .B(n8817), .ZN(n8914) );
  NAND2_X1 U10278 ( .A1(n8914), .A2(n8819), .ZN(n8820) );
  OAI211_X1 U10279 ( .C1(n8916), .C2(n10092), .A(n8821), .B(n8820), .ZN(
        P2_U3213) );
  XNOR2_X1 U10280 ( .A(n8822), .B(n8823), .ZN(n8989) );
  INV_X1 U10281 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n8828) );
  XNOR2_X1 U10282 ( .A(n8824), .B(n8823), .ZN(n8827) );
  AOI222_X1 U10283 ( .A1(n8843), .A2(n8827), .B1(n8826), .B2(n8840), .C1(n8825), .C2(n8838), .ZN(n8984) );
  MUX2_X1 U10284 ( .A(n8828), .B(n8984), .S(n10091), .Z(n8831) );
  AOI22_X1 U10285 ( .A1(n8986), .A2(n10085), .B1(n10087), .B2(n8829), .ZN(
        n8830) );
  OAI211_X1 U10286 ( .C1(n8989), .C2(n8872), .A(n8831), .B(n8830), .ZN(
        P2_U3214) );
  INV_X1 U10287 ( .A(n8832), .ZN(n8835) );
  INV_X1 U10288 ( .A(n8836), .ZN(n8834) );
  OAI21_X1 U10289 ( .B1(n8835), .B2(n8834), .A(n8833), .ZN(n8995) );
  XNOR2_X1 U10290 ( .A(n8837), .B(n8836), .ZN(n8842) );
  AOI222_X1 U10291 ( .A1(n8843), .A2(n8842), .B1(n8841), .B2(n8840), .C1(n8839), .C2(n8838), .ZN(n8990) );
  MUX2_X1 U10292 ( .A(n8844), .B(n8990), .S(n10091), .Z(n8847) );
  AOI22_X1 U10293 ( .A1(n8992), .A2(n10085), .B1(n10087), .B2(n8845), .ZN(
        n8846) );
  OAI211_X1 U10294 ( .C1(n8995), .C2(n8872), .A(n8847), .B(n8846), .ZN(
        P2_U3215) );
  XNOR2_X1 U10295 ( .A(n8848), .B(n8851), .ZN(n9001) );
  AOI211_X1 U10296 ( .C1(n8851), .C2(n8850), .A(n10080), .B(n8849), .ZN(n8855)
         );
  OAI22_X1 U10297 ( .A1(n8853), .A2(n10076), .B1(n8852), .B2(n10074), .ZN(
        n8854) );
  NOR2_X1 U10298 ( .A1(n8855), .A2(n8854), .ZN(n8996) );
  MUX2_X1 U10299 ( .A(n10061), .B(n8996), .S(n8867), .Z(n8858) );
  AOI22_X1 U10300 ( .A1(n8998), .A2(n10085), .B1(n10087), .B2(n8856), .ZN(
        n8857) );
  OAI211_X1 U10301 ( .C1(n9001), .C2(n8872), .A(n8858), .B(n8857), .ZN(
        P2_U3216) );
  XNOR2_X1 U10302 ( .A(n8859), .B(n8862), .ZN(n9009) );
  INV_X1 U10303 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8868) );
  AOI211_X1 U10304 ( .C1(n8862), .C2(n8861), .A(n10080), .B(n8860), .ZN(n8866)
         );
  OAI22_X1 U10305 ( .A1(n8864), .A2(n10074), .B1(n8863), .B2(n10076), .ZN(
        n8865) );
  NOR2_X1 U10306 ( .A1(n8866), .A2(n8865), .ZN(n9002) );
  MUX2_X1 U10307 ( .A(n8868), .B(n9002), .S(n8867), .Z(n8871) );
  AOI22_X1 U10308 ( .A1(n4431), .A2(n10085), .B1(n10087), .B2(n8869), .ZN(
        n8870) );
  OAI211_X1 U10309 ( .C1(n9009), .C2(n8872), .A(n8871), .B(n8870), .ZN(
        P2_U3217) );
  NAND2_X1 U10310 ( .A1(n8933), .A2(n10158), .ZN(n8874) );
  NAND2_X1 U10311 ( .A1(n10156), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n8873) );
  OAI211_X1 U10312 ( .C1(n8932), .C2(n8909), .A(n8874), .B(n8873), .ZN(
        P2_U3490) );
  NAND2_X1 U10313 ( .A1(n10156), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n8875) );
  OAI211_X1 U10314 ( .C1(n8876), .C2(n8909), .A(n8875), .B(n8874), .ZN(
        P2_U3489) );
  INV_X1 U10315 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n8878) );
  MUX2_X1 U10316 ( .A(n8878), .B(n8877), .S(n10158), .Z(n8881) );
  NAND2_X1 U10317 ( .A1(n8879), .A2(n8927), .ZN(n8880) );
  NAND2_X1 U10318 ( .A1(n8881), .A2(n8880), .ZN(P2_U3488) );
  AOI21_X1 U10319 ( .B1(n8927), .B2(n8887), .A(n8886), .ZN(n8888) );
  INV_X1 U10320 ( .A(n8888), .ZN(P2_U3487) );
  INV_X1 U10321 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n8889) );
  MUX2_X1 U10322 ( .A(n8889), .B(n8942), .S(n10158), .Z(n8891) );
  NAND2_X1 U10323 ( .A1(n8944), .A2(n8927), .ZN(n8890) );
  OAI211_X1 U10324 ( .C1(n8947), .C2(n8930), .A(n8891), .B(n8890), .ZN(
        P2_U3486) );
  INV_X1 U10325 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n8892) );
  MUX2_X1 U10326 ( .A(n8892), .B(n8948), .S(n10158), .Z(n8894) );
  NAND2_X1 U10327 ( .A1(n8950), .A2(n8927), .ZN(n8893) );
  OAI211_X1 U10328 ( .C1(n8930), .C2(n8953), .A(n8894), .B(n8893), .ZN(
        P2_U3485) );
  MUX2_X1 U10329 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n8954), .S(n10158), .Z(
        n8896) );
  OAI22_X1 U10330 ( .A1(n8956), .A2(n8930), .B1(n8955), .B2(n8909), .ZN(n8895)
         );
  OR2_X1 U10331 ( .A1(n8896), .A2(n8895), .ZN(P2_U3484) );
  MUX2_X1 U10332 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n8959), .S(n10158), .Z(
        n8900) );
  INV_X1 U10333 ( .A(n8897), .ZN(n8965) );
  OAI22_X1 U10334 ( .A1(n8965), .A2(n8930), .B1(n8898), .B2(n8909), .ZN(n8899)
         );
  OR2_X1 U10335 ( .A1(n8900), .A2(n8899), .ZN(P2_U3483) );
  INV_X1 U10336 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n8903) );
  AOI21_X1 U10337 ( .B1(n10104), .B2(n8902), .A(n8901), .ZN(n8966) );
  MUX2_X1 U10338 ( .A(n8903), .B(n8966), .S(n10158), .Z(n8904) );
  OAI21_X1 U10339 ( .B1(n8970), .B2(n8909), .A(n8904), .ZN(P2_U3482) );
  INV_X1 U10340 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n8905) );
  MUX2_X1 U10341 ( .A(n8905), .B(n8971), .S(n10158), .Z(n8907) );
  NAND2_X1 U10342 ( .A1(n8973), .A2(n8927), .ZN(n8906) );
  OAI211_X1 U10343 ( .C1(n8976), .C2(n8930), .A(n8907), .B(n8906), .ZN(
        P2_U3481) );
  MUX2_X1 U10344 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n8908), .S(n10158), .Z(
        n8912) );
  OAI22_X1 U10345 ( .A1(n8982), .A2(n8930), .B1(n8910), .B2(n8909), .ZN(n8911)
         );
  OR2_X1 U10346 ( .A1(n8912), .A2(n8911), .ZN(P2_U3480) );
  AOI22_X1 U10347 ( .A1(n8914), .A2(n10104), .B1(n10141), .B2(n8913), .ZN(
        n8915) );
  NAND2_X1 U10348 ( .A1(n8916), .A2(n8915), .ZN(n8983) );
  MUX2_X1 U10349 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n8983), .S(n10158), .Z(
        P2_U3479) );
  INV_X1 U10350 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n8917) );
  MUX2_X1 U10351 ( .A(n8917), .B(n8984), .S(n10158), .Z(n8919) );
  NAND2_X1 U10352 ( .A1(n8986), .A2(n8927), .ZN(n8918) );
  OAI211_X1 U10353 ( .C1(n8989), .C2(n8930), .A(n8919), .B(n8918), .ZN(
        P2_U3478) );
  INV_X1 U10354 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8920) );
  MUX2_X1 U10355 ( .A(n8920), .B(n8990), .S(n10158), .Z(n8922) );
  NAND2_X1 U10356 ( .A1(n8992), .A2(n8927), .ZN(n8921) );
  OAI211_X1 U10357 ( .C1(n8930), .C2(n8995), .A(n8922), .B(n8921), .ZN(
        P2_U3477) );
  INV_X1 U10358 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n8923) );
  MUX2_X1 U10359 ( .A(n8923), .B(n8996), .S(n10158), .Z(n8925) );
  NAND2_X1 U10360 ( .A1(n8998), .A2(n8927), .ZN(n8924) );
  OAI211_X1 U10361 ( .C1(n9001), .C2(n8930), .A(n8925), .B(n8924), .ZN(
        P2_U3476) );
  MUX2_X1 U10362 ( .A(n8926), .B(n9002), .S(n10158), .Z(n8929) );
  NAND2_X1 U10363 ( .A1(n4431), .A2(n8927), .ZN(n8928) );
  OAI211_X1 U10364 ( .C1(n9009), .C2(n8930), .A(n8929), .B(n8928), .ZN(
        P2_U3475) );
  MUX2_X1 U10365 ( .A(n8931), .B(P2_REG1_REG_0__SCAN_IN), .S(n10156), .Z(
        P2_U3459) );
  NAND2_X1 U10366 ( .A1(n4523), .A2(n9004), .ZN(n8934) );
  NAND2_X1 U10367 ( .A1(n8933), .A2(n10142), .ZN(n8936) );
  OAI211_X1 U10368 ( .C1(n8413), .C2(n10142), .A(n8934), .B(n8936), .ZN(
        P2_U3458) );
  NAND2_X1 U10369 ( .A1(n8935), .A2(n9004), .ZN(n8937) );
  OAI211_X1 U10370 ( .C1(n8232), .C2(n10142), .A(n8937), .B(n8936), .ZN(
        P2_U3457) );
  INV_X1 U10371 ( .A(n8939), .ZN(n8940) );
  OAI21_X1 U10372 ( .B1(n8941), .B2(n8969), .A(n8940), .ZN(P2_U3455) );
  MUX2_X1 U10373 ( .A(n8943), .B(n8942), .S(n10142), .Z(n8946) );
  NAND2_X1 U10374 ( .A1(n8944), .A2(n9004), .ZN(n8945) );
  OAI211_X1 U10375 ( .C1(n8947), .C2(n9008), .A(n8946), .B(n8945), .ZN(
        P2_U3454) );
  MUX2_X1 U10376 ( .A(n8949), .B(n8948), .S(n10142), .Z(n8952) );
  NAND2_X1 U10377 ( .A1(n8950), .A2(n9004), .ZN(n8951) );
  OAI211_X1 U10378 ( .C1(n8953), .C2(n9008), .A(n8952), .B(n8951), .ZN(
        P2_U3453) );
  MUX2_X1 U10379 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n8954), .S(n10142), .Z(
        n8958) );
  OAI22_X1 U10380 ( .A1(n8956), .A2(n9008), .B1(n8955), .B2(n8969), .ZN(n8957)
         );
  OR2_X1 U10381 ( .A1(n8958), .A2(n8957), .ZN(P2_U3452) );
  INV_X1 U10382 ( .A(n8959), .ZN(n8960) );
  MUX2_X1 U10383 ( .A(n8961), .B(n8960), .S(n10142), .Z(n8964) );
  NAND2_X1 U10384 ( .A1(n8962), .A2(n9004), .ZN(n8963) );
  OAI211_X1 U10385 ( .C1(n8965), .C2(n9008), .A(n8964), .B(n8963), .ZN(
        P2_U3451) );
  MUX2_X1 U10386 ( .A(n8967), .B(n8966), .S(n10142), .Z(n8968) );
  OAI21_X1 U10387 ( .B1(n8970), .B2(n8969), .A(n8968), .ZN(P2_U3450) );
  MUX2_X1 U10388 ( .A(n8972), .B(n8971), .S(n10142), .Z(n8975) );
  NAND2_X1 U10389 ( .A1(n8973), .A2(n9004), .ZN(n8974) );
  OAI211_X1 U10390 ( .C1(n8976), .C2(n9008), .A(n8975), .B(n8974), .ZN(
        P2_U3449) );
  MUX2_X1 U10391 ( .A(n8978), .B(n8977), .S(n10142), .Z(n8981) );
  NAND2_X1 U10392 ( .A1(n8979), .A2(n9004), .ZN(n8980) );
  OAI211_X1 U10393 ( .C1(n8982), .C2(n9008), .A(n8981), .B(n8980), .ZN(
        P2_U3448) );
  MUX2_X1 U10394 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n8983), .S(n10142), .Z(
        P2_U3447) );
  MUX2_X1 U10395 ( .A(n8985), .B(n8984), .S(n10142), .Z(n8988) );
  NAND2_X1 U10396 ( .A1(n8986), .A2(n9004), .ZN(n8987) );
  OAI211_X1 U10397 ( .C1(n8989), .C2(n9008), .A(n8988), .B(n8987), .ZN(
        P2_U3446) );
  INV_X1 U10398 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n8991) );
  MUX2_X1 U10399 ( .A(n8991), .B(n8990), .S(n10142), .Z(n8994) );
  NAND2_X1 U10400 ( .A1(n8992), .A2(n9004), .ZN(n8993) );
  OAI211_X1 U10401 ( .C1(n8995), .C2(n9008), .A(n8994), .B(n8993), .ZN(
        P2_U3444) );
  INV_X1 U10402 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n8997) );
  MUX2_X1 U10403 ( .A(n8997), .B(n8996), .S(n10142), .Z(n9000) );
  NAND2_X1 U10404 ( .A1(n8998), .A2(n9004), .ZN(n8999) );
  OAI211_X1 U10405 ( .C1(n9001), .C2(n9008), .A(n9000), .B(n8999), .ZN(
        P2_U3441) );
  INV_X1 U10406 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n9003) );
  MUX2_X1 U10407 ( .A(n9003), .B(n9002), .S(n10142), .Z(n9007) );
  NAND2_X1 U10408 ( .A1(n4431), .A2(n9004), .ZN(n9006) );
  OAI211_X1 U10409 ( .C1(n9009), .C2(n9008), .A(n9007), .B(n9006), .ZN(
        P2_U3438) );
  INV_X1 U10410 ( .A(n8401), .ZN(n9798) );
  INV_X1 U10411 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n9010) );
  NAND3_X1 U10412 ( .A1(n9010), .A2(P2_STATE_REG_SCAN_IN), .A3(
        P2_IR_REG_31__SCAN_IN), .ZN(n9012) );
  OAI22_X1 U10413 ( .A1(n5869), .A2(n9012), .B1(n9011), .B2(n9015), .ZN(n9013)
         );
  INV_X1 U10414 ( .A(n9013), .ZN(n9014) );
  OAI21_X1 U10415 ( .B1(n9798), .B2(n9022), .A(n9014), .ZN(P2_U3264) );
  OAI222_X1 U10416 ( .A1(P2_U3151), .A2(n9018), .B1(n9022), .B2(n9017), .C1(
        n9016), .C2(n9015), .ZN(P2_U3266) );
  AOI21_X1 U10417 ( .B1(n9020), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n9019), .ZN(
        n9021) );
  OAI21_X1 U10418 ( .B1(n9023), .B2(n9022), .A(n9021), .ZN(P2_U3267) );
  INV_X1 U10419 ( .A(n9024), .ZN(n9025) );
  MUX2_X1 U10420 ( .A(n9025), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  OAI22_X1 U10421 ( .A1(n9458), .A2(n6864), .B1(n9447), .B2(n9113), .ZN(n9037)
         );
  NAND2_X1 U10422 ( .A1(n9762), .A2(n9044), .ZN(n9029) );
  NAND2_X1 U10423 ( .A1(n9665), .A2(n9049), .ZN(n9028) );
  NAND2_X1 U10424 ( .A1(n9029), .A2(n9028), .ZN(n9031) );
  XNOR2_X1 U10425 ( .A(n9031), .B(n9030), .ZN(n9036) );
  XOR2_X1 U10426 ( .A(n9037), .B(n9036), .Z(n9140) );
  OAI22_X1 U10427 ( .A1(n9669), .A2(n4406), .B1(n9657), .B2(n6864), .ZN(n9032)
         );
  XNOR2_X1 U10428 ( .A(n9032), .B(n9111), .ZN(n9041) );
  OR2_X1 U10429 ( .A1(n9669), .A2(n6864), .ZN(n9035) );
  INV_X1 U10430 ( .A(n9657), .ZN(n9262) );
  NAND2_X1 U10431 ( .A1(n9262), .A2(n9033), .ZN(n9034) );
  NAND2_X1 U10432 ( .A1(n9035), .A2(n9034), .ZN(n9042) );
  XNOR2_X1 U10433 ( .A(n9041), .B(n9042), .ZN(n9238) );
  INV_X1 U10434 ( .A(n9036), .ZN(n9039) );
  INV_X1 U10435 ( .A(n9037), .ZN(n9038) );
  NAND2_X1 U10436 ( .A1(n9039), .A2(n9038), .ZN(n9235) );
  INV_X1 U10437 ( .A(n9041), .ZN(n9043) );
  NAND2_X1 U10438 ( .A1(n9043), .A2(n9042), .ZN(n9055) );
  NAND2_X1 U10439 ( .A1(n9661), .A2(n9044), .ZN(n9046) );
  NAND2_X1 U10440 ( .A1(n9666), .A2(n9049), .ZN(n9045) );
  NAND2_X1 U10441 ( .A1(n9046), .A2(n9045), .ZN(n9047) );
  XNOR2_X1 U10442 ( .A(n9047), .B(n9111), .ZN(n9051) );
  INV_X1 U10443 ( .A(n9051), .ZN(n9053) );
  NOR2_X1 U10444 ( .A1(n9242), .A2(n9113), .ZN(n9048) );
  AOI21_X1 U10445 ( .B1(n9661), .B2(n9049), .A(n9048), .ZN(n9050) );
  INV_X1 U10446 ( .A(n9050), .ZN(n9052) );
  AOI21_X1 U10447 ( .B1(n9053), .B2(n9052), .A(n9121), .ZN(n9054) );
  AOI21_X1 U10448 ( .B1(n9236), .B2(n9055), .A(n9054), .ZN(n9059) );
  INV_X1 U10449 ( .A(n9054), .ZN(n9057) );
  INV_X1 U10450 ( .A(n9055), .ZN(n9056) );
  NOR2_X1 U10451 ( .A1(n9057), .A2(n9056), .ZN(n9058) );
  OAI21_X1 U10452 ( .B1(n9059), .B2(n9116), .A(n9237), .ZN(n9065) );
  OAI22_X1 U10453 ( .A1(n9657), .A2(n9255), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9060), .ZN(n9062) );
  NOR2_X1 U10454 ( .A1(n9658), .A2(n9241), .ZN(n9061) );
  AOI211_X1 U10455 ( .C1(n9431), .C2(n9252), .A(n9062), .B(n9061), .ZN(n9064)
         );
  NAND2_X1 U10456 ( .A1(n9661), .A2(n9257), .ZN(n9063) );
  NAND3_X1 U10457 ( .A1(n9065), .A2(n9064), .A3(n9063), .ZN(P1_U3214) );
  XNOR2_X1 U10458 ( .A(n9067), .B(n9066), .ZN(n9068) );
  XNOR2_X1 U10459 ( .A(n9069), .B(n9068), .ZN(n9075) );
  NAND2_X1 U10460 ( .A1(P1_U3086), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n9853) );
  INV_X1 U10461 ( .A(n9853), .ZN(n9070) );
  AOI21_X1 U10462 ( .B1(n9228), .B2(n9881), .A(n9070), .ZN(n9072) );
  NAND2_X1 U10463 ( .A1(n9252), .A2(n9628), .ZN(n9071) );
  OAI211_X1 U10464 ( .C1(n9736), .C2(n9241), .A(n9072), .B(n9071), .ZN(n9073)
         );
  AOI21_X1 U10465 ( .B1(n9749), .B2(n9257), .A(n9073), .ZN(n9074) );
  OAI21_X1 U10466 ( .B1(n9075), .B2(n9259), .A(n9074), .ZN(P1_U3215) );
  INV_X1 U10467 ( .A(n9684), .ZN(n9489) );
  INV_X1 U10468 ( .A(n9076), .ZN(n9078) );
  NOR3_X1 U10469 ( .A1(n4332), .A2(n9078), .A3(n9077), .ZN(n9080) );
  OAI21_X1 U10470 ( .B1(n9080), .B2(n9079), .A(n9237), .ZN(n9085) );
  INV_X1 U10471 ( .A(n9081), .ZN(n9483) );
  AOI22_X1 U10472 ( .A1(n9486), .A2(n9251), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        P1_U3086), .ZN(n9082) );
  OAI21_X1 U10473 ( .B1(n9680), .B2(n9255), .A(n9082), .ZN(n9083) );
  AOI21_X1 U10474 ( .B1(n9483), .B2(n9252), .A(n9083), .ZN(n9084) );
  OAI211_X1 U10475 ( .C1(n9489), .C2(n9247), .A(n9085), .B(n9084), .ZN(
        P1_U3216) );
  XNOR2_X1 U10476 ( .A(n9086), .B(n9209), .ZN(n9087) );
  NAND2_X1 U10477 ( .A1(n9087), .A2(n9088), .ZN(n9210) );
  OAI21_X1 U10478 ( .B1(n9088), .B2(n9087), .A(n9210), .ZN(n9089) );
  NAND2_X1 U10479 ( .A1(n9089), .A2(n9237), .ZN(n9100) );
  NOR2_X1 U10480 ( .A1(n9090), .A2(n9247), .ZN(n9098) );
  AND2_X1 U10481 ( .A1(n9252), .A2(n9091), .ZN(n9097) );
  NOR2_X1 U10482 ( .A1(n9255), .A2(n9092), .ZN(n9096) );
  OAI22_X1 U10483 ( .A1(n9241), .A2(n9094), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9093), .ZN(n9095) );
  NOR4_X1 U10484 ( .A1(n9098), .A2(n9097), .A3(n9096), .A4(n9095), .ZN(n9099)
         );
  NAND2_X1 U10485 ( .A1(n9100), .A2(n9099), .ZN(P1_U3217) );
  XNOR2_X1 U10486 ( .A(n9102), .B(n9101), .ZN(n9103) );
  XNOR2_X1 U10487 ( .A(n9104), .B(n9103), .ZN(n9110) );
  NOR2_X1 U10488 ( .A1(n9105), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9374) );
  AOI21_X1 U10489 ( .B1(n9251), .B2(n9545), .A(n9374), .ZN(n9107) );
  NAND2_X1 U10490 ( .A1(n9252), .A2(n9542), .ZN(n9106) );
  OAI211_X1 U10491 ( .C1(n9708), .C2(n9255), .A(n9107), .B(n9106), .ZN(n9108)
         );
  AOI21_X1 U10492 ( .B1(n9541), .B2(n9257), .A(n9108), .ZN(n9109) );
  OAI21_X1 U10493 ( .B1(n9110), .B2(n9259), .A(n9109), .ZN(P1_U3219) );
  OAI22_X1 U10494 ( .A1(n9651), .A2(n4406), .B1(n9658), .B2(n6864), .ZN(n9112)
         );
  XNOR2_X1 U10495 ( .A(n9112), .B(n9111), .ZN(n9115) );
  OAI22_X1 U10496 ( .A1(n9651), .A2(n6864), .B1(n9658), .B2(n9113), .ZN(n9114)
         );
  XNOR2_X1 U10497 ( .A(n9115), .B(n9114), .ZN(n9122) );
  NAND3_X1 U10498 ( .A1(n9116), .A2(n9237), .A3(n9122), .ZN(n9125) );
  OAI22_X1 U10499 ( .A1(n9261), .A2(n9241), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9117), .ZN(n9118) );
  AOI21_X1 U10500 ( .B1(n9228), .B2(n9666), .A(n9118), .ZN(n9119) );
  OAI21_X1 U10501 ( .B1(n9205), .B2(n9419), .A(n9119), .ZN(n9120) );
  AOI21_X1 U10502 ( .B1(n9401), .B2(n9257), .A(n9120), .ZN(n9124) );
  NAND3_X1 U10503 ( .A1(n9122), .A2(n9237), .A3(n9121), .ZN(n9123) );
  NAND4_X1 U10504 ( .A1(n9126), .A2(n9125), .A3(n9124), .A4(n9123), .ZN(
        P1_U3220) );
  OR2_X1 U10505 ( .A1(n9127), .A2(n9185), .ZN(n9183) );
  NAND2_X1 U10506 ( .A1(n9183), .A2(n9128), .ZN(n9130) );
  OAI21_X1 U10507 ( .B1(n9131), .B2(n9130), .A(n9129), .ZN(n9132) );
  NAND2_X1 U10508 ( .A1(n9132), .A2(n9237), .ZN(n9137) );
  NOR2_X1 U10509 ( .A1(n9241), .A2(n9680), .ZN(n9135) );
  OAI22_X1 U10510 ( .A1(n9255), .A2(n9709), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9133), .ZN(n9134) );
  AOI211_X1 U10511 ( .C1(n9515), .C2(n9252), .A(n9135), .B(n9134), .ZN(n9136)
         );
  OAI211_X1 U10512 ( .C1(n9770), .C2(n9247), .A(n9137), .B(n9136), .ZN(
        P1_U3223) );
  OAI21_X1 U10513 ( .B1(n9140), .B2(n9139), .A(n9138), .ZN(n9141) );
  NAND2_X1 U10514 ( .A1(n9141), .A2(n9237), .ZN(n9146) );
  INV_X1 U10515 ( .A(n9455), .ZN(n9144) );
  AOI22_X1 U10516 ( .A1(n9262), .A2(n9251), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3086), .ZN(n9142) );
  OAI21_X1 U10517 ( .B1(n9681), .B2(n9255), .A(n9142), .ZN(n9143) );
  AOI21_X1 U10518 ( .B1(n9144), .B2(n9252), .A(n9143), .ZN(n9145) );
  OAI211_X1 U10519 ( .C1(n9458), .C2(n9247), .A(n9146), .B(n9145), .ZN(
        P1_U3225) );
  XNOR2_X1 U10520 ( .A(n9147), .B(n9148), .ZN(n9250) );
  NOR2_X1 U10521 ( .A1(n9250), .A2(n9249), .ZN(n9248) );
  AOI21_X1 U10522 ( .B1(n9148), .B2(n9147), .A(n9248), .ZN(n9152) );
  XNOR2_X1 U10523 ( .A(n9150), .B(n9149), .ZN(n9151) );
  XNOR2_X1 U10524 ( .A(n9152), .B(n9151), .ZN(n9158) );
  NAND2_X1 U10525 ( .A1(n9228), .A2(n9263), .ZN(n9154) );
  OAI211_X1 U10526 ( .C1(n9556), .C2(n9241), .A(n9154), .B(n9153), .ZN(n9156)
         );
  NOR2_X1 U10527 ( .A1(n4603), .A2(n9247), .ZN(n9155) );
  AOI211_X1 U10528 ( .C1(n9584), .C2(n9252), .A(n9156), .B(n9155), .ZN(n9157)
         );
  OAI21_X1 U10529 ( .B1(n9158), .B2(n9259), .A(n9157), .ZN(P1_U3226) );
  OAI211_X1 U10530 ( .C1(n9161), .C2(n9160), .A(n9159), .B(n9237), .ZN(n9166)
         );
  AOI21_X1 U10531 ( .B1(n9251), .B2(n9727), .A(n9162), .ZN(n9163) );
  OAI21_X1 U10532 ( .B1(n9571), .B2(n9255), .A(n9163), .ZN(n9164) );
  AOI21_X1 U10533 ( .B1(n9567), .B2(n9252), .A(n9164), .ZN(n9165) );
  OAI211_X1 U10534 ( .C1(n9783), .C2(n9247), .A(n9166), .B(n9165), .ZN(
        P1_U3228) );
  OAI21_X1 U10535 ( .B1(n9169), .B2(n9168), .A(n9167), .ZN(n9173) );
  XNOR2_X1 U10536 ( .A(n9171), .B(n9170), .ZN(n9172) );
  XNOR2_X1 U10537 ( .A(n9173), .B(n9172), .ZN(n9182) );
  OR2_X1 U10538 ( .A1(n9255), .A2(n9174), .ZN(n9177) );
  INV_X1 U10539 ( .A(n9175), .ZN(n9176) );
  OAI211_X1 U10540 ( .C1(n9241), .C2(n9219), .A(n9177), .B(n9176), .ZN(n9179)
         );
  NOR2_X1 U10541 ( .A1(n9940), .A2(n9247), .ZN(n9178) );
  AOI211_X1 U10542 ( .C1(n9180), .C2(n9252), .A(n9179), .B(n9178), .ZN(n9181)
         );
  OAI21_X1 U10543 ( .B1(n9182), .B2(n9259), .A(n9181), .ZN(P1_U3231) );
  INV_X1 U10544 ( .A(n9183), .ZN(n9184) );
  AOI21_X1 U10545 ( .B1(n9185), .B2(n9127), .A(n9184), .ZN(n9191) );
  OAI22_X1 U10546 ( .A1(n9241), .A2(n9531), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9186), .ZN(n9187) );
  AOI21_X1 U10547 ( .B1(n9228), .B2(n9718), .A(n9187), .ZN(n9188) );
  OAI21_X1 U10548 ( .B1(n9205), .B2(n9533), .A(n9188), .ZN(n9189) );
  AOI21_X1 U10549 ( .B1(n9705), .B2(n9257), .A(n9189), .ZN(n9190) );
  OAI21_X1 U10550 ( .B1(n9191), .B2(n9259), .A(n9190), .ZN(P1_U3233) );
  XOR2_X1 U10551 ( .A(n9193), .B(n9192), .Z(n9199) );
  AOI22_X1 U10552 ( .A1(n9251), .A2(n9601), .B1(P1_REG3_REG_13__SCAN_IN), .B2(
        P1_U3086), .ZN(n9196) );
  NAND2_X1 U10553 ( .A1(n9252), .A2(n9194), .ZN(n9195) );
  OAI211_X1 U10554 ( .C1(n9953), .C2(n9255), .A(n9196), .B(n9195), .ZN(n9197)
         );
  AOI21_X1 U10555 ( .B1(n9958), .B2(n9257), .A(n9197), .ZN(n9198) );
  OAI21_X1 U10556 ( .B1(n9199), .B2(n9259), .A(n9198), .ZN(P1_U3234) );
  AOI21_X1 U10557 ( .B1(n9201), .B2(n9200), .A(n4332), .ZN(n9208) );
  OAI22_X1 U10558 ( .A1(n9255), .A2(n9531), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9202), .ZN(n9203) );
  AOI21_X1 U10559 ( .B1(n9251), .B2(n9690), .A(n9203), .ZN(n9204) );
  OAI21_X1 U10560 ( .B1(n9205), .B2(n9495), .A(n9204), .ZN(n9206) );
  AOI21_X1 U10561 ( .B1(n9499), .B2(n9257), .A(n9206), .ZN(n9207) );
  OAI21_X1 U10562 ( .B1(n9208), .B2(n9259), .A(n9207), .ZN(P1_U3235) );
  INV_X1 U10563 ( .A(n9209), .ZN(n9211) );
  OAI21_X1 U10564 ( .B1(n9211), .B2(n9086), .A(n9210), .ZN(n9215) );
  XNOR2_X1 U10565 ( .A(n9213), .B(n9212), .ZN(n9214) );
  XNOR2_X1 U10566 ( .A(n9215), .B(n9214), .ZN(n9223) );
  AOI22_X1 U10567 ( .A1(n9251), .A2(n9264), .B1(P1_REG3_REG_11__SCAN_IN), .B2(
        P1_U3086), .ZN(n9218) );
  NAND2_X1 U10568 ( .A1(n9252), .A2(n9216), .ZN(n9217) );
  OAI211_X1 U10569 ( .C1(n9219), .C2(n9255), .A(n9218), .B(n9217), .ZN(n9220)
         );
  AOI21_X1 U10570 ( .B1(n9221), .B2(n9257), .A(n9220), .ZN(n9222) );
  OAI21_X1 U10571 ( .B1(n9223), .B2(n9259), .A(n9222), .ZN(P1_U3236) );
  NAND2_X1 U10572 ( .A1(n9225), .A2(n9224), .ZN(n9227) );
  XNOR2_X1 U10573 ( .A(n9227), .B(n9226), .ZN(n9234) );
  NAND2_X1 U10574 ( .A1(n9228), .A2(n9719), .ZN(n9230) );
  NAND2_X1 U10575 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9355) );
  OAI211_X1 U10576 ( .C1(n9530), .C2(n9241), .A(n9230), .B(n9355), .ZN(n9232)
         );
  NOR2_X1 U10577 ( .A1(n9779), .A2(n9247), .ZN(n9231) );
  AOI211_X1 U10578 ( .C1(n9553), .C2(n9252), .A(n9232), .B(n9231), .ZN(n9233)
         );
  OAI21_X1 U10579 ( .B1(n9234), .B2(n9259), .A(n9233), .ZN(P1_U3238) );
  AND2_X1 U10580 ( .A1(n9138), .A2(n9235), .ZN(n9239) );
  OAI211_X1 U10581 ( .C1(n9239), .C2(n9238), .A(n9237), .B(n9236), .ZN(n9246)
         );
  OAI22_X1 U10582 ( .A1(n9447), .A2(n9255), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9240), .ZN(n9244) );
  NOR2_X1 U10583 ( .A1(n9242), .A2(n9241), .ZN(n9243) );
  AOI211_X1 U10584 ( .C1(n9445), .C2(n9252), .A(n9244), .B(n9243), .ZN(n9245)
         );
  OAI211_X1 U10585 ( .C1(n9669), .C2(n9247), .A(n9246), .B(n9245), .ZN(
        P1_U3240) );
  AOI21_X1 U10586 ( .B1(n9250), .B2(n9249), .A(n9248), .ZN(n9260) );
  INV_X1 U10587 ( .A(n9571), .ZN(n9728) );
  AOI22_X1 U10588 ( .A1(n9251), .A2(n9728), .B1(P1_REG3_REG_15__SCAN_IN), .B2(
        P1_U3086), .ZN(n9254) );
  NAND2_X1 U10589 ( .A1(n9252), .A2(n9607), .ZN(n9253) );
  OAI211_X1 U10590 ( .C1(n9955), .C2(n9255), .A(n9254), .B(n9253), .ZN(n9256)
         );
  AOI21_X1 U10591 ( .B1(n9606), .B2(n9257), .A(n9256), .ZN(n9258) );
  OAI21_X1 U10592 ( .B1(n9260), .B2(n9259), .A(n9258), .ZN(P1_U3241) );
  INV_X1 U10593 ( .A(n9261), .ZN(n9648) );
  MUX2_X1 U10594 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n9648), .S(P1_U3973), .Z(
        P1_U3583) );
  MUX2_X1 U10595 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9434), .S(P1_U3973), .Z(
        P1_U3582) );
  MUX2_X1 U10596 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9666), .S(P1_U3973), .Z(
        P1_U3581) );
  MUX2_X1 U10597 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9262), .S(P1_U3973), .Z(
        P1_U3580) );
  MUX2_X1 U10598 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9665), .S(P1_U3973), .Z(
        P1_U3579) );
  MUX2_X1 U10599 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9486), .S(P1_U3973), .Z(
        P1_U3578) );
  MUX2_X1 U10600 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9690), .S(P1_U3973), .Z(
        P1_U3577) );
  INV_X1 U10601 ( .A(n9531), .ZN(n9689) );
  MUX2_X1 U10602 ( .A(n9689), .B(P1_DATAO_REG_21__SCAN_IN), .S(n9273), .Z(
        P1_U3575) );
  MUX2_X1 U10603 ( .A(n9545), .B(P1_DATAO_REG_20__SCAN_IN), .S(n9273), .Z(
        P1_U3574) );
  MUX2_X1 U10604 ( .A(n9718), .B(P1_DATAO_REG_19__SCAN_IN), .S(n9273), .Z(
        P1_U3573) );
  MUX2_X1 U10605 ( .A(n9727), .B(P1_DATAO_REG_18__SCAN_IN), .S(n9273), .Z(
        P1_U3572) );
  MUX2_X1 U10606 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9719), .S(P1_U3973), .Z(
        P1_U3571) );
  MUX2_X1 U10607 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9728), .S(P1_U3973), .Z(
        P1_U3570) );
  MUX2_X1 U10608 ( .A(n9263), .B(P1_DATAO_REG_15__SCAN_IN), .S(n9273), .Z(
        P1_U3569) );
  MUX2_X1 U10609 ( .A(n9601), .B(P1_DATAO_REG_14__SCAN_IN), .S(n9273), .Z(
        P1_U3568) );
  MUX2_X1 U10610 ( .A(n9881), .B(P1_DATAO_REG_13__SCAN_IN), .S(n9273), .Z(
        P1_U3567) );
  MUX2_X1 U10611 ( .A(n9264), .B(P1_DATAO_REG_12__SCAN_IN), .S(n9273), .Z(
        P1_U3566) );
  MUX2_X1 U10612 ( .A(n9878), .B(P1_DATAO_REG_11__SCAN_IN), .S(n9273), .Z(
        P1_U3565) );
  MUX2_X1 U10613 ( .A(n9265), .B(P1_DATAO_REG_10__SCAN_IN), .S(n9273), .Z(
        P1_U3564) );
  MUX2_X1 U10614 ( .A(n9266), .B(P1_DATAO_REG_9__SCAN_IN), .S(n9273), .Z(
        P1_U3563) );
  MUX2_X1 U10615 ( .A(n9267), .B(P1_DATAO_REG_8__SCAN_IN), .S(n9273), .Z(
        P1_U3562) );
  MUX2_X1 U10616 ( .A(n9268), .B(P1_DATAO_REG_7__SCAN_IN), .S(n9273), .Z(
        P1_U3561) );
  MUX2_X1 U10617 ( .A(n9269), .B(P1_DATAO_REG_6__SCAN_IN), .S(n9273), .Z(
        P1_U3560) );
  MUX2_X1 U10618 ( .A(n9270), .B(P1_DATAO_REG_5__SCAN_IN), .S(n9273), .Z(
        P1_U3559) );
  MUX2_X1 U10619 ( .A(n9271), .B(P1_DATAO_REG_4__SCAN_IN), .S(n9273), .Z(
        P1_U3558) );
  MUX2_X1 U10620 ( .A(n9272), .B(P1_DATAO_REG_3__SCAN_IN), .S(n9273), .Z(
        P1_U3557) );
  MUX2_X1 U10621 ( .A(n7225), .B(P1_DATAO_REG_2__SCAN_IN), .S(n9273), .Z(
        P1_U3556) );
  MUX2_X1 U10622 ( .A(n9274), .B(P1_DATAO_REG_1__SCAN_IN), .S(n9273), .Z(
        P1_U3555) );
  NAND2_X1 U10623 ( .A1(n9799), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n9277) );
  AOI211_X1 U10624 ( .C1(n9277), .C2(n9276), .A(n9275), .B(n9857), .ZN(n9278)
         );
  INV_X1 U10625 ( .A(n9278), .ZN(n9287) );
  OAI22_X1 U10626 ( .A1(n9872), .A2(n7529), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9279), .ZN(n9280) );
  AOI21_X1 U10627 ( .B1(n9281), .B2(n9868), .A(n9280), .ZN(n9286) );
  OAI211_X1 U10628 ( .C1(n9284), .C2(n9283), .A(n9842), .B(n9282), .ZN(n9285)
         );
  NAND3_X1 U10629 ( .A1(n9287), .A2(n9286), .A3(n9285), .ZN(P1_U3244) );
  AOI211_X1 U10630 ( .C1(n9290), .C2(n9289), .A(n9288), .B(n9857), .ZN(n9291)
         );
  INV_X1 U10631 ( .A(n9291), .ZN(n9301) );
  INV_X1 U10632 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n9293) );
  OAI21_X1 U10633 ( .B1(n9872), .B2(n9293), .A(n9292), .ZN(n9294) );
  AOI21_X1 U10634 ( .B1(n9295), .B2(n9868), .A(n9294), .ZN(n9300) );
  OAI211_X1 U10635 ( .C1(n9298), .C2(n9297), .A(n9842), .B(n9296), .ZN(n9299)
         );
  NAND3_X1 U10636 ( .A1(n9301), .A2(n9300), .A3(n9299), .ZN(P1_U3246) );
  AOI211_X1 U10637 ( .C1(n9304), .C2(n9303), .A(n9857), .B(n9302), .ZN(n9305)
         );
  INV_X1 U10638 ( .A(n9305), .ZN(n9315) );
  INV_X1 U10639 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n9307) );
  OAI21_X1 U10640 ( .B1(n9872), .B2(n9307), .A(n9306), .ZN(n9308) );
  AOI21_X1 U10641 ( .B1(n9309), .B2(n9868), .A(n9308), .ZN(n9314) );
  OAI211_X1 U10642 ( .C1(n9312), .C2(n9311), .A(n9842), .B(n9310), .ZN(n9313)
         );
  NAND3_X1 U10643 ( .A1(n9315), .A2(n9314), .A3(n9313), .ZN(P1_U3248) );
  AOI211_X1 U10644 ( .C1(n9318), .C2(n9317), .A(n9857), .B(n9316), .ZN(n9319)
         );
  INV_X1 U10645 ( .A(n9319), .ZN(n9329) );
  OAI21_X1 U10646 ( .B1(n9872), .B2(n9321), .A(n9320), .ZN(n9322) );
  AOI21_X1 U10647 ( .B1(n9323), .B2(n9868), .A(n9322), .ZN(n9328) );
  OAI211_X1 U10648 ( .C1(n9326), .C2(n9325), .A(n9842), .B(n9324), .ZN(n9327)
         );
  NAND3_X1 U10649 ( .A1(n9329), .A2(n9328), .A3(n9327), .ZN(P1_U3249) );
  AOI211_X1 U10650 ( .C1(n4342), .C2(n9331), .A(n9857), .B(n9330), .ZN(n9332)
         );
  INV_X1 U10651 ( .A(n9332), .ZN(n9342) );
  OAI21_X1 U10652 ( .B1(n9872), .B2(n9334), .A(n9333), .ZN(n9335) );
  AOI21_X1 U10653 ( .B1(n9336), .B2(n9868), .A(n9335), .ZN(n9341) );
  OAI211_X1 U10654 ( .C1(n9339), .C2(n9338), .A(n9842), .B(n9337), .ZN(n9340)
         );
  NAND3_X1 U10655 ( .A1(n9342), .A2(n9341), .A3(n9340), .ZN(P1_U3250) );
  AOI22_X1 U10656 ( .A1(n9345), .A2(n9344), .B1(n9734), .B2(n9343), .ZN(n9348)
         );
  INV_X1 U10657 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9725) );
  AND2_X1 U10658 ( .A1(n9358), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n9362) );
  AOI21_X1 U10659 ( .B1(n9725), .B2(n9346), .A(n9362), .ZN(n9347) );
  NAND2_X1 U10660 ( .A1(n9348), .A2(n9347), .ZN(n9364) );
  OAI211_X1 U10661 ( .C1(n9348), .C2(n9347), .A(n9364), .B(n9847), .ZN(n9361)
         );
  OR2_X1 U10662 ( .A1(n9349), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n9350) );
  AND2_X1 U10663 ( .A1(n9351), .A2(n9350), .ZN(n9354) );
  NAND2_X1 U10664 ( .A1(n9358), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9366) );
  OR2_X1 U10665 ( .A1(n9358), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9352) );
  AND2_X1 U10666 ( .A1(n9366), .A2(n9352), .ZN(n9353) );
  NAND2_X1 U10667 ( .A1(n9354), .A2(n9353), .ZN(n9367) );
  OAI211_X1 U10668 ( .C1(n9354), .C2(n9353), .A(n9367), .B(n9842), .ZN(n9360)
         );
  INV_X1 U10669 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n9356) );
  OAI21_X1 U10670 ( .B1(n9872), .B2(n9356), .A(n9355), .ZN(n9357) );
  AOI21_X1 U10671 ( .B1(n9358), .B2(n9868), .A(n9357), .ZN(n9359) );
  NAND3_X1 U10672 ( .A1(n9361), .A2(n9360), .A3(n9359), .ZN(P1_U3261) );
  INV_X1 U10673 ( .A(n9362), .ZN(n9363) );
  NAND2_X1 U10674 ( .A1(n9364), .A2(n9363), .ZN(n9365) );
  XNOR2_X1 U10675 ( .A(n9365), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n9372) );
  INV_X1 U10676 ( .A(n9372), .ZN(n9370) );
  NAND2_X1 U10677 ( .A1(n9367), .A2(n9366), .ZN(n9368) );
  XNOR2_X1 U10678 ( .A(n9368), .B(P1_REG2_REG_19__SCAN_IN), .ZN(n9371) );
  NAND2_X1 U10679 ( .A1(n9371), .A2(n9842), .ZN(n9369) );
  NOR2_X1 U10680 ( .A1(n4315), .A2(n9637), .ZN(n9380) );
  NOR2_X1 U10681 ( .A1(n9755), .A2(n9630), .ZN(n9377) );
  AOI211_X1 U10682 ( .C1(n4315), .C2(P1_REG2_REG_31__SCAN_IN), .A(n9380), .B(
        n9377), .ZN(n9378) );
  OAI21_X1 U10683 ( .B1(n9638), .B2(n9904), .A(n9378), .ZN(P1_U3263) );
  AND2_X1 U10684 ( .A1(n4315), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n9379) );
  NOR2_X1 U10685 ( .A1(n9380), .A2(n9379), .ZN(n9383) );
  NAND2_X1 U10686 ( .A1(n9381), .A2(n9901), .ZN(n9382) );
  OAI211_X1 U10687 ( .C1(n9384), .C2(n9904), .A(n9383), .B(n9382), .ZN(
        P1_U3264) );
  NAND2_X1 U10688 ( .A1(n9386), .A2(n9385), .ZN(n9461) );
  NAND2_X1 U10689 ( .A1(n9442), .A2(n9441), .ZN(n9440) );
  INV_X1 U10690 ( .A(n9644), .ZN(n9413) );
  NOR2_X1 U10691 ( .A1(n9473), .A2(n9681), .ZN(n9394) );
  NAND2_X1 U10692 ( .A1(n9473), .A2(n9681), .ZN(n9396) );
  NAND2_X1 U10693 ( .A1(n9397), .A2(n9396), .ZN(n9453) );
  NOR2_X1 U10694 ( .A1(n9762), .A2(n9665), .ZN(n9398) );
  NOR2_X1 U10695 ( .A1(n9669), .A2(n9657), .ZN(n9400) );
  NAND2_X1 U10696 ( .A1(n9669), .A2(n9657), .ZN(n9399) );
  NAND2_X1 U10697 ( .A1(n9651), .A2(n9658), .ZN(n9402) );
  XNOR2_X1 U10698 ( .A(n9404), .B(n9403), .ZN(n9641) );
  NAND2_X1 U10699 ( .A1(n9641), .A2(n9907), .ZN(n9412) );
  AOI211_X1 U10700 ( .C1(n6333), .C2(n9417), .A(n9889), .B(n9405), .ZN(n9645)
         );
  INV_X1 U10701 ( .A(n6333), .ZN(n9642) );
  OAI22_X1 U10702 ( .A1(n9407), .A2(n9532), .B1(n9406), .B2(n9611), .ZN(n9408)
         );
  AOI21_X1 U10703 ( .B1(n9434), .B2(n9421), .A(n9408), .ZN(n9409) );
  OAI21_X1 U10704 ( .B1(n9642), .B2(n9630), .A(n9409), .ZN(n9410) );
  AOI21_X1 U10705 ( .B1(n9645), .B2(n9635), .A(n9410), .ZN(n9411) );
  OAI211_X1 U10706 ( .C1(n9413), .C2(n4315), .A(n9412), .B(n9411), .ZN(
        P1_U3356) );
  XNOR2_X1 U10707 ( .A(n9414), .B(n9415), .ZN(n9655) );
  XNOR2_X1 U10708 ( .A(n9416), .B(n9415), .ZN(n9653) );
  OAI211_X1 U10709 ( .C1(n9651), .C2(n9430), .A(n9573), .B(n9417), .ZN(n9650)
         );
  NOR2_X1 U10710 ( .A1(n9650), .A2(n9904), .ZN(n9425) );
  INV_X1 U10711 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n9418) );
  OAI22_X1 U10712 ( .A1(n9419), .A2(n9532), .B1(n9418), .B2(n9611), .ZN(n9420)
         );
  AOI21_X1 U10713 ( .B1(n9648), .B2(n9568), .A(n9420), .ZN(n9423) );
  NAND2_X1 U10714 ( .A1(n9666), .A2(n9421), .ZN(n9422) );
  OAI211_X1 U10715 ( .C1(n9651), .C2(n9630), .A(n9423), .B(n9422), .ZN(n9424)
         );
  AOI211_X1 U10716 ( .C1(n9653), .C2(n9549), .A(n9425), .B(n9424), .ZN(n9426)
         );
  OAI21_X1 U10717 ( .B1(n9655), .B2(n9894), .A(n9426), .ZN(P1_U3265) );
  XNOR2_X1 U10718 ( .A(n9427), .B(n9428), .ZN(n9664) );
  XNOR2_X1 U10719 ( .A(n9429), .B(n9428), .ZN(n9656) );
  NAND2_X1 U10720 ( .A1(n9656), .A2(n9907), .ZN(n9438) );
  AOI211_X1 U10721 ( .C1(n9661), .C2(n9443), .A(n9889), .B(n9430), .ZN(n9659)
         );
  AOI22_X1 U10722 ( .A1(n9431), .A2(n9898), .B1(P1_REG2_REG_27__SCAN_IN), .B2(
        n4315), .ZN(n9432) );
  OAI21_X1 U10723 ( .B1(n9657), .B2(n9587), .A(n9432), .ZN(n9433) );
  AOI21_X1 U10724 ( .B1(n9434), .B2(n9568), .A(n9433), .ZN(n9435) );
  OAI21_X1 U10725 ( .B1(n4606), .B2(n9630), .A(n9435), .ZN(n9436) );
  AOI21_X1 U10726 ( .B1(n9659), .B2(n9635), .A(n9436), .ZN(n9437) );
  OAI211_X1 U10727 ( .C1(n9579), .C2(n9664), .A(n9438), .B(n9437), .ZN(
        P1_U3266) );
  XOR2_X1 U10728 ( .A(n9441), .B(n9439), .Z(n9673) );
  OAI21_X1 U10729 ( .B1(n9442), .B2(n9441), .A(n9440), .ZN(n9671) );
  INV_X1 U10730 ( .A(n9456), .ZN(n9444) );
  OAI211_X1 U10731 ( .C1(n9444), .C2(n9669), .A(n9573), .B(n9443), .ZN(n9668)
         );
  AOI22_X1 U10732 ( .A1(n9445), .A2(n9898), .B1(P1_REG2_REG_26__SCAN_IN), .B2(
        n4315), .ZN(n9446) );
  OAI21_X1 U10733 ( .B1(n9447), .B2(n9587), .A(n9446), .ZN(n9449) );
  NOR2_X1 U10734 ( .A1(n9669), .A2(n9630), .ZN(n9448) );
  AOI211_X1 U10735 ( .C1(n9568), .C2(n9666), .A(n9449), .B(n9448), .ZN(n9450)
         );
  OAI21_X1 U10736 ( .B1(n9904), .B2(n9668), .A(n9450), .ZN(n9451) );
  AOI21_X1 U10737 ( .B1(n9549), .B2(n9671), .A(n9451), .ZN(n9452) );
  OAI21_X1 U10738 ( .B1(n9673), .B2(n9894), .A(n9452), .ZN(P1_U3267) );
  XNOR2_X1 U10739 ( .A(n9453), .B(n9463), .ZN(n9676) );
  OAI22_X1 U10740 ( .A1(n9455), .A2(n9532), .B1(n9454), .B2(n9611), .ZN(n9460)
         );
  OAI211_X1 U10741 ( .C1(n9458), .C2(n9457), .A(n9573), .B(n9456), .ZN(n9674)
         );
  NOR2_X1 U10742 ( .A1(n9674), .A2(n9904), .ZN(n9459) );
  AOI211_X1 U10743 ( .C1(n9901), .C2(n9762), .A(n9460), .B(n9459), .ZN(n9467)
         );
  INV_X1 U10744 ( .A(n9461), .ZN(n9462) );
  XNOR2_X1 U10745 ( .A(n9463), .B(n9462), .ZN(n9465) );
  OAI22_X1 U10746 ( .A1(n9657), .A2(n9954), .B1(n9681), .B2(n9952), .ZN(n9464)
         );
  OR2_X1 U10747 ( .A1(n9675), .A2(n4315), .ZN(n9466) );
  OAI211_X1 U10748 ( .C1(n9676), .C2(n9894), .A(n9467), .B(n9466), .ZN(
        P1_U3268) );
  INV_X1 U10749 ( .A(n9468), .ZN(n9477) );
  NAND2_X1 U10750 ( .A1(n9469), .A2(n9635), .ZN(n9472) );
  AOI22_X1 U10751 ( .A1(n9470), .A2(n9898), .B1(P1_REG2_REG_24__SCAN_IN), .B2(
        n4315), .ZN(n9471) );
  OAI211_X1 U10752 ( .C1(n9473), .C2(n9630), .A(n9472), .B(n9471), .ZN(n9474)
         );
  AOI21_X1 U10753 ( .B1(n9611), .B2(n9475), .A(n9474), .ZN(n9476) );
  OAI21_X1 U10754 ( .B1(n9477), .B2(n9894), .A(n9476), .ZN(P1_U3269) );
  XNOR2_X1 U10755 ( .A(n9478), .B(n9479), .ZN(n9688) );
  XNOR2_X1 U10756 ( .A(n9480), .B(n9479), .ZN(n9685) );
  INV_X1 U10757 ( .A(n9481), .ZN(n9482) );
  AOI211_X1 U10758 ( .C1(n9684), .C2(n9494), .A(n9889), .B(n9482), .ZN(n9682)
         );
  NAND2_X1 U10759 ( .A1(n9682), .A2(n9635), .ZN(n9488) );
  AOI22_X1 U10760 ( .A1(n9483), .A2(n9898), .B1(n4315), .B2(
        P1_REG2_REG_23__SCAN_IN), .ZN(n9484) );
  OAI21_X1 U10761 ( .B1(n9587), .B2(n9680), .A(n9484), .ZN(n9485) );
  AOI21_X1 U10762 ( .B1(n9568), .B2(n9486), .A(n9485), .ZN(n9487) );
  OAI211_X1 U10763 ( .C1(n9489), .C2(n9630), .A(n9488), .B(n9487), .ZN(n9490)
         );
  AOI21_X1 U10764 ( .B1(n9549), .B2(n9685), .A(n9490), .ZN(n9491) );
  OAI21_X1 U10765 ( .B1(n9688), .B2(n9894), .A(n9491), .ZN(P1_U3270) );
  XNOR2_X1 U10766 ( .A(n9492), .B(n4382), .ZN(n9697) );
  XNOR2_X1 U10767 ( .A(n4382), .B(n9493), .ZN(n9695) );
  OAI211_X1 U10768 ( .C1(n9693), .C2(n9513), .A(n9573), .B(n9494), .ZN(n9692)
         );
  OAI22_X1 U10769 ( .A1(n9611), .A2(n9496), .B1(n9495), .B2(n9532), .ZN(n9498)
         );
  NOR2_X1 U10770 ( .A1(n9587), .A2(n9531), .ZN(n9497) );
  AOI211_X1 U10771 ( .C1(n9568), .C2(n9690), .A(n9498), .B(n9497), .ZN(n9501)
         );
  NAND2_X1 U10772 ( .A1(n9499), .A2(n9901), .ZN(n9500) );
  OAI211_X1 U10773 ( .C1(n9692), .C2(n9904), .A(n9501), .B(n9500), .ZN(n9502)
         );
  AOI21_X1 U10774 ( .B1(n9695), .B2(n9549), .A(n9502), .ZN(n9503) );
  OAI21_X1 U10775 ( .B1(n9697), .B2(n9894), .A(n9503), .ZN(P1_U3271) );
  XOR2_X1 U10776 ( .A(n9505), .B(n9508), .Z(n9700) );
  INV_X1 U10777 ( .A(n9700), .ZN(n9520) );
  OAI21_X1 U10778 ( .B1(n9508), .B2(n9507), .A(n9506), .ZN(n9509) );
  NAND2_X1 U10779 ( .A1(n9509), .A2(n9876), .ZN(n9512) );
  OAI22_X1 U10780 ( .A1(n9680), .A2(n9954), .B1(n9709), .B2(n9952), .ZN(n9510)
         );
  INV_X1 U10781 ( .A(n9510), .ZN(n9511) );
  NAND2_X1 U10782 ( .A1(n9512), .A2(n9511), .ZN(n9698) );
  AOI211_X1 U10783 ( .C1(n9514), .C2(n9522), .A(n9889), .B(n9513), .ZN(n9699)
         );
  NAND2_X1 U10784 ( .A1(n9699), .A2(n9635), .ZN(n9517) );
  AOI22_X1 U10785 ( .A1(n4315), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n9515), .B2(
        n9898), .ZN(n9516) );
  OAI211_X1 U10786 ( .C1(n9770), .C2(n9630), .A(n9517), .B(n9516), .ZN(n9518)
         );
  AOI21_X1 U10787 ( .B1(n9611), .B2(n9698), .A(n9518), .ZN(n9519) );
  OAI21_X1 U10788 ( .B1(n9520), .B2(n9894), .A(n9519), .ZN(P1_U3272) );
  XNOR2_X1 U10789 ( .A(n9521), .B(n9527), .ZN(n9707) );
  AOI21_X1 U10790 ( .B1(n9705), .B2(n9540), .A(n9889), .ZN(n9523) );
  AND2_X1 U10791 ( .A1(n9523), .A2(n9522), .ZN(n9704) );
  INV_X1 U10792 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n9524) );
  OAI22_X1 U10793 ( .A1(n9525), .A2(n9630), .B1(n9524), .B2(n9611), .ZN(n9526)
         );
  AOI21_X1 U10794 ( .B1(n9635), .B2(n9704), .A(n9526), .ZN(n9536) );
  XNOR2_X1 U10795 ( .A(n9528), .B(n9527), .ZN(n9529) );
  OAI222_X1 U10796 ( .A1(n9954), .A2(n9531), .B1(n9952), .B2(n9530), .C1(n9529), .C2(n9962), .ZN(n9703) );
  NOR2_X1 U10797 ( .A1(n9533), .A2(n9532), .ZN(n9534) );
  OAI21_X1 U10798 ( .B1(n9703), .B2(n9534), .A(n9611), .ZN(n9535) );
  OAI211_X1 U10799 ( .C1(n9707), .C2(n9894), .A(n9536), .B(n9535), .ZN(
        P1_U3273) );
  XOR2_X1 U10800 ( .A(n9537), .B(n9539), .Z(n9714) );
  XNOR2_X1 U10801 ( .A(n9539), .B(n9538), .ZN(n9712) );
  AOI211_X1 U10802 ( .C1(n9541), .C2(n9557), .A(n9889), .B(n4607), .ZN(n9710)
         );
  NAND2_X1 U10803 ( .A1(n9710), .A2(n9635), .ZN(n9547) );
  AOI22_X1 U10804 ( .A1(n4315), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9542), .B2(
        n9898), .ZN(n9543) );
  OAI21_X1 U10805 ( .B1(n9587), .B2(n9708), .A(n9543), .ZN(n9544) );
  AOI21_X1 U10806 ( .B1(n9568), .B2(n9545), .A(n9544), .ZN(n9546) );
  OAI211_X1 U10807 ( .C1(n9775), .C2(n9630), .A(n9547), .B(n9546), .ZN(n9548)
         );
  AOI21_X1 U10808 ( .B1(n9549), .B2(n9712), .A(n9548), .ZN(n9550) );
  OAI21_X1 U10809 ( .B1(n9714), .B2(n9894), .A(n9550), .ZN(P1_U3274) );
  XOR2_X1 U10810 ( .A(n9552), .B(n9551), .Z(n9722) );
  XOR2_X1 U10811 ( .A(n4381), .B(n9552), .Z(n9724) );
  NAND2_X1 U10812 ( .A1(n9724), .A2(n9907), .ZN(n9562) );
  AOI22_X1 U10813 ( .A1(n4315), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9553), .B2(
        n9898), .ZN(n9555) );
  NAND2_X1 U10814 ( .A1(n9568), .A2(n9718), .ZN(n9554) );
  OAI211_X1 U10815 ( .C1(n9587), .C2(n9556), .A(n9555), .B(n9554), .ZN(n9559)
         );
  OAI211_X1 U10816 ( .C1(n9779), .C2(n9572), .A(n9573), .B(n9557), .ZN(n9720)
         );
  NOR2_X1 U10817 ( .A1(n9720), .A2(n9904), .ZN(n9558) );
  AOI211_X1 U10818 ( .C1(n9901), .C2(n9560), .A(n9559), .B(n9558), .ZN(n9561)
         );
  OAI211_X1 U10819 ( .C1(n9722), .C2(n9579), .A(n9562), .B(n9561), .ZN(
        P1_U3275) );
  XNOR2_X1 U10820 ( .A(n9564), .B(n9563), .ZN(n9731) );
  XNOR2_X1 U10821 ( .A(n9566), .B(n9565), .ZN(n9733) );
  NAND2_X1 U10822 ( .A1(n9733), .A2(n9907), .ZN(n9578) );
  AOI22_X1 U10823 ( .A1(n4315), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9567), .B2(
        n9898), .ZN(n9570) );
  NAND2_X1 U10824 ( .A1(n9568), .A2(n9727), .ZN(n9569) );
  OAI211_X1 U10825 ( .C1(n9587), .C2(n9571), .A(n9570), .B(n9569), .ZN(n9576)
         );
  INV_X1 U10826 ( .A(n9572), .ZN(n9574) );
  OAI211_X1 U10827 ( .C1(n9783), .C2(n4387), .A(n9574), .B(n9573), .ZN(n9729)
         );
  NOR2_X1 U10828 ( .A1(n9729), .A2(n9904), .ZN(n9575) );
  AOI211_X1 U10829 ( .C1(n9901), .C2(n4605), .A(n9576), .B(n9575), .ZN(n9577)
         );
  OAI211_X1 U10830 ( .C1(n9731), .C2(n9579), .A(n9578), .B(n9577), .ZN(
        P1_U3276) );
  OAI21_X1 U10831 ( .B1(n9582), .B2(n9581), .A(n9580), .ZN(n9742) );
  AOI211_X1 U10832 ( .C1(n9583), .C2(n9604), .A(n9889), .B(n4387), .ZN(n9738)
         );
  NAND2_X1 U10833 ( .A1(n9583), .A2(n9901), .ZN(n9586) );
  AOI22_X1 U10834 ( .A1(n4315), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n9584), .B2(
        n9898), .ZN(n9585) );
  OAI211_X1 U10835 ( .C1(n9736), .C2(n9587), .A(n9586), .B(n9585), .ZN(n9593)
         );
  OAI21_X1 U10836 ( .B1(n9590), .B2(n9589), .A(n9588), .ZN(n9591) );
  AOI22_X1 U10837 ( .A1(n9591), .A2(n9876), .B1(n9880), .B2(n9719), .ZN(n9740)
         );
  NOR2_X1 U10838 ( .A1(n9740), .A2(n4315), .ZN(n9592) );
  AOI211_X1 U10839 ( .C1(n9738), .C2(n9635), .A(n9593), .B(n9592), .ZN(n9594)
         );
  OAI21_X1 U10840 ( .B1(n9742), .B2(n9894), .A(n9594), .ZN(P1_U3277) );
  XOR2_X1 U10841 ( .A(n9596), .B(n9595), .Z(n9745) );
  INV_X1 U10842 ( .A(n9745), .ZN(n9613) );
  NAND2_X1 U10843 ( .A1(n9597), .A2(n9596), .ZN(n9598) );
  NAND2_X1 U10844 ( .A1(n9599), .A2(n9598), .ZN(n9600) );
  NAND2_X1 U10845 ( .A1(n9600), .A2(n9876), .ZN(n9603) );
  AOI22_X1 U10846 ( .A1(n9728), .A2(n9880), .B1(n9879), .B2(n9601), .ZN(n9602)
         );
  NAND2_X1 U10847 ( .A1(n9603), .A2(n9602), .ZN(n9743) );
  INV_X1 U10848 ( .A(n9604), .ZN(n9605) );
  AOI211_X1 U10849 ( .C1(n9606), .C2(n9625), .A(n9889), .B(n9605), .ZN(n9744)
         );
  NAND2_X1 U10850 ( .A1(n9744), .A2(n9635), .ZN(n9609) );
  AOI22_X1 U10851 ( .A1(n4315), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n9607), .B2(
        n9898), .ZN(n9608) );
  OAI211_X1 U10852 ( .C1(n9789), .C2(n9630), .A(n9609), .B(n9608), .ZN(n9610)
         );
  AOI21_X1 U10853 ( .B1(n9611), .B2(n9743), .A(n9610), .ZN(n9612) );
  OAI21_X1 U10854 ( .B1(n9613), .B2(n9894), .A(n9612), .ZN(P1_U3278) );
  NAND2_X1 U10855 ( .A1(n9615), .A2(n9614), .ZN(n9616) );
  XNOR2_X1 U10856 ( .A(n9616), .B(n9618), .ZN(n9623) );
  OAI22_X1 U10857 ( .A1(n9736), .A2(n9954), .B1(n9617), .B2(n9952), .ZN(n9622)
         );
  XNOR2_X1 U10858 ( .A(n9619), .B(n9618), .ZN(n9752) );
  NOR2_X1 U10859 ( .A1(n9752), .A2(n9620), .ZN(n9621) );
  AOI211_X1 U10860 ( .C1(n9623), .C2(n9876), .A(n9622), .B(n9621), .ZN(n9751)
         );
  INV_X1 U10861 ( .A(n9624), .ZN(n9627) );
  INV_X1 U10862 ( .A(n9625), .ZN(n9626) );
  AOI211_X1 U10863 ( .C1(n9749), .C2(n9627), .A(n9889), .B(n9626), .ZN(n9748)
         );
  AOI22_X1 U10864 ( .A1(n4315), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n9628), .B2(
        n9898), .ZN(n9629) );
  OAI21_X1 U10865 ( .B1(n9631), .B2(n9630), .A(n9629), .ZN(n9634) );
  NOR2_X1 U10866 ( .A1(n9752), .A2(n9632), .ZN(n9633) );
  AOI211_X1 U10867 ( .C1(n9748), .C2(n9635), .A(n9634), .B(n9633), .ZN(n9636)
         );
  OAI21_X1 U10868 ( .B1(n9751), .B2(n4315), .A(n9636), .ZN(P1_U3279) );
  INV_X1 U10869 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n9639) );
  MUX2_X1 U10870 ( .A(n9639), .B(n9753), .S(n9983), .Z(n9640) );
  OAI21_X1 U10871 ( .B1(n9755), .B2(n9747), .A(n9640), .ZN(P1_U3553) );
  NAND2_X1 U10872 ( .A1(n9641), .A2(n9964), .ZN(n9647) );
  OAI22_X1 U10873 ( .A1(n9642), .A2(n9947), .B1(n9658), .B2(n9952), .ZN(n9643)
         );
  NAND2_X1 U10874 ( .A1(n9647), .A2(n9646), .ZN(n9756) );
  MUX2_X1 U10875 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n9756), .S(n9983), .Z(
        P1_U3551) );
  AOI22_X1 U10876 ( .A1(n9666), .A2(n9879), .B1(n9648), .B2(n9880), .ZN(n9649)
         );
  OAI211_X1 U10877 ( .C1(n9651), .C2(n9947), .A(n9650), .B(n9649), .ZN(n9652)
         );
  AOI21_X1 U10878 ( .B1(n9653), .B2(n9876), .A(n9652), .ZN(n9654) );
  OAI21_X1 U10879 ( .B1(n9655), .B2(n9741), .A(n9654), .ZN(n9757) );
  MUX2_X1 U10880 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9757), .S(n9983), .Z(
        P1_U3550) );
  NAND2_X1 U10881 ( .A1(n9656), .A2(n9964), .ZN(n9663) );
  OAI22_X1 U10882 ( .A1(n9658), .A2(n9954), .B1(n9657), .B2(n9952), .ZN(n9660)
         );
  AOI211_X1 U10883 ( .C1(n9959), .C2(n9661), .A(n9660), .B(n9659), .ZN(n9662)
         );
  OAI211_X1 U10884 ( .C1(n9962), .C2(n9664), .A(n9663), .B(n9662), .ZN(n9758)
         );
  MUX2_X1 U10885 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9758), .S(n9983), .Z(
        P1_U3549) );
  AOI22_X1 U10886 ( .A1(n9666), .A2(n9880), .B1(n9879), .B2(n9665), .ZN(n9667)
         );
  OAI211_X1 U10887 ( .C1(n9669), .C2(n9947), .A(n9668), .B(n9667), .ZN(n9670)
         );
  AOI21_X1 U10888 ( .B1(n9671), .B2(n9876), .A(n9670), .ZN(n9672) );
  OAI21_X1 U10889 ( .B1(n9673), .B2(n9741), .A(n9672), .ZN(n9759) );
  MUX2_X1 U10890 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9759), .S(n9983), .Z(
        P1_U3548) );
  OAI211_X1 U10891 ( .C1(n9676), .C2(n9741), .A(n9675), .B(n9674), .ZN(n9760)
         );
  MUX2_X1 U10892 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9760), .S(n9983), .Z(n9677) );
  AOI21_X1 U10893 ( .B1(n9678), .B2(n9762), .A(n9677), .ZN(n9679) );
  INV_X1 U10894 ( .A(n9679), .ZN(P1_U3547) );
  OAI22_X1 U10895 ( .A1(n9681), .A2(n9954), .B1(n9680), .B2(n9952), .ZN(n9683)
         );
  AOI211_X1 U10896 ( .C1(n9959), .C2(n9684), .A(n9683), .B(n9682), .ZN(n9687)
         );
  NAND2_X1 U10897 ( .A1(n9685), .A2(n9876), .ZN(n9686) );
  OAI211_X1 U10898 ( .C1(n9688), .C2(n9741), .A(n9687), .B(n9686), .ZN(n9765)
         );
  MUX2_X1 U10899 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9765), .S(n9983), .Z(
        P1_U3545) );
  AOI22_X1 U10900 ( .A1(n9690), .A2(n9880), .B1(n9689), .B2(n9879), .ZN(n9691)
         );
  OAI211_X1 U10901 ( .C1(n9693), .C2(n9947), .A(n9692), .B(n9691), .ZN(n9694)
         );
  AOI21_X1 U10902 ( .B1(n9695), .B2(n9876), .A(n9694), .ZN(n9696) );
  OAI21_X1 U10903 ( .B1(n9697), .B2(n9741), .A(n9696), .ZN(n9766) );
  MUX2_X1 U10904 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9766), .S(n9983), .Z(
        P1_U3544) );
  INV_X1 U10905 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n9701) );
  AOI211_X1 U10906 ( .C1(n9700), .C2(n9964), .A(n9699), .B(n9698), .ZN(n9767)
         );
  MUX2_X1 U10907 ( .A(n9701), .B(n9767), .S(n9983), .Z(n9702) );
  OAI21_X1 U10908 ( .B1(n9770), .B2(n9747), .A(n9702), .ZN(P1_U3543) );
  AOI211_X1 U10909 ( .C1(n9959), .C2(n9705), .A(n9704), .B(n9703), .ZN(n9706)
         );
  OAI21_X1 U10910 ( .B1(n9707), .B2(n9741), .A(n9706), .ZN(n9771) );
  MUX2_X1 U10911 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9771), .S(n9983), .Z(
        P1_U3542) );
  INV_X1 U10912 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n9716) );
  OAI22_X1 U10913 ( .A1(n9709), .A2(n9954), .B1(n9708), .B2(n9952), .ZN(n9711)
         );
  AOI211_X1 U10914 ( .C1(n9712), .C2(n9876), .A(n9711), .B(n9710), .ZN(n9713)
         );
  OAI21_X1 U10915 ( .B1(n9714), .B2(n9741), .A(n9713), .ZN(n9715) );
  INV_X1 U10916 ( .A(n9715), .ZN(n9772) );
  MUX2_X1 U10917 ( .A(n9716), .B(n9772), .S(n9983), .Z(n9717) );
  OAI21_X1 U10918 ( .B1(n9775), .B2(n9747), .A(n9717), .ZN(P1_U3541) );
  AOI22_X1 U10919 ( .A1(n9719), .A2(n9879), .B1(n9880), .B2(n9718), .ZN(n9721)
         );
  OAI211_X1 U10920 ( .C1(n9722), .C2(n9962), .A(n9721), .B(n9720), .ZN(n9723)
         );
  AOI21_X1 U10921 ( .B1(n9724), .B2(n9964), .A(n9723), .ZN(n9776) );
  MUX2_X1 U10922 ( .A(n9725), .B(n9776), .S(n9983), .Z(n9726) );
  OAI21_X1 U10923 ( .B1(n9779), .B2(n9747), .A(n9726), .ZN(P1_U3540) );
  AOI22_X1 U10924 ( .A1(n9728), .A2(n9879), .B1(n9880), .B2(n9727), .ZN(n9730)
         );
  OAI211_X1 U10925 ( .C1(n9731), .C2(n9962), .A(n9730), .B(n9729), .ZN(n9732)
         );
  AOI21_X1 U10926 ( .B1(n9733), .B2(n9964), .A(n9732), .ZN(n9780) );
  MUX2_X1 U10927 ( .A(n9734), .B(n9780), .S(n9983), .Z(n9735) );
  OAI21_X1 U10928 ( .B1(n9783), .B2(n9747), .A(n9735), .ZN(P1_U3539) );
  OAI22_X1 U10929 ( .A1(n4603), .A2(n9947), .B1(n9736), .B2(n9952), .ZN(n9737)
         );
  NOR2_X1 U10930 ( .A1(n9738), .A2(n9737), .ZN(n9739) );
  OAI211_X1 U10931 ( .C1(n9742), .C2(n9741), .A(n9740), .B(n9739), .ZN(n9784)
         );
  MUX2_X1 U10932 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9784), .S(n9983), .Z(
        P1_U3538) );
  AOI211_X1 U10933 ( .C1(n9745), .C2(n9964), .A(n9744), .B(n9743), .ZN(n9785)
         );
  MUX2_X1 U10934 ( .A(n9859), .B(n9785), .S(n9983), .Z(n9746) );
  OAI21_X1 U10935 ( .B1(n9789), .B2(n9747), .A(n9746), .ZN(P1_U3537) );
  AOI21_X1 U10936 ( .B1(n9959), .B2(n9749), .A(n9748), .ZN(n9750) );
  OAI211_X1 U10937 ( .C1(n9914), .C2(n9752), .A(n9751), .B(n9750), .ZN(n9790)
         );
  MUX2_X1 U10938 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n9790), .S(n9983), .Z(
        P1_U3536) );
  OAI21_X1 U10939 ( .B1(n9755), .B2(n9788), .A(n9754), .ZN(P1_U3521) );
  MUX2_X1 U10940 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n9756), .S(n9968), .Z(
        P1_U3519) );
  MUX2_X1 U10941 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n9757), .S(n9968), .Z(
        P1_U3518) );
  MUX2_X1 U10942 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9758), .S(n9968), .Z(
        P1_U3517) );
  MUX2_X1 U10943 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9759), .S(n9968), .Z(
        P1_U3516) );
  MUX2_X1 U10944 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9760), .S(n9968), .Z(n9761) );
  AOI21_X1 U10945 ( .B1(n9763), .B2(n9762), .A(n9761), .ZN(n9764) );
  INV_X1 U10946 ( .A(n9764), .ZN(P1_U3515) );
  MUX2_X1 U10947 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9765), .S(n9968), .Z(
        P1_U3513) );
  MUX2_X1 U10948 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9766), .S(n9968), .Z(
        P1_U3512) );
  INV_X1 U10949 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n9768) );
  MUX2_X1 U10950 ( .A(n9768), .B(n9767), .S(n9968), .Z(n9769) );
  OAI21_X1 U10951 ( .B1(n9770), .B2(n9788), .A(n9769), .ZN(P1_U3511) );
  MUX2_X1 U10952 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9771), .S(n9968), .Z(
        P1_U3510) );
  INV_X1 U10953 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n9773) );
  MUX2_X1 U10954 ( .A(n9773), .B(n9772), .S(n9968), .Z(n9774) );
  OAI21_X1 U10955 ( .B1(n9775), .B2(n9788), .A(n9774), .ZN(P1_U3509) );
  INV_X1 U10956 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n9777) );
  MUX2_X1 U10957 ( .A(n9777), .B(n9776), .S(n9968), .Z(n9778) );
  OAI21_X1 U10958 ( .B1(n9779), .B2(n9788), .A(n9778), .ZN(P1_U3507) );
  INV_X1 U10959 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n9781) );
  MUX2_X1 U10960 ( .A(n9781), .B(n9780), .S(n9968), .Z(n9782) );
  OAI21_X1 U10961 ( .B1(n9783), .B2(n9788), .A(n9782), .ZN(P1_U3504) );
  MUX2_X1 U10962 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n9784), .S(n9968), .Z(
        P1_U3501) );
  INV_X1 U10963 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n9786) );
  MUX2_X1 U10964 ( .A(n9786), .B(n9785), .S(n9968), .Z(n9787) );
  OAI21_X1 U10965 ( .B1(n9789), .B2(n9788), .A(n9787), .ZN(P1_U3498) );
  MUX2_X1 U10966 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n9790), .S(n9968), .Z(
        P1_U3495) );
  MUX2_X1 U10967 ( .A(n9791), .B(P1_D_REG_1__SCAN_IN), .S(n9913), .Z(P1_U3440)
         );
  MUX2_X1 U10968 ( .A(n9792), .B(P1_D_REG_0__SCAN_IN), .S(n9913), .Z(P1_U3439)
         );
  NOR4_X1 U10969 ( .A1(n5127), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3086), .A4(
        n9793), .ZN(n9794) );
  AOI21_X1 U10970 ( .B1(n9795), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9794), .ZN(
        n9796) );
  OAI21_X1 U10971 ( .B1(n9798), .B2(n9797), .A(n9796), .ZN(P1_U3324) );
  MUX2_X1 U10972 ( .A(n9800), .B(n9799), .S(P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  AOI211_X1 U10973 ( .C1(n9803), .C2(n9802), .A(n9861), .B(n9801), .ZN(n9808)
         );
  AOI211_X1 U10974 ( .C1(n9806), .C2(n9805), .A(n9857), .B(n9804), .ZN(n9807)
         );
  AOI211_X1 U10975 ( .C1(n9868), .C2(n9809), .A(n9808), .B(n9807), .ZN(n9811)
         );
  NAND2_X1 U10976 ( .A1(P1_REG3_REG_10__SCAN_IN), .A2(P1_U3086), .ZN(n9810) );
  OAI211_X1 U10977 ( .C1(n9872), .C2(n9812), .A(n9811), .B(n9810), .ZN(
        P1_U3253) );
  XNOR2_X1 U10978 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U10979 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  AOI211_X1 U10980 ( .C1(n9815), .C2(n9814), .A(n9813), .B(n9861), .ZN(n9820)
         );
  AOI211_X1 U10981 ( .C1(n9818), .C2(n9817), .A(n9816), .B(n9857), .ZN(n9819)
         );
  AOI211_X1 U10982 ( .C1(n9868), .C2(n9821), .A(n9820), .B(n9819), .ZN(n9823)
         );
  NAND2_X1 U10983 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n9822) );
  OAI211_X1 U10984 ( .C1(n9872), .C2(n9824), .A(n9823), .B(n9822), .ZN(
        P1_U3254) );
  AOI211_X1 U10985 ( .C1(n9827), .C2(n9826), .A(n9825), .B(n9857), .ZN(n9832)
         );
  AOI211_X1 U10986 ( .C1(n9830), .C2(n9829), .A(n9828), .B(n9861), .ZN(n9831)
         );
  AOI211_X1 U10987 ( .C1(n9868), .C2(n9833), .A(n9832), .B(n9831), .ZN(n9835)
         );
  NAND2_X1 U10988 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3086), .ZN(n9834) );
  OAI211_X1 U10989 ( .C1(n9872), .C2(n9836), .A(n9835), .B(n9834), .ZN(
        P1_U3256) );
  INV_X1 U10990 ( .A(n9837), .ZN(n9850) );
  AOI21_X1 U10991 ( .B1(n9840), .B2(n9839), .A(n9838), .ZN(n9841) );
  NAND2_X1 U10992 ( .A1(n9842), .A2(n9841), .ZN(n9849) );
  AOI21_X1 U10993 ( .B1(n9845), .B2(n9844), .A(n9843), .ZN(n9846) );
  NAND2_X1 U10994 ( .A1(n9847), .A2(n9846), .ZN(n9848) );
  OAI211_X1 U10995 ( .C1(n9851), .C2(n9850), .A(n9849), .B(n9848), .ZN(n9852)
         );
  INV_X1 U10996 ( .A(n9852), .ZN(n9854) );
  OAI211_X1 U10997 ( .C1(n9872), .C2(n9855), .A(n9854), .B(n9853), .ZN(
        P1_U3257) );
  INV_X1 U10998 ( .A(n9856), .ZN(n9867) );
  AOI211_X1 U10999 ( .C1(n9860), .C2(n9859), .A(n9858), .B(n9857), .ZN(n9866)
         );
  AOI211_X1 U11000 ( .C1(n9864), .C2(n9863), .A(n9862), .B(n9861), .ZN(n9865)
         );
  AOI211_X1 U11001 ( .C1(n9868), .C2(n9867), .A(n9866), .B(n9865), .ZN(n9870)
         );
  NAND2_X1 U11002 ( .A1(P1_REG3_REG_15__SCAN_IN), .A2(P1_U3086), .ZN(n9869) );
  OAI211_X1 U11003 ( .C1(n9872), .C2(n9871), .A(n9870), .B(n9869), .ZN(
        P1_U3258) );
  NAND2_X1 U11004 ( .A1(n9874), .A2(n9873), .ZN(n9875) );
  XNOR2_X1 U11005 ( .A(n9875), .B(n9885), .ZN(n9877) );
  NAND2_X1 U11006 ( .A1(n9877), .A2(n9876), .ZN(n9883) );
  AOI22_X1 U11007 ( .A1(n9881), .A2(n9880), .B1(n9879), .B2(n9878), .ZN(n9882)
         );
  AOI222_X1 U11008 ( .A1(n9890), .A2(n9901), .B1(P1_REG2_REG_12__SCAN_IN), 
        .B2(n4315), .C1(n9884), .C2(n9898), .ZN(n9897) );
  NOR2_X1 U11009 ( .A1(n9886), .A2(n9885), .ZN(n9887) );
  OR2_X1 U11010 ( .A1(n9888), .A2(n9887), .ZN(n9944) );
  AOI21_X1 U11011 ( .B1(n9891), .B2(n9890), .A(n9889), .ZN(n9893) );
  NAND2_X1 U11012 ( .A1(n9893), .A2(n9892), .ZN(n9945) );
  OAI22_X1 U11013 ( .A1(n9944), .A2(n9894), .B1(n9945), .B2(n9904), .ZN(n9895)
         );
  INV_X1 U11014 ( .A(n9895), .ZN(n9896) );
  OAI211_X1 U11015 ( .C1(n4315), .C2(n9946), .A(n9897), .B(n9896), .ZN(
        P1_U3281) );
  AOI22_X1 U11016 ( .A1(n4315), .A2(P1_REG2_REG_5__SCAN_IN), .B1(n9899), .B2(
        n9898), .ZN(n9903) );
  NAND2_X1 U11017 ( .A1(n9901), .A2(n9900), .ZN(n9902) );
  OAI211_X1 U11018 ( .C1(n9905), .C2(n9904), .A(n9903), .B(n9902), .ZN(n9906)
         );
  AOI21_X1 U11019 ( .B1(n9908), .B2(n9907), .A(n9906), .ZN(n9909) );
  OAI21_X1 U11020 ( .B1(n4315), .B2(n9910), .A(n9909), .ZN(P1_U3288) );
  AND2_X1 U11021 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n9913), .ZN(P1_U3294) );
  AND2_X1 U11022 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n9913), .ZN(P1_U3295) );
  AND2_X1 U11023 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n9913), .ZN(P1_U3296) );
  AND2_X1 U11024 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n9913), .ZN(P1_U3297) );
  AND2_X1 U11025 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n9913), .ZN(P1_U3298) );
  AND2_X1 U11026 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n9913), .ZN(P1_U3299) );
  AND2_X1 U11027 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n9913), .ZN(P1_U3300) );
  AND2_X1 U11028 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9913), .ZN(P1_U3301) );
  AND2_X1 U11029 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n9913), .ZN(P1_U3302) );
  AND2_X1 U11030 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n9913), .ZN(P1_U3303) );
  AND2_X1 U11031 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n9913), .ZN(P1_U3304) );
  AND2_X1 U11032 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n9913), .ZN(P1_U3305) );
  INV_X1 U11033 ( .A(n9913), .ZN(n9912) );
  NOR2_X1 U11034 ( .A1(n9912), .A2(n9911), .ZN(P1_U3306) );
  AND2_X1 U11035 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n9913), .ZN(P1_U3307) );
  AND2_X1 U11036 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n9913), .ZN(P1_U3308) );
  AND2_X1 U11037 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n9913), .ZN(P1_U3309) );
  AND2_X1 U11038 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n9913), .ZN(P1_U3310) );
  AND2_X1 U11039 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n9913), .ZN(P1_U3311) );
  AND2_X1 U11040 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n9913), .ZN(P1_U3312) );
  AND2_X1 U11041 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n9913), .ZN(P1_U3313) );
  AND2_X1 U11042 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n9913), .ZN(P1_U3314) );
  AND2_X1 U11043 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n9913), .ZN(P1_U3315) );
  AND2_X1 U11044 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n9913), .ZN(P1_U3316) );
  AND2_X1 U11045 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n9913), .ZN(P1_U3317) );
  AND2_X1 U11046 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n9913), .ZN(P1_U3318) );
  AND2_X1 U11047 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n9913), .ZN(P1_U3319) );
  AND2_X1 U11048 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n9913), .ZN(P1_U3320) );
  AND2_X1 U11049 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n9913), .ZN(P1_U3321) );
  AND2_X1 U11050 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n9913), .ZN(P1_U3322) );
  AND2_X1 U11051 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n9913), .ZN(P1_U3323) );
  INV_X1 U11052 ( .A(n9914), .ZN(n9936) );
  OAI21_X1 U11053 ( .B1(n7219), .B2(n9947), .A(n9915), .ZN(n9917) );
  AOI211_X1 U11054 ( .C1(n9936), .C2(n9918), .A(n9917), .B(n9916), .ZN(n9970)
         );
  AOI22_X1 U11055 ( .A1(n9968), .A2(n9970), .B1(n9919), .B2(n9966), .ZN(
        P1_U3459) );
  OAI21_X1 U11056 ( .B1(n9921), .B2(n9947), .A(n9920), .ZN(n9923) );
  AOI211_X1 U11057 ( .C1(n9964), .C2(n9924), .A(n9923), .B(n9922), .ZN(n9972)
         );
  INV_X1 U11058 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n9925) );
  AOI22_X1 U11059 ( .A1(n9968), .A2(n9972), .B1(n9925), .B2(n9966), .ZN(
        P1_U3465) );
  OAI21_X1 U11060 ( .B1(n9927), .B2(n9947), .A(n9926), .ZN(n9929) );
  AOI211_X1 U11061 ( .C1(n9964), .C2(n9930), .A(n9929), .B(n9928), .ZN(n9974)
         );
  INV_X1 U11062 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n9931) );
  AOI22_X1 U11063 ( .A1(n9968), .A2(n9974), .B1(n9931), .B2(n9966), .ZN(
        P1_U3471) );
  OAI21_X1 U11064 ( .B1(n4593), .B2(n9947), .A(n9932), .ZN(n9934) );
  AOI211_X1 U11065 ( .C1(n9936), .C2(n9935), .A(n9934), .B(n9933), .ZN(n9976)
         );
  INV_X1 U11066 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n9937) );
  AOI22_X1 U11067 ( .A1(n9968), .A2(n9976), .B1(n9937), .B2(n9966), .ZN(
        P1_U3477) );
  OAI211_X1 U11068 ( .C1(n9940), .C2(n9947), .A(n9939), .B(n9938), .ZN(n9941)
         );
  AOI21_X1 U11069 ( .B1(n9964), .B2(n9942), .A(n9941), .ZN(n9978) );
  INV_X1 U11070 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n9943) );
  AOI22_X1 U11071 ( .A1(n9968), .A2(n9978), .B1(n9943), .B2(n9966), .ZN(
        P1_U3480) );
  INV_X1 U11072 ( .A(n9944), .ZN(n9950) );
  OAI211_X1 U11073 ( .C1(n9948), .C2(n9947), .A(n9946), .B(n9945), .ZN(n9949)
         );
  AOI21_X1 U11074 ( .B1(n9950), .B2(n9964), .A(n9949), .ZN(n9980) );
  INV_X1 U11075 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n9951) );
  AOI22_X1 U11076 ( .A1(n9968), .A2(n9980), .B1(n9951), .B2(n9966), .ZN(
        P1_U3489) );
  OAI22_X1 U11077 ( .A1(n9955), .A2(n9954), .B1(n9953), .B2(n9952), .ZN(n9957)
         );
  AOI211_X1 U11078 ( .C1(n9959), .C2(n9958), .A(n9957), .B(n9956), .ZN(n9960)
         );
  OAI21_X1 U11079 ( .B1(n9962), .B2(n9961), .A(n9960), .ZN(n9963) );
  AOI21_X1 U11080 ( .B1(n9965), .B2(n9964), .A(n9963), .ZN(n9982) );
  INV_X1 U11081 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n9967) );
  AOI22_X1 U11082 ( .A1(n9968), .A2(n9982), .B1(n9967), .B2(n9966), .ZN(
        P1_U3492) );
  INV_X1 U11083 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n9969) );
  AOI22_X1 U11084 ( .A1(n9983), .A2(n9970), .B1(n9969), .B2(n9981), .ZN(
        P1_U3524) );
  INV_X1 U11085 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n9971) );
  AOI22_X1 U11086 ( .A1(n9983), .A2(n9972), .B1(n9971), .B2(n9981), .ZN(
        P1_U3526) );
  AOI22_X1 U11087 ( .A1(n9983), .A2(n9974), .B1(n9973), .B2(n9981), .ZN(
        P1_U3528) );
  INV_X1 U11088 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n9975) );
  AOI22_X1 U11089 ( .A1(n9983), .A2(n9976), .B1(n9975), .B2(n9981), .ZN(
        P1_U3530) );
  INV_X1 U11090 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n9977) );
  AOI22_X1 U11091 ( .A1(n9983), .A2(n9978), .B1(n9977), .B2(n9981), .ZN(
        P1_U3531) );
  AOI22_X1 U11092 ( .A1(n9983), .A2(n9980), .B1(n9979), .B2(n9981), .ZN(
        P1_U3534) );
  AOI22_X1 U11093 ( .A1(n9983), .A2(n9982), .B1(n7903), .B2(n9981), .ZN(
        P1_U3535) );
  AOI22_X1 U11094 ( .A1(n10051), .A2(n9984), .B1(n10049), .B2(
        P2_ADDR_REG_13__SCAN_IN), .ZN(n10001) );
  OAI21_X1 U11095 ( .B1(P2_REG1_REG_13__SCAN_IN), .B2(n9986), .A(n9985), .ZN(
        n9993) );
  NAND2_X1 U11096 ( .A1(n9988), .A2(n9987), .ZN(n9990) );
  AOI21_X1 U11097 ( .B1(n9991), .B2(n9990), .A(n9989), .ZN(n9992) );
  AOI21_X1 U11098 ( .B1(n9993), .B2(n10058), .A(n9992), .ZN(n10000) );
  NAND2_X1 U11099 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(P2_U3151), .ZN(n9999) );
  AOI21_X1 U11100 ( .B1(n9996), .B2(n9995), .A(n9994), .ZN(n9997) );
  OR2_X1 U11101 ( .A1(n9997), .A2(n10064), .ZN(n9998) );
  NAND4_X1 U11102 ( .A1(n10001), .A2(n10000), .A3(n9999), .A4(n9998), .ZN(
        P2_U3195) );
  AOI22_X1 U11103 ( .A1(n10051), .A2(n10002), .B1(n10049), .B2(
        P2_ADDR_REG_14__SCAN_IN), .ZN(n10016) );
  OAI21_X1 U11104 ( .B1(n10005), .B2(n10004), .A(n10003), .ZN(n10009) );
  XNOR2_X1 U11105 ( .A(n10007), .B(n10006), .ZN(n10008) );
  AOI22_X1 U11106 ( .A1(n10009), .A2(n10058), .B1(n10057), .B2(n10008), .ZN(
        n10015) );
  NAND2_X1 U11107 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3151), .ZN(n10014)
         );
  AOI21_X1 U11108 ( .B1(n4390), .B2(n10011), .A(n10010), .ZN(n10012) );
  OR2_X1 U11109 ( .A1(n10012), .A2(n10064), .ZN(n10013) );
  NAND4_X1 U11110 ( .A1(n10016), .A2(n10015), .A3(n10014), .A4(n10013), .ZN(
        P2_U3196) );
  AOI22_X1 U11111 ( .A1(n10051), .A2(n10017), .B1(n10049), .B2(
        P2_ADDR_REG_15__SCAN_IN), .ZN(n10032) );
  OAI21_X1 U11112 ( .B1(P2_REG1_REG_15__SCAN_IN), .B2(n10019), .A(n10018), 
        .ZN(n10023) );
  XNOR2_X1 U11113 ( .A(n10021), .B(n10020), .ZN(n10022) );
  AOI22_X1 U11114 ( .A1(n10023), .A2(n10058), .B1(n10057), .B2(n10022), .ZN(
        n10031) );
  INV_X1 U11115 ( .A(n10024), .ZN(n10025) );
  NOR2_X1 U11116 ( .A1(n10025), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n10027) );
  OAI21_X1 U11117 ( .B1(n10028), .B2(n10027), .A(n10026), .ZN(n10029) );
  NAND4_X1 U11118 ( .A1(n10032), .A2(n10031), .A3(n10030), .A4(n10029), .ZN(
        P2_U3197) );
  AOI22_X1 U11119 ( .A1(n10051), .A2(n10033), .B1(n10049), .B2(
        P2_ADDR_REG_16__SCAN_IN), .ZN(n10048) );
  OAI21_X1 U11120 ( .B1(n10036), .B2(n10035), .A(n10034), .ZN(n10040) );
  XNOR2_X1 U11121 ( .A(n10038), .B(n10037), .ZN(n10039) );
  AOI22_X1 U11122 ( .A1(n10040), .A2(n10058), .B1(n10057), .B2(n10039), .ZN(
        n10047) );
  NAND2_X1 U11123 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(P2_U3151), .ZN(n10046)
         );
  AOI21_X1 U11124 ( .B1(n4348), .B2(n10043), .A(n10042), .ZN(n10044) );
  OR2_X1 U11125 ( .A1(n10044), .A2(n10064), .ZN(n10045) );
  NAND4_X1 U11126 ( .A1(n10048), .A2(n10047), .A3(n10046), .A4(n10045), .ZN(
        P2_U3198) );
  AOI22_X1 U11127 ( .A1(n10051), .A2(n10050), .B1(n10049), .B2(
        P2_ADDR_REG_17__SCAN_IN), .ZN(n10068) );
  OAI21_X1 U11128 ( .B1(P2_REG1_REG_17__SCAN_IN), .B2(n10053), .A(n10052), 
        .ZN(n10059) );
  XNOR2_X1 U11129 ( .A(n10055), .B(n10054), .ZN(n10056) );
  AOI22_X1 U11130 ( .A1(n10059), .A2(n10058), .B1(n10057), .B2(n10056), .ZN(
        n10067) );
  AOI21_X1 U11131 ( .B1(n10062), .B2(n10061), .A(n10060), .ZN(n10063) );
  OR2_X1 U11132 ( .A1(n10064), .A2(n10063), .ZN(n10065) );
  NAND4_X1 U11133 ( .A1(n10068), .A2(n10067), .A3(n10066), .A4(n10065), .ZN(
        P2_U3199) );
  NAND2_X1 U11134 ( .A1(n10070), .A2(n10069), .ZN(n10073) );
  INV_X1 U11135 ( .A(n10071), .ZN(n10072) );
  AOI21_X1 U11136 ( .B1(n10078), .B2(n10073), .A(n10072), .ZN(n10127) );
  OAI22_X1 U11137 ( .A1(n10077), .A2(n10076), .B1(n10075), .B2(n10074), .ZN(
        n10083) );
  XOR2_X1 U11138 ( .A(n10079), .B(n10078), .Z(n10081) );
  NOR2_X1 U11139 ( .A1(n10081), .A2(n10080), .ZN(n10082) );
  AOI211_X1 U11140 ( .C1(n10084), .C2(n10127), .A(n10083), .B(n10082), .ZN(
        n10129) );
  AOI222_X1 U11141 ( .A1(n10088), .A2(n10087), .B1(n10127), .B2(n10086), .C1(
        n10125), .C2(n10085), .ZN(n10089) );
  OAI221_X1 U11142 ( .B1(n10092), .B2(n10129), .C1(n10091), .C2(n10090), .A(
        n10089), .ZN(P2_U3226) );
  INV_X1 U11143 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n10096) );
  INV_X1 U11144 ( .A(n10136), .ZN(n10126) );
  NOR2_X1 U11145 ( .A1(n7055), .A2(n10118), .ZN(n10094) );
  AOI211_X1 U11146 ( .C1(n10126), .C2(n10095), .A(n10094), .B(n10093), .ZN(
        n10146) );
  AOI22_X1 U11147 ( .A1(n10144), .A2(n10096), .B1(n10146), .B2(n10142), .ZN(
        P2_U3393) );
  INV_X1 U11148 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n10101) );
  OAI22_X1 U11149 ( .A1(n10098), .A2(n10136), .B1(n10097), .B2(n10118), .ZN(
        n10099) );
  NOR2_X1 U11150 ( .A1(n10100), .A2(n10099), .ZN(n10147) );
  AOI22_X1 U11151 ( .A1(n10144), .A2(n10101), .B1(n10147), .B2(n10142), .ZN(
        P2_U3396) );
  INV_X1 U11152 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n10106) );
  OAI21_X1 U11153 ( .B1(n7072), .B2(n10118), .A(n10102), .ZN(n10103) );
  AOI21_X1 U11154 ( .B1(n10105), .B2(n10104), .A(n10103), .ZN(n10148) );
  AOI22_X1 U11155 ( .A1(n10144), .A2(n10106), .B1(n10148), .B2(n10142), .ZN(
        P2_U3399) );
  INV_X1 U11156 ( .A(n10107), .ZN(n10110) );
  OAI22_X1 U11157 ( .A1(n10108), .A2(n10120), .B1(n6853), .B2(n10118), .ZN(
        n10109) );
  NOR2_X1 U11158 ( .A1(n10110), .A2(n10109), .ZN(n10150) );
  AOI22_X1 U11159 ( .A1(n10144), .A2(n10111), .B1(n10150), .B2(n10142), .ZN(
        P2_U3402) );
  INV_X1 U11160 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n10116) );
  OAI22_X1 U11161 ( .A1(n10113), .A2(n10136), .B1(n10112), .B2(n10118), .ZN(
        n10115) );
  NOR2_X1 U11162 ( .A1(n10115), .A2(n10114), .ZN(n10152) );
  AOI22_X1 U11163 ( .A1(n10144), .A2(n10116), .B1(n10152), .B2(n10142), .ZN(
        P2_U3405) );
  INV_X1 U11164 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10124) );
  INV_X1 U11165 ( .A(n10117), .ZN(n10123) );
  OAI22_X1 U11166 ( .A1(n10121), .A2(n10120), .B1(n10119), .B2(n10118), .ZN(
        n10122) );
  NOR2_X1 U11167 ( .A1(n10123), .A2(n10122), .ZN(n10153) );
  AOI22_X1 U11168 ( .A1(n10144), .A2(n10124), .B1(n10153), .B2(n10142), .ZN(
        P2_U3408) );
  INV_X1 U11169 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n10130) );
  AOI22_X1 U11170 ( .A1(n10127), .A2(n10126), .B1(n10141), .B2(n10125), .ZN(
        n10128) );
  AND2_X1 U11171 ( .A1(n10129), .A2(n10128), .ZN(n10154) );
  AOI22_X1 U11172 ( .A1(n10144), .A2(n10130), .B1(n10154), .B2(n10142), .ZN(
        P2_U3411) );
  INV_X1 U11173 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n10135) );
  NOR2_X1 U11174 ( .A1(n10131), .A2(n10136), .ZN(n10133) );
  AOI211_X1 U11175 ( .C1(n10141), .C2(n10134), .A(n10133), .B(n10132), .ZN(
        n10155) );
  AOI22_X1 U11176 ( .A1(n10144), .A2(n10135), .B1(n10155), .B2(n10142), .ZN(
        P2_U3417) );
  INV_X1 U11177 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n10143) );
  NOR2_X1 U11178 ( .A1(n10137), .A2(n10136), .ZN(n10139) );
  AOI211_X1 U11179 ( .C1(n10141), .C2(n10140), .A(n10139), .B(n10138), .ZN(
        n10157) );
  AOI22_X1 U11180 ( .A1(n10144), .A2(n10143), .B1(n10157), .B2(n10142), .ZN(
        P2_U3420) );
  INV_X1 U11181 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n10145) );
  AOI22_X1 U11182 ( .A1(n10158), .A2(n10146), .B1(n10145), .B2(n10156), .ZN(
        P2_U3460) );
  AOI22_X1 U11183 ( .A1(n10158), .A2(n10147), .B1(n6619), .B2(n10156), .ZN(
        P2_U3461) );
  AOI22_X1 U11184 ( .A1(n10158), .A2(n10148), .B1(n6671), .B2(n10156), .ZN(
        P2_U3462) );
  AOI22_X1 U11185 ( .A1(n10158), .A2(n10150), .B1(n10149), .B2(n10156), .ZN(
        P2_U3463) );
  INV_X1 U11186 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n10151) );
  AOI22_X1 U11187 ( .A1(n10158), .A2(n10152), .B1(n10151), .B2(n10156), .ZN(
        P2_U3464) );
  AOI22_X1 U11188 ( .A1(n10158), .A2(n10153), .B1(n6774), .B2(n10156), .ZN(
        P2_U3465) );
  AOI22_X1 U11189 ( .A1(n10158), .A2(n10154), .B1(n6996), .B2(n10156), .ZN(
        P2_U3466) );
  AOI22_X1 U11190 ( .A1(n10158), .A2(n10155), .B1(n7106), .B2(n10156), .ZN(
        P2_U3468) );
  AOI22_X1 U11191 ( .A1(n10158), .A2(n10157), .B1(n7193), .B2(n10156), .ZN(
        P2_U3469) );
  NOR2_X1 U11192 ( .A1(n10160), .A2(n10159), .ZN(n10161) );
  XOR2_X1 U11193 ( .A(n10161), .B(P2_ADDR_REG_1__SCAN_IN), .Z(ADD_1068_U5) );
  XOR2_X1 U11194 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1068_U46) );
  NOR2_X1 U11195 ( .A1(n10163), .A2(n10162), .ZN(n10164) );
  XOR2_X1 U11196 ( .A(P2_ADDR_REG_18__SCAN_IN), .B(n10164), .Z(ADD_1068_U55)
         );
  XNOR2_X1 U11197 ( .A(n10166), .B(n10165), .ZN(ADD_1068_U56) );
  XNOR2_X1 U11198 ( .A(n10168), .B(n10167), .ZN(ADD_1068_U57) );
  XNOR2_X1 U11199 ( .A(n10170), .B(n10169), .ZN(ADD_1068_U58) );
  XNOR2_X1 U11200 ( .A(n10172), .B(n10171), .ZN(ADD_1068_U59) );
  XNOR2_X1 U11201 ( .A(n10174), .B(n10173), .ZN(ADD_1068_U60) );
  XNOR2_X1 U11202 ( .A(n10176), .B(n10175), .ZN(ADD_1068_U61) );
  XNOR2_X1 U11203 ( .A(n10178), .B(n10177), .ZN(ADD_1068_U62) );
  XNOR2_X1 U11204 ( .A(n10180), .B(n10179), .ZN(ADD_1068_U63) );
  XNOR2_X1 U11205 ( .A(n10182), .B(n10181), .ZN(ADD_1068_U50) );
  XNOR2_X1 U11206 ( .A(n10184), .B(n10183), .ZN(ADD_1068_U51) );
  XNOR2_X1 U11207 ( .A(n10186), .B(n10185), .ZN(ADD_1068_U47) );
  XNOR2_X1 U11208 ( .A(n10188), .B(n10187), .ZN(ADD_1068_U49) );
  XNOR2_X1 U11209 ( .A(n10190), .B(n10189), .ZN(ADD_1068_U48) );
  XOR2_X1 U11210 ( .A(n10192), .B(n10191), .Z(ADD_1068_U54) );
  XOR2_X1 U11211 ( .A(n10194), .B(n10193), .Z(ADD_1068_U53) );
  XNOR2_X1 U11212 ( .A(n10196), .B(n10195), .ZN(ADD_1068_U52) );
  NAND2_X1 U6145 ( .A1(n5109), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5799) );
  AND4_X1 U6848 ( .A1(n5273), .A2(n5272), .A3(n5271), .A4(n5270), .ZN(n7220)
         );
  CLKBUF_X2 U4890 ( .A(n5948), .Z(n8402) );
  NAND2_X1 U9798 ( .A1(n8187), .A2(n8186), .ZN(n9027) );
endmodule

